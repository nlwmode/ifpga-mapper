module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] , \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] , \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] , \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] , \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] , \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] , \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] , \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] , \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] , \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] , \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] , \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] , \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] , \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] , \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] , \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] , \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] , \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] , \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] , \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] , \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] , \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] , \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] , \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] , \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] , \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] , \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] , \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] , \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] , \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] , \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] , \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127] );
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	input \a[24]  ;
	input \a[25]  ;
	input \a[26]  ;
	input \a[27]  ;
	input \a[28]  ;
	input \a[29]  ;
	input \a[30]  ;
	input \a[31]  ;
	input \a[32]  ;
	input \a[33]  ;
	input \a[34]  ;
	input \a[35]  ;
	input \a[36]  ;
	input \a[37]  ;
	input \a[38]  ;
	input \a[39]  ;
	input \a[40]  ;
	input \a[41]  ;
	input \a[42]  ;
	input \a[43]  ;
	input \a[44]  ;
	input \a[45]  ;
	input \a[46]  ;
	input \a[47]  ;
	input \a[48]  ;
	input \a[49]  ;
	input \a[50]  ;
	input \a[51]  ;
	input \a[52]  ;
	input \a[53]  ;
	input \a[54]  ;
	input \a[55]  ;
	input \a[56]  ;
	input \a[57]  ;
	input \a[58]  ;
	input \a[59]  ;
	input \a[60]  ;
	input \a[61]  ;
	input \a[62]  ;
	input \a[63]  ;
	output \asquared[0]  ;
	output \asquared[1]  ;
	output \asquared[2]  ;
	output \asquared[3]  ;
	output \asquared[4]  ;
	output \asquared[5]  ;
	output \asquared[6]  ;
	output \asquared[7]  ;
	output \asquared[8]  ;
	output \asquared[9]  ;
	output \asquared[10]  ;
	output \asquared[11]  ;
	output \asquared[12]  ;
	output \asquared[13]  ;
	output \asquared[14]  ;
	output \asquared[15]  ;
	output \asquared[16]  ;
	output \asquared[17]  ;
	output \asquared[18]  ;
	output \asquared[19]  ;
	output \asquared[20]  ;
	output \asquared[21]  ;
	output \asquared[22]  ;
	output \asquared[23]  ;
	output \asquared[24]  ;
	output \asquared[25]  ;
	output \asquared[26]  ;
	output \asquared[27]  ;
	output \asquared[28]  ;
	output \asquared[29]  ;
	output \asquared[30]  ;
	output \asquared[31]  ;
	output \asquared[32]  ;
	output \asquared[33]  ;
	output \asquared[34]  ;
	output \asquared[35]  ;
	output \asquared[36]  ;
	output \asquared[37]  ;
	output \asquared[38]  ;
	output \asquared[39]  ;
	output \asquared[40]  ;
	output \asquared[41]  ;
	output \asquared[42]  ;
	output \asquared[43]  ;
	output \asquared[44]  ;
	output \asquared[45]  ;
	output \asquared[46]  ;
	output \asquared[47]  ;
	output \asquared[48]  ;
	output \asquared[49]  ;
	output \asquared[50]  ;
	output \asquared[51]  ;
	output \asquared[52]  ;
	output \asquared[53]  ;
	output \asquared[54]  ;
	output \asquared[55]  ;
	output \asquared[56]  ;
	output \asquared[57]  ;
	output \asquared[58]  ;
	output \asquared[59]  ;
	output \asquared[60]  ;
	output \asquared[61]  ;
	output \asquared[62]  ;
	output \asquared[63]  ;
	output \asquared[64]  ;
	output \asquared[65]  ;
	output \asquared[66]  ;
	output \asquared[67]  ;
	output \asquared[68]  ;
	output \asquared[69]  ;
	output \asquared[70]  ;
	output \asquared[71]  ;
	output \asquared[72]  ;
	output \asquared[73]  ;
	output \asquared[74]  ;
	output \asquared[75]  ;
	output \asquared[76]  ;
	output \asquared[77]  ;
	output \asquared[78]  ;
	output \asquared[79]  ;
	output \asquared[80]  ;
	output \asquared[81]  ;
	output \asquared[82]  ;
	output \asquared[83]  ;
	output \asquared[84]  ;
	output \asquared[85]  ;
	output \asquared[86]  ;
	output \asquared[87]  ;
	output \asquared[88]  ;
	output \asquared[89]  ;
	output \asquared[90]  ;
	output \asquared[91]  ;
	output \asquared[92]  ;
	output \asquared[93]  ;
	output \asquared[94]  ;
	output \asquared[95]  ;
	output \asquared[96]  ;
	output \asquared[97]  ;
	output \asquared[98]  ;
	output \asquared[99]  ;
	output \asquared[100]  ;
	output \asquared[101]  ;
	output \asquared[102]  ;
	output \asquared[103]  ;
	output \asquared[104]  ;
	output \asquared[105]  ;
	output \asquared[106]  ;
	output \asquared[107]  ;
	output \asquared[108]  ;
	output \asquared[109]  ;
	output \asquared[110]  ;
	output \asquared[111]  ;
	output \asquared[112]  ;
	output \asquared[113]  ;
	output \asquared[114]  ;
	output \asquared[115]  ;
	output \asquared[116]  ;
	output \asquared[117]  ;
	output \asquared[118]  ;
	output \asquared[119]  ;
	output \asquared[120]  ;
	output \asquared[121]  ;
	output \asquared[122]  ;
	output \asquared[123]  ;
	output \asquared[124]  ;
	output \asquared[125]  ;
	output \asquared[126]  ;
	output \asquared[127]  ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\a[0] ,
		\a[1] ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\a[1] ,
		\a[2] ,
		_w67_
	);
	LUT3 #(
		.INIT('h28)
	) name2 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w68_
	);
	LUT3 #(
		.INIT('h80)
	) name3 (
		\a[0] ,
		\a[2] ,
		\a[3] ,
		_w69_
	);
	LUT4 #(
		.INIT('h1ab0)
	) name4 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		\a[3] ,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\a[0] ,
		\a[4] ,
		_w71_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6 (
		\a[0] ,
		\a[1] ,
		\a[3] ,
		\a[4] ,
		_w72_
	);
	LUT3 #(
		.INIT('h96)
	) name7 (
		_w67_,
		_w69_,
		_w72_,
		_w73_
	);
	LUT4 #(
		.INIT('h4c00)
	) name8 (
		\a[0] ,
		\a[1] ,
		\a[3] ,
		\a[4] ,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\a[2] ,
		\a[3] ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\a[0] ,
		\a[5] ,
		_w76_
	);
	LUT3 #(
		.INIT('hde)
	) name11 (
		_w74_,
		_w75_,
		_w76_,
		_w77_
	);
	LUT3 #(
		.INIT('hb7)
	) name12 (
		_w74_,
		_w75_,
		_w76_,
		_w78_
	);
	LUT3 #(
		.INIT('h96)
	) name13 (
		_w74_,
		_w75_,
		_w76_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w67_,
		_w72_,
		_w80_
	);
	LUT3 #(
		.INIT('h13)
	) name15 (
		_w67_,
		_w69_,
		_w72_,
		_w81_
	);
	LUT3 #(
		.INIT('he8)
	) name16 (
		_w67_,
		_w69_,
		_w72_,
		_w82_
	);
	LUT2 #(
		.INIT('h6)
	) name17 (
		_w79_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\a[2] ,
		\a[5] ,
		_w84_
	);
	LUT4 #(
		.INIT('h8000)
	) name19 (
		\a[1] ,
		\a[2] ,
		\a[4] ,
		\a[5] ,
		_w85_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name20 (
		\a[1] ,
		\a[2] ,
		\a[4] ,
		\a[5] ,
		_w86_
	);
	LUT4 #(
		.INIT('h153f)
	) name21 (
		\a[0] ,
		\a[2] ,
		\a[3] ,
		\a[6] ,
		_w87_
	);
	LUT4 #(
		.INIT('h8000)
	) name22 (
		\a[0] ,
		\a[2] ,
		\a[3] ,
		\a[6] ,
		_w88_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name23 (
		\a[0] ,
		\a[2] ,
		\a[3] ,
		\a[6] ,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w86_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h6)
	) name25 (
		_w86_,
		_w89_,
		_w91_
	);
	LUT3 #(
		.INIT('h57)
	) name26 (
		\a[1] ,
		\a[3] ,
		\a[5] ,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		_w71_,
		_w92_,
		_w93_
	);
	LUT4 #(
		.INIT('hc341)
	) name28 (
		_w71_,
		_w86_,
		_w89_,
		_w92_,
		_w94_
	);
	LUT4 #(
		.INIT('h0028)
	) name29 (
		_w71_,
		_w86_,
		_w89_,
		_w92_,
		_w95_
	);
	LUT4 #(
		.INIT('h3c96)
	) name30 (
		_w71_,
		_w86_,
		_w89_,
		_w92_,
		_w96_
	);
	LUT4 #(
		.INIT('hccc4)
	) name31 (
		_w77_,
		_w78_,
		_w80_,
		_w81_,
		_w97_
	);
	LUT2 #(
		.INIT('h9)
	) name32 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT3 #(
		.INIT('h0d)
	) name33 (
		_w86_,
		_w87_,
		_w88_,
		_w99_
	);
	LUT3 #(
		.INIT('h9b)
	) name34 (
		\a[1] ,
		\a[4] ,
		\a[6] ,
		_w100_
	);
	LUT4 #(
		.INIT('h004c)
	) name35 (
		\a[2] ,
		\a[4] ,
		\a[5] ,
		\a[6] ,
		_w101_
	);
	LUT4 #(
		.INIT('h8000)
	) name36 (
		\a[1] ,
		\a[2] ,
		\a[5] ,
		\a[6] ,
		_w102_
	);
	LUT3 #(
		.INIT('h02)
	) name37 (
		_w100_,
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\a[0] ,
		\a[7] ,
		_w104_
	);
	LUT4 #(
		.INIT('h153f)
	) name39 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w105_
	);
	LUT4 #(
		.INIT('h8000)
	) name40 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w106_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name41 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w107_
	);
	LUT2 #(
		.INIT('h6)
	) name42 (
		_w104_,
		_w107_,
		_w108_
	);
	LUT3 #(
		.INIT('h09)
	) name43 (
		_w99_,
		_w103_,
		_w108_,
		_w109_
	);
	LUT3 #(
		.INIT('h60)
	) name44 (
		_w99_,
		_w103_,
		_w108_,
		_w110_
	);
	LUT3 #(
		.INIT('h96)
	) name45 (
		_w99_,
		_w103_,
		_w108_,
		_w111_
	);
	LUT4 #(
		.INIT('hba45)
	) name46 (
		_w94_,
		_w95_,
		_w97_,
		_w111_,
		_w112_
	);
	LUT4 #(
		.INIT('h1393)
	) name47 (
		\a[1] ,
		\a[4] ,
		\a[6] ,
		_w84_,
		_w113_
	);
	LUT3 #(
		.INIT('h0b)
	) name48 (
		\a[6] ,
		_w85_,
		_w88_,
		_w114_
	);
	LUT3 #(
		.INIT('h23)
	) name49 (
		_w90_,
		_w113_,
		_w114_,
		_w115_
	);
	LUT4 #(
		.INIT('h8000)
	) name50 (
		\a[1] ,
		\a[3] ,
		\a[5] ,
		\a[7] ,
		_w116_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name51 (
		\a[1] ,
		\a[3] ,
		\a[5] ,
		\a[7] ,
		_w117_
	);
	LUT4 #(
		.INIT('hf200)
	) name52 (
		_w104_,
		_w105_,
		_w106_,
		_w117_,
		_w118_
	);
	LUT4 #(
		.INIT('h000d)
	) name53 (
		_w104_,
		_w105_,
		_w106_,
		_w117_,
		_w119_
	);
	LUT4 #(
		.INIT('h0df2)
	) name54 (
		_w104_,
		_w105_,
		_w106_,
		_w117_,
		_w120_
	);
	LUT3 #(
		.INIT('h80)
	) name55 (
		\a[1] ,
		\a[4] ,
		\a[6] ,
		_w121_
	);
	LUT4 #(
		.INIT('h153f)
	) name56 (
		\a[0] ,
		\a[2] ,
		\a[6] ,
		\a[8] ,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\a[2] ,
		\a[8] ,
		_w123_
	);
	LUT4 #(
		.INIT('h8000)
	) name58 (
		\a[0] ,
		\a[2] ,
		\a[6] ,
		\a[8] ,
		_w124_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name59 (
		\a[0] ,
		\a[2] ,
		\a[6] ,
		\a[8] ,
		_w125_
	);
	LUT2 #(
		.INIT('h6)
	) name60 (
		_w121_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h6)
	) name61 (
		_w120_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w115_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h6)
	) name63 (
		_w115_,
		_w127_,
		_w129_
	);
	LUT4 #(
		.INIT('h0071)
	) name64 (
		_w91_,
		_w93_,
		_w97_,
		_w110_,
		_w130_
	);
	LUT3 #(
		.INIT('hc9)
	) name65 (
		_w109_,
		_w129_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h32)
	) name66 (
		_w118_,
		_w119_,
		_w126_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\a[0] ,
		\a[9] ,
		_w133_
	);
	LUT3 #(
		.INIT('h93)
	) name68 (
		\a[1] ,
		\a[5] ,
		\a[8] ,
		_w134_
	);
	LUT3 #(
		.INIT('h69)
	) name69 (
		_w116_,
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\a[2] ,
		\a[7] ,
		_w136_
	);
	LUT4 #(
		.INIT('h153f)
	) name71 (
		\a[3] ,
		\a[4] ,
		\a[5] ,
		\a[6] ,
		_w137_
	);
	LUT4 #(
		.INIT('h8000)
	) name72 (
		\a[3] ,
		\a[4] ,
		\a[5] ,
		\a[6] ,
		_w138_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name73 (
		\a[3] ,
		\a[4] ,
		\a[5] ,
		\a[6] ,
		_w139_
	);
	LUT2 #(
		.INIT('h6)
	) name74 (
		_w136_,
		_w139_,
		_w140_
	);
	LUT3 #(
		.INIT('h0d)
	) name75 (
		_w121_,
		_w122_,
		_w124_,
		_w141_
	);
	LUT3 #(
		.INIT('h69)
	) name76 (
		_w135_,
		_w140_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h6)
	) name77 (
		_w132_,
		_w142_,
		_w143_
	);
	LUT3 #(
		.INIT('h54)
	) name78 (
		_w109_,
		_w115_,
		_w127_,
		_w144_
	);
	LUT4 #(
		.INIT('h4b5a)
	) name79 (
		_w128_,
		_w130_,
		_w143_,
		_w144_,
		_w145_
	);
	LUT4 #(
		.INIT('h0777)
	) name80 (
		_w115_,
		_w127_,
		_w132_,
		_w142_,
		_w146_
	);
	LUT3 #(
		.INIT('h8e)
	) name81 (
		_w135_,
		_w140_,
		_w141_,
		_w147_
	);
	LUT3 #(
		.INIT('h80)
	) name82 (
		\a[1] ,
		\a[5] ,
		\a[8] ,
		_w148_
	);
	LUT4 #(
		.INIT('h8000)
	) name83 (
		\a[1] ,
		\a[4] ,
		\a[6] ,
		\a[9] ,
		_w149_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name84 (
		\a[1] ,
		\a[4] ,
		\a[6] ,
		\a[9] ,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w148_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w148_,
		_w150_,
		_w152_
	);
	LUT2 #(
		.INIT('h6)
	) name87 (
		_w148_,
		_w150_,
		_w153_
	);
	LUT3 #(
		.INIT('h0d)
	) name88 (
		_w136_,
		_w137_,
		_w138_,
		_w154_
	);
	LUT3 #(
		.INIT('h8e)
	) name89 (
		_w116_,
		_w133_,
		_w134_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\a[3] ,
		\a[7] ,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\a[0] ,
		\a[10] ,
		_w157_
	);
	LUT4 #(
		.INIT('h153f)
	) name92 (
		\a[0] ,
		\a[3] ,
		\a[7] ,
		\a[10] ,
		_w158_
	);
	LUT4 #(
		.INIT('h8000)
	) name93 (
		\a[0] ,
		\a[3] ,
		\a[7] ,
		\a[10] ,
		_w159_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name94 (
		\a[0] ,
		\a[3] ,
		\a[7] ,
		\a[10] ,
		_w160_
	);
	LUT2 #(
		.INIT('h6)
	) name95 (
		_w123_,
		_w160_,
		_w161_
	);
	LUT4 #(
		.INIT('h9669)
	) name96 (
		_w153_,
		_w154_,
		_w155_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w147_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w147_,
		_w162_,
		_w164_
	);
	LUT2 #(
		.INIT('h6)
	) name99 (
		_w147_,
		_w162_,
		_w165_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name100 (
		_w132_,
		_w142_,
		_w147_,
		_w162_,
		_w166_
	);
	LUT4 #(
		.INIT('h4f00)
	) name101 (
		_w130_,
		_w144_,
		_w146_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('h1001)
	) name102 (
		_w132_,
		_w142_,
		_w147_,
		_w162_,
		_w168_
	);
	LUT4 #(
		.INIT('h00b0)
	) name103 (
		_w130_,
		_w144_,
		_w146_,
		_w165_,
		_w169_
	);
	LUT3 #(
		.INIT('h01)
	) name104 (
		_w167_,
		_w168_,
		_w169_,
		_w170_
	);
	LUT4 #(
		.INIT('h0111)
	) name105 (
		_w132_,
		_w142_,
		_w147_,
		_w162_,
		_w171_
	);
	LUT4 #(
		.INIT('h00b0)
	) name106 (
		_w130_,
		_w144_,
		_w146_,
		_w164_,
		_w172_
	);
	LUT4 #(
		.INIT('h066f)
	) name107 (
		_w153_,
		_w154_,
		_w155_,
		_w161_,
		_w173_
	);
	LUT3 #(
		.INIT('h93)
	) name108 (
		\a[1] ,
		\a[6] ,
		\a[10] ,
		_w174_
	);
	LUT3 #(
		.INIT('h32)
	) name109 (
		_w123_,
		_w158_,
		_w159_,
		_w175_
	);
	LUT4 #(
		.INIT('h00e8)
	) name110 (
		_w123_,
		_w156_,
		_w157_,
		_w174_,
		_w176_
	);
	LUT4 #(
		.INIT('h1700)
	) name111 (
		_w123_,
		_w156_,
		_w157_,
		_w174_,
		_w177_
	);
	LUT4 #(
		.INIT('h32cd)
	) name112 (
		_w123_,
		_w158_,
		_w159_,
		_w174_,
		_w178_
	);
	LUT4 #(
		.INIT('h153f)
	) name113 (
		\a[2] ,
		\a[3] ,
		\a[8] ,
		\a[9] ,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\a[3] ,
		\a[9] ,
		_w180_
	);
	LUT4 #(
		.INIT('h8000)
	) name115 (
		\a[2] ,
		\a[3] ,
		\a[8] ,
		\a[9] ,
		_w181_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name116 (
		\a[2] ,
		\a[3] ,
		\a[8] ,
		\a[9] ,
		_w182_
	);
	LUT2 #(
		.INIT('h6)
	) name117 (
		_w149_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h6)
	) name118 (
		_w178_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\a[0] ,
		\a[11] ,
		_w185_
	);
	LUT4 #(
		.INIT('h153f)
	) name120 (
		\a[4] ,
		\a[5] ,
		\a[6] ,
		\a[7] ,
		_w186_
	);
	LUT4 #(
		.INIT('h8000)
	) name121 (
		\a[4] ,
		\a[5] ,
		\a[6] ,
		\a[7] ,
		_w187_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name122 (
		\a[4] ,
		\a[5] ,
		\a[6] ,
		\a[7] ,
		_w188_
	);
	LUT2 #(
		.INIT('h6)
	) name123 (
		_w185_,
		_w188_,
		_w189_
	);
	LUT4 #(
		.INIT('h8e00)
	) name124 (
		_w148_,
		_w150_,
		_w154_,
		_w189_,
		_w190_
	);
	LUT4 #(
		.INIT('h0071)
	) name125 (
		_w148_,
		_w150_,
		_w154_,
		_w189_,
		_w191_
	);
	LUT4 #(
		.INIT('hdc23)
	) name126 (
		_w151_,
		_w152_,
		_w154_,
		_w189_,
		_w192_
	);
	LUT3 #(
		.INIT('h82)
	) name127 (
		_w173_,
		_w184_,
		_w192_,
		_w193_
	);
	LUT3 #(
		.INIT('h14)
	) name128 (
		_w173_,
		_w184_,
		_w192_,
		_w194_
	);
	LUT3 #(
		.INIT('h69)
	) name129 (
		_w173_,
		_w184_,
		_w192_,
		_w195_
	);
	LUT4 #(
		.INIT('hfee0)
	) name130 (
		_w132_,
		_w142_,
		_w147_,
		_w162_,
		_w196_
	);
	LUT4 #(
		.INIT('hfe01)
	) name131 (
		_w163_,
		_w171_,
		_w172_,
		_w195_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w193_,
		_w196_,
		_w198_
	);
	LUT3 #(
		.INIT('h31)
	) name133 (
		_w184_,
		_w190_,
		_w191_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\a[5] ,
		\a[11] ,
		_w200_
	);
	LUT4 #(
		.INIT('h8000)
	) name135 (
		\a[1] ,
		\a[5] ,
		\a[7] ,
		\a[11] ,
		_w201_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name136 (
		\a[1] ,
		\a[5] ,
		\a[7] ,
		\a[11] ,
		_w202_
	);
	LUT3 #(
		.INIT('h80)
	) name137 (
		\a[1] ,
		\a[6] ,
		\a[10] ,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\a[4] ,
		\a[8] ,
		_w204_
	);
	LUT3 #(
		.INIT('h96)
	) name139 (
		_w202_,
		_w203_,
		_w204_,
		_w205_
	);
	LUT4 #(
		.INIT('hd400)
	) name140 (
		_w174_,
		_w175_,
		_w183_,
		_w205_,
		_w206_
	);
	LUT4 #(
		.INIT('h002b)
	) name141 (
		_w174_,
		_w175_,
		_w183_,
		_w205_,
		_w207_
	);
	LUT4 #(
		.INIT('hcd32)
	) name142 (
		_w176_,
		_w177_,
		_w183_,
		_w205_,
		_w208_
	);
	LUT3 #(
		.INIT('h0d)
	) name143 (
		_w149_,
		_w179_,
		_w181_,
		_w209_
	);
	LUT3 #(
		.INIT('h0d)
	) name144 (
		_w185_,
		_w186_,
		_w187_,
		_w210_
	);
	LUT4 #(
		.INIT('h153f)
	) name145 (
		\a[0] ,
		\a[2] ,
		\a[10] ,
		\a[12] ,
		_w211_
	);
	LUT4 #(
		.INIT('h8000)
	) name146 (
		\a[0] ,
		\a[2] ,
		\a[10] ,
		\a[12] ,
		_w212_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name147 (
		\a[0] ,
		\a[2] ,
		\a[10] ,
		\a[12] ,
		_w213_
	);
	LUT2 #(
		.INIT('h6)
	) name148 (
		_w180_,
		_w213_,
		_w214_
	);
	LUT3 #(
		.INIT('h69)
	) name149 (
		_w209_,
		_w210_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h9)
	) name150 (
		_w208_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		_w199_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h9)
	) name152 (
		_w199_,
		_w216_,
		_w218_
	);
	LUT4 #(
		.INIT('h23dc)
	) name153 (
		_w172_,
		_w194_,
		_w198_,
		_w218_,
		_w219_
	);
	LUT3 #(
		.INIT('h45)
	) name154 (
		_w194_,
		_w199_,
		_w216_,
		_w220_
	);
	LUT3 #(
		.INIT('hb0)
	) name155 (
		_w172_,
		_w198_,
		_w220_,
		_w221_
	);
	LUT3 #(
		.INIT('h23)
	) name156 (
		_w206_,
		_w207_,
		_w215_,
		_w222_
	);
	LUT3 #(
		.INIT('he8)
	) name157 (
		_w202_,
		_w203_,
		_w204_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		\a[3] ,
		\a[10] ,
		_w224_
	);
	LUT4 #(
		.INIT('h153f)
	) name159 (
		\a[0] ,
		\a[4] ,
		\a[9] ,
		\a[13] ,
		_w225_
	);
	LUT4 #(
		.INIT('h8000)
	) name160 (
		\a[0] ,
		\a[4] ,
		\a[9] ,
		\a[13] ,
		_w226_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name161 (
		\a[0] ,
		\a[4] ,
		\a[9] ,
		\a[13] ,
		_w227_
	);
	LUT2 #(
		.INIT('h6)
	) name162 (
		_w224_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\a[2] ,
		\a[11] ,
		_w229_
	);
	LUT4 #(
		.INIT('h153f)
	) name164 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w230_
	);
	LUT4 #(
		.INIT('h8000)
	) name165 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w231_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name166 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w232_
	);
	LUT2 #(
		.INIT('h6)
	) name167 (
		_w229_,
		_w232_,
		_w233_
	);
	LUT3 #(
		.INIT('h96)
	) name168 (
		_w223_,
		_w228_,
		_w233_,
		_w234_
	);
	LUT3 #(
		.INIT('h9b)
	) name169 (
		\a[1] ,
		\a[7] ,
		\a[12] ,
		_w235_
	);
	LUT4 #(
		.INIT('h004c)
	) name170 (
		\a[5] ,
		\a[7] ,
		\a[11] ,
		\a[12] ,
		_w236_
	);
	LUT4 #(
		.INIT('h8000)
	) name171 (
		\a[1] ,
		\a[5] ,
		\a[11] ,
		\a[12] ,
		_w237_
	);
	LUT3 #(
		.INIT('h02)
	) name172 (
		_w235_,
		_w236_,
		_w237_,
		_w238_
	);
	LUT3 #(
		.INIT('h0d)
	) name173 (
		_w180_,
		_w211_,
		_w212_,
		_w239_
	);
	LUT2 #(
		.INIT('h6)
	) name174 (
		_w238_,
		_w239_,
		_w240_
	);
	LUT3 #(
		.INIT('h8e)
	) name175 (
		_w209_,
		_w210_,
		_w214_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		_w240_,
		_w241_,
		_w243_
	);
	LUT2 #(
		.INIT('h9)
	) name178 (
		_w240_,
		_w241_,
		_w244_
	);
	LUT3 #(
		.INIT('hde)
	) name179 (
		_w222_,
		_w234_,
		_w244_,
		_w245_
	);
	LUT3 #(
		.INIT('hb7)
	) name180 (
		_w222_,
		_w234_,
		_w244_,
		_w246_
	);
	LUT3 #(
		.INIT('h96)
	) name181 (
		_w222_,
		_w234_,
		_w244_,
		_w247_
	);
	LUT4 #(
		.INIT('h00b0)
	) name182 (
		_w172_,
		_w198_,
		_w220_,
		_w247_,
		_w248_
	);
	LUT4 #(
		.INIT('h00e5)
	) name183 (
		_w217_,
		_w221_,
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w217_,
		_w246_,
		_w250_
	);
	LUT4 #(
		.INIT('hb000)
	) name185 (
		_w172_,
		_w198_,
		_w220_,
		_w246_,
		_w251_
	);
	LUT3 #(
		.INIT('he8)
	) name186 (
		_w223_,
		_w228_,
		_w233_,
		_w252_
	);
	LUT4 #(
		.INIT('h8000)
	) name187 (
		\a[1] ,
		\a[6] ,
		\a[8] ,
		\a[13] ,
		_w253_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name188 (
		\a[1] ,
		\a[6] ,
		\a[8] ,
		\a[13] ,
		_w254_
	);
	LUT4 #(
		.INIT('hf200)
	) name189 (
		_w229_,
		_w230_,
		_w231_,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('h000d)
	) name190 (
		_w229_,
		_w230_,
		_w231_,
		_w254_,
		_w256_
	);
	LUT4 #(
		.INIT('h0df2)
	) name191 (
		_w229_,
		_w230_,
		_w231_,
		_w254_,
		_w257_
	);
	LUT3 #(
		.INIT('h0d)
	) name192 (
		_w224_,
		_w225_,
		_w226_,
		_w258_
	);
	LUT2 #(
		.INIT('h6)
	) name193 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		\a[12] ,
		_w201_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\a[0] ,
		\a[14] ,
		_w261_
	);
	LUT4 #(
		.INIT('h153f)
	) name196 (
		\a[2] ,
		\a[3] ,
		\a[11] ,
		\a[12] ,
		_w262_
	);
	LUT4 #(
		.INIT('h8000)
	) name197 (
		\a[2] ,
		\a[3] ,
		\a[11] ,
		\a[12] ,
		_w263_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name198 (
		\a[2] ,
		\a[3] ,
		\a[11] ,
		\a[12] ,
		_w264_
	);
	LUT3 #(
		.INIT('h80)
	) name199 (
		\a[1] ,
		\a[7] ,
		\a[12] ,
		_w265_
	);
	LUT4 #(
		.INIT('h153f)
	) name200 (
		\a[4] ,
		\a[5] ,
		\a[9] ,
		\a[10] ,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\a[5] ,
		\a[10] ,
		_w267_
	);
	LUT4 #(
		.INIT('h8000)
	) name202 (
		\a[4] ,
		\a[5] ,
		\a[9] ,
		\a[10] ,
		_w268_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name203 (
		\a[4] ,
		\a[5] ,
		\a[9] ,
		\a[10] ,
		_w269_
	);
	LUT4 #(
		.INIT('h0660)
	) name204 (
		_w261_,
		_w264_,
		_w265_,
		_w269_,
		_w270_
	);
	LUT4 #(
		.INIT('h9009)
	) name205 (
		_w261_,
		_w264_,
		_w265_,
		_w269_,
		_w271_
	);
	LUT4 #(
		.INIT('h6996)
	) name206 (
		_w261_,
		_w264_,
		_w265_,
		_w269_,
		_w272_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name207 (
		_w238_,
		_w239_,
		_w260_,
		_w272_,
		_w273_
	);
	LUT3 #(
		.INIT('h69)
	) name208 (
		_w252_,
		_w259_,
		_w273_,
		_w274_
	);
	LUT4 #(
		.INIT('h8e00)
	) name209 (
		_w222_,
		_w240_,
		_w241_,
		_w274_,
		_w275_
	);
	LUT4 #(
		.INIT('h0071)
	) name210 (
		_w222_,
		_w240_,
		_w241_,
		_w274_,
		_w276_
	);
	LUT4 #(
		.INIT('h0df2)
	) name211 (
		_w222_,
		_w242_,
		_w243_,
		_w274_,
		_w277_
	);
	LUT4 #(
		.INIT('hfd02)
	) name212 (
		_w245_,
		_w250_,
		_w251_,
		_w277_,
		_w278_
	);
	LUT4 #(
		.INIT('h004c)
	) name213 (
		_w217_,
		_w245_,
		_w246_,
		_w276_,
		_w279_
	);
	LUT3 #(
		.INIT('hb2)
	) name214 (
		_w252_,
		_w259_,
		_w273_,
		_w280_
	);
	LUT3 #(
		.INIT('h23)
	) name215 (
		_w255_,
		_w256_,
		_w258_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		\a[4] ,
		\a[11] ,
		_w282_
	);
	LUT3 #(
		.INIT('h80)
	) name217 (
		\a[1] ,
		\a[8] ,
		\a[14] ,
		_w283_
	);
	LUT3 #(
		.INIT('h6c)
	) name218 (
		\a[1] ,
		\a[8] ,
		\a[14] ,
		_w284_
	);
	LUT3 #(
		.INIT('h96)
	) name219 (
		_w253_,
		_w282_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\a[2] ,
		\a[13] ,
		_w286_
	);
	LUT4 #(
		.INIT('h153f)
	) name221 (
		\a[6] ,
		\a[7] ,
		\a[8] ,
		\a[9] ,
		_w287_
	);
	LUT4 #(
		.INIT('h8000)
	) name222 (
		\a[6] ,
		\a[7] ,
		\a[8] ,
		\a[9] ,
		_w288_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name223 (
		\a[6] ,
		\a[7] ,
		\a[8] ,
		\a[9] ,
		_w289_
	);
	LUT2 #(
		.INIT('h6)
	) name224 (
		_w286_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		_w285_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		_w285_,
		_w290_,
		_w292_
	);
	LUT2 #(
		.INIT('h6)
	) name227 (
		_w285_,
		_w290_,
		_w293_
	);
	LUT2 #(
		.INIT('h6)
	) name228 (
		_w281_,
		_w293_,
		_w294_
	);
	LUT4 #(
		.INIT('h000e)
	) name229 (
		_w238_,
		_w239_,
		_w260_,
		_w270_,
		_w295_
	);
	LUT3 #(
		.INIT('h0d)
	) name230 (
		_w265_,
		_w266_,
		_w268_,
		_w296_
	);
	LUT3 #(
		.INIT('h0d)
	) name231 (
		_w261_,
		_w262_,
		_w263_,
		_w297_
	);
	LUT4 #(
		.INIT('h153f)
	) name232 (
		\a[0] ,
		\a[3] ,
		\a[12] ,
		\a[15] ,
		_w298_
	);
	LUT4 #(
		.INIT('h8000)
	) name233 (
		\a[0] ,
		\a[3] ,
		\a[12] ,
		\a[15] ,
		_w299_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name234 (
		\a[0] ,
		\a[3] ,
		\a[12] ,
		\a[15] ,
		_w300_
	);
	LUT2 #(
		.INIT('h6)
	) name235 (
		_w267_,
		_w300_,
		_w301_
	);
	LUT3 #(
		.INIT('h69)
	) name236 (
		_w296_,
		_w297_,
		_w301_,
		_w302_
	);
	LUT3 #(
		.INIT('he0)
	) name237 (
		_w271_,
		_w295_,
		_w302_,
		_w303_
	);
	LUT3 #(
		.INIT('h01)
	) name238 (
		_w271_,
		_w295_,
		_w302_,
		_w304_
	);
	LUT3 #(
		.INIT('h1e)
	) name239 (
		_w271_,
		_w295_,
		_w302_,
		_w305_
	);
	LUT3 #(
		.INIT('h28)
	) name240 (
		_w280_,
		_w294_,
		_w305_,
		_w306_
	);
	LUT3 #(
		.INIT('h41)
	) name241 (
		_w280_,
		_w294_,
		_w305_,
		_w307_
	);
	LUT3 #(
		.INIT('h96)
	) name242 (
		_w280_,
		_w294_,
		_w305_,
		_w308_
	);
	LUT4 #(
		.INIT('h23dc)
	) name243 (
		_w251_,
		_w275_,
		_w279_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w275_,
		_w306_,
		_w310_
	);
	LUT3 #(
		.INIT('h0d)
	) name245 (
		_w294_,
		_w303_,
		_w304_,
		_w311_
	);
	LUT3 #(
		.INIT('he8)
	) name246 (
		_w253_,
		_w282_,
		_w284_,
		_w312_
	);
	LUT3 #(
		.INIT('h32)
	) name247 (
		_w267_,
		_w298_,
		_w299_,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w312_,
		_w313_,
		_w314_
	);
	LUT4 #(
		.INIT('h153f)
	) name249 (
		\a[0] ,
		\a[6] ,
		\a[10] ,
		\a[16] ,
		_w315_
	);
	LUT4 #(
		.INIT('h8000)
	) name250 (
		\a[0] ,
		\a[6] ,
		\a[10] ,
		\a[16] ,
		_w316_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name251 (
		\a[0] ,
		\a[6] ,
		\a[10] ,
		\a[16] ,
		_w317_
	);
	LUT2 #(
		.INIT('h6)
	) name252 (
		_w200_,
		_w317_,
		_w318_
	);
	LUT3 #(
		.INIT('h69)
	) name253 (
		_w312_,
		_w313_,
		_w318_,
		_w319_
	);
	LUT4 #(
		.INIT('h1700)
	) name254 (
		_w281_,
		_w285_,
		_w290_,
		_w319_,
		_w320_
	);
	LUT4 #(
		.INIT('h00e8)
	) name255 (
		_w281_,
		_w285_,
		_w290_,
		_w319_,
		_w321_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name256 (
		_w281_,
		_w291_,
		_w292_,
		_w319_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\a[4] ,
		\a[12] ,
		_w323_
	);
	LUT4 #(
		.INIT('h153f)
	) name258 (
		\a[2] ,
		\a[3] ,
		\a[13] ,
		\a[14] ,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\a[3] ,
		\a[14] ,
		_w325_
	);
	LUT4 #(
		.INIT('h8000)
	) name260 (
		\a[2] ,
		\a[3] ,
		\a[13] ,
		\a[14] ,
		_w326_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name261 (
		\a[2] ,
		\a[3] ,
		\a[13] ,
		\a[14] ,
		_w327_
	);
	LUT2 #(
		.INIT('h6)
	) name262 (
		_w323_,
		_w327_,
		_w328_
	);
	LUT4 #(
		.INIT('h7100)
	) name263 (
		_w296_,
		_w297_,
		_w301_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('h8000)
	) name264 (
		\a[1] ,
		\a[7] ,
		\a[9] ,
		\a[15] ,
		_w330_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name265 (
		\a[1] ,
		\a[7] ,
		\a[9] ,
		\a[15] ,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w283_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w283_,
		_w331_,
		_w333_
	);
	LUT2 #(
		.INIT('h6)
	) name268 (
		_w283_,
		_w331_,
		_w334_
	);
	LUT3 #(
		.INIT('h32)
	) name269 (
		_w286_,
		_w287_,
		_w288_,
		_w335_
	);
	LUT2 #(
		.INIT('h6)
	) name270 (
		_w334_,
		_w335_,
		_w336_
	);
	LUT4 #(
		.INIT('h008e)
	) name271 (
		_w296_,
		_w297_,
		_w301_,
		_w328_,
		_w337_
	);
	LUT3 #(
		.INIT('hc9)
	) name272 (
		_w329_,
		_w336_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h6)
	) name273 (
		_w322_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		_w311_,
		_w339_,
		_w340_
	);
	LUT3 #(
		.INIT('h96)
	) name275 (
		_w307_,
		_w311_,
		_w339_,
		_w341_
	);
	LUT4 #(
		.INIT('h4f00)
	) name276 (
		_w251_,
		_w279_,
		_w310_,
		_w341_,
		_w342_
	);
	LUT3 #(
		.INIT('hc3)
	) name277 (
		_w307_,
		_w311_,
		_w339_,
		_w343_
	);
	LUT4 #(
		.INIT('hb000)
	) name278 (
		_w251_,
		_w279_,
		_w310_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('he)
	) name279 (
		_w342_,
		_w344_,
		_w345_
	);
	LUT3 #(
		.INIT('h8a)
	) name280 (
		_w307_,
		_w311_,
		_w339_,
		_w346_
	);
	LUT4 #(
		.INIT('h1011)
	) name281 (
		_w275_,
		_w306_,
		_w311_,
		_w339_,
		_w347_
	);
	LUT3 #(
		.INIT('hb0)
	) name282 (
		_w251_,
		_w279_,
		_w347_,
		_w348_
	);
	LUT4 #(
		.INIT('h040f)
	) name283 (
		_w251_,
		_w279_,
		_w346_,
		_w347_,
		_w349_
	);
	LUT3 #(
		.INIT('h23)
	) name284 (
		_w320_,
		_w321_,
		_w338_,
		_w350_
	);
	LUT4 #(
		.INIT('h153f)
	) name285 (
		\a[0] ,
		\a[5] ,
		\a[12] ,
		\a[17] ,
		_w351_
	);
	LUT4 #(
		.INIT('h8000)
	) name286 (
		\a[0] ,
		\a[5] ,
		\a[12] ,
		\a[17] ,
		_w352_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name287 (
		\a[0] ,
		\a[5] ,
		\a[12] ,
		\a[17] ,
		_w353_
	);
	LUT4 #(
		.INIT('h153f)
	) name288 (
		\a[7] ,
		\a[8] ,
		\a[9] ,
		\a[10] ,
		_w354_
	);
	LUT4 #(
		.INIT('h8000)
	) name289 (
		\a[7] ,
		\a[8] ,
		\a[9] ,
		\a[10] ,
		_w355_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name290 (
		\a[7] ,
		\a[8] ,
		\a[9] ,
		\a[10] ,
		_w356_
	);
	LUT4 #(
		.INIT('h1428)
	) name291 (
		_w325_,
		_w330_,
		_w353_,
		_w356_,
		_w357_
	);
	LUT4 #(
		.INIT('h8241)
	) name292 (
		_w325_,
		_w330_,
		_w353_,
		_w356_,
		_w358_
	);
	LUT4 #(
		.INIT('h6996)
	) name293 (
		_w325_,
		_w330_,
		_w353_,
		_w356_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\a[6] ,
		\a[11] ,
		_w360_
	);
	LUT4 #(
		.INIT('h153f)
	) name295 (
		\a[2] ,
		\a[4] ,
		\a[13] ,
		\a[15] ,
		_w361_
	);
	LUT4 #(
		.INIT('h8000)
	) name296 (
		\a[2] ,
		\a[4] ,
		\a[13] ,
		\a[15] ,
		_w362_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name297 (
		\a[2] ,
		\a[4] ,
		\a[13] ,
		\a[15] ,
		_w363_
	);
	LUT2 #(
		.INIT('h6)
	) name298 (
		_w360_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h6)
	) name299 (
		_w359_,
		_w364_,
		_w365_
	);
	LUT4 #(
		.INIT('h0051)
	) name300 (
		_w329_,
		_w336_,
		_w337_,
		_w365_,
		_w366_
	);
	LUT4 #(
		.INIT('hae00)
	) name301 (
		_w329_,
		_w336_,
		_w337_,
		_w365_,
		_w367_
	);
	LUT4 #(
		.INIT('h51ae)
	) name302 (
		_w329_,
		_w336_,
		_w337_,
		_w365_,
		_w368_
	);
	LUT3 #(
		.INIT('he0)
	) name303 (
		_w312_,
		_w313_,
		_w318_,
		_w369_
	);
	LUT3 #(
		.INIT('h32)
	) name304 (
		_w332_,
		_w333_,
		_w335_,
		_w370_
	);
	LUT3 #(
		.INIT('h17)
	) name305 (
		_w312_,
		_w313_,
		_w318_,
		_w371_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		_w370_,
		_w371_,
		_w372_
	);
	LUT3 #(
		.INIT('h80)
	) name307 (
		\a[1] ,
		\a[9] ,
		\a[16] ,
		_w373_
	);
	LUT3 #(
		.INIT('h6c)
	) name308 (
		\a[1] ,
		\a[9] ,
		\a[16] ,
		_w374_
	);
	LUT4 #(
		.INIT('hf200)
	) name309 (
		_w323_,
		_w324_,
		_w326_,
		_w374_,
		_w375_
	);
	LUT4 #(
		.INIT('h000d)
	) name310 (
		_w323_,
		_w324_,
		_w326_,
		_w374_,
		_w376_
	);
	LUT4 #(
		.INIT('h0df2)
	) name311 (
		_w323_,
		_w324_,
		_w326_,
		_w374_,
		_w377_
	);
	LUT3 #(
		.INIT('h0d)
	) name312 (
		_w200_,
		_w315_,
		_w316_,
		_w378_
	);
	LUT2 #(
		.INIT('h6)
	) name313 (
		_w377_,
		_w378_,
		_w379_
	);
	LUT4 #(
		.INIT('h00fe)
	) name314 (
		_w314_,
		_w369_,
		_w370_,
		_w379_,
		_w380_
	);
	LUT4 #(
		.INIT('h001e)
	) name315 (
		_w314_,
		_w369_,
		_w370_,
		_w379_,
		_w381_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name316 (
		_w314_,
		_w369_,
		_w370_,
		_w379_,
		_w382_
	);
	LUT2 #(
		.INIT('h6)
	) name317 (
		_w368_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w350_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		_w350_,
		_w383_,
		_w385_
	);
	LUT2 #(
		.INIT('h9)
	) name320 (
		_w350_,
		_w383_,
		_w386_
	);
	LUT3 #(
		.INIT('h71)
	) name321 (
		_w307_,
		_w311_,
		_w339_,
		_w387_
	);
	LUT4 #(
		.INIT('h4f00)
	) name322 (
		_w251_,
		_w279_,
		_w347_,
		_w387_,
		_w388_
	);
	LUT4 #(
		.INIT('hbfb0)
	) name323 (
		_w340_,
		_w349_,
		_w386_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		_w385_,
		_w387_,
		_w390_
	);
	LUT3 #(
		.INIT('h23)
	) name325 (
		_w366_,
		_w367_,
		_w382_,
		_w391_
	);
	LUT3 #(
		.INIT('h32)
	) name326 (
		_w330_,
		_w351_,
		_w352_,
		_w392_
	);
	LUT3 #(
		.INIT('h0d)
	) name327 (
		_w325_,
		_w354_,
		_w355_,
		_w393_
	);
	LUT3 #(
		.INIT('h0d)
	) name328 (
		_w360_,
		_w361_,
		_w362_,
		_w394_
	);
	LUT3 #(
		.INIT('h96)
	) name329 (
		_w392_,
		_w393_,
		_w394_,
		_w395_
	);
	LUT3 #(
		.INIT('h23)
	) name330 (
		_w375_,
		_w376_,
		_w378_,
		_w396_
	);
	LUT3 #(
		.INIT('h32)
	) name331 (
		_w357_,
		_w358_,
		_w364_,
		_w397_
	);
	LUT3 #(
		.INIT('h96)
	) name332 (
		_w395_,
		_w396_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		\a[6] ,
		\a[12] ,
		_w399_
	);
	LUT4 #(
		.INIT('h8000)
	) name334 (
		\a[1] ,
		\a[8] ,
		\a[10] ,
		\a[17] ,
		_w400_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name335 (
		\a[1] ,
		\a[8] ,
		\a[10] ,
		\a[17] ,
		_w401_
	);
	LUT3 #(
		.INIT('h96)
	) name336 (
		_w373_,
		_w399_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\a[4] ,
		\a[14] ,
		_w403_
	);
	LUT4 #(
		.INIT('h153f)
	) name338 (
		\a[2] ,
		\a[3] ,
		\a[15] ,
		\a[16] ,
		_w404_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\a[3] ,
		\a[16] ,
		_w405_
	);
	LUT4 #(
		.INIT('h8000)
	) name340 (
		\a[2] ,
		\a[3] ,
		\a[15] ,
		\a[16] ,
		_w406_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name341 (
		\a[2] ,
		\a[3] ,
		\a[15] ,
		\a[16] ,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		\a[7] ,
		\a[11] ,
		_w408_
	);
	LUT4 #(
		.INIT('h153f)
	) name343 (
		\a[0] ,
		\a[5] ,
		\a[13] ,
		\a[18] ,
		_w409_
	);
	LUT4 #(
		.INIT('h8000)
	) name344 (
		\a[0] ,
		\a[5] ,
		\a[13] ,
		\a[18] ,
		_w410_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name345 (
		\a[0] ,
		\a[5] ,
		\a[13] ,
		\a[18] ,
		_w411_
	);
	LUT4 #(
		.INIT('h0660)
	) name346 (
		_w403_,
		_w407_,
		_w408_,
		_w411_,
		_w412_
	);
	LUT4 #(
		.INIT('h9009)
	) name347 (
		_w403_,
		_w407_,
		_w408_,
		_w411_,
		_w413_
	);
	LUT4 #(
		.INIT('h6996)
	) name348 (
		_w403_,
		_w407_,
		_w408_,
		_w411_,
		_w414_
	);
	LUT2 #(
		.INIT('h6)
	) name349 (
		_w402_,
		_w414_,
		_w415_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name350 (
		_w372_,
		_w381_,
		_w398_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h6)
	) name351 (
		_w391_,
		_w416_,
		_w417_
	);
	LUT4 #(
		.INIT('h23dc)
	) name352 (
		_w348_,
		_w384_,
		_w390_,
		_w417_,
		_w418_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name353 (
		_w350_,
		_w383_,
		_w391_,
		_w416_,
		_w419_
	);
	LUT3 #(
		.INIT('h0e)
	) name354 (
		_w402_,
		_w412_,
		_w413_,
		_w420_
	);
	LUT3 #(
		.INIT('h80)
	) name355 (
		\a[1] ,
		\a[10] ,
		\a[18] ,
		_w421_
	);
	LUT3 #(
		.INIT('h6c)
	) name356 (
		\a[1] ,
		\a[10] ,
		\a[18] ,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w400_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		\a[18] ,
		_w400_,
		_w424_
	);
	LUT3 #(
		.INIT('hb8)
	) name359 (
		\a[18] ,
		_w400_,
		_w422_,
		_w425_
	);
	LUT3 #(
		.INIT('h0d)
	) name360 (
		_w403_,
		_w404_,
		_w406_,
		_w426_
	);
	LUT2 #(
		.INIT('h6)
	) name361 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT3 #(
		.INIT('he8)
	) name362 (
		_w373_,
		_w399_,
		_w401_,
		_w428_
	);
	LUT3 #(
		.INIT('h32)
	) name363 (
		_w408_,
		_w409_,
		_w410_,
		_w429_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\a[9] ,
		\a[10] ,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\a[8] ,
		\a[11] ,
		_w431_
	);
	LUT4 #(
		.INIT('h153f)
	) name366 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w432_
	);
	LUT4 #(
		.INIT('h8000)
	) name367 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w433_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name368 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w434_
	);
	LUT2 #(
		.INIT('h6)
	) name369 (
		_w405_,
		_w434_,
		_w435_
	);
	LUT3 #(
		.INIT('h96)
	) name370 (
		_w428_,
		_w429_,
		_w435_,
		_w436_
	);
	LUT3 #(
		.INIT('h69)
	) name371 (
		_w420_,
		_w427_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		\a[5] ,
		\a[14] ,
		_w438_
	);
	LUT4 #(
		.INIT('h153f)
	) name373 (
		\a[6] ,
		\a[7] ,
		\a[12] ,
		\a[13] ,
		_w439_
	);
	LUT4 #(
		.INIT('h8000)
	) name374 (
		\a[6] ,
		\a[7] ,
		\a[12] ,
		\a[13] ,
		_w440_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name375 (
		\a[6] ,
		\a[7] ,
		\a[12] ,
		\a[13] ,
		_w441_
	);
	LUT4 #(
		.INIT('h153f)
	) name376 (
		\a[2] ,
		\a[4] ,
		\a[15] ,
		\a[17] ,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		\a[4] ,
		\a[17] ,
		_w443_
	);
	LUT4 #(
		.INIT('h8000)
	) name378 (
		\a[2] ,
		\a[4] ,
		\a[15] ,
		\a[17] ,
		_w444_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name379 (
		\a[2] ,
		\a[4] ,
		\a[15] ,
		\a[17] ,
		_w445_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		\a[0] ,
		\a[19] ,
		_w446_
	);
	LUT4 #(
		.INIT('h0660)
	) name381 (
		_w438_,
		_w441_,
		_w445_,
		_w446_,
		_w447_
	);
	LUT4 #(
		.INIT('h6996)
	) name382 (
		_w438_,
		_w441_,
		_w445_,
		_w446_,
		_w448_
	);
	LUT4 #(
		.INIT('h2b00)
	) name383 (
		_w392_,
		_w393_,
		_w394_,
		_w448_,
		_w449_
	);
	LUT4 #(
		.INIT('hd42b)
	) name384 (
		_w392_,
		_w393_,
		_w394_,
		_w448_,
		_w450_
	);
	LUT4 #(
		.INIT('he800)
	) name385 (
		_w395_,
		_w396_,
		_w397_,
		_w450_,
		_w451_
	);
	LUT4 #(
		.INIT('h0017)
	) name386 (
		_w395_,
		_w396_,
		_w397_,
		_w450_,
		_w452_
	);
	LUT4 #(
		.INIT('h17e8)
	) name387 (
		_w395_,
		_w396_,
		_w397_,
		_w450_,
		_w453_
	);
	LUT2 #(
		.INIT('h6)
	) name388 (
		_w437_,
		_w453_,
		_w454_
	);
	LUT4 #(
		.INIT('hfee0)
	) name389 (
		_w372_,
		_w380_,
		_w398_,
		_w415_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		_w454_,
		_w455_,
		_w456_
	);
	LUT4 #(
		.INIT('h7887)
	) name391 (
		_w391_,
		_w416_,
		_w454_,
		_w455_,
		_w457_
	);
	LUT4 #(
		.INIT('h4f00)
	) name392 (
		_w348_,
		_w390_,
		_w419_,
		_w457_,
		_w458_
	);
	LUT4 #(
		.INIT('h0ff0)
	) name393 (
		_w391_,
		_w416_,
		_w454_,
		_w455_,
		_w459_
	);
	LUT4 #(
		.INIT('hb000)
	) name394 (
		_w348_,
		_w390_,
		_w419_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('he)
	) name395 (
		_w458_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w419_,
		_w456_,
		_w462_
	);
	LUT4 #(
		.INIT('h0888)
	) name397 (
		_w391_,
		_w416_,
		_w454_,
		_w455_,
		_w463_
	);
	LUT3 #(
		.INIT('h0e)
	) name398 (
		_w437_,
		_w451_,
		_w452_,
		_w464_
	);
	LUT3 #(
		.INIT('h45)
	) name399 (
		_w423_,
		_w424_,
		_w426_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\a[2] ,
		\a[18] ,
		_w466_
	);
	LUT4 #(
		.INIT('h153f)
	) name401 (
		\a[3] ,
		\a[4] ,
		\a[16] ,
		\a[17] ,
		_w467_
	);
	LUT4 #(
		.INIT('h8000)
	) name402 (
		\a[3] ,
		\a[4] ,
		\a[16] ,
		\a[17] ,
		_w468_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name403 (
		\a[3] ,
		\a[4] ,
		\a[16] ,
		\a[17] ,
		_w469_
	);
	LUT2 #(
		.INIT('h6)
	) name404 (
		_w466_,
		_w469_,
		_w470_
	);
	LUT4 #(
		.INIT('h4500)
	) name405 (
		_w423_,
		_w424_,
		_w426_,
		_w470_,
		_w471_
	);
	LUT4 #(
		.INIT('h00ba)
	) name406 (
		_w423_,
		_w424_,
		_w426_,
		_w470_,
		_w472_
	);
	LUT4 #(
		.INIT('hba45)
	) name407 (
		_w423_,
		_w424_,
		_w426_,
		_w470_,
		_w473_
	);
	LUT3 #(
		.INIT('he8)
	) name408 (
		_w428_,
		_w429_,
		_w435_,
		_w474_
	);
	LUT2 #(
		.INIT('h6)
	) name409 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT3 #(
		.INIT('hb2)
	) name410 (
		_w420_,
		_w427_,
		_w436_,
		_w476_
	);
	LUT4 #(
		.INIT('h8000)
	) name411 (
		\a[1] ,
		\a[9] ,
		\a[11] ,
		\a[19] ,
		_w477_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name412 (
		\a[1] ,
		\a[9] ,
		\a[11] ,
		\a[19] ,
		_w478_
	);
	LUT3 #(
		.INIT('h32)
	) name413 (
		_w405_,
		_w432_,
		_w433_,
		_w479_
	);
	LUT4 #(
		.INIT('he800)
	) name414 (
		_w405_,
		_w430_,
		_w431_,
		_w478_,
		_w480_
	);
	LUT4 #(
		.INIT('h0017)
	) name415 (
		_w405_,
		_w430_,
		_w431_,
		_w478_,
		_w481_
	);
	LUT4 #(
		.INIT('hcd32)
	) name416 (
		_w405_,
		_w432_,
		_w433_,
		_w478_,
		_w482_
	);
	LUT3 #(
		.INIT('h23)
	) name417 (
		_w442_,
		_w444_,
		_w446_,
		_w483_
	);
	LUT2 #(
		.INIT('h6)
	) name418 (
		_w482_,
		_w483_,
		_w484_
	);
	LUT4 #(
		.INIT('h153f)
	) name419 (
		\a[0] ,
		\a[7] ,
		\a[13] ,
		\a[20] ,
		_w485_
	);
	LUT4 #(
		.INIT('h8000)
	) name420 (
		\a[0] ,
		\a[7] ,
		\a[13] ,
		\a[20] ,
		_w486_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name421 (
		\a[0] ,
		\a[7] ,
		\a[13] ,
		\a[20] ,
		_w487_
	);
	LUT2 #(
		.INIT('h6)
	) name422 (
		_w421_,
		_w487_,
		_w488_
	);
	LUT3 #(
		.INIT('h0d)
	) name423 (
		_w438_,
		_w439_,
		_w440_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\a[8] ,
		\a[12] ,
		_w490_
	);
	LUT4 #(
		.INIT('h153f)
	) name425 (
		\a[5] ,
		\a[6] ,
		\a[14] ,
		\a[15] ,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\a[6] ,
		\a[15] ,
		_w492_
	);
	LUT4 #(
		.INIT('h8000)
	) name427 (
		\a[5] ,
		\a[6] ,
		\a[14] ,
		\a[15] ,
		_w493_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name428 (
		\a[5] ,
		\a[6] ,
		\a[14] ,
		\a[15] ,
		_w494_
	);
	LUT2 #(
		.INIT('h6)
	) name429 (
		_w490_,
		_w494_,
		_w495_
	);
	LUT3 #(
		.INIT('h69)
	) name430 (
		_w488_,
		_w489_,
		_w495_,
		_w496_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name431 (
		_w447_,
		_w449_,
		_w484_,
		_w496_,
		_w497_
	);
	LUT3 #(
		.INIT('h96)
	) name432 (
		_w475_,
		_w476_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w464_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h6)
	) name434 (
		_w464_,
		_w498_,
		_w500_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name435 (
		_w454_,
		_w455_,
		_w464_,
		_w498_,
		_w501_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		_w463_,
		_w501_,
		_w502_
	);
	LUT4 #(
		.INIT('h4f00)
	) name437 (
		_w348_,
		_w390_,
		_w462_,
		_w502_,
		_w503_
	);
	LUT4 #(
		.INIT('hf770)
	) name438 (
		_w391_,
		_w416_,
		_w454_,
		_w455_,
		_w504_
	);
	LUT4 #(
		.INIT('h4f00)
	) name439 (
		_w348_,
		_w390_,
		_w462_,
		_w504_,
		_w505_
	);
	LUT3 #(
		.INIT('h32)
	) name440 (
		_w500_,
		_w503_,
		_w505_,
		_w506_
	);
	LUT4 #(
		.INIT('heee0)
	) name441 (
		_w454_,
		_w455_,
		_w464_,
		_w498_,
		_w507_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w463_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('h4f00)
	) name443 (
		_w348_,
		_w390_,
		_w462_,
		_w508_,
		_w509_
	);
	LUT3 #(
		.INIT('h17)
	) name444 (
		_w475_,
		_w476_,
		_w497_,
		_w510_
	);
	LUT3 #(
		.INIT('h45)
	) name445 (
		_w471_,
		_w472_,
		_w474_,
		_w511_
	);
	LUT3 #(
		.INIT('h0d)
	) name446 (
		_w466_,
		_w467_,
		_w468_,
		_w512_
	);
	LUT3 #(
		.INIT('h0d)
	) name447 (
		_w490_,
		_w491_,
		_w493_,
		_w513_
	);
	LUT3 #(
		.INIT('h32)
	) name448 (
		_w421_,
		_w485_,
		_w486_,
		_w514_
	);
	LUT3 #(
		.INIT('h96)
	) name449 (
		_w512_,
		_w513_,
		_w514_,
		_w515_
	);
	LUT4 #(
		.INIT('he800)
	) name450 (
		_w465_,
		_w470_,
		_w474_,
		_w515_,
		_w516_
	);
	LUT4 #(
		.INIT('h153f)
	) name451 (
		\a[7] ,
		\a[8] ,
		\a[13] ,
		\a[14] ,
		_w517_
	);
	LUT4 #(
		.INIT('h8000)
	) name452 (
		\a[7] ,
		\a[8] ,
		\a[13] ,
		\a[14] ,
		_w518_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name453 (
		\a[7] ,
		\a[8] ,
		\a[13] ,
		\a[14] ,
		_w519_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\a[5] ,
		\a[16] ,
		_w520_
	);
	LUT4 #(
		.INIT('h153f)
	) name455 (
		\a[2] ,
		\a[3] ,
		\a[18] ,
		\a[19] ,
		_w521_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		\a[3] ,
		\a[19] ,
		_w522_
	);
	LUT4 #(
		.INIT('h8000)
	) name457 (
		\a[2] ,
		\a[3] ,
		\a[18] ,
		\a[19] ,
		_w523_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name458 (
		\a[2] ,
		\a[3] ,
		\a[18] ,
		\a[19] ,
		_w524_
	);
	LUT4 #(
		.INIT('h0660)
	) name459 (
		_w492_,
		_w519_,
		_w520_,
		_w524_,
		_w525_
	);
	LUT4 #(
		.INIT('h9009)
	) name460 (
		_w492_,
		_w519_,
		_w520_,
		_w524_,
		_w526_
	);
	LUT4 #(
		.INIT('h6996)
	) name461 (
		_w492_,
		_w519_,
		_w520_,
		_w524_,
		_w527_
	);
	LUT4 #(
		.INIT('h153f)
	) name462 (
		\a[9] ,
		\a[10] ,
		\a[11] ,
		\a[12] ,
		_w528_
	);
	LUT4 #(
		.INIT('h8000)
	) name463 (
		\a[9] ,
		\a[10] ,
		\a[11] ,
		\a[12] ,
		_w529_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name464 (
		\a[9] ,
		\a[10] ,
		\a[11] ,
		\a[12] ,
		_w530_
	);
	LUT2 #(
		.INIT('h6)
	) name465 (
		_w443_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h6)
	) name466 (
		_w527_,
		_w531_,
		_w532_
	);
	LUT4 #(
		.INIT('h0045)
	) name467 (
		_w471_,
		_w472_,
		_w474_,
		_w515_,
		_w533_
	);
	LUT4 #(
		.INIT('hf949)
	) name468 (
		_w511_,
		_w515_,
		_w532_,
		_w533_,
		_w534_
	);
	LUT3 #(
		.INIT('h23)
	) name469 (
		_w480_,
		_w481_,
		_w483_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		\a[0] ,
		\a[21] ,
		_w536_
	);
	LUT3 #(
		.INIT('h80)
	) name471 (
		\a[1] ,
		\a[11] ,
		\a[20] ,
		_w537_
	);
	LUT3 #(
		.INIT('h6c)
	) name472 (
		\a[1] ,
		\a[11] ,
		\a[20] ,
		_w538_
	);
	LUT3 #(
		.INIT('h96)
	) name473 (
		_w477_,
		_w536_,
		_w538_,
		_w539_
	);
	LUT4 #(
		.INIT('h0071)
	) name474 (
		_w478_,
		_w479_,
		_w483_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('h8e00)
	) name475 (
		_w478_,
		_w479_,
		_w483_,
		_w539_,
		_w541_
	);
	LUT4 #(
		.INIT('hdc23)
	) name476 (
		_w480_,
		_w481_,
		_w483_,
		_w539_,
		_w542_
	);
	LUT3 #(
		.INIT('hb2)
	) name477 (
		_w488_,
		_w489_,
		_w495_,
		_w543_
	);
	LUT2 #(
		.INIT('h6)
	) name478 (
		_w542_,
		_w543_,
		_w544_
	);
	LUT4 #(
		.INIT('hef0e)
	) name479 (
		_w447_,
		_w449_,
		_w484_,
		_w496_,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		_w544_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w544_,
		_w545_,
		_w547_
	);
	LUT2 #(
		.INIT('h6)
	) name482 (
		_w544_,
		_w545_,
		_w548_
	);
	LUT3 #(
		.INIT('h14)
	) name483 (
		_w510_,
		_w534_,
		_w548_,
		_w549_
	);
	LUT3 #(
		.INIT('h82)
	) name484 (
		_w510_,
		_w534_,
		_w548_,
		_w550_
	);
	LUT3 #(
		.INIT('h69)
	) name485 (
		_w510_,
		_w534_,
		_w548_,
		_w551_
	);
	LUT3 #(
		.INIT('h1e)
	) name486 (
		_w499_,
		_w509_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w499_,
		_w549_,
		_w553_
	);
	LUT3 #(
		.INIT('h0e)
	) name488 (
		_w534_,
		_w546_,
		_w547_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\a[0] ,
		\a[22] ,
		_w555_
	);
	LUT4 #(
		.INIT('h153f)
	) name490 (
		\a[7] ,
		\a[8] ,
		\a[14] ,
		\a[15] ,
		_w556_
	);
	LUT4 #(
		.INIT('h8000)
	) name491 (
		\a[7] ,
		\a[8] ,
		\a[14] ,
		\a[15] ,
		_w557_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name492 (
		\a[7] ,
		\a[8] ,
		\a[14] ,
		\a[15] ,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		\a[9] ,
		\a[13] ,
		_w559_
	);
	LUT4 #(
		.INIT('h153f)
	) name494 (
		\a[2] ,
		\a[6] ,
		\a[16] ,
		\a[20] ,
		_w560_
	);
	LUT4 #(
		.INIT('h8000)
	) name495 (
		\a[2] ,
		\a[6] ,
		\a[16] ,
		\a[20] ,
		_w561_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name496 (
		\a[2] ,
		\a[6] ,
		\a[16] ,
		\a[20] ,
		_w562_
	);
	LUT4 #(
		.INIT('h0660)
	) name497 (
		_w555_,
		_w558_,
		_w559_,
		_w562_,
		_w563_
	);
	LUT4 #(
		.INIT('h9009)
	) name498 (
		_w555_,
		_w558_,
		_w559_,
		_w562_,
		_w564_
	);
	LUT4 #(
		.INIT('h6996)
	) name499 (
		_w555_,
		_w558_,
		_w559_,
		_w562_,
		_w565_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\a[4] ,
		\a[19] ,
		_w566_
	);
	LUT4 #(
		.INIT('h8000)
	) name501 (
		\a[3] ,
		\a[4] ,
		\a[18] ,
		\a[19] ,
		_w567_
	);
	LUT4 #(
		.INIT('h8000)
	) name502 (
		\a[3] ,
		\a[5] ,
		\a[17] ,
		\a[19] ,
		_w568_
	);
	LUT4 #(
		.INIT('h8000)
	) name503 (
		\a[4] ,
		\a[5] ,
		\a[17] ,
		\a[18] ,
		_w569_
	);
	LUT3 #(
		.INIT('h0e)
	) name504 (
		_w567_,
		_w568_,
		_w569_,
		_w570_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name505 (
		\a[4] ,
		\a[5] ,
		\a[17] ,
		\a[18] ,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w522_,
		_w571_,
		_w572_
	);
	LUT3 #(
		.INIT('h01)
	) name507 (
		_w565_,
		_w570_,
		_w572_,
		_w573_
	);
	LUT3 #(
		.INIT('h0d)
	) name508 (
		_w520_,
		_w521_,
		_w523_,
		_w574_
	);
	LUT3 #(
		.INIT('h0d)
	) name509 (
		_w492_,
		_w517_,
		_w518_,
		_w575_
	);
	LUT3 #(
		.INIT('he8)
	) name510 (
		_w477_,
		_w536_,
		_w538_,
		_w576_
	);
	LUT3 #(
		.INIT('h96)
	) name511 (
		_w574_,
		_w575_,
		_w576_,
		_w577_
	);
	LUT4 #(
		.INIT('h00e8)
	) name512 (
		_w535_,
		_w539_,
		_w543_,
		_w577_,
		_w578_
	);
	LUT3 #(
		.INIT('ha8)
	) name513 (
		_w565_,
		_w570_,
		_w572_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w577_,
		_w579_,
		_w580_
	);
	LUT4 #(
		.INIT('h00e8)
	) name515 (
		_w535_,
		_w539_,
		_w543_,
		_w579_,
		_w581_
	);
	LUT4 #(
		.INIT('h1110)
	) name516 (
		_w573_,
		_w578_,
		_w580_,
		_w581_,
		_w582_
	);
	LUT3 #(
		.INIT('h54)
	) name517 (
		_w540_,
		_w541_,
		_w543_,
		_w583_
	);
	LUT3 #(
		.INIT('h56)
	) name518 (
		_w565_,
		_w570_,
		_w572_,
		_w584_
	);
	LUT3 #(
		.INIT('hf9)
	) name519 (
		_w577_,
		_w583_,
		_w584_,
		_w585_
	);
	LUT3 #(
		.INIT('h71)
	) name520 (
		_w512_,
		_w513_,
		_w514_,
		_w586_
	);
	LUT4 #(
		.INIT('h8000)
	) name521 (
		\a[1] ,
		\a[10] ,
		\a[12] ,
		\a[21] ,
		_w587_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name522 (
		\a[1] ,
		\a[10] ,
		\a[12] ,
		\a[21] ,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		_w537_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w537_,
		_w588_,
		_w590_
	);
	LUT2 #(
		.INIT('h6)
	) name525 (
		_w537_,
		_w588_,
		_w591_
	);
	LUT3 #(
		.INIT('h0d)
	) name526 (
		_w443_,
		_w528_,
		_w529_,
		_w592_
	);
	LUT2 #(
		.INIT('h6)
	) name527 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT3 #(
		.INIT('h32)
	) name528 (
		_w525_,
		_w526_,
		_w531_,
		_w594_
	);
	LUT3 #(
		.INIT('h69)
	) name529 (
		_w586_,
		_w593_,
		_w594_,
		_w595_
	);
	LUT4 #(
		.INIT('hae00)
	) name530 (
		_w516_,
		_w532_,
		_w533_,
		_w595_,
		_w596_
	);
	LUT4 #(
		.INIT('h0051)
	) name531 (
		_w516_,
		_w532_,
		_w533_,
		_w595_,
		_w597_
	);
	LUT4 #(
		.INIT('h51ae)
	) name532 (
		_w516_,
		_w532_,
		_w533_,
		_w595_,
		_w598_
	);
	LUT3 #(
		.INIT('h0b)
	) name533 (
		_w582_,
		_w585_,
		_w598_,
		_w599_
	);
	LUT4 #(
		.INIT('h0004)
	) name534 (
		_w582_,
		_w585_,
		_w596_,
		_w597_,
		_w600_
	);
	LUT4 #(
		.INIT('h444b)
	) name535 (
		_w582_,
		_w585_,
		_w596_,
		_w597_,
		_w601_
	);
	LUT3 #(
		.INIT('h02)
	) name536 (
		_w554_,
		_w599_,
		_w600_,
		_w602_
	);
	LUT4 #(
		.INIT('h4441)
	) name537 (
		_w550_,
		_w554_,
		_w599_,
		_w600_,
		_w603_
	);
	LUT3 #(
		.INIT('hb0)
	) name538 (
		_w509_,
		_w553_,
		_w603_,
		_w604_
	);
	LUT3 #(
		.INIT('ha9)
	) name539 (
		_w554_,
		_w599_,
		_w600_,
		_w605_
	);
	LUT4 #(
		.INIT('h2228)
	) name540 (
		_w550_,
		_w554_,
		_w599_,
		_w600_,
		_w606_
	);
	LUT4 #(
		.INIT('h00fb)
	) name541 (
		_w509_,
		_w553_,
		_w605_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w604_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		_w553_,
		_w602_,
		_w609_
	);
	LUT4 #(
		.INIT('haaa2)
	) name544 (
		_w550_,
		_w554_,
		_w599_,
		_w600_,
		_w610_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name545 (
		_w582_,
		_w585_,
		_w596_,
		_w597_,
		_w611_
	);
	LUT3 #(
		.INIT('hb2)
	) name546 (
		_w586_,
		_w593_,
		_w594_,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		\a[6] ,
		\a[17] ,
		_w613_
	);
	LUT4 #(
		.INIT('h153f)
	) name548 (
		\a[3] ,
		\a[5] ,
		\a[18] ,
		\a[20] ,
		_w614_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\a[5] ,
		\a[20] ,
		_w615_
	);
	LUT4 #(
		.INIT('h8000)
	) name550 (
		\a[3] ,
		\a[5] ,
		\a[18] ,
		\a[20] ,
		_w616_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name551 (
		\a[3] ,
		\a[5] ,
		\a[18] ,
		\a[20] ,
		_w617_
	);
	LUT4 #(
		.INIT('h153f)
	) name552 (
		\a[10] ,
		\a[11] ,
		\a[12] ,
		\a[13] ,
		_w618_
	);
	LUT4 #(
		.INIT('h8000)
	) name553 (
		\a[10] ,
		\a[11] ,
		\a[12] ,
		\a[13] ,
		_w619_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name554 (
		\a[10] ,
		\a[11] ,
		\a[12] ,
		\a[13] ,
		_w620_
	);
	LUT4 #(
		.INIT('h1428)
	) name555 (
		_w566_,
		_w613_,
		_w617_,
		_w620_,
		_w621_
	);
	LUT4 #(
		.INIT('h8241)
	) name556 (
		_w566_,
		_w613_,
		_w617_,
		_w620_,
		_w622_
	);
	LUT4 #(
		.INIT('h6996)
	) name557 (
		_w566_,
		_w613_,
		_w617_,
		_w620_,
		_w623_
	);
	LUT4 #(
		.INIT('hdc23)
	) name558 (
		_w589_,
		_w590_,
		_w592_,
		_w623_,
		_w624_
	);
	LUT4 #(
		.INIT('h153f)
	) name559 (
		\a[0] ,
		\a[2] ,
		\a[21] ,
		\a[23] ,
		_w625_
	);
	LUT4 #(
		.INIT('h8000)
	) name560 (
		\a[0] ,
		\a[2] ,
		\a[21] ,
		\a[23] ,
		_w626_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name561 (
		\a[0] ,
		\a[2] ,
		\a[21] ,
		\a[23] ,
		_w627_
	);
	LUT2 #(
		.INIT('h6)
	) name562 (
		_w587_,
		_w627_,
		_w628_
	);
	LUT3 #(
		.INIT('h0d)
	) name563 (
		_w555_,
		_w556_,
		_w557_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name564 (
		\a[7] ,
		\a[16] ,
		_w630_
	);
	LUT4 #(
		.INIT('h153f)
	) name565 (
		\a[8] ,
		\a[9] ,
		\a[14] ,
		\a[15] ,
		_w631_
	);
	LUT4 #(
		.INIT('h8000)
	) name566 (
		\a[8] ,
		\a[9] ,
		\a[14] ,
		\a[15] ,
		_w632_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name567 (
		\a[8] ,
		\a[9] ,
		\a[14] ,
		\a[15] ,
		_w633_
	);
	LUT2 #(
		.INIT('h6)
	) name568 (
		_w630_,
		_w633_,
		_w634_
	);
	LUT3 #(
		.INIT('h69)
	) name569 (
		_w628_,
		_w629_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w624_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		_w624_,
		_w635_,
		_w637_
	);
	LUT2 #(
		.INIT('h6)
	) name572 (
		_w624_,
		_w635_,
		_w638_
	);
	LUT2 #(
		.INIT('h6)
	) name573 (
		_w612_,
		_w638_,
		_w639_
	);
	LUT4 #(
		.INIT('hff31)
	) name574 (
		_w577_,
		_w578_,
		_w583_,
		_w584_,
		_w640_
	);
	LUT4 #(
		.INIT('he800)
	) name575 (
		_w535_,
		_w539_,
		_w543_,
		_w577_,
		_w641_
	);
	LUT3 #(
		.INIT('h71)
	) name576 (
		_w574_,
		_w575_,
		_w576_,
		_w642_
	);
	LUT4 #(
		.INIT('h2223)
	) name577 (
		_w563_,
		_w564_,
		_w570_,
		_w572_,
		_w643_
	);
	LUT3 #(
		.INIT('h80)
	) name578 (
		\a[1] ,
		\a[12] ,
		\a[22] ,
		_w644_
	);
	LUT3 #(
		.INIT('h6c)
	) name579 (
		\a[1] ,
		\a[12] ,
		\a[22] ,
		_w645_
	);
	LUT4 #(
		.INIT('h0001)
	) name580 (
		_w567_,
		_w568_,
		_w569_,
		_w645_,
		_w646_
	);
	LUT4 #(
		.INIT('hfe00)
	) name581 (
		_w567_,
		_w568_,
		_w569_,
		_w645_,
		_w647_
	);
	LUT4 #(
		.INIT('h01fe)
	) name582 (
		_w567_,
		_w568_,
		_w569_,
		_w645_,
		_w648_
	);
	LUT3 #(
		.INIT('h32)
	) name583 (
		_w559_,
		_w560_,
		_w561_,
		_w649_
	);
	LUT2 #(
		.INIT('h6)
	) name584 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT3 #(
		.INIT('h96)
	) name585 (
		_w642_,
		_w643_,
		_w650_,
		_w651_
	);
	LUT4 #(
		.INIT('ha659)
	) name586 (
		_w639_,
		_w640_,
		_w641_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		_w611_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		_w611_,
		_w652_,
		_w654_
	);
	LUT2 #(
		.INIT('h9)
	) name589 (
		_w611_,
		_w652_,
		_w655_
	);
	LUT4 #(
		.INIT('he00e)
	) name590 (
		_w554_,
		_w601_,
		_w611_,
		_w652_,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		_w610_,
		_w656_,
		_w657_
	);
	LUT3 #(
		.INIT('hb0)
	) name592 (
		_w509_,
		_w609_,
		_w657_,
		_w658_
	);
	LUT4 #(
		.INIT('h444d)
	) name593 (
		_w550_,
		_w554_,
		_w599_,
		_w600_,
		_w659_
	);
	LUT4 #(
		.INIT('h040f)
	) name594 (
		_w509_,
		_w609_,
		_w655_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w658_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		_w653_,
		_w659_,
		_w662_
	);
	LUT4 #(
		.INIT('hfba2)
	) name597 (
		_w639_,
		_w640_,
		_w641_,
		_w651_,
		_w663_
	);
	LUT3 #(
		.INIT('h54)
	) name598 (
		_w646_,
		_w647_,
		_w649_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		\a[0] ,
		\a[24] ,
		_w665_
	);
	LUT4 #(
		.INIT('h8000)
	) name600 (
		\a[1] ,
		\a[11] ,
		\a[13] ,
		\a[23] ,
		_w666_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name601 (
		\a[1] ,
		\a[11] ,
		\a[13] ,
		\a[23] ,
		_w667_
	);
	LUT3 #(
		.INIT('h96)
	) name602 (
		_w644_,
		_w665_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h8)
	) name603 (
		\a[7] ,
		\a[17] ,
		_w669_
	);
	LUT4 #(
		.INIT('h153f)
	) name604 (
		\a[2] ,
		\a[6] ,
		\a[18] ,
		\a[22] ,
		_w670_
	);
	LUT4 #(
		.INIT('h8000)
	) name605 (
		\a[2] ,
		\a[6] ,
		\a[18] ,
		\a[22] ,
		_w671_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name606 (
		\a[2] ,
		\a[6] ,
		\a[18] ,
		\a[22] ,
		_w672_
	);
	LUT2 #(
		.INIT('h6)
	) name607 (
		_w669_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		_w668_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w668_,
		_w673_,
		_w675_
	);
	LUT2 #(
		.INIT('h6)
	) name610 (
		_w668_,
		_w673_,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		\a[3] ,
		\a[21] ,
		_w677_
	);
	LUT4 #(
		.INIT('h153f)
	) name612 (
		\a[4] ,
		\a[5] ,
		\a[19] ,
		\a[20] ,
		_w678_
	);
	LUT4 #(
		.INIT('h8000)
	) name613 (
		\a[4] ,
		\a[5] ,
		\a[19] ,
		\a[20] ,
		_w679_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name614 (
		\a[4] ,
		\a[5] ,
		\a[19] ,
		\a[20] ,
		_w680_
	);
	LUT2 #(
		.INIT('h6)
	) name615 (
		_w677_,
		_w680_,
		_w681_
	);
	LUT3 #(
		.INIT('h0d)
	) name616 (
		_w587_,
		_w625_,
		_w626_,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\a[8] ,
		\a[16] ,
		_w683_
	);
	LUT4 #(
		.INIT('h153f)
	) name618 (
		\a[9] ,
		\a[10] ,
		\a[14] ,
		\a[15] ,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		\a[10] ,
		\a[15] ,
		_w685_
	);
	LUT4 #(
		.INIT('h8000)
	) name620 (
		\a[9] ,
		\a[10] ,
		\a[14] ,
		\a[15] ,
		_w686_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name621 (
		\a[9] ,
		\a[10] ,
		\a[14] ,
		\a[15] ,
		_w687_
	);
	LUT2 #(
		.INIT('h6)
	) name622 (
		_w683_,
		_w687_,
		_w688_
	);
	LUT3 #(
		.INIT('h69)
	) name623 (
		_w681_,
		_w682_,
		_w688_,
		_w689_
	);
	LUT3 #(
		.INIT('h09)
	) name624 (
		_w664_,
		_w676_,
		_w689_,
		_w690_
	);
	LUT3 #(
		.INIT('h60)
	) name625 (
		_w664_,
		_w676_,
		_w689_,
		_w691_
	);
	LUT3 #(
		.INIT('h96)
	) name626 (
		_w664_,
		_w676_,
		_w689_,
		_w692_
	);
	LUT3 #(
		.INIT('he8)
	) name627 (
		_w642_,
		_w643_,
		_w650_,
		_w693_
	);
	LUT2 #(
		.INIT('h6)
	) name628 (
		_w692_,
		_w693_,
		_w694_
	);
	LUT3 #(
		.INIT('h0d)
	) name629 (
		_w566_,
		_w618_,
		_w619_,
		_w695_
	);
	LUT3 #(
		.INIT('h0d)
	) name630 (
		_w613_,
		_w614_,
		_w616_,
		_w696_
	);
	LUT3 #(
		.INIT('h0d)
	) name631 (
		_w630_,
		_w631_,
		_w632_,
		_w697_
	);
	LUT3 #(
		.INIT('h96)
	) name632 (
		_w695_,
		_w696_,
		_w697_,
		_w698_
	);
	LUT4 #(
		.INIT('h0071)
	) name633 (
		_w537_,
		_w588_,
		_w592_,
		_w621_,
		_w699_
	);
	LUT3 #(
		.INIT('hb2)
	) name634 (
		_w628_,
		_w629_,
		_w634_,
		_w700_
	);
	LUT3 #(
		.INIT('h0e)
	) name635 (
		_w622_,
		_w699_,
		_w700_,
		_w701_
	);
	LUT4 #(
		.INIT('hc936)
	) name636 (
		_w622_,
		_w698_,
		_w699_,
		_w700_,
		_w702_
	);
	LUT4 #(
		.INIT('he800)
	) name637 (
		_w612_,
		_w624_,
		_w635_,
		_w702_,
		_w703_
	);
	LUT4 #(
		.INIT('h0017)
	) name638 (
		_w612_,
		_w624_,
		_w635_,
		_w702_,
		_w704_
	);
	LUT4 #(
		.INIT('hcd32)
	) name639 (
		_w612_,
		_w636_,
		_w637_,
		_w702_,
		_w705_
	);
	LUT2 #(
		.INIT('h6)
	) name640 (
		_w694_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name641 (
		_w663_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h6)
	) name642 (
		_w663_,
		_w706_,
		_w708_
	);
	LUT4 #(
		.INIT('h0bb0)
	) name643 (
		_w611_,
		_w652_,
		_w663_,
		_w706_,
		_w709_
	);
	LUT4 #(
		.INIT('h4f00)
	) name644 (
		_w509_,
		_w609_,
		_w662_,
		_w709_,
		_w710_
	);
	LUT4 #(
		.INIT('h040f)
	) name645 (
		_w509_,
		_w609_,
		_w654_,
		_w662_,
		_w711_
	);
	LUT3 #(
		.INIT('hcd)
	) name646 (
		_w708_,
		_w710_,
		_w711_,
		_w712_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name647 (
		_w611_,
		_w652_,
		_w663_,
		_w706_,
		_w713_
	);
	LUT4 #(
		.INIT('h4f00)
	) name648 (
		_w509_,
		_w609_,
		_w662_,
		_w713_,
		_w714_
	);
	LUT3 #(
		.INIT('h31)
	) name649 (
		_w694_,
		_w703_,
		_w704_,
		_w715_
	);
	LUT3 #(
		.INIT('h0d)
	) name650 (
		_w669_,
		_w670_,
		_w671_,
		_w716_
	);
	LUT3 #(
		.INIT('h0d)
	) name651 (
		_w683_,
		_w684_,
		_w686_,
		_w717_
	);
	LUT3 #(
		.INIT('he8)
	) name652 (
		_w644_,
		_w665_,
		_w667_,
		_w718_
	);
	LUT3 #(
		.INIT('h96)
	) name653 (
		_w716_,
		_w717_,
		_w718_,
		_w719_
	);
	LUT3 #(
		.INIT('hb2)
	) name654 (
		_w681_,
		_w682_,
		_w688_,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		_w719_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h6)
	) name656 (
		_w719_,
		_w720_,
		_w722_
	);
	LUT3 #(
		.INIT('h0e)
	) name657 (
		_w664_,
		_w674_,
		_w675_,
		_w723_
	);
	LUT2 #(
		.INIT('h6)
	) name658 (
		_w722_,
		_w723_,
		_w724_
	);
	LUT3 #(
		.INIT('h54)
	) name659 (
		_w690_,
		_w691_,
		_w693_,
		_w725_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name660 (
		_w622_,
		_w698_,
		_w699_,
		_w700_,
		_w726_
	);
	LUT4 #(
		.INIT('h153f)
	) name661 (
		\a[0] ,
		\a[2] ,
		\a[23] ,
		\a[25] ,
		_w727_
	);
	LUT4 #(
		.INIT('h8000)
	) name662 (
		\a[0] ,
		\a[2] ,
		\a[23] ,
		\a[25] ,
		_w728_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name663 (
		\a[0] ,
		\a[2] ,
		\a[23] ,
		\a[25] ,
		_w729_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		\a[7] ,
		\a[18] ,
		_w730_
	);
	LUT4 #(
		.INIT('h153f)
	) name665 (
		\a[8] ,
		\a[9] ,
		\a[16] ,
		\a[17] ,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		\a[9] ,
		\a[17] ,
		_w732_
	);
	LUT4 #(
		.INIT('h8000)
	) name667 (
		\a[8] ,
		\a[9] ,
		\a[16] ,
		\a[17] ,
		_w733_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name668 (
		\a[8] ,
		\a[9] ,
		\a[16] ,
		\a[17] ,
		_w734_
	);
	LUT4 #(
		.INIT('h0660)
	) name669 (
		_w685_,
		_w729_,
		_w730_,
		_w734_,
		_w735_
	);
	LUT4 #(
		.INIT('h9009)
	) name670 (
		_w685_,
		_w729_,
		_w730_,
		_w734_,
		_w736_
	);
	LUT4 #(
		.INIT('h6996)
	) name671 (
		_w685_,
		_w729_,
		_w730_,
		_w734_,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name672 (
		\a[6] ,
		\a[19] ,
		_w738_
	);
	LUT4 #(
		.INIT('h153f)
	) name673 (
		\a[3] ,
		\a[4] ,
		\a[21] ,
		\a[22] ,
		_w739_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		\a[4] ,
		\a[22] ,
		_w740_
	);
	LUT4 #(
		.INIT('h8000)
	) name675 (
		\a[3] ,
		\a[4] ,
		\a[21] ,
		\a[22] ,
		_w741_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name676 (
		\a[3] ,
		\a[4] ,
		\a[21] ,
		\a[22] ,
		_w742_
	);
	LUT2 #(
		.INIT('h6)
	) name677 (
		_w738_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h6)
	) name678 (
		_w737_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		\a[12] ,
		\a[13] ,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		\a[11] ,
		\a[14] ,
		_w746_
	);
	LUT4 #(
		.INIT('h153f)
	) name681 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w747_
	);
	LUT4 #(
		.INIT('h8000)
	) name682 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w748_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name683 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w749_
	);
	LUT2 #(
		.INIT('h6)
	) name684 (
		_w615_,
		_w749_,
		_w750_
	);
	LUT4 #(
		.INIT('h00e8)
	) name685 (
		_w695_,
		_w696_,
		_w697_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		\a[1] ,
		\a[24] ,
		_w752_
	);
	LUT3 #(
		.INIT('h2d)
	) name687 (
		\a[13] ,
		_w666_,
		_w752_,
		_w753_
	);
	LUT3 #(
		.INIT('h0d)
	) name688 (
		_w677_,
		_w678_,
		_w679_,
		_w754_
	);
	LUT2 #(
		.INIT('h6)
	) name689 (
		_w753_,
		_w754_,
		_w755_
	);
	LUT4 #(
		.INIT('h1700)
	) name690 (
		_w695_,
		_w696_,
		_w697_,
		_w750_,
		_w756_
	);
	LUT3 #(
		.INIT('hc9)
	) name691 (
		_w751_,
		_w755_,
		_w756_,
		_w757_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name692 (
		_w701_,
		_w726_,
		_w744_,
		_w757_,
		_w758_
	);
	LUT3 #(
		.INIT('h96)
	) name693 (
		_w724_,
		_w725_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name694 (
		_w715_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		_w715_,
		_w759_,
		_w761_
	);
	LUT2 #(
		.INIT('h9)
	) name696 (
		_w715_,
		_w759_,
		_w762_
	);
	LUT3 #(
		.INIT('he1)
	) name697 (
		_w707_,
		_w714_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h2)
	) name698 (
		_w713_,
		_w761_,
		_w764_
	);
	LUT4 #(
		.INIT('h4f00)
	) name699 (
		_w509_,
		_w609_,
		_w662_,
		_w764_,
		_w765_
	);
	LUT4 #(
		.INIT('h1011)
	) name700 (
		_w663_,
		_w706_,
		_w715_,
		_w759_,
		_w766_
	);
	LUT3 #(
		.INIT('h17)
	) name701 (
		_w724_,
		_w725_,
		_w758_,
		_w767_
	);
	LUT4 #(
		.INIT('hf110)
	) name702 (
		_w701_,
		_w726_,
		_w744_,
		_w757_,
		_w768_
	);
	LUT3 #(
		.INIT('h54)
	) name703 (
		_w751_,
		_w755_,
		_w756_,
		_w769_
	);
	LUT4 #(
		.INIT('h8000)
	) name704 (
		\a[1] ,
		\a[12] ,
		\a[14] ,
		\a[25] ,
		_w770_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name705 (
		\a[1] ,
		\a[12] ,
		\a[14] ,
		\a[25] ,
		_w771_
	);
	LUT4 #(
		.INIT('he800)
	) name706 (
		_w615_,
		_w745_,
		_w746_,
		_w771_,
		_w772_
	);
	LUT4 #(
		.INIT('h0017)
	) name707 (
		_w615_,
		_w745_,
		_w746_,
		_w771_,
		_w773_
	);
	LUT4 #(
		.INIT('hcd32)
	) name708 (
		_w615_,
		_w747_,
		_w748_,
		_w771_,
		_w774_
	);
	LUT3 #(
		.INIT('h0d)
	) name709 (
		_w738_,
		_w739_,
		_w741_,
		_w775_
	);
	LUT2 #(
		.INIT('h6)
	) name710 (
		_w774_,
		_w775_,
		_w776_
	);
	LUT3 #(
		.INIT('h32)
	) name711 (
		_w735_,
		_w736_,
		_w743_,
		_w777_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		_w776_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h9)
	) name713 (
		_w776_,
		_w777_,
		_w779_
	);
	LUT2 #(
		.INIT('h6)
	) name714 (
		_w769_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		_w768_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		_w768_,
		_w780_,
		_w782_
	);
	LUT2 #(
		.INIT('h6)
	) name717 (
		_w768_,
		_w780_,
		_w783_
	);
	LUT4 #(
		.INIT('h153f)
	) name718 (
		\a[10] ,
		\a[11] ,
		\a[15] ,
		\a[16] ,
		_w784_
	);
	LUT2 #(
		.INIT('h8)
	) name719 (
		\a[11] ,
		\a[16] ,
		_w785_
	);
	LUT4 #(
		.INIT('h8000)
	) name720 (
		\a[10] ,
		\a[11] ,
		\a[15] ,
		\a[16] ,
		_w786_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name721 (
		\a[10] ,
		\a[11] ,
		\a[15] ,
		\a[16] ,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\a[2] ,
		\a[24] ,
		_w788_
	);
	LUT4 #(
		.INIT('h153f)
	) name723 (
		\a[3] ,
		\a[7] ,
		\a[19] ,
		\a[23] ,
		_w789_
	);
	LUT4 #(
		.INIT('h8000)
	) name724 (
		\a[3] ,
		\a[7] ,
		\a[19] ,
		\a[23] ,
		_w790_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name725 (
		\a[3] ,
		\a[7] ,
		\a[19] ,
		\a[23] ,
		_w791_
	);
	LUT4 #(
		.INIT('h0660)
	) name726 (
		_w732_,
		_w787_,
		_w788_,
		_w791_,
		_w792_
	);
	LUT4 #(
		.INIT('h9009)
	) name727 (
		_w732_,
		_w787_,
		_w788_,
		_w791_,
		_w793_
	);
	LUT4 #(
		.INIT('h6996)
	) name728 (
		_w732_,
		_w787_,
		_w788_,
		_w791_,
		_w794_
	);
	LUT4 #(
		.INIT('h153f)
	) name729 (
		\a[5] ,
		\a[6] ,
		\a[20] ,
		\a[21] ,
		_w795_
	);
	LUT4 #(
		.INIT('h8000)
	) name730 (
		\a[5] ,
		\a[6] ,
		\a[20] ,
		\a[21] ,
		_w796_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name731 (
		\a[5] ,
		\a[6] ,
		\a[20] ,
		\a[21] ,
		_w797_
	);
	LUT2 #(
		.INIT('h6)
	) name732 (
		_w740_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h6)
	) name733 (
		_w794_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('h0017)
	) name734 (
		_w719_,
		_w720_,
		_w723_,
		_w799_,
		_w800_
	);
	LUT3 #(
		.INIT('he0)
	) name735 (
		_w719_,
		_w720_,
		_w799_,
		_w801_
	);
	LUT3 #(
		.INIT('he0)
	) name736 (
		_w721_,
		_w723_,
		_w801_,
		_w802_
	);
	LUT3 #(
		.INIT('h71)
	) name737 (
		_w716_,
		_w717_,
		_w718_,
		_w803_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		\a[24] ,
		_w666_,
		_w804_
	);
	LUT4 #(
		.INIT('h5093)
	) name739 (
		\a[1] ,
		\a[13] ,
		\a[24] ,
		_w666_,
		_w805_
	);
	LUT3 #(
		.INIT('h0d)
	) name740 (
		_w754_,
		_w804_,
		_w805_,
		_w806_
	);
	LUT3 #(
		.INIT('h0d)
	) name741 (
		_w730_,
		_w731_,
		_w733_,
		_w807_
	);
	LUT3 #(
		.INIT('h0d)
	) name742 (
		_w685_,
		_w727_,
		_w728_,
		_w808_
	);
	LUT3 #(
		.INIT('h80)
	) name743 (
		\a[1] ,
		\a[13] ,
		\a[24] ,
		_w809_
	);
	LUT4 #(
		.INIT('h153f)
	) name744 (
		\a[0] ,
		\a[8] ,
		\a[18] ,
		\a[26] ,
		_w810_
	);
	LUT4 #(
		.INIT('h8000)
	) name745 (
		\a[0] ,
		\a[8] ,
		\a[18] ,
		\a[26] ,
		_w811_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name746 (
		\a[0] ,
		\a[8] ,
		\a[18] ,
		\a[26] ,
		_w812_
	);
	LUT2 #(
		.INIT('h6)
	) name747 (
		_w809_,
		_w812_,
		_w813_
	);
	LUT3 #(
		.INIT('h69)
	) name748 (
		_w807_,
		_w808_,
		_w813_,
		_w814_
	);
	LUT3 #(
		.INIT('h69)
	) name749 (
		_w803_,
		_w806_,
		_w814_,
		_w815_
	);
	LUT3 #(
		.INIT('he1)
	) name750 (
		_w800_,
		_w802_,
		_w815_,
		_w816_
	);
	LUT3 #(
		.INIT('h14)
	) name751 (
		_w767_,
		_w783_,
		_w816_,
		_w817_
	);
	LUT3 #(
		.INIT('h82)
	) name752 (
		_w767_,
		_w783_,
		_w816_,
		_w818_
	);
	LUT3 #(
		.INIT('h69)
	) name753 (
		_w767_,
		_w783_,
		_w816_,
		_w819_
	);
	LUT4 #(
		.INIT('hfe01)
	) name754 (
		_w760_,
		_w765_,
		_w766_,
		_w819_,
		_w820_
	);
	LUT3 #(
		.INIT('h01)
	) name755 (
		_w760_,
		_w766_,
		_w818_,
		_w821_
	);
	LUT3 #(
		.INIT('h32)
	) name756 (
		_w781_,
		_w782_,
		_w816_,
		_w822_
	);
	LUT4 #(
		.INIT('h001f)
	) name757 (
		_w721_,
		_w723_,
		_w801_,
		_w815_,
		_w823_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w800_,
		_w823_,
		_w824_
	);
	LUT3 #(
		.INIT('h8e)
	) name759 (
		_w803_,
		_w806_,
		_w814_,
		_w825_
	);
	LUT3 #(
		.INIT('h0d)
	) name760 (
		_w732_,
		_w784_,
		_w786_,
		_w826_
	);
	LUT3 #(
		.INIT('h0d)
	) name761 (
		_w740_,
		_w795_,
		_w796_,
		_w827_
	);
	LUT3 #(
		.INIT('h32)
	) name762 (
		_w788_,
		_w789_,
		_w790_,
		_w828_
	);
	LUT3 #(
		.INIT('h96)
	) name763 (
		_w826_,
		_w827_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		\a[0] ,
		\a[27] ,
		_w830_
	);
	LUT3 #(
		.INIT('h93)
	) name765 (
		\a[1] ,
		\a[14] ,
		\a[26] ,
		_w831_
	);
	LUT3 #(
		.INIT('h69)
	) name766 (
		_w770_,
		_w830_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name767 (
		\a[5] ,
		\a[22] ,
		_w833_
	);
	LUT4 #(
		.INIT('h153f)
	) name768 (
		\a[12] ,
		\a[13] ,
		\a[14] ,
		\a[15] ,
		_w834_
	);
	LUT4 #(
		.INIT('h8000)
	) name769 (
		\a[12] ,
		\a[13] ,
		\a[14] ,
		\a[15] ,
		_w835_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name770 (
		\a[12] ,
		\a[13] ,
		\a[14] ,
		\a[15] ,
		_w836_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		\a[3] ,
		\a[24] ,
		_w837_
	);
	LUT4 #(
		.INIT('h153f)
	) name772 (
		\a[4] ,
		\a[6] ,
		\a[21] ,
		\a[23] ,
		_w838_
	);
	LUT4 #(
		.INIT('h8000)
	) name773 (
		\a[4] ,
		\a[6] ,
		\a[21] ,
		\a[23] ,
		_w839_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name774 (
		\a[4] ,
		\a[6] ,
		\a[21] ,
		\a[23] ,
		_w840_
	);
	LUT4 #(
		.INIT('h0660)
	) name775 (
		_w833_,
		_w836_,
		_w837_,
		_w840_,
		_w841_
	);
	LUT4 #(
		.INIT('h9009)
	) name776 (
		_w833_,
		_w836_,
		_w837_,
		_w840_,
		_w842_
	);
	LUT4 #(
		.INIT('h6996)
	) name777 (
		_w833_,
		_w836_,
		_w837_,
		_w840_,
		_w843_
	);
	LUT2 #(
		.INIT('h6)
	) name778 (
		_w832_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		_w829_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		_w829_,
		_w844_,
		_w846_
	);
	LUT3 #(
		.INIT('h9f)
	) name781 (
		_w825_,
		_w829_,
		_w844_,
		_w847_
	);
	LUT3 #(
		.INIT('h96)
	) name782 (
		_w825_,
		_w829_,
		_w844_,
		_w848_
	);
	LUT3 #(
		.INIT('h10)
	) name783 (
		_w800_,
		_w823_,
		_w848_,
		_w849_
	);
	LUT3 #(
		.INIT('h0e)
	) name784 (
		_w800_,
		_w823_,
		_w848_,
		_w850_
	);
	LUT3 #(
		.INIT('he1)
	) name785 (
		_w800_,
		_w823_,
		_w848_,
		_w851_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w776_,
		_w777_,
		_w852_
	);
	LUT3 #(
		.INIT('h0e)
	) name787 (
		_w769_,
		_w778_,
		_w852_,
		_w853_
	);
	LUT4 #(
		.INIT('h153f)
	) name788 (
		\a[2] ,
		\a[7] ,
		\a[20] ,
		\a[25] ,
		_w854_
	);
	LUT4 #(
		.INIT('h8000)
	) name789 (
		\a[2] ,
		\a[7] ,
		\a[20] ,
		\a[25] ,
		_w855_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name790 (
		\a[2] ,
		\a[7] ,
		\a[20] ,
		\a[25] ,
		_w856_
	);
	LUT2 #(
		.INIT('h6)
	) name791 (
		_w785_,
		_w856_,
		_w857_
	);
	LUT3 #(
		.INIT('h32)
	) name792 (
		_w809_,
		_w810_,
		_w811_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		\a[8] ,
		\a[19] ,
		_w859_
	);
	LUT4 #(
		.INIT('h153f)
	) name794 (
		\a[9] ,
		\a[10] ,
		\a[17] ,
		\a[18] ,
		_w860_
	);
	LUT4 #(
		.INIT('h8000)
	) name795 (
		\a[9] ,
		\a[10] ,
		\a[17] ,
		\a[18] ,
		_w861_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name796 (
		\a[9] ,
		\a[10] ,
		\a[17] ,
		\a[18] ,
		_w862_
	);
	LUT2 #(
		.INIT('h6)
	) name797 (
		_w859_,
		_w862_,
		_w863_
	);
	LUT3 #(
		.INIT('h96)
	) name798 (
		_w857_,
		_w858_,
		_w863_,
		_w864_
	);
	LUT4 #(
		.INIT('h004d)
	) name799 (
		_w769_,
		_w776_,
		_w777_,
		_w864_,
		_w865_
	);
	LUT4 #(
		.INIT('hb200)
	) name800 (
		_w769_,
		_w776_,
		_w777_,
		_w864_,
		_w866_
	);
	LUT3 #(
		.INIT('h23)
	) name801 (
		_w772_,
		_w773_,
		_w775_,
		_w867_
	);
	LUT3 #(
		.INIT('h8e)
	) name802 (
		_w807_,
		_w808_,
		_w813_,
		_w868_
	);
	LUT3 #(
		.INIT('h32)
	) name803 (
		_w792_,
		_w793_,
		_w798_,
		_w869_
	);
	LUT3 #(
		.INIT('h69)
	) name804 (
		_w867_,
		_w868_,
		_w869_,
		_w870_
	);
	LUT3 #(
		.INIT('h96)
	) name805 (
		_w853_,
		_w864_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h6)
	) name806 (
		_w851_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		_w822_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		_w822_,
		_w872_,
		_w874_
	);
	LUT2 #(
		.INIT('h6)
	) name809 (
		_w822_,
		_w872_,
		_w875_
	);
	LUT4 #(
		.INIT('h23dc)
	) name810 (
		_w765_,
		_w817_,
		_w821_,
		_w875_,
		_w876_
	);
	LUT3 #(
		.INIT('h15)
	) name811 (
		_w817_,
		_w822_,
		_w872_,
		_w877_
	);
	LUT3 #(
		.INIT('h32)
	) name812 (
		_w849_,
		_w850_,
		_w871_,
		_w878_
	);
	LUT4 #(
		.INIT('h8e00)
	) name813 (
		_w803_,
		_w806_,
		_w814_,
		_w829_,
		_w879_
	);
	LUT4 #(
		.INIT('h0027)
	) name814 (
		_w825_,
		_w845_,
		_w846_,
		_w879_,
		_w880_
	);
	LUT3 #(
		.INIT('h8e)
	) name815 (
		_w770_,
		_w830_,
		_w831_,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		\a[8] ,
		\a[20] ,
		_w882_
	);
	LUT4 #(
		.INIT('h153f)
	) name817 (
		\a[3] ,
		\a[4] ,
		\a[24] ,
		\a[25] ,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		\a[4] ,
		\a[25] ,
		_w884_
	);
	LUT4 #(
		.INIT('h8000)
	) name819 (
		\a[3] ,
		\a[4] ,
		\a[24] ,
		\a[25] ,
		_w885_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name820 (
		\a[3] ,
		\a[4] ,
		\a[24] ,
		\a[25] ,
		_w886_
	);
	LUT2 #(
		.INIT('h6)
	) name821 (
		_w882_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		\a[7] ,
		\a[21] ,
		_w888_
	);
	LUT4 #(
		.INIT('h153f)
	) name823 (
		\a[5] ,
		\a[6] ,
		\a[22] ,
		\a[23] ,
		_w889_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\a[6] ,
		\a[23] ,
		_w890_
	);
	LUT4 #(
		.INIT('h8000)
	) name825 (
		\a[5] ,
		\a[6] ,
		\a[22] ,
		\a[23] ,
		_w891_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name826 (
		\a[5] ,
		\a[6] ,
		\a[22] ,
		\a[23] ,
		_w892_
	);
	LUT2 #(
		.INIT('h6)
	) name827 (
		_w888_,
		_w892_,
		_w893_
	);
	LUT3 #(
		.INIT('h96)
	) name828 (
		_w881_,
		_w887_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		_w880_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w879_,
		_w894_,
		_w896_
	);
	LUT3 #(
		.INIT('h0e)
	) name831 (
		_w832_,
		_w841_,
		_w842_,
		_w897_
	);
	LUT3 #(
		.INIT('he8)
	) name832 (
		_w857_,
		_w858_,
		_w863_,
		_w898_
	);
	LUT3 #(
		.INIT('h80)
	) name833 (
		\a[1] ,
		\a[14] ,
		\a[26] ,
		_w899_
	);
	LUT4 #(
		.INIT('h8000)
	) name834 (
		\a[1] ,
		\a[13] ,
		\a[15] ,
		\a[27] ,
		_w900_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name835 (
		\a[1] ,
		\a[13] ,
		\a[15] ,
		\a[27] ,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name836 (
		_w899_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w899_,
		_w901_,
		_w903_
	);
	LUT2 #(
		.INIT('h6)
	) name838 (
		_w899_,
		_w901_,
		_w904_
	);
	LUT3 #(
		.INIT('h0d)
	) name839 (
		_w833_,
		_w834_,
		_w835_,
		_w905_
	);
	LUT2 #(
		.INIT('h6)
	) name840 (
		_w904_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('h69)
	) name841 (
		_w897_,
		_w898_,
		_w906_,
		_w907_
	);
	LUT3 #(
		.INIT('h70)
	) name842 (
		_w847_,
		_w896_,
		_w907_,
		_w908_
	);
	LUT4 #(
		.INIT('h2d00)
	) name843 (
		_w847_,
		_w879_,
		_w894_,
		_w907_,
		_w909_
	);
	LUT3 #(
		.INIT('h08)
	) name844 (
		_w847_,
		_w896_,
		_w907_,
		_w910_
	);
	LUT4 #(
		.INIT('h7dd7)
	) name845 (
		_w894_,
		_w897_,
		_w898_,
		_w906_,
		_w911_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w880_,
		_w911_,
		_w912_
	);
	LUT3 #(
		.INIT('h01)
	) name847 (
		_w909_,
		_w910_,
		_w912_,
		_w913_
	);
	LUT3 #(
		.INIT('hb2)
	) name848 (
		_w867_,
		_w868_,
		_w869_,
		_w914_
	);
	LUT3 #(
		.INIT('h32)
	) name849 (
		_w837_,
		_w838_,
		_w839_,
		_w915_
	);
	LUT3 #(
		.INIT('h0d)
	) name850 (
		_w859_,
		_w860_,
		_w861_,
		_w916_
	);
	LUT3 #(
		.INIT('h0d)
	) name851 (
		_w785_,
		_w854_,
		_w855_,
		_w917_
	);
	LUT3 #(
		.INIT('h69)
	) name852 (
		_w915_,
		_w916_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h8)
	) name853 (
		\a[2] ,
		\a[26] ,
		_w919_
	);
	LUT4 #(
		.INIT('h153f)
	) name854 (
		\a[9] ,
		\a[10] ,
		\a[18] ,
		\a[19] ,
		_w920_
	);
	LUT4 #(
		.INIT('h8000)
	) name855 (
		\a[9] ,
		\a[10] ,
		\a[18] ,
		\a[19] ,
		_w921_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name856 (
		\a[9] ,
		\a[10] ,
		\a[18] ,
		\a[19] ,
		_w922_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		\a[11] ,
		\a[17] ,
		_w923_
	);
	LUT4 #(
		.INIT('h153f)
	) name858 (
		\a[0] ,
		\a[12] ,
		\a[16] ,
		\a[28] ,
		_w924_
	);
	LUT4 #(
		.INIT('h8000)
	) name859 (
		\a[0] ,
		\a[12] ,
		\a[16] ,
		\a[28] ,
		_w925_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name860 (
		\a[0] ,
		\a[12] ,
		\a[16] ,
		\a[28] ,
		_w926_
	);
	LUT4 #(
		.INIT('h0660)
	) name861 (
		_w919_,
		_w922_,
		_w923_,
		_w926_,
		_w927_
	);
	LUT4 #(
		.INIT('h6996)
	) name862 (
		_w919_,
		_w922_,
		_w923_,
		_w926_,
		_w928_
	);
	LUT4 #(
		.INIT('h7100)
	) name863 (
		_w826_,
		_w827_,
		_w828_,
		_w928_,
		_w929_
	);
	LUT4 #(
		.INIT('h8e71)
	) name864 (
		_w826_,
		_w827_,
		_w828_,
		_w928_,
		_w930_
	);
	LUT3 #(
		.INIT('h6f)
	) name865 (
		_w914_,
		_w918_,
		_w930_,
		_w931_
	);
	LUT3 #(
		.INIT('h69)
	) name866 (
		_w914_,
		_w918_,
		_w930_,
		_w932_
	);
	LUT4 #(
		.INIT('hdc00)
	) name867 (
		_w865_,
		_w866_,
		_w870_,
		_w932_,
		_w933_
	);
	LUT4 #(
		.INIT('h17e8)
	) name868 (
		_w853_,
		_w864_,
		_w870_,
		_w932_,
		_w934_
	);
	LUT3 #(
		.INIT('hde)
	) name869 (
		_w878_,
		_w913_,
		_w934_,
		_w935_
	);
	LUT3 #(
		.INIT('hb7)
	) name870 (
		_w878_,
		_w913_,
		_w934_,
		_w936_
	);
	LUT3 #(
		.INIT('h96)
	) name871 (
		_w878_,
		_w913_,
		_w934_,
		_w937_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w874_,
		_w937_,
		_w938_
	);
	LUT4 #(
		.INIT('h4f00)
	) name873 (
		_w765_,
		_w821_,
		_w877_,
		_w938_,
		_w939_
	);
	LUT3 #(
		.INIT('h04)
	) name874 (
		_w873_,
		_w874_,
		_w937_,
		_w940_
	);
	LUT3 #(
		.INIT('h01)
	) name875 (
		_w817_,
		_w873_,
		_w937_,
		_w941_
	);
	LUT4 #(
		.INIT('h040f)
	) name876 (
		_w765_,
		_w821_,
		_w940_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h4)
	) name877 (
		_w939_,
		_w942_,
		_w943_
	);
	LUT3 #(
		.INIT('h40)
	) name878 (
		_w873_,
		_w874_,
		_w936_,
		_w944_
	);
	LUT3 #(
		.INIT('h10)
	) name879 (
		_w817_,
		_w873_,
		_w936_,
		_w945_
	);
	LUT4 #(
		.INIT('h040f)
	) name880 (
		_w765_,
		_w821_,
		_w944_,
		_w945_,
		_w946_
	);
	LUT3 #(
		.INIT('h2b)
	) name881 (
		_w915_,
		_w916_,
		_w917_,
		_w947_
	);
	LUT3 #(
		.INIT('h23)
	) name882 (
		_w902_,
		_w903_,
		_w905_,
		_w948_
	);
	LUT4 #(
		.INIT('h153f)
	) name883 (
		\a[13] ,
		\a[14] ,
		\a[15] ,
		\a[16] ,
		_w949_
	);
	LUT4 #(
		.INIT('h8000)
	) name884 (
		\a[13] ,
		\a[14] ,
		\a[15] ,
		\a[16] ,
		_w950_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name885 (
		\a[13] ,
		\a[14] ,
		\a[15] ,
		\a[16] ,
		_w951_
	);
	LUT2 #(
		.INIT('h6)
	) name886 (
		_w890_,
		_w951_,
		_w952_
	);
	LUT4 #(
		.INIT('h8e00)
	) name887 (
		_w899_,
		_w901_,
		_w905_,
		_w952_,
		_w953_
	);
	LUT4 #(
		.INIT('h0071)
	) name888 (
		_w899_,
		_w901_,
		_w905_,
		_w952_,
		_w954_
	);
	LUT4 #(
		.INIT('hdc23)
	) name889 (
		_w902_,
		_w903_,
		_w905_,
		_w952_,
		_w955_
	);
	LUT3 #(
		.INIT('h80)
	) name890 (
		\a[1] ,
		\a[15] ,
		\a[28] ,
		_w956_
	);
	LUT3 #(
		.INIT('h6c)
	) name891 (
		\a[1] ,
		\a[15] ,
		\a[28] ,
		_w957_
	);
	LUT3 #(
		.INIT('h0d)
	) name892 (
		_w888_,
		_w889_,
		_w891_,
		_w958_
	);
	LUT4 #(
		.INIT('h000d)
	) name893 (
		_w888_,
		_w889_,
		_w891_,
		_w957_,
		_w959_
	);
	LUT4 #(
		.INIT('hf200)
	) name894 (
		_w888_,
		_w889_,
		_w891_,
		_w957_,
		_w960_
	);
	LUT4 #(
		.INIT('h0df2)
	) name895 (
		_w888_,
		_w889_,
		_w891_,
		_w957_,
		_w961_
	);
	LUT3 #(
		.INIT('h0d)
	) name896 (
		_w882_,
		_w883_,
		_w885_,
		_w962_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		\a[12] ,
		\a[17] ,
		_w963_
	);
	LUT4 #(
		.INIT('h153f)
	) name898 (
		\a[3] ,
		\a[8] ,
		\a[21] ,
		\a[26] ,
		_w964_
	);
	LUT4 #(
		.INIT('h8000)
	) name899 (
		\a[3] ,
		\a[8] ,
		\a[21] ,
		\a[26] ,
		_w965_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name900 (
		\a[3] ,
		\a[8] ,
		\a[21] ,
		\a[26] ,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		\a[9] ,
		\a[20] ,
		_w967_
	);
	LUT4 #(
		.INIT('h153f)
	) name902 (
		\a[10] ,
		\a[11] ,
		\a[18] ,
		\a[19] ,
		_w968_
	);
	LUT4 #(
		.INIT('h8000)
	) name903 (
		\a[10] ,
		\a[11] ,
		\a[18] ,
		\a[19] ,
		_w969_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name904 (
		\a[10] ,
		\a[11] ,
		\a[18] ,
		\a[19] ,
		_w970_
	);
	LUT4 #(
		.INIT('h0660)
	) name905 (
		_w963_,
		_w966_,
		_w967_,
		_w970_,
		_w971_
	);
	LUT4 #(
		.INIT('h9009)
	) name906 (
		_w963_,
		_w966_,
		_w967_,
		_w970_,
		_w972_
	);
	LUT4 #(
		.INIT('h6996)
	) name907 (
		_w963_,
		_w966_,
		_w967_,
		_w970_,
		_w973_
	);
	LUT4 #(
		.INIT('h153f)
	) name908 (
		\a[5] ,
		\a[7] ,
		\a[22] ,
		\a[24] ,
		_w974_
	);
	LUT4 #(
		.INIT('h8000)
	) name909 (
		\a[5] ,
		\a[7] ,
		\a[22] ,
		\a[24] ,
		_w975_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name910 (
		\a[5] ,
		\a[7] ,
		\a[22] ,
		\a[24] ,
		_w976_
	);
	LUT2 #(
		.INIT('h6)
	) name911 (
		_w884_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('h0990)
	) name912 (
		_w961_,
		_w962_,
		_w973_,
		_w977_,
		_w978_
	);
	LUT4 #(
		.INIT('h6006)
	) name913 (
		_w961_,
		_w962_,
		_w973_,
		_w977_,
		_w979_
	);
	LUT4 #(
		.INIT('h9669)
	) name914 (
		_w961_,
		_w962_,
		_w973_,
		_w977_,
		_w980_
	);
	LUT3 #(
		.INIT('h96)
	) name915 (
		_w947_,
		_w955_,
		_w980_,
		_w981_
	);
	LUT4 #(
		.INIT('h00b2)
	) name916 (
		_w867_,
		_w868_,
		_w869_,
		_w918_,
		_w982_
	);
	LUT3 #(
		.INIT('h8e)
	) name917 (
		_w897_,
		_w898_,
		_w906_,
		_w983_
	);
	LUT3 #(
		.INIT('h32)
	) name918 (
		_w923_,
		_w924_,
		_w925_,
		_w984_
	);
	LUT3 #(
		.INIT('h0d)
	) name919 (
		_w919_,
		_w920_,
		_w921_,
		_w985_
	);
	LUT4 #(
		.INIT('h153f)
	) name920 (
		\a[0] ,
		\a[2] ,
		\a[27] ,
		\a[29] ,
		_w986_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		\a[2] ,
		\a[29] ,
		_w987_
	);
	LUT4 #(
		.INIT('h8000)
	) name922 (
		\a[0] ,
		\a[2] ,
		\a[27] ,
		\a[29] ,
		_w988_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name923 (
		\a[0] ,
		\a[2] ,
		\a[27] ,
		\a[29] ,
		_w989_
	);
	LUT2 #(
		.INIT('h6)
	) name924 (
		_w900_,
		_w989_,
		_w990_
	);
	LUT3 #(
		.INIT('h69)
	) name925 (
		_w984_,
		_w985_,
		_w990_,
		_w991_
	);
	LUT3 #(
		.INIT('he8)
	) name926 (
		_w881_,
		_w887_,
		_w893_,
		_w992_
	);
	LUT4 #(
		.INIT('hef1f)
	) name927 (
		_w927_,
		_w929_,
		_w991_,
		_w992_,
		_w993_
	);
	LUT4 #(
		.INIT('he11e)
	) name928 (
		_w927_,
		_w929_,
		_w991_,
		_w992_,
		_w994_
	);
	LUT4 #(
		.INIT('hd22d)
	) name929 (
		_w931_,
		_w982_,
		_w983_,
		_w994_,
		_w995_
	);
	LUT4 #(
		.INIT('he11e)
	) name930 (
		_w895_,
		_w908_,
		_w981_,
		_w995_,
		_w996_
	);
	LUT4 #(
		.INIT('he800)
	) name931 (
		_w824_,
		_w848_,
		_w871_,
		_w934_,
		_w997_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w933_,
		_w997_,
		_w998_
	);
	LUT3 #(
		.INIT('h7d)
	) name933 (
		_w935_,
		_w996_,
		_w998_,
		_w999_
	);
	LUT3 #(
		.INIT('hc8)
	) name934 (
		_w933_,
		_w996_,
		_w997_,
		_w1000_
	);
	LUT3 #(
		.INIT('h01)
	) name935 (
		_w933_,
		_w996_,
		_w997_,
		_w1001_
	);
	LUT3 #(
		.INIT('h36)
	) name936 (
		_w933_,
		_w996_,
		_w997_,
		_w1002_
	);
	LUT4 #(
		.INIT('hf380)
	) name937 (
		_w935_,
		_w946_,
		_w999_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		_w935_,
		_w1001_,
		_w1004_
	);
	LUT4 #(
		.INIT('h011f)
	) name939 (
		_w895_,
		_w909_,
		_w981_,
		_w995_,
		_w1005_
	);
	LUT4 #(
		.INIT('h022f)
	) name940 (
		_w931_,
		_w982_,
		_w983_,
		_w994_,
		_w1006_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		\a[5] ,
		\a[25] ,
		_w1007_
	);
	LUT4 #(
		.INIT('h153f)
	) name942 (
		\a[6] ,
		\a[7] ,
		\a[23] ,
		\a[24] ,
		_w1008_
	);
	LUT4 #(
		.INIT('h8000)
	) name943 (
		\a[6] ,
		\a[7] ,
		\a[23] ,
		\a[24] ,
		_w1009_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name944 (
		\a[6] ,
		\a[7] ,
		\a[23] ,
		\a[24] ,
		_w1010_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\a[3] ,
		\a[27] ,
		_w1011_
	);
	LUT4 #(
		.INIT('h153f)
	) name946 (
		\a[4] ,
		\a[8] ,
		\a[22] ,
		\a[26] ,
		_w1012_
	);
	LUT4 #(
		.INIT('h8000)
	) name947 (
		\a[4] ,
		\a[8] ,
		\a[22] ,
		\a[26] ,
		_w1013_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name948 (
		\a[4] ,
		\a[8] ,
		\a[22] ,
		\a[26] ,
		_w1014_
	);
	LUT4 #(
		.INIT('h0660)
	) name949 (
		_w1007_,
		_w1010_,
		_w1011_,
		_w1014_,
		_w1015_
	);
	LUT4 #(
		.INIT('h9009)
	) name950 (
		_w1007_,
		_w1010_,
		_w1011_,
		_w1014_,
		_w1016_
	);
	LUT4 #(
		.INIT('h6996)
	) name951 (
		_w1007_,
		_w1010_,
		_w1011_,
		_w1014_,
		_w1017_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		\a[10] ,
		\a[20] ,
		_w1018_
	);
	LUT4 #(
		.INIT('h153f)
	) name953 (
		\a[11] ,
		\a[12] ,
		\a[18] ,
		\a[19] ,
		_w1019_
	);
	LUT4 #(
		.INIT('h8000)
	) name954 (
		\a[11] ,
		\a[12] ,
		\a[18] ,
		\a[19] ,
		_w1020_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name955 (
		\a[11] ,
		\a[12] ,
		\a[18] ,
		\a[19] ,
		_w1021_
	);
	LUT2 #(
		.INIT('h6)
	) name956 (
		_w1018_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h6)
	) name957 (
		_w1017_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('h0017)
	) name958 (
		_w947_,
		_w948_,
		_w952_,
		_w1023_,
		_w1024_
	);
	LUT4 #(
		.INIT('he800)
	) name959 (
		_w947_,
		_w948_,
		_w952_,
		_w1023_,
		_w1025_
	);
	LUT4 #(
		.INIT('hf10e)
	) name960 (
		_w947_,
		_w953_,
		_w954_,
		_w1023_,
		_w1026_
	);
	LUT3 #(
		.INIT('he0)
	) name961 (
		_w927_,
		_w929_,
		_w992_,
		_w1027_
	);
	LUT4 #(
		.INIT('h011f)
	) name962 (
		_w927_,
		_w929_,
		_w991_,
		_w992_,
		_w1028_
	);
	LUT2 #(
		.INIT('h6)
	) name963 (
		_w1026_,
		_w1028_,
		_w1029_
	);
	LUT4 #(
		.INIT('h8000)
	) name964 (
		\a[1] ,
		\a[14] ,
		\a[16] ,
		\a[29] ,
		_w1030_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name965 (
		\a[1] ,
		\a[14] ,
		\a[16] ,
		\a[29] ,
		_w1031_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		\a[0] ,
		\a[30] ,
		_w1032_
	);
	LUT3 #(
		.INIT('h96)
	) name967 (
		_w956_,
		_w1031_,
		_w1032_,
		_w1033_
	);
	LUT4 #(
		.INIT('h00d4)
	) name968 (
		_w957_,
		_w958_,
		_w962_,
		_w1033_,
		_w1034_
	);
	LUT4 #(
		.INIT('h2b00)
	) name969 (
		_w957_,
		_w958_,
		_w962_,
		_w1033_,
		_w1035_
	);
	LUT4 #(
		.INIT('hba45)
	) name970 (
		_w959_,
		_w960_,
		_w962_,
		_w1033_,
		_w1036_
	);
	LUT3 #(
		.INIT('hb2)
	) name971 (
		_w984_,
		_w985_,
		_w990_,
		_w1037_
	);
	LUT2 #(
		.INIT('h6)
	) name972 (
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('h00f6)
	) name973 (
		_w947_,
		_w955_,
		_w978_,
		_w979_,
		_w1039_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT3 #(
		.INIT('h32)
	) name975 (
		_w971_,
		_w972_,
		_w977_,
		_w1041_
	);
	LUT3 #(
		.INIT('h32)
	) name976 (
		_w890_,
		_w949_,
		_w950_,
		_w1042_
	);
	LUT3 #(
		.INIT('h0d)
	) name977 (
		_w884_,
		_w974_,
		_w975_,
		_w1043_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		\a[13] ,
		\a[17] ,
		_w1044_
	);
	LUT4 #(
		.INIT('h153f)
	) name979 (
		\a[2] ,
		\a[9] ,
		\a[21] ,
		\a[28] ,
		_w1045_
	);
	LUT4 #(
		.INIT('h8000)
	) name980 (
		\a[2] ,
		\a[9] ,
		\a[21] ,
		\a[28] ,
		_w1046_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name981 (
		\a[2] ,
		\a[9] ,
		\a[21] ,
		\a[28] ,
		_w1047_
	);
	LUT2 #(
		.INIT('h6)
	) name982 (
		_w1044_,
		_w1047_,
		_w1048_
	);
	LUT3 #(
		.INIT('h69)
	) name983 (
		_w1042_,
		_w1043_,
		_w1048_,
		_w1049_
	);
	LUT3 #(
		.INIT('h0d)
	) name984 (
		_w967_,
		_w968_,
		_w969_,
		_w1050_
	);
	LUT3 #(
		.INIT('h0d)
	) name985 (
		_w963_,
		_w964_,
		_w965_,
		_w1051_
	);
	LUT3 #(
		.INIT('h0d)
	) name986 (
		_w900_,
		_w986_,
		_w988_,
		_w1052_
	);
	LUT3 #(
		.INIT('h96)
	) name987 (
		_w1050_,
		_w1051_,
		_w1052_,
		_w1053_
	);
	LUT3 #(
		.INIT('h69)
	) name988 (
		_w1041_,
		_w1049_,
		_w1053_,
		_w1054_
	);
	LUT3 #(
		.INIT('h96)
	) name989 (
		_w1038_,
		_w1039_,
		_w1054_,
		_w1055_
	);
	LUT3 #(
		.INIT('h96)
	) name990 (
		_w1006_,
		_w1029_,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		_w1005_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h9)
	) name992 (
		_w1005_,
		_w1056_,
		_w1058_
	);
	LUT4 #(
		.INIT('h13ec)
	) name993 (
		_w946_,
		_w1000_,
		_w1004_,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w1000_,
		_w1057_,
		_w1060_
	);
	LUT3 #(
		.INIT('h8e)
	) name995 (
		_w1006_,
		_w1029_,
		_w1055_,
		_w1061_
	);
	LUT3 #(
		.INIT('h07)
	) name996 (
		_w1038_,
		_w1039_,
		_w1054_,
		_w1062_
	);
	LUT3 #(
		.INIT('h8e)
	) name997 (
		_w1041_,
		_w1049_,
		_w1053_,
		_w1063_
	);
	LUT3 #(
		.INIT('he8)
	) name998 (
		_w956_,
		_w1031_,
		_w1032_,
		_w1064_
	);
	LUT2 #(
		.INIT('h8)
	) name999 (
		\a[11] ,
		\a[20] ,
		_w1065_
	);
	LUT4 #(
		.INIT('h153f)
	) name1000 (
		\a[12] ,
		\a[13] ,
		\a[18] ,
		\a[19] ,
		_w1066_
	);
	LUT4 #(
		.INIT('h8000)
	) name1001 (
		\a[12] ,
		\a[13] ,
		\a[18] ,
		\a[19] ,
		_w1067_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1002 (
		\a[12] ,
		\a[13] ,
		\a[18] ,
		\a[19] ,
		_w1068_
	);
	LUT2 #(
		.INIT('h6)
	) name1003 (
		_w1065_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name1004 (
		\a[10] ,
		\a[21] ,
		_w1070_
	);
	LUT4 #(
		.INIT('h153f)
	) name1005 (
		\a[0] ,
		\a[9] ,
		\a[22] ,
		\a[31] ,
		_w1071_
	);
	LUT4 #(
		.INIT('h8000)
	) name1006 (
		\a[0] ,
		\a[9] ,
		\a[22] ,
		\a[31] ,
		_w1072_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1007 (
		\a[0] ,
		\a[9] ,
		\a[22] ,
		\a[31] ,
		_w1073_
	);
	LUT2 #(
		.INIT('h6)
	) name1008 (
		_w1070_,
		_w1073_,
		_w1074_
	);
	LUT3 #(
		.INIT('h96)
	) name1009 (
		_w1064_,
		_w1069_,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		\a[8] ,
		\a[23] ,
		_w1076_
	);
	LUT4 #(
		.INIT('h153f)
	) name1011 (
		\a[5] ,
		\a[7] ,
		\a[24] ,
		\a[26] ,
		_w1077_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		\a[7] ,
		\a[26] ,
		_w1078_
	);
	LUT4 #(
		.INIT('h8000)
	) name1013 (
		\a[5] ,
		\a[7] ,
		\a[24] ,
		\a[26] ,
		_w1079_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1014 (
		\a[5] ,
		\a[7] ,
		\a[24] ,
		\a[26] ,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		\a[6] ,
		\a[25] ,
		_w1081_
	);
	LUT4 #(
		.INIT('h153f)
	) name1016 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w1082_
	);
	LUT4 #(
		.INIT('h8000)
	) name1017 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w1083_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1018 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w1084_
	);
	LUT4 #(
		.INIT('h0660)
	) name1019 (
		_w1076_,
		_w1080_,
		_w1081_,
		_w1084_,
		_w1085_
	);
	LUT4 #(
		.INIT('h9009)
	) name1020 (
		_w1076_,
		_w1080_,
		_w1081_,
		_w1084_,
		_w1086_
	);
	LUT4 #(
		.INIT('h6996)
	) name1021 (
		_w1076_,
		_w1080_,
		_w1081_,
		_w1084_,
		_w1087_
	);
	LUT4 #(
		.INIT('h153f)
	) name1022 (
		\a[3] ,
		\a[4] ,
		\a[27] ,
		\a[28] ,
		_w1088_
	);
	LUT4 #(
		.INIT('h8000)
	) name1023 (
		\a[3] ,
		\a[4] ,
		\a[27] ,
		\a[28] ,
		_w1089_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1024 (
		\a[3] ,
		\a[4] ,
		\a[27] ,
		\a[28] ,
		_w1090_
	);
	LUT2 #(
		.INIT('h6)
	) name1025 (
		_w987_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h6)
	) name1026 (
		_w1087_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		_w1075_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		_w1075_,
		_w1092_,
		_w1094_
	);
	LUT2 #(
		.INIT('h6)
	) name1029 (
		_w1075_,
		_w1092_,
		_w1095_
	);
	LUT2 #(
		.INIT('h6)
	) name1030 (
		_w1063_,
		_w1095_,
		_w1096_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name1031 (
		_w1038_,
		_w1039_,
		_w1063_,
		_w1095_,
		_w1097_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		_w1062_,
		_w1097_,
		_w1098_
	);
	LUT3 #(
		.INIT('he8)
	) name1033 (
		_w1038_,
		_w1039_,
		_w1054_,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w1096_,
		_w1099_,
		_w1100_
	);
	LUT3 #(
		.INIT('he1)
	) name1035 (
		_w1040_,
		_w1062_,
		_w1096_,
		_w1101_
	);
	LUT3 #(
		.INIT('h02)
	) name1036 (
		_w993_,
		_w1025_,
		_w1027_,
		_w1102_
	);
	LUT4 #(
		.INIT('h3331)
	) name1037 (
		_w993_,
		_w1024_,
		_w1025_,
		_w1027_,
		_w1103_
	);
	LUT3 #(
		.INIT('h32)
	) name1038 (
		_w1044_,
		_w1045_,
		_w1046_,
		_w1104_
	);
	LUT3 #(
		.INIT('h32)
	) name1039 (
		_w1011_,
		_w1012_,
		_w1013_,
		_w1105_
	);
	LUT3 #(
		.INIT('h0d)
	) name1040 (
		_w1018_,
		_w1019_,
		_w1020_,
		_w1106_
	);
	LUT3 #(
		.INIT('h96)
	) name1041 (
		_w1104_,
		_w1105_,
		_w1106_,
		_w1107_
	);
	LUT3 #(
		.INIT('h32)
	) name1042 (
		_w1015_,
		_w1016_,
		_w1022_,
		_w1108_
	);
	LUT2 #(
		.INIT('h2)
	) name1043 (
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name1044 (
		_w1107_,
		_w1108_,
		_w1110_
	);
	LUT2 #(
		.INIT('h9)
	) name1045 (
		_w1107_,
		_w1108_,
		_w1111_
	);
	LUT3 #(
		.INIT('h54)
	) name1046 (
		_w1034_,
		_w1035_,
		_w1037_,
		_w1112_
	);
	LUT2 #(
		.INIT('h8)
	) name1047 (
		_w1111_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h6)
	) name1048 (
		_w1111_,
		_w1112_,
		_w1114_
	);
	LUT3 #(
		.INIT('h17)
	) name1049 (
		_w1050_,
		_w1051_,
		_w1052_,
		_w1115_
	);
	LUT3 #(
		.INIT('hb2)
	) name1050 (
		_w1042_,
		_w1043_,
		_w1048_,
		_w1116_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		\a[1] ,
		\a[30] ,
		_w1117_
	);
	LUT3 #(
		.INIT('h2d)
	) name1052 (
		\a[16] ,
		_w1030_,
		_w1117_,
		_w1118_
	);
	LUT3 #(
		.INIT('h0d)
	) name1053 (
		_w1007_,
		_w1008_,
		_w1009_,
		_w1119_
	);
	LUT2 #(
		.INIT('h6)
	) name1054 (
		_w1118_,
		_w1119_,
		_w1120_
	);
	LUT3 #(
		.INIT('h96)
	) name1055 (
		_w1115_,
		_w1116_,
		_w1120_,
		_w1121_
	);
	LUT3 #(
		.INIT('h09)
	) name1056 (
		_w1111_,
		_w1112_,
		_w1121_,
		_w1122_
	);
	LUT3 #(
		.INIT('h90)
	) name1057 (
		_w1111_,
		_w1112_,
		_w1121_,
		_w1123_
	);
	LUT3 #(
		.INIT('h27)
	) name1058 (
		_w1103_,
		_w1122_,
		_w1123_,
		_w1124_
	);
	LUT4 #(
		.INIT('h10e0)
	) name1059 (
		_w1024_,
		_w1102_,
		_w1114_,
		_w1121_,
		_w1125_
	);
	LUT3 #(
		.INIT('h59)
	) name1060 (
		_w1101_,
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h4)
	) name1061 (
		_w1061_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h2)
	) name1062 (
		_w1061_,
		_w1126_,
		_w1128_
	);
	LUT4 #(
		.INIT('h2dd2)
	) name1063 (
		_w1005_,
		_w1056_,
		_w1061_,
		_w1126_,
		_w1129_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1064 (
		_w946_,
		_w1004_,
		_w1060_,
		_w1129_,
		_w1130_
	);
	LUT4 #(
		.INIT('hf00f)
	) name1065 (
		_w1005_,
		_w1056_,
		_w1061_,
		_w1126_,
		_w1131_
	);
	LUT4 #(
		.INIT('h7000)
	) name1066 (
		_w946_,
		_w1004_,
		_w1060_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('he)
	) name1067 (
		_w1130_,
		_w1132_,
		_w1133_
	);
	LUT4 #(
		.INIT('h0070)
	) name1068 (
		_w946_,
		_w1004_,
		_w1060_,
		_w1127_,
		_w1134_
	);
	LUT4 #(
		.INIT('h2022)
	) name1069 (
		_w1005_,
		_w1056_,
		_w1061_,
		_w1126_,
		_w1135_
	);
	LUT4 #(
		.INIT('h3323)
	) name1070 (
		_w1098_,
		_w1100_,
		_w1124_,
		_w1125_,
		_w1136_
	);
	LUT2 #(
		.INIT('h4)
	) name1071 (
		_w1024_,
		_w1121_,
		_w1137_
	);
	LUT2 #(
		.INIT('h4)
	) name1072 (
		_w1102_,
		_w1137_,
		_w1138_
	);
	LUT3 #(
		.INIT('h23)
	) name1073 (
		_w1102_,
		_w1113_,
		_w1137_,
		_w1139_
	);
	LUT3 #(
		.INIT('he0)
	) name1074 (
		_w1111_,
		_w1112_,
		_w1121_,
		_w1140_
	);
	LUT3 #(
		.INIT('h54)
	) name1075 (
		_w1024_,
		_w1111_,
		_w1112_,
		_w1141_
	);
	LUT3 #(
		.INIT('h23)
	) name1076 (
		_w1102_,
		_w1140_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h4)
	) name1077 (
		\a[30] ,
		_w1030_,
		_w1143_
	);
	LUT4 #(
		.INIT('h5093)
	) name1078 (
		\a[1] ,
		\a[16] ,
		\a[30] ,
		_w1030_,
		_w1144_
	);
	LUT2 #(
		.INIT('h8)
	) name1079 (
		\a[9] ,
		\a[23] ,
		_w1145_
	);
	LUT4 #(
		.INIT('h153f)
	) name1080 (
		\a[4] ,
		\a[5] ,
		\a[27] ,
		\a[28] ,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name1081 (
		\a[5] ,
		\a[28] ,
		_w1147_
	);
	LUT4 #(
		.INIT('h8000)
	) name1082 (
		\a[4] ,
		\a[5] ,
		\a[27] ,
		\a[28] ,
		_w1148_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1083 (
		\a[4] ,
		\a[5] ,
		\a[27] ,
		\a[28] ,
		_w1149_
	);
	LUT2 #(
		.INIT('h8)
	) name1084 (
		\a[8] ,
		\a[24] ,
		_w1150_
	);
	LUT4 #(
		.INIT('h153f)
	) name1085 (
		\a[6] ,
		\a[7] ,
		\a[25] ,
		\a[26] ,
		_w1151_
	);
	LUT4 #(
		.INIT('h8000)
	) name1086 (
		\a[6] ,
		\a[7] ,
		\a[25] ,
		\a[26] ,
		_w1152_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1087 (
		\a[6] ,
		\a[7] ,
		\a[25] ,
		\a[26] ,
		_w1153_
	);
	LUT4 #(
		.INIT('h0660)
	) name1088 (
		_w1145_,
		_w1149_,
		_w1150_,
		_w1153_,
		_w1154_
	);
	LUT4 #(
		.INIT('h9009)
	) name1089 (
		_w1145_,
		_w1149_,
		_w1150_,
		_w1153_,
		_w1155_
	);
	LUT4 #(
		.INIT('h6996)
	) name1090 (
		_w1145_,
		_w1149_,
		_w1150_,
		_w1153_,
		_w1156_
	);
	LUT4 #(
		.INIT('hf20d)
	) name1091 (
		_w1119_,
		_w1143_,
		_w1144_,
		_w1156_,
		_w1157_
	);
	LUT3 #(
		.INIT('h80)
	) name1092 (
		\a[1] ,
		\a[16] ,
		\a[30] ,
		_w1158_
	);
	LUT4 #(
		.INIT('h153f)
	) name1093 (
		\a[0] ,
		\a[2] ,
		\a[30] ,
		\a[32] ,
		_w1159_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		\a[2] ,
		\a[32] ,
		_w1160_
	);
	LUT4 #(
		.INIT('h8000)
	) name1095 (
		\a[0] ,
		\a[2] ,
		\a[30] ,
		\a[32] ,
		_w1161_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1096 (
		\a[0] ,
		\a[2] ,
		\a[30] ,
		\a[32] ,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name1097 (
		\a[11] ,
		\a[21] ,
		_w1163_
	);
	LUT4 #(
		.INIT('h153f)
	) name1098 (
		\a[12] ,
		\a[13] ,
		\a[19] ,
		\a[20] ,
		_w1164_
	);
	LUT4 #(
		.INIT('h8000)
	) name1099 (
		\a[12] ,
		\a[13] ,
		\a[19] ,
		\a[20] ,
		_w1165_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1100 (
		\a[12] ,
		\a[13] ,
		\a[19] ,
		\a[20] ,
		_w1166_
	);
	LUT4 #(
		.INIT('h0660)
	) name1101 (
		_w1158_,
		_w1162_,
		_w1163_,
		_w1166_,
		_w1167_
	);
	LUT4 #(
		.INIT('h9009)
	) name1102 (
		_w1158_,
		_w1162_,
		_w1163_,
		_w1166_,
		_w1168_
	);
	LUT4 #(
		.INIT('h6996)
	) name1103 (
		_w1158_,
		_w1162_,
		_w1163_,
		_w1166_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name1104 (
		\a[14] ,
		\a[18] ,
		_w1170_
	);
	LUT4 #(
		.INIT('h153f)
	) name1105 (
		\a[3] ,
		\a[10] ,
		\a[22] ,
		\a[29] ,
		_w1171_
	);
	LUT4 #(
		.INIT('h8000)
	) name1106 (
		\a[3] ,
		\a[10] ,
		\a[22] ,
		\a[29] ,
		_w1172_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1107 (
		\a[3] ,
		\a[10] ,
		\a[22] ,
		\a[29] ,
		_w1173_
	);
	LUT2 #(
		.INIT('h6)
	) name1108 (
		_w1170_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h6)
	) name1109 (
		_w1169_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name1110 (
		_w1157_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h6)
	) name1111 (
		_w1157_,
		_w1175_,
		_w1177_
	);
	LUT4 #(
		.INIT('h23dc)
	) name1112 (
		_w1109_,
		_w1110_,
		_w1112_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('hae00)
	) name1113 (
		_w1138_,
		_w1139_,
		_w1142_,
		_w1178_,
		_w1179_
	);
	LUT3 #(
		.INIT('h0b)
	) name1114 (
		_w1102_,
		_w1137_,
		_w1178_,
		_w1180_
	);
	LUT3 #(
		.INIT('hd0)
	) name1115 (
		_w1139_,
		_w1142_,
		_w1180_,
		_w1181_
	);
	LUT3 #(
		.INIT('h31)
	) name1116 (
		_w1063_,
		_w1093_,
		_w1094_,
		_w1182_
	);
	LUT3 #(
		.INIT('he8)
	) name1117 (
		_w1064_,
		_w1069_,
		_w1074_,
		_w1183_
	);
	LUT3 #(
		.INIT('h8e)
	) name1118 (
		_w1104_,
		_w1105_,
		_w1106_,
		_w1184_
	);
	LUT3 #(
		.INIT('h32)
	) name1119 (
		_w1085_,
		_w1086_,
		_w1091_,
		_w1185_
	);
	LUT3 #(
		.INIT('h96)
	) name1120 (
		_w1183_,
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT3 #(
		.INIT('he8)
	) name1121 (
		_w1115_,
		_w1116_,
		_w1120_,
		_w1187_
	);
	LUT3 #(
		.INIT('h0d)
	) name1122 (
		_w1065_,
		_w1066_,
		_w1067_,
		_w1188_
	);
	LUT3 #(
		.INIT('h0d)
	) name1123 (
		_w1070_,
		_w1071_,
		_w1072_,
		_w1189_
	);
	LUT3 #(
		.INIT('h0d)
	) name1124 (
		_w987_,
		_w1088_,
		_w1089_,
		_w1190_
	);
	LUT3 #(
		.INIT('h96)
	) name1125 (
		_w1188_,
		_w1189_,
		_w1190_,
		_w1191_
	);
	LUT4 #(
		.INIT('h8000)
	) name1126 (
		\a[1] ,
		\a[15] ,
		\a[17] ,
		\a[31] ,
		_w1192_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1127 (
		\a[1] ,
		\a[15] ,
		\a[17] ,
		\a[31] ,
		_w1193_
	);
	LUT4 #(
		.INIT('h000d)
	) name1128 (
		_w1081_,
		_w1082_,
		_w1083_,
		_w1193_,
		_w1194_
	);
	LUT4 #(
		.INIT('hf200)
	) name1129 (
		_w1081_,
		_w1082_,
		_w1083_,
		_w1193_,
		_w1195_
	);
	LUT4 #(
		.INIT('h0df2)
	) name1130 (
		_w1081_,
		_w1082_,
		_w1083_,
		_w1193_,
		_w1196_
	);
	LUT3 #(
		.INIT('h0d)
	) name1131 (
		_w1076_,
		_w1077_,
		_w1079_,
		_w1197_
	);
	LUT2 #(
		.INIT('h6)
	) name1132 (
		_w1196_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h1)
	) name1133 (
		_w1191_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name1134 (
		_w1191_,
		_w1198_,
		_w1200_
	);
	LUT2 #(
		.INIT('h6)
	) name1135 (
		_w1191_,
		_w1198_,
		_w1201_
	);
	LUT4 #(
		.INIT('h9669)
	) name1136 (
		_w1182_,
		_w1186_,
		_w1187_,
		_w1201_,
		_w1202_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1137 (
		_w1139_,
		_w1142_,
		_w1180_,
		_w1202_,
		_w1203_
	);
	LUT4 #(
		.INIT('h0154)
	) name1138 (
		_w1136_,
		_w1179_,
		_w1181_,
		_w1202_,
		_w1204_
	);
	LUT4 #(
		.INIT('ha802)
	) name1139 (
		_w1136_,
		_w1179_,
		_w1181_,
		_w1202_,
		_w1205_
	);
	LUT4 #(
		.INIT('h0001)
	) name1140 (
		_w1128_,
		_w1135_,
		_w1204_,
		_w1205_,
		_w1206_
	);
	LUT4 #(
		.INIT('h56a9)
	) name1141 (
		_w1136_,
		_w1179_,
		_w1181_,
		_w1202_,
		_w1207_
	);
	LUT4 #(
		.INIT('hdf0d)
	) name1142 (
		_w1005_,
		_w1056_,
		_w1061_,
		_w1126_,
		_w1208_
	);
	LUT4 #(
		.INIT('hb1b0)
	) name1143 (
		_w1134_,
		_w1206_,
		_w1207_,
		_w1208_,
		_w1209_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name1144 (
		_w1107_,
		_w1108_,
		_w1157_,
		_w1175_,
		_w1210_
	);
	LUT4 #(
		.INIT('h080f)
	) name1145 (
		_w1111_,
		_w1112_,
		_w1176_,
		_w1210_,
		_w1211_
	);
	LUT3 #(
		.INIT('h17)
	) name1146 (
		_w1188_,
		_w1189_,
		_w1190_,
		_w1212_
	);
	LUT3 #(
		.INIT('h32)
	) name1147 (
		_w1167_,
		_w1168_,
		_w1174_,
		_w1213_
	);
	LUT4 #(
		.INIT('h00f2)
	) name1148 (
		_w1119_,
		_w1143_,
		_w1144_,
		_w1154_,
		_w1214_
	);
	LUT4 #(
		.INIT('h3c69)
	) name1149 (
		_w1155_,
		_w1212_,
		_w1213_,
		_w1214_,
		_w1215_
	);
	LUT3 #(
		.INIT('h0d)
	) name1150 (
		_w1163_,
		_w1164_,
		_w1165_,
		_w1216_
	);
	LUT3 #(
		.INIT('h0d)
	) name1151 (
		_w1158_,
		_w1159_,
		_w1161_,
		_w1217_
	);
	LUT3 #(
		.INIT('h32)
	) name1152 (
		_w1170_,
		_w1171_,
		_w1172_,
		_w1218_
	);
	LUT3 #(
		.INIT('h96)
	) name1153 (
		_w1216_,
		_w1217_,
		_w1218_,
		_w1219_
	);
	LUT3 #(
		.INIT('h0d)
	) name1154 (
		_w1150_,
		_w1151_,
		_w1152_,
		_w1220_
	);
	LUT3 #(
		.INIT('h0d)
	) name1155 (
		_w1145_,
		_w1146_,
		_w1148_,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		\a[2] ,
		\a[31] ,
		_w1222_
	);
	LUT4 #(
		.INIT('h153f)
	) name1157 (
		\a[0] ,
		\a[11] ,
		\a[22] ,
		\a[33] ,
		_w1223_
	);
	LUT4 #(
		.INIT('h8000)
	) name1158 (
		\a[0] ,
		\a[11] ,
		\a[22] ,
		\a[33] ,
		_w1224_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1159 (
		\a[0] ,
		\a[11] ,
		\a[22] ,
		\a[33] ,
		_w1225_
	);
	LUT2 #(
		.INIT('h6)
	) name1160 (
		_w1222_,
		_w1225_,
		_w1226_
	);
	LUT3 #(
		.INIT('h69)
	) name1161 (
		_w1220_,
		_w1221_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name1162 (
		\a[6] ,
		\a[28] ,
		_w1228_
	);
	LUT4 #(
		.INIT('h8000)
	) name1163 (
		\a[5] ,
		\a[6] ,
		\a[27] ,
		\a[28] ,
		_w1229_
	);
	LUT4 #(
		.INIT('h8000)
	) name1164 (
		\a[5] ,
		\a[8] ,
		\a[25] ,
		\a[28] ,
		_w1230_
	);
	LUT4 #(
		.INIT('h8000)
	) name1165 (
		\a[6] ,
		\a[8] ,
		\a[25] ,
		\a[27] ,
		_w1231_
	);
	LUT3 #(
		.INIT('h0e)
	) name1166 (
		_w1229_,
		_w1230_,
		_w1231_,
		_w1232_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1167 (
		\a[6] ,
		\a[8] ,
		\a[25] ,
		\a[27] ,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w1147_,
		_w1233_,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name1169 (
		\a[3] ,
		\a[30] ,
		_w1235_
	);
	LUT4 #(
		.INIT('h153f)
	) name1170 (
		\a[4] ,
		\a[9] ,
		\a[24] ,
		\a[29] ,
		_w1236_
	);
	LUT4 #(
		.INIT('h8000)
	) name1171 (
		\a[4] ,
		\a[9] ,
		\a[24] ,
		\a[29] ,
		_w1237_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1172 (
		\a[4] ,
		\a[9] ,
		\a[24] ,
		\a[29] ,
		_w1238_
	);
	LUT2 #(
		.INIT('h6)
	) name1173 (
		_w1235_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('h153f)
	) name1174 (
		\a[15] ,
		\a[16] ,
		\a[17] ,
		\a[18] ,
		_w1240_
	);
	LUT4 #(
		.INIT('h8000)
	) name1175 (
		\a[15] ,
		\a[16] ,
		\a[17] ,
		\a[18] ,
		_w1241_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1176 (
		\a[15] ,
		\a[16] ,
		\a[17] ,
		\a[18] ,
		_w1242_
	);
	LUT2 #(
		.INIT('h6)
	) name1177 (
		_w1078_,
		_w1242_,
		_w1243_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name1178 (
		_w1232_,
		_w1234_,
		_w1239_,
		_w1243_,
		_w1244_
	);
	LUT3 #(
		.INIT('h69)
	) name1179 (
		_w1219_,
		_w1227_,
		_w1244_,
		_w1245_
	);
	LUT3 #(
		.INIT('h96)
	) name1180 (
		_w1211_,
		_w1215_,
		_w1245_,
		_w1246_
	);
	LUT3 #(
		.INIT('h45)
	) name1181 (
		_w1194_,
		_w1195_,
		_w1197_,
		_w1247_
	);
	LUT2 #(
		.INIT('h8)
	) name1182 (
		\a[10] ,
		\a[23] ,
		_w1248_
	);
	LUT3 #(
		.INIT('h80)
	) name1183 (
		\a[1] ,
		\a[17] ,
		\a[32] ,
		_w1249_
	);
	LUT3 #(
		.INIT('h6c)
	) name1184 (
		\a[1] ,
		\a[17] ,
		\a[32] ,
		_w1250_
	);
	LUT3 #(
		.INIT('h96)
	) name1185 (
		_w1192_,
		_w1248_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h8)
	) name1186 (
		\a[12] ,
		\a[21] ,
		_w1252_
	);
	LUT4 #(
		.INIT('h153f)
	) name1187 (
		\a[13] ,
		\a[14] ,
		\a[19] ,
		\a[20] ,
		_w1253_
	);
	LUT4 #(
		.INIT('h8000)
	) name1188 (
		\a[13] ,
		\a[14] ,
		\a[19] ,
		\a[20] ,
		_w1254_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1189 (
		\a[13] ,
		\a[14] ,
		\a[19] ,
		\a[20] ,
		_w1255_
	);
	LUT2 #(
		.INIT('h6)
	) name1190 (
		_w1252_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		_w1251_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		_w1251_,
		_w1256_,
		_w1258_
	);
	LUT2 #(
		.INIT('h6)
	) name1193 (
		_w1251_,
		_w1256_,
		_w1259_
	);
	LUT2 #(
		.INIT('h6)
	) name1194 (
		_w1247_,
		_w1259_,
		_w1260_
	);
	LUT3 #(
		.INIT('he8)
	) name1195 (
		_w1183_,
		_w1184_,
		_w1185_,
		_w1261_
	);
	LUT2 #(
		.INIT('h1)
	) name1196 (
		_w1260_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		_w1260_,
		_w1261_,
		_w1263_
	);
	LUT2 #(
		.INIT('h6)
	) name1198 (
		_w1260_,
		_w1261_,
		_w1264_
	);
	LUT3 #(
		.INIT('h31)
	) name1199 (
		_w1187_,
		_w1199_,
		_w1200_,
		_w1265_
	);
	LUT2 #(
		.INIT('h6)
	) name1200 (
		_w1264_,
		_w1265_,
		_w1266_
	);
	LUT4 #(
		.INIT('hb22b)
	) name1201 (
		_w1182_,
		_w1186_,
		_w1187_,
		_w1201_,
		_w1267_
	);
	LUT3 #(
		.INIT('h96)
	) name1202 (
		_w1246_,
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT3 #(
		.INIT('h01)
	) name1203 (
		_w1179_,
		_w1203_,
		_w1268_,
		_w1269_
	);
	LUT3 #(
		.INIT('he0)
	) name1204 (
		_w1179_,
		_w1203_,
		_w1268_,
		_w1270_
	);
	LUT3 #(
		.INIT('h1e)
	) name1205 (
		_w1179_,
		_w1203_,
		_w1268_,
		_w1271_
	);
	LUT2 #(
		.INIT('h4)
	) name1206 (
		_w1204_,
		_w1208_,
		_w1272_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name1207 (
		_w1134_,
		_w1205_,
		_w1271_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name1208 (
		_w1205_,
		_w1270_,
		_w1274_
	);
	LUT3 #(
		.INIT('h2b)
	) name1209 (
		_w1246_,
		_w1266_,
		_w1267_,
		_w1275_
	);
	LUT3 #(
		.INIT('h32)
	) name1210 (
		_w1235_,
		_w1236_,
		_w1237_,
		_w1276_
	);
	LUT3 #(
		.INIT('h0d)
	) name1211 (
		_w1222_,
		_w1223_,
		_w1224_,
		_w1277_
	);
	LUT3 #(
		.INIT('h01)
	) name1212 (
		_w1229_,
		_w1230_,
		_w1231_,
		_w1278_
	);
	LUT3 #(
		.INIT('h69)
	) name1213 (
		_w1276_,
		_w1277_,
		_w1278_,
		_w1279_
	);
	LUT4 #(
		.INIT('hf110)
	) name1214 (
		_w1232_,
		_w1234_,
		_w1239_,
		_w1243_,
		_w1280_
	);
	LUT4 #(
		.INIT('h8000)
	) name1215 (
		\a[1] ,
		\a[16] ,
		\a[18] ,
		\a[33] ,
		_w1281_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1216 (
		\a[1] ,
		\a[16] ,
		\a[18] ,
		\a[33] ,
		_w1282_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		_w1249_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1249_,
		_w1282_,
		_w1284_
	);
	LUT2 #(
		.INIT('h6)
	) name1219 (
		_w1249_,
		_w1282_,
		_w1285_
	);
	LUT3 #(
		.INIT('h0d)
	) name1220 (
		_w1078_,
		_w1240_,
		_w1241_,
		_w1286_
	);
	LUT2 #(
		.INIT('h6)
	) name1221 (
		_w1285_,
		_w1286_,
		_w1287_
	);
	LUT3 #(
		.INIT('h96)
	) name1222 (
		_w1279_,
		_w1280_,
		_w1287_,
		_w1288_
	);
	LUT3 #(
		.INIT('he8)
	) name1223 (
		_w1192_,
		_w1248_,
		_w1250_,
		_w1289_
	);
	LUT3 #(
		.INIT('h0d)
	) name1224 (
		_w1252_,
		_w1253_,
		_w1254_,
		_w1290_
	);
	LUT4 #(
		.INIT('h153f)
	) name1225 (
		\a[11] ,
		\a[12] ,
		\a[22] ,
		\a[23] ,
		_w1291_
	);
	LUT4 #(
		.INIT('h8000)
	) name1226 (
		\a[11] ,
		\a[12] ,
		\a[22] ,
		\a[23] ,
		_w1292_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1227 (
		\a[11] ,
		\a[12] ,
		\a[22] ,
		\a[23] ,
		_w1293_
	);
	LUT2 #(
		.INIT('h6)
	) name1228 (
		_w1160_,
		_w1293_,
		_w1294_
	);
	LUT3 #(
		.INIT('h69)
	) name1229 (
		_w1289_,
		_w1290_,
		_w1294_,
		_w1295_
	);
	LUT4 #(
		.INIT('h0017)
	) name1230 (
		_w1247_,
		_w1251_,
		_w1256_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('he800)
	) name1231 (
		_w1247_,
		_w1251_,
		_w1256_,
		_w1295_,
		_w1297_
	);
	LUT4 #(
		.INIT('hf10e)
	) name1232 (
		_w1247_,
		_w1257_,
		_w1258_,
		_w1295_,
		_w1298_
	);
	LUT2 #(
		.INIT('h8)
	) name1233 (
		\a[13] ,
		\a[21] ,
		_w1299_
	);
	LUT4 #(
		.INIT('h153f)
	) name1234 (
		\a[14] ,
		\a[15] ,
		\a[19] ,
		\a[20] ,
		_w1300_
	);
	LUT4 #(
		.INIT('h8000)
	) name1235 (
		\a[14] ,
		\a[15] ,
		\a[19] ,
		\a[20] ,
		_w1301_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1236 (
		\a[14] ,
		\a[15] ,
		\a[19] ,
		\a[20] ,
		_w1302_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		\a[10] ,
		\a[24] ,
		_w1303_
	);
	LUT4 #(
		.INIT('h153f)
	) name1238 (
		\a[5] ,
		\a[9] ,
		\a[25] ,
		\a[29] ,
		_w1304_
	);
	LUT4 #(
		.INIT('h8000)
	) name1239 (
		\a[5] ,
		\a[9] ,
		\a[25] ,
		\a[29] ,
		_w1305_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1240 (
		\a[5] ,
		\a[9] ,
		\a[25] ,
		\a[29] ,
		_w1306_
	);
	LUT4 #(
		.INIT('h0660)
	) name1241 (
		_w1299_,
		_w1302_,
		_w1303_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('h9009)
	) name1242 (
		_w1299_,
		_w1302_,
		_w1303_,
		_w1306_,
		_w1308_
	);
	LUT4 #(
		.INIT('h6996)
	) name1243 (
		_w1299_,
		_w1302_,
		_w1303_,
		_w1306_,
		_w1309_
	);
	LUT4 #(
		.INIT('h153f)
	) name1244 (
		\a[7] ,
		\a[8] ,
		\a[26] ,
		\a[27] ,
		_w1310_
	);
	LUT4 #(
		.INIT('h8000)
	) name1245 (
		\a[7] ,
		\a[8] ,
		\a[26] ,
		\a[27] ,
		_w1311_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1246 (
		\a[7] ,
		\a[8] ,
		\a[26] ,
		\a[27] ,
		_w1312_
	);
	LUT2 #(
		.INIT('h6)
	) name1247 (
		_w1228_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h6)
	) name1248 (
		_w1309_,
		_w1313_,
		_w1314_
	);
	LUT3 #(
		.INIT('h28)
	) name1249 (
		_w1288_,
		_w1298_,
		_w1314_,
		_w1315_
	);
	LUT3 #(
		.INIT('h41)
	) name1250 (
		_w1288_,
		_w1298_,
		_w1314_,
		_w1316_
	);
	LUT3 #(
		.INIT('h96)
	) name1251 (
		_w1288_,
		_w1298_,
		_w1314_,
		_w1317_
	);
	LUT4 #(
		.INIT('hba45)
	) name1252 (
		_w1262_,
		_w1263_,
		_w1265_,
		_w1317_,
		_w1318_
	);
	LUT3 #(
		.INIT('hb2)
	) name1253 (
		_w1219_,
		_w1227_,
		_w1244_,
		_w1319_
	);
	LUT4 #(
		.INIT('hc0d4)
	) name1254 (
		_w1155_,
		_w1212_,
		_w1213_,
		_w1214_,
		_w1320_
	);
	LUT4 #(
		.INIT('h153f)
	) name1255 (
		\a[3] ,
		\a[4] ,
		\a[30] ,
		\a[31] ,
		_w1321_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		\a[4] ,
		\a[31] ,
		_w1322_
	);
	LUT4 #(
		.INIT('h8000)
	) name1257 (
		\a[3] ,
		\a[4] ,
		\a[30] ,
		\a[31] ,
		_w1323_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1258 (
		\a[3] ,
		\a[4] ,
		\a[30] ,
		\a[31] ,
		_w1324_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		\a[0] ,
		\a[34] ,
		_w1325_
	);
	LUT2 #(
		.INIT('h6)
	) name1260 (
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT4 #(
		.INIT('h008e)
	) name1261 (
		_w1216_,
		_w1217_,
		_w1218_,
		_w1326_,
		_w1327_
	);
	LUT4 #(
		.INIT('h7100)
	) name1262 (
		_w1216_,
		_w1217_,
		_w1218_,
		_w1326_,
		_w1328_
	);
	LUT3 #(
		.INIT('h8e)
	) name1263 (
		_w1220_,
		_w1221_,
		_w1226_,
		_w1329_
	);
	LUT3 #(
		.INIT('he1)
	) name1264 (
		_w1327_,
		_w1328_,
		_w1329_,
		_w1330_
	);
	LUT3 #(
		.INIT('h69)
	) name1265 (
		_w1319_,
		_w1320_,
		_w1330_,
		_w1331_
	);
	LUT4 #(
		.INIT('h0017)
	) name1266 (
		_w1211_,
		_w1215_,
		_w1245_,
		_w1331_,
		_w1332_
	);
	LUT4 #(
		.INIT('he800)
	) name1267 (
		_w1211_,
		_w1215_,
		_w1245_,
		_w1331_,
		_w1333_
	);
	LUT4 #(
		.INIT('h17e8)
	) name1268 (
		_w1211_,
		_w1215_,
		_w1245_,
		_w1331_,
		_w1334_
	);
	LUT2 #(
		.INIT('h6)
	) name1269 (
		_w1318_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		_w1275_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w1275_,
		_w1335_,
		_w1337_
	);
	LUT2 #(
		.INIT('h6)
	) name1272 (
		_w1275_,
		_w1335_,
		_w1338_
	);
	LUT2 #(
		.INIT('h9)
	) name1273 (
		_w1269_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1274 (
		_w1134_,
		_w1272_,
		_w1274_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('hc)
	) name1275 (
		_w1269_,
		_w1338_,
		_w1341_
	);
	LUT4 #(
		.INIT('hb000)
	) name1276 (
		_w1134_,
		_w1272_,
		_w1274_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('he)
	) name1277 (
		_w1340_,
		_w1342_,
		_w1343_
	);
	LUT3 #(
		.INIT('h32)
	) name1278 (
		_w1318_,
		_w1332_,
		_w1333_,
		_w1344_
	);
	LUT4 #(
		.INIT('h0071)
	) name1279 (
		_w1260_,
		_w1261_,
		_w1265_,
		_w1315_,
		_w1345_
	);
	LUT3 #(
		.INIT('h2b)
	) name1280 (
		_w1276_,
		_w1277_,
		_w1278_,
		_w1346_
	);
	LUT3 #(
		.INIT('h23)
	) name1281 (
		_w1283_,
		_w1284_,
		_w1286_,
		_w1347_
	);
	LUT3 #(
		.INIT('hb2)
	) name1282 (
		_w1289_,
		_w1290_,
		_w1294_,
		_w1348_
	);
	LUT3 #(
		.INIT('h96)
	) name1283 (
		_w1346_,
		_w1347_,
		_w1348_,
		_w1349_
	);
	LUT3 #(
		.INIT('h4d)
	) name1284 (
		_w1279_,
		_w1280_,
		_w1287_,
		_w1350_
	);
	LUT2 #(
		.INIT('h1)
	) name1285 (
		_w1349_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		_w1349_,
		_w1350_,
		_w1352_
	);
	LUT2 #(
		.INIT('h6)
	) name1287 (
		_w1349_,
		_w1350_,
		_w1353_
	);
	LUT3 #(
		.INIT('h54)
	) name1288 (
		_w1296_,
		_w1297_,
		_w1314_,
		_w1354_
	);
	LUT2 #(
		.INIT('h6)
	) name1289 (
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT3 #(
		.INIT('h8e)
	) name1290 (
		_w1319_,
		_w1320_,
		_w1330_,
		_w1356_
	);
	LUT3 #(
		.INIT('h0d)
	) name1291 (
		_w1160_,
		_w1291_,
		_w1292_,
		_w1357_
	);
	LUT3 #(
		.INIT('h0d)
	) name1292 (
		_w1299_,
		_w1300_,
		_w1301_,
		_w1358_
	);
	LUT3 #(
		.INIT('h23)
	) name1293 (
		_w1321_,
		_w1323_,
		_w1325_,
		_w1359_
	);
	LUT3 #(
		.INIT('h96)
	) name1294 (
		_w1357_,
		_w1358_,
		_w1359_,
		_w1360_
	);
	LUT3 #(
		.INIT('h80)
	) name1295 (
		\a[1] ,
		\a[18] ,
		\a[34] ,
		_w1361_
	);
	LUT3 #(
		.INIT('h6c)
	) name1296 (
		\a[1] ,
		\a[18] ,
		\a[34] ,
		_w1362_
	);
	LUT4 #(
		.INIT('h000d)
	) name1297 (
		_w1228_,
		_w1310_,
		_w1311_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('hf200)
	) name1298 (
		_w1228_,
		_w1310_,
		_w1311_,
		_w1362_,
		_w1364_
	);
	LUT4 #(
		.INIT('h0df2)
	) name1299 (
		_w1228_,
		_w1310_,
		_w1311_,
		_w1362_,
		_w1365_
	);
	LUT3 #(
		.INIT('h32)
	) name1300 (
		_w1303_,
		_w1304_,
		_w1305_,
		_w1366_
	);
	LUT2 #(
		.INIT('h6)
	) name1301 (
		_w1365_,
		_w1366_,
		_w1367_
	);
	LUT3 #(
		.INIT('h32)
	) name1302 (
		_w1307_,
		_w1308_,
		_w1313_,
		_w1368_
	);
	LUT3 #(
		.INIT('h69)
	) name1303 (
		_w1360_,
		_w1367_,
		_w1368_,
		_w1369_
	);
	LUT3 #(
		.INIT('h45)
	) name1304 (
		_w1327_,
		_w1328_,
		_w1329_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		\a[5] ,
		\a[30] ,
		_w1371_
	);
	LUT4 #(
		.INIT('h153f)
	) name1306 (
		\a[6] ,
		\a[8] ,
		\a[27] ,
		\a[29] ,
		_w1372_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		\a[8] ,
		\a[29] ,
		_w1373_
	);
	LUT4 #(
		.INIT('h8000)
	) name1308 (
		\a[6] ,
		\a[8] ,
		\a[27] ,
		\a[29] ,
		_w1374_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1309 (
		\a[6] ,
		\a[8] ,
		\a[27] ,
		\a[29] ,
		_w1375_
	);
	LUT2 #(
		.INIT('h8)
	) name1310 (
		\a[7] ,
		\a[28] ,
		_w1376_
	);
	LUT4 #(
		.INIT('h153f)
	) name1311 (
		\a[16] ,
		\a[17] ,
		\a[18] ,
		\a[19] ,
		_w1377_
	);
	LUT4 #(
		.INIT('h8000)
	) name1312 (
		\a[16] ,
		\a[17] ,
		\a[18] ,
		\a[19] ,
		_w1378_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1313 (
		\a[16] ,
		\a[17] ,
		\a[18] ,
		\a[19] ,
		_w1379_
	);
	LUT4 #(
		.INIT('h0660)
	) name1314 (
		_w1371_,
		_w1375_,
		_w1376_,
		_w1379_,
		_w1380_
	);
	LUT4 #(
		.INIT('h9009)
	) name1315 (
		_w1371_,
		_w1375_,
		_w1376_,
		_w1379_,
		_w1381_
	);
	LUT4 #(
		.INIT('h6996)
	) name1316 (
		_w1371_,
		_w1375_,
		_w1376_,
		_w1379_,
		_w1382_
	);
	LUT4 #(
		.INIT('h153f)
	) name1317 (
		\a[9] ,
		\a[10] ,
		\a[25] ,
		\a[26] ,
		_w1383_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		\a[10] ,
		\a[26] ,
		_w1384_
	);
	LUT4 #(
		.INIT('h8000)
	) name1319 (
		\a[9] ,
		\a[10] ,
		\a[25] ,
		\a[26] ,
		_w1385_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1320 (
		\a[9] ,
		\a[10] ,
		\a[25] ,
		\a[26] ,
		_w1386_
	);
	LUT2 #(
		.INIT('h6)
	) name1321 (
		_w1322_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h6)
	) name1322 (
		_w1382_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h153f)
	) name1323 (
		\a[0] ,
		\a[2] ,
		\a[33] ,
		\a[35] ,
		_w1389_
	);
	LUT4 #(
		.INIT('h8000)
	) name1324 (
		\a[0] ,
		\a[2] ,
		\a[33] ,
		\a[35] ,
		_w1390_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1325 (
		\a[0] ,
		\a[2] ,
		\a[33] ,
		\a[35] ,
		_w1391_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		\a[3] ,
		\a[32] ,
		_w1392_
	);
	LUT4 #(
		.INIT('h153f)
	) name1327 (
		\a[11] ,
		\a[12] ,
		\a[23] ,
		\a[24] ,
		_w1393_
	);
	LUT4 #(
		.INIT('h8000)
	) name1328 (
		\a[11] ,
		\a[12] ,
		\a[23] ,
		\a[24] ,
		_w1394_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1329 (
		\a[11] ,
		\a[12] ,
		\a[23] ,
		\a[24] ,
		_w1395_
	);
	LUT4 #(
		.INIT('h0660)
	) name1330 (
		_w1281_,
		_w1391_,
		_w1392_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('h9009)
	) name1331 (
		_w1281_,
		_w1391_,
		_w1392_,
		_w1395_,
		_w1397_
	);
	LUT4 #(
		.INIT('h6996)
	) name1332 (
		_w1281_,
		_w1391_,
		_w1392_,
		_w1395_,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name1333 (
		\a[13] ,
		\a[22] ,
		_w1399_
	);
	LUT4 #(
		.INIT('h153f)
	) name1334 (
		\a[14] ,
		\a[15] ,
		\a[20] ,
		\a[21] ,
		_w1400_
	);
	LUT4 #(
		.INIT('h8000)
	) name1335 (
		\a[14] ,
		\a[15] ,
		\a[20] ,
		\a[21] ,
		_w1401_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1336 (
		\a[14] ,
		\a[15] ,
		\a[20] ,
		\a[21] ,
		_w1402_
	);
	LUT2 #(
		.INIT('h6)
	) name1337 (
		_w1399_,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h6)
	) name1338 (
		_w1398_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1339 (
		_w1327_,
		_w1328_,
		_w1329_,
		_w1388_,
		_w1405_
	);
	LUT3 #(
		.INIT('h96)
	) name1340 (
		_w1370_,
		_w1388_,
		_w1404_,
		_w1406_
	);
	LUT4 #(
		.INIT('h4114)
	) name1341 (
		_w1369_,
		_w1370_,
		_w1388_,
		_w1404_,
		_w1407_
	);
	LUT4 #(
		.INIT('h8228)
	) name1342 (
		_w1369_,
		_w1370_,
		_w1388_,
		_w1404_,
		_w1408_
	);
	LUT3 #(
		.INIT('h9f)
	) name1343 (
		_w1356_,
		_w1369_,
		_w1406_,
		_w1409_
	);
	LUT3 #(
		.INIT('h96)
	) name1344 (
		_w1356_,
		_w1369_,
		_w1406_,
		_w1410_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name1345 (
		_w1316_,
		_w1345_,
		_w1355_,
		_w1410_,
		_w1411_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		_w1344_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h6)
	) name1347 (
		_w1344_,
		_w1411_,
		_w1413_
	);
	LUT3 #(
		.INIT('h01)
	) name1348 (
		_w1205_,
		_w1270_,
		_w1336_,
		_w1414_
	);
	LUT3 #(
		.INIT('hb0)
	) name1349 (
		_w1134_,
		_w1272_,
		_w1414_,
		_w1415_
	);
	LUT3 #(
		.INIT('h0d)
	) name1350 (
		_w1269_,
		_w1336_,
		_w1337_,
		_w1416_
	);
	LUT3 #(
		.INIT('h9a)
	) name1351 (
		_w1413_,
		_w1415_,
		_w1416_,
		_w1417_
	);
	LUT4 #(
		.INIT('heee0)
	) name1352 (
		_w1275_,
		_w1335_,
		_w1344_,
		_w1411_,
		_w1418_
	);
	LUT3 #(
		.INIT('hd0)
	) name1353 (
		_w1269_,
		_w1336_,
		_w1418_,
		_w1419_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1354 (
		_w1134_,
		_w1272_,
		_w1414_,
		_w1419_,
		_w1420_
	);
	LUT4 #(
		.INIT('hf110)
	) name1355 (
		_w1316_,
		_w1345_,
		_w1355_,
		_w1410_,
		_w1421_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1356 (
		_w1319_,
		_w1320_,
		_w1330_,
		_w1369_,
		_w1422_
	);
	LUT4 #(
		.INIT('h0027)
	) name1357 (
		_w1356_,
		_w1407_,
		_w1408_,
		_w1422_,
		_w1423_
	);
	LUT3 #(
		.INIT('h17)
	) name1358 (
		_w1357_,
		_w1358_,
		_w1359_,
		_w1424_
	);
	LUT3 #(
		.INIT('h54)
	) name1359 (
		_w1363_,
		_w1364_,
		_w1366_,
		_w1425_
	);
	LUT3 #(
		.INIT('h32)
	) name1360 (
		_w1396_,
		_w1397_,
		_w1403_,
		_w1426_
	);
	LUT3 #(
		.INIT('h96)
	) name1361 (
		_w1424_,
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT3 #(
		.INIT('hd4)
	) name1362 (
		_w1360_,
		_w1367_,
		_w1368_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		_w1427_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		_w1427_,
		_w1428_,
		_w1430_
	);
	LUT2 #(
		.INIT('h6)
	) name1365 (
		_w1427_,
		_w1428_,
		_w1431_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1366 (
		_w1327_,
		_w1328_,
		_w1329_,
		_w1404_,
		_w1432_
	);
	LUT4 #(
		.INIT('h9009)
	) name1367 (
		_w1382_,
		_w1387_,
		_w1398_,
		_w1403_,
		_w1433_
	);
	LUT3 #(
		.INIT('h01)
	) name1368 (
		_w1405_,
		_w1432_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h6)
	) name1369 (
		_w1431_,
		_w1434_,
		_w1435_
	);
	LUT2 #(
		.INIT('h4)
	) name1370 (
		_w1423_,
		_w1435_,
		_w1436_
	);
	LUT3 #(
		.INIT('h41)
	) name1371 (
		_w1422_,
		_w1431_,
		_w1434_,
		_w1437_
	);
	LUT2 #(
		.INIT('h8)
	) name1372 (
		_w1409_,
		_w1437_,
		_w1438_
	);
	LUT3 #(
		.INIT('h54)
	) name1373 (
		_w1351_,
		_w1352_,
		_w1354_,
		_w1439_
	);
	LUT3 #(
		.INIT('h0d)
	) name1374 (
		_w1322_,
		_w1383_,
		_w1385_,
		_w1440_
	);
	LUT3 #(
		.INIT('h0d)
	) name1375 (
		_w1371_,
		_w1372_,
		_w1374_,
		_w1441_
	);
	LUT3 #(
		.INIT('h32)
	) name1376 (
		_w1376_,
		_w1377_,
		_w1378_,
		_w1442_
	);
	LUT3 #(
		.INIT('h96)
	) name1377 (
		_w1440_,
		_w1441_,
		_w1442_,
		_w1443_
	);
	LUT3 #(
		.INIT('h0d)
	) name1378 (
		_w1392_,
		_w1393_,
		_w1394_,
		_w1444_
	);
	LUT3 #(
		.INIT('h0d)
	) name1379 (
		_w1399_,
		_w1400_,
		_w1401_,
		_w1445_
	);
	LUT3 #(
		.INIT('h0d)
	) name1380 (
		_w1281_,
		_w1389_,
		_w1390_,
		_w1446_
	);
	LUT3 #(
		.INIT('h96)
	) name1381 (
		_w1444_,
		_w1445_,
		_w1446_,
		_w1447_
	);
	LUT3 #(
		.INIT('h32)
	) name1382 (
		_w1380_,
		_w1381_,
		_w1387_,
		_w1448_
	);
	LUT3 #(
		.INIT('h69)
	) name1383 (
		_w1443_,
		_w1447_,
		_w1448_,
		_w1449_
	);
	LUT3 #(
		.INIT('he8)
	) name1384 (
		_w1346_,
		_w1347_,
		_w1348_,
		_w1450_
	);
	LUT4 #(
		.INIT('h8000)
	) name1385 (
		\a[1] ,
		\a[17] ,
		\a[19] ,
		\a[35] ,
		_w1451_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1386 (
		\a[1] ,
		\a[17] ,
		\a[19] ,
		\a[35] ,
		_w1452_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		\a[0] ,
		\a[36] ,
		_w1453_
	);
	LUT3 #(
		.INIT('h96)
	) name1388 (
		_w1361_,
		_w1452_,
		_w1453_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		\a[14] ,
		\a[22] ,
		_w1455_
	);
	LUT4 #(
		.INIT('h153f)
	) name1390 (
		\a[15] ,
		\a[16] ,
		\a[20] ,
		\a[21] ,
		_w1456_
	);
	LUT2 #(
		.INIT('h8)
	) name1391 (
		\a[16] ,
		\a[21] ,
		_w1457_
	);
	LUT4 #(
		.INIT('h8000)
	) name1392 (
		\a[15] ,
		\a[16] ,
		\a[20] ,
		\a[21] ,
		_w1458_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1393 (
		\a[15] ,
		\a[16] ,
		\a[20] ,
		\a[21] ,
		_w1459_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		\a[3] ,
		\a[33] ,
		_w1460_
	);
	LUT4 #(
		.INIT('h153f)
	) name1395 (
		\a[4] ,
		\a[11] ,
		\a[25] ,
		\a[32] ,
		_w1461_
	);
	LUT4 #(
		.INIT('h8000)
	) name1396 (
		\a[4] ,
		\a[11] ,
		\a[25] ,
		\a[32] ,
		_w1462_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1397 (
		\a[4] ,
		\a[11] ,
		\a[25] ,
		\a[32] ,
		_w1463_
	);
	LUT4 #(
		.INIT('h0660)
	) name1398 (
		_w1455_,
		_w1459_,
		_w1460_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('h9009)
	) name1399 (
		_w1455_,
		_w1459_,
		_w1460_,
		_w1463_,
		_w1465_
	);
	LUT4 #(
		.INIT('h6996)
	) name1400 (
		_w1455_,
		_w1459_,
		_w1460_,
		_w1463_,
		_w1466_
	);
	LUT2 #(
		.INIT('h6)
	) name1401 (
		_w1454_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h8)
	) name1402 (
		\a[2] ,
		\a[34] ,
		_w1468_
	);
	LUT4 #(
		.INIT('h153f)
	) name1403 (
		\a[12] ,
		\a[13] ,
		\a[23] ,
		\a[24] ,
		_w1469_
	);
	LUT2 #(
		.INIT('h8)
	) name1404 (
		\a[13] ,
		\a[24] ,
		_w1470_
	);
	LUT4 #(
		.INIT('h8000)
	) name1405 (
		\a[12] ,
		\a[13] ,
		\a[23] ,
		\a[24] ,
		_w1471_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1406 (
		\a[12] ,
		\a[13] ,
		\a[23] ,
		\a[24] ,
		_w1472_
	);
	LUT4 #(
		.INIT('h153f)
	) name1407 (
		\a[5] ,
		\a[9] ,
		\a[27] ,
		\a[31] ,
		_w1473_
	);
	LUT4 #(
		.INIT('h8000)
	) name1408 (
		\a[5] ,
		\a[9] ,
		\a[27] ,
		\a[31] ,
		_w1474_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1409 (
		\a[5] ,
		\a[9] ,
		\a[27] ,
		\a[31] ,
		_w1475_
	);
	LUT4 #(
		.INIT('h1428)
	) name1410 (
		_w1384_,
		_w1468_,
		_w1472_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h8241)
	) name1411 (
		_w1384_,
		_w1468_,
		_w1472_,
		_w1475_,
		_w1477_
	);
	LUT4 #(
		.INIT('h6996)
	) name1412 (
		_w1384_,
		_w1468_,
		_w1472_,
		_w1475_,
		_w1478_
	);
	LUT2 #(
		.INIT('h8)
	) name1413 (
		\a[6] ,
		\a[30] ,
		_w1479_
	);
	LUT4 #(
		.INIT('h153f)
	) name1414 (
		\a[7] ,
		\a[8] ,
		\a[28] ,
		\a[29] ,
		_w1480_
	);
	LUT4 #(
		.INIT('h8000)
	) name1415 (
		\a[7] ,
		\a[8] ,
		\a[28] ,
		\a[29] ,
		_w1481_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1416 (
		\a[7] ,
		\a[8] ,
		\a[28] ,
		\a[29] ,
		_w1482_
	);
	LUT2 #(
		.INIT('h6)
	) name1417 (
		_w1479_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('h6)
	) name1418 (
		_w1478_,
		_w1483_,
		_w1484_
	);
	LUT3 #(
		.INIT('h96)
	) name1419 (
		_w1450_,
		_w1467_,
		_w1484_,
		_w1485_
	);
	LUT4 #(
		.INIT('h4114)
	) name1420 (
		_w1449_,
		_w1450_,
		_w1467_,
		_w1484_,
		_w1486_
	);
	LUT4 #(
		.INIT('he800)
	) name1421 (
		_w1349_,
		_w1350_,
		_w1354_,
		_w1486_,
		_w1487_
	);
	LUT4 #(
		.INIT('h8228)
	) name1422 (
		_w1449_,
		_w1450_,
		_w1467_,
		_w1484_,
		_w1488_
	);
	LUT4 #(
		.INIT('h1700)
	) name1423 (
		_w1349_,
		_w1350_,
		_w1354_,
		_w1488_,
		_w1489_
	);
	LUT3 #(
		.INIT('h96)
	) name1424 (
		_w1439_,
		_w1449_,
		_w1485_,
		_w1490_
	);
	LUT4 #(
		.INIT('h0154)
	) name1425 (
		_w1421_,
		_w1436_,
		_w1438_,
		_w1490_,
		_w1491_
	);
	LUT4 #(
		.INIT('ha802)
	) name1426 (
		_w1421_,
		_w1436_,
		_w1438_,
		_w1490_,
		_w1492_
	);
	LUT4 #(
		.INIT('h56a9)
	) name1427 (
		_w1421_,
		_w1436_,
		_w1438_,
		_w1490_,
		_w1493_
	);
	LUT3 #(
		.INIT('h1e)
	) name1428 (
		_w1412_,
		_w1420_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h1)
	) name1429 (
		_w1412_,
		_w1492_,
		_w1495_
	);
	LUT3 #(
		.INIT('he8)
	) name1430 (
		_w1427_,
		_w1428_,
		_w1434_,
		_w1496_
	);
	LUT3 #(
		.INIT('h32)
	) name1431 (
		_w1460_,
		_w1461_,
		_w1462_,
		_w1497_
	);
	LUT3 #(
		.INIT('h0d)
	) name1432 (
		_w1455_,
		_w1456_,
		_w1458_,
		_w1498_
	);
	LUT3 #(
		.INIT('h0d)
	) name1433 (
		_w1468_,
		_w1469_,
		_w1471_,
		_w1499_
	);
	LUT3 #(
		.INIT('h69)
	) name1434 (
		_w1497_,
		_w1498_,
		_w1499_,
		_w1500_
	);
	LUT3 #(
		.INIT('h0e)
	) name1435 (
		_w1454_,
		_w1464_,
		_w1465_,
		_w1501_
	);
	LUT3 #(
		.INIT('he8)
	) name1436 (
		_w1361_,
		_w1452_,
		_w1453_,
		_w1502_
	);
	LUT3 #(
		.INIT('h0d)
	) name1437 (
		_w1384_,
		_w1473_,
		_w1474_,
		_w1503_
	);
	LUT4 #(
		.INIT('h153f)
	) name1438 (
		\a[14] ,
		\a[15] ,
		\a[22] ,
		\a[23] ,
		_w1504_
	);
	LUT2 #(
		.INIT('h8)
	) name1439 (
		\a[15] ,
		\a[23] ,
		_w1505_
	);
	LUT4 #(
		.INIT('h8000)
	) name1440 (
		\a[14] ,
		\a[15] ,
		\a[22] ,
		\a[23] ,
		_w1506_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1441 (
		\a[14] ,
		\a[15] ,
		\a[22] ,
		\a[23] ,
		_w1507_
	);
	LUT2 #(
		.INIT('h6)
	) name1442 (
		_w1470_,
		_w1507_,
		_w1508_
	);
	LUT3 #(
		.INIT('h69)
	) name1443 (
		_w1502_,
		_w1503_,
		_w1508_,
		_w1509_
	);
	LUT3 #(
		.INIT('h69)
	) name1444 (
		_w1500_,
		_w1501_,
		_w1509_,
		_w1510_
	);
	LUT3 #(
		.INIT('he8)
	) name1445 (
		_w1424_,
		_w1425_,
		_w1426_,
		_w1511_
	);
	LUT2 #(
		.INIT('h8)
	) name1446 (
		\a[11] ,
		\a[26] ,
		_w1512_
	);
	LUT4 #(
		.INIT('h153f)
	) name1447 (
		\a[5] ,
		\a[10] ,
		\a[27] ,
		\a[32] ,
		_w1513_
	);
	LUT2 #(
		.INIT('h8)
	) name1448 (
		\a[10] ,
		\a[32] ,
		_w1514_
	);
	LUT4 #(
		.INIT('h8000)
	) name1449 (
		\a[5] ,
		\a[10] ,
		\a[27] ,
		\a[32] ,
		_w1515_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1450 (
		\a[5] ,
		\a[10] ,
		\a[27] ,
		\a[32] ,
		_w1516_
	);
	LUT4 #(
		.INIT('h153f)
	) name1451 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w1517_
	);
	LUT4 #(
		.INIT('h8000)
	) name1452 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w1518_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1453 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w1519_
	);
	LUT4 #(
		.INIT('h1428)
	) name1454 (
		_w1373_,
		_w1512_,
		_w1516_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h6996)
	) name1455 (
		_w1373_,
		_w1512_,
		_w1516_,
		_w1519_,
		_w1521_
	);
	LUT4 #(
		.INIT('h1700)
	) name1456 (
		_w1444_,
		_w1445_,
		_w1446_,
		_w1521_,
		_w1522_
	);
	LUT4 #(
		.INIT('he817)
	) name1457 (
		_w1444_,
		_w1445_,
		_w1446_,
		_w1521_,
		_w1523_
	);
	LUT4 #(
		.INIT('h153f)
	) name1458 (
		\a[2] ,
		\a[3] ,
		\a[34] ,
		\a[35] ,
		_w1524_
	);
	LUT2 #(
		.INIT('h8)
	) name1459 (
		\a[3] ,
		\a[35] ,
		_w1525_
	);
	LUT4 #(
		.INIT('h8000)
	) name1460 (
		\a[2] ,
		\a[3] ,
		\a[34] ,
		\a[35] ,
		_w1526_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1461 (
		\a[2] ,
		\a[3] ,
		\a[34] ,
		\a[35] ,
		_w1527_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		\a[0] ,
		\a[37] ,
		_w1528_
	);
	LUT4 #(
		.INIT('h153f)
	) name1463 (
		\a[4] ,
		\a[12] ,
		\a[25] ,
		\a[33] ,
		_w1529_
	);
	LUT2 #(
		.INIT('h8)
	) name1464 (
		\a[12] ,
		\a[33] ,
		_w1530_
	);
	LUT4 #(
		.INIT('h8000)
	) name1465 (
		\a[4] ,
		\a[12] ,
		\a[25] ,
		\a[33] ,
		_w1531_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1466 (
		\a[4] ,
		\a[12] ,
		\a[25] ,
		\a[33] ,
		_w1532_
	);
	LUT4 #(
		.INIT('h0660)
	) name1467 (
		_w1457_,
		_w1527_,
		_w1528_,
		_w1532_,
		_w1533_
	);
	LUT4 #(
		.INIT('h9009)
	) name1468 (
		_w1457_,
		_w1527_,
		_w1528_,
		_w1532_,
		_w1534_
	);
	LUT4 #(
		.INIT('h6996)
	) name1469 (
		_w1457_,
		_w1527_,
		_w1528_,
		_w1532_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name1470 (
		\a[9] ,
		\a[28] ,
		_w1536_
	);
	LUT4 #(
		.INIT('h153f)
	) name1471 (
		\a[6] ,
		\a[7] ,
		\a[30] ,
		\a[31] ,
		_w1537_
	);
	LUT4 #(
		.INIT('h8000)
	) name1472 (
		\a[6] ,
		\a[7] ,
		\a[30] ,
		\a[31] ,
		_w1538_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1473 (
		\a[6] ,
		\a[7] ,
		\a[30] ,
		\a[31] ,
		_w1539_
	);
	LUT2 #(
		.INIT('h6)
	) name1474 (
		_w1536_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h6)
	) name1475 (
		_w1535_,
		_w1540_,
		_w1541_
	);
	LUT3 #(
		.INIT('h96)
	) name1476 (
		_w1511_,
		_w1523_,
		_w1541_,
		_w1542_
	);
	LUT4 #(
		.INIT('h4114)
	) name1477 (
		_w1510_,
		_w1511_,
		_w1523_,
		_w1541_,
		_w1543_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1478 (
		_w1429_,
		_w1430_,
		_w1434_,
		_w1543_,
		_w1544_
	);
	LUT4 #(
		.INIT('h8228)
	) name1479 (
		_w1510_,
		_w1511_,
		_w1523_,
		_w1541_,
		_w1545_
	);
	LUT4 #(
		.INIT('h2300)
	) name1480 (
		_w1429_,
		_w1430_,
		_w1434_,
		_w1545_,
		_w1546_
	);
	LUT3 #(
		.INIT('h96)
	) name1481 (
		_w1496_,
		_w1510_,
		_w1542_,
		_w1547_
	);
	LUT3 #(
		.INIT('he0)
	) name1482 (
		_w1349_,
		_w1350_,
		_w1449_,
		_w1548_
	);
	LUT3 #(
		.INIT('he0)
	) name1483 (
		_w1352_,
		_w1354_,
		_w1548_,
		_w1549_
	);
	LUT3 #(
		.INIT('hb2)
	) name1484 (
		_w1443_,
		_w1447_,
		_w1448_,
		_w1550_
	);
	LUT3 #(
		.INIT('h71)
	) name1485 (
		_w1440_,
		_w1441_,
		_w1442_,
		_w1551_
	);
	LUT2 #(
		.INIT('h4)
	) name1486 (
		\a[36] ,
		_w1451_,
		_w1552_
	);
	LUT3 #(
		.INIT('h80)
	) name1487 (
		\a[1] ,
		\a[19] ,
		\a[36] ,
		_w1553_
	);
	LUT3 #(
		.INIT('h6c)
	) name1488 (
		\a[1] ,
		\a[19] ,
		\a[36] ,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w1451_,
		_w1554_,
		_w1555_
	);
	LUT3 #(
		.INIT('hb8)
	) name1490 (
		\a[36] ,
		_w1451_,
		_w1554_,
		_w1556_
	);
	LUT3 #(
		.INIT('h0d)
	) name1491 (
		_w1479_,
		_w1480_,
		_w1481_,
		_w1557_
	);
	LUT2 #(
		.INIT('h6)
	) name1492 (
		_w1556_,
		_w1557_,
		_w1558_
	);
	LUT3 #(
		.INIT('h32)
	) name1493 (
		_w1476_,
		_w1477_,
		_w1483_,
		_w1559_
	);
	LUT3 #(
		.INIT('h69)
	) name1494 (
		_w1551_,
		_w1558_,
		_w1559_,
		_w1560_
	);
	LUT2 #(
		.INIT('h6)
	) name1495 (
		_w1550_,
		_w1560_,
		_w1561_
	);
	LUT4 #(
		.INIT('h0017)
	) name1496 (
		_w1346_,
		_w1347_,
		_w1348_,
		_w1467_,
		_w1562_
	);
	LUT4 #(
		.INIT('he800)
	) name1497 (
		_w1346_,
		_w1347_,
		_w1348_,
		_w1467_,
		_w1563_
	);
	LUT3 #(
		.INIT('h32)
	) name1498 (
		_w1484_,
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h6)
	) name1499 (
		_w1561_,
		_w1564_,
		_w1565_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1500 (
		_w1487_,
		_w1489_,
		_w1549_,
		_w1565_,
		_w1566_
	);
	LUT4 #(
		.INIT('h0001)
	) name1501 (
		_w1487_,
		_w1489_,
		_w1549_,
		_w1565_,
		_w1567_
	);
	LUT4 #(
		.INIT('h01fe)
	) name1502 (
		_w1487_,
		_w1489_,
		_w1549_,
		_w1565_,
		_w1568_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w1547_,
		_w1568_,
		_w1569_
	);
	LUT3 #(
		.INIT('h45)
	) name1504 (
		_w1436_,
		_w1438_,
		_w1490_,
		_w1570_
	);
	LUT3 #(
		.INIT('h02)
	) name1505 (
		_w1547_,
		_w1566_,
		_w1567_,
		_w1571_
	);
	LUT3 #(
		.INIT('h01)
	) name1506 (
		_w1569_,
		_w1570_,
		_w1571_,
		_w1572_
	);
	LUT3 #(
		.INIT('ha9)
	) name1507 (
		_w1547_,
		_w1566_,
		_w1567_,
		_w1573_
	);
	LUT2 #(
		.INIT('h2)
	) name1508 (
		_w1570_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h36)
	) name1509 (
		_w1569_,
		_w1570_,
		_w1571_,
		_w1575_
	);
	LUT4 #(
		.INIT('hdc23)
	) name1510 (
		_w1420_,
		_w1491_,
		_w1495_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1511 (
		_w1420_,
		_w1491_,
		_w1495_,
		_w1572_,
		_w1577_
	);
	LUT3 #(
		.INIT('h0e)
	) name1512 (
		_w1547_,
		_w1566_,
		_w1567_,
		_w1578_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1513 (
		_w1429_,
		_w1430_,
		_w1434_,
		_w1510_,
		_w1579_
	);
	LUT3 #(
		.INIT('hd4)
	) name1514 (
		_w1500_,
		_w1501_,
		_w1509_,
		_w1580_
	);
	LUT4 #(
		.INIT('he800)
	) name1515 (
		_w1511_,
		_w1523_,
		_w1541_,
		_w1580_,
		_w1581_
	);
	LUT3 #(
		.INIT('h0d)
	) name1516 (
		_w1528_,
		_w1529_,
		_w1531_,
		_w1582_
	);
	LUT3 #(
		.INIT('h0d)
	) name1517 (
		_w1457_,
		_w1524_,
		_w1526_,
		_w1583_
	);
	LUT3 #(
		.INIT('h0d)
	) name1518 (
		_w1470_,
		_w1504_,
		_w1506_,
		_w1584_
	);
	LUT3 #(
		.INIT('h96)
	) name1519 (
		_w1582_,
		_w1583_,
		_w1584_,
		_w1585_
	);
	LUT4 #(
		.INIT('h153f)
	) name1520 (
		\a[16] ,
		\a[17] ,
		\a[21] ,
		\a[22] ,
		_w1586_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		\a[17] ,
		\a[22] ,
		_w1587_
	);
	LUT4 #(
		.INIT('h8000)
	) name1522 (
		\a[16] ,
		\a[17] ,
		\a[21] ,
		\a[22] ,
		_w1588_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1523 (
		\a[16] ,
		\a[17] ,
		\a[21] ,
		\a[22] ,
		_w1589_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		\a[5] ,
		\a[33] ,
		_w1590_
	);
	LUT4 #(
		.INIT('h153f)
	) name1525 (
		\a[6] ,
		\a[10] ,
		\a[28] ,
		\a[32] ,
		_w1591_
	);
	LUT4 #(
		.INIT('h8000)
	) name1526 (
		\a[6] ,
		\a[10] ,
		\a[28] ,
		\a[32] ,
		_w1592_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1527 (
		\a[6] ,
		\a[10] ,
		\a[28] ,
		\a[32] ,
		_w1593_
	);
	LUT4 #(
		.INIT('h0660)
	) name1528 (
		_w1505_,
		_w1589_,
		_w1590_,
		_w1593_,
		_w1594_
	);
	LUT4 #(
		.INIT('h9009)
	) name1529 (
		_w1505_,
		_w1589_,
		_w1590_,
		_w1593_,
		_w1595_
	);
	LUT4 #(
		.INIT('h6996)
	) name1530 (
		_w1505_,
		_w1589_,
		_w1590_,
		_w1593_,
		_w1596_
	);
	LUT2 #(
		.INIT('h8)
	) name1531 (
		\a[9] ,
		\a[29] ,
		_w1597_
	);
	LUT4 #(
		.INIT('h153f)
	) name1532 (
		\a[7] ,
		\a[8] ,
		\a[30] ,
		\a[31] ,
		_w1598_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		\a[8] ,
		\a[31] ,
		_w1599_
	);
	LUT4 #(
		.INIT('h8000)
	) name1534 (
		\a[7] ,
		\a[8] ,
		\a[30] ,
		\a[31] ,
		_w1600_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1535 (
		\a[7] ,
		\a[8] ,
		\a[30] ,
		\a[31] ,
		_w1601_
	);
	LUT2 #(
		.INIT('h6)
	) name1536 (
		_w1597_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h6)
	) name1537 (
		_w1596_,
		_w1602_,
		_w1603_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name1538 (
		_w1520_,
		_w1522_,
		_w1585_,
		_w1603_,
		_w1604_
	);
	LUT4 #(
		.INIT('h0017)
	) name1539 (
		_w1511_,
		_w1523_,
		_w1541_,
		_w1580_,
		_w1605_
	);
	LUT3 #(
		.INIT('hc9)
	) name1540 (
		_w1581_,
		_w1604_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('h0001)
	) name1541 (
		_w1544_,
		_w1546_,
		_w1579_,
		_w1606_,
		_w1607_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1542 (
		_w1544_,
		_w1546_,
		_w1579_,
		_w1606_,
		_w1608_
	);
	LUT4 #(
		.INIT('h17e8)
	) name1543 (
		_w1496_,
		_w1510_,
		_w1542_,
		_w1606_,
		_w1609_
	);
	LUT3 #(
		.INIT('h32)
	) name1544 (
		_w1533_,
		_w1534_,
		_w1540_,
		_w1610_
	);
	LUT3 #(
		.INIT('hb2)
	) name1545 (
		_w1502_,
		_w1503_,
		_w1508_,
		_w1611_
	);
	LUT4 #(
		.INIT('h8000)
	) name1546 (
		\a[1] ,
		\a[18] ,
		\a[20] ,
		\a[37] ,
		_w1612_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1547 (
		\a[1] ,
		\a[18] ,
		\a[20] ,
		\a[37] ,
		_w1613_
	);
	LUT3 #(
		.INIT('h0d)
	) name1548 (
		_w1373_,
		_w1517_,
		_w1518_,
		_w1614_
	);
	LUT4 #(
		.INIT('h000d)
	) name1549 (
		_w1373_,
		_w1517_,
		_w1518_,
		_w1613_,
		_w1615_
	);
	LUT4 #(
		.INIT('hf200)
	) name1550 (
		_w1373_,
		_w1517_,
		_w1518_,
		_w1613_,
		_w1616_
	);
	LUT4 #(
		.INIT('h0df2)
	) name1551 (
		_w1373_,
		_w1517_,
		_w1518_,
		_w1613_,
		_w1617_
	);
	LUT3 #(
		.INIT('h0d)
	) name1552 (
		_w1536_,
		_w1537_,
		_w1538_,
		_w1618_
	);
	LUT2 #(
		.INIT('h6)
	) name1553 (
		_w1617_,
		_w1618_,
		_w1619_
	);
	LUT3 #(
		.INIT('h69)
	) name1554 (
		_w1610_,
		_w1611_,
		_w1619_,
		_w1620_
	);
	LUT4 #(
		.INIT('he800)
	) name1555 (
		_w1550_,
		_w1560_,
		_w1564_,
		_w1620_,
		_w1621_
	);
	LUT3 #(
		.INIT('h07)
	) name1556 (
		_w1550_,
		_w1560_,
		_w1620_,
		_w1622_
	);
	LUT3 #(
		.INIT('h70)
	) name1557 (
		_w1561_,
		_w1564_,
		_w1622_,
		_w1623_
	);
	LUT3 #(
		.INIT('h2b)
	) name1558 (
		_w1497_,
		_w1498_,
		_w1499_,
		_w1624_
	);
	LUT3 #(
		.INIT('h23)
	) name1559 (
		_w1552_,
		_w1555_,
		_w1557_,
		_w1625_
	);
	LUT2 #(
		.INIT('h8)
	) name1560 (
		\a[12] ,
		\a[26] ,
		_w1626_
	);
	LUT4 #(
		.INIT('h153f)
	) name1561 (
		\a[4] ,
		\a[11] ,
		\a[27] ,
		\a[34] ,
		_w1627_
	);
	LUT4 #(
		.INIT('h8000)
	) name1562 (
		\a[4] ,
		\a[11] ,
		\a[27] ,
		\a[34] ,
		_w1628_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1563 (
		\a[4] ,
		\a[11] ,
		\a[27] ,
		\a[34] ,
		_w1629_
	);
	LUT2 #(
		.INIT('h6)
	) name1564 (
		_w1626_,
		_w1629_,
		_w1630_
	);
	LUT4 #(
		.INIT('h2300)
	) name1565 (
		_w1552_,
		_w1555_,
		_w1557_,
		_w1630_,
		_w1631_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1566 (
		_w1552_,
		_w1555_,
		_w1557_,
		_w1630_,
		_w1632_
	);
	LUT4 #(
		.INIT('hdc23)
	) name1567 (
		_w1552_,
		_w1555_,
		_w1557_,
		_w1630_,
		_w1633_
	);
	LUT2 #(
		.INIT('h6)
	) name1568 (
		_w1624_,
		_w1633_,
		_w1634_
	);
	LUT3 #(
		.INIT('h0d)
	) name1569 (
		_w1512_,
		_w1513_,
		_w1515_,
		_w1635_
	);
	LUT4 #(
		.INIT('h153f)
	) name1570 (
		\a[0] ,
		\a[2] ,
		\a[36] ,
		\a[38] ,
		_w1636_
	);
	LUT4 #(
		.INIT('h8000)
	) name1571 (
		\a[0] ,
		\a[2] ,
		\a[36] ,
		\a[38] ,
		_w1637_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1572 (
		\a[0] ,
		\a[2] ,
		\a[36] ,
		\a[38] ,
		_w1638_
	);
	LUT2 #(
		.INIT('h6)
	) name1573 (
		_w1553_,
		_w1638_,
		_w1639_
	);
	LUT4 #(
		.INIT('h153f)
	) name1574 (
		\a[13] ,
		\a[14] ,
		\a[24] ,
		\a[25] ,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name1575 (
		\a[14] ,
		\a[25] ,
		_w1641_
	);
	LUT4 #(
		.INIT('h8000)
	) name1576 (
		\a[13] ,
		\a[14] ,
		\a[24] ,
		\a[25] ,
		_w1642_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1577 (
		\a[13] ,
		\a[14] ,
		\a[24] ,
		\a[25] ,
		_w1643_
	);
	LUT2 #(
		.INIT('h6)
	) name1578 (
		_w1525_,
		_w1643_,
		_w1644_
	);
	LUT3 #(
		.INIT('h69)
	) name1579 (
		_w1635_,
		_w1639_,
		_w1644_,
		_w1645_
	);
	LUT4 #(
		.INIT('h004d)
	) name1580 (
		_w1551_,
		_w1558_,
		_w1559_,
		_w1645_,
		_w1646_
	);
	LUT4 #(
		.INIT('hb200)
	) name1581 (
		_w1551_,
		_w1558_,
		_w1559_,
		_w1645_,
		_w1647_
	);
	LUT4 #(
		.INIT('h4db2)
	) name1582 (
		_w1551_,
		_w1558_,
		_w1559_,
		_w1645_,
		_w1648_
	);
	LUT2 #(
		.INIT('h6)
	) name1583 (
		_w1634_,
		_w1648_,
		_w1649_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1584 (
		_w1561_,
		_w1564_,
		_w1622_,
		_w1649_,
		_w1650_
	);
	LUT3 #(
		.INIT('h82)
	) name1585 (
		_w1620_,
		_w1634_,
		_w1648_,
		_w1651_
	);
	LUT4 #(
		.INIT('he800)
	) name1586 (
		_w1550_,
		_w1560_,
		_w1564_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h00e3)
	) name1587 (
		_w1621_,
		_w1623_,
		_w1649_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h6)
	) name1588 (
		_w1609_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name1589 (
		_w1578_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w1578_,
		_w1654_,
		_w1656_
	);
	LUT2 #(
		.INIT('h6)
	) name1591 (
		_w1578_,
		_w1654_,
		_w1657_
	);
	LUT3 #(
		.INIT('h51)
	) name1592 (
		_w1491_,
		_w1570_,
		_w1573_,
		_w1658_
	);
	LUT4 #(
		.INIT('h040f)
	) name1593 (
		_w1420_,
		_w1495_,
		_w1572_,
		_w1658_,
		_w1659_
	);
	LUT4 #(
		.INIT('he0ef)
	) name1594 (
		_w1574_,
		_w1577_,
		_w1657_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h2)
	) name1595 (
		_w1572_,
		_w1656_,
		_w1661_
	);
	LUT3 #(
		.INIT('h54)
	) name1596 (
		_w1491_,
		_w1578_,
		_w1654_,
		_w1662_
	);
	LUT4 #(
		.INIT('h040f)
	) name1597 (
		_w1420_,
		_w1495_,
		_w1661_,
		_w1662_,
		_w1663_
	);
	LUT3 #(
		.INIT('h54)
	) name1598 (
		_w1607_,
		_w1608_,
		_w1653_,
		_w1664_
	);
	LUT3 #(
		.INIT('h32)
	) name1599 (
		_w1634_,
		_w1646_,
		_w1647_,
		_w1665_
	);
	LUT3 #(
		.INIT('h45)
	) name1600 (
		_w1615_,
		_w1616_,
		_w1618_,
		_w1666_
	);
	LUT2 #(
		.INIT('h8)
	) name1601 (
		\a[0] ,
		\a[39] ,
		_w1667_
	);
	LUT3 #(
		.INIT('h93)
	) name1602 (
		\a[1] ,
		\a[20] ,
		\a[38] ,
		_w1668_
	);
	LUT3 #(
		.INIT('h69)
	) name1603 (
		_w1612_,
		_w1667_,
		_w1668_,
		_w1669_
	);
	LUT4 #(
		.INIT('h00d4)
	) name1604 (
		_w1613_,
		_w1614_,
		_w1618_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('h2b00)
	) name1605 (
		_w1613_,
		_w1614_,
		_w1618_,
		_w1669_,
		_w1671_
	);
	LUT4 #(
		.INIT('hba45)
	) name1606 (
		_w1615_,
		_w1616_,
		_w1618_,
		_w1669_,
		_w1672_
	);
	LUT3 #(
		.INIT('h17)
	) name1607 (
		_w1582_,
		_w1583_,
		_w1584_,
		_w1673_
	);
	LUT2 #(
		.INIT('h6)
	) name1608 (
		_w1672_,
		_w1673_,
		_w1674_
	);
	LUT3 #(
		.INIT('h32)
	) name1609 (
		_w1553_,
		_w1636_,
		_w1637_,
		_w1675_
	);
	LUT3 #(
		.INIT('h0d)
	) name1610 (
		_w1525_,
		_w1640_,
		_w1642_,
		_w1676_
	);
	LUT3 #(
		.INIT('h0d)
	) name1611 (
		_w1505_,
		_w1586_,
		_w1588_,
		_w1677_
	);
	LUT3 #(
		.INIT('h69)
	) name1612 (
		_w1675_,
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT3 #(
		.INIT('h32)
	) name1613 (
		_w1594_,
		_w1595_,
		_w1602_,
		_w1679_
	);
	LUT3 #(
		.INIT('hd4)
	) name1614 (
		_w1635_,
		_w1639_,
		_w1644_,
		_w1680_
	);
	LUT3 #(
		.INIT('h69)
	) name1615 (
		_w1678_,
		_w1679_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h6)
	) name1616 (
		_w1674_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h6)
	) name1617 (
		_w1665_,
		_w1682_,
		_w1683_
	);
	LUT3 #(
		.INIT('h01)
	) name1618 (
		_w1621_,
		_w1650_,
		_w1683_,
		_w1684_
	);
	LUT3 #(
		.INIT('he0)
	) name1619 (
		_w1621_,
		_w1650_,
		_w1683_,
		_w1685_
	);
	LUT3 #(
		.INIT('h1e)
	) name1620 (
		_w1621_,
		_w1650_,
		_w1683_,
		_w1686_
	);
	LUT3 #(
		.INIT('h51)
	) name1621 (
		_w1581_,
		_w1604_,
		_w1605_,
		_w1687_
	);
	LUT3 #(
		.INIT('h0d)
	) name1622 (
		_w1597_,
		_w1598_,
		_w1600_,
		_w1688_
	);
	LUT3 #(
		.INIT('h0d)
	) name1623 (
		_w1626_,
		_w1627_,
		_w1628_,
		_w1689_
	);
	LUT3 #(
		.INIT('h32)
	) name1624 (
		_w1590_,
		_w1591_,
		_w1592_,
		_w1690_
	);
	LUT3 #(
		.INIT('h96)
	) name1625 (
		_w1688_,
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h0e)
	) name1626 (
		_w1624_,
		_w1631_,
		_w1632_,
		_w1692_
	);
	LUT4 #(
		.INIT('h0017)
	) name1627 (
		_w1624_,
		_w1625_,
		_w1630_,
		_w1691_,
		_w1693_
	);
	LUT4 #(
		.INIT('he800)
	) name1628 (
		_w1624_,
		_w1625_,
		_w1630_,
		_w1691_,
		_w1694_
	);
	LUT4 #(
		.INIT('hf10e)
	) name1629 (
		_w1624_,
		_w1631_,
		_w1632_,
		_w1691_,
		_w1695_
	);
	LUT4 #(
		.INIT('h153f)
	) name1630 (
		\a[4] ,
		\a[12] ,
		\a[27] ,
		\a[35] ,
		_w1696_
	);
	LUT4 #(
		.INIT('h8000)
	) name1631 (
		\a[4] ,
		\a[12] ,
		\a[27] ,
		\a[35] ,
		_w1697_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1632 (
		\a[4] ,
		\a[12] ,
		\a[27] ,
		\a[35] ,
		_w1698_
	);
	LUT4 #(
		.INIT('h153f)
	) name1633 (
		\a[18] ,
		\a[19] ,
		\a[20] ,
		\a[21] ,
		_w1699_
	);
	LUT4 #(
		.INIT('h8000)
	) name1634 (
		\a[18] ,
		\a[19] ,
		\a[20] ,
		\a[21] ,
		_w1700_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1635 (
		\a[18] ,
		\a[19] ,
		\a[20] ,
		\a[21] ,
		_w1701_
	);
	LUT4 #(
		.INIT('h1248)
	) name1636 (
		_w1587_,
		_w1599_,
		_w1698_,
		_w1701_,
		_w1702_
	);
	LUT4 #(
		.INIT('h8421)
	) name1637 (
		_w1587_,
		_w1599_,
		_w1698_,
		_w1701_,
		_w1703_
	);
	LUT4 #(
		.INIT('h6996)
	) name1638 (
		_w1587_,
		_w1599_,
		_w1698_,
		_w1701_,
		_w1704_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		\a[11] ,
		\a[28] ,
		_w1705_
	);
	LUT4 #(
		.INIT('h153f)
	) name1640 (
		\a[5] ,
		\a[10] ,
		\a[29] ,
		\a[34] ,
		_w1706_
	);
	LUT4 #(
		.INIT('h8000)
	) name1641 (
		\a[5] ,
		\a[10] ,
		\a[29] ,
		\a[34] ,
		_w1707_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1642 (
		\a[5] ,
		\a[10] ,
		\a[29] ,
		\a[34] ,
		_w1708_
	);
	LUT2 #(
		.INIT('h6)
	) name1643 (
		_w1705_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h6)
	) name1644 (
		_w1704_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h6)
	) name1645 (
		_w1695_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('hae00)
	) name1646 (
		_w1581_,
		_w1604_,
		_w1605_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h153f)
	) name1647 (
		\a[15] ,
		\a[16] ,
		\a[23] ,
		\a[24] ,
		_w1713_
	);
	LUT4 #(
		.INIT('h8000)
	) name1648 (
		\a[15] ,
		\a[16] ,
		\a[23] ,
		\a[24] ,
		_w1714_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1649 (
		\a[15] ,
		\a[16] ,
		\a[23] ,
		\a[24] ,
		_w1715_
	);
	LUT2 #(
		.INIT('h8)
	) name1650 (
		\a[2] ,
		\a[37] ,
		_w1716_
	);
	LUT4 #(
		.INIT('h153f)
	) name1651 (
		\a[3] ,
		\a[13] ,
		\a[26] ,
		\a[36] ,
		_w1717_
	);
	LUT4 #(
		.INIT('h8000)
	) name1652 (
		\a[3] ,
		\a[13] ,
		\a[26] ,
		\a[36] ,
		_w1718_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1653 (
		\a[3] ,
		\a[13] ,
		\a[26] ,
		\a[36] ,
		_w1719_
	);
	LUT4 #(
		.INIT('h0660)
	) name1654 (
		_w1641_,
		_w1715_,
		_w1716_,
		_w1719_,
		_w1720_
	);
	LUT4 #(
		.INIT('h9009)
	) name1655 (
		_w1641_,
		_w1715_,
		_w1716_,
		_w1719_,
		_w1721_
	);
	LUT4 #(
		.INIT('h6996)
	) name1656 (
		_w1641_,
		_w1715_,
		_w1716_,
		_w1719_,
		_w1722_
	);
	LUT2 #(
		.INIT('h8)
	) name1657 (
		\a[7] ,
		\a[33] ,
		_w1723_
	);
	LUT4 #(
		.INIT('h8000)
	) name1658 (
		\a[6] ,
		\a[7] ,
		\a[32] ,
		\a[33] ,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		\a[6] ,
		\a[33] ,
		_w1725_
	);
	LUT4 #(
		.INIT('h8000)
	) name1660 (
		\a[6] ,
		\a[9] ,
		\a[30] ,
		\a[33] ,
		_w1726_
	);
	LUT4 #(
		.INIT('h8000)
	) name1661 (
		\a[7] ,
		\a[9] ,
		\a[30] ,
		\a[32] ,
		_w1727_
	);
	LUT3 #(
		.INIT('h0e)
	) name1662 (
		_w1724_,
		_w1726_,
		_w1727_,
		_w1728_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1663 (
		\a[7] ,
		\a[9] ,
		\a[30] ,
		\a[32] ,
		_w1729_
	);
	LUT2 #(
		.INIT('h1)
	) name1664 (
		_w1725_,
		_w1729_,
		_w1730_
	);
	LUT3 #(
		.INIT('ha9)
	) name1665 (
		_w1722_,
		_w1728_,
		_w1730_,
		_w1731_
	);
	LUT4 #(
		.INIT('h0071)
	) name1666 (
		_w1610_,
		_w1611_,
		_w1619_,
		_w1731_,
		_w1732_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1667 (
		_w1610_,
		_w1611_,
		_w1619_,
		_w1731_,
		_w1733_
	);
	LUT4 #(
		.INIT('h718e)
	) name1668 (
		_w1610_,
		_w1611_,
		_w1619_,
		_w1731_,
		_w1734_
	);
	LUT4 #(
		.INIT('hef0e)
	) name1669 (
		_w1520_,
		_w1522_,
		_w1585_,
		_w1603_,
		_w1735_
	);
	LUT2 #(
		.INIT('h6)
	) name1670 (
		_w1734_,
		_w1735_,
		_w1736_
	);
	LUT4 #(
		.INIT('h0051)
	) name1671 (
		_w1581_,
		_w1604_,
		_w1605_,
		_w1711_,
		_w1737_
	);
	LUT3 #(
		.INIT('h69)
	) name1672 (
		_w1687_,
		_w1711_,
		_w1736_,
		_w1738_
	);
	LUT2 #(
		.INIT('h6)
	) name1673 (
		_w1686_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h6)
	) name1674 (
		_w1664_,
		_w1739_,
		_w1740_
	);
	LUT4 #(
		.INIT('h32cd)
	) name1675 (
		_w1574_,
		_w1655_,
		_w1663_,
		_w1740_,
		_w1741_
	);
	LUT4 #(
		.INIT('h0777)
	) name1676 (
		_w1578_,
		_w1654_,
		_w1664_,
		_w1739_,
		_w1742_
	);
	LUT3 #(
		.INIT('h54)
	) name1677 (
		_w1684_,
		_w1685_,
		_w1738_,
		_w1743_
	);
	LUT3 #(
		.INIT('h54)
	) name1678 (
		_w1670_,
		_w1671_,
		_w1673_,
		_w1744_
	);
	LUT2 #(
		.INIT('h8)
	) name1679 (
		\a[18] ,
		\a[22] ,
		_w1745_
	);
	LUT4 #(
		.INIT('h153f)
	) name1680 (
		\a[0] ,
		\a[2] ,
		\a[38] ,
		\a[40] ,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1681 (
		\a[2] ,
		\a[40] ,
		_w1747_
	);
	LUT4 #(
		.INIT('h8000)
	) name1682 (
		\a[0] ,
		\a[2] ,
		\a[38] ,
		\a[40] ,
		_w1748_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1683 (
		\a[0] ,
		\a[2] ,
		\a[38] ,
		\a[40] ,
		_w1749_
	);
	LUT4 #(
		.INIT('h153f)
	) name1684 (
		\a[8] ,
		\a[9] ,
		\a[31] ,
		\a[32] ,
		_w1750_
	);
	LUT4 #(
		.INIT('h8000)
	) name1685 (
		\a[8] ,
		\a[9] ,
		\a[31] ,
		\a[32] ,
		_w1751_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1686 (
		\a[8] ,
		\a[9] ,
		\a[31] ,
		\a[32] ,
		_w1752_
	);
	LUT4 #(
		.INIT('h1428)
	) name1687 (
		_w1723_,
		_w1745_,
		_w1749_,
		_w1752_,
		_w1753_
	);
	LUT4 #(
		.INIT('h8241)
	) name1688 (
		_w1723_,
		_w1745_,
		_w1749_,
		_w1752_,
		_w1754_
	);
	LUT4 #(
		.INIT('h6996)
	) name1689 (
		_w1723_,
		_w1745_,
		_w1749_,
		_w1752_,
		_w1755_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		\a[4] ,
		\a[36] ,
		_w1756_
	);
	LUT4 #(
		.INIT('h153f)
	) name1691 (
		\a[5] ,
		\a[12] ,
		\a[28] ,
		\a[35] ,
		_w1757_
	);
	LUT4 #(
		.INIT('h8000)
	) name1692 (
		\a[5] ,
		\a[12] ,
		\a[28] ,
		\a[35] ,
		_w1758_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1693 (
		\a[5] ,
		\a[12] ,
		\a[28] ,
		\a[35] ,
		_w1759_
	);
	LUT2 #(
		.INIT('h6)
	) name1694 (
		_w1756_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h6)
	) name1695 (
		_w1755_,
		_w1760_,
		_w1761_
	);
	LUT3 #(
		.INIT('h01)
	) name1696 (
		_w1724_,
		_w1726_,
		_w1727_,
		_w1762_
	);
	LUT3 #(
		.INIT('h0d)
	) name1697 (
		_w1641_,
		_w1713_,
		_w1714_,
		_w1763_
	);
	LUT3 #(
		.INIT('h8e)
	) name1698 (
		_w1612_,
		_w1667_,
		_w1668_,
		_w1764_
	);
	LUT3 #(
		.INIT('h96)
	) name1699 (
		_w1762_,
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1700 (
		_w1666_,
		_w1669_,
		_w1673_,
		_w1765_,
		_w1766_
	);
	LUT4 #(
		.INIT('hed61)
	) name1701 (
		_w1744_,
		_w1761_,
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT4 #(
		.INIT('h1700)
	) name1702 (
		_w1665_,
		_w1674_,
		_w1681_,
		_w1767_,
		_w1768_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1703 (
		_w1665_,
		_w1674_,
		_w1681_,
		_w1767_,
		_w1769_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		\a[3] ,
		\a[37] ,
		_w1770_
	);
	LUT4 #(
		.INIT('h153f)
	) name1705 (
		\a[13] ,
		\a[14] ,
		\a[26] ,
		\a[27] ,
		_w1771_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		\a[14] ,
		\a[27] ,
		_w1772_
	);
	LUT4 #(
		.INIT('h8000)
	) name1707 (
		\a[13] ,
		\a[14] ,
		\a[26] ,
		\a[27] ,
		_w1773_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1708 (
		\a[13] ,
		\a[14] ,
		\a[26] ,
		\a[27] ,
		_w1774_
	);
	LUT2 #(
		.INIT('h8)
	) name1709 (
		\a[15] ,
		\a[25] ,
		_w1775_
	);
	LUT4 #(
		.INIT('h153f)
	) name1710 (
		\a[16] ,
		\a[17] ,
		\a[23] ,
		\a[24] ,
		_w1776_
	);
	LUT4 #(
		.INIT('h8000)
	) name1711 (
		\a[16] ,
		\a[17] ,
		\a[23] ,
		\a[24] ,
		_w1777_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1712 (
		\a[16] ,
		\a[17] ,
		\a[23] ,
		\a[24] ,
		_w1778_
	);
	LUT4 #(
		.INIT('h0660)
	) name1713 (
		_w1770_,
		_w1774_,
		_w1775_,
		_w1778_,
		_w1779_
	);
	LUT4 #(
		.INIT('h9009)
	) name1714 (
		_w1770_,
		_w1774_,
		_w1775_,
		_w1778_,
		_w1780_
	);
	LUT4 #(
		.INIT('h6996)
	) name1715 (
		_w1770_,
		_w1774_,
		_w1775_,
		_w1778_,
		_w1781_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		\a[11] ,
		\a[29] ,
		_w1782_
	);
	LUT4 #(
		.INIT('h153f)
	) name1717 (
		\a[6] ,
		\a[10] ,
		\a[30] ,
		\a[34] ,
		_w1783_
	);
	LUT4 #(
		.INIT('h8000)
	) name1718 (
		\a[6] ,
		\a[10] ,
		\a[30] ,
		\a[34] ,
		_w1784_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1719 (
		\a[6] ,
		\a[10] ,
		\a[30] ,
		\a[34] ,
		_w1785_
	);
	LUT2 #(
		.INIT('h6)
	) name1720 (
		_w1782_,
		_w1785_,
		_w1786_
	);
	LUT2 #(
		.INIT('h6)
	) name1721 (
		_w1781_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h002b)
	) name1722 (
		_w1678_,
		_w1679_,
		_w1680_,
		_w1787_,
		_w1788_
	);
	LUT4 #(
		.INIT('hd400)
	) name1723 (
		_w1678_,
		_w1679_,
		_w1680_,
		_w1787_,
		_w1789_
	);
	LUT3 #(
		.INIT('h71)
	) name1724 (
		_w1688_,
		_w1689_,
		_w1690_,
		_w1790_
	);
	LUT3 #(
		.INIT('h2b)
	) name1725 (
		_w1675_,
		_w1676_,
		_w1677_,
		_w1791_
	);
	LUT3 #(
		.INIT('h80)
	) name1726 (
		\a[1] ,
		\a[20] ,
		\a[38] ,
		_w1792_
	);
	LUT4 #(
		.INIT('h8000)
	) name1727 (
		\a[1] ,
		\a[19] ,
		\a[21] ,
		\a[39] ,
		_w1793_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1728 (
		\a[1] ,
		\a[19] ,
		\a[21] ,
		\a[39] ,
		_w1794_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		_w1792_,
		_w1794_,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name1730 (
		_w1792_,
		_w1794_,
		_w1796_
	);
	LUT2 #(
		.INIT('h6)
	) name1731 (
		_w1792_,
		_w1794_,
		_w1797_
	);
	LUT3 #(
		.INIT('h0d)
	) name1732 (
		_w1599_,
		_w1699_,
		_w1700_,
		_w1798_
	);
	LUT2 #(
		.INIT('h6)
	) name1733 (
		_w1797_,
		_w1798_,
		_w1799_
	);
	LUT3 #(
		.INIT('h69)
	) name1734 (
		_w1790_,
		_w1791_,
		_w1799_,
		_w1800_
	);
	LUT3 #(
		.INIT('he1)
	) name1735 (
		_w1788_,
		_w1789_,
		_w1800_,
		_w1801_
	);
	LUT3 #(
		.INIT('he1)
	) name1736 (
		_w1768_,
		_w1769_,
		_w1801_,
		_w1802_
	);
	LUT3 #(
		.INIT('h54)
	) name1737 (
		_w1732_,
		_w1733_,
		_w1735_,
		_w1803_
	);
	LUT3 #(
		.INIT('h54)
	) name1738 (
		_w1693_,
		_w1694_,
		_w1710_,
		_w1804_
	);
	LUT3 #(
		.INIT('h32)
	) name1739 (
		_w1587_,
		_w1696_,
		_w1697_,
		_w1805_
	);
	LUT3 #(
		.INIT('h32)
	) name1740 (
		_w1716_,
		_w1717_,
		_w1718_,
		_w1806_
	);
	LUT3 #(
		.INIT('h0d)
	) name1741 (
		_w1705_,
		_w1706_,
		_w1707_,
		_w1807_
	);
	LUT3 #(
		.INIT('h69)
	) name1742 (
		_w1805_,
		_w1806_,
		_w1807_,
		_w1808_
	);
	LUT3 #(
		.INIT('h32)
	) name1743 (
		_w1702_,
		_w1703_,
		_w1709_,
		_w1809_
	);
	LUT4 #(
		.INIT('h2223)
	) name1744 (
		_w1720_,
		_w1721_,
		_w1728_,
		_w1730_,
		_w1810_
	);
	LUT3 #(
		.INIT('h96)
	) name1745 (
		_w1808_,
		_w1809_,
		_w1810_,
		_w1811_
	);
	LUT4 #(
		.INIT('he800)
	) name1746 (
		_w1691_,
		_w1692_,
		_w1710_,
		_w1811_,
		_w1812_
	);
	LUT4 #(
		.INIT('h0017)
	) name1747 (
		_w1691_,
		_w1692_,
		_w1710_,
		_w1811_,
		_w1813_
	);
	LUT4 #(
		.INIT('hab54)
	) name1748 (
		_w1693_,
		_w1694_,
		_w1710_,
		_w1811_,
		_w1814_
	);
	LUT2 #(
		.INIT('h6)
	) name1749 (
		_w1803_,
		_w1814_,
		_w1815_
	);
	LUT4 #(
		.INIT('h2bff)
	) name1750 (
		_w1687_,
		_w1711_,
		_w1736_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h002b)
	) name1751 (
		_w1687_,
		_w1711_,
		_w1736_,
		_w1815_,
		_w1817_
	);
	LUT4 #(
		.INIT('h51ae)
	) name1752 (
		_w1712_,
		_w1736_,
		_w1737_,
		_w1815_,
		_w1818_
	);
	LUT2 #(
		.INIT('h9)
	) name1753 (
		_w1802_,
		_w1818_,
		_w1819_
	);
	LUT2 #(
		.INIT('h2)
	) name1754 (
		_w1743_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name1755 (
		_w1664_,
		_w1739_,
		_w1743_,
		_w1819_,
		_w1821_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1756 (
		_w1574_,
		_w1663_,
		_w1742_,
		_w1821_,
		_w1822_
	);
	LUT4 #(
		.INIT('hf00f)
	) name1757 (
		_w1664_,
		_w1739_,
		_w1743_,
		_w1819_,
		_w1823_
	);
	LUT4 #(
		.INIT('he000)
	) name1758 (
		_w1574_,
		_w1663_,
		_w1742_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('he)
	) name1759 (
		_w1822_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h2)
	) name1760 (
		_w1742_,
		_w1820_,
		_w1826_
	);
	LUT4 #(
		.INIT('h1101)
	) name1761 (
		_w1664_,
		_w1739_,
		_w1743_,
		_w1819_,
		_w1827_
	);
	LUT3 #(
		.INIT('h0b)
	) name1762 (
		_w1802_,
		_w1816_,
		_w1817_,
		_w1828_
	);
	LUT3 #(
		.INIT('h54)
	) name1763 (
		_w1788_,
		_w1789_,
		_w1800_,
		_w1829_
	);
	LUT2 #(
		.INIT('h2)
	) name1764 (
		_w1761_,
		_w1765_,
		_w1830_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w1761_,
		_w1765_,
		_w1831_
	);
	LUT4 #(
		.INIT('he800)
	) name1766 (
		_w1666_,
		_w1669_,
		_w1673_,
		_w1765_,
		_w1832_
	);
	LUT4 #(
		.INIT('h0027)
	) name1767 (
		_w1744_,
		_w1830_,
		_w1831_,
		_w1832_,
		_w1833_
	);
	LUT3 #(
		.INIT('h0d)
	) name1768 (
		_w1775_,
		_w1776_,
		_w1777_,
		_w1834_
	);
	LUT3 #(
		.INIT('h0d)
	) name1769 (
		_w1745_,
		_w1746_,
		_w1748_,
		_w1835_
	);
	LUT3 #(
		.INIT('h0d)
	) name1770 (
		_w1770_,
		_w1771_,
		_w1773_,
		_w1836_
	);
	LUT3 #(
		.INIT('h96)
	) name1771 (
		_w1834_,
		_w1835_,
		_w1836_,
		_w1837_
	);
	LUT3 #(
		.INIT('h32)
	) name1772 (
		_w1753_,
		_w1754_,
		_w1760_,
		_w1838_
	);
	LUT3 #(
		.INIT('h80)
	) name1773 (
		\a[1] ,
		\a[21] ,
		\a[40] ,
		_w1839_
	);
	LUT3 #(
		.INIT('h6c)
	) name1774 (
		\a[1] ,
		\a[21] ,
		\a[40] ,
		_w1840_
	);
	LUT4 #(
		.INIT('h000d)
	) name1775 (
		_w1723_,
		_w1750_,
		_w1751_,
		_w1840_,
		_w1841_
	);
	LUT4 #(
		.INIT('hf200)
	) name1776 (
		_w1723_,
		_w1750_,
		_w1751_,
		_w1840_,
		_w1842_
	);
	LUT4 #(
		.INIT('h0df2)
	) name1777 (
		_w1723_,
		_w1750_,
		_w1751_,
		_w1840_,
		_w1843_
	);
	LUT3 #(
		.INIT('h32)
	) name1778 (
		_w1782_,
		_w1783_,
		_w1784_,
		_w1844_
	);
	LUT2 #(
		.INIT('h6)
	) name1779 (
		_w1843_,
		_w1844_,
		_w1845_
	);
	LUT3 #(
		.INIT('h69)
	) name1780 (
		_w1837_,
		_w1838_,
		_w1845_,
		_w1846_
	);
	LUT3 #(
		.INIT('h69)
	) name1781 (
		_w1829_,
		_w1833_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1782 (
		_w1768_,
		_w1769_,
		_w1801_,
		_w1847_,
		_w1848_
	);
	LUT4 #(
		.INIT('h5400)
	) name1783 (
		_w1768_,
		_w1769_,
		_w1801_,
		_w1847_,
		_w1849_
	);
	LUT4 #(
		.INIT('hab54)
	) name1784 (
		_w1768_,
		_w1769_,
		_w1801_,
		_w1847_,
		_w1850_
	);
	LUT3 #(
		.INIT('h8e)
	) name1785 (
		_w1790_,
		_w1791_,
		_w1799_,
		_w1851_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		\a[5] ,
		\a[36] ,
		_w1852_
	);
	LUT4 #(
		.INIT('h153f)
	) name1787 (
		\a[6] ,
		\a[11] ,
		\a[30] ,
		\a[35] ,
		_w1853_
	);
	LUT4 #(
		.INIT('h8000)
	) name1788 (
		\a[6] ,
		\a[11] ,
		\a[30] ,
		\a[35] ,
		_w1854_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1789 (
		\a[6] ,
		\a[11] ,
		\a[30] ,
		\a[35] ,
		_w1855_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		\a[8] ,
		\a[33] ,
		_w1856_
	);
	LUT4 #(
		.INIT('h153f)
	) name1791 (
		\a[19] ,
		\a[20] ,
		\a[21] ,
		\a[22] ,
		_w1857_
	);
	LUT4 #(
		.INIT('h8000)
	) name1792 (
		\a[19] ,
		\a[20] ,
		\a[21] ,
		\a[22] ,
		_w1858_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1793 (
		\a[19] ,
		\a[20] ,
		\a[21] ,
		\a[22] ,
		_w1859_
	);
	LUT4 #(
		.INIT('h0660)
	) name1794 (
		_w1852_,
		_w1855_,
		_w1856_,
		_w1859_,
		_w1860_
	);
	LUT4 #(
		.INIT('h9009)
	) name1795 (
		_w1852_,
		_w1855_,
		_w1856_,
		_w1859_,
		_w1861_
	);
	LUT4 #(
		.INIT('h6996)
	) name1796 (
		_w1852_,
		_w1855_,
		_w1856_,
		_w1859_,
		_w1862_
	);
	LUT4 #(
		.INIT('hdc23)
	) name1797 (
		_w1795_,
		_w1796_,
		_w1798_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		\a[16] ,
		\a[25] ,
		_w1864_
	);
	LUT4 #(
		.INIT('h153f)
	) name1799 (
		\a[17] ,
		\a[18] ,
		\a[23] ,
		\a[24] ,
		_w1865_
	);
	LUT4 #(
		.INIT('h8000)
	) name1800 (
		\a[17] ,
		\a[18] ,
		\a[23] ,
		\a[24] ,
		_w1866_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1801 (
		\a[17] ,
		\a[18] ,
		\a[23] ,
		\a[24] ,
		_w1867_
	);
	LUT4 #(
		.INIT('h153f)
	) name1802 (
		\a[4] ,
		\a[12] ,
		\a[29] ,
		\a[37] ,
		_w1868_
	);
	LUT4 #(
		.INIT('h8000)
	) name1803 (
		\a[4] ,
		\a[12] ,
		\a[29] ,
		\a[37] ,
		_w1869_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1804 (
		\a[4] ,
		\a[12] ,
		\a[29] ,
		\a[37] ,
		_w1870_
	);
	LUT4 #(
		.INIT('h1428)
	) name1805 (
		_w1772_,
		_w1864_,
		_w1867_,
		_w1870_,
		_w1871_
	);
	LUT4 #(
		.INIT('h8241)
	) name1806 (
		_w1772_,
		_w1864_,
		_w1867_,
		_w1870_,
		_w1872_
	);
	LUT4 #(
		.INIT('h6996)
	) name1807 (
		_w1772_,
		_w1864_,
		_w1867_,
		_w1870_,
		_w1873_
	);
	LUT2 #(
		.INIT('h8)
	) name1808 (
		\a[10] ,
		\a[31] ,
		_w1874_
	);
	LUT4 #(
		.INIT('h153f)
	) name1809 (
		\a[7] ,
		\a[9] ,
		\a[32] ,
		\a[34] ,
		_w1875_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		\a[9] ,
		\a[34] ,
		_w1876_
	);
	LUT4 #(
		.INIT('h8000)
	) name1811 (
		\a[7] ,
		\a[9] ,
		\a[32] ,
		\a[34] ,
		_w1877_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1812 (
		\a[7] ,
		\a[9] ,
		\a[32] ,
		\a[34] ,
		_w1878_
	);
	LUT2 #(
		.INIT('h6)
	) name1813 (
		_w1874_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h6)
	) name1814 (
		_w1873_,
		_w1879_,
		_w1880_
	);
	LUT3 #(
		.INIT('h96)
	) name1815 (
		_w1851_,
		_w1863_,
		_w1880_,
		_w1881_
	);
	LUT4 #(
		.INIT('he800)
	) name1816 (
		_w1803_,
		_w1804_,
		_w1811_,
		_w1881_,
		_w1882_
	);
	LUT3 #(
		.INIT('h71)
	) name1817 (
		_w1762_,
		_w1763_,
		_w1764_,
		_w1883_
	);
	LUT3 #(
		.INIT('h8e)
	) name1818 (
		_w1805_,
		_w1806_,
		_w1807_,
		_w1884_
	);
	LUT3 #(
		.INIT('h32)
	) name1819 (
		_w1779_,
		_w1780_,
		_w1786_,
		_w1885_
	);
	LUT3 #(
		.INIT('h96)
	) name1820 (
		_w1883_,
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h8)
	) name1821 (
		\a[2] ,
		\a[41] ,
		_w1887_
	);
	LUT4 #(
		.INIT('h8000)
	) name1822 (
		\a[0] ,
		\a[2] ,
		\a[39] ,
		\a[41] ,
		_w1888_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1823 (
		\a[0] ,
		\a[2] ,
		\a[39] ,
		\a[41] ,
		_w1889_
	);
	LUT2 #(
		.INIT('h6)
	) name1824 (
		_w1793_,
		_w1889_,
		_w1890_
	);
	LUT3 #(
		.INIT('h32)
	) name1825 (
		_w1756_,
		_w1757_,
		_w1758_,
		_w1891_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		\a[3] ,
		\a[38] ,
		_w1892_
	);
	LUT4 #(
		.INIT('h153f)
	) name1827 (
		\a[13] ,
		\a[15] ,
		\a[26] ,
		\a[28] ,
		_w1893_
	);
	LUT4 #(
		.INIT('h8000)
	) name1828 (
		\a[13] ,
		\a[15] ,
		\a[26] ,
		\a[28] ,
		_w1894_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1829 (
		\a[13] ,
		\a[15] ,
		\a[26] ,
		\a[28] ,
		_w1895_
	);
	LUT2 #(
		.INIT('h6)
	) name1830 (
		_w1892_,
		_w1895_,
		_w1896_
	);
	LUT3 #(
		.INIT('h96)
	) name1831 (
		_w1890_,
		_w1891_,
		_w1896_,
		_w1897_
	);
	LUT4 #(
		.INIT('he800)
	) name1832 (
		_w1808_,
		_w1809_,
		_w1810_,
		_w1897_,
		_w1898_
	);
	LUT4 #(
		.INIT('h0017)
	) name1833 (
		_w1808_,
		_w1809_,
		_w1810_,
		_w1897_,
		_w1899_
	);
	LUT3 #(
		.INIT('ha9)
	) name1834 (
		_w1886_,
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT4 #(
		.INIT('h0031)
	) name1835 (
		_w1803_,
		_w1812_,
		_w1813_,
		_w1881_,
		_w1901_
	);
	LUT3 #(
		.INIT('h04)
	) name1836 (
		_w1882_,
		_w1900_,
		_w1901_,
		_w1902_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1837 (
		_w1803_,
		_w1804_,
		_w1811_,
		_w1881_,
		_w1903_
	);
	LUT4 #(
		.INIT('h3100)
	) name1838 (
		_w1803_,
		_w1812_,
		_w1813_,
		_w1881_,
		_w1904_
	);
	LUT3 #(
		.INIT('h01)
	) name1839 (
		_w1900_,
		_w1903_,
		_w1904_,
		_w1905_
	);
	LUT3 #(
		.INIT('ha9)
	) name1840 (
		_w1850_,
		_w1902_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h8)
	) name1841 (
		_w1828_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h6)
	) name1842 (
		_w1828_,
		_w1906_,
		_w1908_
	);
	LUT4 #(
		.INIT('h0bb0)
	) name1843 (
		_w1743_,
		_w1819_,
		_w1828_,
		_w1906_,
		_w1909_
	);
	LUT2 #(
		.INIT('h4)
	) name1844 (
		_w1827_,
		_w1909_,
		_w1910_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1845 (
		_w1574_,
		_w1663_,
		_w1826_,
		_w1910_,
		_w1911_
	);
	LUT4 #(
		.INIT('he0fe)
	) name1846 (
		_w1664_,
		_w1739_,
		_w1743_,
		_w1819_,
		_w1912_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1847 (
		_w1574_,
		_w1663_,
		_w1826_,
		_w1912_,
		_w1913_
	);
	LUT3 #(
		.INIT('h32)
	) name1848 (
		_w1908_,
		_w1911_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name1849 (
		_w1743_,
		_w1819_,
		_w1828_,
		_w1906_,
		_w1915_
	);
	LUT2 #(
		.INIT('h4)
	) name1850 (
		_w1827_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1851 (
		_w1574_,
		_w1663_,
		_w1826_,
		_w1916_,
		_w1917_
	);
	LUT3 #(
		.INIT('h0e)
	) name1852 (
		_w1886_,
		_w1898_,
		_w1899_,
		_w1918_
	);
	LUT3 #(
		.INIT('h17)
	) name1853 (
		_w1834_,
		_w1835_,
		_w1836_,
		_w1919_
	);
	LUT3 #(
		.INIT('he8)
	) name1854 (
		_w1890_,
		_w1891_,
		_w1896_,
		_w1920_
	);
	LUT3 #(
		.INIT('h32)
	) name1855 (
		_w1871_,
		_w1872_,
		_w1879_,
		_w1921_
	);
	LUT3 #(
		.INIT('h96)
	) name1856 (
		_w1919_,
		_w1920_,
		_w1921_,
		_w1922_
	);
	LUT3 #(
		.INIT('h17)
	) name1857 (
		_w1851_,
		_w1863_,
		_w1880_,
		_w1923_
	);
	LUT4 #(
		.INIT('he800)
	) name1858 (
		_w1851_,
		_w1863_,
		_w1880_,
		_w1922_,
		_w1924_
	);
	LUT4 #(
		.INIT('h0017)
	) name1859 (
		_w1851_,
		_w1863_,
		_w1880_,
		_w1922_,
		_w1925_
	);
	LUT4 #(
		.INIT('h17e8)
	) name1860 (
		_w1851_,
		_w1863_,
		_w1880_,
		_w1922_,
		_w1926_
	);
	LUT2 #(
		.INIT('h6)
	) name1861 (
		_w1918_,
		_w1926_,
		_w1927_
	);
	LUT4 #(
		.INIT('hae00)
	) name1862 (
		_w1882_,
		_w1900_,
		_w1901_,
		_w1927_,
		_w1928_
	);
	LUT4 #(
		.INIT('h0051)
	) name1863 (
		_w1882_,
		_w1900_,
		_w1901_,
		_w1927_,
		_w1929_
	);
	LUT4 #(
		.INIT('h51ae)
	) name1864 (
		_w1882_,
		_w1900_,
		_w1901_,
		_w1927_,
		_w1930_
	);
	LUT3 #(
		.INIT('hb2)
	) name1865 (
		_w1829_,
		_w1833_,
		_w1846_,
		_w1931_
	);
	LUT3 #(
		.INIT('h54)
	) name1866 (
		_w1841_,
		_w1842_,
		_w1844_,
		_w1932_
	);
	LUT4 #(
		.INIT('h8000)
	) name1867 (
		\a[1] ,
		\a[20] ,
		\a[22] ,
		\a[41] ,
		_w1933_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1868 (
		\a[1] ,
		\a[20] ,
		\a[22] ,
		\a[41] ,
		_w1934_
	);
	LUT2 #(
		.INIT('h8)
	) name1869 (
		\a[0] ,
		\a[42] ,
		_w1935_
	);
	LUT3 #(
		.INIT('h96)
	) name1870 (
		_w1839_,
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		\a[13] ,
		\a[29] ,
		_w1937_
	);
	LUT4 #(
		.INIT('h153f)
	) name1872 (
		\a[5] ,
		\a[12] ,
		\a[30] ,
		\a[37] ,
		_w1938_
	);
	LUT4 #(
		.INIT('h8000)
	) name1873 (
		\a[5] ,
		\a[12] ,
		\a[30] ,
		\a[37] ,
		_w1939_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1874 (
		\a[5] ,
		\a[12] ,
		\a[30] ,
		\a[37] ,
		_w1940_
	);
	LUT2 #(
		.INIT('h6)
	) name1875 (
		_w1937_,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		_w1936_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w1936_,
		_w1941_,
		_w1943_
	);
	LUT2 #(
		.INIT('h6)
	) name1878 (
		_w1936_,
		_w1941_,
		_w1944_
	);
	LUT2 #(
		.INIT('h6)
	) name1879 (
		_w1932_,
		_w1944_,
		_w1945_
	);
	LUT3 #(
		.INIT('hd4)
	) name1880 (
		_w1837_,
		_w1838_,
		_w1845_,
		_w1946_
	);
	LUT3 #(
		.INIT('h32)
	) name1881 (
		_w1856_,
		_w1857_,
		_w1858_,
		_w1947_
	);
	LUT3 #(
		.INIT('h32)
	) name1882 (
		_w1772_,
		_w1868_,
		_w1869_,
		_w1948_
	);
	LUT3 #(
		.INIT('h0d)
	) name1883 (
		_w1852_,
		_w1853_,
		_w1854_,
		_w1949_
	);
	LUT3 #(
		.INIT('h96)
	) name1884 (
		_w1947_,
		_w1948_,
		_w1949_,
		_w1950_
	);
	LUT4 #(
		.INIT('h0071)
	) name1885 (
		_w1792_,
		_w1794_,
		_w1798_,
		_w1860_,
		_w1951_
	);
	LUT3 #(
		.INIT('h0d)
	) name1886 (
		_w1892_,
		_w1893_,
		_w1894_,
		_w1952_
	);
	LUT3 #(
		.INIT('h0d)
	) name1887 (
		_w1864_,
		_w1865_,
		_w1866_,
		_w1953_
	);
	LUT4 #(
		.INIT('h153f)
	) name1888 (
		\a[0] ,
		\a[2] ,
		\a[39] ,
		\a[41] ,
		_w1954_
	);
	LUT3 #(
		.INIT('h0e)
	) name1889 (
		_w1793_,
		_w1888_,
		_w1954_,
		_w1955_
	);
	LUT3 #(
		.INIT('h96)
	) name1890 (
		_w1952_,
		_w1953_,
		_w1955_,
		_w1956_
	);
	LUT4 #(
		.INIT('hc936)
	) name1891 (
		_w1861_,
		_w1950_,
		_w1951_,
		_w1956_,
		_w1957_
	);
	LUT3 #(
		.INIT('h96)
	) name1892 (
		_w1945_,
		_w1946_,
		_w1957_,
		_w1958_
	);
	LUT3 #(
		.INIT('he8)
	) name1893 (
		_w1883_,
		_w1884_,
		_w1885_,
		_w1959_
	);
	LUT2 #(
		.INIT('h8)
	) name1894 (
		\a[17] ,
		\a[25] ,
		_w1960_
	);
	LUT4 #(
		.INIT('h153f)
	) name1895 (
		\a[18] ,
		\a[19] ,
		\a[23] ,
		\a[24] ,
		_w1961_
	);
	LUT4 #(
		.INIT('h8000)
	) name1896 (
		\a[18] ,
		\a[19] ,
		\a[23] ,
		\a[24] ,
		_w1962_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1897 (
		\a[18] ,
		\a[19] ,
		\a[23] ,
		\a[24] ,
		_w1963_
	);
	LUT4 #(
		.INIT('h153f)
	) name1898 (
		\a[3] ,
		\a[16] ,
		\a[26] ,
		\a[39] ,
		_w1964_
	);
	LUT4 #(
		.INIT('h8000)
	) name1899 (
		\a[3] ,
		\a[16] ,
		\a[26] ,
		\a[39] ,
		_w1965_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1900 (
		\a[3] ,
		\a[16] ,
		\a[26] ,
		\a[39] ,
		_w1966_
	);
	LUT4 #(
		.INIT('h1428)
	) name1901 (
		_w1747_,
		_w1960_,
		_w1963_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h8241)
	) name1902 (
		_w1747_,
		_w1960_,
		_w1963_,
		_w1966_,
		_w1968_
	);
	LUT4 #(
		.INIT('h6996)
	) name1903 (
		_w1747_,
		_w1960_,
		_w1963_,
		_w1966_,
		_w1969_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		\a[15] ,
		\a[27] ,
		_w1970_
	);
	LUT4 #(
		.INIT('h153f)
	) name1905 (
		\a[4] ,
		\a[14] ,
		\a[28] ,
		\a[38] ,
		_w1971_
	);
	LUT2 #(
		.INIT('h8)
	) name1906 (
		\a[14] ,
		\a[38] ,
		_w1972_
	);
	LUT4 #(
		.INIT('h8000)
	) name1907 (
		\a[4] ,
		\a[14] ,
		\a[28] ,
		\a[38] ,
		_w1973_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1908 (
		\a[4] ,
		\a[14] ,
		\a[28] ,
		\a[38] ,
		_w1974_
	);
	LUT2 #(
		.INIT('h6)
	) name1909 (
		_w1970_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h1)
	) name1910 (
		_w1969_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w1969_,
		_w1975_,
		_w1977_
	);
	LUT2 #(
		.INIT('h6)
	) name1912 (
		_w1969_,
		_w1975_,
		_w1978_
	);
	LUT3 #(
		.INIT('h0d)
	) name1913 (
		_w1874_,
		_w1875_,
		_w1877_,
		_w1979_
	);
	LUT2 #(
		.INIT('h8)
	) name1914 (
		\a[6] ,
		\a[36] ,
		_w1980_
	);
	LUT4 #(
		.INIT('h153f)
	) name1915 (
		\a[7] ,
		\a[11] ,
		\a[31] ,
		\a[35] ,
		_w1981_
	);
	LUT4 #(
		.INIT('h8000)
	) name1916 (
		\a[7] ,
		\a[11] ,
		\a[31] ,
		\a[35] ,
		_w1982_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1917 (
		\a[7] ,
		\a[11] ,
		\a[31] ,
		\a[35] ,
		_w1983_
	);
	LUT2 #(
		.INIT('h6)
	) name1918 (
		_w1980_,
		_w1983_,
		_w1984_
	);
	LUT4 #(
		.INIT('h153f)
	) name1919 (
		\a[8] ,
		\a[9] ,
		\a[33] ,
		\a[34] ,
		_w1985_
	);
	LUT4 #(
		.INIT('h8000)
	) name1920 (
		\a[8] ,
		\a[9] ,
		\a[33] ,
		\a[34] ,
		_w1986_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1921 (
		\a[8] ,
		\a[9] ,
		\a[33] ,
		\a[34] ,
		_w1987_
	);
	LUT2 #(
		.INIT('h6)
	) name1922 (
		_w1514_,
		_w1987_,
		_w1988_
	);
	LUT3 #(
		.INIT('h69)
	) name1923 (
		_w1979_,
		_w1984_,
		_w1988_,
		_w1989_
	);
	LUT3 #(
		.INIT('h69)
	) name1924 (
		_w1959_,
		_w1978_,
		_w1989_,
		_w1990_
	);
	LUT3 #(
		.INIT('h7b)
	) name1925 (
		_w1931_,
		_w1958_,
		_w1990_,
		_w1991_
	);
	LUT3 #(
		.INIT('h69)
	) name1926 (
		_w1931_,
		_w1958_,
		_w1990_,
		_w1992_
	);
	LUT2 #(
		.INIT('h1)
	) name1927 (
		_w1930_,
		_w1992_,
		_w1993_
	);
	LUT4 #(
		.INIT('h4445)
	) name1928 (
		_w1848_,
		_w1849_,
		_w1902_,
		_w1905_,
		_w1994_
	);
	LUT3 #(
		.INIT('h10)
	) name1929 (
		_w1928_,
		_w1929_,
		_w1992_,
		_w1995_
	);
	LUT3 #(
		.INIT('h04)
	) name1930 (
		_w1993_,
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT3 #(
		.INIT('he1)
	) name1931 (
		_w1928_,
		_w1929_,
		_w1992_,
		_w1997_
	);
	LUT2 #(
		.INIT('h1)
	) name1932 (
		_w1994_,
		_w1997_,
		_w1998_
	);
	LUT3 #(
		.INIT('hc9)
	) name1933 (
		_w1993_,
		_w1994_,
		_w1995_,
		_w1999_
	);
	LUT3 #(
		.INIT('h1e)
	) name1934 (
		_w1907_,
		_w1917_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w1907_,
		_w1996_,
		_w2001_
	);
	LUT3 #(
		.INIT('h45)
	) name1936 (
		_w1928_,
		_w1929_,
		_w1992_,
		_w2002_
	);
	LUT4 #(
		.INIT('h00b2)
	) name1937 (
		_w1829_,
		_w1833_,
		_w1846_,
		_w1990_,
		_w2003_
	);
	LUT3 #(
		.INIT('he8)
	) name1938 (
		_w1945_,
		_w1946_,
		_w1957_,
		_w2004_
	);
	LUT4 #(
		.INIT('he800)
	) name1939 (
		_w1883_,
		_w1884_,
		_w1885_,
		_w1989_,
		_w2005_
	);
	LUT2 #(
		.INIT('h4)
	) name1940 (
		_w1976_,
		_w1989_,
		_w2006_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1941 (
		_w1883_,
		_w1884_,
		_w1885_,
		_w1976_,
		_w2007_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1942 (
		_w1977_,
		_w2005_,
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT3 #(
		.INIT('hd4)
	) name1943 (
		_w1979_,
		_w1984_,
		_w1988_,
		_w2009_
	);
	LUT3 #(
		.INIT('h80)
	) name1944 (
		\a[1] ,
		\a[22] ,
		\a[42] ,
		_w2010_
	);
	LUT3 #(
		.INIT('h6c)
	) name1945 (
		\a[1] ,
		\a[22] ,
		\a[42] ,
		_w2011_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w1933_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h4)
	) name1947 (
		\a[42] ,
		_w1933_,
		_w2013_
	);
	LUT3 #(
		.INIT('hb8)
	) name1948 (
		\a[42] ,
		_w1933_,
		_w2011_,
		_w2014_
	);
	LUT3 #(
		.INIT('h0d)
	) name1949 (
		_w1514_,
		_w1985_,
		_w1986_,
		_w2015_
	);
	LUT2 #(
		.INIT('h6)
	) name1950 (
		_w2014_,
		_w2015_,
		_w2016_
	);
	LUT3 #(
		.INIT('h32)
	) name1951 (
		_w1967_,
		_w1968_,
		_w1975_,
		_w2017_
	);
	LUT3 #(
		.INIT('h69)
	) name1952 (
		_w2009_,
		_w2016_,
		_w2017_,
		_w2018_
	);
	LUT3 #(
		.INIT('h96)
	) name1953 (
		_w2004_,
		_w2008_,
		_w2018_,
		_w2019_
	);
	LUT3 #(
		.INIT('h0e)
	) name1954 (
		_w1918_,
		_w1924_,
		_w1925_,
		_w2020_
	);
	LUT2 #(
		.INIT('h8)
	) name1955 (
		\a[14] ,
		\a[29] ,
		_w2021_
	);
	LUT4 #(
		.INIT('h153f)
	) name1956 (
		\a[15] ,
		\a[16] ,
		\a[27] ,
		\a[28] ,
		_w2022_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		\a[16] ,
		\a[28] ,
		_w2023_
	);
	LUT4 #(
		.INIT('h8000)
	) name1958 (
		\a[15] ,
		\a[16] ,
		\a[27] ,
		\a[28] ,
		_w2024_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1959 (
		\a[15] ,
		\a[16] ,
		\a[27] ,
		\a[28] ,
		_w2025_
	);
	LUT2 #(
		.INIT('h8)
	) name1960 (
		\a[4] ,
		\a[39] ,
		_w2026_
	);
	LUT4 #(
		.INIT('h153f)
	) name1961 (
		\a[0] ,
		\a[3] ,
		\a[40] ,
		\a[43] ,
		_w2027_
	);
	LUT4 #(
		.INIT('h8000)
	) name1962 (
		\a[0] ,
		\a[3] ,
		\a[40] ,
		\a[43] ,
		_w2028_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1963 (
		\a[0] ,
		\a[3] ,
		\a[40] ,
		\a[43] ,
		_w2029_
	);
	LUT4 #(
		.INIT('h0660)
	) name1964 (
		_w2021_,
		_w2025_,
		_w2026_,
		_w2029_,
		_w2030_
	);
	LUT4 #(
		.INIT('h9009)
	) name1965 (
		_w2021_,
		_w2025_,
		_w2026_,
		_w2029_,
		_w2031_
	);
	LUT4 #(
		.INIT('h6996)
	) name1966 (
		_w2021_,
		_w2025_,
		_w2026_,
		_w2029_,
		_w2032_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		\a[17] ,
		\a[26] ,
		_w2033_
	);
	LUT4 #(
		.INIT('h153f)
	) name1968 (
		\a[18] ,
		\a[19] ,
		\a[24] ,
		\a[25] ,
		_w2034_
	);
	LUT4 #(
		.INIT('h8000)
	) name1969 (
		\a[18] ,
		\a[19] ,
		\a[24] ,
		\a[25] ,
		_w2035_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1970 (
		\a[18] ,
		\a[19] ,
		\a[24] ,
		\a[25] ,
		_w2036_
	);
	LUT2 #(
		.INIT('h6)
	) name1971 (
		_w2033_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h8)
	) name1972 (
		\a[7] ,
		\a[36] ,
		_w2038_
	);
	LUT4 #(
		.INIT('h153f)
	) name1973 (
		\a[8] ,
		\a[10] ,
		\a[33] ,
		\a[35] ,
		_w2039_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		\a[10] ,
		\a[35] ,
		_w2040_
	);
	LUT4 #(
		.INIT('h8000)
	) name1975 (
		\a[8] ,
		\a[10] ,
		\a[33] ,
		\a[35] ,
		_w2041_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1976 (
		\a[8] ,
		\a[10] ,
		\a[33] ,
		\a[35] ,
		_w2042_
	);
	LUT4 #(
		.INIT('h153f)
	) name1977 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w2043_
	);
	LUT4 #(
		.INIT('h8000)
	) name1978 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w2044_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1979 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w2045_
	);
	LUT4 #(
		.INIT('h1428)
	) name1980 (
		_w1876_,
		_w2038_,
		_w2042_,
		_w2045_,
		_w2046_
	);
	LUT4 #(
		.INIT('h8241)
	) name1981 (
		_w1876_,
		_w2038_,
		_w2042_,
		_w2045_,
		_w2047_
	);
	LUT4 #(
		.INIT('h6996)
	) name1982 (
		_w1876_,
		_w2038_,
		_w2042_,
		_w2045_,
		_w2048_
	);
	LUT4 #(
		.INIT('h153f)
	) name1983 (
		\a[5] ,
		\a[13] ,
		\a[30] ,
		\a[38] ,
		_w2049_
	);
	LUT4 #(
		.INIT('h8000)
	) name1984 (
		\a[5] ,
		\a[13] ,
		\a[30] ,
		\a[38] ,
		_w2050_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name1985 (
		\a[5] ,
		\a[13] ,
		\a[30] ,
		\a[38] ,
		_w2051_
	);
	LUT2 #(
		.INIT('h6)
	) name1986 (
		_w1887_,
		_w2051_,
		_w2052_
	);
	LUT4 #(
		.INIT('h0660)
	) name1987 (
		_w2032_,
		_w2037_,
		_w2048_,
		_w2052_,
		_w2053_
	);
	LUT4 #(
		.INIT('h6996)
	) name1988 (
		_w2032_,
		_w2037_,
		_w2048_,
		_w2052_,
		_w2054_
	);
	LUT4 #(
		.INIT('he800)
	) name1989 (
		_w1919_,
		_w1920_,
		_w1921_,
		_w2054_,
		_w2055_
	);
	LUT4 #(
		.INIT('h17e8)
	) name1990 (
		_w1919_,
		_w1920_,
		_w1921_,
		_w2054_,
		_w2056_
	);
	LUT3 #(
		.INIT('h0e)
	) name1991 (
		_w1932_,
		_w1942_,
		_w1943_,
		_w2057_
	);
	LUT3 #(
		.INIT('h32)
	) name1992 (
		_w1980_,
		_w1981_,
		_w1982_,
		_w2058_
	);
	LUT3 #(
		.INIT('h0d)
	) name1993 (
		_w1970_,
		_w1971_,
		_w1973_,
		_w2059_
	);
	LUT3 #(
		.INIT('h0d)
	) name1994 (
		_w1960_,
		_w1961_,
		_w1962_,
		_w2060_
	);
	LUT3 #(
		.INIT('h69)
	) name1995 (
		_w2058_,
		_w2059_,
		_w2060_,
		_w2061_
	);
	LUT3 #(
		.INIT('h32)
	) name1996 (
		_w1937_,
		_w1938_,
		_w1939_,
		_w2062_
	);
	LUT3 #(
		.INIT('h32)
	) name1997 (
		_w1747_,
		_w1964_,
		_w1965_,
		_w2063_
	);
	LUT3 #(
		.INIT('he8)
	) name1998 (
		_w1839_,
		_w1934_,
		_w1935_,
		_w2064_
	);
	LUT3 #(
		.INIT('h96)
	) name1999 (
		_w2062_,
		_w2063_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h2)
	) name2000 (
		_w2061_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h4)
	) name2001 (
		_w2061_,
		_w2065_,
		_w2067_
	);
	LUT2 #(
		.INIT('h9)
	) name2002 (
		_w2061_,
		_w2065_,
		_w2068_
	);
	LUT3 #(
		.INIT('h71)
	) name2003 (
		_w1952_,
		_w1953_,
		_w1955_,
		_w2069_
	);
	LUT2 #(
		.INIT('h8)
	) name2004 (
		\a[12] ,
		\a[31] ,
		_w2070_
	);
	LUT4 #(
		.INIT('h153f)
	) name2005 (
		\a[6] ,
		\a[11] ,
		\a[32] ,
		\a[37] ,
		_w2071_
	);
	LUT4 #(
		.INIT('h8000)
	) name2006 (
		\a[6] ,
		\a[11] ,
		\a[32] ,
		\a[37] ,
		_w2072_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2007 (
		\a[6] ,
		\a[11] ,
		\a[32] ,
		\a[37] ,
		_w2073_
	);
	LUT2 #(
		.INIT('h6)
	) name2008 (
		_w2070_,
		_w2073_,
		_w2074_
	);
	LUT4 #(
		.INIT('h8e00)
	) name2009 (
		_w1947_,
		_w1948_,
		_w1949_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('h0071)
	) name2010 (
		_w1947_,
		_w1948_,
		_w1949_,
		_w2074_,
		_w2076_
	);
	LUT3 #(
		.INIT('ha9)
	) name2011 (
		_w2069_,
		_w2075_,
		_w2076_,
		_w2077_
	);
	LUT4 #(
		.INIT('h3701)
	) name2012 (
		_w1861_,
		_w1950_,
		_w1951_,
		_w1956_,
		_w2078_
	);
	LUT4 #(
		.INIT('h6996)
	) name2013 (
		_w2057_,
		_w2068_,
		_w2077_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h4)
	) name2014 (
		_w2056_,
		_w2079_,
		_w2080_
	);
	LUT2 #(
		.INIT('h8)
	) name2015 (
		_w2056_,
		_w2079_,
		_w2081_
	);
	LUT3 #(
		.INIT('h9f)
	) name2016 (
		_w2020_,
		_w2056_,
		_w2079_,
		_w2082_
	);
	LUT3 #(
		.INIT('h96)
	) name2017 (
		_w2020_,
		_w2056_,
		_w2079_,
		_w2083_
	);
	LUT4 #(
		.INIT('hd22d)
	) name2018 (
		_w1991_,
		_w2003_,
		_w2019_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		_w2002_,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h2)
	) name2020 (
		_w2002_,
		_w2084_,
		_w2086_
	);
	LUT2 #(
		.INIT('h9)
	) name2021 (
		_w2002_,
		_w2084_,
		_w2087_
	);
	LUT4 #(
		.INIT('hdc23)
	) name2022 (
		_w1917_,
		_w1998_,
		_w2001_,
		_w2087_,
		_w2088_
	);
	LUT3 #(
		.INIT('h01)
	) name2023 (
		_w1907_,
		_w1996_,
		_w2085_,
		_w2089_
	);
	LUT4 #(
		.INIT('h1011)
	) name2024 (
		_w1994_,
		_w1997_,
		_w2002_,
		_w2084_,
		_w2090_
	);
	LUT3 #(
		.INIT('h15)
	) name2025 (
		_w2004_,
		_w2008_,
		_w2018_,
		_w2091_
	);
	LUT3 #(
		.INIT('he8)
	) name2026 (
		_w2004_,
		_w2008_,
		_w2018_,
		_w2092_
	);
	LUT3 #(
		.INIT('h0e)
	) name2027 (
		_w2069_,
		_w2075_,
		_w2076_,
		_w2093_
	);
	LUT4 #(
		.INIT('h8000)
	) name2028 (
		\a[1] ,
		\a[21] ,
		\a[23] ,
		\a[43] ,
		_w2094_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2029 (
		\a[1] ,
		\a[21] ,
		\a[23] ,
		\a[43] ,
		_w2095_
	);
	LUT4 #(
		.INIT('h000d)
	) name2030 (
		_w1876_,
		_w2043_,
		_w2044_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('hf200)
	) name2031 (
		_w1876_,
		_w2043_,
		_w2044_,
		_w2095_,
		_w2097_
	);
	LUT4 #(
		.INIT('h0df2)
	) name2032 (
		_w1876_,
		_w2043_,
		_w2044_,
		_w2095_,
		_w2098_
	);
	LUT3 #(
		.INIT('h0d)
	) name2033 (
		_w2038_,
		_w2039_,
		_w2041_,
		_w2099_
	);
	LUT2 #(
		.INIT('h6)
	) name2034 (
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT3 #(
		.INIT('h32)
	) name2035 (
		_w2070_,
		_w2071_,
		_w2072_,
		_w2101_
	);
	LUT3 #(
		.INIT('h0d)
	) name2036 (
		_w2021_,
		_w2022_,
		_w2024_,
		_w2102_
	);
	LUT4 #(
		.INIT('h153f)
	) name2037 (
		\a[0] ,
		\a[2] ,
		\a[42] ,
		\a[44] ,
		_w2103_
	);
	LUT2 #(
		.INIT('h8)
	) name2038 (
		\a[2] ,
		\a[44] ,
		_w2104_
	);
	LUT4 #(
		.INIT('h8000)
	) name2039 (
		\a[0] ,
		\a[2] ,
		\a[42] ,
		\a[44] ,
		_w2105_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2040 (
		\a[0] ,
		\a[2] ,
		\a[42] ,
		\a[44] ,
		_w2106_
	);
	LUT2 #(
		.INIT('h6)
	) name2041 (
		_w2010_,
		_w2106_,
		_w2107_
	);
	LUT3 #(
		.INIT('h69)
	) name2042 (
		_w2101_,
		_w2102_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h4)
	) name2043 (
		_w2100_,
		_w2108_,
		_w2109_
	);
	LUT2 #(
		.INIT('h2)
	) name2044 (
		_w2100_,
		_w2108_,
		_w2110_
	);
	LUT2 #(
		.INIT('h9)
	) name2045 (
		_w2100_,
		_w2108_,
		_w2111_
	);
	LUT2 #(
		.INIT('h6)
	) name2046 (
		_w2093_,
		_w2111_,
		_w2112_
	);
	LUT3 #(
		.INIT('he8)
	) name2047 (
		_w2062_,
		_w2063_,
		_w2064_,
		_w2113_
	);
	LUT3 #(
		.INIT('h45)
	) name2048 (
		_w2012_,
		_w2013_,
		_w2015_,
		_w2114_
	);
	LUT3 #(
		.INIT('h2b)
	) name2049 (
		_w2058_,
		_w2059_,
		_w2060_,
		_w2115_
	);
	LUT3 #(
		.INIT('h96)
	) name2050 (
		_w2113_,
		_w2114_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('hb200)
	) name2051 (
		_w2057_,
		_w2061_,
		_w2065_,
		_w2116_,
		_w2117_
	);
	LUT4 #(
		.INIT('h004d)
	) name2052 (
		_w2057_,
		_w2061_,
		_w2065_,
		_w2116_,
		_w2118_
	);
	LUT4 #(
		.INIT('hcd32)
	) name2053 (
		_w2057_,
		_w2066_,
		_w2067_,
		_w2116_,
		_w2119_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w2112_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h6)
	) name2055 (
		_w2112_,
		_w2119_,
		_w2121_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		\a[3] ,
		\a[41] ,
		_w2122_
	);
	LUT4 #(
		.INIT('h153f)
	) name2057 (
		\a[15] ,
		\a[17] ,
		\a[27] ,
		\a[29] ,
		_w2123_
	);
	LUT4 #(
		.INIT('h8000)
	) name2058 (
		\a[15] ,
		\a[17] ,
		\a[27] ,
		\a[29] ,
		_w2124_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2059 (
		\a[15] ,
		\a[17] ,
		\a[27] ,
		\a[29] ,
		_w2125_
	);
	LUT2 #(
		.INIT('h8)
	) name2060 (
		\a[18] ,
		\a[26] ,
		_w2126_
	);
	LUT4 #(
		.INIT('h153f)
	) name2061 (
		\a[19] ,
		\a[20] ,
		\a[24] ,
		\a[25] ,
		_w2127_
	);
	LUT4 #(
		.INIT('h8000)
	) name2062 (
		\a[19] ,
		\a[20] ,
		\a[24] ,
		\a[25] ,
		_w2128_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2063 (
		\a[19] ,
		\a[20] ,
		\a[24] ,
		\a[25] ,
		_w2129_
	);
	LUT4 #(
		.INIT('h0660)
	) name2064 (
		_w2122_,
		_w2125_,
		_w2126_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('h9009)
	) name2065 (
		_w2122_,
		_w2125_,
		_w2126_,
		_w2129_,
		_w2131_
	);
	LUT4 #(
		.INIT('h6996)
	) name2066 (
		_w2122_,
		_w2125_,
		_w2126_,
		_w2129_,
		_w2132_
	);
	LUT2 #(
		.INIT('h8)
	) name2067 (
		\a[6] ,
		\a[38] ,
		_w2133_
	);
	LUT4 #(
		.INIT('h153f)
	) name2068 (
		\a[7] ,
		\a[11] ,
		\a[33] ,
		\a[37] ,
		_w2134_
	);
	LUT4 #(
		.INIT('h8000)
	) name2069 (
		\a[7] ,
		\a[11] ,
		\a[33] ,
		\a[37] ,
		_w2135_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2070 (
		\a[7] ,
		\a[11] ,
		\a[33] ,
		\a[37] ,
		_w2136_
	);
	LUT2 #(
		.INIT('h6)
	) name2071 (
		_w2133_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		\a[8] ,
		\a[36] ,
		_w2138_
	);
	LUT4 #(
		.INIT('h153f)
	) name2073 (
		\a[9] ,
		\a[10] ,
		\a[34] ,
		\a[35] ,
		_w2139_
	);
	LUT4 #(
		.INIT('h8000)
	) name2074 (
		\a[9] ,
		\a[10] ,
		\a[34] ,
		\a[35] ,
		_w2140_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2075 (
		\a[9] ,
		\a[10] ,
		\a[34] ,
		\a[35] ,
		_w2141_
	);
	LUT4 #(
		.INIT('h153f)
	) name2076 (
		\a[4] ,
		\a[14] ,
		\a[30] ,
		\a[40] ,
		_w2142_
	);
	LUT4 #(
		.INIT('h8000)
	) name2077 (
		\a[4] ,
		\a[14] ,
		\a[30] ,
		\a[40] ,
		_w2143_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2078 (
		\a[4] ,
		\a[14] ,
		\a[30] ,
		\a[40] ,
		_w2144_
	);
	LUT4 #(
		.INIT('h1428)
	) name2079 (
		_w2023_,
		_w2138_,
		_w2141_,
		_w2144_,
		_w2145_
	);
	LUT4 #(
		.INIT('h8241)
	) name2080 (
		_w2023_,
		_w2138_,
		_w2141_,
		_w2144_,
		_w2146_
	);
	LUT4 #(
		.INIT('h6996)
	) name2081 (
		_w2023_,
		_w2138_,
		_w2141_,
		_w2144_,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		\a[5] ,
		\a[39] ,
		_w2148_
	);
	LUT4 #(
		.INIT('h153f)
	) name2083 (
		\a[12] ,
		\a[13] ,
		\a[31] ,
		\a[32] ,
		_w2149_
	);
	LUT4 #(
		.INIT('h8000)
	) name2084 (
		\a[12] ,
		\a[13] ,
		\a[31] ,
		\a[32] ,
		_w2150_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2085 (
		\a[12] ,
		\a[13] ,
		\a[31] ,
		\a[32] ,
		_w2151_
	);
	LUT2 #(
		.INIT('h6)
	) name2086 (
		_w2148_,
		_w2151_,
		_w2152_
	);
	LUT4 #(
		.INIT('h0660)
	) name2087 (
		_w2132_,
		_w2137_,
		_w2147_,
		_w2152_,
		_w2153_
	);
	LUT4 #(
		.INIT('h6996)
	) name2088 (
		_w2132_,
		_w2137_,
		_w2147_,
		_w2152_,
		_w2154_
	);
	LUT4 #(
		.INIT('hb200)
	) name2089 (
		_w2009_,
		_w2016_,
		_w2017_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('h4db2)
	) name2090 (
		_w2009_,
		_w2016_,
		_w2017_,
		_w2154_,
		_w2156_
	);
	LUT3 #(
		.INIT('h09)
	) name2091 (
		_w2112_,
		_w2119_,
		_w2156_,
		_w2157_
	);
	LUT3 #(
		.INIT('h90)
	) name2092 (
		_w2112_,
		_w2119_,
		_w2156_,
		_w2158_
	);
	LUT3 #(
		.INIT('h27)
	) name2093 (
		_w2092_,
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT4 #(
		.INIT('h1700)
	) name2094 (
		_w2004_,
		_w2008_,
		_w2018_,
		_w2156_,
		_w2160_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2095 (
		_w2004_,
		_w2008_,
		_w2018_,
		_w2156_,
		_w2161_
	);
	LUT3 #(
		.INIT('h02)
	) name2096 (
		_w2121_,
		_w2160_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h2)
	) name2097 (
		_w2159_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('h8e00)
	) name2098 (
		_w1918_,
		_w1922_,
		_w1923_,
		_w2056_,
		_w2164_
	);
	LUT4 #(
		.INIT('h0027)
	) name2099 (
		_w2020_,
		_w2080_,
		_w2081_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('hf660)
	) name2100 (
		_w2057_,
		_w2068_,
		_w2077_,
		_w2078_,
		_w2166_
	);
	LUT3 #(
		.INIT('h32)
	) name2101 (
		_w2026_,
		_w2027_,
		_w2028_,
		_w2167_
	);
	LUT3 #(
		.INIT('h32)
	) name2102 (
		_w1887_,
		_w2049_,
		_w2050_,
		_w2168_
	);
	LUT3 #(
		.INIT('h0d)
	) name2103 (
		_w2033_,
		_w2034_,
		_w2035_,
		_w2169_
	);
	LUT3 #(
		.INIT('h96)
	) name2104 (
		_w2167_,
		_w2168_,
		_w2169_,
		_w2170_
	);
	LUT3 #(
		.INIT('h32)
	) name2105 (
		_w2030_,
		_w2031_,
		_w2037_,
		_w2171_
	);
	LUT3 #(
		.INIT('h32)
	) name2106 (
		_w2046_,
		_w2047_,
		_w2052_,
		_w2172_
	);
	LUT3 #(
		.INIT('h69)
	) name2107 (
		_w2170_,
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT3 #(
		.INIT('he0)
	) name2108 (
		_w2053_,
		_w2055_,
		_w2173_,
		_w2174_
	);
	LUT3 #(
		.INIT('h01)
	) name2109 (
		_w2053_,
		_w2055_,
		_w2173_,
		_w2175_
	);
	LUT3 #(
		.INIT('h1e)
	) name2110 (
		_w2053_,
		_w2055_,
		_w2173_,
		_w2176_
	);
	LUT2 #(
		.INIT('h6)
	) name2111 (
		_w2166_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h4)
	) name2112 (
		_w2165_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name2113 (
		_w2164_,
		_w2177_,
		_w2179_
	);
	LUT2 #(
		.INIT('h8)
	) name2114 (
		_w2082_,
		_w2179_,
		_w2180_
	);
	LUT4 #(
		.INIT('h022f)
	) name2115 (
		_w1991_,
		_w2003_,
		_w2019_,
		_w2083_,
		_w2181_
	);
	LUT4 #(
		.INIT('h51f3)
	) name2116 (
		_w2082_,
		_w2159_,
		_w2162_,
		_w2179_,
		_w2182_
	);
	LUT4 #(
		.INIT('h0056)
	) name2117 (
		_w2163_,
		_w2178_,
		_w2180_,
		_w2181_,
		_w2183_
	);
	LUT4 #(
		.INIT('ha900)
	) name2118 (
		_w2163_,
		_w2178_,
		_w2180_,
		_w2181_,
		_w2184_
	);
	LUT4 #(
		.INIT('h56a9)
	) name2119 (
		_w2163_,
		_w2178_,
		_w2180_,
		_w2181_,
		_w2185_
	);
	LUT3 #(
		.INIT('h10)
	) name2120 (
		_w2086_,
		_w2090_,
		_w2185_,
		_w2186_
	);
	LUT3 #(
		.INIT('hb0)
	) name2121 (
		_w1917_,
		_w2089_,
		_w2186_,
		_w2187_
	);
	LUT4 #(
		.INIT('hef0e)
	) name2122 (
		_w1994_,
		_w1997_,
		_w2002_,
		_w2084_,
		_w2188_
	);
	LUT4 #(
		.INIT('h040f)
	) name2123 (
		_w1917_,
		_w2089_,
		_w2185_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w2187_,
		_w2189_,
		_w2190_
	);
	LUT3 #(
		.INIT('h01)
	) name2125 (
		_w2086_,
		_w2090_,
		_w2184_,
		_w2191_
	);
	LUT4 #(
		.INIT('he800)
	) name2126 (
		_w2004_,
		_w2008_,
		_w2018_,
		_w2156_,
		_w2192_
	);
	LUT2 #(
		.INIT('h1)
	) name2127 (
		_w2120_,
		_w2192_,
		_w2193_
	);
	LUT3 #(
		.INIT('he0)
	) name2128 (
		_w2112_,
		_w2119_,
		_w2156_,
		_w2194_
	);
	LUT4 #(
		.INIT('heee0)
	) name2129 (
		_w2008_,
		_w2018_,
		_w2112_,
		_w2119_,
		_w2195_
	);
	LUT3 #(
		.INIT('h23)
	) name2130 (
		_w2091_,
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT3 #(
		.INIT('h0e)
	) name2131 (
		_w2112_,
		_w2117_,
		_w2118_,
		_w2197_
	);
	LUT2 #(
		.INIT('h1)
	) name2132 (
		_w2153_,
		_w2155_,
		_w2198_
	);
	LUT3 #(
		.INIT('he8)
	) name2133 (
		_w2113_,
		_w2114_,
		_w2115_,
		_w2199_
	);
	LUT3 #(
		.INIT('h32)
	) name2134 (
		_w2010_,
		_w2103_,
		_w2105_,
		_w2200_
	);
	LUT3 #(
		.INIT('h0d)
	) name2135 (
		_w2122_,
		_w2123_,
		_w2124_,
		_w2201_
	);
	LUT3 #(
		.INIT('h0d)
	) name2136 (
		_w2126_,
		_w2127_,
		_w2128_,
		_w2202_
	);
	LUT3 #(
		.INIT('h69)
	) name2137 (
		_w2200_,
		_w2201_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h8)
	) name2138 (
		\a[3] ,
		\a[42] ,
		_w2204_
	);
	LUT3 #(
		.INIT('h93)
	) name2139 (
		\a[1] ,
		\a[23] ,
		\a[44] ,
		_w2205_
	);
	LUT3 #(
		.INIT('h69)
	) name2140 (
		_w2094_,
		_w2204_,
		_w2205_,
		_w2206_
	);
	LUT4 #(
		.INIT('h153f)
	) name2141 (
		\a[6] ,
		\a[11] ,
		\a[34] ,
		\a[39] ,
		_w2207_
	);
	LUT4 #(
		.INIT('h8000)
	) name2142 (
		\a[6] ,
		\a[11] ,
		\a[34] ,
		\a[39] ,
		_w2208_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2143 (
		\a[6] ,
		\a[11] ,
		\a[34] ,
		\a[39] ,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name2144 (
		\a[15] ,
		\a[30] ,
		_w2210_
	);
	LUT4 #(
		.INIT('h153f)
	) name2145 (
		\a[16] ,
		\a[17] ,
		\a[28] ,
		\a[29] ,
		_w2211_
	);
	LUT4 #(
		.INIT('h8000)
	) name2146 (
		\a[16] ,
		\a[17] ,
		\a[28] ,
		\a[29] ,
		_w2212_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2147 (
		\a[16] ,
		\a[17] ,
		\a[28] ,
		\a[29] ,
		_w2213_
	);
	LUT4 #(
		.INIT('h0660)
	) name2148 (
		_w1530_,
		_w2209_,
		_w2210_,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('h9009)
	) name2149 (
		_w1530_,
		_w2209_,
		_w2210_,
		_w2213_,
		_w2215_
	);
	LUT4 #(
		.INIT('h6996)
	) name2150 (
		_w1530_,
		_w2209_,
		_w2210_,
		_w2213_,
		_w2216_
	);
	LUT2 #(
		.INIT('h6)
	) name2151 (
		_w2206_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name2152 (
		_w2203_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h4)
	) name2153 (
		_w2203_,
		_w2217_,
		_w2219_
	);
	LUT3 #(
		.INIT('h6f)
	) name2154 (
		_w2199_,
		_w2203_,
		_w2217_,
		_w2220_
	);
	LUT3 #(
		.INIT('h69)
	) name2155 (
		_w2199_,
		_w2203_,
		_w2217_,
		_w2221_
	);
	LUT3 #(
		.INIT('h69)
	) name2156 (
		_w2197_,
		_w2198_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('h4114)
	) name2157 (
		_w2192_,
		_w2197_,
		_w2198_,
		_w2221_,
		_w2223_
	);
	LUT3 #(
		.INIT('hd0)
	) name2158 (
		_w2193_,
		_w2196_,
		_w2223_,
		_w2224_
	);
	LUT4 #(
		.INIT('hae00)
	) name2159 (
		_w2192_,
		_w2193_,
		_w2196_,
		_w2222_,
		_w2225_
	);
	LUT4 #(
		.INIT('h51ae)
	) name2160 (
		_w2192_,
		_w2193_,
		_w2196_,
		_w2222_,
		_w2226_
	);
	LUT3 #(
		.INIT('h0e)
	) name2161 (
		_w2166_,
		_w2174_,
		_w2175_,
		_w2227_
	);
	LUT3 #(
		.INIT('hd4)
	) name2162 (
		_w2170_,
		_w2171_,
		_w2172_,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		\a[0] ,
		\a[45] ,
		_w2229_
	);
	LUT4 #(
		.INIT('h153f)
	) name2164 (
		\a[2] ,
		\a[4] ,
		\a[41] ,
		\a[43] ,
		_w2230_
	);
	LUT4 #(
		.INIT('h8000)
	) name2165 (
		\a[2] ,
		\a[4] ,
		\a[41] ,
		\a[43] ,
		_w2231_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2166 (
		\a[2] ,
		\a[4] ,
		\a[41] ,
		\a[43] ,
		_w2232_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		\a[7] ,
		\a[38] ,
		_w2233_
	);
	LUT4 #(
		.INIT('h153f)
	) name2168 (
		\a[8] ,
		\a[9] ,
		\a[36] ,
		\a[37] ,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		\a[9] ,
		\a[37] ,
		_w2235_
	);
	LUT4 #(
		.INIT('h8000)
	) name2170 (
		\a[8] ,
		\a[9] ,
		\a[36] ,
		\a[37] ,
		_w2236_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2171 (
		\a[8] ,
		\a[9] ,
		\a[36] ,
		\a[37] ,
		_w2237_
	);
	LUT4 #(
		.INIT('h0660)
	) name2172 (
		_w2229_,
		_w2232_,
		_w2233_,
		_w2237_,
		_w2238_
	);
	LUT4 #(
		.INIT('h9009)
	) name2173 (
		_w2229_,
		_w2232_,
		_w2233_,
		_w2237_,
		_w2239_
	);
	LUT4 #(
		.INIT('h6996)
	) name2174 (
		_w2229_,
		_w2232_,
		_w2233_,
		_w2237_,
		_w2240_
	);
	LUT4 #(
		.INIT('h153f)
	) name2175 (
		\a[21] ,
		\a[22] ,
		\a[23] ,
		\a[24] ,
		_w2241_
	);
	LUT4 #(
		.INIT('h8000)
	) name2176 (
		\a[21] ,
		\a[22] ,
		\a[23] ,
		\a[24] ,
		_w2242_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2177 (
		\a[21] ,
		\a[22] ,
		\a[23] ,
		\a[24] ,
		_w2243_
	);
	LUT2 #(
		.INIT('h6)
	) name2178 (
		_w2040_,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h6)
	) name2179 (
		_w2240_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		\a[18] ,
		\a[27] ,
		_w2246_
	);
	LUT4 #(
		.INIT('h153f)
	) name2181 (
		\a[19] ,
		\a[20] ,
		\a[25] ,
		\a[26] ,
		_w2247_
	);
	LUT4 #(
		.INIT('h8000)
	) name2182 (
		\a[19] ,
		\a[20] ,
		\a[25] ,
		\a[26] ,
		_w2248_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2183 (
		\a[19] ,
		\a[20] ,
		\a[25] ,
		\a[26] ,
		_w2249_
	);
	LUT2 #(
		.INIT('h6)
	) name2184 (
		_w2246_,
		_w2249_,
		_w2250_
	);
	LUT3 #(
		.INIT('h0d)
	) name2185 (
		_w2138_,
		_w2139_,
		_w2140_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name2186 (
		\a[14] ,
		\a[31] ,
		_w2252_
	);
	LUT4 #(
		.INIT('h153f)
	) name2187 (
		\a[5] ,
		\a[13] ,
		\a[32] ,
		\a[40] ,
		_w2253_
	);
	LUT4 #(
		.INIT('h8000)
	) name2188 (
		\a[5] ,
		\a[13] ,
		\a[32] ,
		\a[40] ,
		_w2254_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2189 (
		\a[5] ,
		\a[13] ,
		\a[32] ,
		\a[40] ,
		_w2255_
	);
	LUT2 #(
		.INIT('h6)
	) name2190 (
		_w2252_,
		_w2255_,
		_w2256_
	);
	LUT3 #(
		.INIT('h96)
	) name2191 (
		_w2250_,
		_w2251_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h2)
	) name2192 (
		_w2245_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h4)
	) name2193 (
		_w2245_,
		_w2257_,
		_w2259_
	);
	LUT2 #(
		.INIT('h9)
	) name2194 (
		_w2245_,
		_w2257_,
		_w2260_
	);
	LUT2 #(
		.INIT('h6)
	) name2195 (
		_w2228_,
		_w2260_,
		_w2261_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2196 (
		_w2166_,
		_w2174_,
		_w2175_,
		_w2261_,
		_w2262_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2197 (
		_w2166_,
		_w2174_,
		_w2175_,
		_w2261_,
		_w2263_
	);
	LUT3 #(
		.INIT('h8e)
	) name2198 (
		_w2167_,
		_w2168_,
		_w2169_,
		_w2264_
	);
	LUT3 #(
		.INIT('hb2)
	) name2199 (
		_w2101_,
		_w2102_,
		_w2107_,
		_w2265_
	);
	LUT3 #(
		.INIT('h45)
	) name2200 (
		_w2096_,
		_w2097_,
		_w2099_,
		_w2266_
	);
	LUT3 #(
		.INIT('h96)
	) name2201 (
		_w2264_,
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('h0031)
	) name2202 (
		_w2093_,
		_w2109_,
		_w2110_,
		_w2267_,
		_w2268_
	);
	LUT4 #(
		.INIT('hce00)
	) name2203 (
		_w2093_,
		_w2109_,
		_w2110_,
		_w2267_,
		_w2269_
	);
	LUT4 #(
		.INIT('h4db2)
	) name2204 (
		_w2093_,
		_w2100_,
		_w2108_,
		_w2267_,
		_w2270_
	);
	LUT3 #(
		.INIT('h32)
	) name2205 (
		_w2023_,
		_w2142_,
		_w2143_,
		_w2271_
	);
	LUT3 #(
		.INIT('h0d)
	) name2206 (
		_w2133_,
		_w2134_,
		_w2135_,
		_w2272_
	);
	LUT3 #(
		.INIT('h0d)
	) name2207 (
		_w2148_,
		_w2149_,
		_w2150_,
		_w2273_
	);
	LUT3 #(
		.INIT('h69)
	) name2208 (
		_w2271_,
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT3 #(
		.INIT('h32)
	) name2209 (
		_w2145_,
		_w2146_,
		_w2152_,
		_w2275_
	);
	LUT3 #(
		.INIT('h32)
	) name2210 (
		_w2130_,
		_w2131_,
		_w2137_,
		_w2276_
	);
	LUT3 #(
		.INIT('h69)
	) name2211 (
		_w2274_,
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('h6)
	) name2212 (
		_w2270_,
		_w2277_,
		_w2278_
	);
	LUT3 #(
		.INIT('h10)
	) name2213 (
		_w2262_,
		_w2263_,
		_w2278_,
		_w2279_
	);
	LUT3 #(
		.INIT('h41)
	) name2214 (
		_w2261_,
		_w2270_,
		_w2277_,
		_w2280_
	);
	LUT3 #(
		.INIT('h82)
	) name2215 (
		_w2261_,
		_w2270_,
		_w2277_,
		_w2281_
	);
	LUT3 #(
		.INIT('h1b)
	) name2216 (
		_w2227_,
		_w2280_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h4)
	) name2217 (
		_w2279_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w2226_,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h1)
	) name2219 (
		_w2178_,
		_w2182_,
		_w2285_
	);
	LUT3 #(
		.INIT('h10)
	) name2220 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2286_
	);
	LUT3 #(
		.INIT('he1)
	) name2221 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name2222 (
		_w2285_,
		_w2287_,
		_w2288_
	);
	LUT3 #(
		.INIT('h36)
	) name2223 (
		_w2284_,
		_w2285_,
		_w2286_,
		_w2289_
	);
	LUT4 #(
		.INIT('h0514)
	) name2224 (
		_w2183_,
		_w2284_,
		_w2285_,
		_w2286_,
		_w2290_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2225 (
		_w1917_,
		_w2089_,
		_w2191_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('h040f)
	) name2226 (
		_w1917_,
		_w2089_,
		_w2183_,
		_w2191_,
		_w2292_
	);
	LUT3 #(
		.INIT('hcd)
	) name2227 (
		_w2289_,
		_w2291_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('h5554)
	) name2228 (
		_w2183_,
		_w2284_,
		_w2285_,
		_w2286_,
		_w2294_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2229 (
		_w1917_,
		_w2089_,
		_w2191_,
		_w2294_,
		_w2295_
	);
	LUT3 #(
		.INIT('h23)
	) name2230 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2296_
	);
	LUT3 #(
		.INIT('hd4)
	) name2231 (
		_w2274_,
		_w2275_,
		_w2276_,
		_w2297_
	);
	LUT3 #(
		.INIT('h8e)
	) name2232 (
		_w2094_,
		_w2204_,
		_w2205_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name2233 (
		\a[16] ,
		\a[30] ,
		_w2299_
	);
	LUT4 #(
		.INIT('h153f)
	) name2234 (
		\a[17] ,
		\a[18] ,
		\a[28] ,
		\a[29] ,
		_w2300_
	);
	LUT4 #(
		.INIT('h8000)
	) name2235 (
		\a[17] ,
		\a[18] ,
		\a[28] ,
		\a[29] ,
		_w2301_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2236 (
		\a[17] ,
		\a[18] ,
		\a[28] ,
		\a[29] ,
		_w2302_
	);
	LUT2 #(
		.INIT('h6)
	) name2237 (
		_w2299_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h8)
	) name2238 (
		\a[12] ,
		\a[34] ,
		_w2304_
	);
	LUT4 #(
		.INIT('h153f)
	) name2239 (
		\a[7] ,
		\a[8] ,
		\a[38] ,
		\a[39] ,
		_w2305_
	);
	LUT2 #(
		.INIT('h8)
	) name2240 (
		\a[8] ,
		\a[39] ,
		_w2306_
	);
	LUT4 #(
		.INIT('h8000)
	) name2241 (
		\a[7] ,
		\a[8] ,
		\a[38] ,
		\a[39] ,
		_w2307_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2242 (
		\a[7] ,
		\a[8] ,
		\a[38] ,
		\a[39] ,
		_w2308_
	);
	LUT2 #(
		.INIT('h6)
	) name2243 (
		_w2304_,
		_w2308_,
		_w2309_
	);
	LUT3 #(
		.INIT('h96)
	) name2244 (
		_w2298_,
		_w2303_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('h153f)
	) name2245 (
		\a[10] ,
		\a[11] ,
		\a[35] ,
		\a[36] ,
		_w2311_
	);
	LUT4 #(
		.INIT('h8000)
	) name2246 (
		\a[10] ,
		\a[11] ,
		\a[35] ,
		\a[36] ,
		_w2312_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2247 (
		\a[10] ,
		\a[11] ,
		\a[35] ,
		\a[36] ,
		_w2313_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		\a[3] ,
		\a[43] ,
		_w2314_
	);
	LUT4 #(
		.INIT('h153f)
	) name2249 (
		\a[0] ,
		\a[4] ,
		\a[42] ,
		\a[46] ,
		_w2315_
	);
	LUT4 #(
		.INIT('h8000)
	) name2250 (
		\a[0] ,
		\a[4] ,
		\a[42] ,
		\a[46] ,
		_w2316_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2251 (
		\a[0] ,
		\a[4] ,
		\a[42] ,
		\a[46] ,
		_w2317_
	);
	LUT4 #(
		.INIT('h0660)
	) name2252 (
		_w2235_,
		_w2313_,
		_w2314_,
		_w2317_,
		_w2318_
	);
	LUT4 #(
		.INIT('h9009)
	) name2253 (
		_w2235_,
		_w2313_,
		_w2314_,
		_w2317_,
		_w2319_
	);
	LUT4 #(
		.INIT('h6996)
	) name2254 (
		_w2235_,
		_w2313_,
		_w2314_,
		_w2317_,
		_w2320_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		\a[19] ,
		\a[27] ,
		_w2321_
	);
	LUT4 #(
		.INIT('h153f)
	) name2256 (
		\a[20] ,
		\a[21] ,
		\a[25] ,
		\a[26] ,
		_w2322_
	);
	LUT4 #(
		.INIT('h8000)
	) name2257 (
		\a[20] ,
		\a[21] ,
		\a[25] ,
		\a[26] ,
		_w2323_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2258 (
		\a[20] ,
		\a[21] ,
		\a[25] ,
		\a[26] ,
		_w2324_
	);
	LUT2 #(
		.INIT('h6)
	) name2259 (
		_w2321_,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h6)
	) name2260 (
		_w2320_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name2261 (
		_w2310_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h1)
	) name2262 (
		_w2310_,
		_w2326_,
		_w2328_
	);
	LUT2 #(
		.INIT('h6)
	) name2263 (
		_w2310_,
		_w2326_,
		_w2329_
	);
	LUT2 #(
		.INIT('h6)
	) name2264 (
		_w2297_,
		_w2329_,
		_w2330_
	);
	LUT3 #(
		.INIT('h40)
	) name2265 (
		_w2198_,
		_w2221_,
		_w2330_,
		_w2331_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name2266 (
		_w2153_,
		_w2155_,
		_w2297_,
		_w2329_,
		_w2332_
	);
	LUT2 #(
		.INIT('h8)
	) name2267 (
		_w2221_,
		_w2330_,
		_w2333_
	);
	LUT4 #(
		.INIT('h1113)
	) name2268 (
		_w2197_,
		_w2331_,
		_w2332_,
		_w2333_,
		_w2334_
	);
	LUT4 #(
		.INIT('h004d)
	) name2269 (
		_w2197_,
		_w2198_,
		_w2221_,
		_w2330_,
		_w2335_
	);
	LUT4 #(
		.INIT('h4db2)
	) name2270 (
		_w2197_,
		_w2198_,
		_w2221_,
		_w2330_,
		_w2336_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2271 (
		_w2113_,
		_w2114_,
		_w2115_,
		_w2203_,
		_w2337_
	);
	LUT4 #(
		.INIT('h0027)
	) name2272 (
		_w2199_,
		_w2218_,
		_w2219_,
		_w2337_,
		_w2338_
	);
	LUT3 #(
		.INIT('h32)
	) name2273 (
		_w2252_,
		_w2253_,
		_w2254_,
		_w2339_
	);
	LUT3 #(
		.INIT('h0d)
	) name2274 (
		_w2229_,
		_w2230_,
		_w2231_,
		_w2340_
	);
	LUT3 #(
		.INIT('h0d)
	) name2275 (
		_w2233_,
		_w2234_,
		_w2236_,
		_w2341_
	);
	LUT3 #(
		.INIT('h69)
	) name2276 (
		_w2339_,
		_w2340_,
		_w2341_,
		_w2342_
	);
	LUT3 #(
		.INIT('h2b)
	) name2277 (
		_w2200_,
		_w2201_,
		_w2202_,
		_w2343_
	);
	LUT3 #(
		.INIT('h80)
	) name2278 (
		\a[1] ,
		\a[23] ,
		\a[44] ,
		_w2344_
	);
	LUT4 #(
		.INIT('h8000)
	) name2279 (
		\a[1] ,
		\a[22] ,
		\a[24] ,
		\a[45] ,
		_w2345_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2280 (
		\a[1] ,
		\a[22] ,
		\a[24] ,
		\a[45] ,
		_w2346_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		_w2344_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w2344_,
		_w2346_,
		_w2348_
	);
	LUT2 #(
		.INIT('h6)
	) name2283 (
		_w2344_,
		_w2346_,
		_w2349_
	);
	LUT3 #(
		.INIT('h0d)
	) name2284 (
		_w2040_,
		_w2241_,
		_w2242_,
		_w2350_
	);
	LUT2 #(
		.INIT('h6)
	) name2285 (
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT3 #(
		.INIT('h96)
	) name2286 (
		_w2342_,
		_w2343_,
		_w2351_,
		_w2352_
	);
	LUT3 #(
		.INIT('h32)
	) name2287 (
		_w2238_,
		_w2239_,
		_w2244_,
		_w2353_
	);
	LUT3 #(
		.INIT('h4d)
	) name2288 (
		_w2250_,
		_w2251_,
		_w2256_,
		_w2354_
	);
	LUT3 #(
		.INIT('h0e)
	) name2289 (
		_w2206_,
		_w2214_,
		_w2215_,
		_w2355_
	);
	LUT3 #(
		.INIT('h69)
	) name2290 (
		_w2353_,
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w2337_,
		_w2352_,
		_w2357_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2292 (
		_w2220_,
		_w2337_,
		_w2352_,
		_w2356_,
		_w2358_
	);
	LUT3 #(
		.INIT('h20)
	) name2293 (
		_w2220_,
		_w2356_,
		_w2357_,
		_w2359_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w2352_,
		_w2356_,
		_w2360_
	);
	LUT2 #(
		.INIT('h4)
	) name2295 (
		_w2338_,
		_w2360_,
		_w2361_
	);
	LUT3 #(
		.INIT('h01)
	) name2296 (
		_w2358_,
		_w2359_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h6)
	) name2297 (
		_w2336_,
		_w2362_,
		_w2363_
	);
	LUT3 #(
		.INIT('h54)
	) name2298 (
		_w2262_,
		_w2263_,
		_w2278_,
		_w2364_
	);
	LUT3 #(
		.INIT('h54)
	) name2299 (
		_w2268_,
		_w2269_,
		_w2277_,
		_w2365_
	);
	LUT3 #(
		.INIT('h31)
	) name2300 (
		_w2228_,
		_w2258_,
		_w2259_,
		_w2366_
	);
	LUT3 #(
		.INIT('he8)
	) name2301 (
		_w2264_,
		_w2265_,
		_w2266_,
		_w2367_
	);
	LUT3 #(
		.INIT('h0d)
	) name2302 (
		_w2210_,
		_w2211_,
		_w2212_,
		_w2368_
	);
	LUT3 #(
		.INIT('h0d)
	) name2303 (
		_w2246_,
		_w2247_,
		_w2248_,
		_w2369_
	);
	LUT3 #(
		.INIT('h0d)
	) name2304 (
		_w1530_,
		_w2207_,
		_w2208_,
		_w2370_
	);
	LUT3 #(
		.INIT('h96)
	) name2305 (
		_w2368_,
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('h153f)
	) name2306 (
		\a[5] ,
		\a[15] ,
		\a[31] ,
		\a[41] ,
		_w2372_
	);
	LUT4 #(
		.INIT('h8000)
	) name2307 (
		\a[5] ,
		\a[15] ,
		\a[31] ,
		\a[41] ,
		_w2373_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2308 (
		\a[5] ,
		\a[15] ,
		\a[31] ,
		\a[41] ,
		_w2374_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		\a[14] ,
		\a[32] ,
		_w2375_
	);
	LUT4 #(
		.INIT('h153f)
	) name2310 (
		\a[6] ,
		\a[13] ,
		\a[33] ,
		\a[40] ,
		_w2376_
	);
	LUT4 #(
		.INIT('h8000)
	) name2311 (
		\a[6] ,
		\a[13] ,
		\a[33] ,
		\a[40] ,
		_w2377_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2312 (
		\a[6] ,
		\a[13] ,
		\a[33] ,
		\a[40] ,
		_w2378_
	);
	LUT4 #(
		.INIT('h0660)
	) name2313 (
		_w2104_,
		_w2374_,
		_w2375_,
		_w2378_,
		_w2379_
	);
	LUT4 #(
		.INIT('h6996)
	) name2314 (
		_w2104_,
		_w2374_,
		_w2375_,
		_w2378_,
		_w2380_
	);
	LUT4 #(
		.INIT('h2b00)
	) name2315 (
		_w2271_,
		_w2272_,
		_w2273_,
		_w2380_,
		_w2381_
	);
	LUT4 #(
		.INIT('hd42b)
	) name2316 (
		_w2271_,
		_w2272_,
		_w2273_,
		_w2380_,
		_w2382_
	);
	LUT2 #(
		.INIT('h8)
	) name2317 (
		_w2371_,
		_w2382_,
		_w2383_
	);
	LUT2 #(
		.INIT('h4)
	) name2318 (
		_w2371_,
		_w2382_,
		_w2384_
	);
	LUT3 #(
		.INIT('h69)
	) name2319 (
		_w2367_,
		_w2371_,
		_w2382_,
		_w2385_
	);
	LUT3 #(
		.INIT('h69)
	) name2320 (
		_w2365_,
		_w2366_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w2364_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h6)
	) name2322 (
		_w2364_,
		_w2386_,
		_w2388_
	);
	LUT4 #(
		.INIT('h9009)
	) name2323 (
		_w2336_,
		_w2362_,
		_w2364_,
		_w2386_,
		_w2389_
	);
	LUT4 #(
		.INIT('h2300)
	) name2324 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2389_,
		_w2390_
	);
	LUT4 #(
		.INIT('h0990)
	) name2325 (
		_w2336_,
		_w2362_,
		_w2364_,
		_w2386_,
		_w2391_
	);
	LUT4 #(
		.INIT('hdc00)
	) name2326 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w2390_,
		_w2392_,
		_w2393_
	);
	LUT4 #(
		.INIT('h6006)
	) name2328 (
		_w2336_,
		_w2362_,
		_w2364_,
		_w2386_,
		_w2394_
	);
	LUT4 #(
		.INIT('hdc00)
	) name2329 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2394_,
		_w2395_
	);
	LUT4 #(
		.INIT('h0660)
	) name2330 (
		_w2336_,
		_w2362_,
		_w2364_,
		_w2386_,
		_w2396_
	);
	LUT4 #(
		.INIT('h2300)
	) name2331 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2396_,
		_w2397_
	);
	LUT2 #(
		.INIT('h1)
	) name2332 (
		_w2395_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('h69)
	) name2333 (
		_w2296_,
		_w2363_,
		_w2388_,
		_w2399_
	);
	LUT3 #(
		.INIT('he1)
	) name2334 (
		_w2288_,
		_w2295_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h8)
	) name2335 (
		_w2294_,
		_w2398_,
		_w2401_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2336 (
		_w1917_,
		_w2089_,
		_w2191_,
		_w2401_,
		_w2402_
	);
	LUT4 #(
		.INIT('h0002)
	) name2337 (
		_w2285_,
		_w2287_,
		_w2395_,
		_w2397_,
		_w2403_
	);
	LUT4 #(
		.INIT('hdc00)
	) name2338 (
		_w2224_,
		_w2225_,
		_w2283_,
		_w2388_,
		_w2404_
	);
	LUT3 #(
		.INIT('h4d)
	) name2339 (
		_w2365_,
		_w2366_,
		_w2385_,
		_w2405_
	);
	LUT4 #(
		.INIT('h022f)
	) name2340 (
		_w2220_,
		_w2337_,
		_w2352_,
		_w2356_,
		_w2406_
	);
	LUT3 #(
		.INIT('h0d)
	) name2341 (
		_w2321_,
		_w2322_,
		_w2323_,
		_w2407_
	);
	LUT3 #(
		.INIT('h0d)
	) name2342 (
		_w2104_,
		_w2372_,
		_w2373_,
		_w2408_
	);
	LUT3 #(
		.INIT('h32)
	) name2343 (
		_w2314_,
		_w2315_,
		_w2316_,
		_w2409_
	);
	LUT3 #(
		.INIT('h96)
	) name2344 (
		_w2407_,
		_w2408_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('h32)
	) name2345 (
		_w2318_,
		_w2319_,
		_w2325_,
		_w2411_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2346 (
		_w2379_,
		_w2381_,
		_w2410_,
		_w2411_,
		_w2412_
	);
	LUT3 #(
		.INIT('h31)
	) name2347 (
		_w2297_,
		_w2327_,
		_w2328_,
		_w2413_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2348 (
		_w2264_,
		_w2265_,
		_w2266_,
		_w2371_,
		_w2414_
	);
	LUT4 #(
		.INIT('h0027)
	) name2349 (
		_w2367_,
		_w2383_,
		_w2384_,
		_w2414_,
		_w2415_
	);
	LUT3 #(
		.INIT('h69)
	) name2350 (
		_w2412_,
		_w2413_,
		_w2415_,
		_w2416_
	);
	LUT3 #(
		.INIT('h96)
	) name2351 (
		_w2405_,
		_w2406_,
		_w2416_,
		_w2417_
	);
	LUT3 #(
		.INIT('h17)
	) name2352 (
		_w2368_,
		_w2369_,
		_w2370_,
		_w2418_
	);
	LUT3 #(
		.INIT('h23)
	) name2353 (
		_w2347_,
		_w2348_,
		_w2350_,
		_w2419_
	);
	LUT2 #(
		.INIT('h8)
	) name2354 (
		\a[13] ,
		\a[34] ,
		_w2420_
	);
	LUT4 #(
		.INIT('h153f)
	) name2355 (
		\a[7] ,
		\a[12] ,
		\a[35] ,
		\a[40] ,
		_w2421_
	);
	LUT4 #(
		.INIT('h8000)
	) name2356 (
		\a[7] ,
		\a[12] ,
		\a[35] ,
		\a[40] ,
		_w2422_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2357 (
		\a[7] ,
		\a[12] ,
		\a[35] ,
		\a[40] ,
		_w2423_
	);
	LUT2 #(
		.INIT('h6)
	) name2358 (
		_w2420_,
		_w2423_,
		_w2424_
	);
	LUT4 #(
		.INIT('h8e00)
	) name2359 (
		_w2344_,
		_w2346_,
		_w2350_,
		_w2424_,
		_w2425_
	);
	LUT4 #(
		.INIT('h0071)
	) name2360 (
		_w2344_,
		_w2346_,
		_w2350_,
		_w2424_,
		_w2426_
	);
	LUT4 #(
		.INIT('hdc23)
	) name2361 (
		_w2347_,
		_w2348_,
		_w2350_,
		_w2424_,
		_w2427_
	);
	LUT2 #(
		.INIT('h6)
	) name2362 (
		_w2418_,
		_w2427_,
		_w2428_
	);
	LUT3 #(
		.INIT('h4d)
	) name2363 (
		_w2342_,
		_w2343_,
		_w2351_,
		_w2429_
	);
	LUT3 #(
		.INIT('hb2)
	) name2364 (
		_w2353_,
		_w2354_,
		_w2355_,
		_w2430_
	);
	LUT3 #(
		.INIT('h96)
	) name2365 (
		_w2428_,
		_w2429_,
		_w2430_,
		_w2431_
	);
	LUT3 #(
		.INIT('h32)
	) name2366 (
		_w2375_,
		_w2376_,
		_w2377_,
		_w2432_
	);
	LUT3 #(
		.INIT('h0d)
	) name2367 (
		_w2299_,
		_w2300_,
		_w2301_,
		_w2433_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		\a[3] ,
		\a[44] ,
		_w2434_
	);
	LUT4 #(
		.INIT('h153f)
	) name2369 (
		\a[4] ,
		\a[15] ,
		\a[32] ,
		\a[43] ,
		_w2435_
	);
	LUT4 #(
		.INIT('h8000)
	) name2370 (
		\a[4] ,
		\a[15] ,
		\a[32] ,
		\a[43] ,
		_w2436_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2371 (
		\a[4] ,
		\a[15] ,
		\a[32] ,
		\a[43] ,
		_w2437_
	);
	LUT2 #(
		.INIT('h6)
	) name2372 (
		_w2434_,
		_w2437_,
		_w2438_
	);
	LUT3 #(
		.INIT('h69)
	) name2373 (
		_w2432_,
		_w2433_,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('h153f)
	) name2374 (
		\a[9] ,
		\a[11] ,
		\a[36] ,
		\a[38] ,
		_w2440_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		\a[11] ,
		\a[38] ,
		_w2441_
	);
	LUT4 #(
		.INIT('h8000)
	) name2376 (
		\a[9] ,
		\a[11] ,
		\a[36] ,
		\a[38] ,
		_w2442_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2377 (
		\a[9] ,
		\a[11] ,
		\a[36] ,
		\a[38] ,
		_w2443_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		\a[10] ,
		\a[37] ,
		_w2444_
	);
	LUT4 #(
		.INIT('h153f)
	) name2379 (
		\a[22] ,
		\a[23] ,
		\a[24] ,
		\a[25] ,
		_w2445_
	);
	LUT4 #(
		.INIT('h8000)
	) name2380 (
		\a[22] ,
		\a[23] ,
		\a[24] ,
		\a[25] ,
		_w2446_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2381 (
		\a[22] ,
		\a[23] ,
		\a[24] ,
		\a[25] ,
		_w2447_
	);
	LUT4 #(
		.INIT('h0660)
	) name2382 (
		_w2306_,
		_w2443_,
		_w2444_,
		_w2447_,
		_w2448_
	);
	LUT4 #(
		.INIT('h9009)
	) name2383 (
		_w2306_,
		_w2443_,
		_w2444_,
		_w2447_,
		_w2449_
	);
	LUT4 #(
		.INIT('h6996)
	) name2384 (
		_w2306_,
		_w2443_,
		_w2444_,
		_w2447_,
		_w2450_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		\a[5] ,
		\a[42] ,
		_w2451_
	);
	LUT4 #(
		.INIT('h153f)
	) name2386 (
		\a[6] ,
		\a[14] ,
		\a[33] ,
		\a[41] ,
		_w2452_
	);
	LUT4 #(
		.INIT('h8000)
	) name2387 (
		\a[6] ,
		\a[14] ,
		\a[33] ,
		\a[41] ,
		_w2453_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2388 (
		\a[6] ,
		\a[14] ,
		\a[33] ,
		\a[41] ,
		_w2454_
	);
	LUT2 #(
		.INIT('h6)
	) name2389 (
		_w2451_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h6)
	) name2390 (
		_w2450_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h153f)
	) name2391 (
		\a[0] ,
		\a[2] ,
		\a[45] ,
		\a[47] ,
		_w2457_
	);
	LUT4 #(
		.INIT('h8000)
	) name2392 (
		\a[0] ,
		\a[2] ,
		\a[45] ,
		\a[47] ,
		_w2458_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2393 (
		\a[0] ,
		\a[2] ,
		\a[45] ,
		\a[47] ,
		_w2459_
	);
	LUT2 #(
		.INIT('h8)
	) name2394 (
		\a[16] ,
		\a[31] ,
		_w2460_
	);
	LUT4 #(
		.INIT('h153f)
	) name2395 (
		\a[17] ,
		\a[18] ,
		\a[29] ,
		\a[30] ,
		_w2461_
	);
	LUT4 #(
		.INIT('h8000)
	) name2396 (
		\a[17] ,
		\a[18] ,
		\a[29] ,
		\a[30] ,
		_w2462_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2397 (
		\a[17] ,
		\a[18] ,
		\a[29] ,
		\a[30] ,
		_w2463_
	);
	LUT4 #(
		.INIT('h0660)
	) name2398 (
		_w2345_,
		_w2459_,
		_w2460_,
		_w2463_,
		_w2464_
	);
	LUT4 #(
		.INIT('h9009)
	) name2399 (
		_w2345_,
		_w2459_,
		_w2460_,
		_w2463_,
		_w2465_
	);
	LUT4 #(
		.INIT('h6996)
	) name2400 (
		_w2345_,
		_w2459_,
		_w2460_,
		_w2463_,
		_w2466_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		\a[19] ,
		\a[28] ,
		_w2467_
	);
	LUT4 #(
		.INIT('h153f)
	) name2402 (
		\a[20] ,
		\a[21] ,
		\a[26] ,
		\a[27] ,
		_w2468_
	);
	LUT4 #(
		.INIT('h8000)
	) name2403 (
		\a[20] ,
		\a[21] ,
		\a[26] ,
		\a[27] ,
		_w2469_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2404 (
		\a[20] ,
		\a[21] ,
		\a[26] ,
		\a[27] ,
		_w2470_
	);
	LUT2 #(
		.INIT('h6)
	) name2405 (
		_w2467_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h6)
	) name2406 (
		_w2466_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('h96)
	) name2407 (
		_w2439_,
		_w2456_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('he8)
	) name2408 (
		_w2298_,
		_w2303_,
		_w2309_,
		_w2474_
	);
	LUT3 #(
		.INIT('h2b)
	) name2409 (
		_w2339_,
		_w2340_,
		_w2341_,
		_w2475_
	);
	LUT3 #(
		.INIT('h80)
	) name2410 (
		\a[1] ,
		\a[24] ,
		\a[46] ,
		_w2476_
	);
	LUT3 #(
		.INIT('h6c)
	) name2411 (
		\a[1] ,
		\a[24] ,
		\a[46] ,
		_w2477_
	);
	LUT4 #(
		.INIT('hf200)
	) name2412 (
		_w2235_,
		_w2311_,
		_w2312_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('h000d)
	) name2413 (
		_w2235_,
		_w2311_,
		_w2312_,
		_w2477_,
		_w2479_
	);
	LUT4 #(
		.INIT('h0df2)
	) name2414 (
		_w2235_,
		_w2311_,
		_w2312_,
		_w2477_,
		_w2480_
	);
	LUT3 #(
		.INIT('h0d)
	) name2415 (
		_w2304_,
		_w2305_,
		_w2307_,
		_w2481_
	);
	LUT2 #(
		.INIT('h6)
	) name2416 (
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT3 #(
		.INIT('h69)
	) name2417 (
		_w2474_,
		_w2475_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		_w2473_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name2419 (
		_w2473_,
		_w2483_,
		_w2485_
	);
	LUT2 #(
		.INIT('h6)
	) name2420 (
		_w2473_,
		_w2483_,
		_w2486_
	);
	LUT2 #(
		.INIT('h6)
	) name2421 (
		_w2431_,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('h7500)
	) name2422 (
		_w2334_,
		_w2335_,
		_w2362_,
		_w2487_,
		_w2488_
	);
	LUT4 #(
		.INIT('h008a)
	) name2423 (
		_w2334_,
		_w2335_,
		_w2362_,
		_w2487_,
		_w2489_
	);
	LUT4 #(
		.INIT('hf20d)
	) name2424 (
		_w2334_,
		_w2362_,
		_w2335_,
		_w2487_,
		_w2490_
	);
	LUT2 #(
		.INIT('h6)
	) name2425 (
		_w2417_,
		_w2490_,
		_w2491_
	);
	LUT3 #(
		.INIT('he0)
	) name2426 (
		_w2387_,
		_w2404_,
		_w2491_,
		_w2492_
	);
	LUT3 #(
		.INIT('h01)
	) name2427 (
		_w2387_,
		_w2404_,
		_w2491_,
		_w2493_
	);
	LUT3 #(
		.INIT('h1e)
	) name2428 (
		_w2387_,
		_w2404_,
		_w2491_,
		_w2494_
	);
	LUT4 #(
		.INIT('hfd02)
	) name2429 (
		_w2393_,
		_w2402_,
		_w2403_,
		_w2494_,
		_w2495_
	);
	LUT3 #(
		.INIT('h02)
	) name2430 (
		_w2393_,
		_w2403_,
		_w2493_,
		_w2496_
	);
	LUT3 #(
		.INIT('h31)
	) name2431 (
		_w2417_,
		_w2488_,
		_w2489_,
		_w2497_
	);
	LUT3 #(
		.INIT('h71)
	) name2432 (
		_w2405_,
		_w2406_,
		_w2416_,
		_w2498_
	);
	LUT3 #(
		.INIT('h17)
	) name2433 (
		_w2412_,
		_w2413_,
		_w2415_,
		_w2499_
	);
	LUT3 #(
		.INIT('he8)
	) name2434 (
		_w2428_,
		_w2429_,
		_w2430_,
		_w2500_
	);
	LUT2 #(
		.INIT('h8)
	) name2435 (
		\a[7] ,
		\a[41] ,
		_w2501_
	);
	LUT4 #(
		.INIT('h153f)
	) name2436 (
		\a[8] ,
		\a[12] ,
		\a[36] ,
		\a[40] ,
		_w2502_
	);
	LUT4 #(
		.INIT('h8000)
	) name2437 (
		\a[8] ,
		\a[12] ,
		\a[36] ,
		\a[40] ,
		_w2503_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2438 (
		\a[8] ,
		\a[12] ,
		\a[36] ,
		\a[40] ,
		_w2504_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		\a[14] ,
		\a[34] ,
		_w2505_
	);
	LUT4 #(
		.INIT('h153f)
	) name2440 (
		\a[6] ,
		\a[13] ,
		\a[35] ,
		\a[42] ,
		_w2506_
	);
	LUT4 #(
		.INIT('h8000)
	) name2441 (
		\a[6] ,
		\a[13] ,
		\a[35] ,
		\a[42] ,
		_w2507_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2442 (
		\a[6] ,
		\a[13] ,
		\a[35] ,
		\a[42] ,
		_w2508_
	);
	LUT4 #(
		.INIT('h0660)
	) name2443 (
		_w2501_,
		_w2504_,
		_w2505_,
		_w2508_,
		_w2509_
	);
	LUT4 #(
		.INIT('h9009)
	) name2444 (
		_w2501_,
		_w2504_,
		_w2505_,
		_w2508_,
		_w2510_
	);
	LUT4 #(
		.INIT('h6996)
	) name2445 (
		_w2501_,
		_w2504_,
		_w2505_,
		_w2508_,
		_w2511_
	);
	LUT2 #(
		.INIT('h8)
	) name2446 (
		\a[9] ,
		\a[39] ,
		_w2512_
	);
	LUT4 #(
		.INIT('h153f)
	) name2447 (
		\a[10] ,
		\a[11] ,
		\a[37] ,
		\a[38] ,
		_w2513_
	);
	LUT4 #(
		.INIT('h8000)
	) name2448 (
		\a[10] ,
		\a[11] ,
		\a[37] ,
		\a[38] ,
		_w2514_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2449 (
		\a[10] ,
		\a[11] ,
		\a[37] ,
		\a[38] ,
		_w2515_
	);
	LUT2 #(
		.INIT('h6)
	) name2450 (
		_w2512_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h6)
	) name2451 (
		_w2511_,
		_w2516_,
		_w2517_
	);
	LUT4 #(
		.INIT('h0017)
	) name2452 (
		_w2418_,
		_w2419_,
		_w2424_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('he800)
	) name2453 (
		_w2418_,
		_w2419_,
		_w2424_,
		_w2517_,
		_w2519_
	);
	LUT4 #(
		.INIT('hf10e)
	) name2454 (
		_w2418_,
		_w2425_,
		_w2426_,
		_w2517_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name2455 (
		\a[4] ,
		\a[44] ,
		_w2521_
	);
	LUT4 #(
		.INIT('h153f)
	) name2456 (
		\a[5] ,
		\a[15] ,
		\a[33] ,
		\a[43] ,
		_w2522_
	);
	LUT4 #(
		.INIT('h8000)
	) name2457 (
		\a[5] ,
		\a[15] ,
		\a[33] ,
		\a[43] ,
		_w2523_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2458 (
		\a[5] ,
		\a[15] ,
		\a[33] ,
		\a[43] ,
		_w2524_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		\a[20] ,
		\a[28] ,
		_w2525_
	);
	LUT4 #(
		.INIT('h153f)
	) name2460 (
		\a[21] ,
		\a[22] ,
		\a[26] ,
		\a[27] ,
		_w2526_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		\a[22] ,
		\a[27] ,
		_w2527_
	);
	LUT4 #(
		.INIT('h8000)
	) name2462 (
		\a[21] ,
		\a[22] ,
		\a[26] ,
		\a[27] ,
		_w2528_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2463 (
		\a[21] ,
		\a[22] ,
		\a[26] ,
		\a[27] ,
		_w2529_
	);
	LUT4 #(
		.INIT('h0660)
	) name2464 (
		_w2521_,
		_w2524_,
		_w2525_,
		_w2529_,
		_w2530_
	);
	LUT4 #(
		.INIT('h9009)
	) name2465 (
		_w2521_,
		_w2524_,
		_w2525_,
		_w2529_,
		_w2531_
	);
	LUT4 #(
		.INIT('h6996)
	) name2466 (
		_w2521_,
		_w2524_,
		_w2525_,
		_w2529_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name2467 (
		\a[17] ,
		\a[31] ,
		_w2533_
	);
	LUT4 #(
		.INIT('h153f)
	) name2468 (
		\a[18] ,
		\a[19] ,
		\a[29] ,
		\a[30] ,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		\a[19] ,
		\a[30] ,
		_w2535_
	);
	LUT4 #(
		.INIT('h8000)
	) name2470 (
		\a[18] ,
		\a[19] ,
		\a[29] ,
		\a[30] ,
		_w2536_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2471 (
		\a[18] ,
		\a[19] ,
		\a[29] ,
		\a[30] ,
		_w2537_
	);
	LUT2 #(
		.INIT('h6)
	) name2472 (
		_w2533_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h6)
	) name2473 (
		_w2532_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h6)
	) name2474 (
		_w2520_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h6)
	) name2475 (
		_w2500_,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h6)
	) name2476 (
		_w2499_,
		_w2541_,
		_w2542_
	);
	LUT3 #(
		.INIT('h0d)
	) name2477 (
		_w2467_,
		_w2468_,
		_w2469_,
		_w2543_
	);
	LUT3 #(
		.INIT('h0d)
	) name2478 (
		_w2306_,
		_w2440_,
		_w2442_,
		_w2544_
	);
	LUT3 #(
		.INIT('h0d)
	) name2479 (
		_w2451_,
		_w2452_,
		_w2453_,
		_w2545_
	);
	LUT3 #(
		.INIT('h96)
	) name2480 (
		_w2543_,
		_w2544_,
		_w2545_,
		_w2546_
	);
	LUT3 #(
		.INIT('h32)
	) name2481 (
		_w2448_,
		_w2449_,
		_w2455_,
		_w2547_
	);
	LUT3 #(
		.INIT('h0d)
	) name2482 (
		_w2420_,
		_w2421_,
		_w2422_,
		_w2548_
	);
	LUT3 #(
		.INIT('h0d)
	) name2483 (
		_w2444_,
		_w2445_,
		_w2446_,
		_w2549_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		\a[2] ,
		\a[46] ,
		_w2550_
	);
	LUT4 #(
		.INIT('h153f)
	) name2485 (
		\a[3] ,
		\a[16] ,
		\a[32] ,
		\a[45] ,
		_w2551_
	);
	LUT4 #(
		.INIT('h8000)
	) name2486 (
		\a[3] ,
		\a[16] ,
		\a[32] ,
		\a[45] ,
		_w2552_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2487 (
		\a[3] ,
		\a[16] ,
		\a[32] ,
		\a[45] ,
		_w2553_
	);
	LUT2 #(
		.INIT('h6)
	) name2488 (
		_w2550_,
		_w2553_,
		_w2554_
	);
	LUT3 #(
		.INIT('h69)
	) name2489 (
		_w2548_,
		_w2549_,
		_w2554_,
		_w2555_
	);
	LUT3 #(
		.INIT('h96)
	) name2490 (
		_w2546_,
		_w2547_,
		_w2555_,
		_w2556_
	);
	LUT3 #(
		.INIT('he8)
	) name2491 (
		_w2439_,
		_w2456_,
		_w2472_,
		_w2557_
	);
	LUT3 #(
		.INIT('h0d)
	) name2492 (
		_w2460_,
		_w2461_,
		_w2462_,
		_w2558_
	);
	LUT3 #(
		.INIT('h0d)
	) name2493 (
		_w2434_,
		_w2435_,
		_w2436_,
		_w2559_
	);
	LUT3 #(
		.INIT('h0d)
	) name2494 (
		_w2345_,
		_w2457_,
		_w2458_,
		_w2560_
	);
	LUT3 #(
		.INIT('h96)
	) name2495 (
		_w2558_,
		_w2559_,
		_w2560_,
		_w2561_
	);
	LUT3 #(
		.INIT('h23)
	) name2496 (
		_w2478_,
		_w2479_,
		_w2481_,
		_w2562_
	);
	LUT3 #(
		.INIT('h32)
	) name2497 (
		_w2464_,
		_w2465_,
		_w2471_,
		_w2563_
	);
	LUT3 #(
		.INIT('h69)
	) name2498 (
		_w2561_,
		_w2562_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h96)
	) name2499 (
		_w2556_,
		_w2557_,
		_w2564_,
		_w2565_
	);
	LUT3 #(
		.INIT('h0e)
	) name2500 (
		_w2431_,
		_w2484_,
		_w2485_,
		_w2566_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2501 (
		_w2379_,
		_w2381_,
		_w2410_,
		_w2411_,
		_w2567_
	);
	LUT3 #(
		.INIT('h8e)
	) name2502 (
		_w2474_,
		_w2475_,
		_w2482_,
		_w2568_
	);
	LUT4 #(
		.INIT('h8000)
	) name2503 (
		\a[1] ,
		\a[23] ,
		\a[25] ,
		\a[47] ,
		_w2569_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2504 (
		\a[1] ,
		\a[23] ,
		\a[25] ,
		\a[47] ,
		_w2570_
	);
	LUT2 #(
		.INIT('h8)
	) name2505 (
		\a[0] ,
		\a[48] ,
		_w2571_
	);
	LUT3 #(
		.INIT('h96)
	) name2506 (
		_w2476_,
		_w2570_,
		_w2571_,
		_w2572_
	);
	LUT4 #(
		.INIT('h008e)
	) name2507 (
		_w2407_,
		_w2408_,
		_w2409_,
		_w2572_,
		_w2573_
	);
	LUT4 #(
		.INIT('h7100)
	) name2508 (
		_w2407_,
		_w2408_,
		_w2409_,
		_w2572_,
		_w2574_
	);
	LUT4 #(
		.INIT('h8e71)
	) name2509 (
		_w2407_,
		_w2408_,
		_w2409_,
		_w2572_,
		_w2575_
	);
	LUT3 #(
		.INIT('hb2)
	) name2510 (
		_w2432_,
		_w2433_,
		_w2438_,
		_w2576_
	);
	LUT2 #(
		.INIT('h6)
	) name2511 (
		_w2575_,
		_w2576_,
		_w2577_
	);
	LUT3 #(
		.INIT('h96)
	) name2512 (
		_w2567_,
		_w2568_,
		_w2577_,
		_w2578_
	);
	LUT4 #(
		.INIT('he800)
	) name2513 (
		_w2431_,
		_w2473_,
		_w2483_,
		_w2578_,
		_w2579_
	);
	LUT4 #(
		.INIT('h0017)
	) name2514 (
		_w2431_,
		_w2473_,
		_w2483_,
		_w2578_,
		_w2580_
	);
	LUT4 #(
		.INIT('hf10e)
	) name2515 (
		_w2431_,
		_w2484_,
		_w2485_,
		_w2578_,
		_w2581_
	);
	LUT2 #(
		.INIT('h6)
	) name2516 (
		_w2565_,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('h96)
	) name2517 (
		_w2498_,
		_w2542_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h4)
	) name2518 (
		_w2497_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h9)
	) name2519 (
		_w2497_,
		_w2583_,
		_w2585_
	);
	LUT4 #(
		.INIT('h23dc)
	) name2520 (
		_w2402_,
		_w2492_,
		_w2496_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name2521 (
		_w2492_,
		_w2584_,
		_w2587_
	);
	LUT3 #(
		.INIT('he8)
	) name2522 (
		_w2556_,
		_w2557_,
		_w2564_,
		_w2588_
	);
	LUT3 #(
		.INIT('he8)
	) name2523 (
		_w2567_,
		_w2568_,
		_w2577_,
		_w2589_
	);
	LUT3 #(
		.INIT('he8)
	) name2524 (
		_w2476_,
		_w2570_,
		_w2571_,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		\a[0] ,
		\a[49] ,
		_w2591_
	);
	LUT4 #(
		.INIT('h153f)
	) name2526 (
		\a[4] ,
		\a[5] ,
		\a[44] ,
		\a[45] ,
		_w2592_
	);
	LUT4 #(
		.INIT('h8000)
	) name2527 (
		\a[4] ,
		\a[5] ,
		\a[44] ,
		\a[45] ,
		_w2593_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2528 (
		\a[4] ,
		\a[5] ,
		\a[44] ,
		\a[45] ,
		_w2594_
	);
	LUT2 #(
		.INIT('h6)
	) name2529 (
		_w2591_,
		_w2594_,
		_w2595_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		\a[16] ,
		\a[33] ,
		_w2596_
	);
	LUT4 #(
		.INIT('h153f)
	) name2531 (
		\a[17] ,
		\a[18] ,
		\a[31] ,
		\a[32] ,
		_w2597_
	);
	LUT4 #(
		.INIT('h8000)
	) name2532 (
		\a[17] ,
		\a[18] ,
		\a[31] ,
		\a[32] ,
		_w2598_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2533 (
		\a[17] ,
		\a[18] ,
		\a[31] ,
		\a[32] ,
		_w2599_
	);
	LUT2 #(
		.INIT('h6)
	) name2534 (
		_w2596_,
		_w2599_,
		_w2600_
	);
	LUT3 #(
		.INIT('h96)
	) name2535 (
		_w2590_,
		_w2595_,
		_w2600_,
		_w2601_
	);
	LUT4 #(
		.INIT('h153f)
	) name2536 (
		\a[2] ,
		\a[3] ,
		\a[46] ,
		\a[47] ,
		_w2602_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		\a[3] ,
		\a[47] ,
		_w2603_
	);
	LUT4 #(
		.INIT('h8000)
	) name2538 (
		\a[2] ,
		\a[3] ,
		\a[46] ,
		\a[47] ,
		_w2604_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2539 (
		\a[2] ,
		\a[3] ,
		\a[46] ,
		\a[47] ,
		_w2605_
	);
	LUT4 #(
		.INIT('h153f)
	) name2540 (
		\a[20] ,
		\a[21] ,
		\a[28] ,
		\a[29] ,
		_w2606_
	);
	LUT4 #(
		.INIT('h8000)
	) name2541 (
		\a[20] ,
		\a[21] ,
		\a[28] ,
		\a[29] ,
		_w2607_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2542 (
		\a[20] ,
		\a[21] ,
		\a[28] ,
		\a[29] ,
		_w2608_
	);
	LUT4 #(
		.INIT('h1248)
	) name2543 (
		_w2527_,
		_w2535_,
		_w2605_,
		_w2608_,
		_w2609_
	);
	LUT4 #(
		.INIT('h8421)
	) name2544 (
		_w2527_,
		_w2535_,
		_w2605_,
		_w2608_,
		_w2610_
	);
	LUT4 #(
		.INIT('h6996)
	) name2545 (
		_w2527_,
		_w2535_,
		_w2605_,
		_w2608_,
		_w2611_
	);
	LUT2 #(
		.INIT('h8)
	) name2546 (
		\a[9] ,
		\a[40] ,
		_w2612_
	);
	LUT4 #(
		.INIT('h153f)
	) name2547 (
		\a[10] ,
		\a[12] ,
		\a[37] ,
		\a[39] ,
		_w2613_
	);
	LUT4 #(
		.INIT('h8000)
	) name2548 (
		\a[10] ,
		\a[12] ,
		\a[37] ,
		\a[39] ,
		_w2614_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2549 (
		\a[10] ,
		\a[12] ,
		\a[37] ,
		\a[39] ,
		_w2615_
	);
	LUT2 #(
		.INIT('h6)
	) name2550 (
		_w2612_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h6)
	) name2551 (
		_w2611_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h8)
	) name2552 (
		\a[13] ,
		\a[36] ,
		_w2618_
	);
	LUT4 #(
		.INIT('h153f)
	) name2553 (
		\a[7] ,
		\a[8] ,
		\a[41] ,
		\a[42] ,
		_w2619_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		\a[8] ,
		\a[42] ,
		_w2620_
	);
	LUT4 #(
		.INIT('h8000)
	) name2555 (
		\a[7] ,
		\a[8] ,
		\a[41] ,
		\a[42] ,
		_w2621_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2556 (
		\a[7] ,
		\a[8] ,
		\a[41] ,
		\a[42] ,
		_w2622_
	);
	LUT2 #(
		.INIT('h8)
	) name2557 (
		\a[24] ,
		\a[25] ,
		_w2623_
	);
	LUT2 #(
		.INIT('h8)
	) name2558 (
		\a[23] ,
		\a[26] ,
		_w2624_
	);
	LUT4 #(
		.INIT('h153f)
	) name2559 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w2625_
	);
	LUT4 #(
		.INIT('h8000)
	) name2560 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w2626_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2561 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w2627_
	);
	LUT4 #(
		.INIT('h1428)
	) name2562 (
		_w2441_,
		_w2618_,
		_w2622_,
		_w2627_,
		_w2628_
	);
	LUT4 #(
		.INIT('h8241)
	) name2563 (
		_w2441_,
		_w2618_,
		_w2622_,
		_w2627_,
		_w2629_
	);
	LUT4 #(
		.INIT('h6996)
	) name2564 (
		_w2441_,
		_w2618_,
		_w2622_,
		_w2627_,
		_w2630_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		\a[15] ,
		\a[34] ,
		_w2631_
	);
	LUT4 #(
		.INIT('h153f)
	) name2566 (
		\a[6] ,
		\a[14] ,
		\a[35] ,
		\a[43] ,
		_w2632_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		\a[14] ,
		\a[43] ,
		_w2633_
	);
	LUT4 #(
		.INIT('h8000)
	) name2568 (
		\a[6] ,
		\a[14] ,
		\a[35] ,
		\a[43] ,
		_w2634_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2569 (
		\a[6] ,
		\a[14] ,
		\a[35] ,
		\a[43] ,
		_w2635_
	);
	LUT2 #(
		.INIT('h6)
	) name2570 (
		_w2631_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h6)
	) name2571 (
		_w2630_,
		_w2636_,
		_w2637_
	);
	LUT3 #(
		.INIT('h96)
	) name2572 (
		_w2601_,
		_w2617_,
		_w2637_,
		_w2638_
	);
	LUT4 #(
		.INIT('he800)
	) name2573 (
		_w2567_,
		_w2568_,
		_w2577_,
		_w2638_,
		_w2639_
	);
	LUT4 #(
		.INIT('h0017)
	) name2574 (
		_w2567_,
		_w2568_,
		_w2577_,
		_w2638_,
		_w2640_
	);
	LUT4 #(
		.INIT('h17e8)
	) name2575 (
		_w2567_,
		_w2568_,
		_w2577_,
		_w2638_,
		_w2641_
	);
	LUT2 #(
		.INIT('h6)
	) name2576 (
		_w2588_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('he800)
	) name2577 (
		_w2565_,
		_w2566_,
		_w2578_,
		_w2642_,
		_w2643_
	);
	LUT4 #(
		.INIT('h0017)
	) name2578 (
		_w2565_,
		_w2566_,
		_w2578_,
		_w2642_,
		_w2644_
	);
	LUT4 #(
		.INIT('hf10e)
	) name2579 (
		_w2565_,
		_w2579_,
		_w2580_,
		_w2642_,
		_w2645_
	);
	LUT3 #(
		.INIT('h17)
	) name2580 (
		_w2543_,
		_w2544_,
		_w2545_,
		_w2646_
	);
	LUT3 #(
		.INIT('h8e)
	) name2581 (
		_w2548_,
		_w2549_,
		_w2554_,
		_w2647_
	);
	LUT3 #(
		.INIT('h17)
	) name2582 (
		_w2558_,
		_w2559_,
		_w2560_,
		_w2648_
	);
	LUT3 #(
		.INIT('h69)
	) name2583 (
		_w2646_,
		_w2647_,
		_w2648_,
		_w2649_
	);
	LUT3 #(
		.INIT('h4d)
	) name2584 (
		_w2546_,
		_w2547_,
		_w2555_,
		_w2650_
	);
	LUT3 #(
		.INIT('hd4)
	) name2585 (
		_w2561_,
		_w2562_,
		_w2563_,
		_w2651_
	);
	LUT3 #(
		.INIT('h96)
	) name2586 (
		_w2649_,
		_w2650_,
		_w2651_,
		_w2652_
	);
	LUT4 #(
		.INIT('he800)
	) name2587 (
		_w2499_,
		_w2500_,
		_w2540_,
		_w2652_,
		_w2653_
	);
	LUT3 #(
		.INIT('h32)
	) name2588 (
		_w2505_,
		_w2506_,
		_w2507_,
		_w2654_
	);
	LUT3 #(
		.INIT('h0d)
	) name2589 (
		_w2533_,
		_w2534_,
		_w2536_,
		_w2655_
	);
	LUT3 #(
		.INIT('h0d)
	) name2590 (
		_w2501_,
		_w2502_,
		_w2503_,
		_w2656_
	);
	LUT3 #(
		.INIT('h69)
	) name2591 (
		_w2654_,
		_w2655_,
		_w2656_,
		_w2657_
	);
	LUT3 #(
		.INIT('h32)
	) name2592 (
		_w2530_,
		_w2531_,
		_w2538_,
		_w2658_
	);
	LUT2 #(
		.INIT('h2)
	) name2593 (
		_w2657_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h4)
	) name2594 (
		_w2657_,
		_w2658_,
		_w2660_
	);
	LUT2 #(
		.INIT('h9)
	) name2595 (
		_w2657_,
		_w2658_,
		_w2661_
	);
	LUT3 #(
		.INIT('h54)
	) name2596 (
		_w2573_,
		_w2574_,
		_w2576_,
		_w2662_
	);
	LUT2 #(
		.INIT('h6)
	) name2597 (
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT3 #(
		.INIT('h54)
	) name2598 (
		_w2518_,
		_w2519_,
		_w2539_,
		_w2664_
	);
	LUT3 #(
		.INIT('h32)
	) name2599 (
		_w2550_,
		_w2551_,
		_w2552_,
		_w2665_
	);
	LUT3 #(
		.INIT('h0d)
	) name2600 (
		_w2521_,
		_w2522_,
		_w2523_,
		_w2666_
	);
	LUT3 #(
		.INIT('h0d)
	) name2601 (
		_w2525_,
		_w2526_,
		_w2528_,
		_w2667_
	);
	LUT3 #(
		.INIT('h69)
	) name2602 (
		_w2665_,
		_w2666_,
		_w2667_,
		_w2668_
	);
	LUT3 #(
		.INIT('h32)
	) name2603 (
		_w2509_,
		_w2510_,
		_w2516_,
		_w2669_
	);
	LUT3 #(
		.INIT('h80)
	) name2604 (
		\a[1] ,
		\a[25] ,
		\a[48] ,
		_w2670_
	);
	LUT3 #(
		.INIT('h6c)
	) name2605 (
		\a[1] ,
		\a[25] ,
		\a[48] ,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w2569_,
		_w2671_,
		_w2672_
	);
	LUT2 #(
		.INIT('h4)
	) name2607 (
		\a[48] ,
		_w2569_,
		_w2673_
	);
	LUT3 #(
		.INIT('hb8)
	) name2608 (
		\a[48] ,
		_w2569_,
		_w2671_,
		_w2674_
	);
	LUT3 #(
		.INIT('h0d)
	) name2609 (
		_w2512_,
		_w2513_,
		_w2514_,
		_w2675_
	);
	LUT2 #(
		.INIT('h6)
	) name2610 (
		_w2674_,
		_w2675_,
		_w2676_
	);
	LUT3 #(
		.INIT('h96)
	) name2611 (
		_w2668_,
		_w2669_,
		_w2676_,
		_w2677_
	);
	LUT3 #(
		.INIT('h96)
	) name2612 (
		_w2663_,
		_w2664_,
		_w2677_,
		_w2678_
	);
	LUT3 #(
		.INIT('h07)
	) name2613 (
		_w2500_,
		_w2540_,
		_w2652_,
		_w2679_
	);
	LUT4 #(
		.INIT('h80f0)
	) name2614 (
		_w2499_,
		_w2541_,
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT4 #(
		.INIT('h0700)
	) name2615 (
		_w2499_,
		_w2541_,
		_w2678_,
		_w2679_,
		_w2681_
	);
	LUT4 #(
		.INIT('h2882)
	) name2616 (
		_w2652_,
		_w2663_,
		_w2664_,
		_w2677_,
		_w2682_
	);
	LUT4 #(
		.INIT('he800)
	) name2617 (
		_w2499_,
		_w2500_,
		_w2540_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('h000b)
	) name2618 (
		_w2653_,
		_w2680_,
		_w2681_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h6)
	) name2619 (
		_w2645_,
		_w2684_,
		_w2685_
	);
	LUT3 #(
		.INIT('he8)
	) name2620 (
		_w2498_,
		_w2542_,
		_w2582_,
		_w2686_
	);
	LUT2 #(
		.INIT('h8)
	) name2621 (
		_w2685_,
		_w2686_,
		_w2687_
	);
	LUT4 #(
		.INIT('hd22d)
	) name2622 (
		_w2497_,
		_w2583_,
		_w2685_,
		_w2686_,
		_w2688_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2623 (
		_w2402_,
		_w2496_,
		_w2587_,
		_w2688_,
		_w2689_
	);
	LUT4 #(
		.INIT('h0ff0)
	) name2624 (
		_w2497_,
		_w2583_,
		_w2685_,
		_w2686_,
		_w2690_
	);
	LUT4 #(
		.INIT('hb000)
	) name2625 (
		_w2402_,
		_w2496_,
		_w2587_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('he)
	) name2626 (
		_w2689_,
		_w2691_,
		_w2692_
	);
	LUT3 #(
		.INIT('h01)
	) name2627 (
		_w2492_,
		_w2584_,
		_w2687_,
		_w2693_
	);
	LUT4 #(
		.INIT('h0222)
	) name2628 (
		_w2497_,
		_w2583_,
		_w2685_,
		_w2686_,
		_w2694_
	);
	LUT3 #(
		.INIT('h45)
	) name2629 (
		_w2643_,
		_w2644_,
		_w2684_,
		_w2695_
	);
	LUT2 #(
		.INIT('h1)
	) name2630 (
		_w2653_,
		_w2680_,
		_w2696_
	);
	LUT2 #(
		.INIT('h8)
	) name2631 (
		\a[16] ,
		\a[34] ,
		_w2697_
	);
	LUT4 #(
		.INIT('h153f)
	) name2632 (
		\a[5] ,
		\a[15] ,
		\a[35] ,
		\a[45] ,
		_w2698_
	);
	LUT4 #(
		.INIT('h8000)
	) name2633 (
		\a[5] ,
		\a[15] ,
		\a[35] ,
		\a[45] ,
		_w2699_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2634 (
		\a[5] ,
		\a[15] ,
		\a[35] ,
		\a[45] ,
		_w2700_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		\a[22] ,
		\a[28] ,
		_w2701_
	);
	LUT4 #(
		.INIT('h153f)
	) name2636 (
		\a[18] ,
		\a[23] ,
		\a[27] ,
		\a[32] ,
		_w2702_
	);
	LUT4 #(
		.INIT('h8000)
	) name2637 (
		\a[18] ,
		\a[23] ,
		\a[27] ,
		\a[32] ,
		_w2703_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2638 (
		\a[18] ,
		\a[23] ,
		\a[27] ,
		\a[32] ,
		_w2704_
	);
	LUT4 #(
		.INIT('h0660)
	) name2639 (
		_w2697_,
		_w2700_,
		_w2701_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('h9009)
	) name2640 (
		_w2697_,
		_w2700_,
		_w2701_,
		_w2704_,
		_w2706_
	);
	LUT4 #(
		.INIT('h6996)
	) name2641 (
		_w2697_,
		_w2700_,
		_w2701_,
		_w2704_,
		_w2707_
	);
	LUT4 #(
		.INIT('hba45)
	) name2642 (
		_w2672_,
		_w2673_,
		_w2675_,
		_w2707_,
		_w2708_
	);
	LUT4 #(
		.INIT('h153f)
	) name2643 (
		\a[4] ,
		\a[17] ,
		\a[33] ,
		\a[46] ,
		_w2709_
	);
	LUT4 #(
		.INIT('h8000)
	) name2644 (
		\a[4] ,
		\a[17] ,
		\a[33] ,
		\a[46] ,
		_w2710_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2645 (
		\a[4] ,
		\a[17] ,
		\a[33] ,
		\a[46] ,
		_w2711_
	);
	LUT4 #(
		.INIT('h153f)
	) name2646 (
		\a[0] ,
		\a[2] ,
		\a[48] ,
		\a[50] ,
		_w2712_
	);
	LUT4 #(
		.INIT('h8000)
	) name2647 (
		\a[0] ,
		\a[2] ,
		\a[48] ,
		\a[50] ,
		_w2713_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2648 (
		\a[0] ,
		\a[2] ,
		\a[48] ,
		\a[50] ,
		_w2714_
	);
	LUT4 #(
		.INIT('h1248)
	) name2649 (
		_w2603_,
		_w2670_,
		_w2711_,
		_w2714_,
		_w2715_
	);
	LUT4 #(
		.INIT('h8421)
	) name2650 (
		_w2603_,
		_w2670_,
		_w2711_,
		_w2714_,
		_w2716_
	);
	LUT4 #(
		.INIT('h6996)
	) name2651 (
		_w2603_,
		_w2670_,
		_w2711_,
		_w2714_,
		_w2717_
	);
	LUT2 #(
		.INIT('h8)
	) name2652 (
		\a[19] ,
		\a[31] ,
		_w2718_
	);
	LUT4 #(
		.INIT('h153f)
	) name2653 (
		\a[20] ,
		\a[21] ,
		\a[29] ,
		\a[30] ,
		_w2719_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		\a[21] ,
		\a[30] ,
		_w2720_
	);
	LUT4 #(
		.INIT('h8000)
	) name2655 (
		\a[20] ,
		\a[21] ,
		\a[29] ,
		\a[30] ,
		_w2721_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2656 (
		\a[20] ,
		\a[21] ,
		\a[29] ,
		\a[30] ,
		_w2722_
	);
	LUT2 #(
		.INIT('h6)
	) name2657 (
		_w2718_,
		_w2722_,
		_w2723_
	);
	LUT4 #(
		.INIT('h153f)
	) name2658 (
		\a[9] ,
		\a[13] ,
		\a[37] ,
		\a[41] ,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name2659 (
		\a[13] ,
		\a[41] ,
		_w2725_
	);
	LUT4 #(
		.INIT('h8000)
	) name2660 (
		\a[9] ,
		\a[13] ,
		\a[37] ,
		\a[41] ,
		_w2726_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2661 (
		\a[9] ,
		\a[13] ,
		\a[37] ,
		\a[41] ,
		_w2727_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		\a[6] ,
		\a[44] ,
		_w2728_
	);
	LUT4 #(
		.INIT('h153f)
	) name2663 (
		\a[7] ,
		\a[14] ,
		\a[36] ,
		\a[43] ,
		_w2729_
	);
	LUT4 #(
		.INIT('h8000)
	) name2664 (
		\a[7] ,
		\a[14] ,
		\a[36] ,
		\a[43] ,
		_w2730_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2665 (
		\a[7] ,
		\a[14] ,
		\a[36] ,
		\a[43] ,
		_w2731_
	);
	LUT4 #(
		.INIT('h0660)
	) name2666 (
		_w2620_,
		_w2727_,
		_w2728_,
		_w2731_,
		_w2732_
	);
	LUT4 #(
		.INIT('h9009)
	) name2667 (
		_w2620_,
		_w2727_,
		_w2728_,
		_w2731_,
		_w2733_
	);
	LUT4 #(
		.INIT('h6996)
	) name2668 (
		_w2620_,
		_w2727_,
		_w2728_,
		_w2731_,
		_w2734_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		\a[12] ,
		\a[38] ,
		_w2735_
	);
	LUT4 #(
		.INIT('h153f)
	) name2670 (
		\a[10] ,
		\a[11] ,
		\a[39] ,
		\a[40] ,
		_w2736_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		\a[11] ,
		\a[40] ,
		_w2737_
	);
	LUT4 #(
		.INIT('h8000)
	) name2672 (
		\a[10] ,
		\a[11] ,
		\a[39] ,
		\a[40] ,
		_w2738_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2673 (
		\a[10] ,
		\a[11] ,
		\a[39] ,
		\a[40] ,
		_w2739_
	);
	LUT2 #(
		.INIT('h6)
	) name2674 (
		_w2735_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('h0660)
	) name2675 (
		_w2717_,
		_w2723_,
		_w2734_,
		_w2740_,
		_w2741_
	);
	LUT4 #(
		.INIT('h9009)
	) name2676 (
		_w2717_,
		_w2723_,
		_w2734_,
		_w2740_,
		_w2742_
	);
	LUT4 #(
		.INIT('h6996)
	) name2677 (
		_w2717_,
		_w2723_,
		_w2734_,
		_w2740_,
		_w2743_
	);
	LUT2 #(
		.INIT('h6)
	) name2678 (
		_w2708_,
		_w2743_,
		_w2744_
	);
	LUT4 #(
		.INIT('he800)
	) name2679 (
		_w2649_,
		_w2650_,
		_w2651_,
		_w2744_,
		_w2745_
	);
	LUT4 #(
		.INIT('h0017)
	) name2680 (
		_w2649_,
		_w2650_,
		_w2651_,
		_w2744_,
		_w2746_
	);
	LUT4 #(
		.INIT('h17e8)
	) name2681 (
		_w2649_,
		_w2650_,
		_w2651_,
		_w2744_,
		_w2747_
	);
	LUT4 #(
		.INIT('h17e8)
	) name2682 (
		_w2663_,
		_w2664_,
		_w2677_,
		_w2747_,
		_w2748_
	);
	LUT3 #(
		.INIT('he0)
	) name2683 (
		_w2653_,
		_w2680_,
		_w2748_,
		_w2749_
	);
	LUT3 #(
		.INIT('h01)
	) name2684 (
		_w2653_,
		_w2680_,
		_w2748_,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w2588_,
		_w2639_,
		_w2751_
	);
	LUT3 #(
		.INIT('h0e)
	) name2686 (
		_w2588_,
		_w2639_,
		_w2640_,
		_w2752_
	);
	LUT3 #(
		.INIT('he8)
	) name2687 (
		_w2590_,
		_w2595_,
		_w2600_,
		_w2753_
	);
	LUT3 #(
		.INIT('h32)
	) name2688 (
		_w2609_,
		_w2610_,
		_w2616_,
		_w2754_
	);
	LUT4 #(
		.INIT('h8000)
	) name2689 (
		\a[1] ,
		\a[24] ,
		\a[26] ,
		\a[49] ,
		_w2755_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2690 (
		\a[1] ,
		\a[24] ,
		\a[26] ,
		\a[49] ,
		_w2756_
	);
	LUT4 #(
		.INIT('h0017)
	) name2691 (
		_w2441_,
		_w2623_,
		_w2624_,
		_w2756_,
		_w2757_
	);
	LUT4 #(
		.INIT('he800)
	) name2692 (
		_w2441_,
		_w2623_,
		_w2624_,
		_w2756_,
		_w2758_
	);
	LUT4 #(
		.INIT('hcd32)
	) name2693 (
		_w2441_,
		_w2625_,
		_w2626_,
		_w2756_,
		_w2759_
	);
	LUT3 #(
		.INIT('h0d)
	) name2694 (
		_w2612_,
		_w2613_,
		_w2614_,
		_w2760_
	);
	LUT2 #(
		.INIT('h6)
	) name2695 (
		_w2759_,
		_w2760_,
		_w2761_
	);
	LUT3 #(
		.INIT('h69)
	) name2696 (
		_w2753_,
		_w2754_,
		_w2761_,
		_w2762_
	);
	LUT3 #(
		.INIT('h0d)
	) name2697 (
		_w2535_,
		_w2606_,
		_w2607_,
		_w2763_
	);
	LUT3 #(
		.INIT('h0d)
	) name2698 (
		_w2596_,
		_w2597_,
		_w2598_,
		_w2764_
	);
	LUT3 #(
		.INIT('h0d)
	) name2699 (
		_w2618_,
		_w2619_,
		_w2621_,
		_w2765_
	);
	LUT3 #(
		.INIT('h96)
	) name2700 (
		_w2763_,
		_w2764_,
		_w2765_,
		_w2766_
	);
	LUT3 #(
		.INIT('h32)
	) name2701 (
		_w2628_,
		_w2629_,
		_w2636_,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name2702 (
		_w2766_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h4)
	) name2703 (
		_w2766_,
		_w2767_,
		_w2769_
	);
	LUT2 #(
		.INIT('h9)
	) name2704 (
		_w2766_,
		_w2767_,
		_w2770_
	);
	LUT3 #(
		.INIT('hb2)
	) name2705 (
		_w2646_,
		_w2647_,
		_w2648_,
		_w2771_
	);
	LUT3 #(
		.INIT('he8)
	) name2706 (
		_w2601_,
		_w2617_,
		_w2637_,
		_w2772_
	);
	LUT4 #(
		.INIT('h8228)
	) name2707 (
		_w2762_,
		_w2770_,
		_w2771_,
		_w2772_,
		_w2773_
	);
	LUT4 #(
		.INIT('h1441)
	) name2708 (
		_w2762_,
		_w2770_,
		_w2771_,
		_w2772_,
		_w2774_
	);
	LUT4 #(
		.INIT('h6996)
	) name2709 (
		_w2762_,
		_w2770_,
		_w2771_,
		_w2772_,
		_w2775_
	);
	LUT3 #(
		.INIT('h23)
	) name2710 (
		_w2659_,
		_w2660_,
		_w2662_,
		_w2776_
	);
	LUT3 #(
		.INIT('h4d)
	) name2711 (
		_w2668_,
		_w2669_,
		_w2676_,
		_w2777_
	);
	LUT3 #(
		.INIT('h2b)
	) name2712 (
		_w2654_,
		_w2655_,
		_w2656_,
		_w2778_
	);
	LUT3 #(
		.INIT('h2b)
	) name2713 (
		_w2665_,
		_w2666_,
		_w2667_,
		_w2779_
	);
	LUT3 #(
		.INIT('h0d)
	) name2714 (
		_w2591_,
		_w2592_,
		_w2593_,
		_w2780_
	);
	LUT3 #(
		.INIT('h0d)
	) name2715 (
		_w2527_,
		_w2602_,
		_w2604_,
		_w2781_
	);
	LUT3 #(
		.INIT('h0d)
	) name2716 (
		_w2631_,
		_w2632_,
		_w2634_,
		_w2782_
	);
	LUT3 #(
		.INIT('h96)
	) name2717 (
		_w2780_,
		_w2781_,
		_w2782_,
		_w2783_
	);
	LUT3 #(
		.INIT('h69)
	) name2718 (
		_w2778_,
		_w2779_,
		_w2783_,
		_w2784_
	);
	LUT3 #(
		.INIT('h69)
	) name2719 (
		_w2776_,
		_w2777_,
		_w2784_,
		_w2785_
	);
	LUT3 #(
		.INIT('hed)
	) name2720 (
		_w2752_,
		_w2775_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h10e0)
	) name2721 (
		_w2640_,
		_w2751_,
		_w2775_,
		_w2785_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2722 (
		_w2786_,
		_w2787_,
		_w2788_
	);
	LUT4 #(
		.INIT('h0bf4)
	) name2723 (
		_w2696_,
		_w2748_,
		_w2750_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h4)
	) name2724 (
		_w2695_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h9)
	) name2725 (
		_w2695_,
		_w2789_,
		_w2791_
	);
	LUT4 #(
		.INIT('he00e)
	) name2726 (
		_w2685_,
		_w2686_,
		_w2695_,
		_w2789_,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name2727 (
		_w2694_,
		_w2792_,
		_w2793_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2728 (
		_w2402_,
		_w2496_,
		_w2693_,
		_w2793_,
		_w2794_
	);
	LUT4 #(
		.INIT('hfdd0)
	) name2729 (
		_w2497_,
		_w2583_,
		_w2685_,
		_w2686_,
		_w2795_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2730 (
		_w2402_,
		_w2496_,
		_w2693_,
		_w2795_,
		_w2796_
	);
	LUT3 #(
		.INIT('h32)
	) name2731 (
		_w2791_,
		_w2794_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('hee0e)
	) name2732 (
		_w2685_,
		_w2686_,
		_w2695_,
		_w2789_,
		_w2798_
	);
	LUT2 #(
		.INIT('h4)
	) name2733 (
		_w2694_,
		_w2798_,
		_w2799_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2734 (
		_w2402_,
		_w2496_,
		_w2693_,
		_w2799_,
		_w2800_
	);
	LUT3 #(
		.INIT('h54)
	) name2735 (
		_w2749_,
		_w2750_,
		_w2788_,
		_w2801_
	);
	LUT4 #(
		.INIT('h1441)
	) name2736 (
		_w2640_,
		_w2776_,
		_w2777_,
		_w2784_,
		_w2802_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w2751_,
		_w2802_,
		_w2803_
	);
	LUT3 #(
		.INIT('h23)
	) name2738 (
		_w2751_,
		_w2773_,
		_w2802_,
		_w2804_
	);
	LUT4 #(
		.INIT('h1441)
	) name2739 (
		_w2774_,
		_w2776_,
		_w2777_,
		_w2784_,
		_w2805_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2740 (
		_w2588_,
		_w2589_,
		_w2638_,
		_w2774_,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w2805_,
		_w2806_,
		_w2807_
	);
	LUT3 #(
		.INIT('h17)
	) name2742 (
		_w2763_,
		_w2764_,
		_w2765_,
		_w2808_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		\a[0] ,
		\a[51] ,
		_w2809_
	);
	LUT3 #(
		.INIT('h80)
	) name2744 (
		\a[1] ,
		\a[26] ,
		\a[50] ,
		_w2810_
	);
	LUT3 #(
		.INIT('h6c)
	) name2745 (
		\a[1] ,
		\a[26] ,
		\a[50] ,
		_w2811_
	);
	LUT3 #(
		.INIT('h96)
	) name2746 (
		_w2755_,
		_w2809_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h8)
	) name2747 (
		\a[17] ,
		\a[34] ,
		_w2813_
	);
	LUT4 #(
		.INIT('h153f)
	) name2748 (
		\a[19] ,
		\a[20] ,
		\a[31] ,
		\a[32] ,
		_w2814_
	);
	LUT4 #(
		.INIT('h8000)
	) name2749 (
		\a[19] ,
		\a[20] ,
		\a[31] ,
		\a[32] ,
		_w2815_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2750 (
		\a[19] ,
		\a[20] ,
		\a[31] ,
		\a[32] ,
		_w2816_
	);
	LUT2 #(
		.INIT('h6)
	) name2751 (
		_w2813_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h8)
	) name2752 (
		_w2812_,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		_w2812_,
		_w2817_,
		_w2819_
	);
	LUT2 #(
		.INIT('h6)
	) name2754 (
		_w2812_,
		_w2817_,
		_w2820_
	);
	LUT4 #(
		.INIT('h153f)
	) name2755 (
		\a[22] ,
		\a[23] ,
		\a[28] ,
		\a[29] ,
		_w2821_
	);
	LUT4 #(
		.INIT('h8000)
	) name2756 (
		\a[22] ,
		\a[23] ,
		\a[28] ,
		\a[29] ,
		_w2822_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2757 (
		\a[22] ,
		\a[23] ,
		\a[28] ,
		\a[29] ,
		_w2823_
	);
	LUT2 #(
		.INIT('h8)
	) name2758 (
		\a[18] ,
		\a[33] ,
		_w2824_
	);
	LUT4 #(
		.INIT('h153f)
	) name2759 (
		\a[5] ,
		\a[16] ,
		\a[35] ,
		\a[46] ,
		_w2825_
	);
	LUT4 #(
		.INIT('h8000)
	) name2760 (
		\a[5] ,
		\a[16] ,
		\a[35] ,
		\a[46] ,
		_w2826_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2761 (
		\a[5] ,
		\a[16] ,
		\a[35] ,
		\a[46] ,
		_w2827_
	);
	LUT4 #(
		.INIT('h0660)
	) name2762 (
		_w2720_,
		_w2823_,
		_w2824_,
		_w2827_,
		_w2828_
	);
	LUT4 #(
		.INIT('h9009)
	) name2763 (
		_w2720_,
		_w2823_,
		_w2824_,
		_w2827_,
		_w2829_
	);
	LUT4 #(
		.INIT('h6996)
	) name2764 (
		_w2720_,
		_w2823_,
		_w2824_,
		_w2827_,
		_w2830_
	);
	LUT2 #(
		.INIT('h8)
	) name2765 (
		\a[15] ,
		\a[36] ,
		_w2831_
	);
	LUT4 #(
		.INIT('h153f)
	) name2766 (
		\a[6] ,
		\a[14] ,
		\a[37] ,
		\a[45] ,
		_w2832_
	);
	LUT4 #(
		.INIT('h8000)
	) name2767 (
		\a[6] ,
		\a[14] ,
		\a[37] ,
		\a[45] ,
		_w2833_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2768 (
		\a[6] ,
		\a[14] ,
		\a[37] ,
		\a[45] ,
		_w2834_
	);
	LUT2 #(
		.INIT('h6)
	) name2769 (
		_w2831_,
		_w2834_,
		_w2835_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		\a[7] ,
		\a[44] ,
		_w2836_
	);
	LUT4 #(
		.INIT('h153f)
	) name2771 (
		\a[8] ,
		\a[13] ,
		\a[38] ,
		\a[43] ,
		_w2837_
	);
	LUT4 #(
		.INIT('h8000)
	) name2772 (
		\a[8] ,
		\a[13] ,
		\a[38] ,
		\a[43] ,
		_w2838_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2773 (
		\a[8] ,
		\a[13] ,
		\a[38] ,
		\a[43] ,
		_w2839_
	);
	LUT2 #(
		.INIT('h8)
	) name2774 (
		\a[9] ,
		\a[42] ,
		_w2840_
	);
	LUT4 #(
		.INIT('h153f)
	) name2775 (
		\a[10] ,
		\a[12] ,
		\a[39] ,
		\a[41] ,
		_w2841_
	);
	LUT4 #(
		.INIT('h8000)
	) name2776 (
		\a[10] ,
		\a[12] ,
		\a[39] ,
		\a[41] ,
		_w2842_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2777 (
		\a[10] ,
		\a[12] ,
		\a[39] ,
		\a[41] ,
		_w2843_
	);
	LUT4 #(
		.INIT('h0660)
	) name2778 (
		_w2836_,
		_w2839_,
		_w2840_,
		_w2843_,
		_w2844_
	);
	LUT4 #(
		.INIT('h9009)
	) name2779 (
		_w2836_,
		_w2839_,
		_w2840_,
		_w2843_,
		_w2845_
	);
	LUT4 #(
		.INIT('h6996)
	) name2780 (
		_w2836_,
		_w2839_,
		_w2840_,
		_w2843_,
		_w2846_
	);
	LUT4 #(
		.INIT('h153f)
	) name2781 (
		\a[24] ,
		\a[25] ,
		\a[26] ,
		\a[27] ,
		_w2847_
	);
	LUT4 #(
		.INIT('h8000)
	) name2782 (
		\a[24] ,
		\a[25] ,
		\a[26] ,
		\a[27] ,
		_w2848_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2783 (
		\a[24] ,
		\a[25] ,
		\a[26] ,
		\a[27] ,
		_w2849_
	);
	LUT2 #(
		.INIT('h6)
	) name2784 (
		_w2737_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h0660)
	) name2785 (
		_w2830_,
		_w2835_,
		_w2846_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('h9009)
	) name2786 (
		_w2830_,
		_w2835_,
		_w2846_,
		_w2850_,
		_w2852_
	);
	LUT4 #(
		.INIT('h6996)
	) name2787 (
		_w2830_,
		_w2835_,
		_w2846_,
		_w2850_,
		_w2853_
	);
	LUT3 #(
		.INIT('h96)
	) name2788 (
		_w2808_,
		_w2820_,
		_w2853_,
		_w2854_
	);
	LUT4 #(
		.INIT('hd400)
	) name2789 (
		_w2776_,
		_w2777_,
		_w2784_,
		_w2854_,
		_w2855_
	);
	LUT4 #(
		.INIT('hbe28)
	) name2790 (
		_w2762_,
		_w2770_,
		_w2771_,
		_w2772_,
		_w2856_
	);
	LUT4 #(
		.INIT('h002b)
	) name2791 (
		_w2776_,
		_w2777_,
		_w2784_,
		_w2854_,
		_w2857_
	);
	LUT3 #(
		.INIT('hc9)
	) name2792 (
		_w2855_,
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT4 #(
		.INIT('hae00)
	) name2793 (
		_w2803_,
		_w2804_,
		_w2807_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h0051)
	) name2794 (
		_w2803_,
		_w2804_,
		_w2807_,
		_w2858_,
		_w2860_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2795 (
		_w2773_,
		_w2803_,
		_w2807_,
		_w2858_,
		_w2861_
	);
	LUT4 #(
		.INIT('h0017)
	) name2796 (
		_w2663_,
		_w2664_,
		_w2677_,
		_w2745_,
		_w2862_
	);
	LUT3 #(
		.INIT('h0e)
	) name2797 (
		_w2708_,
		_w2741_,
		_w2742_,
		_w2863_
	);
	LUT4 #(
		.INIT('h00ba)
	) name2798 (
		_w2672_,
		_w2673_,
		_w2675_,
		_w2705_,
		_w2864_
	);
	LUT3 #(
		.INIT('h0d)
	) name2799 (
		_w2735_,
		_w2736_,
		_w2738_,
		_w2865_
	);
	LUT3 #(
		.INIT('h0d)
	) name2800 (
		_w2697_,
		_w2698_,
		_w2699_,
		_w2866_
	);
	LUT2 #(
		.INIT('h8)
	) name2801 (
		\a[2] ,
		\a[49] ,
		_w2867_
	);
	LUT4 #(
		.INIT('h153f)
	) name2802 (
		\a[3] ,
		\a[4] ,
		\a[47] ,
		\a[48] ,
		_w2868_
	);
	LUT4 #(
		.INIT('h8000)
	) name2803 (
		\a[3] ,
		\a[4] ,
		\a[47] ,
		\a[48] ,
		_w2869_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2804 (
		\a[3] ,
		\a[4] ,
		\a[47] ,
		\a[48] ,
		_w2870_
	);
	LUT2 #(
		.INIT('h6)
	) name2805 (
		_w2867_,
		_w2870_,
		_w2871_
	);
	LUT3 #(
		.INIT('h69)
	) name2806 (
		_w2865_,
		_w2866_,
		_w2871_,
		_w2872_
	);
	LUT3 #(
		.INIT('he0)
	) name2807 (
		_w2706_,
		_w2864_,
		_w2872_,
		_w2873_
	);
	LUT3 #(
		.INIT('h01)
	) name2808 (
		_w2706_,
		_w2864_,
		_w2872_,
		_w2874_
	);
	LUT3 #(
		.INIT('h1e)
	) name2809 (
		_w2706_,
		_w2864_,
		_w2872_,
		_w2875_
	);
	LUT3 #(
		.INIT('h8e)
	) name2810 (
		_w2778_,
		_w2779_,
		_w2783_,
		_w2876_
	);
	LUT3 #(
		.INIT('h32)
	) name2811 (
		_w2728_,
		_w2729_,
		_w2730_,
		_w2877_
	);
	LUT3 #(
		.INIT('h0d)
	) name2812 (
		_w2620_,
		_w2724_,
		_w2726_,
		_w2878_
	);
	LUT3 #(
		.INIT('h32)
	) name2813 (
		_w2701_,
		_w2702_,
		_w2703_,
		_w2879_
	);
	LUT3 #(
		.INIT('h69)
	) name2814 (
		_w2877_,
		_w2878_,
		_w2879_,
		_w2880_
	);
	LUT3 #(
		.INIT('h32)
	) name2815 (
		_w2732_,
		_w2733_,
		_w2740_,
		_w2881_
	);
	LUT3 #(
		.INIT('h0d)
	) name2816 (
		_w2603_,
		_w2709_,
		_w2710_,
		_w2882_
	);
	LUT3 #(
		.INIT('h0d)
	) name2817 (
		_w2718_,
		_w2719_,
		_w2721_,
		_w2883_
	);
	LUT3 #(
		.INIT('h32)
	) name2818 (
		_w2670_,
		_w2712_,
		_w2713_,
		_w2884_
	);
	LUT3 #(
		.INIT('h96)
	) name2819 (
		_w2882_,
		_w2883_,
		_w2884_,
		_w2885_
	);
	LUT3 #(
		.INIT('h96)
	) name2820 (
		_w2880_,
		_w2881_,
		_w2885_,
		_w2886_
	);
	LUT4 #(
		.INIT('h6996)
	) name2821 (
		_w2863_,
		_w2875_,
		_w2876_,
		_w2886_,
		_w2887_
	);
	LUT3 #(
		.INIT('h23)
	) name2822 (
		_w2768_,
		_w2769_,
		_w2771_,
		_w2888_
	);
	LUT3 #(
		.INIT('h8e)
	) name2823 (
		_w2753_,
		_w2754_,
		_w2761_,
		_w2889_
	);
	LUT3 #(
		.INIT('h17)
	) name2824 (
		_w2780_,
		_w2781_,
		_w2782_,
		_w2890_
	);
	LUT3 #(
		.INIT('h45)
	) name2825 (
		_w2757_,
		_w2758_,
		_w2760_,
		_w2891_
	);
	LUT3 #(
		.INIT('h32)
	) name2826 (
		_w2715_,
		_w2716_,
		_w2723_,
		_w2892_
	);
	LUT3 #(
		.INIT('h96)
	) name2827 (
		_w2890_,
		_w2891_,
		_w2892_,
		_w2893_
	);
	LUT3 #(
		.INIT('h69)
	) name2828 (
		_w2888_,
		_w2889_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('he11e)
	) name2829 (
		_w2746_,
		_w2862_,
		_w2887_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h9)
	) name2830 (
		_w2861_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h4)
	) name2831 (
		_w2801_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name2832 (
		_w2801_,
		_w2896_,
		_w2898_
	);
	LUT2 #(
		.INIT('h9)
	) name2833 (
		_w2801_,
		_w2896_,
		_w2899_
	);
	LUT3 #(
		.INIT('h1e)
	) name2834 (
		_w2790_,
		_w2800_,
		_w2899_,
		_w2900_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2835 (
		_w2695_,
		_w2789_,
		_w2801_,
		_w2896_,
		_w2901_
	);
	LUT3 #(
		.INIT('h23)
	) name2836 (
		_w2859_,
		_w2860_,
		_w2895_,
		_w2902_
	);
	LUT4 #(
		.INIT('hbe28)
	) name2837 (
		_w2863_,
		_w2875_,
		_w2876_,
		_w2886_,
		_w2903_
	);
	LUT2 #(
		.INIT('h8)
	) name2838 (
		\a[10] ,
		\a[42] ,
		_w2904_
	);
	LUT4 #(
		.INIT('h153f)
	) name2839 (
		\a[11] ,
		\a[12] ,
		\a[40] ,
		\a[41] ,
		_w2905_
	);
	LUT4 #(
		.INIT('h8000)
	) name2840 (
		\a[11] ,
		\a[12] ,
		\a[40] ,
		\a[41] ,
		_w2906_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2841 (
		\a[11] ,
		\a[12] ,
		\a[40] ,
		\a[41] ,
		_w2907_
	);
	LUT2 #(
		.INIT('h8)
	) name2842 (
		\a[5] ,
		\a[47] ,
		_w2908_
	);
	LUT4 #(
		.INIT('h153f)
	) name2843 (
		\a[6] ,
		\a[16] ,
		\a[36] ,
		\a[46] ,
		_w2909_
	);
	LUT2 #(
		.INIT('h8)
	) name2844 (
		\a[16] ,
		\a[46] ,
		_w2910_
	);
	LUT4 #(
		.INIT('h8000)
	) name2845 (
		\a[6] ,
		\a[16] ,
		\a[36] ,
		\a[46] ,
		_w2911_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2846 (
		\a[6] ,
		\a[16] ,
		\a[36] ,
		\a[46] ,
		_w2912_
	);
	LUT4 #(
		.INIT('h0660)
	) name2847 (
		_w2904_,
		_w2907_,
		_w2908_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('h9009)
	) name2848 (
		_w2904_,
		_w2907_,
		_w2908_,
		_w2912_,
		_w2914_
	);
	LUT4 #(
		.INIT('h6996)
	) name2849 (
		_w2904_,
		_w2907_,
		_w2908_,
		_w2912_,
		_w2915_
	);
	LUT2 #(
		.INIT('h8)
	) name2850 (
		\a[15] ,
		\a[37] ,
		_w2916_
	);
	LUT4 #(
		.INIT('h153f)
	) name2851 (
		\a[7] ,
		\a[8] ,
		\a[44] ,
		\a[45] ,
		_w2917_
	);
	LUT2 #(
		.INIT('h8)
	) name2852 (
		\a[8] ,
		\a[45] ,
		_w2918_
	);
	LUT4 #(
		.INIT('h8000)
	) name2853 (
		\a[7] ,
		\a[8] ,
		\a[44] ,
		\a[45] ,
		_w2919_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2854 (
		\a[7] ,
		\a[8] ,
		\a[44] ,
		\a[45] ,
		_w2920_
	);
	LUT2 #(
		.INIT('h6)
	) name2855 (
		_w2916_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name2856 (
		\a[18] ,
		\a[34] ,
		_w2922_
	);
	LUT4 #(
		.INIT('h153f)
	) name2857 (
		\a[20] ,
		\a[21] ,
		\a[31] ,
		\a[32] ,
		_w2923_
	);
	LUT4 #(
		.INIT('h8000)
	) name2858 (
		\a[20] ,
		\a[21] ,
		\a[31] ,
		\a[32] ,
		_w2924_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2859 (
		\a[20] ,
		\a[21] ,
		\a[31] ,
		\a[32] ,
		_w2925_
	);
	LUT2 #(
		.INIT('h8)
	) name2860 (
		\a[22] ,
		\a[30] ,
		_w2926_
	);
	LUT4 #(
		.INIT('h153f)
	) name2861 (
		\a[23] ,
		\a[24] ,
		\a[28] ,
		\a[29] ,
		_w2927_
	);
	LUT4 #(
		.INIT('h8000)
	) name2862 (
		\a[23] ,
		\a[24] ,
		\a[28] ,
		\a[29] ,
		_w2928_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2863 (
		\a[23] ,
		\a[24] ,
		\a[28] ,
		\a[29] ,
		_w2929_
	);
	LUT4 #(
		.INIT('h0660)
	) name2864 (
		_w2922_,
		_w2925_,
		_w2926_,
		_w2929_,
		_w2930_
	);
	LUT4 #(
		.INIT('h9009)
	) name2865 (
		_w2922_,
		_w2925_,
		_w2926_,
		_w2929_,
		_w2931_
	);
	LUT4 #(
		.INIT('h6996)
	) name2866 (
		_w2922_,
		_w2925_,
		_w2926_,
		_w2929_,
		_w2932_
	);
	LUT4 #(
		.INIT('h153f)
	) name2867 (
		\a[9] ,
		\a[13] ,
		\a[39] ,
		\a[43] ,
		_w2933_
	);
	LUT4 #(
		.INIT('h8000)
	) name2868 (
		\a[9] ,
		\a[13] ,
		\a[39] ,
		\a[43] ,
		_w2934_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2869 (
		\a[9] ,
		\a[13] ,
		\a[39] ,
		\a[43] ,
		_w2935_
	);
	LUT2 #(
		.INIT('h6)
	) name2870 (
		_w1972_,
		_w2935_,
		_w2936_
	);
	LUT4 #(
		.INIT('h0660)
	) name2871 (
		_w2915_,
		_w2921_,
		_w2932_,
		_w2936_,
		_w2937_
	);
	LUT4 #(
		.INIT('h6996)
	) name2872 (
		_w2915_,
		_w2921_,
		_w2932_,
		_w2936_,
		_w2938_
	);
	LUT4 #(
		.INIT('he800)
	) name2873 (
		_w2880_,
		_w2881_,
		_w2885_,
		_w2938_,
		_w2939_
	);
	LUT4 #(
		.INIT('h17e8)
	) name2874 (
		_w2880_,
		_w2881_,
		_w2885_,
		_w2938_,
		_w2940_
	);
	LUT4 #(
		.INIT('hd400)
	) name2875 (
		_w2888_,
		_w2889_,
		_w2893_,
		_w2940_,
		_w2941_
	);
	LUT4 #(
		.INIT('h002b)
	) name2876 (
		_w2888_,
		_w2889_,
		_w2893_,
		_w2940_,
		_w2942_
	);
	LUT3 #(
		.INIT('ha9)
	) name2877 (
		_w2903_,
		_w2941_,
		_w2942_,
		_w2943_
	);
	LUT4 #(
		.INIT('hf110)
	) name2878 (
		_w2746_,
		_w2862_,
		_w2887_,
		_w2894_,
		_w2944_
	);
	LUT2 #(
		.INIT('h8)
	) name2879 (
		_w2943_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h1)
	) name2880 (
		_w2943_,
		_w2944_,
		_w2946_
	);
	LUT2 #(
		.INIT('h6)
	) name2881 (
		_w2943_,
		_w2944_,
		_w2947_
	);
	LUT3 #(
		.INIT('h23)
	) name2882 (
		_w2873_,
		_w2874_,
		_w2876_,
		_w2948_
	);
	LUT3 #(
		.INIT('hb2)
	) name2883 (
		_w2877_,
		_w2878_,
		_w2879_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name2884 (
		\a[19] ,
		\a[33] ,
		_w2950_
	);
	LUT4 #(
		.INIT('h153f)
	) name2885 (
		\a[2] ,
		\a[3] ,
		\a[49] ,
		\a[50] ,
		_w2951_
	);
	LUT4 #(
		.INIT('h8000)
	) name2886 (
		\a[2] ,
		\a[3] ,
		\a[49] ,
		\a[50] ,
		_w2952_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2887 (
		\a[2] ,
		\a[3] ,
		\a[49] ,
		\a[50] ,
		_w2953_
	);
	LUT2 #(
		.INIT('h6)
	) name2888 (
		_w2950_,
		_w2953_,
		_w2954_
	);
	LUT4 #(
		.INIT('h7100)
	) name2889 (
		_w2882_,
		_w2883_,
		_w2884_,
		_w2954_,
		_w2955_
	);
	LUT4 #(
		.INIT('h008e)
	) name2890 (
		_w2882_,
		_w2883_,
		_w2884_,
		_w2954_,
		_w2956_
	);
	LUT3 #(
		.INIT('ha9)
	) name2891 (
		_w2949_,
		_w2955_,
		_w2956_,
		_w2957_
	);
	LUT3 #(
		.INIT('h32)
	) name2892 (
		_w2844_,
		_w2845_,
		_w2850_,
		_w2958_
	);
	LUT4 #(
		.INIT('h8000)
	) name2893 (
		\a[1] ,
		\a[25] ,
		\a[27] ,
		\a[51] ,
		_w2959_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2894 (
		\a[1] ,
		\a[25] ,
		\a[27] ,
		\a[51] ,
		_w2960_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		_w2810_,
		_w2960_,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name2896 (
		_w2810_,
		_w2960_,
		_w2962_
	);
	LUT2 #(
		.INIT('h6)
	) name2897 (
		_w2810_,
		_w2960_,
		_w2963_
	);
	LUT3 #(
		.INIT('h0d)
	) name2898 (
		_w2737_,
		_w2847_,
		_w2848_,
		_w2964_
	);
	LUT2 #(
		.INIT('h6)
	) name2899 (
		_w2963_,
		_w2964_,
		_w2965_
	);
	LUT3 #(
		.INIT('h8e)
	) name2900 (
		_w2865_,
		_w2866_,
		_w2871_,
		_w2966_
	);
	LUT3 #(
		.INIT('h96)
	) name2901 (
		_w2958_,
		_w2965_,
		_w2966_,
		_w2967_
	);
	LUT3 #(
		.INIT('h69)
	) name2902 (
		_w2948_,
		_w2957_,
		_w2967_,
		_w2968_
	);
	LUT4 #(
		.INIT('h0051)
	) name2903 (
		_w2855_,
		_w2856_,
		_w2857_,
		_w2968_,
		_w2969_
	);
	LUT3 #(
		.INIT('h0e)
	) name2904 (
		_w2808_,
		_w2818_,
		_w2819_,
		_w2970_
	);
	LUT3 #(
		.INIT('he8)
	) name2905 (
		_w2755_,
		_w2809_,
		_w2811_,
		_w2971_
	);
	LUT3 #(
		.INIT('h0d)
	) name2906 (
		_w2840_,
		_w2841_,
		_w2842_,
		_w2972_
	);
	LUT4 #(
		.INIT('h153f)
	) name2907 (
		\a[4] ,
		\a[17] ,
		\a[35] ,
		\a[48] ,
		_w2973_
	);
	LUT4 #(
		.INIT('h8000)
	) name2908 (
		\a[4] ,
		\a[17] ,
		\a[35] ,
		\a[48] ,
		_w2974_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2909 (
		\a[4] ,
		\a[17] ,
		\a[35] ,
		\a[48] ,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		\a[0] ,
		\a[52] ,
		_w2976_
	);
	LUT2 #(
		.INIT('h6)
	) name2911 (
		_w2975_,
		_w2976_,
		_w2977_
	);
	LUT3 #(
		.INIT('h96)
	) name2912 (
		_w2971_,
		_w2972_,
		_w2977_,
		_w2978_
	);
	LUT4 #(
		.INIT('h1700)
	) name2913 (
		_w2808_,
		_w2812_,
		_w2817_,
		_w2978_,
		_w2979_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2914 (
		_w2808_,
		_w2812_,
		_w2817_,
		_w2978_,
		_w2980_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name2915 (
		_w2808_,
		_w2818_,
		_w2819_,
		_w2978_,
		_w2981_
	);
	LUT3 #(
		.INIT('he8)
	) name2916 (
		_w2890_,
		_w2891_,
		_w2892_,
		_w2982_
	);
	LUT4 #(
		.INIT('h00f6)
	) name2917 (
		_w2808_,
		_w2820_,
		_w2851_,
		_w2852_,
		_w2983_
	);
	LUT3 #(
		.INIT('h32)
	) name2918 (
		_w2824_,
		_w2825_,
		_w2826_,
		_w2984_
	);
	LUT3 #(
		.INIT('h0d)
	) name2919 (
		_w2836_,
		_w2837_,
		_w2838_,
		_w2985_
	);
	LUT3 #(
		.INIT('h0d)
	) name2920 (
		_w2720_,
		_w2821_,
		_w2822_,
		_w2986_
	);
	LUT3 #(
		.INIT('h69)
	) name2921 (
		_w2984_,
		_w2985_,
		_w2986_,
		_w2987_
	);
	LUT3 #(
		.INIT('h0d)
	) name2922 (
		_w2813_,
		_w2814_,
		_w2815_,
		_w2988_
	);
	LUT3 #(
		.INIT('h0d)
	) name2923 (
		_w2867_,
		_w2868_,
		_w2869_,
		_w2989_
	);
	LUT3 #(
		.INIT('h0d)
	) name2924 (
		_w2831_,
		_w2832_,
		_w2833_,
		_w2990_
	);
	LUT3 #(
		.INIT('h96)
	) name2925 (
		_w2988_,
		_w2989_,
		_w2990_,
		_w2991_
	);
	LUT3 #(
		.INIT('h32)
	) name2926 (
		_w2828_,
		_w2829_,
		_w2835_,
		_w2992_
	);
	LUT3 #(
		.INIT('h96)
	) name2927 (
		_w2987_,
		_w2991_,
		_w2992_,
		_w2993_
	);
	LUT4 #(
		.INIT('h6996)
	) name2928 (
		_w2981_,
		_w2982_,
		_w2983_,
		_w2993_,
		_w2994_
	);
	LUT3 #(
		.INIT('h51)
	) name2929 (
		_w2855_,
		_w2856_,
		_w2857_,
		_w2995_
	);
	LUT4 #(
		.INIT('hae00)
	) name2930 (
		_w2855_,
		_w2856_,
		_w2857_,
		_w2968_,
		_w2996_
	);
	LUT4 #(
		.INIT('hcae5)
	) name2931 (
		_w2968_,
		_w2969_,
		_w2994_,
		_w2995_,
		_w2997_
	);
	LUT2 #(
		.INIT('h6)
	) name2932 (
		_w2947_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h6)
	) name2933 (
		_w2902_,
		_w2998_,
		_w2999_
	);
	LUT4 #(
		.INIT('hdc23)
	) name2934 (
		_w2800_,
		_w2898_,
		_w2901_,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('h0e)
	) name2935 (
		_w2994_,
		_w2996_,
		_w2969_,
		_w3001_
	);
	LUT4 #(
		.INIT('hf660)
	) name2936 (
		_w2981_,
		_w2982_,
		_w2983_,
		_w2993_,
		_w3002_
	);
	LUT3 #(
		.INIT('h0e)
	) name2937 (
		_w2949_,
		_w2955_,
		_w2956_,
		_w3003_
	);
	LUT4 #(
		.INIT('h153f)
	) name2938 (
		\a[2] ,
		\a[3] ,
		\a[50] ,
		\a[51] ,
		_w3004_
	);
	LUT4 #(
		.INIT('h8000)
	) name2939 (
		\a[2] ,
		\a[3] ,
		\a[50] ,
		\a[51] ,
		_w3005_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2940 (
		\a[2] ,
		\a[3] ,
		\a[50] ,
		\a[51] ,
		_w3006_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		\a[4] ,
		\a[49] ,
		_w3007_
	);
	LUT4 #(
		.INIT('h153f)
	) name2942 (
		\a[17] ,
		\a[18] ,
		\a[35] ,
		\a[36] ,
		_w3008_
	);
	LUT4 #(
		.INIT('h8000)
	) name2943 (
		\a[17] ,
		\a[18] ,
		\a[35] ,
		\a[36] ,
		_w3009_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2944 (
		\a[17] ,
		\a[18] ,
		\a[35] ,
		\a[36] ,
		_w3010_
	);
	LUT4 #(
		.INIT('h0660)
	) name2945 (
		_w2959_,
		_w3006_,
		_w3007_,
		_w3010_,
		_w3011_
	);
	LUT4 #(
		.INIT('h9009)
	) name2946 (
		_w2959_,
		_w3006_,
		_w3007_,
		_w3010_,
		_w3012_
	);
	LUT4 #(
		.INIT('h6996)
	) name2947 (
		_w2959_,
		_w3006_,
		_w3007_,
		_w3010_,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name2948 (
		\a[19] ,
		\a[34] ,
		_w3014_
	);
	LUT4 #(
		.INIT('h153f)
	) name2949 (
		\a[20] ,
		\a[21] ,
		\a[32] ,
		\a[33] ,
		_w3015_
	);
	LUT4 #(
		.INIT('h8000)
	) name2950 (
		\a[20] ,
		\a[21] ,
		\a[32] ,
		\a[33] ,
		_w3016_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2951 (
		\a[20] ,
		\a[21] ,
		\a[32] ,
		\a[33] ,
		_w3017_
	);
	LUT2 #(
		.INIT('h6)
	) name2952 (
		_w3014_,
		_w3017_,
		_w3018_
	);
	LUT2 #(
		.INIT('h6)
	) name2953 (
		_w3013_,
		_w3018_,
		_w3019_
	);
	LUT4 #(
		.INIT('h153f)
	) name2954 (
		\a[9] ,
		\a[14] ,
		\a[39] ,
		\a[44] ,
		_w3020_
	);
	LUT2 #(
		.INIT('h8)
	) name2955 (
		\a[14] ,
		\a[44] ,
		_w3021_
	);
	LUT4 #(
		.INIT('h8000)
	) name2956 (
		\a[9] ,
		\a[14] ,
		\a[39] ,
		\a[44] ,
		_w3022_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2957 (
		\a[9] ,
		\a[14] ,
		\a[39] ,
		\a[44] ,
		_w3023_
	);
	LUT2 #(
		.INIT('h8)
	) name2958 (
		\a[6] ,
		\a[47] ,
		_w3024_
	);
	LUT4 #(
		.INIT('h153f)
	) name2959 (
		\a[7] ,
		\a[15] ,
		\a[38] ,
		\a[46] ,
		_w3025_
	);
	LUT4 #(
		.INIT('h8000)
	) name2960 (
		\a[7] ,
		\a[15] ,
		\a[38] ,
		\a[46] ,
		_w3026_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2961 (
		\a[7] ,
		\a[15] ,
		\a[38] ,
		\a[46] ,
		_w3027_
	);
	LUT4 #(
		.INIT('h0660)
	) name2962 (
		_w2918_,
		_w3023_,
		_w3024_,
		_w3027_,
		_w3028_
	);
	LUT4 #(
		.INIT('h9009)
	) name2963 (
		_w2918_,
		_w3023_,
		_w3024_,
		_w3027_,
		_w3029_
	);
	LUT4 #(
		.INIT('h6996)
	) name2964 (
		_w2918_,
		_w3023_,
		_w3024_,
		_w3027_,
		_w3030_
	);
	LUT2 #(
		.INIT('h8)
	) name2965 (
		\a[0] ,
		\a[53] ,
		_w3031_
	);
	LUT4 #(
		.INIT('h153f)
	) name2966 (
		\a[5] ,
		\a[16] ,
		\a[37] ,
		\a[48] ,
		_w3032_
	);
	LUT4 #(
		.INIT('h8000)
	) name2967 (
		\a[5] ,
		\a[16] ,
		\a[37] ,
		\a[48] ,
		_w3033_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2968 (
		\a[5] ,
		\a[16] ,
		\a[37] ,
		\a[48] ,
		_w3034_
	);
	LUT2 #(
		.INIT('h6)
	) name2969 (
		_w3031_,
		_w3034_,
		_w3035_
	);
	LUT2 #(
		.INIT('h6)
	) name2970 (
		_w3030_,
		_w3035_,
		_w3036_
	);
	LUT4 #(
		.INIT('h9009)
	) name2971 (
		_w3013_,
		_w3018_,
		_w3030_,
		_w3035_,
		_w3037_
	);
	LUT3 #(
		.INIT('h96)
	) name2972 (
		_w3003_,
		_w3019_,
		_w3036_,
		_w3038_
	);
	LUT3 #(
		.INIT('h2b)
	) name2973 (
		_w2958_,
		_w2965_,
		_w2966_,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name2974 (
		\a[13] ,
		\a[40] ,
		_w3040_
	);
	LUT4 #(
		.INIT('h153f)
	) name2975 (
		\a[10] ,
		\a[12] ,
		\a[41] ,
		\a[43] ,
		_w3041_
	);
	LUT2 #(
		.INIT('h8)
	) name2976 (
		\a[12] ,
		\a[43] ,
		_w3042_
	);
	LUT4 #(
		.INIT('h8000)
	) name2977 (
		\a[10] ,
		\a[12] ,
		\a[41] ,
		\a[43] ,
		_w3043_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2978 (
		\a[10] ,
		\a[12] ,
		\a[41] ,
		\a[43] ,
		_w3044_
	);
	LUT2 #(
		.INIT('h8)
	) name2979 (
		\a[22] ,
		\a[31] ,
		_w3045_
	);
	LUT4 #(
		.INIT('h153f)
	) name2980 (
		\a[23] ,
		\a[24] ,
		\a[29] ,
		\a[30] ,
		_w3046_
	);
	LUT4 #(
		.INIT('h8000)
	) name2981 (
		\a[23] ,
		\a[24] ,
		\a[29] ,
		\a[30] ,
		_w3047_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2982 (
		\a[23] ,
		\a[24] ,
		\a[29] ,
		\a[30] ,
		_w3048_
	);
	LUT4 #(
		.INIT('h0660)
	) name2983 (
		_w3040_,
		_w3044_,
		_w3045_,
		_w3048_,
		_w3049_
	);
	LUT4 #(
		.INIT('h9009)
	) name2984 (
		_w3040_,
		_w3044_,
		_w3045_,
		_w3048_,
		_w3050_
	);
	LUT4 #(
		.INIT('h6996)
	) name2985 (
		_w3040_,
		_w3044_,
		_w3045_,
		_w3048_,
		_w3051_
	);
	LUT2 #(
		.INIT('h8)
	) name2986 (
		\a[11] ,
		\a[42] ,
		_w3052_
	);
	LUT4 #(
		.INIT('h153f)
	) name2987 (
		\a[25] ,
		\a[26] ,
		\a[27] ,
		\a[28] ,
		_w3053_
	);
	LUT4 #(
		.INIT('h8000)
	) name2988 (
		\a[25] ,
		\a[26] ,
		\a[27] ,
		\a[28] ,
		_w3054_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2989 (
		\a[25] ,
		\a[26] ,
		\a[27] ,
		\a[28] ,
		_w3055_
	);
	LUT2 #(
		.INIT('h6)
	) name2990 (
		_w3052_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h6)
	) name2991 (
		_w3051_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('h00d4)
	) name2992 (
		_w2958_,
		_w2965_,
		_w2966_,
		_w3057_,
		_w3058_
	);
	LUT4 #(
		.INIT('h2b00)
	) name2993 (
		_w2958_,
		_w2965_,
		_w2966_,
		_w3057_,
		_w3059_
	);
	LUT4 #(
		.INIT('hd42b)
	) name2994 (
		_w2958_,
		_w2965_,
		_w2966_,
		_w3057_,
		_w3060_
	);
	LUT3 #(
		.INIT('h71)
	) name2995 (
		_w2987_,
		_w2991_,
		_w2992_,
		_w3061_
	);
	LUT2 #(
		.INIT('h6)
	) name2996 (
		_w3060_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('h96)
	) name2997 (
		_w3002_,
		_w3038_,
		_w3062_,
		_w3063_
	);
	LUT4 #(
		.INIT('hf10e)
	) name2998 (
		_w2994_,
		_w2996_,
		_w2969_,
		_w3063_,
		_w3064_
	);
	LUT3 #(
		.INIT('h54)
	) name2999 (
		_w2973_,
		_w2974_,
		_w2976_,
		_w3065_
	);
	LUT3 #(
		.INIT('h0d)
	) name3000 (
		_w2950_,
		_w2951_,
		_w2952_,
		_w3066_
	);
	LUT3 #(
		.INIT('h0d)
	) name3001 (
		_w2926_,
		_w2927_,
		_w2928_,
		_w3067_
	);
	LUT3 #(
		.INIT('h69)
	) name3002 (
		_w3065_,
		_w3066_,
		_w3067_,
		_w3068_
	);
	LUT3 #(
		.INIT('h32)
	) name3003 (
		_w2930_,
		_w2931_,
		_w2936_,
		_w3069_
	);
	LUT3 #(
		.INIT('h4d)
	) name3004 (
		_w2971_,
		_w2972_,
		_w2977_,
		_w3070_
	);
	LUT3 #(
		.INIT('h96)
	) name3005 (
		_w3068_,
		_w3069_,
		_w3070_,
		_w3071_
	);
	LUT3 #(
		.INIT('h0d)
	) name3006 (
		_w2908_,
		_w2909_,
		_w2911_,
		_w3072_
	);
	LUT3 #(
		.INIT('h0d)
	) name3007 (
		_w2922_,
		_w2923_,
		_w2924_,
		_w3073_
	);
	LUT3 #(
		.INIT('h0d)
	) name3008 (
		_w2916_,
		_w2917_,
		_w2919_,
		_w3074_
	);
	LUT3 #(
		.INIT('h96)
	) name3009 (
		_w3072_,
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT3 #(
		.INIT('h32)
	) name3010 (
		_w2913_,
		_w2914_,
		_w2921_,
		_w3076_
	);
	LUT3 #(
		.INIT('h80)
	) name3011 (
		\a[1] ,
		\a[27] ,
		\a[52] ,
		_w3077_
	);
	LUT3 #(
		.INIT('h6c)
	) name3012 (
		\a[1] ,
		\a[27] ,
		\a[52] ,
		_w3078_
	);
	LUT4 #(
		.INIT('h000d)
	) name3013 (
		_w2904_,
		_w2905_,
		_w2906_,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('hf200)
	) name3014 (
		_w2904_,
		_w2905_,
		_w2906_,
		_w3078_,
		_w3080_
	);
	LUT4 #(
		.INIT('h0df2)
	) name3015 (
		_w2904_,
		_w2905_,
		_w2906_,
		_w3078_,
		_w3081_
	);
	LUT3 #(
		.INIT('h0d)
	) name3016 (
		_w1972_,
		_w2933_,
		_w2934_,
		_w3082_
	);
	LUT2 #(
		.INIT('h6)
	) name3017 (
		_w3081_,
		_w3082_,
		_w3083_
	);
	LUT3 #(
		.INIT('h96)
	) name3018 (
		_w3075_,
		_w3076_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h8)
	) name3019 (
		_w3071_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h1)
	) name3020 (
		_w3071_,
		_w3084_,
		_w3086_
	);
	LUT2 #(
		.INIT('h6)
	) name3021 (
		_w3071_,
		_w3084_,
		_w3087_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name3022 (
		_w2948_,
		_w2957_,
		_w2967_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h1)
	) name3023 (
		_w2937_,
		_w2939_,
		_w3089_
	);
	LUT3 #(
		.INIT('h2b)
	) name3024 (
		_w2984_,
		_w2985_,
		_w2986_,
		_w3090_
	);
	LUT3 #(
		.INIT('h23)
	) name3025 (
		_w2961_,
		_w2962_,
		_w2964_,
		_w3091_
	);
	LUT3 #(
		.INIT('h17)
	) name3026 (
		_w2988_,
		_w2989_,
		_w2990_,
		_w3092_
	);
	LUT3 #(
		.INIT('h96)
	) name3027 (
		_w3090_,
		_w3091_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h004d)
	) name3028 (
		_w2970_,
		_w2978_,
		_w2982_,
		_w3093_,
		_w3094_
	);
	LUT4 #(
		.INIT('hb200)
	) name3029 (
		_w2970_,
		_w2978_,
		_w2982_,
		_w3093_,
		_w3095_
	);
	LUT4 #(
		.INIT('hab54)
	) name3030 (
		_w2979_,
		_w2980_,
		_w2982_,
		_w3093_,
		_w3096_
	);
	LUT2 #(
		.INIT('h9)
	) name3031 (
		_w3089_,
		_w3096_,
		_w3097_
	);
	LUT4 #(
		.INIT('h0031)
	) name3032 (
		_w2903_,
		_w2941_,
		_w2942_,
		_w3097_,
		_w3098_
	);
	LUT4 #(
		.INIT('h31ff)
	) name3033 (
		_w2903_,
		_w2941_,
		_w2942_,
		_w3097_,
		_w3099_
	);
	LUT4 #(
		.INIT('h31ce)
	) name3034 (
		_w2903_,
		_w2941_,
		_w2942_,
		_w3097_,
		_w3100_
	);
	LUT2 #(
		.INIT('h6)
	) name3035 (
		_w3088_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name3036 (
		_w3064_,
		_w3101_,
		_w3102_
	);
	LUT3 #(
		.INIT('h32)
	) name3037 (
		_w2945_,
		_w2946_,
		_w2997_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name3038 (
		_w3064_,
		_w3101_,
		_w3104_
	);
	LUT3 #(
		.INIT('h04)
	) name3039 (
		_w3102_,
		_w3103_,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('h6)
	) name3040 (
		_w3064_,
		_w3101_,
		_w3106_
	);
	LUT3 #(
		.INIT('h96)
	) name3041 (
		_w3064_,
		_w3101_,
		_w3103_,
		_w3107_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3042 (
		_w2695_,
		_w2789_,
		_w2902_,
		_w2998_,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name3043 (
		_w2897_,
		_w3108_,
		_w3109_
	);
	LUT4 #(
		.INIT('h0222)
	) name3044 (
		_w2801_,
		_w2896_,
		_w2902_,
		_w2998_,
		_w3110_
	);
	LUT4 #(
		.INIT('hfdd0)
	) name3045 (
		_w2801_,
		_w2896_,
		_w2902_,
		_w2998_,
		_w3111_
	);
	LUT4 #(
		.INIT('h63cc)
	) name3046 (
		_w2800_,
		_w3107_,
		_w3109_,
		_w3111_,
		_w3112_
	);
	LUT3 #(
		.INIT('he8)
	) name3047 (
		_w3001_,
		_w3063_,
		_w3101_,
		_w3113_
	);
	LUT4 #(
		.INIT('h002b)
	) name3048 (
		_w2948_,
		_w2957_,
		_w2967_,
		_w3085_,
		_w3114_
	);
	LUT3 #(
		.INIT('h31)
	) name3049 (
		_w3089_,
		_w3094_,
		_w3095_,
		_w3115_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		\a[19] ,
		\a[35] ,
		_w3116_
	);
	LUT4 #(
		.INIT('h153f)
	) name3051 (
		\a[21] ,
		\a[22] ,
		\a[32] ,
		\a[33] ,
		_w3117_
	);
	LUT4 #(
		.INIT('h8000)
	) name3052 (
		\a[21] ,
		\a[22] ,
		\a[32] ,
		\a[33] ,
		_w3118_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3053 (
		\a[21] ,
		\a[22] ,
		\a[32] ,
		\a[33] ,
		_w3119_
	);
	LUT2 #(
		.INIT('h8)
	) name3054 (
		\a[23] ,
		\a[31] ,
		_w3120_
	);
	LUT4 #(
		.INIT('h153f)
	) name3055 (
		\a[24] ,
		\a[25] ,
		\a[29] ,
		\a[30] ,
		_w3121_
	);
	LUT4 #(
		.INIT('h8000)
	) name3056 (
		\a[24] ,
		\a[25] ,
		\a[29] ,
		\a[30] ,
		_w3122_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3057 (
		\a[24] ,
		\a[25] ,
		\a[29] ,
		\a[30] ,
		_w3123_
	);
	LUT4 #(
		.INIT('h0660)
	) name3058 (
		_w3116_,
		_w3119_,
		_w3120_,
		_w3123_,
		_w3124_
	);
	LUT4 #(
		.INIT('h9009)
	) name3059 (
		_w3116_,
		_w3119_,
		_w3120_,
		_w3123_,
		_w3125_
	);
	LUT4 #(
		.INIT('h6996)
	) name3060 (
		_w3116_,
		_w3119_,
		_w3120_,
		_w3123_,
		_w3126_
	);
	LUT4 #(
		.INIT('h8000)
	) name3061 (
		\a[1] ,
		\a[26] ,
		\a[28] ,
		\a[53] ,
		_w3127_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3062 (
		\a[1] ,
		\a[26] ,
		\a[28] ,
		\a[53] ,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name3063 (
		\a[0] ,
		\a[54] ,
		_w3129_
	);
	LUT3 #(
		.INIT('h96)
	) name3064 (
		_w3077_,
		_w3128_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h6)
	) name3065 (
		_w3126_,
		_w3130_,
		_w3131_
	);
	LUT4 #(
		.INIT('h00b2)
	) name3066 (
		_w3068_,
		_w3069_,
		_w3070_,
		_w3131_,
		_w3132_
	);
	LUT3 #(
		.INIT('h4d)
	) name3067 (
		_w3075_,
		_w3076_,
		_w3083_,
		_w3133_
	);
	LUT4 #(
		.INIT('h4d00)
	) name3068 (
		_w3068_,
		_w3069_,
		_w3070_,
		_w3131_,
		_w3134_
	);
	LUT3 #(
		.INIT('hc9)
	) name3069 (
		_w3132_,
		_w3133_,
		_w3134_,
		_w3135_
	);
	LUT4 #(
		.INIT('h1eff)
	) name3070 (
		_w3086_,
		_w3114_,
		_w3115_,
		_w3135_,
		_w3136_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name3071 (
		_w3086_,
		_w3114_,
		_w3115_,
		_w3135_,
		_w3137_
	);
	LUT4 #(
		.INIT('h2300)
	) name3072 (
		_w3088_,
		_w3098_,
		_w3099_,
		_w3137_,
		_w3138_
	);
	LUT4 #(
		.INIT('h00dc)
	) name3073 (
		_w3088_,
		_w3098_,
		_w3099_,
		_w3137_,
		_w3139_
	);
	LUT4 #(
		.INIT('hdc23)
	) name3074 (
		_w3088_,
		_w3098_,
		_w3099_,
		_w3137_,
		_w3140_
	);
	LUT3 #(
		.INIT('he8)
	) name3075 (
		_w3002_,
		_w3038_,
		_w3062_,
		_w3141_
	);
	LUT3 #(
		.INIT('h17)
	) name3076 (
		_w3072_,
		_w3073_,
		_w3074_,
		_w3142_
	);
	LUT3 #(
		.INIT('h2b)
	) name3077 (
		_w3065_,
		_w3066_,
		_w3067_,
		_w3143_
	);
	LUT3 #(
		.INIT('h45)
	) name3078 (
		_w3079_,
		_w3080_,
		_w3082_,
		_w3144_
	);
	LUT3 #(
		.INIT('h96)
	) name3079 (
		_w3142_,
		_w3143_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3080 (
		_w2949_,
		_w2955_,
		_w2956_,
		_w3019_,
		_w3146_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3081 (
		_w2949_,
		_w2955_,
		_w2956_,
		_w3036_,
		_w3147_
	);
	LUT3 #(
		.INIT('h01)
	) name3082 (
		_w3037_,
		_w3146_,
		_w3147_,
		_w3148_
	);
	LUT4 #(
		.INIT('h0017)
	) name3083 (
		_w3003_,
		_w3019_,
		_w3036_,
		_w3145_,
		_w3149_
	);
	LUT4 #(
		.INIT('he800)
	) name3084 (
		_w3003_,
		_w3019_,
		_w3036_,
		_w3145_,
		_w3150_
	);
	LUT3 #(
		.INIT('h32)
	) name3085 (
		_w3024_,
		_w3025_,
		_w3026_,
		_w3151_
	);
	LUT3 #(
		.INIT('h0d)
	) name3086 (
		_w3031_,
		_w3032_,
		_w3033_,
		_w3152_
	);
	LUT3 #(
		.INIT('h0d)
	) name3087 (
		_w3052_,
		_w3053_,
		_w3054_,
		_w3153_
	);
	LUT3 #(
		.INIT('h69)
	) name3088 (
		_w3151_,
		_w3152_,
		_w3153_,
		_w3154_
	);
	LUT3 #(
		.INIT('h0d)
	) name3089 (
		_w3007_,
		_w3008_,
		_w3009_,
		_w3155_
	);
	LUT3 #(
		.INIT('h0d)
	) name3090 (
		_w3014_,
		_w3015_,
		_w3016_,
		_w3156_
	);
	LUT3 #(
		.INIT('h0d)
	) name3091 (
		_w3045_,
		_w3046_,
		_w3047_,
		_w3157_
	);
	LUT3 #(
		.INIT('h96)
	) name3092 (
		_w3155_,
		_w3156_,
		_w3157_,
		_w3158_
	);
	LUT3 #(
		.INIT('h32)
	) name3093 (
		_w3028_,
		_w3029_,
		_w3035_,
		_w3159_
	);
	LUT3 #(
		.INIT('h96)
	) name3094 (
		_w3154_,
		_w3158_,
		_w3159_,
		_w3160_
	);
	LUT3 #(
		.INIT('h96)
	) name3095 (
		_w3145_,
		_w3148_,
		_w3160_,
		_w3161_
	);
	LUT3 #(
		.INIT('he8)
	) name3096 (
		_w3090_,
		_w3091_,
		_w3092_,
		_w3162_
	);
	LUT4 #(
		.INIT('h153f)
	) name3097 (
		\a[11] ,
		\a[12] ,
		\a[42] ,
		\a[43] ,
		_w3163_
	);
	LUT4 #(
		.INIT('h8000)
	) name3098 (
		\a[11] ,
		\a[12] ,
		\a[42] ,
		\a[43] ,
		_w3164_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3099 (
		\a[11] ,
		\a[12] ,
		\a[42] ,
		\a[43] ,
		_w3165_
	);
	LUT2 #(
		.INIT('h8)
	) name3100 (
		\a[20] ,
		\a[34] ,
		_w3166_
	);
	LUT4 #(
		.INIT('h153f)
	) name3101 (
		\a[5] ,
		\a[18] ,
		\a[36] ,
		\a[49] ,
		_w3167_
	);
	LUT4 #(
		.INIT('h8000)
	) name3102 (
		\a[5] ,
		\a[18] ,
		\a[36] ,
		\a[49] ,
		_w3168_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3103 (
		\a[5] ,
		\a[18] ,
		\a[36] ,
		\a[49] ,
		_w3169_
	);
	LUT4 #(
		.INIT('h0660)
	) name3104 (
		_w2725_,
		_w3165_,
		_w3166_,
		_w3169_,
		_w3170_
	);
	LUT4 #(
		.INIT('h9009)
	) name3105 (
		_w2725_,
		_w3165_,
		_w3166_,
		_w3169_,
		_w3171_
	);
	LUT4 #(
		.INIT('h6996)
	) name3106 (
		_w2725_,
		_w3165_,
		_w3166_,
		_w3169_,
		_w3172_
	);
	LUT2 #(
		.INIT('h8)
	) name3107 (
		\a[17] ,
		\a[37] ,
		_w3173_
	);
	LUT4 #(
		.INIT('h153f)
	) name3108 (
		\a[6] ,
		\a[16] ,
		\a[38] ,
		\a[48] ,
		_w3174_
	);
	LUT4 #(
		.INIT('h8000)
	) name3109 (
		\a[6] ,
		\a[16] ,
		\a[38] ,
		\a[48] ,
		_w3175_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3110 (
		\a[6] ,
		\a[16] ,
		\a[38] ,
		\a[48] ,
		_w3176_
	);
	LUT2 #(
		.INIT('h6)
	) name3111 (
		_w3173_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h6)
	) name3112 (
		_w3172_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h8)
	) name3113 (
		\a[2] ,
		\a[52] ,
		_w3179_
	);
	LUT4 #(
		.INIT('h153f)
	) name3114 (
		\a[3] ,
		\a[4] ,
		\a[50] ,
		\a[51] ,
		_w3180_
	);
	LUT4 #(
		.INIT('h8000)
	) name3115 (
		\a[3] ,
		\a[4] ,
		\a[50] ,
		\a[51] ,
		_w3181_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3116 (
		\a[3] ,
		\a[4] ,
		\a[50] ,
		\a[51] ,
		_w3182_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		\a[7] ,
		\a[47] ,
		_w3183_
	);
	LUT4 #(
		.INIT('h153f)
	) name3118 (
		\a[8] ,
		\a[15] ,
		\a[39] ,
		\a[46] ,
		_w3184_
	);
	LUT4 #(
		.INIT('h8000)
	) name3119 (
		\a[8] ,
		\a[15] ,
		\a[39] ,
		\a[46] ,
		_w3185_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3120 (
		\a[8] ,
		\a[15] ,
		\a[39] ,
		\a[46] ,
		_w3186_
	);
	LUT4 #(
		.INIT('h0660)
	) name3121 (
		_w3179_,
		_w3182_,
		_w3183_,
		_w3186_,
		_w3187_
	);
	LUT4 #(
		.INIT('h9009)
	) name3122 (
		_w3179_,
		_w3182_,
		_w3183_,
		_w3186_,
		_w3188_
	);
	LUT4 #(
		.INIT('h6996)
	) name3123 (
		_w3179_,
		_w3182_,
		_w3183_,
		_w3186_,
		_w3189_
	);
	LUT2 #(
		.INIT('h8)
	) name3124 (
		\a[9] ,
		\a[45] ,
		_w3190_
	);
	LUT4 #(
		.INIT('h153f)
	) name3125 (
		\a[10] ,
		\a[14] ,
		\a[40] ,
		\a[44] ,
		_w3191_
	);
	LUT4 #(
		.INIT('h8000)
	) name3126 (
		\a[10] ,
		\a[14] ,
		\a[40] ,
		\a[44] ,
		_w3192_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3127 (
		\a[10] ,
		\a[14] ,
		\a[40] ,
		\a[44] ,
		_w3193_
	);
	LUT2 #(
		.INIT('h6)
	) name3128 (
		_w3190_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h6)
	) name3129 (
		_w3189_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h0990)
	) name3130 (
		_w3172_,
		_w3177_,
		_w3189_,
		_w3194_,
		_w3196_
	);
	LUT4 #(
		.INIT('he800)
	) name3131 (
		_w3090_,
		_w3091_,
		_w3092_,
		_w3196_,
		_w3197_
	);
	LUT4 #(
		.INIT('h0660)
	) name3132 (
		_w3172_,
		_w3177_,
		_w3189_,
		_w3194_,
		_w3198_
	);
	LUT4 #(
		.INIT('h1700)
	) name3133 (
		_w3090_,
		_w3091_,
		_w3092_,
		_w3198_,
		_w3199_
	);
	LUT3 #(
		.INIT('h96)
	) name3134 (
		_w3162_,
		_w3178_,
		_w3195_,
		_w3200_
	);
	LUT3 #(
		.INIT('h0d)
	) name3135 (
		_w2918_,
		_w3020_,
		_w3022_,
		_w3201_
	);
	LUT3 #(
		.INIT('h0d)
	) name3136 (
		_w2959_,
		_w3004_,
		_w3005_,
		_w3202_
	);
	LUT3 #(
		.INIT('h0d)
	) name3137 (
		_w3040_,
		_w3041_,
		_w3043_,
		_w3203_
	);
	LUT3 #(
		.INIT('h96)
	) name3138 (
		_w3201_,
		_w3202_,
		_w3203_,
		_w3204_
	);
	LUT3 #(
		.INIT('h32)
	) name3139 (
		_w3049_,
		_w3050_,
		_w3056_,
		_w3205_
	);
	LUT3 #(
		.INIT('h32)
	) name3140 (
		_w3011_,
		_w3012_,
		_w3018_,
		_w3206_
	);
	LUT3 #(
		.INIT('h69)
	) name3141 (
		_w3204_,
		_w3205_,
		_w3206_,
		_w3207_
	);
	LUT4 #(
		.INIT('he800)
	) name3142 (
		_w3039_,
		_w3057_,
		_w3061_,
		_w3207_,
		_w3208_
	);
	LUT4 #(
		.INIT('h0017)
	) name3143 (
		_w3039_,
		_w3057_,
		_w3061_,
		_w3207_,
		_w3209_
	);
	LUT4 #(
		.INIT('hab54)
	) name3144 (
		_w3058_,
		_w3059_,
		_w3061_,
		_w3207_,
		_w3210_
	);
	LUT2 #(
		.INIT('h6)
	) name3145 (
		_w3200_,
		_w3210_,
		_w3211_
	);
	LUT3 #(
		.INIT('h96)
	) name3146 (
		_w3141_,
		_w3161_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h6)
	) name3147 (
		_w3140_,
		_w3212_,
		_w3213_
	);
	LUT2 #(
		.INIT('h8)
	) name3148 (
		_w3113_,
		_w3213_,
		_w3214_
	);
	LUT2 #(
		.INIT('h1)
	) name3149 (
		_w3113_,
		_w3213_,
		_w3215_
	);
	LUT2 #(
		.INIT('h6)
	) name3150 (
		_w3113_,
		_w3213_,
		_w3216_
	);
	LUT4 #(
		.INIT('heee0)
	) name3151 (
		_w2902_,
		_w2998_,
		_w3103_,
		_w3106_,
		_w3217_
	);
	LUT2 #(
		.INIT('h4)
	) name3152 (
		_w3110_,
		_w3217_,
		_w3218_
	);
	LUT3 #(
		.INIT('hb0)
	) name3153 (
		_w2800_,
		_w3109_,
		_w3218_,
		_w3219_
	);
	LUT3 #(
		.INIT('h36)
	) name3154 (
		_w3105_,
		_w3216_,
		_w3219_,
		_w3220_
	);
	LUT2 #(
		.INIT('h1)
	) name3155 (
		_w3105_,
		_w3214_,
		_w3221_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3156 (
		_w2800_,
		_w3109_,
		_w3218_,
		_w3221_,
		_w3222_
	);
	LUT3 #(
		.INIT('h32)
	) name3157 (
		_w3138_,
		_w3139_,
		_w3212_,
		_w3223_
	);
	LUT3 #(
		.INIT('h10)
	) name3158 (
		_w3086_,
		_w3114_,
		_w3115_,
		_w3224_
	);
	LUT4 #(
		.INIT('h0eef)
	) name3159 (
		_w3086_,
		_w3114_,
		_w3115_,
		_w3135_,
		_w3225_
	);
	LUT4 #(
		.INIT('he800)
	) name3160 (
		_w3090_,
		_w3091_,
		_w3092_,
		_w3178_,
		_w3226_
	);
	LUT3 #(
		.INIT('h17)
	) name3161 (
		_w3162_,
		_w3178_,
		_w3195_,
		_w3227_
	);
	LUT3 #(
		.INIT('h2b)
	) name3162 (
		_w3151_,
		_w3152_,
		_w3153_,
		_w3228_
	);
	LUT3 #(
		.INIT('h17)
	) name3163 (
		_w3201_,
		_w3202_,
		_w3203_,
		_w3229_
	);
	LUT2 #(
		.INIT('h4)
	) name3164 (
		\a[54] ,
		_w3127_,
		_w3230_
	);
	LUT2 #(
		.INIT('h8)
	) name3165 (
		\a[28] ,
		\a[54] ,
		_w3231_
	);
	LUT3 #(
		.INIT('h80)
	) name3166 (
		\a[1] ,
		\a[28] ,
		\a[54] ,
		_w3232_
	);
	LUT3 #(
		.INIT('h6c)
	) name3167 (
		\a[1] ,
		\a[28] ,
		\a[54] ,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name3168 (
		_w3127_,
		_w3233_,
		_w3234_
	);
	LUT3 #(
		.INIT('hb8)
	) name3169 (
		\a[54] ,
		_w3127_,
		_w3233_,
		_w3235_
	);
	LUT3 #(
		.INIT('h0d)
	) name3170 (
		_w2725_,
		_w3163_,
		_w3164_,
		_w3236_
	);
	LUT2 #(
		.INIT('h6)
	) name3171 (
		_w3235_,
		_w3236_,
		_w3237_
	);
	LUT3 #(
		.INIT('h69)
	) name3172 (
		_w3228_,
		_w3229_,
		_w3237_,
		_w3238_
	);
	LUT4 #(
		.INIT('hfe00)
	) name3173 (
		_w3197_,
		_w3199_,
		_w3226_,
		_w3238_,
		_w3239_
	);
	LUT4 #(
		.INIT('h0017)
	) name3174 (
		_w3162_,
		_w3178_,
		_w3195_,
		_w3238_,
		_w3240_
	);
	LUT3 #(
		.INIT('h0d)
	) name3175 (
		_w3190_,
		_w3191_,
		_w3192_,
		_w3241_
	);
	LUT3 #(
		.INIT('h0d)
	) name3176 (
		_w3179_,
		_w3180_,
		_w3181_,
		_w3242_
	);
	LUT3 #(
		.INIT('h32)
	) name3177 (
		_w3166_,
		_w3167_,
		_w3168_,
		_w3243_
	);
	LUT3 #(
		.INIT('h96)
	) name3178 (
		_w3241_,
		_w3242_,
		_w3243_,
		_w3244_
	);
	LUT3 #(
		.INIT('h32)
	) name3179 (
		_w3124_,
		_w3125_,
		_w3130_,
		_w3245_
	);
	LUT3 #(
		.INIT('he8)
	) name3180 (
		_w3077_,
		_w3128_,
		_w3129_,
		_w3246_
	);
	LUT3 #(
		.INIT('h32)
	) name3181 (
		_w3183_,
		_w3184_,
		_w3185_,
		_w3247_
	);
	LUT2 #(
		.INIT('h8)
	) name3182 (
		\a[5] ,
		\a[50] ,
		_w3248_
	);
	LUT4 #(
		.INIT('h153f)
	) name3183 (
		\a[18] ,
		\a[19] ,
		\a[36] ,
		\a[37] ,
		_w3249_
	);
	LUT4 #(
		.INIT('h8000)
	) name3184 (
		\a[18] ,
		\a[19] ,
		\a[36] ,
		\a[37] ,
		_w3250_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3185 (
		\a[18] ,
		\a[19] ,
		\a[36] ,
		\a[37] ,
		_w3251_
	);
	LUT2 #(
		.INIT('h6)
	) name3186 (
		_w3248_,
		_w3251_,
		_w3252_
	);
	LUT3 #(
		.INIT('h96)
	) name3187 (
		_w3246_,
		_w3247_,
		_w3252_,
		_w3253_
	);
	LUT3 #(
		.INIT('h96)
	) name3188 (
		_w3244_,
		_w3245_,
		_w3253_,
		_w3254_
	);
	LUT4 #(
		.INIT('hf40b)
	) name3189 (
		_w3227_,
		_w3238_,
		_w3240_,
		_w3254_,
		_w3255_
	);
	LUT3 #(
		.INIT('he8)
	) name3190 (
		_w3142_,
		_w3143_,
		_w3144_,
		_w3256_
	);
	LUT2 #(
		.INIT('h8)
	) name3191 (
		\a[10] ,
		\a[45] ,
		_w3257_
	);
	LUT4 #(
		.INIT('h153f)
	) name3192 (
		\a[11] ,
		\a[13] ,
		\a[42] ,
		\a[44] ,
		_w3258_
	);
	LUT4 #(
		.INIT('h8000)
	) name3193 (
		\a[11] ,
		\a[13] ,
		\a[42] ,
		\a[44] ,
		_w3259_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3194 (
		\a[11] ,
		\a[13] ,
		\a[42] ,
		\a[44] ,
		_w3260_
	);
	LUT2 #(
		.INIT('h8)
	) name3195 (
		\a[27] ,
		\a[28] ,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name3196 (
		\a[26] ,
		\a[29] ,
		_w3262_
	);
	LUT4 #(
		.INIT('h153f)
	) name3197 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w3263_
	);
	LUT4 #(
		.INIT('h8000)
	) name3198 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w3264_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3199 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w3265_
	);
	LUT4 #(
		.INIT('h1428)
	) name3200 (
		_w3042_,
		_w3257_,
		_w3260_,
		_w3265_,
		_w3266_
	);
	LUT4 #(
		.INIT('h8241)
	) name3201 (
		_w3042_,
		_w3257_,
		_w3260_,
		_w3265_,
		_w3267_
	);
	LUT4 #(
		.INIT('h6996)
	) name3202 (
		_w3042_,
		_w3257_,
		_w3260_,
		_w3265_,
		_w3268_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		\a[16] ,
		\a[39] ,
		_w3269_
	);
	LUT4 #(
		.INIT('h153f)
	) name3204 (
		\a[7] ,
		\a[8] ,
		\a[47] ,
		\a[48] ,
		_w3270_
	);
	LUT4 #(
		.INIT('h8000)
	) name3205 (
		\a[7] ,
		\a[8] ,
		\a[47] ,
		\a[48] ,
		_w3271_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3206 (
		\a[7] ,
		\a[8] ,
		\a[47] ,
		\a[48] ,
		_w3272_
	);
	LUT2 #(
		.INIT('h6)
	) name3207 (
		_w3269_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('h6)
	) name3208 (
		_w3268_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		\a[20] ,
		\a[35] ,
		_w3275_
	);
	LUT4 #(
		.INIT('h153f)
	) name3210 (
		\a[21] ,
		\a[22] ,
		\a[33] ,
		\a[34] ,
		_w3276_
	);
	LUT4 #(
		.INIT('h8000)
	) name3211 (
		\a[21] ,
		\a[22] ,
		\a[33] ,
		\a[34] ,
		_w3277_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3212 (
		\a[21] ,
		\a[22] ,
		\a[33] ,
		\a[34] ,
		_w3278_
	);
	LUT4 #(
		.INIT('h153f)
	) name3213 (
		\a[2] ,
		\a[4] ,
		\a[51] ,
		\a[53] ,
		_w3279_
	);
	LUT4 #(
		.INIT('h8000)
	) name3214 (
		\a[2] ,
		\a[4] ,
		\a[51] ,
		\a[53] ,
		_w3280_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3215 (
		\a[2] ,
		\a[4] ,
		\a[51] ,
		\a[53] ,
		_w3281_
	);
	LUT2 #(
		.INIT('h8)
	) name3216 (
		\a[0] ,
		\a[55] ,
		_w3282_
	);
	LUT4 #(
		.INIT('h0660)
	) name3217 (
		_w3275_,
		_w3278_,
		_w3281_,
		_w3282_,
		_w3283_
	);
	LUT4 #(
		.INIT('h9009)
	) name3218 (
		_w3275_,
		_w3278_,
		_w3281_,
		_w3282_,
		_w3284_
	);
	LUT4 #(
		.INIT('h6996)
	) name3219 (
		_w3275_,
		_w3278_,
		_w3281_,
		_w3282_,
		_w3285_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		\a[23] ,
		\a[32] ,
		_w3286_
	);
	LUT4 #(
		.INIT('h153f)
	) name3221 (
		\a[24] ,
		\a[25] ,
		\a[30] ,
		\a[31] ,
		_w3287_
	);
	LUT4 #(
		.INIT('h8000)
	) name3222 (
		\a[24] ,
		\a[25] ,
		\a[30] ,
		\a[31] ,
		_w3288_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3223 (
		\a[24] ,
		\a[25] ,
		\a[30] ,
		\a[31] ,
		_w3289_
	);
	LUT2 #(
		.INIT('h6)
	) name3224 (
		_w3286_,
		_w3289_,
		_w3290_
	);
	LUT2 #(
		.INIT('h6)
	) name3225 (
		_w3285_,
		_w3290_,
		_w3291_
	);
	LUT4 #(
		.INIT('h9009)
	) name3226 (
		_w3268_,
		_w3273_,
		_w3285_,
		_w3290_,
		_w3292_
	);
	LUT4 #(
		.INIT('h1700)
	) name3227 (
		_w3142_,
		_w3143_,
		_w3144_,
		_w3292_,
		_w3293_
	);
	LUT4 #(
		.INIT('h6006)
	) name3228 (
		_w3268_,
		_w3273_,
		_w3285_,
		_w3290_,
		_w3294_
	);
	LUT4 #(
		.INIT('he800)
	) name3229 (
		_w3142_,
		_w3143_,
		_w3144_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		_w3293_,
		_w3295_,
		_w3296_
	);
	LUT3 #(
		.INIT('h54)
	) name3231 (
		_w3132_,
		_w3133_,
		_w3134_,
		_w3297_
	);
	LUT3 #(
		.INIT('h0d)
	) name3232 (
		_w3120_,
		_w3121_,
		_w3122_,
		_w3298_
	);
	LUT3 #(
		.INIT('h0d)
	) name3233 (
		_w3116_,
		_w3117_,
		_w3118_,
		_w3299_
	);
	LUT3 #(
		.INIT('h0d)
	) name3234 (
		_w3173_,
		_w3174_,
		_w3175_,
		_w3300_
	);
	LUT3 #(
		.INIT('h96)
	) name3235 (
		_w3298_,
		_w3299_,
		_w3300_,
		_w3301_
	);
	LUT3 #(
		.INIT('h32)
	) name3236 (
		_w3187_,
		_w3188_,
		_w3194_,
		_w3302_
	);
	LUT3 #(
		.INIT('h32)
	) name3237 (
		_w3170_,
		_w3171_,
		_w3177_,
		_w3303_
	);
	LUT3 #(
		.INIT('h69)
	) name3238 (
		_w3301_,
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT4 #(
		.INIT('h0990)
	) name3239 (
		_w3268_,
		_w3273_,
		_w3285_,
		_w3290_,
		_w3305_
	);
	LUT4 #(
		.INIT('he800)
	) name3240 (
		_w3142_,
		_w3143_,
		_w3144_,
		_w3305_,
		_w3306_
	);
	LUT4 #(
		.INIT('h0660)
	) name3241 (
		_w3268_,
		_w3273_,
		_w3285_,
		_w3290_,
		_w3307_
	);
	LUT4 #(
		.INIT('h1700)
	) name3242 (
		_w3142_,
		_w3143_,
		_w3144_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h1)
	) name3243 (
		_w3306_,
		_w3308_,
		_w3309_
	);
	LUT3 #(
		.INIT('h02)
	) name3244 (
		_w3304_,
		_w3306_,
		_w3308_,
		_w3310_
	);
	LUT3 #(
		.INIT('h01)
	) name3245 (
		_w3304_,
		_w3306_,
		_w3308_,
		_w3311_
	);
	LUT4 #(
		.INIT('ha820)
	) name3246 (
		_w3296_,
		_w3297_,
		_w3310_,
		_w3311_,
		_w3312_
	);
	LUT3 #(
		.INIT('h96)
	) name3247 (
		_w3256_,
		_w3274_,
		_w3291_,
		_w3313_
	);
	LUT3 #(
		.INIT('hf6)
	) name3248 (
		_w3297_,
		_w3304_,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h4)
	) name3249 (
		_w3312_,
		_w3314_,
		_w3315_
	);
	LUT3 #(
		.INIT('hf9)
	) name3250 (
		_w3225_,
		_w3255_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h4)
	) name3251 (
		_w3225_,
		_w3255_,
		_w3317_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3252 (
		_w3086_,
		_w3114_,
		_w3115_,
		_w3255_,
		_w3318_
	);
	LUT3 #(
		.INIT('h4c)
	) name3253 (
		_w3136_,
		_w3315_,
		_w3318_,
		_w3319_
	);
	LUT4 #(
		.INIT('h2d00)
	) name3254 (
		_w3136_,
		_w3224_,
		_w3255_,
		_w3315_,
		_w3320_
	);
	LUT3 #(
		.INIT('he8)
	) name3255 (
		_w3141_,
		_w3161_,
		_w3211_,
		_w3321_
	);
	LUT3 #(
		.INIT('h0e)
	) name3256 (
		_w3200_,
		_w3208_,
		_w3209_,
		_w3322_
	);
	LUT2 #(
		.INIT('h8)
	) name3257 (
		\a[3] ,
		\a[52] ,
		_w3323_
	);
	LUT4 #(
		.INIT('h153f)
	) name3258 (
		\a[6] ,
		\a[17] ,
		\a[38] ,
		\a[49] ,
		_w3324_
	);
	LUT4 #(
		.INIT('h8000)
	) name3259 (
		\a[6] ,
		\a[17] ,
		\a[38] ,
		\a[49] ,
		_w3325_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3260 (
		\a[6] ,
		\a[17] ,
		\a[38] ,
		\a[49] ,
		_w3326_
	);
	LUT2 #(
		.INIT('h8)
	) name3261 (
		\a[15] ,
		\a[40] ,
		_w3327_
	);
	LUT4 #(
		.INIT('h153f)
	) name3262 (
		\a[9] ,
		\a[14] ,
		\a[41] ,
		\a[46] ,
		_w3328_
	);
	LUT4 #(
		.INIT('h8000)
	) name3263 (
		\a[9] ,
		\a[14] ,
		\a[41] ,
		\a[46] ,
		_w3329_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3264 (
		\a[9] ,
		\a[14] ,
		\a[41] ,
		\a[46] ,
		_w3330_
	);
	LUT4 #(
		.INIT('h0660)
	) name3265 (
		_w3323_,
		_w3326_,
		_w3327_,
		_w3330_,
		_w3331_
	);
	LUT4 #(
		.INIT('h6996)
	) name3266 (
		_w3323_,
		_w3326_,
		_w3327_,
		_w3330_,
		_w3332_
	);
	LUT4 #(
		.INIT('h1700)
	) name3267 (
		_w3155_,
		_w3156_,
		_w3157_,
		_w3332_,
		_w3333_
	);
	LUT4 #(
		.INIT('he817)
	) name3268 (
		_w3155_,
		_w3156_,
		_w3157_,
		_w3332_,
		_w3334_
	);
	LUT4 #(
		.INIT('h002b)
	) name3269 (
		_w3204_,
		_w3205_,
		_w3206_,
		_w3334_,
		_w3335_
	);
	LUT3 #(
		.INIT('h71)
	) name3270 (
		_w3154_,
		_w3158_,
		_w3159_,
		_w3336_
	);
	LUT4 #(
		.INIT('hd400)
	) name3271 (
		_w3204_,
		_w3205_,
		_w3206_,
		_w3334_,
		_w3337_
	);
	LUT3 #(
		.INIT('hc9)
	) name3272 (
		_w3335_,
		_w3336_,
		_w3337_,
		_w3338_
	);
	LUT4 #(
		.INIT('hdc00)
	) name3273 (
		_w3149_,
		_w3150_,
		_w3160_,
		_w3338_,
		_w3339_
	);
	LUT4 #(
		.INIT('h0023)
	) name3274 (
		_w3149_,
		_w3150_,
		_w3160_,
		_w3338_,
		_w3340_
	);
	LUT4 #(
		.INIT('h17e8)
	) name3275 (
		_w3145_,
		_w3148_,
		_w3160_,
		_w3338_,
		_w3341_
	);
	LUT2 #(
		.INIT('h6)
	) name3276 (
		_w3322_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name3277 (
		_w3321_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name3278 (
		_w3321_,
		_w3342_,
		_w3344_
	);
	LUT2 #(
		.INIT('h6)
	) name3279 (
		_w3321_,
		_w3342_,
		_w3345_
	);
	LUT3 #(
		.INIT('hd2)
	) name3280 (
		_w3316_,
		_w3320_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h8)
	) name3281 (
		_w3223_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h1)
	) name3282 (
		_w3223_,
		_w3346_,
		_w3348_
	);
	LUT2 #(
		.INIT('h6)
	) name3283 (
		_w3223_,
		_w3346_,
		_w3349_
	);
	LUT3 #(
		.INIT('he1)
	) name3284 (
		_w3215_,
		_w3222_,
		_w3349_,
		_w3350_
	);
	LUT3 #(
		.INIT('h01)
	) name3285 (
		_w3105_,
		_w3214_,
		_w3347_,
		_w3351_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3286 (
		_w2800_,
		_w3109_,
		_w3218_,
		_w3351_,
		_w3352_
	);
	LUT4 #(
		.INIT('h0111)
	) name3287 (
		_w3113_,
		_w3213_,
		_w3223_,
		_w3346_,
		_w3353_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3288 (
		_w3316_,
		_w3320_,
		_w3343_,
		_w3344_,
		_w3354_
	);
	LUT3 #(
		.INIT('h0e)
	) name3289 (
		_w3322_,
		_w3339_,
		_w3340_,
		_w3355_
	);
	LUT2 #(
		.INIT('h8)
	) name3290 (
		\a[11] ,
		\a[45] ,
		_w3356_
	);
	LUT4 #(
		.INIT('h153f)
	) name3291 (
		\a[12] ,
		\a[13] ,
		\a[43] ,
		\a[44] ,
		_w3357_
	);
	LUT4 #(
		.INIT('h8000)
	) name3292 (
		\a[12] ,
		\a[13] ,
		\a[43] ,
		\a[44] ,
		_w3358_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3293 (
		\a[12] ,
		\a[13] ,
		\a[43] ,
		\a[44] ,
		_w3359_
	);
	LUT2 #(
		.INIT('h8)
	) name3294 (
		\a[6] ,
		\a[50] ,
		_w3360_
	);
	LUT4 #(
		.INIT('h153f)
	) name3295 (
		\a[7] ,
		\a[17] ,
		\a[39] ,
		\a[49] ,
		_w3361_
	);
	LUT4 #(
		.INIT('h8000)
	) name3296 (
		\a[7] ,
		\a[17] ,
		\a[39] ,
		\a[49] ,
		_w3362_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3297 (
		\a[7] ,
		\a[17] ,
		\a[39] ,
		\a[49] ,
		_w3363_
	);
	LUT4 #(
		.INIT('h0660)
	) name3298 (
		_w3356_,
		_w3359_,
		_w3360_,
		_w3363_,
		_w3364_
	);
	LUT4 #(
		.INIT('h9009)
	) name3299 (
		_w3356_,
		_w3359_,
		_w3360_,
		_w3363_,
		_w3365_
	);
	LUT4 #(
		.INIT('h6996)
	) name3300 (
		_w3356_,
		_w3359_,
		_w3360_,
		_w3363_,
		_w3366_
	);
	LUT2 #(
		.INIT('h8)
	) name3301 (
		\a[16] ,
		\a[40] ,
		_w3367_
	);
	LUT4 #(
		.INIT('h153f)
	) name3302 (
		\a[8] ,
		\a[15] ,
		\a[41] ,
		\a[48] ,
		_w3368_
	);
	LUT2 #(
		.INIT('h8)
	) name3303 (
		\a[15] ,
		\a[48] ,
		_w3369_
	);
	LUT4 #(
		.INIT('h8000)
	) name3304 (
		\a[8] ,
		\a[15] ,
		\a[41] ,
		\a[48] ,
		_w3370_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3305 (
		\a[8] ,
		\a[15] ,
		\a[41] ,
		\a[48] ,
		_w3371_
	);
	LUT2 #(
		.INIT('h6)
	) name3306 (
		_w3367_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h8)
	) name3307 (
		\a[20] ,
		\a[36] ,
		_w3373_
	);
	LUT4 #(
		.INIT('h153f)
	) name3308 (
		\a[22] ,
		\a[23] ,
		\a[33] ,
		\a[34] ,
		_w3374_
	);
	LUT4 #(
		.INIT('h8000)
	) name3309 (
		\a[22] ,
		\a[23] ,
		\a[33] ,
		\a[34] ,
		_w3375_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3310 (
		\a[22] ,
		\a[23] ,
		\a[33] ,
		\a[34] ,
		_w3376_
	);
	LUT2 #(
		.INIT('h8)
	) name3311 (
		\a[24] ,
		\a[32] ,
		_w3377_
	);
	LUT4 #(
		.INIT('h153f)
	) name3312 (
		\a[25] ,
		\a[26] ,
		\a[30] ,
		\a[31] ,
		_w3378_
	);
	LUT4 #(
		.INIT('h8000)
	) name3313 (
		\a[25] ,
		\a[26] ,
		\a[30] ,
		\a[31] ,
		_w3379_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3314 (
		\a[25] ,
		\a[26] ,
		\a[30] ,
		\a[31] ,
		_w3380_
	);
	LUT4 #(
		.INIT('h0660)
	) name3315 (
		_w3373_,
		_w3376_,
		_w3377_,
		_w3380_,
		_w3381_
	);
	LUT4 #(
		.INIT('h9009)
	) name3316 (
		_w3373_,
		_w3376_,
		_w3377_,
		_w3380_,
		_w3382_
	);
	LUT4 #(
		.INIT('h6996)
	) name3317 (
		_w3373_,
		_w3376_,
		_w3377_,
		_w3380_,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name3318 (
		\a[9] ,
		\a[47] ,
		_w3384_
	);
	LUT4 #(
		.INIT('h153f)
	) name3319 (
		\a[10] ,
		\a[14] ,
		\a[42] ,
		\a[46] ,
		_w3385_
	);
	LUT2 #(
		.INIT('h8)
	) name3320 (
		\a[14] ,
		\a[46] ,
		_w3386_
	);
	LUT4 #(
		.INIT('h8000)
	) name3321 (
		\a[10] ,
		\a[14] ,
		\a[42] ,
		\a[46] ,
		_w3387_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3322 (
		\a[10] ,
		\a[14] ,
		\a[42] ,
		\a[46] ,
		_w3388_
	);
	LUT2 #(
		.INIT('h6)
	) name3323 (
		_w3384_,
		_w3388_,
		_w3389_
	);
	LUT4 #(
		.INIT('h0660)
	) name3324 (
		_w3366_,
		_w3372_,
		_w3383_,
		_w3389_,
		_w3390_
	);
	LUT4 #(
		.INIT('h9009)
	) name3325 (
		_w3366_,
		_w3372_,
		_w3383_,
		_w3389_,
		_w3391_
	);
	LUT4 #(
		.INIT('h6996)
	) name3326 (
		_w3366_,
		_w3372_,
		_w3383_,
		_w3389_,
		_w3392_
	);
	LUT4 #(
		.INIT('h153f)
	) name3327 (
		\a[0] ,
		\a[2] ,
		\a[54] ,
		\a[56] ,
		_w3393_
	);
	LUT2 #(
		.INIT('h8)
	) name3328 (
		\a[2] ,
		\a[56] ,
		_w3394_
	);
	LUT4 #(
		.INIT('h8000)
	) name3329 (
		\a[0] ,
		\a[2] ,
		\a[54] ,
		\a[56] ,
		_w3395_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3330 (
		\a[0] ,
		\a[2] ,
		\a[54] ,
		\a[56] ,
		_w3396_
	);
	LUT2 #(
		.INIT('h6)
	) name3331 (
		_w3232_,
		_w3396_,
		_w3397_
	);
	LUT3 #(
		.INIT('h0d)
	) name3332 (
		_w3269_,
		_w3270_,
		_w3271_,
		_w3398_
	);
	LUT2 #(
		.INIT('h8)
	) name3333 (
		\a[3] ,
		\a[53] ,
		_w3399_
	);
	LUT4 #(
		.INIT('h153f)
	) name3334 (
		\a[4] ,
		\a[19] ,
		\a[37] ,
		\a[52] ,
		_w3400_
	);
	LUT4 #(
		.INIT('h8000)
	) name3335 (
		\a[4] ,
		\a[19] ,
		\a[37] ,
		\a[52] ,
		_w3401_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3336 (
		\a[4] ,
		\a[19] ,
		\a[37] ,
		\a[52] ,
		_w3402_
	);
	LUT2 #(
		.INIT('h6)
	) name3337 (
		_w3399_,
		_w3402_,
		_w3403_
	);
	LUT3 #(
		.INIT('h69)
	) name3338 (
		_w3397_,
		_w3398_,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h6)
	) name3339 (
		_w3392_,
		_w3404_,
		_w3405_
	);
	LUT3 #(
		.INIT('h54)
	) name3340 (
		_w3335_,
		_w3336_,
		_w3337_,
		_w3406_
	);
	LUT3 #(
		.INIT('h0d)
	) name3341 (
		_w3275_,
		_w3276_,
		_w3277_,
		_w3407_
	);
	LUT3 #(
		.INIT('h0d)
	) name3342 (
		_w3286_,
		_w3287_,
		_w3288_,
		_w3408_
	);
	LUT3 #(
		.INIT('h0d)
	) name3343 (
		_w3323_,
		_w3324_,
		_w3325_,
		_w3409_
	);
	LUT3 #(
		.INIT('h96)
	) name3344 (
		_w3407_,
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('h8000)
	) name3345 (
		\a[1] ,
		\a[27] ,
		\a[29] ,
		\a[55] ,
		_w3411_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3346 (
		\a[1] ,
		\a[27] ,
		\a[29] ,
		\a[55] ,
		_w3412_
	);
	LUT4 #(
		.INIT('he800)
	) name3347 (
		_w3042_,
		_w3261_,
		_w3262_,
		_w3412_,
		_w3413_
	);
	LUT4 #(
		.INIT('h0017)
	) name3348 (
		_w3042_,
		_w3261_,
		_w3262_,
		_w3412_,
		_w3414_
	);
	LUT4 #(
		.INIT('hcd32)
	) name3349 (
		_w3042_,
		_w3263_,
		_w3264_,
		_w3412_,
		_w3415_
	);
	LUT3 #(
		.INIT('h0d)
	) name3350 (
		_w3257_,
		_w3258_,
		_w3259_,
		_w3416_
	);
	LUT2 #(
		.INIT('h6)
	) name3351 (
		_w3415_,
		_w3416_,
		_w3417_
	);
	LUT3 #(
		.INIT('h32)
	) name3352 (
		_w3266_,
		_w3267_,
		_w3273_,
		_w3418_
	);
	LUT3 #(
		.INIT('h96)
	) name3353 (
		_w3410_,
		_w3417_,
		_w3418_,
		_w3419_
	);
	LUT4 #(
		.INIT('h5400)
	) name3354 (
		_w3335_,
		_w3336_,
		_w3337_,
		_w3419_,
		_w3420_
	);
	LUT3 #(
		.INIT('h96)
	) name3355 (
		_w3405_,
		_w3406_,
		_w3419_,
		_w3421_
	);
	LUT3 #(
		.INIT('h23)
	) name3356 (
		_w3279_,
		_w3280_,
		_w3282_,
		_w3422_
	);
	LUT3 #(
		.INIT('h0d)
	) name3357 (
		_w3248_,
		_w3249_,
		_w3250_,
		_w3423_
	);
	LUT3 #(
		.INIT('h32)
	) name3358 (
		_w3327_,
		_w3328_,
		_w3329_,
		_w3424_
	);
	LUT3 #(
		.INIT('h96)
	) name3359 (
		_w3422_,
		_w3423_,
		_w3424_,
		_w3425_
	);
	LUT3 #(
		.INIT('h01)
	) name3360 (
		_w3331_,
		_w3333_,
		_w3425_,
		_w3426_
	);
	LUT3 #(
		.INIT('he0)
	) name3361 (
		_w3331_,
		_w3333_,
		_w3425_,
		_w3427_
	);
	LUT3 #(
		.INIT('h1e)
	) name3362 (
		_w3331_,
		_w3333_,
		_w3425_,
		_w3428_
	);
	LUT3 #(
		.INIT('h8e)
	) name3363 (
		_w3228_,
		_w3229_,
		_w3237_,
		_w3429_
	);
	LUT2 #(
		.INIT('h6)
	) name3364 (
		_w3428_,
		_w3429_,
		_w3430_
	);
	LUT3 #(
		.INIT('h17)
	) name3365 (
		_w3298_,
		_w3299_,
		_w3300_,
		_w3431_
	);
	LUT3 #(
		.INIT('he8)
	) name3366 (
		_w3246_,
		_w3247_,
		_w3252_,
		_w3432_
	);
	LUT3 #(
		.INIT('h32)
	) name3367 (
		_w3283_,
		_w3284_,
		_w3290_,
		_w3433_
	);
	LUT3 #(
		.INIT('h96)
	) name3368 (
		_w3431_,
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT4 #(
		.INIT('he800)
	) name3369 (
		_w3142_,
		_w3143_,
		_w3144_,
		_w3274_,
		_w3435_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name3370 (
		_w3306_,
		_w3308_,
		_w3434_,
		_w3435_,
		_w3436_
	);
	LUT4 #(
		.INIT('h0001)
	) name3371 (
		_w3306_,
		_w3308_,
		_w3434_,
		_w3435_,
		_w3437_
	);
	LUT4 #(
		.INIT('h17e8)
	) name3372 (
		_w3256_,
		_w3274_,
		_w3291_,
		_w3434_,
		_w3438_
	);
	LUT2 #(
		.INIT('h6)
	) name3373 (
		_w3430_,
		_w3438_,
		_w3439_
	);
	LUT3 #(
		.INIT('h96)
	) name3374 (
		_w3355_,
		_w3421_,
		_w3439_,
		_w3440_
	);
	LUT3 #(
		.INIT('h71)
	) name3375 (
		_w3241_,
		_w3242_,
		_w3243_,
		_w3441_
	);
	LUT3 #(
		.INIT('h23)
	) name3376 (
		_w3230_,
		_w3234_,
		_w3236_,
		_w3442_
	);
	LUT2 #(
		.INIT('h8)
	) name3377 (
		\a[21] ,
		\a[35] ,
		_w3443_
	);
	LUT4 #(
		.INIT('h153f)
	) name3378 (
		\a[5] ,
		\a[18] ,
		\a[38] ,
		\a[51] ,
		_w3444_
	);
	LUT4 #(
		.INIT('h8000)
	) name3379 (
		\a[5] ,
		\a[18] ,
		\a[38] ,
		\a[51] ,
		_w3445_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3380 (
		\a[5] ,
		\a[18] ,
		\a[38] ,
		\a[51] ,
		_w3446_
	);
	LUT2 #(
		.INIT('h6)
	) name3381 (
		_w3443_,
		_w3446_,
		_w3447_
	);
	LUT4 #(
		.INIT('h2300)
	) name3382 (
		_w3230_,
		_w3234_,
		_w3236_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('h00dc)
	) name3383 (
		_w3230_,
		_w3234_,
		_w3236_,
		_w3447_,
		_w3449_
	);
	LUT4 #(
		.INIT('hdc23)
	) name3384 (
		_w3230_,
		_w3234_,
		_w3236_,
		_w3447_,
		_w3450_
	);
	LUT2 #(
		.INIT('h6)
	) name3385 (
		_w3441_,
		_w3450_,
		_w3451_
	);
	LUT3 #(
		.INIT('hd4)
	) name3386 (
		_w3301_,
		_w3302_,
		_w3303_,
		_w3452_
	);
	LUT3 #(
		.INIT('he8)
	) name3387 (
		_w3244_,
		_w3245_,
		_w3253_,
		_w3453_
	);
	LUT3 #(
		.INIT('h96)
	) name3388 (
		_w3451_,
		_w3452_,
		_w3453_,
		_w3454_
	);
	LUT4 #(
		.INIT('h00cd)
	) name3389 (
		_w3239_,
		_w3240_,
		_w3254_,
		_w3454_,
		_w3455_
	);
	LUT4 #(
		.INIT('h3200)
	) name3390 (
		_w3239_,
		_w3240_,
		_w3254_,
		_w3454_,
		_w3456_
	);
	LUT4 #(
		.INIT('hcd32)
	) name3391 (
		_w3239_,
		_w3240_,
		_w3254_,
		_w3454_,
		_w3457_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3392 (
		_w3132_,
		_w3133_,
		_w3134_,
		_w3304_,
		_w3458_
	);
	LUT3 #(
		.INIT('h0e)
	) name3393 (
		_w3297_,
		_w3309_,
		_w3458_,
		_w3459_
	);
	LUT4 #(
		.INIT('hff96)
	) name3394 (
		_w3256_,
		_w3274_,
		_w3291_,
		_w3304_,
		_w3460_
	);
	LUT3 #(
		.INIT('he0)
	) name3395 (
		_w3296_,
		_w3297_,
		_w3460_,
		_w3461_
	);
	LUT3 #(
		.INIT('h95)
	) name3396 (
		_w3457_,
		_w3459_,
		_w3461_,
		_w3462_
	);
	LUT4 #(
		.INIT('he11e)
	) name3397 (
		_w3317_,
		_w3319_,
		_w3440_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w3354_,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h6)
	) name3399 (
		_w3354_,
		_w3463_,
		_w3465_
	);
	LUT4 #(
		.INIT('hfe01)
	) name3400 (
		_w3348_,
		_w3352_,
		_w3353_,
		_w3465_,
		_w3466_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3401 (
		_w3223_,
		_w3346_,
		_w3354_,
		_w3463_,
		_w3467_
	);
	LUT2 #(
		.INIT('h4)
	) name3402 (
		_w3353_,
		_w3467_,
		_w3468_
	);
	LUT3 #(
		.INIT('h15)
	) name3403 (
		_w3456_,
		_w3459_,
		_w3461_,
		_w3469_
	);
	LUT4 #(
		.INIT('h5444)
	) name3404 (
		_w3455_,
		_w3456_,
		_w3459_,
		_w3461_,
		_w3470_
	);
	LUT3 #(
		.INIT('h23)
	) name3405 (
		_w3413_,
		_w3414_,
		_w3416_,
		_w3471_
	);
	LUT3 #(
		.INIT('hb2)
	) name3406 (
		_w3397_,
		_w3398_,
		_w3403_,
		_w3472_
	);
	LUT3 #(
		.INIT('h32)
	) name3407 (
		_w3381_,
		_w3382_,
		_w3389_,
		_w3473_
	);
	LUT3 #(
		.INIT('h96)
	) name3408 (
		_w3471_,
		_w3472_,
		_w3473_,
		_w3474_
	);
	LUT3 #(
		.INIT('h32)
	) name3409 (
		_w3390_,
		_w3391_,
		_w3404_,
		_w3475_
	);
	LUT3 #(
		.INIT('h0d)
	) name3410 (
		_w3367_,
		_w3368_,
		_w3370_,
		_w3476_
	);
	LUT3 #(
		.INIT('h0d)
	) name3411 (
		_w3377_,
		_w3378_,
		_w3379_,
		_w3477_
	);
	LUT3 #(
		.INIT('h32)
	) name3412 (
		_w3360_,
		_w3361_,
		_w3362_,
		_w3478_
	);
	LUT3 #(
		.INIT('h96)
	) name3413 (
		_w3476_,
		_w3477_,
		_w3478_,
		_w3479_
	);
	LUT3 #(
		.INIT('h32)
	) name3414 (
		_w3399_,
		_w3400_,
		_w3401_,
		_w3480_
	);
	LUT3 #(
		.INIT('h0d)
	) name3415 (
		_w3373_,
		_w3374_,
		_w3375_,
		_w3481_
	);
	LUT3 #(
		.INIT('h0d)
	) name3416 (
		_w3232_,
		_w3393_,
		_w3395_,
		_w3482_
	);
	LUT3 #(
		.INIT('h69)
	) name3417 (
		_w3480_,
		_w3481_,
		_w3482_,
		_w3483_
	);
	LUT3 #(
		.INIT('h32)
	) name3418 (
		_w3364_,
		_w3365_,
		_w3372_,
		_w3484_
	);
	LUT3 #(
		.INIT('h69)
	) name3419 (
		_w3479_,
		_w3483_,
		_w3484_,
		_w3485_
	);
	LUT3 #(
		.INIT('h96)
	) name3420 (
		_w3474_,
		_w3475_,
		_w3485_,
		_w3486_
	);
	LUT3 #(
		.INIT('he8)
	) name3421 (
		_w3451_,
		_w3452_,
		_w3453_,
		_w3487_
	);
	LUT2 #(
		.INIT('h8)
	) name3422 (
		\a[3] ,
		\a[54] ,
		_w3488_
	);
	LUT4 #(
		.INIT('h153f)
	) name3423 (
		\a[2] ,
		\a[4] ,
		\a[53] ,
		\a[55] ,
		_w3489_
	);
	LUT2 #(
		.INIT('h8)
	) name3424 (
		\a[4] ,
		\a[55] ,
		_w3490_
	);
	LUT4 #(
		.INIT('h8000)
	) name3425 (
		\a[2] ,
		\a[4] ,
		\a[53] ,
		\a[55] ,
		_w3491_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3426 (
		\a[2] ,
		\a[4] ,
		\a[53] ,
		\a[55] ,
		_w3492_
	);
	LUT2 #(
		.INIT('h8)
	) name3427 (
		\a[5] ,
		\a[52] ,
		_w3493_
	);
	LUT4 #(
		.INIT('h153f)
	) name3428 (
		\a[19] ,
		\a[20] ,
		\a[37] ,
		\a[38] ,
		_w3494_
	);
	LUT4 #(
		.INIT('h8000)
	) name3429 (
		\a[19] ,
		\a[20] ,
		\a[37] ,
		\a[38] ,
		_w3495_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3430 (
		\a[19] ,
		\a[20] ,
		\a[37] ,
		\a[38] ,
		_w3496_
	);
	LUT4 #(
		.INIT('h0660)
	) name3431 (
		_w3488_,
		_w3492_,
		_w3493_,
		_w3496_,
		_w3497_
	);
	LUT4 #(
		.INIT('h9009)
	) name3432 (
		_w3488_,
		_w3492_,
		_w3493_,
		_w3496_,
		_w3498_
	);
	LUT4 #(
		.INIT('h6996)
	) name3433 (
		_w3488_,
		_w3492_,
		_w3493_,
		_w3496_,
		_w3499_
	);
	LUT2 #(
		.INIT('h8)
	) name3434 (
		\a[15] ,
		\a[42] ,
		_w3500_
	);
	LUT4 #(
		.INIT('h153f)
	) name3435 (
		\a[9] ,
		\a[10] ,
		\a[47] ,
		\a[48] ,
		_w3501_
	);
	LUT2 #(
		.INIT('h8)
	) name3436 (
		\a[10] ,
		\a[48] ,
		_w3502_
	);
	LUT4 #(
		.INIT('h8000)
	) name3437 (
		\a[9] ,
		\a[10] ,
		\a[47] ,
		\a[48] ,
		_w3503_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3438 (
		\a[9] ,
		\a[10] ,
		\a[47] ,
		\a[48] ,
		_w3504_
	);
	LUT2 #(
		.INIT('h6)
	) name3439 (
		_w3500_,
		_w3504_,
		_w3505_
	);
	LUT4 #(
		.INIT('h153f)
	) name3440 (
		\a[11] ,
		\a[13] ,
		\a[44] ,
		\a[46] ,
		_w3506_
	);
	LUT2 #(
		.INIT('h8)
	) name3441 (
		\a[13] ,
		\a[46] ,
		_w3507_
	);
	LUT4 #(
		.INIT('h8000)
	) name3442 (
		\a[11] ,
		\a[13] ,
		\a[44] ,
		\a[46] ,
		_w3508_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3443 (
		\a[11] ,
		\a[13] ,
		\a[44] ,
		\a[46] ,
		_w3509_
	);
	LUT2 #(
		.INIT('h8)
	) name3444 (
		\a[12] ,
		\a[45] ,
		_w3510_
	);
	LUT4 #(
		.INIT('h153f)
	) name3445 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w3511_
	);
	LUT4 #(
		.INIT('h8000)
	) name3446 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w3512_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3447 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w3513_
	);
	LUT4 #(
		.INIT('h0660)
	) name3448 (
		_w2633_,
		_w3509_,
		_w3510_,
		_w3513_,
		_w3514_
	);
	LUT4 #(
		.INIT('h9009)
	) name3449 (
		_w2633_,
		_w3509_,
		_w3510_,
		_w3513_,
		_w3515_
	);
	LUT4 #(
		.INIT('h6996)
	) name3450 (
		_w2633_,
		_w3509_,
		_w3510_,
		_w3513_,
		_w3516_
	);
	LUT2 #(
		.INIT('h8)
	) name3451 (
		\a[18] ,
		\a[39] ,
		_w3517_
	);
	LUT4 #(
		.INIT('h153f)
	) name3452 (
		\a[6] ,
		\a[17] ,
		\a[40] ,
		\a[51] ,
		_w3518_
	);
	LUT4 #(
		.INIT('h8000)
	) name3453 (
		\a[6] ,
		\a[17] ,
		\a[40] ,
		\a[51] ,
		_w3519_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3454 (
		\a[6] ,
		\a[17] ,
		\a[40] ,
		\a[51] ,
		_w3520_
	);
	LUT2 #(
		.INIT('h6)
	) name3455 (
		_w3517_,
		_w3520_,
		_w3521_
	);
	LUT4 #(
		.INIT('h0660)
	) name3456 (
		_w3499_,
		_w3505_,
		_w3516_,
		_w3521_,
		_w3522_
	);
	LUT4 #(
		.INIT('h6996)
	) name3457 (
		_w3499_,
		_w3505_,
		_w3516_,
		_w3521_,
		_w3523_
	);
	LUT4 #(
		.INIT('he800)
	) name3458 (
		_w3431_,
		_w3432_,
		_w3433_,
		_w3523_,
		_w3524_
	);
	LUT4 #(
		.INIT('h17e8)
	) name3459 (
		_w3431_,
		_w3432_,
		_w3433_,
		_w3523_,
		_w3525_
	);
	LUT3 #(
		.INIT('h0d)
	) name3460 (
		_w3443_,
		_w3444_,
		_w3445_,
		_w3526_
	);
	LUT3 #(
		.INIT('h0d)
	) name3461 (
		_w3384_,
		_w3385_,
		_w3387_,
		_w3527_
	);
	LUT3 #(
		.INIT('h0d)
	) name3462 (
		_w3356_,
		_w3357_,
		_w3358_,
		_w3528_
	);
	LUT3 #(
		.INIT('h96)
	) name3463 (
		_w3526_,
		_w3527_,
		_w3528_,
		_w3529_
	);
	LUT4 #(
		.INIT('h1700)
	) name3464 (
		_w3441_,
		_w3442_,
		_w3447_,
		_w3529_,
		_w3530_
	);
	LUT4 #(
		.INIT('h00e8)
	) name3465 (
		_w3441_,
		_w3442_,
		_w3447_,
		_w3529_,
		_w3531_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name3466 (
		_w3441_,
		_w3448_,
		_w3449_,
		_w3529_,
		_w3532_
	);
	LUT2 #(
		.INIT('h8)
	) name3467 (
		\a[7] ,
		\a[50] ,
		_w3533_
	);
	LUT4 #(
		.INIT('h153f)
	) name3468 (
		\a[8] ,
		\a[16] ,
		\a[41] ,
		\a[49] ,
		_w3534_
	);
	LUT2 #(
		.INIT('h8)
	) name3469 (
		\a[16] ,
		\a[49] ,
		_w3535_
	);
	LUT4 #(
		.INIT('h8000)
	) name3470 (
		\a[8] ,
		\a[16] ,
		\a[41] ,
		\a[49] ,
		_w3536_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3471 (
		\a[8] ,
		\a[16] ,
		\a[41] ,
		\a[49] ,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name3472 (
		\a[21] ,
		\a[36] ,
		_w3538_
	);
	LUT4 #(
		.INIT('h153f)
	) name3473 (
		\a[22] ,
		\a[23] ,
		\a[34] ,
		\a[35] ,
		_w3539_
	);
	LUT4 #(
		.INIT('h8000)
	) name3474 (
		\a[22] ,
		\a[23] ,
		\a[34] ,
		\a[35] ,
		_w3540_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3475 (
		\a[22] ,
		\a[23] ,
		\a[34] ,
		\a[35] ,
		_w3541_
	);
	LUT4 #(
		.INIT('h0660)
	) name3476 (
		_w3533_,
		_w3537_,
		_w3538_,
		_w3541_,
		_w3542_
	);
	LUT4 #(
		.INIT('h9009)
	) name3477 (
		_w3533_,
		_w3537_,
		_w3538_,
		_w3541_,
		_w3543_
	);
	LUT4 #(
		.INIT('h6996)
	) name3478 (
		_w3533_,
		_w3537_,
		_w3538_,
		_w3541_,
		_w3544_
	);
	LUT2 #(
		.INIT('h8)
	) name3479 (
		\a[24] ,
		\a[33] ,
		_w3545_
	);
	LUT4 #(
		.INIT('h153f)
	) name3480 (
		\a[25] ,
		\a[26] ,
		\a[31] ,
		\a[32] ,
		_w3546_
	);
	LUT4 #(
		.INIT('h8000)
	) name3481 (
		\a[25] ,
		\a[26] ,
		\a[31] ,
		\a[32] ,
		_w3547_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3482 (
		\a[25] ,
		\a[26] ,
		\a[31] ,
		\a[32] ,
		_w3548_
	);
	LUT2 #(
		.INIT('h6)
	) name3483 (
		_w3545_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h6)
	) name3484 (
		_w3544_,
		_w3549_,
		_w3550_
	);
	LUT4 #(
		.INIT('h6996)
	) name3485 (
		_w3487_,
		_w3525_,
		_w3532_,
		_w3550_,
		_w3551_
	);
	LUT3 #(
		.INIT('h9f)
	) name3486 (
		_w3470_,
		_w3486_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h1)
	) name3487 (
		_w3455_,
		_w3551_,
		_w3553_
	);
	LUT3 #(
		.INIT('h40)
	) name3488 (
		_w3469_,
		_w3486_,
		_w3553_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name3489 (
		_w3486_,
		_w3551_,
		_w3555_
	);
	LUT2 #(
		.INIT('h4)
	) name3490 (
		_w3470_,
		_w3555_,
		_w3556_
	);
	LUT3 #(
		.INIT('h02)
	) name3491 (
		_w3552_,
		_w3554_,
		_w3556_,
		_w3557_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3492 (
		_w3335_,
		_w3336_,
		_w3337_,
		_w3419_,
		_w3558_
	);
	LUT3 #(
		.INIT('h0e)
	) name3493 (
		_w3405_,
		_w3420_,
		_w3558_,
		_w3559_
	);
	LUT3 #(
		.INIT('h0e)
	) name3494 (
		_w3430_,
		_w3436_,
		_w3437_,
		_w3560_
	);
	LUT3 #(
		.INIT('h54)
	) name3495 (
		_w3426_,
		_w3427_,
		_w3429_,
		_w3561_
	);
	LUT3 #(
		.INIT('h17)
	) name3496 (
		_w3407_,
		_w3408_,
		_w3409_,
		_w3562_
	);
	LUT2 #(
		.INIT('h8)
	) name3497 (
		\a[0] ,
		\a[57] ,
		_w3563_
	);
	LUT3 #(
		.INIT('h80)
	) name3498 (
		\a[1] ,
		\a[29] ,
		\a[56] ,
		_w3564_
	);
	LUT3 #(
		.INIT('h6c)
	) name3499 (
		\a[1] ,
		\a[29] ,
		\a[56] ,
		_w3565_
	);
	LUT3 #(
		.INIT('h96)
	) name3500 (
		_w3411_,
		_w3563_,
		_w3565_,
		_w3566_
	);
	LUT4 #(
		.INIT('h00e8)
	) name3501 (
		_w3407_,
		_w3408_,
		_w3409_,
		_w3566_,
		_w3567_
	);
	LUT4 #(
		.INIT('h1700)
	) name3502 (
		_w3407_,
		_w3408_,
		_w3409_,
		_w3566_,
		_w3568_
	);
	LUT4 #(
		.INIT('he817)
	) name3503 (
		_w3407_,
		_w3408_,
		_w3409_,
		_w3566_,
		_w3569_
	);
	LUT3 #(
		.INIT('h71)
	) name3504 (
		_w3422_,
		_w3423_,
		_w3424_,
		_w3570_
	);
	LUT2 #(
		.INIT('h6)
	) name3505 (
		_w3569_,
		_w3570_,
		_w3571_
	);
	LUT3 #(
		.INIT('h71)
	) name3506 (
		_w3410_,
		_w3417_,
		_w3418_,
		_w3572_
	);
	LUT3 #(
		.INIT('h69)
	) name3507 (
		_w3561_,
		_w3571_,
		_w3572_,
		_w3573_
	);
	LUT3 #(
		.INIT('h69)
	) name3508 (
		_w3559_,
		_w3560_,
		_w3573_,
		_w3574_
	);
	LUT4 #(
		.INIT('he800)
	) name3509 (
		_w3355_,
		_w3421_,
		_w3439_,
		_w3574_,
		_w3575_
	);
	LUT4 #(
		.INIT('h17e8)
	) name3510 (
		_w3355_,
		_w3421_,
		_w3439_,
		_w3574_,
		_w3576_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3511 (
		_w3552_,
		_w3554_,
		_w3556_,
		_w3576_,
		_w3577_
	);
	LUT4 #(
		.INIT('he0fe)
	) name3512 (
		_w3317_,
		_w3319_,
		_w3440_,
		_w3462_,
		_w3578_
	);
	LUT4 #(
		.INIT('h0200)
	) name3513 (
		_w3552_,
		_w3554_,
		_w3556_,
		_w3576_,
		_w3579_
	);
	LUT3 #(
		.INIT('h04)
	) name3514 (
		_w3577_,
		_w3578_,
		_w3579_,
		_w3580_
	);
	LUT4 #(
		.INIT('hfd02)
	) name3515 (
		_w3552_,
		_w3554_,
		_w3556_,
		_w3576_,
		_w3581_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		_w3578_,
		_w3581_,
		_w3582_
	);
	LUT3 #(
		.INIT('h96)
	) name3517 (
		_w3557_,
		_w3576_,
		_w3578_,
		_w3583_
	);
	LUT4 #(
		.INIT('h23dc)
	) name3518 (
		_w3352_,
		_w3464_,
		_w3468_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h1)
	) name3519 (
		_w3464_,
		_w3580_,
		_w3585_
	);
	LUT4 #(
		.INIT('h0017)
	) name3520 (
		_w3355_,
		_w3421_,
		_w3439_,
		_w3574_,
		_w3586_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3521 (
		_w3552_,
		_w3554_,
		_w3556_,
		_w3575_,
		_w3587_
	);
	LUT2 #(
		.INIT('h4)
	) name3522 (
		_w3455_,
		_w3486_,
		_w3588_
	);
	LUT2 #(
		.INIT('h4)
	) name3523 (
		_w3469_,
		_w3588_,
		_w3589_
	);
	LUT3 #(
		.INIT('he8)
	) name3524 (
		_w3474_,
		_w3475_,
		_w3485_,
		_w3590_
	);
	LUT3 #(
		.INIT('h54)
	) name3525 (
		_w3530_,
		_w3531_,
		_w3550_,
		_w3591_
	);
	LUT3 #(
		.INIT('h17)
	) name3526 (
		_w3526_,
		_w3527_,
		_w3528_,
		_w3592_
	);
	LUT3 #(
		.INIT('h2b)
	) name3527 (
		_w3480_,
		_w3481_,
		_w3482_,
		_w3593_
	);
	LUT3 #(
		.INIT('h71)
	) name3528 (
		_w3476_,
		_w3477_,
		_w3478_,
		_w3594_
	);
	LUT3 #(
		.INIT('h96)
	) name3529 (
		_w3592_,
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT3 #(
		.INIT('hb2)
	) name3530 (
		_w3479_,
		_w3483_,
		_w3484_,
		_w3596_
	);
	LUT2 #(
		.INIT('h8)
	) name3531 (
		_w3595_,
		_w3596_,
		_w3597_
	);
	LUT2 #(
		.INIT('h1)
	) name3532 (
		_w3595_,
		_w3596_,
		_w3598_
	);
	LUT2 #(
		.INIT('h6)
	) name3533 (
		_w3595_,
		_w3596_,
		_w3599_
	);
	LUT2 #(
		.INIT('h6)
	) name3534 (
		_w3591_,
		_w3599_,
		_w3600_
	);
	LUT3 #(
		.INIT('h41)
	) name3535 (
		_w3590_,
		_w3591_,
		_w3599_,
		_w3601_
	);
	LUT3 #(
		.INIT('h28)
	) name3536 (
		_w3590_,
		_w3591_,
		_w3599_,
		_w3602_
	);
	LUT3 #(
		.INIT('h96)
	) name3537 (
		_w3590_,
		_w3591_,
		_w3599_,
		_w3603_
	);
	LUT4 #(
		.INIT('h7117)
	) name3538 (
		_w3487_,
		_w3525_,
		_w3532_,
		_w3550_,
		_w3604_
	);
	LUT2 #(
		.INIT('h2)
	) name3539 (
		_w3603_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h9)
	) name3540 (
		_w3603_,
		_w3604_,
		_w3606_
	);
	LUT3 #(
		.INIT('h8e)
	) name3541 (
		_w3559_,
		_w3560_,
		_w3573_,
		_w3607_
	);
	LUT4 #(
		.INIT('h8000)
	) name3542 (
		\a[1] ,
		\a[28] ,
		\a[30] ,
		\a[57] ,
		_w3608_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3543 (
		\a[1] ,
		\a[28] ,
		\a[30] ,
		\a[57] ,
		_w3609_
	);
	LUT2 #(
		.INIT('h1)
	) name3544 (
		_w3564_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		_w3564_,
		_w3609_,
		_w3611_
	);
	LUT2 #(
		.INIT('h6)
	) name3546 (
		_w3564_,
		_w3609_,
		_w3612_
	);
	LUT3 #(
		.INIT('h0d)
	) name3547 (
		_w3510_,
		_w3511_,
		_w3512_,
		_w3613_
	);
	LUT2 #(
		.INIT('h6)
	) name3548 (
		_w3612_,
		_w3613_,
		_w3614_
	);
	LUT3 #(
		.INIT('h32)
	) name3549 (
		_w3497_,
		_w3498_,
		_w3505_,
		_w3615_
	);
	LUT3 #(
		.INIT('h32)
	) name3550 (
		_w3514_,
		_w3515_,
		_w3521_,
		_w3616_
	);
	LUT3 #(
		.INIT('h69)
	) name3551 (
		_w3614_,
		_w3615_,
		_w3616_,
		_w3617_
	);
	LUT3 #(
		.INIT('h0d)
	) name3552 (
		_w3500_,
		_w3501_,
		_w3503_,
		_w3618_
	);
	LUT3 #(
		.INIT('h0d)
	) name3553 (
		_w3545_,
		_w3546_,
		_w3547_,
		_w3619_
	);
	LUT3 #(
		.INIT('h0d)
	) name3554 (
		_w3538_,
		_w3539_,
		_w3540_,
		_w3620_
	);
	LUT3 #(
		.INIT('h96)
	) name3555 (
		_w3618_,
		_w3619_,
		_w3620_,
		_w3621_
	);
	LUT3 #(
		.INIT('h0d)
	) name3556 (
		_w3493_,
		_w3494_,
		_w3495_,
		_w3622_
	);
	LUT3 #(
		.INIT('h0d)
	) name3557 (
		_w3488_,
		_w3489_,
		_w3491_,
		_w3623_
	);
	LUT3 #(
		.INIT('h0d)
	) name3558 (
		_w2633_,
		_w3506_,
		_w3508_,
		_w3624_
	);
	LUT3 #(
		.INIT('h96)
	) name3559 (
		_w3622_,
		_w3623_,
		_w3624_,
		_w3625_
	);
	LUT3 #(
		.INIT('h32)
	) name3560 (
		_w3542_,
		_w3543_,
		_w3549_,
		_w3626_
	);
	LUT3 #(
		.INIT('h96)
	) name3561 (
		_w3621_,
		_w3625_,
		_w3626_,
		_w3627_
	);
	LUT4 #(
		.INIT('he11e)
	) name3562 (
		_w3522_,
		_w3524_,
		_w3617_,
		_w3627_,
		_w3628_
	);
	LUT3 #(
		.INIT('h17)
	) name3563 (
		_w3561_,
		_w3571_,
		_w3572_,
		_w3629_
	);
	LUT3 #(
		.INIT('h54)
	) name3564 (
		_w3567_,
		_w3568_,
		_w3570_,
		_w3630_
	);
	LUT4 #(
		.INIT('h153f)
	) name3565 (
		\a[11] ,
		\a[15] ,
		\a[43] ,
		\a[47] ,
		_w3631_
	);
	LUT4 #(
		.INIT('h8000)
	) name3566 (
		\a[11] ,
		\a[15] ,
		\a[43] ,
		\a[47] ,
		_w3632_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3567 (
		\a[11] ,
		\a[15] ,
		\a[43] ,
		\a[47] ,
		_w3633_
	);
	LUT4 #(
		.INIT('h153f)
	) name3568 (
		\a[12] ,
		\a[13] ,
		\a[45] ,
		\a[46] ,
		_w3634_
	);
	LUT4 #(
		.INIT('h8000)
	) name3569 (
		\a[12] ,
		\a[13] ,
		\a[45] ,
		\a[46] ,
		_w3635_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3570 (
		\a[12] ,
		\a[13] ,
		\a[45] ,
		\a[46] ,
		_w3636_
	);
	LUT4 #(
		.INIT('h1428)
	) name3571 (
		_w3021_,
		_w3502_,
		_w3633_,
		_w3636_,
		_w3637_
	);
	LUT4 #(
		.INIT('h8241)
	) name3572 (
		_w3021_,
		_w3502_,
		_w3633_,
		_w3636_,
		_w3638_
	);
	LUT4 #(
		.INIT('h6996)
	) name3573 (
		_w3021_,
		_w3502_,
		_w3633_,
		_w3636_,
		_w3639_
	);
	LUT2 #(
		.INIT('h8)
	) name3574 (
		\a[3] ,
		\a[55] ,
		_w3640_
	);
	LUT4 #(
		.INIT('h153f)
	) name3575 (
		\a[6] ,
		\a[19] ,
		\a[39] ,
		\a[52] ,
		_w3641_
	);
	LUT4 #(
		.INIT('h8000)
	) name3576 (
		\a[6] ,
		\a[19] ,
		\a[39] ,
		\a[52] ,
		_w3642_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3577 (
		\a[6] ,
		\a[19] ,
		\a[39] ,
		\a[52] ,
		_w3643_
	);
	LUT2 #(
		.INIT('h6)
	) name3578 (
		_w3640_,
		_w3643_,
		_w3644_
	);
	LUT2 #(
		.INIT('h6)
	) name3579 (
		_w3639_,
		_w3644_,
		_w3645_
	);
	LUT3 #(
		.INIT('h0d)
	) name3580 (
		_w3517_,
		_w3518_,
		_w3519_,
		_w3646_
	);
	LUT3 #(
		.INIT('h0d)
	) name3581 (
		_w3533_,
		_w3534_,
		_w3536_,
		_w3647_
	);
	LUT3 #(
		.INIT('he8)
	) name3582 (
		_w3411_,
		_w3563_,
		_w3565_,
		_w3648_
	);
	LUT3 #(
		.INIT('h96)
	) name3583 (
		_w3646_,
		_w3647_,
		_w3648_,
		_w3649_
	);
	LUT4 #(
		.INIT('h00e8)
	) name3584 (
		_w3562_,
		_w3566_,
		_w3570_,
		_w3649_,
		_w3650_
	);
	LUT4 #(
		.INIT('hed61)
	) name3585 (
		_w3630_,
		_w3645_,
		_w3649_,
		_w3650_,
		_w3651_
	);
	LUT4 #(
		.INIT('h00e8)
	) name3586 (
		_w3561_,
		_w3571_,
		_w3572_,
		_w3651_,
		_w3652_
	);
	LUT2 #(
		.INIT('h8)
	) name3587 (
		\a[5] ,
		\a[53] ,
		_w3653_
	);
	LUT4 #(
		.INIT('h153f)
	) name3588 (
		\a[20] ,
		\a[21] ,
		\a[37] ,
		\a[38] ,
		_w3654_
	);
	LUT4 #(
		.INIT('h8000)
	) name3589 (
		\a[20] ,
		\a[21] ,
		\a[37] ,
		\a[38] ,
		_w3655_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3590 (
		\a[20] ,
		\a[21] ,
		\a[37] ,
		\a[38] ,
		_w3656_
	);
	LUT4 #(
		.INIT('h153f)
	) name3591 (
		\a[0] ,
		\a[4] ,
		\a[54] ,
		\a[58] ,
		_w3657_
	);
	LUT4 #(
		.INIT('h8000)
	) name3592 (
		\a[0] ,
		\a[4] ,
		\a[54] ,
		\a[58] ,
		_w3658_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3593 (
		\a[0] ,
		\a[4] ,
		\a[54] ,
		\a[58] ,
		_w3659_
	);
	LUT4 #(
		.INIT('h1428)
	) name3594 (
		_w3394_,
		_w3653_,
		_w3656_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('h8241)
	) name3595 (
		_w3394_,
		_w3653_,
		_w3656_,
		_w3659_,
		_w3661_
	);
	LUT4 #(
		.INIT('h6996)
	) name3596 (
		_w3394_,
		_w3653_,
		_w3656_,
		_w3659_,
		_w3662_
	);
	LUT2 #(
		.INIT('h8)
	) name3597 (
		\a[17] ,
		\a[41] ,
		_w3663_
	);
	LUT4 #(
		.INIT('h153f)
	) name3598 (
		\a[9] ,
		\a[16] ,
		\a[42] ,
		\a[49] ,
		_w3664_
	);
	LUT4 #(
		.INIT('h8000)
	) name3599 (
		\a[9] ,
		\a[16] ,
		\a[42] ,
		\a[49] ,
		_w3665_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3600 (
		\a[9] ,
		\a[16] ,
		\a[42] ,
		\a[49] ,
		_w3666_
	);
	LUT2 #(
		.INIT('h6)
	) name3601 (
		_w3663_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h8)
	) name3602 (
		\a[18] ,
		\a[40] ,
		_w3668_
	);
	LUT4 #(
		.INIT('h153f)
	) name3603 (
		\a[7] ,
		\a[8] ,
		\a[50] ,
		\a[51] ,
		_w3669_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		\a[8] ,
		\a[51] ,
		_w3670_
	);
	LUT4 #(
		.INIT('h8000)
	) name3605 (
		\a[7] ,
		\a[8] ,
		\a[50] ,
		\a[51] ,
		_w3671_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3606 (
		\a[7] ,
		\a[8] ,
		\a[50] ,
		\a[51] ,
		_w3672_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		\a[22] ,
		\a[36] ,
		_w3673_
	);
	LUT4 #(
		.INIT('h153f)
	) name3608 (
		\a[23] ,
		\a[24] ,
		\a[34] ,
		\a[35] ,
		_w3674_
	);
	LUT4 #(
		.INIT('h8000)
	) name3609 (
		\a[23] ,
		\a[24] ,
		\a[34] ,
		\a[35] ,
		_w3675_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3610 (
		\a[23] ,
		\a[24] ,
		\a[34] ,
		\a[35] ,
		_w3676_
	);
	LUT4 #(
		.INIT('h0660)
	) name3611 (
		_w3668_,
		_w3672_,
		_w3673_,
		_w3676_,
		_w3677_
	);
	LUT4 #(
		.INIT('h9009)
	) name3612 (
		_w3668_,
		_w3672_,
		_w3673_,
		_w3676_,
		_w3678_
	);
	LUT4 #(
		.INIT('h6996)
	) name3613 (
		_w3668_,
		_w3672_,
		_w3673_,
		_w3676_,
		_w3679_
	);
	LUT2 #(
		.INIT('h8)
	) name3614 (
		\a[25] ,
		\a[33] ,
		_w3680_
	);
	LUT4 #(
		.INIT('h153f)
	) name3615 (
		\a[26] ,
		\a[27] ,
		\a[31] ,
		\a[32] ,
		_w3681_
	);
	LUT4 #(
		.INIT('h8000)
	) name3616 (
		\a[26] ,
		\a[27] ,
		\a[31] ,
		\a[32] ,
		_w3682_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3617 (
		\a[26] ,
		\a[27] ,
		\a[31] ,
		\a[32] ,
		_w3683_
	);
	LUT2 #(
		.INIT('h6)
	) name3618 (
		_w3680_,
		_w3683_,
		_w3684_
	);
	LUT4 #(
		.INIT('h0660)
	) name3619 (
		_w3662_,
		_w3667_,
		_w3679_,
		_w3684_,
		_w3685_
	);
	LUT4 #(
		.INIT('h6996)
	) name3620 (
		_w3662_,
		_w3667_,
		_w3679_,
		_w3684_,
		_w3686_
	);
	LUT4 #(
		.INIT('he800)
	) name3621 (
		_w3471_,
		_w3472_,
		_w3473_,
		_w3686_,
		_w3687_
	);
	LUT4 #(
		.INIT('h17e8)
	) name3622 (
		_w3471_,
		_w3472_,
		_w3473_,
		_w3686_,
		_w3688_
	);
	LUT4 #(
		.INIT('h1700)
	) name3623 (
		_w3561_,
		_w3571_,
		_w3572_,
		_w3651_,
		_w3689_
	);
	LUT4 #(
		.INIT('hf616)
	) name3624 (
		_w3629_,
		_w3651_,
		_w3688_,
		_w3689_,
		_w3690_
	);
	LUT3 #(
		.INIT('h69)
	) name3625 (
		_w3607_,
		_w3628_,
		_w3690_,
		_w3691_
	);
	LUT4 #(
		.INIT('hd200)
	) name3626 (
		_w3552_,
		_w3589_,
		_w3606_,
		_w3691_,
		_w3692_
	);
	LUT4 #(
		.INIT('h002d)
	) name3627 (
		_w3552_,
		_w3589_,
		_w3606_,
		_w3691_,
		_w3693_
	);
	LUT4 #(
		.INIT('h2dd2)
	) name3628 (
		_w3552_,
		_w3589_,
		_w3606_,
		_w3691_,
		_w3694_
	);
	LUT3 #(
		.INIT('h0e)
	) name3629 (
		_w3586_,
		_w3587_,
		_w3694_,
		_w3695_
	);
	LUT4 #(
		.INIT('h0001)
	) name3630 (
		_w3586_,
		_w3587_,
		_w3692_,
		_w3693_,
		_w3696_
	);
	LUT3 #(
		.INIT('h56)
	) name3631 (
		_w3582_,
		_w3695_,
		_w3696_,
		_w3697_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3632 (
		_w3352_,
		_w3468_,
		_w3585_,
		_w3697_,
		_w3698_
	);
	LUT3 #(
		.INIT('h03)
	) name3633 (
		_w3582_,
		_w3695_,
		_w3696_,
		_w3699_
	);
	LUT4 #(
		.INIT('hb000)
	) name3634 (
		_w3352_,
		_w3468_,
		_w3585_,
		_w3699_,
		_w3700_
	);
	LUT2 #(
		.INIT('he)
	) name3635 (
		_w3698_,
		_w3700_,
		_w3701_
	);
	LUT4 #(
		.INIT('h040f)
	) name3636 (
		_w3352_,
		_w3468_,
		_w3582_,
		_w3585_,
		_w3702_
	);
	LUT4 #(
		.INIT('h8e00)
	) name3637 (
		_w3559_,
		_w3560_,
		_w3573_,
		_w3628_,
		_w3703_
	);
	LUT4 #(
		.INIT('hff8e)
	) name3638 (
		_w3559_,
		_w3560_,
		_w3573_,
		_w3628_,
		_w3704_
	);
	LUT4 #(
		.INIT('h0071)
	) name3639 (
		_w3559_,
		_w3560_,
		_w3573_,
		_w3628_,
		_w3705_
	);
	LUT3 #(
		.INIT('h0e)
	) name3640 (
		_w3690_,
		_w3703_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('h011f)
	) name3641 (
		_w3522_,
		_w3524_,
		_w3617_,
		_w3627_,
		_w3707_
	);
	LUT2 #(
		.INIT('h2)
	) name3642 (
		_w3645_,
		_w3649_,
		_w3708_
	);
	LUT2 #(
		.INIT('h8)
	) name3643 (
		_w3645_,
		_w3649_,
		_w3709_
	);
	LUT4 #(
		.INIT('he800)
	) name3644 (
		_w3562_,
		_w3566_,
		_w3570_,
		_w3649_,
		_w3710_
	);
	LUT4 #(
		.INIT('h0027)
	) name3645 (
		_w3630_,
		_w3708_,
		_w3709_,
		_w3710_,
		_w3711_
	);
	LUT3 #(
		.INIT('h71)
	) name3646 (
		_w3646_,
		_w3647_,
		_w3648_,
		_w3712_
	);
	LUT3 #(
		.INIT('h17)
	) name3647 (
		_w3622_,
		_w3623_,
		_w3624_,
		_w3713_
	);
	LUT3 #(
		.INIT('h17)
	) name3648 (
		_w3618_,
		_w3619_,
		_w3620_,
		_w3714_
	);
	LUT3 #(
		.INIT('h96)
	) name3649 (
		_w3712_,
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT3 #(
		.INIT('h71)
	) name3650 (
		_w3621_,
		_w3625_,
		_w3626_,
		_w3716_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		_w3715_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h1)
	) name3652 (
		_w3715_,
		_w3716_,
		_w3718_
	);
	LUT2 #(
		.INIT('h6)
	) name3653 (
		_w3715_,
		_w3716_,
		_w3719_
	);
	LUT3 #(
		.INIT('h41)
	) name3654 (
		_w3707_,
		_w3711_,
		_w3719_,
		_w3720_
	);
	LUT3 #(
		.INIT('h96)
	) name3655 (
		_w3707_,
		_w3711_,
		_w3719_,
		_w3721_
	);
	LUT4 #(
		.INIT('hae00)
	) name3656 (
		_w3652_,
		_w3688_,
		_w3689_,
		_w3721_,
		_w3722_
	);
	LUT4 #(
		.INIT('h51ae)
	) name3657 (
		_w3652_,
		_w3688_,
		_w3689_,
		_w3721_,
		_w3723_
	);
	LUT4 #(
		.INIT('hec00)
	) name3658 (
		_w3690_,
		_w3703_,
		_w3704_,
		_w3723_,
		_w3724_
	);
	LUT4 #(
		.INIT('h0013)
	) name3659 (
		_w3690_,
		_w3703_,
		_w3704_,
		_w3723_,
		_w3725_
	);
	LUT3 #(
		.INIT('h32)
	) name3660 (
		_w3601_,
		_w3602_,
		_w3604_,
		_w3726_
	);
	LUT3 #(
		.INIT('h32)
	) name3661 (
		_w3394_,
		_w3657_,
		_w3658_,
		_w3727_
	);
	LUT3 #(
		.INIT('h32)
	) name3662 (
		_w3640_,
		_w3641_,
		_w3642_,
		_w3728_
	);
	LUT3 #(
		.INIT('h0d)
	) name3663 (
		_w3663_,
		_w3664_,
		_w3665_,
		_w3729_
	);
	LUT3 #(
		.INIT('h96)
	) name3664 (
		_w3727_,
		_w3728_,
		_w3729_,
		_w3730_
	);
	LUT3 #(
		.INIT('h0d)
	) name3665 (
		_w3653_,
		_w3654_,
		_w3655_,
		_w3731_
	);
	LUT3 #(
		.INIT('h0d)
	) name3666 (
		_w3673_,
		_w3674_,
		_w3675_,
		_w3732_
	);
	LUT3 #(
		.INIT('h0d)
	) name3667 (
		_w3668_,
		_w3669_,
		_w3671_,
		_w3733_
	);
	LUT3 #(
		.INIT('h96)
	) name3668 (
		_w3731_,
		_w3732_,
		_w3733_,
		_w3734_
	);
	LUT3 #(
		.INIT('h80)
	) name3669 (
		\a[1] ,
		\a[30] ,
		\a[58] ,
		_w3735_
	);
	LUT3 #(
		.INIT('h6c)
	) name3670 (
		\a[1] ,
		\a[30] ,
		\a[58] ,
		_w3736_
	);
	LUT4 #(
		.INIT('h000d)
	) name3671 (
		_w3021_,
		_w3634_,
		_w3635_,
		_w3736_,
		_w3737_
	);
	LUT4 #(
		.INIT('hf200)
	) name3672 (
		_w3021_,
		_w3634_,
		_w3635_,
		_w3736_,
		_w3738_
	);
	LUT4 #(
		.INIT('h0df2)
	) name3673 (
		_w3021_,
		_w3634_,
		_w3635_,
		_w3736_,
		_w3739_
	);
	LUT3 #(
		.INIT('h0d)
	) name3674 (
		_w3502_,
		_w3631_,
		_w3632_,
		_w3740_
	);
	LUT2 #(
		.INIT('h6)
	) name3675 (
		_w3739_,
		_w3740_,
		_w3741_
	);
	LUT3 #(
		.INIT('h69)
	) name3676 (
		_w3730_,
		_w3734_,
		_w3741_,
		_w3742_
	);
	LUT3 #(
		.INIT('h32)
	) name3677 (
		_w3677_,
		_w3678_,
		_w3684_,
		_w3743_
	);
	LUT3 #(
		.INIT('h32)
	) name3678 (
		_w3637_,
		_w3638_,
		_w3644_,
		_w3744_
	);
	LUT3 #(
		.INIT('h32)
	) name3679 (
		_w3660_,
		_w3661_,
		_w3667_,
		_w3745_
	);
	LUT3 #(
		.INIT('h96)
	) name3680 (
		_w3743_,
		_w3744_,
		_w3745_,
		_w3746_
	);
	LUT4 #(
		.INIT('he11e)
	) name3681 (
		_w3685_,
		_w3687_,
		_w3742_,
		_w3746_,
		_w3747_
	);
	LUT4 #(
		.INIT('h8e00)
	) name3682 (
		_w3590_,
		_w3600_,
		_w3604_,
		_w3747_,
		_w3748_
	);
	LUT3 #(
		.INIT('h0e)
	) name3683 (
		_w3591_,
		_w3597_,
		_w3598_,
		_w3749_
	);
	LUT3 #(
		.INIT('hd4)
	) name3684 (
		_w3614_,
		_w3615_,
		_w3616_,
		_w3750_
	);
	LUT4 #(
		.INIT('h153f)
	) name3685 (
		\a[2] ,
		\a[3] ,
		\a[56] ,
		\a[57] ,
		_w3751_
	);
	LUT4 #(
		.INIT('h8000)
	) name3686 (
		\a[2] ,
		\a[3] ,
		\a[56] ,
		\a[57] ,
		_w3752_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3687 (
		\a[2] ,
		\a[3] ,
		\a[56] ,
		\a[57] ,
		_w3753_
	);
	LUT2 #(
		.INIT('h6)
	) name3688 (
		_w3608_,
		_w3753_,
		_w3754_
	);
	LUT3 #(
		.INIT('h0d)
	) name3689 (
		_w3680_,
		_w3681_,
		_w3682_,
		_w3755_
	);
	LUT4 #(
		.INIT('h153f)
	) name3690 (
		\a[5] ,
		\a[19] ,
		\a[40] ,
		\a[54] ,
		_w3756_
	);
	LUT4 #(
		.INIT('h8000)
	) name3691 (
		\a[5] ,
		\a[19] ,
		\a[40] ,
		\a[54] ,
		_w3757_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3692 (
		\a[5] ,
		\a[19] ,
		\a[40] ,
		\a[54] ,
		_w3758_
	);
	LUT2 #(
		.INIT('h6)
	) name3693 (
		_w3490_,
		_w3758_,
		_w3759_
	);
	LUT3 #(
		.INIT('h69)
	) name3694 (
		_w3754_,
		_w3755_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('h8)
	) name3695 (
		\a[11] ,
		\a[48] ,
		_w3761_
	);
	LUT4 #(
		.INIT('h153f)
	) name3696 (
		\a[12] ,
		\a[14] ,
		\a[45] ,
		\a[47] ,
		_w3762_
	);
	LUT4 #(
		.INIT('h8000)
	) name3697 (
		\a[12] ,
		\a[14] ,
		\a[45] ,
		\a[47] ,
		_w3763_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3698 (
		\a[12] ,
		\a[14] ,
		\a[45] ,
		\a[47] ,
		_w3764_
	);
	LUT4 #(
		.INIT('h153f)
	) name3699 (
		\a[28] ,
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w3765_
	);
	LUT4 #(
		.INIT('h8000)
	) name3700 (
		\a[28] ,
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w3766_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3701 (
		\a[28] ,
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w3767_
	);
	LUT4 #(
		.INIT('h1428)
	) name3702 (
		_w3507_,
		_w3761_,
		_w3764_,
		_w3767_,
		_w3768_
	);
	LUT4 #(
		.INIT('h8241)
	) name3703 (
		_w3507_,
		_w3761_,
		_w3764_,
		_w3767_,
		_w3769_
	);
	LUT4 #(
		.INIT('h6996)
	) name3704 (
		_w3507_,
		_w3761_,
		_w3764_,
		_w3767_,
		_w3770_
	);
	LUT4 #(
		.INIT('h153f)
	) name3705 (
		\a[16] ,
		\a[17] ,
		\a[42] ,
		\a[43] ,
		_w3771_
	);
	LUT2 #(
		.INIT('h8)
	) name3706 (
		\a[17] ,
		\a[43] ,
		_w3772_
	);
	LUT4 #(
		.INIT('h8000)
	) name3707 (
		\a[16] ,
		\a[17] ,
		\a[42] ,
		\a[43] ,
		_w3773_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3708 (
		\a[16] ,
		\a[17] ,
		\a[42] ,
		\a[43] ,
		_w3774_
	);
	LUT2 #(
		.INIT('h6)
	) name3709 (
		_w3670_,
		_w3774_,
		_w3775_
	);
	LUT2 #(
		.INIT('h6)
	) name3710 (
		_w3770_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h1)
	) name3711 (
		_w3760_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h8)
	) name3712 (
		_w3760_,
		_w3776_,
		_w3778_
	);
	LUT2 #(
		.INIT('h6)
	) name3713 (
		_w3760_,
		_w3776_,
		_w3779_
	);
	LUT2 #(
		.INIT('h6)
	) name3714 (
		_w3750_,
		_w3779_,
		_w3780_
	);
	LUT3 #(
		.INIT('he8)
	) name3715 (
		_w3592_,
		_w3593_,
		_w3594_,
		_w3781_
	);
	LUT2 #(
		.INIT('h8)
	) name3716 (
		\a[6] ,
		\a[53] ,
		_w3782_
	);
	LUT4 #(
		.INIT('h153f)
	) name3717 (
		\a[7] ,
		\a[18] ,
		\a[41] ,
		\a[52] ,
		_w3783_
	);
	LUT2 #(
		.INIT('h8)
	) name3718 (
		\a[18] ,
		\a[52] ,
		_w3784_
	);
	LUT4 #(
		.INIT('h8000)
	) name3719 (
		\a[7] ,
		\a[18] ,
		\a[41] ,
		\a[52] ,
		_w3785_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3720 (
		\a[7] ,
		\a[18] ,
		\a[41] ,
		\a[52] ,
		_w3786_
	);
	LUT2 #(
		.INIT('h8)
	) name3721 (
		\a[9] ,
		\a[50] ,
		_w3787_
	);
	LUT4 #(
		.INIT('h153f)
	) name3722 (
		\a[10] ,
		\a[15] ,
		\a[44] ,
		\a[49] ,
		_w3788_
	);
	LUT4 #(
		.INIT('h8000)
	) name3723 (
		\a[10] ,
		\a[15] ,
		\a[44] ,
		\a[49] ,
		_w3789_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3724 (
		\a[10] ,
		\a[15] ,
		\a[44] ,
		\a[49] ,
		_w3790_
	);
	LUT4 #(
		.INIT('h0660)
	) name3725 (
		_w3782_,
		_w3786_,
		_w3787_,
		_w3790_,
		_w3791_
	);
	LUT4 #(
		.INIT('h9009)
	) name3726 (
		_w3782_,
		_w3786_,
		_w3787_,
		_w3790_,
		_w3792_
	);
	LUT4 #(
		.INIT('h6996)
	) name3727 (
		_w3782_,
		_w3786_,
		_w3787_,
		_w3790_,
		_w3793_
	);
	LUT4 #(
		.INIT('hba45)
	) name3728 (
		_w3610_,
		_w3611_,
		_w3613_,
		_w3793_,
		_w3794_
	);
	LUT2 #(
		.INIT('h8)
	) name3729 (
		\a[20] ,
		\a[39] ,
		_w3795_
	);
	LUT4 #(
		.INIT('h153f)
	) name3730 (
		\a[21] ,
		\a[22] ,
		\a[37] ,
		\a[38] ,
		_w3796_
	);
	LUT4 #(
		.INIT('h8000)
	) name3731 (
		\a[21] ,
		\a[22] ,
		\a[37] ,
		\a[38] ,
		_w3797_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3732 (
		\a[21] ,
		\a[22] ,
		\a[37] ,
		\a[38] ,
		_w3798_
	);
	LUT2 #(
		.INIT('h8)
	) name3733 (
		\a[23] ,
		\a[36] ,
		_w3799_
	);
	LUT4 #(
		.INIT('h153f)
	) name3734 (
		\a[24] ,
		\a[25] ,
		\a[34] ,
		\a[35] ,
		_w3800_
	);
	LUT4 #(
		.INIT('h8000)
	) name3735 (
		\a[24] ,
		\a[25] ,
		\a[34] ,
		\a[35] ,
		_w3801_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3736 (
		\a[24] ,
		\a[25] ,
		\a[34] ,
		\a[35] ,
		_w3802_
	);
	LUT4 #(
		.INIT('h0660)
	) name3737 (
		_w3795_,
		_w3798_,
		_w3799_,
		_w3802_,
		_w3803_
	);
	LUT4 #(
		.INIT('h9009)
	) name3738 (
		_w3795_,
		_w3798_,
		_w3799_,
		_w3802_,
		_w3804_
	);
	LUT4 #(
		.INIT('h6996)
	) name3739 (
		_w3795_,
		_w3798_,
		_w3799_,
		_w3802_,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name3740 (
		\a[26] ,
		\a[33] ,
		_w3806_
	);
	LUT4 #(
		.INIT('h153f)
	) name3741 (
		\a[0] ,
		\a[27] ,
		\a[32] ,
		\a[59] ,
		_w3807_
	);
	LUT4 #(
		.INIT('h8000)
	) name3742 (
		\a[0] ,
		\a[27] ,
		\a[32] ,
		\a[59] ,
		_w3808_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3743 (
		\a[0] ,
		\a[27] ,
		\a[32] ,
		\a[59] ,
		_w3809_
	);
	LUT2 #(
		.INIT('h6)
	) name3744 (
		_w3806_,
		_w3809_,
		_w3810_
	);
	LUT2 #(
		.INIT('h6)
	) name3745 (
		_w3805_,
		_w3810_,
		_w3811_
	);
	LUT3 #(
		.INIT('h96)
	) name3746 (
		_w3781_,
		_w3794_,
		_w3811_,
		_w3812_
	);
	LUT3 #(
		.INIT('h96)
	) name3747 (
		_w3749_,
		_w3780_,
		_w3812_,
		_w3813_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3748 (
		_w3590_,
		_w3591_,
		_w3599_,
		_w3747_,
		_w3814_
	);
	LUT3 #(
		.INIT('hd0)
	) name3749 (
		_w3603_,
		_w3604_,
		_w3814_,
		_w3815_
	);
	LUT4 #(
		.INIT('h1441)
	) name3750 (
		_w3747_,
		_w3749_,
		_w3780_,
		_w3812_,
		_w3816_
	);
	LUT4 #(
		.INIT('hf949)
	) name3751 (
		_w3726_,
		_w3747_,
		_w3813_,
		_w3815_,
		_w3817_
	);
	LUT3 #(
		.INIT('h96)
	) name3752 (
		_w3706_,
		_w3723_,
		_w3817_,
		_w3818_
	);
	LUT4 #(
		.INIT('h2f02)
	) name3753 (
		_w3552_,
		_w3589_,
		_w3606_,
		_w3691_,
		_w3819_
	);
	LUT2 #(
		.INIT('h4)
	) name3754 (
		_w3818_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h9)
	) name3755 (
		_w3818_,
		_w3819_,
		_w3821_
	);
	LUT2 #(
		.INIT('h4)
	) name3756 (
		_w3695_,
		_w3821_,
		_w3822_
	);
	LUT3 #(
		.INIT('he0)
	) name3757 (
		_w3696_,
		_w3702_,
		_w3822_,
		_w3823_
	);
	LUT2 #(
		.INIT('h4)
	) name3758 (
		_w3695_,
		_w3696_,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name3759 (
		_w3582_,
		_w3695_,
		_w3825_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3760 (
		_w3352_,
		_w3468_,
		_w3585_,
		_w3825_,
		_w3826_
	);
	LUT3 #(
		.INIT('h01)
	) name3761 (
		_w3821_,
		_w3824_,
		_w3826_,
		_w3827_
	);
	LUT2 #(
		.INIT('h1)
	) name3762 (
		_w3823_,
		_w3827_,
		_w3828_
	);
	LUT3 #(
		.INIT('h45)
	) name3763 (
		_w3724_,
		_w3725_,
		_w3817_,
		_w3829_
	);
	LUT4 #(
		.INIT('h011f)
	) name3764 (
		_w3685_,
		_w3687_,
		_w3742_,
		_w3746_,
		_w3830_
	);
	LUT3 #(
		.INIT('h17)
	) name3765 (
		_w3731_,
		_w3732_,
		_w3733_,
		_w3831_
	);
	LUT3 #(
		.INIT('h8e)
	) name3766 (
		_w3727_,
		_w3728_,
		_w3729_,
		_w3832_
	);
	LUT3 #(
		.INIT('hb2)
	) name3767 (
		_w3754_,
		_w3755_,
		_w3759_,
		_w3833_
	);
	LUT3 #(
		.INIT('h96)
	) name3768 (
		_w3831_,
		_w3832_,
		_w3833_,
		_w3834_
	);
	LUT3 #(
		.INIT('he8)
	) name3769 (
		_w3743_,
		_w3744_,
		_w3745_,
		_w3835_
	);
	LUT2 #(
		.INIT('h1)
	) name3770 (
		_w3834_,
		_w3835_,
		_w3836_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		_w3834_,
		_w3835_,
		_w3837_
	);
	LUT2 #(
		.INIT('h6)
	) name3772 (
		_w3834_,
		_w3835_,
		_w3838_
	);
	LUT3 #(
		.INIT('h17)
	) name3773 (
		_w3781_,
		_w3794_,
		_w3811_,
		_w3839_
	);
	LUT3 #(
		.INIT('h41)
	) name3774 (
		_w3830_,
		_w3838_,
		_w3839_,
		_w3840_
	);
	LUT3 #(
		.INIT('h28)
	) name3775 (
		_w3830_,
		_w3838_,
		_w3839_,
		_w3841_
	);
	LUT3 #(
		.INIT('h96)
	) name3776 (
		_w3830_,
		_w3838_,
		_w3839_,
		_w3842_
	);
	LUT4 #(
		.INIT('h17e8)
	) name3777 (
		_w3749_,
		_w3780_,
		_w3812_,
		_w3842_,
		_w3843_
	);
	LUT4 #(
		.INIT('h0051)
	) name3778 (
		_w3748_,
		_w3813_,
		_w3815_,
		_w3843_,
		_w3844_
	);
	LUT4 #(
		.INIT('h1441)
	) name3779 (
		_w3602_,
		_w3749_,
		_w3780_,
		_w3812_,
		_w3845_
	);
	LUT4 #(
		.INIT('h0203)
	) name3780 (
		_w3605_,
		_w3815_,
		_w3816_,
		_w3845_,
		_w3846_
	);
	LUT3 #(
		.INIT('h0d)
	) name3781 (
		_w3750_,
		_w3777_,
		_w3778_,
		_w3847_
	);
	LUT4 #(
		.INIT('h0071)
	) name3782 (
		_w3564_,
		_w3609_,
		_w3613_,
		_w3791_,
		_w3848_
	);
	LUT3 #(
		.INIT('h32)
	) name3783 (
		_w3490_,
		_w3756_,
		_w3757_,
		_w3849_
	);
	LUT3 #(
		.INIT('h0d)
	) name3784 (
		_w3795_,
		_w3796_,
		_w3797_,
		_w3850_
	);
	LUT3 #(
		.INIT('h0d)
	) name3785 (
		_w3799_,
		_w3800_,
		_w3801_,
		_w3851_
	);
	LUT3 #(
		.INIT('h69)
	) name3786 (
		_w3849_,
		_w3850_,
		_w3851_,
		_w3852_
	);
	LUT3 #(
		.INIT('h0d)
	) name3787 (
		_w3806_,
		_w3807_,
		_w3808_,
		_w3853_
	);
	LUT3 #(
		.INIT('h0d)
	) name3788 (
		_w3608_,
		_w3751_,
		_w3752_,
		_w3854_
	);
	LUT3 #(
		.INIT('h0d)
	) name3789 (
		_w3787_,
		_w3788_,
		_w3789_,
		_w3855_
	);
	LUT3 #(
		.INIT('h96)
	) name3790 (
		_w3853_,
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name3791 (
		_w3792_,
		_w3848_,
		_w3852_,
		_w3856_,
		_w3857_
	);
	LUT3 #(
		.INIT('h0d)
	) name3792 (
		_w3670_,
		_w3771_,
		_w3773_,
		_w3858_
	);
	LUT3 #(
		.INIT('h0d)
	) name3793 (
		_w3782_,
		_w3783_,
		_w3785_,
		_w3859_
	);
	LUT3 #(
		.INIT('h32)
	) name3794 (
		_w3507_,
		_w3765_,
		_w3766_,
		_w3860_
	);
	LUT3 #(
		.INIT('h96)
	) name3795 (
		_w3858_,
		_w3859_,
		_w3860_,
		_w3861_
	);
	LUT3 #(
		.INIT('h32)
	) name3796 (
		_w3803_,
		_w3804_,
		_w3810_,
		_w3862_
	);
	LUT3 #(
		.INIT('h32)
	) name3797 (
		_w3768_,
		_w3769_,
		_w3775_,
		_w3863_
	);
	LUT3 #(
		.INIT('h96)
	) name3798 (
		_w3861_,
		_w3862_,
		_w3863_,
		_w3864_
	);
	LUT3 #(
		.INIT('h69)
	) name3799 (
		_w3847_,
		_w3857_,
		_w3864_,
		_w3865_
	);
	LUT3 #(
		.INIT('h32)
	) name3800 (
		_w3711_,
		_w3717_,
		_w3718_,
		_w3866_
	);
	LUT3 #(
		.INIT('he8)
	) name3801 (
		_w3712_,
		_w3713_,
		_w3714_,
		_w3867_
	);
	LUT2 #(
		.INIT('h8)
	) name3802 (
		\a[2] ,
		\a[58] ,
		_w3868_
	);
	LUT4 #(
		.INIT('h153f)
	) name3803 (
		\a[3] ,
		\a[4] ,
		\a[56] ,
		\a[57] ,
		_w3869_
	);
	LUT4 #(
		.INIT('h8000)
	) name3804 (
		\a[3] ,
		\a[4] ,
		\a[56] ,
		\a[57] ,
		_w3870_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3805 (
		\a[3] ,
		\a[4] ,
		\a[56] ,
		\a[57] ,
		_w3871_
	);
	LUT2 #(
		.INIT('h8)
	) name3806 (
		\a[20] ,
		\a[40] ,
		_w3872_
	);
	LUT4 #(
		.INIT('h153f)
	) name3807 (
		\a[21] ,
		\a[22] ,
		\a[38] ,
		\a[39] ,
		_w3873_
	);
	LUT2 #(
		.INIT('h8)
	) name3808 (
		\a[22] ,
		\a[39] ,
		_w3874_
	);
	LUT4 #(
		.INIT('h8000)
	) name3809 (
		\a[21] ,
		\a[22] ,
		\a[38] ,
		\a[39] ,
		_w3875_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3810 (
		\a[21] ,
		\a[22] ,
		\a[38] ,
		\a[39] ,
		_w3876_
	);
	LUT4 #(
		.INIT('h0660)
	) name3811 (
		_w3868_,
		_w3871_,
		_w3872_,
		_w3876_,
		_w3877_
	);
	LUT4 #(
		.INIT('h9009)
	) name3812 (
		_w3868_,
		_w3871_,
		_w3872_,
		_w3876_,
		_w3878_
	);
	LUT4 #(
		.INIT('h6996)
	) name3813 (
		_w3868_,
		_w3871_,
		_w3872_,
		_w3876_,
		_w3879_
	);
	LUT2 #(
		.INIT('h8)
	) name3814 (
		\a[24] ,
		\a[36] ,
		_w3880_
	);
	LUT4 #(
		.INIT('h153f)
	) name3815 (
		\a[25] ,
		\a[26] ,
		\a[34] ,
		\a[35] ,
		_w3881_
	);
	LUT2 #(
		.INIT('h8)
	) name3816 (
		\a[26] ,
		\a[35] ,
		_w3882_
	);
	LUT4 #(
		.INIT('h8000)
	) name3817 (
		\a[25] ,
		\a[26] ,
		\a[34] ,
		\a[35] ,
		_w3883_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3818 (
		\a[25] ,
		\a[26] ,
		\a[34] ,
		\a[35] ,
		_w3884_
	);
	LUT2 #(
		.INIT('h6)
	) name3819 (
		_w3880_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h6)
	) name3820 (
		_w3879_,
		_w3885_,
		_w3886_
	);
	LUT4 #(
		.INIT('h153f)
	) name3821 (
		\a[9] ,
		\a[16] ,
		\a[44] ,
		\a[51] ,
		_w3887_
	);
	LUT4 #(
		.INIT('h8000)
	) name3822 (
		\a[9] ,
		\a[16] ,
		\a[44] ,
		\a[51] ,
		_w3888_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3823 (
		\a[9] ,
		\a[16] ,
		\a[44] ,
		\a[51] ,
		_w3889_
	);
	LUT2 #(
		.INIT('h6)
	) name3824 (
		_w3772_,
		_w3889_,
		_w3890_
	);
	LUT3 #(
		.INIT('h0d)
	) name3825 (
		_w3761_,
		_w3762_,
		_w3763_,
		_w3891_
	);
	LUT2 #(
		.INIT('h8)
	) name3826 (
		\a[10] ,
		\a[50] ,
		_w3892_
	);
	LUT4 #(
		.INIT('h153f)
	) name3827 (
		\a[11] ,
		\a[15] ,
		\a[45] ,
		\a[49] ,
		_w3893_
	);
	LUT4 #(
		.INIT('h8000)
	) name3828 (
		\a[11] ,
		\a[15] ,
		\a[45] ,
		\a[49] ,
		_w3894_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3829 (
		\a[11] ,
		\a[15] ,
		\a[45] ,
		\a[49] ,
		_w3895_
	);
	LUT2 #(
		.INIT('h6)
	) name3830 (
		_w3892_,
		_w3895_,
		_w3896_
	);
	LUT3 #(
		.INIT('h69)
	) name3831 (
		_w3890_,
		_w3891_,
		_w3896_,
		_w3897_
	);
	LUT3 #(
		.INIT('h96)
	) name3832 (
		_w3867_,
		_w3886_,
		_w3897_,
		_w3898_
	);
	LUT4 #(
		.INIT('hd400)
	) name3833 (
		_w3711_,
		_w3715_,
		_w3716_,
		_w3898_,
		_w3899_
	);
	LUT3 #(
		.INIT('h17)
	) name3834 (
		_w3730_,
		_w3734_,
		_w3741_,
		_w3900_
	);
	LUT3 #(
		.INIT('h45)
	) name3835 (
		_w3737_,
		_w3738_,
		_w3740_,
		_w3901_
	);
	LUT4 #(
		.INIT('h8000)
	) name3836 (
		\a[1] ,
		\a[29] ,
		\a[31] ,
		\a[59] ,
		_w3902_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3837 (
		\a[1] ,
		\a[29] ,
		\a[31] ,
		\a[59] ,
		_w3903_
	);
	LUT2 #(
		.INIT('h8)
	) name3838 (
		\a[0] ,
		\a[60] ,
		_w3904_
	);
	LUT3 #(
		.INIT('h96)
	) name3839 (
		_w3735_,
		_w3903_,
		_w3904_,
		_w3905_
	);
	LUT2 #(
		.INIT('h8)
	) name3840 (
		\a[27] ,
		\a[33] ,
		_w3906_
	);
	LUT4 #(
		.INIT('h153f)
	) name3841 (
		\a[23] ,
		\a[28] ,
		\a[32] ,
		\a[37] ,
		_w3907_
	);
	LUT4 #(
		.INIT('h8000)
	) name3842 (
		\a[23] ,
		\a[28] ,
		\a[32] ,
		\a[37] ,
		_w3908_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3843 (
		\a[23] ,
		\a[28] ,
		\a[32] ,
		\a[37] ,
		_w3909_
	);
	LUT2 #(
		.INIT('h6)
	) name3844 (
		_w3906_,
		_w3909_,
		_w3910_
	);
	LUT2 #(
		.INIT('h8)
	) name3845 (
		_w3905_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h1)
	) name3846 (
		_w3905_,
		_w3910_,
		_w3912_
	);
	LUT2 #(
		.INIT('h6)
	) name3847 (
		_w3905_,
		_w3910_,
		_w3913_
	);
	LUT4 #(
		.INIT('h153f)
	) name3848 (
		\a[12] ,
		\a[13] ,
		\a[47] ,
		\a[48] ,
		_w3914_
	);
	LUT2 #(
		.INIT('h8)
	) name3849 (
		\a[13] ,
		\a[48] ,
		_w3915_
	);
	LUT4 #(
		.INIT('h8000)
	) name3850 (
		\a[12] ,
		\a[13] ,
		\a[47] ,
		\a[48] ,
		_w3916_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3851 (
		\a[12] ,
		\a[13] ,
		\a[47] ,
		\a[48] ,
		_w3917_
	);
	LUT2 #(
		.INIT('h8)
	) name3852 (
		\a[7] ,
		\a[53] ,
		_w3918_
	);
	LUT4 #(
		.INIT('h153f)
	) name3853 (
		\a[8] ,
		\a[18] ,
		\a[42] ,
		\a[52] ,
		_w3919_
	);
	LUT4 #(
		.INIT('h8000)
	) name3854 (
		\a[8] ,
		\a[18] ,
		\a[42] ,
		\a[52] ,
		_w3920_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3855 (
		\a[8] ,
		\a[18] ,
		\a[42] ,
		\a[52] ,
		_w3921_
	);
	LUT4 #(
		.INIT('h0660)
	) name3856 (
		_w3386_,
		_w3917_,
		_w3918_,
		_w3921_,
		_w3922_
	);
	LUT4 #(
		.INIT('h9009)
	) name3857 (
		_w3386_,
		_w3917_,
		_w3918_,
		_w3921_,
		_w3923_
	);
	LUT4 #(
		.INIT('h6996)
	) name3858 (
		_w3386_,
		_w3917_,
		_w3918_,
		_w3921_,
		_w3924_
	);
	LUT2 #(
		.INIT('h8)
	) name3859 (
		\a[5] ,
		\a[55] ,
		_w3925_
	);
	LUT4 #(
		.INIT('h153f)
	) name3860 (
		\a[6] ,
		\a[19] ,
		\a[41] ,
		\a[54] ,
		_w3926_
	);
	LUT4 #(
		.INIT('h8000)
	) name3861 (
		\a[6] ,
		\a[19] ,
		\a[41] ,
		\a[54] ,
		_w3927_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3862 (
		\a[6] ,
		\a[19] ,
		\a[41] ,
		\a[54] ,
		_w3928_
	);
	LUT2 #(
		.INIT('h6)
	) name3863 (
		_w3925_,
		_w3928_,
		_w3929_
	);
	LUT2 #(
		.INIT('h6)
	) name3864 (
		_w3924_,
		_w3929_,
		_w3930_
	);
	LUT3 #(
		.INIT('h09)
	) name3865 (
		_w3901_,
		_w3913_,
		_w3930_,
		_w3931_
	);
	LUT3 #(
		.INIT('h60)
	) name3866 (
		_w3901_,
		_w3913_,
		_w3930_,
		_w3932_
	);
	LUT3 #(
		.INIT('h96)
	) name3867 (
		_w3901_,
		_w3913_,
		_w3930_,
		_w3933_
	);
	LUT2 #(
		.INIT('h6)
	) name3868 (
		_w3900_,
		_w3933_,
		_w3934_
	);
	LUT4 #(
		.INIT('h002b)
	) name3869 (
		_w3711_,
		_w3715_,
		_w3716_,
		_w3898_,
		_w3935_
	);
	LUT3 #(
		.INIT('h04)
	) name3870 (
		_w3899_,
		_w3934_,
		_w3935_,
		_w3936_
	);
	LUT4 #(
		.INIT('hf04b)
	) name3871 (
		_w3866_,
		_w3898_,
		_w3934_,
		_w3935_,
		_w3937_
	);
	LUT4 #(
		.INIT('he11e)
	) name3872 (
		_w3720_,
		_w3722_,
		_w3865_,
		_w3937_,
		_w3938_
	);
	LUT4 #(
		.INIT('hec13)
	) name3873 (
		_w3843_,
		_w3844_,
		_w3846_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h2)
	) name3874 (
		_w3829_,
		_w3939_,
		_w3940_
	);
	LUT4 #(
		.INIT('hd00d)
	) name3875 (
		_w3818_,
		_w3819_,
		_w3829_,
		_w3939_,
		_w3941_
	);
	LUT4 #(
		.INIT('hab00)
	) name3876 (
		_w3820_,
		_w3824_,
		_w3826_,
		_w3941_,
		_w3942_
	);
	LUT4 #(
		.INIT('h0220)
	) name3877 (
		_w3818_,
		_w3819_,
		_w3829_,
		_w3939_,
		_w3943_
	);
	LUT4 #(
		.INIT('h0bb0)
	) name3878 (
		_w3818_,
		_w3819_,
		_w3829_,
		_w3939_,
		_w3944_
	);
	LUT4 #(
		.INIT('h010f)
	) name3879 (
		_w3824_,
		_w3826_,
		_w3943_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('hb)
	) name3880 (
		_w3942_,
		_w3945_,
		_w3946_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3881 (
		_w3818_,
		_w3819_,
		_w3829_,
		_w3939_,
		_w3947_
	);
	LUT4 #(
		.INIT('hab00)
	) name3882 (
		_w3820_,
		_w3824_,
		_w3826_,
		_w3947_,
		_w3948_
	);
	LUT4 #(
		.INIT('h0017)
	) name3883 (
		_w3749_,
		_w3780_,
		_w3812_,
		_w3840_,
		_w3949_
	);
	LUT3 #(
		.INIT('h32)
	) name3884 (
		_w3900_,
		_w3931_,
		_w3932_,
		_w3950_
	);
	LUT3 #(
		.INIT('h32)
	) name3885 (
		_w3918_,
		_w3919_,
		_w3920_,
		_w3951_
	);
	LUT3 #(
		.INIT('h0d)
	) name3886 (
		_w3772_,
		_w3887_,
		_w3888_,
		_w3952_
	);
	LUT3 #(
		.INIT('he8)
	) name3887 (
		_w3735_,
		_w3903_,
		_w3904_,
		_w3953_
	);
	LUT3 #(
		.INIT('h69)
	) name3888 (
		_w3951_,
		_w3952_,
		_w3953_,
		_w3954_
	);
	LUT3 #(
		.INIT('h32)
	) name3889 (
		_w3922_,
		_w3923_,
		_w3929_,
		_w3955_
	);
	LUT2 #(
		.INIT('h1)
	) name3890 (
		_w3954_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h8)
	) name3891 (
		_w3954_,
		_w3955_,
		_w3957_
	);
	LUT2 #(
		.INIT('h6)
	) name3892 (
		_w3954_,
		_w3955_,
		_w3958_
	);
	LUT3 #(
		.INIT('h0e)
	) name3893 (
		_w3901_,
		_w3911_,
		_w3912_,
		_w3959_
	);
	LUT3 #(
		.INIT('h32)
	) name3894 (
		_w3906_,
		_w3907_,
		_w3908_,
		_w3960_
	);
	LUT3 #(
		.INIT('h0d)
	) name3895 (
		_w3880_,
		_w3881_,
		_w3883_,
		_w3961_
	);
	LUT3 #(
		.INIT('h0d)
	) name3896 (
		_w3872_,
		_w3873_,
		_w3875_,
		_w3962_
	);
	LUT3 #(
		.INIT('h69)
	) name3897 (
		_w3960_,
		_w3961_,
		_w3962_,
		_w3963_
	);
	LUT3 #(
		.INIT('h32)
	) name3898 (
		_w3925_,
		_w3926_,
		_w3927_,
		_w3964_
	);
	LUT3 #(
		.INIT('h0d)
	) name3899 (
		_w3868_,
		_w3869_,
		_w3870_,
		_w3965_
	);
	LUT3 #(
		.INIT('h0d)
	) name3900 (
		_w3892_,
		_w3893_,
		_w3894_,
		_w3966_
	);
	LUT3 #(
		.INIT('h69)
	) name3901 (
		_w3964_,
		_w3965_,
		_w3966_,
		_w3967_
	);
	LUT3 #(
		.INIT('h32)
	) name3902 (
		_w3877_,
		_w3878_,
		_w3885_,
		_w3968_
	);
	LUT3 #(
		.INIT('h96)
	) name3903 (
		_w3963_,
		_w3967_,
		_w3968_,
		_w3969_
	);
	LUT3 #(
		.INIT('h09)
	) name3904 (
		_w3958_,
		_w3959_,
		_w3969_,
		_w3970_
	);
	LUT3 #(
		.INIT('h60)
	) name3905 (
		_w3958_,
		_w3959_,
		_w3969_,
		_w3971_
	);
	LUT3 #(
		.INIT('h96)
	) name3906 (
		_w3958_,
		_w3959_,
		_w3969_,
		_w3972_
	);
	LUT2 #(
		.INIT('h9)
	) name3907 (
		_w3950_,
		_w3972_,
		_w3973_
	);
	LUT3 #(
		.INIT('h2b)
	) name3908 (
		_w3847_,
		_w3857_,
		_w3864_,
		_w3974_
	);
	LUT3 #(
		.INIT('he8)
	) name3909 (
		_w3831_,
		_w3832_,
		_w3833_,
		_w3975_
	);
	LUT2 #(
		.INIT('h8)
	) name3910 (
		\a[11] ,
		\a[50] ,
		_w3976_
	);
	LUT4 #(
		.INIT('h153f)
	) name3911 (
		\a[12] ,
		\a[14] ,
		\a[47] ,
		\a[49] ,
		_w3977_
	);
	LUT2 #(
		.INIT('h8)
	) name3912 (
		\a[14] ,
		\a[49] ,
		_w3978_
	);
	LUT4 #(
		.INIT('h8000)
	) name3913 (
		\a[12] ,
		\a[14] ,
		\a[47] ,
		\a[49] ,
		_w3979_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3914 (
		\a[12] ,
		\a[14] ,
		\a[47] ,
		\a[49] ,
		_w3980_
	);
	LUT2 #(
		.INIT('h8)
	) name3915 (
		\a[16] ,
		\a[45] ,
		_w3981_
	);
	LUT4 #(
		.INIT('h153f)
	) name3916 (
		\a[10] ,
		\a[15] ,
		\a[46] ,
		\a[51] ,
		_w3982_
	);
	LUT4 #(
		.INIT('h8000)
	) name3917 (
		\a[10] ,
		\a[15] ,
		\a[46] ,
		\a[51] ,
		_w3983_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3918 (
		\a[10] ,
		\a[15] ,
		\a[46] ,
		\a[51] ,
		_w3984_
	);
	LUT4 #(
		.INIT('h0660)
	) name3919 (
		_w3976_,
		_w3980_,
		_w3981_,
		_w3984_,
		_w3985_
	);
	LUT4 #(
		.INIT('h9009)
	) name3920 (
		_w3976_,
		_w3980_,
		_w3981_,
		_w3984_,
		_w3986_
	);
	LUT4 #(
		.INIT('h6996)
	) name3921 (
		_w3976_,
		_w3980_,
		_w3981_,
		_w3984_,
		_w3987_
	);
	LUT4 #(
		.INIT('h153f)
	) name3922 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		\a[32] ,
		_w3988_
	);
	LUT4 #(
		.INIT('h8000)
	) name3923 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		\a[32] ,
		_w3989_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3924 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		\a[32] ,
		_w3990_
	);
	LUT2 #(
		.INIT('h6)
	) name3925 (
		_w3915_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h6)
	) name3926 (
		_w3987_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h8)
	) name3927 (
		\a[0] ,
		\a[61] ,
		_w3993_
	);
	LUT4 #(
		.INIT('h153f)
	) name3928 (
		\a[2] ,
		\a[5] ,
		\a[56] ,
		\a[59] ,
		_w3994_
	);
	LUT2 #(
		.INIT('h8)
	) name3929 (
		\a[5] ,
		\a[59] ,
		_w3995_
	);
	LUT4 #(
		.INIT('h8000)
	) name3930 (
		\a[2] ,
		\a[5] ,
		\a[56] ,
		\a[59] ,
		_w3996_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3931 (
		\a[2] ,
		\a[5] ,
		\a[56] ,
		\a[59] ,
		_w3997_
	);
	LUT2 #(
		.INIT('h8)
	) name3932 (
		\a[6] ,
		\a[55] ,
		_w3998_
	);
	LUT4 #(
		.INIT('h153f)
	) name3933 (
		\a[20] ,
		\a[21] ,
		\a[40] ,
		\a[41] ,
		_w3999_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		\a[21] ,
		\a[41] ,
		_w4000_
	);
	LUT4 #(
		.INIT('h8000)
	) name3935 (
		\a[20] ,
		\a[21] ,
		\a[40] ,
		\a[41] ,
		_w4001_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3936 (
		\a[20] ,
		\a[21] ,
		\a[40] ,
		\a[41] ,
		_w4002_
	);
	LUT4 #(
		.INIT('h0660)
	) name3937 (
		_w3993_,
		_w3997_,
		_w3998_,
		_w4002_,
		_w4003_
	);
	LUT4 #(
		.INIT('h9009)
	) name3938 (
		_w3993_,
		_w3997_,
		_w3998_,
		_w4002_,
		_w4004_
	);
	LUT4 #(
		.INIT('h6996)
	) name3939 (
		_w3993_,
		_w3997_,
		_w3998_,
		_w4002_,
		_w4005_
	);
	LUT4 #(
		.INIT('h153f)
	) name3940 (
		\a[24] ,
		\a[25] ,
		\a[36] ,
		\a[37] ,
		_w4006_
	);
	LUT4 #(
		.INIT('h8000)
	) name3941 (
		\a[24] ,
		\a[25] ,
		\a[36] ,
		\a[37] ,
		_w4007_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3942 (
		\a[24] ,
		\a[25] ,
		\a[36] ,
		\a[37] ,
		_w4008_
	);
	LUT2 #(
		.INIT('h6)
	) name3943 (
		_w3874_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h6)
	) name3944 (
		_w4005_,
		_w4009_,
		_w4010_
	);
	LUT4 #(
		.INIT('h0990)
	) name3945 (
		_w3987_,
		_w3991_,
		_w4005_,
		_w4009_,
		_w4011_
	);
	LUT4 #(
		.INIT('he800)
	) name3946 (
		_w3831_,
		_w3832_,
		_w3833_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('h0660)
	) name3947 (
		_w3987_,
		_w3991_,
		_w4005_,
		_w4009_,
		_w4013_
	);
	LUT4 #(
		.INIT('h1700)
	) name3948 (
		_w3831_,
		_w3832_,
		_w3833_,
		_w4013_,
		_w4014_
	);
	LUT3 #(
		.INIT('h96)
	) name3949 (
		_w3975_,
		_w3992_,
		_w4010_,
		_w4015_
	);
	LUT4 #(
		.INIT('h8e00)
	) name3950 (
		_w3834_,
		_w3835_,
		_w3839_,
		_w4015_,
		_w4016_
	);
	LUT4 #(
		.INIT('h0071)
	) name3951 (
		_w3834_,
		_w3835_,
		_w3839_,
		_w4015_,
		_w4017_
	);
	LUT4 #(
		.INIT('h32cd)
	) name3952 (
		_w3836_,
		_w3837_,
		_w3839_,
		_w4015_,
		_w4018_
	);
	LUT2 #(
		.INIT('h9)
	) name3953 (
		_w3974_,
		_w4018_,
		_w4019_
	);
	LUT4 #(
		.INIT('he11e)
	) name3954 (
		_w3841_,
		_w3949_,
		_w3973_,
		_w4019_,
		_w4020_
	);
	LUT4 #(
		.INIT('hfee0)
	) name3955 (
		_w3720_,
		_w3722_,
		_w3865_,
		_w3937_,
		_w4021_
	);
	LUT3 #(
		.INIT('h51)
	) name3956 (
		_w3899_,
		_w3934_,
		_w3935_,
		_w4022_
	);
	LUT3 #(
		.INIT('h17)
	) name3957 (
		_w3867_,
		_w3886_,
		_w3897_,
		_w4023_
	);
	LUT3 #(
		.INIT('hb2)
	) name3958 (
		_w3890_,
		_w3891_,
		_w3896_,
		_w4024_
	);
	LUT3 #(
		.INIT('h2b)
	) name3959 (
		_w3849_,
		_w3850_,
		_w3851_,
		_w4025_
	);
	LUT2 #(
		.INIT('h8)
	) name3960 (
		\a[1] ,
		\a[60] ,
		_w4026_
	);
	LUT3 #(
		.INIT('h2d)
	) name3961 (
		\a[31] ,
		_w3902_,
		_w4026_,
		_w4027_
	);
	LUT3 #(
		.INIT('h0d)
	) name3962 (
		_w3386_,
		_w3914_,
		_w3916_,
		_w4028_
	);
	LUT2 #(
		.INIT('h6)
	) name3963 (
		_w4027_,
		_w4028_,
		_w4029_
	);
	LUT3 #(
		.INIT('h96)
	) name3964 (
		_w4024_,
		_w4025_,
		_w4029_,
		_w4030_
	);
	LUT2 #(
		.INIT('h8)
	) name3965 (
		\a[23] ,
		\a[38] ,
		_w4031_
	);
	LUT4 #(
		.INIT('h153f)
	) name3966 (
		\a[3] ,
		\a[4] ,
		\a[57] ,
		\a[58] ,
		_w4032_
	);
	LUT4 #(
		.INIT('h8000)
	) name3967 (
		\a[3] ,
		\a[4] ,
		\a[57] ,
		\a[58] ,
		_w4033_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3968 (
		\a[3] ,
		\a[4] ,
		\a[57] ,
		\a[58] ,
		_w4034_
	);
	LUT2 #(
		.INIT('h6)
	) name3969 (
		_w4031_,
		_w4034_,
		_w4035_
	);
	LUT4 #(
		.INIT('h008e)
	) name3970 (
		_w3858_,
		_w3859_,
		_w3860_,
		_w4035_,
		_w4036_
	);
	LUT3 #(
		.INIT('h17)
	) name3971 (
		_w3853_,
		_w3854_,
		_w3855_,
		_w4037_
	);
	LUT4 #(
		.INIT('h7100)
	) name3972 (
		_w3858_,
		_w3859_,
		_w3860_,
		_w4035_,
		_w4038_
	);
	LUT3 #(
		.INIT('hc9)
	) name3973 (
		_w4036_,
		_w4037_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h6)
	) name3974 (
		_w4030_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h9)
	) name3975 (
		_w4023_,
		_w4040_,
		_w4041_
	);
	LUT4 #(
		.INIT('heee0)
	) name3976 (
		_w3792_,
		_w3848_,
		_w3852_,
		_w3856_,
		_w4042_
	);
	LUT4 #(
		.INIT('h011f)
	) name3977 (
		_w3792_,
		_w3848_,
		_w3852_,
		_w3856_,
		_w4043_
	);
	LUT2 #(
		.INIT('h8)
	) name3978 (
		\a[19] ,
		\a[42] ,
		_w4044_
	);
	LUT4 #(
		.INIT('h153f)
	) name3979 (
		\a[7] ,
		\a[8] ,
		\a[53] ,
		\a[54] ,
		_w4045_
	);
	LUT4 #(
		.INIT('h8000)
	) name3980 (
		\a[7] ,
		\a[8] ,
		\a[53] ,
		\a[54] ,
		_w4046_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3981 (
		\a[7] ,
		\a[8] ,
		\a[53] ,
		\a[54] ,
		_w4047_
	);
	LUT2 #(
		.INIT('h8)
	) name3982 (
		\a[18] ,
		\a[43] ,
		_w4048_
	);
	LUT4 #(
		.INIT('h153f)
	) name3983 (
		\a[9] ,
		\a[17] ,
		\a[44] ,
		\a[52] ,
		_w4049_
	);
	LUT4 #(
		.INIT('h8000)
	) name3984 (
		\a[9] ,
		\a[17] ,
		\a[44] ,
		\a[52] ,
		_w4050_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3985 (
		\a[9] ,
		\a[17] ,
		\a[44] ,
		\a[52] ,
		_w4051_
	);
	LUT4 #(
		.INIT('h0660)
	) name3986 (
		_w4044_,
		_w4047_,
		_w4048_,
		_w4051_,
		_w4052_
	);
	LUT4 #(
		.INIT('h9009)
	) name3987 (
		_w4044_,
		_w4047_,
		_w4048_,
		_w4051_,
		_w4053_
	);
	LUT4 #(
		.INIT('h6996)
	) name3988 (
		_w4044_,
		_w4047_,
		_w4048_,
		_w4051_,
		_w4054_
	);
	LUT4 #(
		.INIT('h153f)
	) name3989 (
		\a[27] ,
		\a[28] ,
		\a[33] ,
		\a[34] ,
		_w4055_
	);
	LUT4 #(
		.INIT('h8000)
	) name3990 (
		\a[27] ,
		\a[28] ,
		\a[33] ,
		\a[34] ,
		_w4056_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name3991 (
		\a[27] ,
		\a[28] ,
		\a[33] ,
		\a[34] ,
		_w4057_
	);
	LUT2 #(
		.INIT('h6)
	) name3992 (
		_w3882_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h6)
	) name3993 (
		_w4054_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h1)
	) name3994 (
		_w4043_,
		_w4059_,
		_w4060_
	);
	LUT3 #(
		.INIT('he8)
	) name3995 (
		_w3861_,
		_w3862_,
		_w3863_,
		_w4061_
	);
	LUT3 #(
		.INIT('h70)
	) name3996 (
		_w3852_,
		_w3856_,
		_w4059_,
		_w4062_
	);
	LUT2 #(
		.INIT('h4)
	) name3997 (
		_w4042_,
		_w4062_,
		_w4063_
	);
	LUT3 #(
		.INIT('hc9)
	) name3998 (
		_w4060_,
		_w4061_,
		_w4063_,
		_w4064_
	);
	LUT2 #(
		.INIT('h1)
	) name3999 (
		_w4041_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h6)
	) name4000 (
		_w4041_,
		_w4064_,
		_w4066_
	);
	LUT2 #(
		.INIT('h9)
	) name4001 (
		_w4022_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h6)
	) name4002 (
		_w4021_,
		_w4067_,
		_w4068_
	);
	LUT3 #(
		.INIT('h41)
	) name4003 (
		_w4020_,
		_w4021_,
		_w4067_,
		_w4069_
	);
	LUT4 #(
		.INIT('h3320)
	) name4004 (
		_w3843_,
		_w3844_,
		_w3846_,
		_w3938_,
		_w4070_
	);
	LUT3 #(
		.INIT('h28)
	) name4005 (
		_w4020_,
		_w4021_,
		_w4067_,
		_w4071_
	);
	LUT3 #(
		.INIT('h04)
	) name4006 (
		_w4069_,
		_w4070_,
		_w4071_,
		_w4072_
	);
	LUT3 #(
		.INIT('h96)
	) name4007 (
		_w4020_,
		_w4021_,
		_w4067_,
		_w4073_
	);
	LUT2 #(
		.INIT('h1)
	) name4008 (
		_w4070_,
		_w4073_,
		_w4074_
	);
	LUT3 #(
		.INIT('h96)
	) name4009 (
		_w4020_,
		_w4068_,
		_w4070_,
		_w4075_
	);
	LUT3 #(
		.INIT('he1)
	) name4010 (
		_w3940_,
		_w3948_,
		_w4075_,
		_w4076_
	);
	LUT2 #(
		.INIT('h2)
	) name4011 (
		_w3947_,
		_w4072_,
		_w4077_
	);
	LUT4 #(
		.INIT('hab00)
	) name4012 (
		_w3820_,
		_w3824_,
		_w3826_,
		_w4077_,
		_w4078_
	);
	LUT3 #(
		.INIT('he8)
	) name4013 (
		_w4020_,
		_w4021_,
		_w4067_,
		_w4079_
	);
	LUT3 #(
		.INIT('h15)
	) name4014 (
		_w3899_,
		_w4041_,
		_w4064_,
		_w4080_
	);
	LUT3 #(
		.INIT('hb2)
	) name4015 (
		_w3951_,
		_w3952_,
		_w3953_,
		_w4081_
	);
	LUT2 #(
		.INIT('h4)
	) name4016 (
		\a[60] ,
		_w3902_,
		_w4082_
	);
	LUT4 #(
		.INIT('h5093)
	) name4017 (
		\a[1] ,
		\a[31] ,
		\a[60] ,
		_w3902_,
		_w4083_
	);
	LUT3 #(
		.INIT('h0d)
	) name4018 (
		_w4028_,
		_w4082_,
		_w4083_,
		_w4084_
	);
	LUT3 #(
		.INIT('h2b)
	) name4019 (
		_w3960_,
		_w3961_,
		_w3962_,
		_w4085_
	);
	LUT3 #(
		.INIT('h96)
	) name4020 (
		_w4081_,
		_w4084_,
		_w4085_,
		_w4086_
	);
	LUT4 #(
		.INIT('he800)
	) name4021 (
		_w3831_,
		_w3832_,
		_w3833_,
		_w3992_,
		_w4087_
	);
	LUT3 #(
		.INIT('h17)
	) name4022 (
		_w3975_,
		_w3992_,
		_w4010_,
		_w4088_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name4023 (
		_w4012_,
		_w4014_,
		_w4086_,
		_w4087_,
		_w4089_
	);
	LUT3 #(
		.INIT('h32)
	) name4024 (
		_w4052_,
		_w4053_,
		_w4058_,
		_w4090_
	);
	LUT3 #(
		.INIT('h0d)
	) name4025 (
		_w4048_,
		_w4049_,
		_w4050_,
		_w4091_
	);
	LUT3 #(
		.INIT('h0d)
	) name4026 (
		_w3981_,
		_w3982_,
		_w3983_,
		_w4092_
	);
	LUT2 #(
		.INIT('h8)
	) name4027 (
		\a[3] ,
		\a[59] ,
		_w4093_
	);
	LUT4 #(
		.INIT('h153f)
	) name4028 (
		\a[4] ,
		\a[5] ,
		\a[57] ,
		\a[58] ,
		_w4094_
	);
	LUT2 #(
		.INIT('h8)
	) name4029 (
		\a[5] ,
		\a[58] ,
		_w4095_
	);
	LUT4 #(
		.INIT('h8000)
	) name4030 (
		\a[4] ,
		\a[5] ,
		\a[57] ,
		\a[58] ,
		_w4096_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4031 (
		\a[4] ,
		\a[5] ,
		\a[57] ,
		\a[58] ,
		_w4097_
	);
	LUT2 #(
		.INIT('h6)
	) name4032 (
		_w4093_,
		_w4097_,
		_w4098_
	);
	LUT3 #(
		.INIT('h69)
	) name4033 (
		_w4091_,
		_w4092_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h9)
	) name4034 (
		_w4090_,
		_w4099_,
		_w4100_
	);
	LUT3 #(
		.INIT('h54)
	) name4035 (
		_w4036_,
		_w4037_,
		_w4038_,
		_w4101_
	);
	LUT2 #(
		.INIT('h6)
	) name4036 (
		_w4100_,
		_w4101_,
		_w4102_
	);
	LUT4 #(
		.INIT('h0017)
	) name4037 (
		_w3975_,
		_w3992_,
		_w4010_,
		_w4086_,
		_w4103_
	);
	LUT3 #(
		.INIT('h04)
	) name4038 (
		_w4089_,
		_w4102_,
		_w4103_,
		_w4104_
	);
	LUT3 #(
		.INIT('h82)
	) name4039 (
		_w4086_,
		_w4100_,
		_w4101_,
		_w4105_
	);
	LUT3 #(
		.INIT('h41)
	) name4040 (
		_w4086_,
		_w4100_,
		_w4101_,
		_w4106_
	);
	LUT3 #(
		.INIT('h1b)
	) name4041 (
		_w4088_,
		_w4105_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h4)
	) name4042 (
		_w4104_,
		_w4107_,
		_w4108_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4043 (
		_w4041_,
		_w4064_,
		_w4104_,
		_w4107_,
		_w4109_
	);
	LUT3 #(
		.INIT('hb0)
	) name4044 (
		_w3936_,
		_w4080_,
		_w4109_,
		_w4110_
	);
	LUT4 #(
		.INIT('h00dc)
	) name4045 (
		_w3936_,
		_w4065_,
		_w4080_,
		_w4108_,
		_w4111_
	);
	LUT3 #(
		.INIT('h80)
	) name4046 (
		\a[1] ,
		\a[31] ,
		\a[60] ,
		_w4112_
	);
	LUT4 #(
		.INIT('h153f)
	) name4047 (
		\a[0] ,
		\a[2] ,
		\a[60] ,
		\a[62] ,
		_w4113_
	);
	LUT2 #(
		.INIT('h8)
	) name4048 (
		\a[2] ,
		\a[62] ,
		_w4114_
	);
	LUT4 #(
		.INIT('h8000)
	) name4049 (
		\a[0] ,
		\a[2] ,
		\a[60] ,
		\a[62] ,
		_w4115_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4050 (
		\a[0] ,
		\a[2] ,
		\a[60] ,
		\a[62] ,
		_w4116_
	);
	LUT4 #(
		.INIT('h153f)
	) name4051 (
		\a[25] ,
		\a[26] ,
		\a[36] ,
		\a[37] ,
		_w4117_
	);
	LUT4 #(
		.INIT('h8000)
	) name4052 (
		\a[25] ,
		\a[26] ,
		\a[36] ,
		\a[37] ,
		_w4118_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4053 (
		\a[25] ,
		\a[26] ,
		\a[36] ,
		\a[37] ,
		_w4119_
	);
	LUT4 #(
		.INIT('h1428)
	) name4054 (
		_w4000_,
		_w4112_,
		_w4116_,
		_w4119_,
		_w4120_
	);
	LUT4 #(
		.INIT('h8241)
	) name4055 (
		_w4000_,
		_w4112_,
		_w4116_,
		_w4119_,
		_w4121_
	);
	LUT4 #(
		.INIT('h6996)
	) name4056 (
		_w4000_,
		_w4112_,
		_w4116_,
		_w4119_,
		_w4122_
	);
	LUT2 #(
		.INIT('h8)
	) name4057 (
		\a[9] ,
		\a[53] ,
		_w4123_
	);
	LUT4 #(
		.INIT('h153f)
	) name4058 (
		\a[10] ,
		\a[17] ,
		\a[45] ,
		\a[52] ,
		_w4124_
	);
	LUT4 #(
		.INIT('h8000)
	) name4059 (
		\a[10] ,
		\a[17] ,
		\a[45] ,
		\a[52] ,
		_w4125_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4060 (
		\a[10] ,
		\a[17] ,
		\a[45] ,
		\a[52] ,
		_w4126_
	);
	LUT2 #(
		.INIT('h6)
	) name4061 (
		_w4123_,
		_w4126_,
		_w4127_
	);
	LUT4 #(
		.INIT('h153f)
	) name4062 (
		\a[11] ,
		\a[15] ,
		\a[47] ,
		\a[51] ,
		_w4128_
	);
	LUT4 #(
		.INIT('h8000)
	) name4063 (
		\a[11] ,
		\a[15] ,
		\a[47] ,
		\a[51] ,
		_w4129_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4064 (
		\a[11] ,
		\a[15] ,
		\a[47] ,
		\a[51] ,
		_w4130_
	);
	LUT2 #(
		.INIT('h8)
	) name4065 (
		\a[12] ,
		\a[50] ,
		_w4131_
	);
	LUT4 #(
		.INIT('h153f)
	) name4066 (
		\a[13] ,
		\a[14] ,
		\a[48] ,
		\a[49] ,
		_w4132_
	);
	LUT4 #(
		.INIT('h8000)
	) name4067 (
		\a[13] ,
		\a[14] ,
		\a[48] ,
		\a[49] ,
		_w4133_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4068 (
		\a[13] ,
		\a[14] ,
		\a[48] ,
		\a[49] ,
		_w4134_
	);
	LUT4 #(
		.INIT('h0660)
	) name4069 (
		_w2910_,
		_w4130_,
		_w4131_,
		_w4134_,
		_w4135_
	);
	LUT4 #(
		.INIT('h9009)
	) name4070 (
		_w2910_,
		_w4130_,
		_w4131_,
		_w4134_,
		_w4136_
	);
	LUT4 #(
		.INIT('h6996)
	) name4071 (
		_w2910_,
		_w4130_,
		_w4131_,
		_w4134_,
		_w4137_
	);
	LUT2 #(
		.INIT('h8)
	) name4072 (
		\a[20] ,
		\a[42] ,
		_w4138_
	);
	LUT4 #(
		.INIT('h153f)
	) name4073 (
		\a[6] ,
		\a[7] ,
		\a[55] ,
		\a[56] ,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name4074 (
		\a[7] ,
		\a[56] ,
		_w4140_
	);
	LUT4 #(
		.INIT('h8000)
	) name4075 (
		\a[6] ,
		\a[7] ,
		\a[55] ,
		\a[56] ,
		_w4141_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4076 (
		\a[6] ,
		\a[7] ,
		\a[55] ,
		\a[56] ,
		_w4142_
	);
	LUT2 #(
		.INIT('h6)
	) name4077 (
		_w4138_,
		_w4142_,
		_w4143_
	);
	LUT4 #(
		.INIT('h0660)
	) name4078 (
		_w4122_,
		_w4127_,
		_w4137_,
		_w4143_,
		_w4144_
	);
	LUT4 #(
		.INIT('h9009)
	) name4079 (
		_w4122_,
		_w4127_,
		_w4137_,
		_w4143_,
		_w4145_
	);
	LUT4 #(
		.INIT('h6996)
	) name4080 (
		_w4122_,
		_w4127_,
		_w4137_,
		_w4143_,
		_w4146_
	);
	LUT2 #(
		.INIT('h8)
	) name4081 (
		\a[19] ,
		\a[43] ,
		_w4147_
	);
	LUT4 #(
		.INIT('h153f)
	) name4082 (
		\a[8] ,
		\a[18] ,
		\a[44] ,
		\a[54] ,
		_w4148_
	);
	LUT4 #(
		.INIT('h8000)
	) name4083 (
		\a[8] ,
		\a[18] ,
		\a[44] ,
		\a[54] ,
		_w4149_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4084 (
		\a[8] ,
		\a[18] ,
		\a[44] ,
		\a[54] ,
		_w4150_
	);
	LUT2 #(
		.INIT('h8)
	) name4085 (
		\a[27] ,
		\a[35] ,
		_w4151_
	);
	LUT4 #(
		.INIT('h153f)
	) name4086 (
		\a[28] ,
		\a[29] ,
		\a[33] ,
		\a[34] ,
		_w4152_
	);
	LUT4 #(
		.INIT('h8000)
	) name4087 (
		\a[28] ,
		\a[29] ,
		\a[33] ,
		\a[34] ,
		_w4153_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4088 (
		\a[28] ,
		\a[29] ,
		\a[33] ,
		\a[34] ,
		_w4154_
	);
	LUT4 #(
		.INIT('h0660)
	) name4089 (
		_w4147_,
		_w4150_,
		_w4151_,
		_w4154_,
		_w4155_
	);
	LUT4 #(
		.INIT('h9009)
	) name4090 (
		_w4147_,
		_w4150_,
		_w4151_,
		_w4154_,
		_w4156_
	);
	LUT4 #(
		.INIT('h6996)
	) name4091 (
		_w4147_,
		_w4150_,
		_w4151_,
		_w4154_,
		_w4157_
	);
	LUT2 #(
		.INIT('h8)
	) name4092 (
		\a[22] ,
		\a[40] ,
		_w4158_
	);
	LUT4 #(
		.INIT('h153f)
	) name4093 (
		\a[23] ,
		\a[24] ,
		\a[38] ,
		\a[39] ,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name4094 (
		\a[24] ,
		\a[39] ,
		_w4160_
	);
	LUT4 #(
		.INIT('h8000)
	) name4095 (
		\a[23] ,
		\a[24] ,
		\a[38] ,
		\a[39] ,
		_w4161_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4096 (
		\a[23] ,
		\a[24] ,
		\a[38] ,
		\a[39] ,
		_w4162_
	);
	LUT2 #(
		.INIT('h6)
	) name4097 (
		_w4158_,
		_w4162_,
		_w4163_
	);
	LUT2 #(
		.INIT('h6)
	) name4098 (
		_w4157_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h6)
	) name4099 (
		_w4146_,
		_w4164_,
		_w4165_
	);
	LUT4 #(
		.INIT('hd400)
	) name4100 (
		_w4023_,
		_w4030_,
		_w4039_,
		_w4165_,
		_w4166_
	);
	LUT3 #(
		.INIT('h07)
	) name4101 (
		_w4030_,
		_w4039_,
		_w4165_,
		_w4167_
	);
	LUT3 #(
		.INIT('hb0)
	) name4102 (
		_w4023_,
		_w4040_,
		_w4167_,
		_w4168_
	);
	LUT3 #(
		.INIT('h32)
	) name4103 (
		_w3950_,
		_w3970_,
		_w3971_,
		_w4169_
	);
	LUT3 #(
		.INIT('he1)
	) name4104 (
		_w4166_,
		_w4168_,
		_w4169_,
		_w4170_
	);
	LUT3 #(
		.INIT('he1)
	) name4105 (
		_w4110_,
		_w4111_,
		_w4170_,
		_w4171_
	);
	LUT4 #(
		.INIT('h1f01)
	) name4106 (
		_w3841_,
		_w3949_,
		_w3973_,
		_w4019_,
		_w4172_
	);
	LUT3 #(
		.INIT('h71)
	) name4107 (
		_w3963_,
		_w3967_,
		_w3968_,
		_w4173_
	);
	LUT3 #(
		.INIT('he8)
	) name4108 (
		_w4024_,
		_w4025_,
		_w4029_,
		_w4174_
	);
	LUT2 #(
		.INIT('h1)
	) name4109 (
		_w4173_,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h8)
	) name4110 (
		_w4173_,
		_w4174_,
		_w4176_
	);
	LUT2 #(
		.INIT('h6)
	) name4111 (
		_w4173_,
		_w4174_,
		_w4177_
	);
	LUT3 #(
		.INIT('h54)
	) name4112 (
		_w3956_,
		_w3957_,
		_w3959_,
		_w4178_
	);
	LUT2 #(
		.INIT('h6)
	) name4113 (
		_w4177_,
		_w4178_,
		_w4179_
	);
	LUT3 #(
		.INIT('h0d)
	) name4114 (
		_w3974_,
		_w4016_,
		_w4017_,
		_w4180_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4115 (
		_w3974_,
		_w4016_,
		_w4017_,
		_w4179_,
		_w4181_
	);
	LUT3 #(
		.INIT('h23)
	) name4116 (
		_w4042_,
		_w4061_,
		_w4062_,
		_w4182_
	);
	LUT3 #(
		.INIT('h2b)
	) name4117 (
		_w3964_,
		_w3965_,
		_w3966_,
		_w4183_
	);
	LUT3 #(
		.INIT('h32)
	) name4118 (
		_w4003_,
		_w4004_,
		_w4009_,
		_w4184_
	);
	LUT3 #(
		.INIT('h32)
	) name4119 (
		_w3985_,
		_w3986_,
		_w3991_,
		_w4185_
	);
	LUT3 #(
		.INIT('h96)
	) name4120 (
		_w4183_,
		_w4184_,
		_w4185_,
		_w4186_
	);
	LUT3 #(
		.INIT('h0d)
	) name4121 (
		_w3998_,
		_w3999_,
		_w4001_,
		_w4187_
	);
	LUT3 #(
		.INIT('h0d)
	) name4122 (
		_w3993_,
		_w3994_,
		_w3996_,
		_w4188_
	);
	LUT3 #(
		.INIT('h0d)
	) name4123 (
		_w4044_,
		_w4045_,
		_w4046_,
		_w4189_
	);
	LUT3 #(
		.INIT('h96)
	) name4124 (
		_w4187_,
		_w4188_,
		_w4189_,
		_w4190_
	);
	LUT3 #(
		.INIT('h0d)
	) name4125 (
		_w3882_,
		_w4055_,
		_w4056_,
		_w4191_
	);
	LUT3 #(
		.INIT('h0d)
	) name4126 (
		_w4031_,
		_w4032_,
		_w4033_,
		_w4192_
	);
	LUT3 #(
		.INIT('h0d)
	) name4127 (
		_w3874_,
		_w4006_,
		_w4007_,
		_w4193_
	);
	LUT3 #(
		.INIT('h96)
	) name4128 (
		_w4191_,
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT4 #(
		.INIT('h8000)
	) name4129 (
		\a[1] ,
		\a[30] ,
		\a[32] ,
		\a[61] ,
		_w4195_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4130 (
		\a[1] ,
		\a[30] ,
		\a[32] ,
		\a[61] ,
		_w4196_
	);
	LUT4 #(
		.INIT('h000d)
	) name4131 (
		_w3915_,
		_w3988_,
		_w3989_,
		_w4196_,
		_w4197_
	);
	LUT4 #(
		.INIT('hf200)
	) name4132 (
		_w3915_,
		_w3988_,
		_w3989_,
		_w4196_,
		_w4198_
	);
	LUT4 #(
		.INIT('h0df2)
	) name4133 (
		_w3915_,
		_w3988_,
		_w3989_,
		_w4196_,
		_w4199_
	);
	LUT3 #(
		.INIT('h0d)
	) name4134 (
		_w3976_,
		_w3977_,
		_w3979_,
		_w4200_
	);
	LUT2 #(
		.INIT('h6)
	) name4135 (
		_w4199_,
		_w4200_,
		_w4201_
	);
	LUT3 #(
		.INIT('h69)
	) name4136 (
		_w4190_,
		_w4194_,
		_w4201_,
		_w4202_
	);
	LUT2 #(
		.INIT('h8)
	) name4137 (
		_w4186_,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h6)
	) name4138 (
		_w4186_,
		_w4202_,
		_w4204_
	);
	LUT3 #(
		.INIT('he1)
	) name4139 (
		_w4060_,
		_w4182_,
		_w4204_,
		_w4205_
	);
	LUT4 #(
		.INIT('h32ff)
	) name4140 (
		_w3974_,
		_w4016_,
		_w4017_,
		_w4179_,
		_w4206_
	);
	LUT3 #(
		.INIT('h40)
	) name4141 (
		_w4181_,
		_w4205_,
		_w4206_,
		_w4207_
	);
	LUT4 #(
		.INIT('hf200)
	) name4142 (
		_w3974_,
		_w4016_,
		_w4017_,
		_w4179_,
		_w4208_
	);
	LUT4 #(
		.INIT('h000d)
	) name4143 (
		_w3974_,
		_w4016_,
		_w4017_,
		_w4179_,
		_w4209_
	);
	LUT3 #(
		.INIT('h01)
	) name4144 (
		_w4205_,
		_w4208_,
		_w4209_,
		_w4210_
	);
	LUT3 #(
		.INIT('h02)
	) name4145 (
		_w4172_,
		_w4207_,
		_w4210_,
		_w4211_
	);
	LUT3 #(
		.INIT('h54)
	) name4146 (
		_w4172_,
		_w4207_,
		_w4210_,
		_w4212_
	);
	LUT3 #(
		.INIT('ha9)
	) name4147 (
		_w4172_,
		_w4207_,
		_w4210_,
		_w4213_
	);
	LUT3 #(
		.INIT('h28)
	) name4148 (
		_w4079_,
		_w4171_,
		_w4213_,
		_w4214_
	);
	LUT3 #(
		.INIT('h41)
	) name4149 (
		_w4079_,
		_w4171_,
		_w4213_,
		_w4215_
	);
	LUT3 #(
		.INIT('h96)
	) name4150 (
		_w4079_,
		_w4171_,
		_w4213_,
		_w4216_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4151 (
		_w3940_,
		_w4072_,
		_w4074_,
		_w4216_,
		_w4217_
	);
	LUT3 #(
		.INIT('h0d)
	) name4152 (
		_w3940_,
		_w4072_,
		_w4074_,
		_w4218_
	);
	LUT4 #(
		.INIT('h8d8c)
	) name4153 (
		_w4078_,
		_w4216_,
		_w4217_,
		_w4218_,
		_w4219_
	);
	LUT4 #(
		.INIT('h000d)
	) name4154 (
		_w3940_,
		_w4072_,
		_w4074_,
		_w4215_,
		_w4220_
	);
	LUT3 #(
		.INIT('h0e)
	) name4155 (
		_w4171_,
		_w4211_,
		_w4212_,
		_w4221_
	);
	LUT4 #(
		.INIT('h004f)
	) name4156 (
		_w3936_,
		_w4080_,
		_w4109_,
		_w4170_,
		_w4222_
	);
	LUT3 #(
		.INIT('h45)
	) name4157 (
		_w4166_,
		_w4168_,
		_w4169_,
		_w4223_
	);
	LUT3 #(
		.INIT('h17)
	) name4158 (
		_w4190_,
		_w4194_,
		_w4201_,
		_w4224_
	);
	LUT3 #(
		.INIT('he8)
	) name4159 (
		_w4183_,
		_w4184_,
		_w4185_,
		_w4225_
	);
	LUT2 #(
		.INIT('h1)
	) name4160 (
		_w4224_,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h8)
	) name4161 (
		_w4224_,
		_w4225_,
		_w4227_
	);
	LUT2 #(
		.INIT('h6)
	) name4162 (
		_w4224_,
		_w4225_,
		_w4228_
	);
	LUT3 #(
		.INIT('hb2)
	) name4163 (
		_w4090_,
		_w4099_,
		_w4101_,
		_w4229_
	);
	LUT2 #(
		.INIT('h9)
	) name4164 (
		_w4228_,
		_w4229_,
		_w4230_
	);
	LUT3 #(
		.INIT('h17)
	) name4165 (
		_w4191_,
		_w4192_,
		_w4193_,
		_w4231_
	);
	LUT3 #(
		.INIT('h8e)
	) name4166 (
		_w4091_,
		_w4092_,
		_w4098_,
		_w4232_
	);
	LUT3 #(
		.INIT('h45)
	) name4167 (
		_w4197_,
		_w4198_,
		_w4200_,
		_w4233_
	);
	LUT3 #(
		.INIT('h69)
	) name4168 (
		_w4231_,
		_w4232_,
		_w4233_,
		_w4234_
	);
	LUT3 #(
		.INIT('h32)
	) name4169 (
		_w4144_,
		_w4145_,
		_w4164_,
		_w4235_
	);
	LUT3 #(
		.INIT('h0d)
	) name4170 (
		_w4158_,
		_w4159_,
		_w4161_,
		_w4236_
	);
	LUT3 #(
		.INIT('h0d)
	) name4171 (
		_w4138_,
		_w4139_,
		_w4141_,
		_w4237_
	);
	LUT3 #(
		.INIT('h0d)
	) name4172 (
		_w4131_,
		_w4132_,
		_w4133_,
		_w4238_
	);
	LUT3 #(
		.INIT('h96)
	) name4173 (
		_w4236_,
		_w4237_,
		_w4238_,
		_w4239_
	);
	LUT3 #(
		.INIT('h0d)
	) name4174 (
		_w4093_,
		_w4094_,
		_w4096_,
		_w4240_
	);
	LUT3 #(
		.INIT('h0d)
	) name4175 (
		_w4000_,
		_w4117_,
		_w4118_,
		_w4241_
	);
	LUT3 #(
		.INIT('h0d)
	) name4176 (
		_w4112_,
		_w4113_,
		_w4115_,
		_w4242_
	);
	LUT3 #(
		.INIT('h96)
	) name4177 (
		_w4240_,
		_w4241_,
		_w4242_,
		_w4243_
	);
	LUT3 #(
		.INIT('h17)
	) name4178 (
		_w4187_,
		_w4188_,
		_w4189_,
		_w4244_
	);
	LUT3 #(
		.INIT('h96)
	) name4179 (
		_w4239_,
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT3 #(
		.INIT('h96)
	) name4180 (
		_w4234_,
		_w4235_,
		_w4245_,
		_w4246_
	);
	LUT3 #(
		.INIT('h60)
	) name4181 (
		_w4228_,
		_w4229_,
		_w4246_,
		_w4247_
	);
	LUT3 #(
		.INIT('h96)
	) name4182 (
		_w4228_,
		_w4229_,
		_w4246_,
		_w4248_
	);
	LUT4 #(
		.INIT('hba00)
	) name4183 (
		_w4166_,
		_w4168_,
		_w4169_,
		_w4248_,
		_w4249_
	);
	LUT4 #(
		.INIT('h45ba)
	) name4184 (
		_w4166_,
		_w4168_,
		_w4169_,
		_w4248_,
		_w4250_
	);
	LUT3 #(
		.INIT('h0e)
	) name4185 (
		_w4111_,
		_w4222_,
		_w4250_,
		_w4251_
	);
	LUT3 #(
		.INIT('h10)
	) name4186 (
		_w4111_,
		_w4222_,
		_w4250_,
		_w4252_
	);
	LUT3 #(
		.INIT('he1)
	) name4187 (
		_w4111_,
		_w4222_,
		_w4250_,
		_w4253_
	);
	LUT3 #(
		.INIT('h0d)
	) name4188 (
		_w4151_,
		_w4152_,
		_w4153_,
		_w4254_
	);
	LUT3 #(
		.INIT('h0d)
	) name4189 (
		_w4123_,
		_w4124_,
		_w4125_,
		_w4255_
	);
	LUT3 #(
		.INIT('h0d)
	) name4190 (
		_w4147_,
		_w4148_,
		_w4149_,
		_w4256_
	);
	LUT3 #(
		.INIT('h96)
	) name4191 (
		_w4254_,
		_w4255_,
		_w4256_,
		_w4257_
	);
	LUT3 #(
		.INIT('h32)
	) name4192 (
		_w4155_,
		_w4156_,
		_w4163_,
		_w4258_
	);
	LUT3 #(
		.INIT('h32)
	) name4193 (
		_w4135_,
		_w4136_,
		_w4143_,
		_w4259_
	);
	LUT3 #(
		.INIT('h69)
	) name4194 (
		_w4257_,
		_w4258_,
		_w4259_,
		_w4260_
	);
	LUT3 #(
		.INIT('he8)
	) name4195 (
		_w4081_,
		_w4084_,
		_w4085_,
		_w4261_
	);
	LUT3 #(
		.INIT('h32)
	) name4196 (
		_w4120_,
		_w4121_,
		_w4127_,
		_w4262_
	);
	LUT3 #(
		.INIT('h93)
	) name4197 (
		\a[1] ,
		\a[32] ,
		\a[62] ,
		_w4263_
	);
	LUT2 #(
		.INIT('h8)
	) name4198 (
		\a[0] ,
		\a[63] ,
		_w4264_
	);
	LUT3 #(
		.INIT('h69)
	) name4199 (
		_w4195_,
		_w4263_,
		_w4264_,
		_w4265_
	);
	LUT4 #(
		.INIT('h153f)
	) name4200 (
		\a[25] ,
		\a[26] ,
		\a[37] ,
		\a[38] ,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name4201 (
		\a[26] ,
		\a[38] ,
		_w4267_
	);
	LUT4 #(
		.INIT('h8000)
	) name4202 (
		\a[25] ,
		\a[26] ,
		\a[37] ,
		\a[38] ,
		_w4268_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4203 (
		\a[25] ,
		\a[26] ,
		\a[37] ,
		\a[38] ,
		_w4269_
	);
	LUT2 #(
		.INIT('h8)
	) name4204 (
		\a[27] ,
		\a[36] ,
		_w4270_
	);
	LUT4 #(
		.INIT('h153f)
	) name4205 (
		\a[28] ,
		\a[29] ,
		\a[34] ,
		\a[35] ,
		_w4271_
	);
	LUT4 #(
		.INIT('h8000)
	) name4206 (
		\a[28] ,
		\a[29] ,
		\a[34] ,
		\a[35] ,
		_w4272_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4207 (
		\a[28] ,
		\a[29] ,
		\a[34] ,
		\a[35] ,
		_w4273_
	);
	LUT4 #(
		.INIT('h0660)
	) name4208 (
		_w4160_,
		_w4269_,
		_w4270_,
		_w4273_,
		_w4274_
	);
	LUT4 #(
		.INIT('h9009)
	) name4209 (
		_w4160_,
		_w4269_,
		_w4270_,
		_w4273_,
		_w4275_
	);
	LUT4 #(
		.INIT('h6996)
	) name4210 (
		_w4160_,
		_w4269_,
		_w4270_,
		_w4273_,
		_w4276_
	);
	LUT2 #(
		.INIT('h6)
	) name4211 (
		_w4265_,
		_w4276_,
		_w4277_
	);
	LUT4 #(
		.INIT('h1441)
	) name4212 (
		_w4260_,
		_w4261_,
		_w4262_,
		_w4277_,
		_w4278_
	);
	LUT4 #(
		.INIT('h8228)
	) name4213 (
		_w4260_,
		_w4261_,
		_w4262_,
		_w4277_,
		_w4279_
	);
	LUT4 #(
		.INIT('h6996)
	) name4214 (
		_w4260_,
		_w4261_,
		_w4262_,
		_w4277_,
		_w4280_
	);
	LUT4 #(
		.INIT('hab54)
	) name4215 (
		_w4175_,
		_w4176_,
		_w4178_,
		_w4280_,
		_w4281_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4216 (
		_w4181_,
		_w4205_,
		_w4206_,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h8)
	) name4217 (
		_w4205_,
		_w4281_,
		_w4283_
	);
	LUT3 #(
		.INIT('h80)
	) name4218 (
		_w4179_,
		_w4205_,
		_w4281_,
		_w4284_
	);
	LUT3 #(
		.INIT('h07)
	) name4219 (
		_w4180_,
		_w4283_,
		_w4284_,
		_w4285_
	);
	LUT4 #(
		.INIT('ha140)
	) name4220 (
		_w4175_,
		_w4176_,
		_w4178_,
		_w4280_,
		_w4286_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4221 (
		_w3974_,
		_w4016_,
		_w4017_,
		_w4286_,
		_w4287_
	);
	LUT3 #(
		.INIT('h51)
	) name4222 (
		_w4089_,
		_w4102_,
		_w4103_,
		_w4288_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		\a[18] ,
		\a[45] ,
		_w4289_
	);
	LUT4 #(
		.INIT('h153f)
	) name4224 (
		\a[9] ,
		\a[17] ,
		\a[46] ,
		\a[54] ,
		_w4290_
	);
	LUT4 #(
		.INIT('h8000)
	) name4225 (
		\a[9] ,
		\a[17] ,
		\a[46] ,
		\a[54] ,
		_w4291_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4226 (
		\a[9] ,
		\a[17] ,
		\a[46] ,
		\a[54] ,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		\a[10] ,
		\a[53] ,
		_w4293_
	);
	LUT4 #(
		.INIT('h153f)
	) name4228 (
		\a[11] ,
		\a[16] ,
		\a[47] ,
		\a[52] ,
		_w4294_
	);
	LUT4 #(
		.INIT('h8000)
	) name4229 (
		\a[11] ,
		\a[16] ,
		\a[47] ,
		\a[52] ,
		_w4295_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4230 (
		\a[11] ,
		\a[16] ,
		\a[47] ,
		\a[52] ,
		_w4296_
	);
	LUT4 #(
		.INIT('h0660)
	) name4231 (
		_w4289_,
		_w4292_,
		_w4293_,
		_w4296_,
		_w4297_
	);
	LUT4 #(
		.INIT('h9009)
	) name4232 (
		_w4289_,
		_w4292_,
		_w4293_,
		_w4296_,
		_w4298_
	);
	LUT4 #(
		.INIT('h6996)
	) name4233 (
		_w4289_,
		_w4292_,
		_w4293_,
		_w4296_,
		_w4299_
	);
	LUT4 #(
		.INIT('h153f)
	) name4234 (
		\a[12] ,
		\a[13] ,
		\a[50] ,
		\a[51] ,
		_w4300_
	);
	LUT2 #(
		.INIT('h8)
	) name4235 (
		\a[13] ,
		\a[51] ,
		_w4301_
	);
	LUT4 #(
		.INIT('h8000)
	) name4236 (
		\a[12] ,
		\a[13] ,
		\a[50] ,
		\a[51] ,
		_w4302_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4237 (
		\a[12] ,
		\a[13] ,
		\a[50] ,
		\a[51] ,
		_w4303_
	);
	LUT2 #(
		.INIT('h6)
	) name4238 (
		_w3369_,
		_w4303_,
		_w4304_
	);
	LUT2 #(
		.INIT('h6)
	) name4239 (
		_w4299_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name4240 (
		\a[2] ,
		\a[61] ,
		_w4306_
	);
	LUT4 #(
		.INIT('h153f)
	) name4241 (
		\a[3] ,
		\a[4] ,
		\a[59] ,
		\a[60] ,
		_w4307_
	);
	LUT4 #(
		.INIT('h8000)
	) name4242 (
		\a[3] ,
		\a[4] ,
		\a[59] ,
		\a[60] ,
		_w4308_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4243 (
		\a[3] ,
		\a[4] ,
		\a[59] ,
		\a[60] ,
		_w4309_
	);
	LUT2 #(
		.INIT('h6)
	) name4244 (
		_w4306_,
		_w4309_,
		_w4310_
	);
	LUT3 #(
		.INIT('h0d)
	) name4245 (
		_w2910_,
		_w4128_,
		_w4129_,
		_w4311_
	);
	LUT4 #(
		.INIT('h153f)
	) name4246 (
		\a[21] ,
		\a[22] ,
		\a[41] ,
		\a[42] ,
		_w4312_
	);
	LUT4 #(
		.INIT('h8000)
	) name4247 (
		\a[21] ,
		\a[22] ,
		\a[41] ,
		\a[42] ,
		_w4313_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4248 (
		\a[21] ,
		\a[22] ,
		\a[41] ,
		\a[42] ,
		_w4314_
	);
	LUT2 #(
		.INIT('h6)
	) name4249 (
		_w4095_,
		_w4314_,
		_w4315_
	);
	LUT3 #(
		.INIT('h69)
	) name4250 (
		_w4310_,
		_w4311_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name4251 (
		\a[23] ,
		\a[40] ,
		_w4317_
	);
	LUT4 #(
		.INIT('h153f)
	) name4252 (
		\a[6] ,
		\a[20] ,
		\a[43] ,
		\a[57] ,
		_w4318_
	);
	LUT4 #(
		.INIT('h8000)
	) name4253 (
		\a[6] ,
		\a[20] ,
		\a[43] ,
		\a[57] ,
		_w4319_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4254 (
		\a[6] ,
		\a[20] ,
		\a[43] ,
		\a[57] ,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name4255 (
		\a[31] ,
		\a[32] ,
		_w4321_
	);
	LUT2 #(
		.INIT('h8)
	) name4256 (
		\a[30] ,
		\a[33] ,
		_w4322_
	);
	LUT4 #(
		.INIT('h153f)
	) name4257 (
		\a[30] ,
		\a[31] ,
		\a[32] ,
		\a[33] ,
		_w4323_
	);
	LUT4 #(
		.INIT('h8000)
	) name4258 (
		\a[30] ,
		\a[31] ,
		\a[32] ,
		\a[33] ,
		_w4324_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4259 (
		\a[30] ,
		\a[31] ,
		\a[32] ,
		\a[33] ,
		_w4325_
	);
	LUT4 #(
		.INIT('h1428)
	) name4260 (
		_w3978_,
		_w4317_,
		_w4320_,
		_w4325_,
		_w4326_
	);
	LUT4 #(
		.INIT('h8241)
	) name4261 (
		_w3978_,
		_w4317_,
		_w4320_,
		_w4325_,
		_w4327_
	);
	LUT4 #(
		.INIT('h6996)
	) name4262 (
		_w3978_,
		_w4317_,
		_w4320_,
		_w4325_,
		_w4328_
	);
	LUT4 #(
		.INIT('h153f)
	) name4263 (
		\a[8] ,
		\a[19] ,
		\a[44] ,
		\a[55] ,
		_w4329_
	);
	LUT4 #(
		.INIT('h8000)
	) name4264 (
		\a[8] ,
		\a[19] ,
		\a[44] ,
		\a[55] ,
		_w4330_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4265 (
		\a[8] ,
		\a[19] ,
		\a[44] ,
		\a[55] ,
		_w4331_
	);
	LUT2 #(
		.INIT('h6)
	) name4266 (
		_w4140_,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h6)
	) name4267 (
		_w4328_,
		_w4332_,
		_w4333_
	);
	LUT3 #(
		.INIT('h96)
	) name4268 (
		_w4305_,
		_w4316_,
		_w4333_,
		_w4334_
	);
	LUT4 #(
		.INIT('hae00)
	) name4269 (
		_w4089_,
		_w4102_,
		_w4103_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w4186_,
		_w4202_,
		_w4336_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4271 (
		_w4060_,
		_w4182_,
		_w4203_,
		_w4336_,
		_w4337_
	);
	LUT4 #(
		.INIT('h0051)
	) name4272 (
		_w4089_,
		_w4102_,
		_w4103_,
		_w4334_,
		_w4338_
	);
	LUT4 #(
		.INIT('hf949)
	) name4273 (
		_w4288_,
		_w4334_,
		_w4337_,
		_w4338_,
		_w4339_
	);
	LUT4 #(
		.INIT('h17ff)
	) name4274 (
		_w4179_,
		_w4180_,
		_w4205_,
		_w4281_,
		_w4340_
	);
	LUT4 #(
		.INIT('hfb04)
	) name4275 (
		_w4282_,
		_w4285_,
		_w4287_,
		_w4339_,
		_w4341_
	);
	LUT2 #(
		.INIT('h6)
	) name4276 (
		_w4253_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h6)
	) name4277 (
		_w4221_,
		_w4342_,
		_w4343_
	);
	LUT4 #(
		.INIT('h23dc)
	) name4278 (
		_w4078_,
		_w4214_,
		_w4220_,
		_w4343_,
		_w4344_
	);
	LUT3 #(
		.INIT('h15)
	) name4279 (
		_w4214_,
		_w4221_,
		_w4342_,
		_w4345_
	);
	LUT2 #(
		.INIT('h1)
	) name4280 (
		_w4287_,
		_w4339_,
		_w4346_
	);
	LUT2 #(
		.INIT('h8)
	) name4281 (
		_w4285_,
		_w4346_,
		_w4347_
	);
	LUT2 #(
		.INIT('h8)
	) name4282 (
		_w4282_,
		_w4340_,
		_w4348_
	);
	LUT4 #(
		.INIT('h0017)
	) name4283 (
		_w4173_,
		_w4174_,
		_w4178_,
		_w4279_,
		_w4349_
	);
	LUT2 #(
		.INIT('h1)
	) name4284 (
		_w4278_,
		_w4349_,
		_w4350_
	);
	LUT4 #(
		.INIT('h0017)
	) name4285 (
		_w4081_,
		_w4084_,
		_w4085_,
		_w4262_,
		_w4351_
	);
	LUT4 #(
		.INIT('he800)
	) name4286 (
		_w4081_,
		_w4084_,
		_w4085_,
		_w4262_,
		_w4352_
	);
	LUT3 #(
		.INIT('h32)
	) name4287 (
		_w4277_,
		_w4351_,
		_w4352_,
		_w4353_
	);
	LUT3 #(
		.INIT('he8)
	) name4288 (
		_w4305_,
		_w4316_,
		_w4333_,
		_w4354_
	);
	LUT3 #(
		.INIT('h0e)
	) name4289 (
		_w4265_,
		_w4274_,
		_w4275_,
		_w4355_
	);
	LUT3 #(
		.INIT('h32)
	) name4290 (
		_w4317_,
		_w4318_,
		_w4319_,
		_w4356_
	);
	LUT3 #(
		.INIT('h0d)
	) name4291 (
		_w4289_,
		_w4290_,
		_w4291_,
		_w4357_
	);
	LUT3 #(
		.INIT('h0d)
	) name4292 (
		_w4270_,
		_w4271_,
		_w4272_,
		_w4358_
	);
	LUT3 #(
		.INIT('h69)
	) name4293 (
		_w4356_,
		_w4357_,
		_w4358_,
		_w4359_
	);
	LUT3 #(
		.INIT('h0d)
	) name4294 (
		_w4306_,
		_w4307_,
		_w4308_,
		_w4360_
	);
	LUT3 #(
		.INIT('h0d)
	) name4295 (
		_w4095_,
		_w4312_,
		_w4313_,
		_w4361_
	);
	LUT3 #(
		.INIT('h0d)
	) name4296 (
		_w4140_,
		_w4329_,
		_w4330_,
		_w4362_
	);
	LUT3 #(
		.INIT('h96)
	) name4297 (
		_w4360_,
		_w4361_,
		_w4362_,
		_w4363_
	);
	LUT3 #(
		.INIT('h96)
	) name4298 (
		_w4355_,
		_w4359_,
		_w4363_,
		_w4364_
	);
	LUT2 #(
		.INIT('h1)
	) name4299 (
		_w4354_,
		_w4364_,
		_w4365_
	);
	LUT3 #(
		.INIT('h96)
	) name4300 (
		_w4353_,
		_w4354_,
		_w4364_,
		_w4366_
	);
	LUT3 #(
		.INIT('h10)
	) name4301 (
		_w4278_,
		_w4349_,
		_w4366_,
		_w4367_
	);
	LUT3 #(
		.INIT('h0e)
	) name4302 (
		_w4278_,
		_w4349_,
		_w4366_,
		_w4368_
	);
	LUT3 #(
		.INIT('he1)
	) name4303 (
		_w4278_,
		_w4349_,
		_w4366_,
		_w4369_
	);
	LUT3 #(
		.INIT('h51)
	) name4304 (
		_w4335_,
		_w4337_,
		_w4338_,
		_w4370_
	);
	LUT2 #(
		.INIT('h6)
	) name4305 (
		_w4369_,
		_w4370_,
		_w4371_
	);
	LUT3 #(
		.INIT('h54)
	) name4306 (
		_w4226_,
		_w4227_,
		_w4229_,
		_w4372_
	);
	LUT3 #(
		.INIT('h0d)
	) name4307 (
		_w3369_,
		_w4300_,
		_w4302_,
		_w4373_
	);
	LUT3 #(
		.INIT('h0d)
	) name4308 (
		_w4160_,
		_w4266_,
		_w4268_,
		_w4374_
	);
	LUT3 #(
		.INIT('h0d)
	) name4309 (
		_w4293_,
		_w4294_,
		_w4295_,
		_w4375_
	);
	LUT3 #(
		.INIT('h96)
	) name4310 (
		_w4373_,
		_w4374_,
		_w4375_,
		_w4376_
	);
	LUT3 #(
		.INIT('h32)
	) name4311 (
		_w4326_,
		_w4327_,
		_w4332_,
		_w4377_
	);
	LUT3 #(
		.INIT('h32)
	) name4312 (
		_w4297_,
		_w4298_,
		_w4304_,
		_w4378_
	);
	LUT3 #(
		.INIT('h69)
	) name4313 (
		_w4376_,
		_w4377_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('hb2)
	) name4314 (
		_w4231_,
		_w4232_,
		_w4233_,
		_w4380_
	);
	LUT4 #(
		.INIT('h8000)
	) name4315 (
		\a[1] ,
		\a[32] ,
		\a[62] ,
		\a[63] ,
		_w4381_
	);
	LUT2 #(
		.INIT('h8)
	) name4316 (
		\a[32] ,
		\a[62] ,
		_w4382_
	);
	LUT4 #(
		.INIT('h2a80)
	) name4317 (
		\a[1] ,
		\a[32] ,
		\a[62] ,
		\a[63] ,
		_w4383_
	);
	LUT4 #(
		.INIT('he800)
	) name4318 (
		_w3978_,
		_w4321_,
		_w4322_,
		_w4383_,
		_w4384_
	);
	LUT4 #(
		.INIT('hcd32)
	) name4319 (
		_w3978_,
		_w4323_,
		_w4324_,
		_w4383_,
		_w4385_
	);
	LUT4 #(
		.INIT('h153f)
	) name4320 (
		\a[11] ,
		\a[12] ,
		\a[52] ,
		\a[53] ,
		_w4386_
	);
	LUT2 #(
		.INIT('h8)
	) name4321 (
		\a[12] ,
		\a[53] ,
		_w4387_
	);
	LUT4 #(
		.INIT('h8000)
	) name4322 (
		\a[11] ,
		\a[12] ,
		\a[52] ,
		\a[53] ,
		_w4388_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4323 (
		\a[11] ,
		\a[12] ,
		\a[52] ,
		\a[53] ,
		_w4389_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		\a[9] ,
		\a[55] ,
		_w4390_
	);
	LUT4 #(
		.INIT('h153f)
	) name4325 (
		\a[10] ,
		\a[15] ,
		\a[49] ,
		\a[54] ,
		_w4391_
	);
	LUT4 #(
		.INIT('h8000)
	) name4326 (
		\a[10] ,
		\a[15] ,
		\a[49] ,
		\a[54] ,
		_w4392_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4327 (
		\a[10] ,
		\a[15] ,
		\a[49] ,
		\a[54] ,
		_w4393_
	);
	LUT4 #(
		.INIT('h0660)
	) name4328 (
		_w4301_,
		_w4389_,
		_w4390_,
		_w4393_,
		_w4394_
	);
	LUT4 #(
		.INIT('h9009)
	) name4329 (
		_w4301_,
		_w4389_,
		_w4390_,
		_w4393_,
		_w4395_
	);
	LUT4 #(
		.INIT('h6996)
	) name4330 (
		_w4301_,
		_w4389_,
		_w4390_,
		_w4393_,
		_w4396_
	);
	LUT2 #(
		.INIT('h6)
	) name4331 (
		_w4385_,
		_w4396_,
		_w4397_
	);
	LUT3 #(
		.INIT('hb2)
	) name4332 (
		_w4310_,
		_w4311_,
		_w4315_,
		_w4398_
	);
	LUT4 #(
		.INIT('h00b2)
	) name4333 (
		_w4231_,
		_w4232_,
		_w4233_,
		_w4398_,
		_w4399_
	);
	LUT4 #(
		.INIT('hed61)
	) name4334 (
		_w4380_,
		_w4397_,
		_w4398_,
		_w4399_,
		_w4400_
	);
	LUT3 #(
		.INIT('h0e)
	) name4335 (
		_w4224_,
		_w4225_,
		_w4379_,
		_w4401_
	);
	LUT3 #(
		.INIT('he0)
	) name4336 (
		_w4227_,
		_w4229_,
		_w4401_,
		_w4402_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4337 (
		_w4227_,
		_w4229_,
		_w4400_,
		_w4401_,
		_w4403_
	);
	LUT2 #(
		.INIT('h2)
	) name4338 (
		_w4379_,
		_w4400_,
		_w4404_
	);
	LUT4 #(
		.INIT('h606b)
	) name4339 (
		_w4372_,
		_w4379_,
		_w4400_,
		_w4402_,
		_w4405_
	);
	LUT3 #(
		.INIT('h01)
	) name4340 (
		_w4247_,
		_w4249_,
		_w4405_,
		_w4406_
	);
	LUT4 #(
		.INIT('h0045)
	) name4341 (
		_w4166_,
		_w4168_,
		_w4169_,
		_w4247_,
		_w4407_
	);
	LUT3 #(
		.INIT('h09)
	) name4342 (
		_w4228_,
		_w4229_,
		_w4246_,
		_w4408_
	);
	LUT3 #(
		.INIT('hb2)
	) name4343 (
		_w4195_,
		_w4263_,
		_w4264_,
		_w4409_
	);
	LUT4 #(
		.INIT('h153f)
	) name4344 (
		\a[18] ,
		\a[19] ,
		\a[45] ,
		\a[46] ,
		_w4410_
	);
	LUT4 #(
		.INIT('h8000)
	) name4345 (
		\a[18] ,
		\a[19] ,
		\a[45] ,
		\a[46] ,
		_w4411_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4346 (
		\a[18] ,
		\a[19] ,
		\a[45] ,
		\a[46] ,
		_w4412_
	);
	LUT2 #(
		.INIT('h6)
	) name4347 (
		_w3995_,
		_w4412_,
		_w4413_
	);
	LUT4 #(
		.INIT('h153f)
	) name4348 (
		\a[3] ,
		\a[4] ,
		\a[60] ,
		\a[61] ,
		_w4414_
	);
	LUT4 #(
		.INIT('h8000)
	) name4349 (
		\a[3] ,
		\a[4] ,
		\a[60] ,
		\a[61] ,
		_w4415_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4350 (
		\a[3] ,
		\a[4] ,
		\a[60] ,
		\a[61] ,
		_w4416_
	);
	LUT2 #(
		.INIT('h6)
	) name4351 (
		_w4114_,
		_w4416_,
		_w4417_
	);
	LUT3 #(
		.INIT('h96)
	) name4352 (
		_w4409_,
		_w4413_,
		_w4417_,
		_w4418_
	);
	LUT4 #(
		.INIT('h153f)
	) name4353 (
		\a[8] ,
		\a[16] ,
		\a[48] ,
		\a[56] ,
		_w4419_
	);
	LUT4 #(
		.INIT('h8000)
	) name4354 (
		\a[8] ,
		\a[16] ,
		\a[48] ,
		\a[56] ,
		_w4420_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4355 (
		\a[8] ,
		\a[16] ,
		\a[48] ,
		\a[56] ,
		_w4421_
	);
	LUT2 #(
		.INIT('h8)
	) name4356 (
		\a[27] ,
		\a[37] ,
		_w4422_
	);
	LUT4 #(
		.INIT('h153f)
	) name4357 (
		\a[28] ,
		\a[29] ,
		\a[35] ,
		\a[36] ,
		_w4423_
	);
	LUT2 #(
		.INIT('h8)
	) name4358 (
		\a[29] ,
		\a[36] ,
		_w4424_
	);
	LUT4 #(
		.INIT('h8000)
	) name4359 (
		\a[28] ,
		\a[29] ,
		\a[35] ,
		\a[36] ,
		_w4425_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4360 (
		\a[28] ,
		\a[29] ,
		\a[35] ,
		\a[36] ,
		_w4426_
	);
	LUT4 #(
		.INIT('h0660)
	) name4361 (
		_w4267_,
		_w4421_,
		_w4422_,
		_w4426_,
		_w4427_
	);
	LUT4 #(
		.INIT('h9009)
	) name4362 (
		_w4267_,
		_w4421_,
		_w4422_,
		_w4426_,
		_w4428_
	);
	LUT4 #(
		.INIT('h6996)
	) name4363 (
		_w4267_,
		_w4421_,
		_w4422_,
		_w4426_,
		_w4429_
	);
	LUT2 #(
		.INIT('h8)
	) name4364 (
		\a[14] ,
		\a[50] ,
		_w4430_
	);
	LUT4 #(
		.INIT('h153f)
	) name4365 (
		\a[30] ,
		\a[31] ,
		\a[33] ,
		\a[34] ,
		_w4431_
	);
	LUT4 #(
		.INIT('h8000)
	) name4366 (
		\a[30] ,
		\a[31] ,
		\a[33] ,
		\a[34] ,
		_w4432_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4367 (
		\a[30] ,
		\a[31] ,
		\a[33] ,
		\a[34] ,
		_w4433_
	);
	LUT2 #(
		.INIT('h6)
	) name4368 (
		_w4430_,
		_w4433_,
		_w4434_
	);
	LUT2 #(
		.INIT('h6)
	) name4369 (
		_w4429_,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('h8)
	) name4370 (
		\a[6] ,
		\a[58] ,
		_w4436_
	);
	LUT4 #(
		.INIT('h153f)
	) name4371 (
		\a[7] ,
		\a[17] ,
		\a[47] ,
		\a[57] ,
		_w4437_
	);
	LUT4 #(
		.INIT('h8000)
	) name4372 (
		\a[7] ,
		\a[17] ,
		\a[47] ,
		\a[57] ,
		_w4438_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4373 (
		\a[7] ,
		\a[17] ,
		\a[47] ,
		\a[57] ,
		_w4439_
	);
	LUT2 #(
		.INIT('h8)
	) name4374 (
		\a[20] ,
		\a[44] ,
		_w4440_
	);
	LUT4 #(
		.INIT('h153f)
	) name4375 (
		\a[21] ,
		\a[22] ,
		\a[42] ,
		\a[43] ,
		_w4441_
	);
	LUT4 #(
		.INIT('h8000)
	) name4376 (
		\a[21] ,
		\a[22] ,
		\a[42] ,
		\a[43] ,
		_w4442_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4377 (
		\a[21] ,
		\a[22] ,
		\a[42] ,
		\a[43] ,
		_w4443_
	);
	LUT4 #(
		.INIT('h0660)
	) name4378 (
		_w4436_,
		_w4439_,
		_w4440_,
		_w4443_,
		_w4444_
	);
	LUT4 #(
		.INIT('h9009)
	) name4379 (
		_w4436_,
		_w4439_,
		_w4440_,
		_w4443_,
		_w4445_
	);
	LUT4 #(
		.INIT('h6996)
	) name4380 (
		_w4436_,
		_w4439_,
		_w4440_,
		_w4443_,
		_w4446_
	);
	LUT2 #(
		.INIT('h8)
	) name4381 (
		\a[23] ,
		\a[41] ,
		_w4447_
	);
	LUT4 #(
		.INIT('h153f)
	) name4382 (
		\a[24] ,
		\a[25] ,
		\a[39] ,
		\a[40] ,
		_w4448_
	);
	LUT4 #(
		.INIT('h8000)
	) name4383 (
		\a[24] ,
		\a[25] ,
		\a[39] ,
		\a[40] ,
		_w4449_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4384 (
		\a[24] ,
		\a[25] ,
		\a[39] ,
		\a[40] ,
		_w4450_
	);
	LUT2 #(
		.INIT('h6)
	) name4385 (
		_w4447_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h6)
	) name4386 (
		_w4446_,
		_w4451_,
		_w4452_
	);
	LUT3 #(
		.INIT('h96)
	) name4387 (
		_w4418_,
		_w4435_,
		_w4452_,
		_w4453_
	);
	LUT4 #(
		.INIT('h0017)
	) name4388 (
		_w4234_,
		_w4235_,
		_w4245_,
		_w4453_,
		_w4454_
	);
	LUT4 #(
		.INIT('he800)
	) name4389 (
		_w4234_,
		_w4235_,
		_w4245_,
		_w4453_,
		_w4455_
	);
	LUT3 #(
		.INIT('h17)
	) name4390 (
		_w4236_,
		_w4237_,
		_w4238_,
		_w4456_
	);
	LUT3 #(
		.INIT('h17)
	) name4391 (
		_w4254_,
		_w4255_,
		_w4256_,
		_w4457_
	);
	LUT3 #(
		.INIT('h17)
	) name4392 (
		_w4240_,
		_w4241_,
		_w4242_,
		_w4458_
	);
	LUT3 #(
		.INIT('h96)
	) name4393 (
		_w4456_,
		_w4457_,
		_w4458_,
		_w4459_
	);
	LUT3 #(
		.INIT('hd4)
	) name4394 (
		_w4257_,
		_w4258_,
		_w4259_,
		_w4460_
	);
	LUT3 #(
		.INIT('h71)
	) name4395 (
		_w4239_,
		_w4243_,
		_w4244_,
		_w4461_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		_w4460_,
		_w4461_,
		_w4462_
	);
	LUT3 #(
		.INIT('h96)
	) name4397 (
		_w4459_,
		_w4460_,
		_w4461_,
		_w4463_
	);
	LUT3 #(
		.INIT('he1)
	) name4398 (
		_w4454_,
		_w4455_,
		_w4463_,
		_w4464_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4399 (
		_w4405_,
		_w4407_,
		_w4408_,
		_w4464_,
		_w4465_
	);
	LUT4 #(
		.INIT('hffa9)
	) name4400 (
		_w4405_,
		_w4407_,
		_w4408_,
		_w4464_,
		_w4466_
	);
	LUT3 #(
		.INIT('hb0)
	) name4401 (
		_w4406_,
		_w4465_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('he11e)
	) name4402 (
		_w4347_,
		_w4348_,
		_w4371_,
		_w4467_,
		_w4468_
	);
	LUT3 #(
		.INIT('h23)
	) name4403 (
		_w4251_,
		_w4252_,
		_w4341_,
		_w4469_
	);
	LUT2 #(
		.INIT('h4)
	) name4404 (
		_w4468_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('he00e)
	) name4405 (
		_w4221_,
		_w4342_,
		_w4468_,
		_w4469_,
		_w4471_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4406 (
		_w4078_,
		_w4220_,
		_w4345_,
		_w4471_,
		_w4472_
	);
	LUT4 #(
		.INIT('h0770)
	) name4407 (
		_w4221_,
		_w4342_,
		_w4468_,
		_w4469_,
		_w4473_
	);
	LUT4 #(
		.INIT('h0110)
	) name4408 (
		_w4221_,
		_w4342_,
		_w4468_,
		_w4469_,
		_w4474_
	);
	LUT2 #(
		.INIT('h4)
	) name4409 (
		_w4214_,
		_w4473_,
		_w4475_
	);
	LUT4 #(
		.INIT('h040f)
	) name4410 (
		_w4078_,
		_w4220_,
		_w4474_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h4)
	) name4411 (
		_w4472_,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('h1f01)
	) name4412 (
		_w4347_,
		_w4348_,
		_w4371_,
		_w4467_,
		_w4478_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4413 (
		_w4405_,
		_w4407_,
		_w4408_,
		_w4464_,
		_w4479_
	);
	LUT4 #(
		.INIT('h008e)
	) name4414 (
		_w4223_,
		_w4230_,
		_w4246_,
		_w4405_,
		_w4480_
	);
	LUT3 #(
		.INIT('h54)
	) name4415 (
		_w4454_,
		_w4455_,
		_w4463_,
		_w4481_
	);
	LUT3 #(
		.INIT('he0)
	) name4416 (
		_w4224_,
		_w4225_,
		_w4379_,
		_w4482_
	);
	LUT3 #(
		.INIT('he0)
	) name4417 (
		_w4227_,
		_w4229_,
		_w4482_,
		_w4483_
	);
	LUT4 #(
		.INIT('h0023)
	) name4418 (
		_w4372_,
		_w4403_,
		_w4404_,
		_w4483_,
		_w4484_
	);
	LUT2 #(
		.INIT('h8)
	) name4419 (
		_w4397_,
		_w4398_,
		_w4485_
	);
	LUT2 #(
		.INIT('h2)
	) name4420 (
		_w4397_,
		_w4398_,
		_w4486_
	);
	LUT4 #(
		.INIT('hb200)
	) name4421 (
		_w4231_,
		_w4232_,
		_w4233_,
		_w4398_,
		_w4487_
	);
	LUT4 #(
		.INIT('h001b)
	) name4422 (
		_w4380_,
		_w4485_,
		_w4486_,
		_w4487_,
		_w4488_
	);
	LUT3 #(
		.INIT('he8)
	) name4423 (
		_w4418_,
		_w4435_,
		_w4452_,
		_w4489_
	);
	LUT3 #(
		.INIT('h0e)
	) name4424 (
		_w4385_,
		_w4394_,
		_w4395_,
		_w4490_
	);
	LUT3 #(
		.INIT('h32)
	) name4425 (
		_w4390_,
		_w4391_,
		_w4392_,
		_w4491_
	);
	LUT3 #(
		.INIT('h0d)
	) name4426 (
		_w4447_,
		_w4448_,
		_w4449_,
		_w4492_
	);
	LUT3 #(
		.INIT('h0d)
	) name4427 (
		_w4436_,
		_w4437_,
		_w4438_,
		_w4493_
	);
	LUT3 #(
		.INIT('h69)
	) name4428 (
		_w4491_,
		_w4492_,
		_w4493_,
		_w4494_
	);
	LUT3 #(
		.INIT('h0d)
	) name4429 (
		_w3995_,
		_w4410_,
		_w4411_,
		_w4495_
	);
	LUT3 #(
		.INIT('h0d)
	) name4430 (
		_w4114_,
		_w4414_,
		_w4415_,
		_w4496_
	);
	LUT3 #(
		.INIT('h0d)
	) name4431 (
		_w4267_,
		_w4419_,
		_w4420_,
		_w4497_
	);
	LUT3 #(
		.INIT('h96)
	) name4432 (
		_w4495_,
		_w4496_,
		_w4497_,
		_w4498_
	);
	LUT3 #(
		.INIT('h96)
	) name4433 (
		_w4490_,
		_w4494_,
		_w4498_,
		_w4499_
	);
	LUT3 #(
		.INIT('h69)
	) name4434 (
		_w4488_,
		_w4489_,
		_w4499_,
		_w4500_
	);
	LUT3 #(
		.INIT('h69)
	) name4435 (
		_w4481_,
		_w4484_,
		_w4500_,
		_w4501_
	);
	LUT3 #(
		.INIT('h10)
	) name4436 (
		_w4479_,
		_w4480_,
		_w4501_,
		_w4502_
	);
	LUT3 #(
		.INIT('h0e)
	) name4437 (
		_w4479_,
		_w4480_,
		_w4501_,
		_w4503_
	);
	LUT3 #(
		.INIT('h23)
	) name4438 (
		_w4367_,
		_w4368_,
		_w4370_,
		_w4504_
	);
	LUT3 #(
		.INIT('h15)
	) name4439 (
		_w4459_,
		_w4460_,
		_w4461_,
		_w4505_
	);
	LUT3 #(
		.INIT('he8)
	) name4440 (
		_w4459_,
		_w4460_,
		_w4461_,
		_w4506_
	);
	LUT3 #(
		.INIT('he8)
	) name4441 (
		_w4456_,
		_w4457_,
		_w4458_,
		_w4507_
	);
	LUT2 #(
		.INIT('h8)
	) name4442 (
		\a[4] ,
		\a[63] ,
		_w4508_
	);
	LUT4 #(
		.INIT('h8000)
	) name4443 (
		\a[2] ,
		\a[4] ,
		\a[61] ,
		\a[63] ,
		_w4509_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4444 (
		\a[2] ,
		\a[4] ,
		\a[61] ,
		\a[63] ,
		_w4510_
	);
	LUT4 #(
		.INIT('hf20d)
	) name4445 (
		_w4430_,
		_w4431_,
		_w4432_,
		_w4510_,
		_w4511_
	);
	LUT4 #(
		.INIT('h153f)
	) name4446 (
		\a[14] ,
		\a[15] ,
		\a[50] ,
		\a[51] ,
		_w4512_
	);
	LUT4 #(
		.INIT('h8000)
	) name4447 (
		\a[14] ,
		\a[15] ,
		\a[50] ,
		\a[51] ,
		_w4513_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4448 (
		\a[14] ,
		\a[15] ,
		\a[50] ,
		\a[51] ,
		_w4514_
	);
	LUT4 #(
		.INIT('h153f)
	) name4449 (
		\a[13] ,
		\a[18] ,
		\a[47] ,
		\a[52] ,
		_w4515_
	);
	LUT4 #(
		.INIT('h8000)
	) name4450 (
		\a[13] ,
		\a[18] ,
		\a[47] ,
		\a[52] ,
		_w4516_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4451 (
		\a[13] ,
		\a[18] ,
		\a[47] ,
		\a[52] ,
		_w4517_
	);
	LUT4 #(
		.INIT('h1248)
	) name4452 (
		_w3535_,
		_w4387_,
		_w4514_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('h8421)
	) name4453 (
		_w3535_,
		_w4387_,
		_w4514_,
		_w4517_,
		_w4519_
	);
	LUT4 #(
		.INIT('h6996)
	) name4454 (
		_w3535_,
		_w4387_,
		_w4514_,
		_w4517_,
		_w4520_
	);
	LUT2 #(
		.INIT('h9)
	) name4455 (
		_w4511_,
		_w4520_,
		_w4521_
	);
	LUT3 #(
		.INIT('he8)
	) name4456 (
		_w4409_,
		_w4413_,
		_w4417_,
		_w4522_
	);
	LUT4 #(
		.INIT('h00e8)
	) name4457 (
		_w4456_,
		_w4457_,
		_w4458_,
		_w4522_,
		_w4523_
	);
	LUT4 #(
		.INIT('hed61)
	) name4458 (
		_w4507_,
		_w4521_,
		_w4522_,
		_w4523_,
		_w4524_
	);
	LUT3 #(
		.INIT('h0d)
	) name4459 (
		_w4440_,
		_w4441_,
		_w4442_,
		_w4525_
	);
	LUT3 #(
		.INIT('h0d)
	) name4460 (
		_w4422_,
		_w4423_,
		_w4425_,
		_w4526_
	);
	LUT3 #(
		.INIT('h0d)
	) name4461 (
		_w4301_,
		_w4386_,
		_w4388_,
		_w4527_
	);
	LUT3 #(
		.INIT('h96)
	) name4462 (
		_w4525_,
		_w4526_,
		_w4527_,
		_w4528_
	);
	LUT3 #(
		.INIT('h32)
	) name4463 (
		_w4427_,
		_w4428_,
		_w4434_,
		_w4529_
	);
	LUT3 #(
		.INIT('h32)
	) name4464 (
		_w4444_,
		_w4445_,
		_w4451_,
		_w4530_
	);
	LUT3 #(
		.INIT('h69)
	) name4465 (
		_w4528_,
		_w4529_,
		_w4530_,
		_w4531_
	);
	LUT3 #(
		.INIT('h69)
	) name4466 (
		_w4506_,
		_w4524_,
		_w4531_,
		_w4532_
	);
	LUT3 #(
		.INIT('h17)
	) name4467 (
		_w4373_,
		_w4374_,
		_w4375_,
		_w4533_
	);
	LUT3 #(
		.INIT('h2b)
	) name4468 (
		_w4356_,
		_w4357_,
		_w4358_,
		_w4534_
	);
	LUT3 #(
		.INIT('h17)
	) name4469 (
		_w4360_,
		_w4361_,
		_w4362_,
		_w4535_
	);
	LUT3 #(
		.INIT('h96)
	) name4470 (
		_w4533_,
		_w4534_,
		_w4535_,
		_w4536_
	);
	LUT3 #(
		.INIT('h2b)
	) name4471 (
		_w4355_,
		_w4359_,
		_w4363_,
		_w4537_
	);
	LUT3 #(
		.INIT('hd4)
	) name4472 (
		_w4376_,
		_w4377_,
		_w4378_,
		_w4538_
	);
	LUT3 #(
		.INIT('h96)
	) name4473 (
		_w4536_,
		_w4537_,
		_w4538_,
		_w4539_
	);
	LUT4 #(
		.INIT('h00cd)
	) name4474 (
		_w4277_,
		_w4351_,
		_w4352_,
		_w4354_,
		_w4540_
	);
	LUT4 #(
		.INIT('h00cd)
	) name4475 (
		_w4277_,
		_w4351_,
		_w4352_,
		_w4364_,
		_w4541_
	);
	LUT3 #(
		.INIT('h01)
	) name4476 (
		_w4365_,
		_w4540_,
		_w4541_,
		_w4542_
	);
	LUT2 #(
		.INIT('h8)
	) name4477 (
		\a[8] ,
		\a[57] ,
		_w4543_
	);
	LUT4 #(
		.INIT('h153f)
	) name4478 (
		\a[21] ,
		\a[22] ,
		\a[43] ,
		\a[44] ,
		_w4544_
	);
	LUT4 #(
		.INIT('h8000)
	) name4479 (
		\a[21] ,
		\a[22] ,
		\a[43] ,
		\a[44] ,
		_w4545_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4480 (
		\a[21] ,
		\a[22] ,
		\a[43] ,
		\a[44] ,
		_w4546_
	);
	LUT2 #(
		.INIT('h6)
	) name4481 (
		_w4543_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		\a[5] ,
		\a[60] ,
		_w4548_
	);
	LUT4 #(
		.INIT('h153f)
	) name4483 (
		\a[6] ,
		\a[7] ,
		\a[58] ,
		\a[59] ,
		_w4549_
	);
	LUT4 #(
		.INIT('h8000)
	) name4484 (
		\a[6] ,
		\a[7] ,
		\a[58] ,
		\a[59] ,
		_w4550_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4485 (
		\a[6] ,
		\a[7] ,
		\a[58] ,
		\a[59] ,
		_w4551_
	);
	LUT2 #(
		.INIT('h6)
	) name4486 (
		_w4548_,
		_w4551_,
		_w4552_
	);
	LUT4 #(
		.INIT('he11e)
	) name4487 (
		_w4381_,
		_w4384_,
		_w4547_,
		_w4552_,
		_w4553_
	);
	LUT4 #(
		.INIT('h153f)
	) name4488 (
		\a[11] ,
		\a[19] ,
		\a[46] ,
		\a[54] ,
		_w4554_
	);
	LUT4 #(
		.INIT('h8000)
	) name4489 (
		\a[11] ,
		\a[19] ,
		\a[46] ,
		\a[54] ,
		_w4555_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4490 (
		\a[11] ,
		\a[19] ,
		\a[46] ,
		\a[54] ,
		_w4556_
	);
	LUT2 #(
		.INIT('h8)
	) name4491 (
		\a[30] ,
		\a[35] ,
		_w4557_
	);
	LUT4 #(
		.INIT('h153f)
	) name4492 (
		\a[31] ,
		\a[32] ,
		\a[33] ,
		\a[34] ,
		_w4558_
	);
	LUT2 #(
		.INIT('h8)
	) name4493 (
		\a[32] ,
		\a[34] ,
		_w4559_
	);
	LUT4 #(
		.INIT('h8000)
	) name4494 (
		\a[31] ,
		\a[32] ,
		\a[33] ,
		\a[34] ,
		_w4560_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4495 (
		\a[31] ,
		\a[32] ,
		\a[33] ,
		\a[34] ,
		_w4561_
	);
	LUT4 #(
		.INIT('h0660)
	) name4496 (
		_w4424_,
		_w4556_,
		_w4557_,
		_w4561_,
		_w4562_
	);
	LUT4 #(
		.INIT('h9009)
	) name4497 (
		_w4424_,
		_w4556_,
		_w4557_,
		_w4561_,
		_w4563_
	);
	LUT4 #(
		.INIT('h6996)
	) name4498 (
		_w4424_,
		_w4556_,
		_w4557_,
		_w4561_,
		_w4564_
	);
	LUT2 #(
		.INIT('h8)
	) name4499 (
		\a[17] ,
		\a[48] ,
		_w4565_
	);
	LUT2 #(
		.INIT('h8)
	) name4500 (
		\a[3] ,
		\a[62] ,
		_w4566_
	);
	LUT3 #(
		.INIT('h6c)
	) name4501 (
		\a[3] ,
		\a[33] ,
		\a[62] ,
		_w4567_
	);
	LUT2 #(
		.INIT('h6)
	) name4502 (
		_w4565_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h6)
	) name4503 (
		_w4564_,
		_w4568_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name4504 (
		\a[23] ,
		\a[42] ,
		_w4570_
	);
	LUT4 #(
		.INIT('h153f)
	) name4505 (
		\a[24] ,
		\a[25] ,
		\a[40] ,
		\a[41] ,
		_w4571_
	);
	LUT4 #(
		.INIT('h8000)
	) name4506 (
		\a[24] ,
		\a[25] ,
		\a[40] ,
		\a[41] ,
		_w4572_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4507 (
		\a[24] ,
		\a[25] ,
		\a[40] ,
		\a[41] ,
		_w4573_
	);
	LUT2 #(
		.INIT('h8)
	) name4508 (
		\a[9] ,
		\a[56] ,
		_w4574_
	);
	LUT4 #(
		.INIT('h153f)
	) name4509 (
		\a[10] ,
		\a[20] ,
		\a[45] ,
		\a[55] ,
		_w4575_
	);
	LUT4 #(
		.INIT('h8000)
	) name4510 (
		\a[10] ,
		\a[20] ,
		\a[45] ,
		\a[55] ,
		_w4576_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4511 (
		\a[10] ,
		\a[20] ,
		\a[45] ,
		\a[55] ,
		_w4577_
	);
	LUT4 #(
		.INIT('h0660)
	) name4512 (
		_w4570_,
		_w4573_,
		_w4574_,
		_w4577_,
		_w4578_
	);
	LUT4 #(
		.INIT('h9009)
	) name4513 (
		_w4570_,
		_w4573_,
		_w4574_,
		_w4577_,
		_w4579_
	);
	LUT4 #(
		.INIT('h6996)
	) name4514 (
		_w4570_,
		_w4573_,
		_w4574_,
		_w4577_,
		_w4580_
	);
	LUT2 #(
		.INIT('h8)
	) name4515 (
		\a[26] ,
		\a[39] ,
		_w4581_
	);
	LUT4 #(
		.INIT('h153f)
	) name4516 (
		\a[27] ,
		\a[28] ,
		\a[37] ,
		\a[38] ,
		_w4582_
	);
	LUT4 #(
		.INIT('h8000)
	) name4517 (
		\a[27] ,
		\a[28] ,
		\a[37] ,
		\a[38] ,
		_w4583_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4518 (
		\a[27] ,
		\a[28] ,
		\a[37] ,
		\a[38] ,
		_w4584_
	);
	LUT2 #(
		.INIT('h6)
	) name4519 (
		_w4581_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h6)
	) name4520 (
		_w4580_,
		_w4585_,
		_w4586_
	);
	LUT3 #(
		.INIT('h96)
	) name4521 (
		_w4553_,
		_w4569_,
		_w4586_,
		_w4587_
	);
	LUT4 #(
		.INIT('he800)
	) name4522 (
		_w4353_,
		_w4354_,
		_w4364_,
		_w4587_,
		_w4588_
	);
	LUT3 #(
		.INIT('h96)
	) name4523 (
		_w4539_,
		_w4542_,
		_w4587_,
		_w4589_
	);
	LUT4 #(
		.INIT('h4114)
	) name4524 (
		_w4532_,
		_w4539_,
		_w4542_,
		_w4587_,
		_w4590_
	);
	LUT4 #(
		.INIT('h8e00)
	) name4525 (
		_w4350_,
		_w4366_,
		_w4370_,
		_w4590_,
		_w4591_
	);
	LUT4 #(
		.INIT('h8228)
	) name4526 (
		_w4532_,
		_w4539_,
		_w4542_,
		_w4587_,
		_w4592_
	);
	LUT4 #(
		.INIT('h7100)
	) name4527 (
		_w4350_,
		_w4366_,
		_w4370_,
		_w4592_,
		_w4593_
	);
	LUT3 #(
		.INIT('h96)
	) name4528 (
		_w4504_,
		_w4532_,
		_w4589_,
		_w4594_
	);
	LUT3 #(
		.INIT('he1)
	) name4529 (
		_w4502_,
		_w4503_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h8)
	) name4530 (
		_w4478_,
		_w4595_,
		_w4596_
	);
	LUT2 #(
		.INIT('h6)
	) name4531 (
		_w4478_,
		_w4595_,
		_w4597_
	);
	LUT4 #(
		.INIT('h7707)
	) name4532 (
		_w4221_,
		_w4342_,
		_w4468_,
		_w4469_,
		_w4598_
	);
	LUT4 #(
		.INIT('h1101)
	) name4533 (
		_w4221_,
		_w4342_,
		_w4468_,
		_w4469_,
		_w4599_
	);
	LUT2 #(
		.INIT('h4)
	) name4534 (
		_w4214_,
		_w4598_,
		_w4600_
	);
	LUT4 #(
		.INIT('h040f)
	) name4535 (
		_w4078_,
		_w4220_,
		_w4599_,
		_w4600_,
		_w4601_
	);
	LUT3 #(
		.INIT('h9c)
	) name4536 (
		_w4470_,
		_w4597_,
		_w4601_,
		_w4602_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name4537 (
		_w4468_,
		_w4469_,
		_w4478_,
		_w4595_,
		_w4603_
	);
	LUT3 #(
		.INIT('hb2)
	) name4538 (
		_w4481_,
		_w4484_,
		_w4500_,
		_w4604_
	);
	LUT2 #(
		.INIT('h8)
	) name4539 (
		\a[23] ,
		\a[43] ,
		_w4605_
	);
	LUT4 #(
		.INIT('h153f)
	) name4540 (
		\a[9] ,
		\a[24] ,
		\a[42] ,
		\a[57] ,
		_w4606_
	);
	LUT2 #(
		.INIT('h8)
	) name4541 (
		\a[24] ,
		\a[57] ,
		_w4607_
	);
	LUT4 #(
		.INIT('h8000)
	) name4542 (
		\a[9] ,
		\a[24] ,
		\a[42] ,
		\a[57] ,
		_w4608_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4543 (
		\a[9] ,
		\a[24] ,
		\a[42] ,
		\a[57] ,
		_w4609_
	);
	LUT2 #(
		.INIT('h8)
	) name4544 (
		\a[20] ,
		\a[46] ,
		_w4610_
	);
	LUT4 #(
		.INIT('h153f)
	) name4545 (
		\a[21] ,
		\a[22] ,
		\a[44] ,
		\a[45] ,
		_w4611_
	);
	LUT2 #(
		.INIT('h8)
	) name4546 (
		\a[22] ,
		\a[45] ,
		_w4612_
	);
	LUT4 #(
		.INIT('h8000)
	) name4547 (
		\a[21] ,
		\a[22] ,
		\a[44] ,
		\a[45] ,
		_w4613_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4548 (
		\a[21] ,
		\a[22] ,
		\a[44] ,
		\a[45] ,
		_w4614_
	);
	LUT4 #(
		.INIT('h0660)
	) name4549 (
		_w4605_,
		_w4609_,
		_w4610_,
		_w4614_,
		_w4615_
	);
	LUT4 #(
		.INIT('h9009)
	) name4550 (
		_w4605_,
		_w4609_,
		_w4610_,
		_w4614_,
		_w4616_
	);
	LUT4 #(
		.INIT('h6996)
	) name4551 (
		_w4605_,
		_w4609_,
		_w4610_,
		_w4614_,
		_w4617_
	);
	LUT2 #(
		.INIT('h8)
	) name4552 (
		\a[10] ,
		\a[56] ,
		_w4618_
	);
	LUT4 #(
		.INIT('h153f)
	) name4553 (
		\a[25] ,
		\a[26] ,
		\a[40] ,
		\a[41] ,
		_w4619_
	);
	LUT4 #(
		.INIT('h8000)
	) name4554 (
		\a[25] ,
		\a[26] ,
		\a[40] ,
		\a[41] ,
		_w4620_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4555 (
		\a[25] ,
		\a[26] ,
		\a[40] ,
		\a[41] ,
		_w4621_
	);
	LUT2 #(
		.INIT('h6)
	) name4556 (
		_w4618_,
		_w4621_,
		_w4622_
	);
	LUT2 #(
		.INIT('h8)
	) name4557 (
		\a[18] ,
		\a[48] ,
		_w4623_
	);
	LUT4 #(
		.INIT('h153f)
	) name4558 (
		\a[13] ,
		\a[15] ,
		\a[51] ,
		\a[53] ,
		_w4624_
	);
	LUT4 #(
		.INIT('h8000)
	) name4559 (
		\a[13] ,
		\a[15] ,
		\a[51] ,
		\a[53] ,
		_w4625_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4560 (
		\a[13] ,
		\a[15] ,
		\a[51] ,
		\a[53] ,
		_w4626_
	);
	LUT2 #(
		.INIT('h8)
	) name4561 (
		\a[14] ,
		\a[52] ,
		_w4627_
	);
	LUT4 #(
		.INIT('h153f)
	) name4562 (
		\a[30] ,
		\a[31] ,
		\a[35] ,
		\a[36] ,
		_w4628_
	);
	LUT2 #(
		.INIT('h8)
	) name4563 (
		\a[31] ,
		\a[36] ,
		_w4629_
	);
	LUT4 #(
		.INIT('h8000)
	) name4564 (
		\a[30] ,
		\a[31] ,
		\a[35] ,
		\a[36] ,
		_w4630_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4565 (
		\a[30] ,
		\a[31] ,
		\a[35] ,
		\a[36] ,
		_w4631_
	);
	LUT4 #(
		.INIT('h0660)
	) name4566 (
		_w4623_,
		_w4626_,
		_w4627_,
		_w4631_,
		_w4632_
	);
	LUT4 #(
		.INIT('h9009)
	) name4567 (
		_w4623_,
		_w4626_,
		_w4627_,
		_w4631_,
		_w4633_
	);
	LUT4 #(
		.INIT('h6996)
	) name4568 (
		_w4623_,
		_w4626_,
		_w4627_,
		_w4631_,
		_w4634_
	);
	LUT4 #(
		.INIT('h153f)
	) name4569 (
		\a[16] ,
		\a[17] ,
		\a[49] ,
		\a[50] ,
		_w4635_
	);
	LUT4 #(
		.INIT('h8000)
	) name4570 (
		\a[16] ,
		\a[17] ,
		\a[49] ,
		\a[50] ,
		_w4636_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4571 (
		\a[16] ,
		\a[17] ,
		\a[49] ,
		\a[50] ,
		_w4637_
	);
	LUT2 #(
		.INIT('h6)
	) name4572 (
		_w4559_,
		_w4637_,
		_w4638_
	);
	LUT4 #(
		.INIT('h0660)
	) name4573 (
		_w4617_,
		_w4622_,
		_w4634_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h9009)
	) name4574 (
		_w4617_,
		_w4622_,
		_w4634_,
		_w4638_,
		_w4640_
	);
	LUT4 #(
		.INIT('h6996)
	) name4575 (
		_w4617_,
		_w4622_,
		_w4634_,
		_w4638_,
		_w4641_
	);
	LUT2 #(
		.INIT('h8)
	) name4576 (
		\a[3] ,
		\a[63] ,
		_w4642_
	);
	LUT4 #(
		.INIT('h153f)
	) name4577 (
		\a[4] ,
		\a[5] ,
		\a[61] ,
		\a[62] ,
		_w4643_
	);
	LUT4 #(
		.INIT('h8000)
	) name4578 (
		\a[4] ,
		\a[5] ,
		\a[61] ,
		\a[62] ,
		_w4644_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4579 (
		\a[4] ,
		\a[5] ,
		\a[61] ,
		\a[62] ,
		_w4645_
	);
	LUT2 #(
		.INIT('h8)
	) name4580 (
		\a[27] ,
		\a[39] ,
		_w4646_
	);
	LUT4 #(
		.INIT('h153f)
	) name4581 (
		\a[28] ,
		\a[29] ,
		\a[37] ,
		\a[38] ,
		_w4647_
	);
	LUT2 #(
		.INIT('h8)
	) name4582 (
		\a[29] ,
		\a[38] ,
		_w4648_
	);
	LUT4 #(
		.INIT('h8000)
	) name4583 (
		\a[28] ,
		\a[29] ,
		\a[37] ,
		\a[38] ,
		_w4649_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4584 (
		\a[28] ,
		\a[29] ,
		\a[37] ,
		\a[38] ,
		_w4650_
	);
	LUT4 #(
		.INIT('h0660)
	) name4585 (
		_w4642_,
		_w4645_,
		_w4646_,
		_w4650_,
		_w4651_
	);
	LUT4 #(
		.INIT('h9009)
	) name4586 (
		_w4642_,
		_w4645_,
		_w4646_,
		_w4650_,
		_w4652_
	);
	LUT4 #(
		.INIT('h6996)
	) name4587 (
		_w4642_,
		_w4645_,
		_w4646_,
		_w4650_,
		_w4653_
	);
	LUT2 #(
		.INIT('h8)
	) name4588 (
		\a[11] ,
		\a[55] ,
		_w4654_
	);
	LUT4 #(
		.INIT('h153f)
	) name4589 (
		\a[12] ,
		\a[19] ,
		\a[47] ,
		\a[54] ,
		_w4655_
	);
	LUT4 #(
		.INIT('h8000)
	) name4590 (
		\a[12] ,
		\a[19] ,
		\a[47] ,
		\a[54] ,
		_w4656_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4591 (
		\a[12] ,
		\a[19] ,
		\a[47] ,
		\a[54] ,
		_w4657_
	);
	LUT2 #(
		.INIT('h6)
	) name4592 (
		_w4654_,
		_w4657_,
		_w4658_
	);
	LUT2 #(
		.INIT('h6)
	) name4593 (
		_w4653_,
		_w4658_,
		_w4659_
	);
	LUT2 #(
		.INIT('h6)
	) name4594 (
		_w4641_,
		_w4659_,
		_w4660_
	);
	LUT4 #(
		.INIT('h002b)
	) name4595 (
		_w4488_,
		_w4489_,
		_w4499_,
		_w4660_,
		_w4661_
	);
	LUT3 #(
		.INIT('h2b)
	) name4596 (
		_w4491_,
		_w4492_,
		_w4493_,
		_w4662_
	);
	LUT3 #(
		.INIT('h17)
	) name4597 (
		_w4495_,
		_w4496_,
		_w4497_,
		_w4663_
	);
	LUT3 #(
		.INIT('h17)
	) name4598 (
		_w4525_,
		_w4526_,
		_w4527_,
		_w4664_
	);
	LUT3 #(
		.INIT('h96)
	) name4599 (
		_w4662_,
		_w4663_,
		_w4664_,
		_w4665_
	);
	LUT3 #(
		.INIT('h2b)
	) name4600 (
		_w4490_,
		_w4494_,
		_w4498_,
		_w4666_
	);
	LUT3 #(
		.INIT('hd4)
	) name4601 (
		_w4528_,
		_w4529_,
		_w4530_,
		_w4667_
	);
	LUT3 #(
		.INIT('h96)
	) name4602 (
		_w4665_,
		_w4666_,
		_w4667_,
		_w4668_
	);
	LUT4 #(
		.INIT('h2882)
	) name4603 (
		_w4660_,
		_w4665_,
		_w4666_,
		_w4667_,
		_w4669_
	);
	LUT4 #(
		.INIT('hd400)
	) name4604 (
		_w4488_,
		_w4489_,
		_w4499_,
		_w4669_,
		_w4670_
	);
	LUT3 #(
		.INIT('h0d)
	) name4605 (
		_w4661_,
		_w4668_,
		_w4670_,
		_w4671_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4606 (
		_w4365_,
		_w4540_,
		_w4541_,
		_w4587_,
		_w4672_
	);
	LUT3 #(
		.INIT('h0e)
	) name4607 (
		_w4539_,
		_w4588_,
		_w4672_,
		_w4673_
	);
	LUT4 #(
		.INIT('hd400)
	) name4608 (
		_w4488_,
		_w4489_,
		_w4499_,
		_w4660_,
		_w4674_
	);
	LUT3 #(
		.INIT('h04)
	) name4609 (
		_w4661_,
		_w4668_,
		_w4674_,
		_w4675_
	);
	LUT3 #(
		.INIT('h08)
	) name4610 (
		_w4671_,
		_w4673_,
		_w4675_,
		_w4676_
	);
	LUT3 #(
		.INIT('h02)
	) name4611 (
		_w4671_,
		_w4673_,
		_w4675_,
		_w4677_
	);
	LUT3 #(
		.INIT('h1b)
	) name4612 (
		_w4604_,
		_w4676_,
		_w4677_,
		_w4678_
	);
	LUT4 #(
		.INIT('h5a96)
	) name4613 (
		_w4604_,
		_w4671_,
		_w4673_,
		_w4675_,
		_w4679_
	);
	LUT4 #(
		.INIT('hf100)
	) name4614 (
		_w4278_,
		_w4349_,
		_w4366_,
		_w4532_,
		_w4680_
	);
	LUT3 #(
		.INIT('hb0)
	) name4615 (
		_w4367_,
		_w4370_,
		_w4680_,
		_w4681_
	);
	LUT3 #(
		.INIT('he8)
	) name4616 (
		_w4536_,
		_w4537_,
		_w4538_,
		_w4682_
	);
	LUT3 #(
		.INIT('he8)
	) name4617 (
		_w4533_,
		_w4534_,
		_w4535_,
		_w4683_
	);
	LUT3 #(
		.INIT('h0d)
	) name4618 (
		_w4511_,
		_w4518_,
		_w4519_,
		_w4684_
	);
	LUT4 #(
		.INIT('h153f)
	) name4619 (
		\a[2] ,
		\a[4] ,
		\a[61] ,
		\a[63] ,
		_w4685_
	);
	LUT4 #(
		.INIT('h000d)
	) name4620 (
		_w4430_,
		_w4431_,
		_w4432_,
		_w4509_,
		_w4686_
	);
	LUT3 #(
		.INIT('h0d)
	) name4621 (
		_w4581_,
		_w4582_,
		_w4583_,
		_w4687_
	);
	LUT2 #(
		.INIT('h8)
	) name4622 (
		\a[6] ,
		\a[60] ,
		_w4688_
	);
	LUT4 #(
		.INIT('h153f)
	) name4623 (
		\a[7] ,
		\a[8] ,
		\a[58] ,
		\a[59] ,
		_w4689_
	);
	LUT4 #(
		.INIT('h8000)
	) name4624 (
		\a[7] ,
		\a[8] ,
		\a[58] ,
		\a[59] ,
		_w4690_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4625 (
		\a[7] ,
		\a[8] ,
		\a[58] ,
		\a[59] ,
		_w4691_
	);
	LUT2 #(
		.INIT('h6)
	) name4626 (
		_w4688_,
		_w4691_,
		_w4692_
	);
	LUT4 #(
		.INIT('he11e)
	) name4627 (
		_w4685_,
		_w4686_,
		_w4687_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		_w4684_,
		_w4693_,
		_w4694_
	);
	LUT2 #(
		.INIT('h1)
	) name4629 (
		_w4684_,
		_w4693_,
		_w4695_
	);
	LUT2 #(
		.INIT('h6)
	) name4630 (
		_w4684_,
		_w4693_,
		_w4696_
	);
	LUT3 #(
		.INIT('h0d)
	) name4631 (
		_w4557_,
		_w4558_,
		_w4560_,
		_w4697_
	);
	LUT3 #(
		.INIT('he8)
	) name4632 (
		\a[33] ,
		_w4565_,
		_w4566_,
		_w4698_
	);
	LUT3 #(
		.INIT('h0d)
	) name4633 (
		_w3535_,
		_w4512_,
		_w4513_,
		_w4699_
	);
	LUT3 #(
		.INIT('h69)
	) name4634 (
		_w4697_,
		_w4698_,
		_w4699_,
		_w4700_
	);
	LUT3 #(
		.INIT('h32)
	) name4635 (
		_w4424_,
		_w4554_,
		_w4555_,
		_w4701_
	);
	LUT3 #(
		.INIT('h0d)
	) name4636 (
		_w4543_,
		_w4544_,
		_w4545_,
		_w4702_
	);
	LUT3 #(
		.INIT('h0d)
	) name4637 (
		_w4548_,
		_w4549_,
		_w4550_,
		_w4703_
	);
	LUT3 #(
		.INIT('h96)
	) name4638 (
		_w4701_,
		_w4702_,
		_w4703_,
		_w4704_
	);
	LUT3 #(
		.INIT('h32)
	) name4639 (
		_w4562_,
		_w4563_,
		_w4568_,
		_w4705_
	);
	LUT3 #(
		.INIT('h69)
	) name4640 (
		_w4700_,
		_w4704_,
		_w4705_,
		_w4706_
	);
	LUT3 #(
		.INIT('h60)
	) name4641 (
		_w4683_,
		_w4696_,
		_w4706_,
		_w4707_
	);
	LUT3 #(
		.INIT('h09)
	) name4642 (
		_w4683_,
		_w4696_,
		_w4706_,
		_w4708_
	);
	LUT3 #(
		.INIT('h96)
	) name4643 (
		_w4683_,
		_w4696_,
		_w4706_,
		_w4709_
	);
	LUT2 #(
		.INIT('h6)
	) name4644 (
		_w4682_,
		_w4709_,
		_w4710_
	);
	LUT4 #(
		.INIT('he0fe)
	) name4645 (
		_w4462_,
		_w4505_,
		_w4524_,
		_w4531_,
		_w4711_
	);
	LUT2 #(
		.INIT('h2)
	) name4646 (
		_w4521_,
		_w4522_,
		_w4712_
	);
	LUT2 #(
		.INIT('h8)
	) name4647 (
		_w4521_,
		_w4522_,
		_w4713_
	);
	LUT4 #(
		.INIT('he800)
	) name4648 (
		_w4456_,
		_w4457_,
		_w4458_,
		_w4522_,
		_w4714_
	);
	LUT4 #(
		.INIT('h0027)
	) name4649 (
		_w4507_,
		_w4712_,
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT4 #(
		.INIT('h011f)
	) name4650 (
		_w4381_,
		_w4384_,
		_w4547_,
		_w4552_,
		_w4716_
	);
	LUT3 #(
		.INIT('h32)
	) name4651 (
		_w4387_,
		_w4515_,
		_w4516_,
		_w4717_
	);
	LUT3 #(
		.INIT('h32)
	) name4652 (
		_w4574_,
		_w4575_,
		_w4576_,
		_w4718_
	);
	LUT3 #(
		.INIT('h0d)
	) name4653 (
		_w4570_,
		_w4571_,
		_w4572_,
		_w4719_
	);
	LUT3 #(
		.INIT('h96)
	) name4654 (
		_w4717_,
		_w4718_,
		_w4719_,
		_w4720_
	);
	LUT3 #(
		.INIT('h32)
	) name4655 (
		_w4578_,
		_w4579_,
		_w4585_,
		_w4721_
	);
	LUT3 #(
		.INIT('h96)
	) name4656 (
		_w4716_,
		_w4720_,
		_w4721_,
		_w4722_
	);
	LUT3 #(
		.INIT('he8)
	) name4657 (
		_w4553_,
		_w4569_,
		_w4586_,
		_w4723_
	);
	LUT3 #(
		.INIT('h69)
	) name4658 (
		_w4715_,
		_w4722_,
		_w4723_,
		_w4724_
	);
	LUT3 #(
		.INIT('h69)
	) name4659 (
		_w4710_,
		_w4711_,
		_w4724_,
		_w4725_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4660 (
		_w4591_,
		_w4593_,
		_w4681_,
		_w4725_,
		_w4726_
	);
	LUT4 #(
		.INIT('h004f)
	) name4661 (
		_w4367_,
		_w4370_,
		_w4680_,
		_w4725_,
		_w4727_
	);
	LUT3 #(
		.INIT('h10)
	) name4662 (
		_w4591_,
		_w4593_,
		_w4727_,
		_w4728_
	);
	LUT4 #(
		.INIT('h01fe)
	) name4663 (
		_w4591_,
		_w4593_,
		_w4681_,
		_w4725_,
		_w4729_
	);
	LUT2 #(
		.INIT('h1)
	) name4664 (
		_w4679_,
		_w4729_,
		_w4730_
	);
	LUT3 #(
		.INIT('h45)
	) name4665 (
		_w4502_,
		_w4503_,
		_w4594_,
		_w4731_
	);
	LUT3 #(
		.INIT('h02)
	) name4666 (
		_w4679_,
		_w4726_,
		_w4728_,
		_w4732_
	);
	LUT3 #(
		.INIT('h01)
	) name4667 (
		_w4730_,
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT3 #(
		.INIT('ha9)
	) name4668 (
		_w4679_,
		_w4726_,
		_w4728_,
		_w4734_
	);
	LUT2 #(
		.INIT('h2)
	) name4669 (
		_w4731_,
		_w4734_,
		_w4735_
	);
	LUT3 #(
		.INIT('h36)
	) name4670 (
		_w4730_,
		_w4731_,
		_w4732_,
		_w4736_
	);
	LUT4 #(
		.INIT('h15ea)
	) name4671 (
		_w4596_,
		_w4601_,
		_w4603_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h1)
	) name4672 (
		_w4596_,
		_w4733_,
		_w4738_
	);
	LUT3 #(
		.INIT('hb2)
	) name4673 (
		_w4710_,
		_w4711_,
		_w4724_,
		_w4739_
	);
	LUT3 #(
		.INIT('h0b)
	) name4674 (
		_w4661_,
		_w4668_,
		_w4674_,
		_w4740_
	);
	LUT3 #(
		.INIT('h2b)
	) name4675 (
		_w4715_,
		_w4722_,
		_w4723_,
		_w4741_
	);
	LUT2 #(
		.INIT('h8)
	) name4676 (
		\a[25] ,
		\a[42] ,
		_w4742_
	);
	LUT4 #(
		.INIT('h153f)
	) name4677 (
		\a[21] ,
		\a[26] ,
		\a[41] ,
		\a[46] ,
		_w4743_
	);
	LUT4 #(
		.INIT('h8000)
	) name4678 (
		\a[21] ,
		\a[26] ,
		\a[41] ,
		\a[46] ,
		_w4744_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4679 (
		\a[21] ,
		\a[26] ,
		\a[41] ,
		\a[46] ,
		_w4745_
	);
	LUT2 #(
		.INIT('h8)
	) name4680 (
		\a[19] ,
		\a[48] ,
		_w4746_
	);
	LUT4 #(
		.INIT('h153f)
	) name4681 (
		\a[14] ,
		\a[17] ,
		\a[50] ,
		\a[53] ,
		_w4747_
	);
	LUT4 #(
		.INIT('h8000)
	) name4682 (
		\a[14] ,
		\a[17] ,
		\a[50] ,
		\a[53] ,
		_w4748_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4683 (
		\a[14] ,
		\a[17] ,
		\a[50] ,
		\a[53] ,
		_w4749_
	);
	LUT4 #(
		.INIT('h0660)
	) name4684 (
		_w4742_,
		_w4745_,
		_w4746_,
		_w4749_,
		_w4750_
	);
	LUT4 #(
		.INIT('h9009)
	) name4685 (
		_w4742_,
		_w4745_,
		_w4746_,
		_w4749_,
		_w4751_
	);
	LUT4 #(
		.INIT('h6996)
	) name4686 (
		_w4742_,
		_w4745_,
		_w4746_,
		_w4749_,
		_w4752_
	);
	LUT4 #(
		.INIT('h153f)
	) name4687 (
		\a[27] ,
		\a[28] ,
		\a[39] ,
		\a[40] ,
		_w4753_
	);
	LUT4 #(
		.INIT('h8000)
	) name4688 (
		\a[27] ,
		\a[28] ,
		\a[39] ,
		\a[40] ,
		_w4754_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4689 (
		\a[27] ,
		\a[28] ,
		\a[39] ,
		\a[40] ,
		_w4755_
	);
	LUT2 #(
		.INIT('h6)
	) name4690 (
		_w4508_,
		_w4755_,
		_w4756_
	);
	LUT2 #(
		.INIT('h6)
	) name4691 (
		_w4752_,
		_w4756_,
		_w4757_
	);
	LUT4 #(
		.INIT('h153f)
	) name4692 (
		\a[32] ,
		\a[33] ,
		\a[34] ,
		\a[35] ,
		_w4758_
	);
	LUT2 #(
		.INIT('h8)
	) name4693 (
		\a[33] ,
		\a[35] ,
		_w4759_
	);
	LUT4 #(
		.INIT('h8000)
	) name4694 (
		\a[32] ,
		\a[33] ,
		\a[34] ,
		\a[35] ,
		_w4760_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4695 (
		\a[32] ,
		\a[33] ,
		\a[34] ,
		\a[35] ,
		_w4761_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		\a[18] ,
		\a[49] ,
		_w4762_
	);
	LUT3 #(
		.INIT('h13)
	) name4697 (
		\a[5] ,
		\a[34] ,
		\a[62] ,
		_w4763_
	);
	LUT3 #(
		.INIT('h80)
	) name4698 (
		\a[5] ,
		\a[34] ,
		\a[62] ,
		_w4764_
	);
	LUT3 #(
		.INIT('h6c)
	) name4699 (
		\a[5] ,
		\a[34] ,
		\a[62] ,
		_w4765_
	);
	LUT4 #(
		.INIT('h0660)
	) name4700 (
		_w4629_,
		_w4761_,
		_w4762_,
		_w4765_,
		_w4766_
	);
	LUT4 #(
		.INIT('h9009)
	) name4701 (
		_w4629_,
		_w4761_,
		_w4762_,
		_w4765_,
		_w4767_
	);
	LUT4 #(
		.INIT('h6996)
	) name4702 (
		_w4629_,
		_w4761_,
		_w4762_,
		_w4765_,
		_w4768_
	);
	LUT4 #(
		.INIT('h153f)
	) name4703 (
		\a[12] ,
		\a[13] ,
		\a[54] ,
		\a[55] ,
		_w4769_
	);
	LUT4 #(
		.INIT('h8000)
	) name4704 (
		\a[12] ,
		\a[13] ,
		\a[54] ,
		\a[55] ,
		_w4770_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4705 (
		\a[12] ,
		\a[13] ,
		\a[54] ,
		\a[55] ,
		_w4771_
	);
	LUT2 #(
		.INIT('h6)
	) name4706 (
		_w4648_,
		_w4771_,
		_w4772_
	);
	LUT2 #(
		.INIT('h8)
	) name4707 (
		\a[7] ,
		\a[60] ,
		_w4773_
	);
	LUT4 #(
		.INIT('h153f)
	) name4708 (
		\a[8] ,
		\a[9] ,
		\a[58] ,
		\a[59] ,
		_w4774_
	);
	LUT2 #(
		.INIT('h8)
	) name4709 (
		\a[9] ,
		\a[59] ,
		_w4775_
	);
	LUT4 #(
		.INIT('h8000)
	) name4710 (
		\a[8] ,
		\a[9] ,
		\a[58] ,
		\a[59] ,
		_w4776_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4711 (
		\a[8] ,
		\a[9] ,
		\a[58] ,
		\a[59] ,
		_w4777_
	);
	LUT4 #(
		.INIT('h153f)
	) name4712 (
		\a[23] ,
		\a[24] ,
		\a[43] ,
		\a[44] ,
		_w4778_
	);
	LUT2 #(
		.INIT('h8)
	) name4713 (
		\a[24] ,
		\a[44] ,
		_w4779_
	);
	LUT4 #(
		.INIT('h8000)
	) name4714 (
		\a[23] ,
		\a[24] ,
		\a[43] ,
		\a[44] ,
		_w4780_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4715 (
		\a[23] ,
		\a[24] ,
		\a[43] ,
		\a[44] ,
		_w4781_
	);
	LUT4 #(
		.INIT('h1428)
	) name4716 (
		_w4612_,
		_w4773_,
		_w4777_,
		_w4781_,
		_w4782_
	);
	LUT4 #(
		.INIT('h8241)
	) name4717 (
		_w4612_,
		_w4773_,
		_w4777_,
		_w4781_,
		_w4783_
	);
	LUT4 #(
		.INIT('h6996)
	) name4718 (
		_w4612_,
		_w4773_,
		_w4777_,
		_w4781_,
		_w4784_
	);
	LUT2 #(
		.INIT('h8)
	) name4719 (
		\a[15] ,
		\a[52] ,
		_w4785_
	);
	LUT4 #(
		.INIT('h153f)
	) name4720 (
		\a[16] ,
		\a[30] ,
		\a[37] ,
		\a[51] ,
		_w4786_
	);
	LUT4 #(
		.INIT('h8000)
	) name4721 (
		\a[16] ,
		\a[30] ,
		\a[37] ,
		\a[51] ,
		_w4787_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4722 (
		\a[16] ,
		\a[30] ,
		\a[37] ,
		\a[51] ,
		_w4788_
	);
	LUT2 #(
		.INIT('h6)
	) name4723 (
		_w4785_,
		_w4788_,
		_w4789_
	);
	LUT4 #(
		.INIT('h0660)
	) name4724 (
		_w4768_,
		_w4772_,
		_w4784_,
		_w4789_,
		_w4790_
	);
	LUT4 #(
		.INIT('h9009)
	) name4725 (
		_w4768_,
		_w4772_,
		_w4784_,
		_w4789_,
		_w4791_
	);
	LUT4 #(
		.INIT('h6996)
	) name4726 (
		_w4768_,
		_w4772_,
		_w4784_,
		_w4789_,
		_w4792_
	);
	LUT2 #(
		.INIT('h6)
	) name4727 (
		_w4757_,
		_w4792_,
		_w4793_
	);
	LUT4 #(
		.INIT('hd400)
	) name4728 (
		_w4715_,
		_w4722_,
		_w4723_,
		_w4793_,
		_w4794_
	);
	LUT4 #(
		.INIT('h002b)
	) name4729 (
		_w4715_,
		_w4722_,
		_w4723_,
		_w4793_,
		_w4795_
	);
	LUT3 #(
		.INIT('h8e)
	) name4730 (
		_w4716_,
		_w4720_,
		_w4721_,
		_w4796_
	);
	LUT3 #(
		.INIT('hd4)
	) name4731 (
		_w4700_,
		_w4704_,
		_w4705_,
		_w4797_
	);
	LUT3 #(
		.INIT('h2b)
	) name4732 (
		_w4701_,
		_w4702_,
		_w4703_,
		_w4798_
	);
	LUT3 #(
		.INIT('h8e)
	) name4733 (
		_w4717_,
		_w4718_,
		_w4719_,
		_w4799_
	);
	LUT3 #(
		.INIT('h4d)
	) name4734 (
		_w4697_,
		_w4698_,
		_w4699_,
		_w4800_
	);
	LUT3 #(
		.INIT('h96)
	) name4735 (
		_w4798_,
		_w4799_,
		_w4800_,
		_w4801_
	);
	LUT3 #(
		.INIT('h6f)
	) name4736 (
		_w4796_,
		_w4797_,
		_w4801_,
		_w4802_
	);
	LUT3 #(
		.INIT('h69)
	) name4737 (
		_w4796_,
		_w4797_,
		_w4801_,
		_w4803_
	);
	LUT4 #(
		.INIT('hf40b)
	) name4738 (
		_w4741_,
		_w4793_,
		_w4795_,
		_w4803_,
		_w4804_
	);
	LUT3 #(
		.INIT('h69)
	) name4739 (
		_w4739_,
		_w4740_,
		_w4804_,
		_w4805_
	);
	LUT4 #(
		.INIT('hb200)
	) name4740 (
		_w4481_,
		_w4484_,
		_w4500_,
		_w4673_,
		_w4806_
	);
	LUT3 #(
		.INIT('h0e)
	) name4741 (
		_w4682_,
		_w4707_,
		_w4708_,
		_w4807_
	);
	LUT3 #(
		.INIT('he8)
	) name4742 (
		_w4665_,
		_w4666_,
		_w4667_,
		_w4808_
	);
	LUT3 #(
		.INIT('h32)
	) name4743 (
		_w4615_,
		_w4616_,
		_w4622_,
		_w4809_
	);
	LUT4 #(
		.INIT('h1f01)
	) name4744 (
		_w4685_,
		_w4686_,
		_w4687_,
		_w4692_,
		_w4810_
	);
	LUT3 #(
		.INIT('h32)
	) name4745 (
		_w4651_,
		_w4652_,
		_w4658_,
		_w4811_
	);
	LUT3 #(
		.INIT('h96)
	) name4746 (
		_w4809_,
		_w4810_,
		_w4811_,
		_w4812_
	);
	LUT3 #(
		.INIT('h0d)
	) name4747 (
		_w4688_,
		_w4689_,
		_w4690_,
		_w4813_
	);
	LUT3 #(
		.INIT('h0d)
	) name4748 (
		_w4642_,
		_w4643_,
		_w4644_,
		_w4814_
	);
	LUT3 #(
		.INIT('h0d)
	) name4749 (
		_w4646_,
		_w4647_,
		_w4649_,
		_w4815_
	);
	LUT3 #(
		.INIT('h96)
	) name4750 (
		_w4813_,
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT3 #(
		.INIT('h0d)
	) name4751 (
		_w4618_,
		_w4619_,
		_w4620_,
		_w4817_
	);
	LUT3 #(
		.INIT('h0d)
	) name4752 (
		_w4605_,
		_w4606_,
		_w4608_,
		_w4818_
	);
	LUT3 #(
		.INIT('h0d)
	) name4753 (
		_w4610_,
		_w4611_,
		_w4613_,
		_w4819_
	);
	LUT3 #(
		.INIT('h96)
	) name4754 (
		_w4817_,
		_w4818_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h8)
	) name4755 (
		\a[6] ,
		\a[61] ,
		_w4821_
	);
	LUT4 #(
		.INIT('h0dff)
	) name4756 (
		_w4559_,
		_w4635_,
		_w4636_,
		_w4821_,
		_w4822_
	);
	LUT4 #(
		.INIT('h000d)
	) name4757 (
		_w4559_,
		_w4635_,
		_w4636_,
		_w4821_,
		_w4823_
	);
	LUT4 #(
		.INIT('h0df2)
	) name4758 (
		_w4559_,
		_w4635_,
		_w4636_,
		_w4821_,
		_w4824_
	);
	LUT3 #(
		.INIT('h0d)
	) name4759 (
		_w4627_,
		_w4628_,
		_w4630_,
		_w4825_
	);
	LUT2 #(
		.INIT('h6)
	) name4760 (
		_w4824_,
		_w4825_,
		_w4826_
	);
	LUT3 #(
		.INIT('h69)
	) name4761 (
		_w4816_,
		_w4820_,
		_w4826_,
		_w4827_
	);
	LUT2 #(
		.INIT('h8)
	) name4762 (
		_w4812_,
		_w4827_,
		_w4828_
	);
	LUT2 #(
		.INIT('h1)
	) name4763 (
		_w4812_,
		_w4827_,
		_w4829_
	);
	LUT2 #(
		.INIT('h6)
	) name4764 (
		_w4812_,
		_w4827_,
		_w4830_
	);
	LUT2 #(
		.INIT('h6)
	) name4765 (
		_w4808_,
		_w4830_,
		_w4831_
	);
	LUT3 #(
		.INIT('h32)
	) name4766 (
		_w4632_,
		_w4633_,
		_w4638_,
		_w4832_
	);
	LUT3 #(
		.INIT('h32)
	) name4767 (
		_w4654_,
		_w4655_,
		_w4656_,
		_w4833_
	);
	LUT3 #(
		.INIT('h0d)
	) name4768 (
		_w4623_,
		_w4624_,
		_w4625_,
		_w4834_
	);
	LUT2 #(
		.INIT('h8)
	) name4769 (
		\a[10] ,
		\a[57] ,
		_w4835_
	);
	LUT4 #(
		.INIT('h153f)
	) name4770 (
		\a[11] ,
		\a[20] ,
		\a[47] ,
		\a[56] ,
		_w4836_
	);
	LUT2 #(
		.INIT('h8)
	) name4771 (
		\a[20] ,
		\a[56] ,
		_w4837_
	);
	LUT4 #(
		.INIT('h8000)
	) name4772 (
		\a[11] ,
		\a[20] ,
		\a[47] ,
		\a[56] ,
		_w4838_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4773 (
		\a[11] ,
		\a[20] ,
		\a[47] ,
		\a[56] ,
		_w4839_
	);
	LUT2 #(
		.INIT('h6)
	) name4774 (
		_w4835_,
		_w4839_,
		_w4840_
	);
	LUT3 #(
		.INIT('h96)
	) name4775 (
		_w4833_,
		_w4834_,
		_w4840_,
		_w4841_
	);
	LUT2 #(
		.INIT('h4)
	) name4776 (
		_w4832_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h2)
	) name4777 (
		_w4832_,
		_w4841_,
		_w4843_
	);
	LUT2 #(
		.INIT('h9)
	) name4778 (
		_w4832_,
		_w4841_,
		_w4844_
	);
	LUT3 #(
		.INIT('he8)
	) name4779 (
		_w4662_,
		_w4663_,
		_w4664_,
		_w4845_
	);
	LUT2 #(
		.INIT('h6)
	) name4780 (
		_w4844_,
		_w4845_,
		_w4846_
	);
	LUT3 #(
		.INIT('h32)
	) name4781 (
		_w4639_,
		_w4640_,
		_w4659_,
		_w4847_
	);
	LUT4 #(
		.INIT('h0017)
	) name4782 (
		_w4683_,
		_w4684_,
		_w4693_,
		_w4847_,
		_w4848_
	);
	LUT4 #(
		.INIT('he800)
	) name4783 (
		_w4683_,
		_w4684_,
		_w4693_,
		_w4847_,
		_w4849_
	);
	LUT4 #(
		.INIT('hf10e)
	) name4784 (
		_w4683_,
		_w4694_,
		_w4695_,
		_w4847_,
		_w4850_
	);
	LUT2 #(
		.INIT('h6)
	) name4785 (
		_w4846_,
		_w4850_,
		_w4851_
	);
	LUT3 #(
		.INIT('h96)
	) name4786 (
		_w4807_,
		_w4831_,
		_w4851_,
		_w4852_
	);
	LUT4 #(
		.INIT('h3102)
	) name4787 (
		_w4678_,
		_w4805_,
		_w4806_,
		_w4852_,
		_w4853_
	);
	LUT3 #(
		.INIT('h31)
	) name4788 (
		_w4679_,
		_w4726_,
		_w4728_,
		_w4854_
	);
	LUT4 #(
		.INIT('h08c4)
	) name4789 (
		_w4678_,
		_w4805_,
		_w4806_,
		_w4852_,
		_w4855_
	);
	LUT3 #(
		.INIT('h01)
	) name4790 (
		_w4853_,
		_w4854_,
		_w4855_,
		_w4856_
	);
	LUT4 #(
		.INIT('hc639)
	) name4791 (
		_w4678_,
		_w4805_,
		_w4806_,
		_w4852_,
		_w4857_
	);
	LUT2 #(
		.INIT('h2)
	) name4792 (
		_w4854_,
		_w4857_,
		_w4858_
	);
	LUT3 #(
		.INIT('h36)
	) name4793 (
		_w4853_,
		_w4854_,
		_w4855_,
		_w4859_
	);
	LUT2 #(
		.INIT('h9)
	) name4794 (
		_w4735_,
		_w4859_,
		_w4860_
	);
	LUT4 #(
		.INIT('h8f00)
	) name4795 (
		_w4601_,
		_w4603_,
		_w4738_,
		_w4860_,
		_w4861_
	);
	LUT2 #(
		.INIT('hc)
	) name4796 (
		_w4735_,
		_w4859_,
		_w4862_
	);
	LUT4 #(
		.INIT('h7000)
	) name4797 (
		_w4601_,
		_w4603_,
		_w4738_,
		_w4862_,
		_w4863_
	);
	LUT2 #(
		.INIT('he)
	) name4798 (
		_w4861_,
		_w4863_,
		_w4864_
	);
	LUT3 #(
		.INIT('h01)
	) name4799 (
		_w4596_,
		_w4733_,
		_w4856_,
		_w4865_
	);
	LUT4 #(
		.INIT('h023b)
	) name4800 (
		_w4678_,
		_w4805_,
		_w4806_,
		_w4852_,
		_w4866_
	);
	LUT2 #(
		.INIT('h4)
	) name4801 (
		_w4796_,
		_w4797_,
		_w4867_
	);
	LUT3 #(
		.INIT('h2b)
	) name4802 (
		_w4796_,
		_w4797_,
		_w4801_,
		_w4868_
	);
	LUT3 #(
		.INIT('h32)
	) name4803 (
		_w4746_,
		_w4747_,
		_w4748_,
		_w4869_
	);
	LUT3 #(
		.INIT('h32)
	) name4804 (
		_w4742_,
		_w4743_,
		_w4744_,
		_w4870_
	);
	LUT3 #(
		.INIT('h0d)
	) name4805 (
		_w4648_,
		_w4769_,
		_w4770_,
		_w4871_
	);
	LUT3 #(
		.INIT('h96)
	) name4806 (
		_w4869_,
		_w4870_,
		_w4871_,
		_w4872_
	);
	LUT3 #(
		.INIT('h32)
	) name4807 (
		_w4750_,
		_w4751_,
		_w4756_,
		_w4873_
	);
	LUT3 #(
		.INIT('h32)
	) name4808 (
		_w4766_,
		_w4767_,
		_w4772_,
		_w4874_
	);
	LUT3 #(
		.INIT('h69)
	) name4809 (
		_w4872_,
		_w4873_,
		_w4874_,
		_w4875_
	);
	LUT3 #(
		.INIT('he8)
	) name4810 (
		_w4798_,
		_w4799_,
		_w4800_,
		_w4876_
	);
	LUT3 #(
		.INIT('h0d)
	) name4811 (
		_w4835_,
		_w4836_,
		_w4838_,
		_w4877_
	);
	LUT3 #(
		.INIT('h0d)
	) name4812 (
		_w4612_,
		_w4778_,
		_w4780_,
		_w4878_
	);
	LUT3 #(
		.INIT('h0d)
	) name4813 (
		_w4773_,
		_w4774_,
		_w4776_,
		_w4879_
	);
	LUT3 #(
		.INIT('h96)
	) name4814 (
		_w4877_,
		_w4878_,
		_w4879_,
		_w4880_
	);
	LUT3 #(
		.INIT('h0d)
	) name4815 (
		_w4508_,
		_w4753_,
		_w4754_,
		_w4881_
	);
	LUT3 #(
		.INIT('h0d)
	) name4816 (
		_w4629_,
		_w4758_,
		_w4760_,
		_w4882_
	);
	LUT3 #(
		.INIT('h32)
	) name4817 (
		_w4785_,
		_w4786_,
		_w4787_,
		_w4883_
	);
	LUT3 #(
		.INIT('h96)
	) name4818 (
		_w4881_,
		_w4882_,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h4)
	) name4819 (
		_w4880_,
		_w4884_,
		_w4885_
	);
	LUT2 #(
		.INIT('h2)
	) name4820 (
		_w4880_,
		_w4884_,
		_w4886_
	);
	LUT2 #(
		.INIT('h9)
	) name4821 (
		_w4880_,
		_w4884_,
		_w4887_
	);
	LUT3 #(
		.INIT('h28)
	) name4822 (
		_w4875_,
		_w4876_,
		_w4887_,
		_w4888_
	);
	LUT3 #(
		.INIT('h41)
	) name4823 (
		_w4875_,
		_w4876_,
		_w4887_,
		_w4889_
	);
	LUT3 #(
		.INIT('h96)
	) name4824 (
		_w4875_,
		_w4876_,
		_w4887_,
		_w4890_
	);
	LUT2 #(
		.INIT('h9)
	) name4825 (
		_w4868_,
		_w4890_,
		_w4891_
	);
	LUT3 #(
		.INIT('h0e)
	) name4826 (
		_w4757_,
		_w4790_,
		_w4791_,
		_w4892_
	);
	LUT3 #(
		.INIT('h17)
	) name4827 (
		_w4817_,
		_w4818_,
		_w4819_,
		_w4893_
	);
	LUT3 #(
		.INIT('h4d)
	) name4828 (
		_w4833_,
		_w4834_,
		_w4840_,
		_w4894_
	);
	LUT3 #(
		.INIT('h32)
	) name4829 (
		_w4782_,
		_w4783_,
		_w4789_,
		_w4895_
	);
	LUT3 #(
		.INIT('h69)
	) name4830 (
		_w4893_,
		_w4894_,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h8)
	) name4831 (
		\a[8] ,
		\a[61] ,
		_w4897_
	);
	LUT4 #(
		.INIT('h8000)
	) name4832 (
		\a[7] ,
		\a[8] ,
		\a[60] ,
		\a[61] ,
		_w4898_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4833 (
		\a[7] ,
		\a[8] ,
		\a[60] ,
		\a[61] ,
		_w4899_
	);
	LUT4 #(
		.INIT('hf20d)
	) name4834 (
		_w4762_,
		_w4763_,
		_w4764_,
		_w4899_,
		_w4900_
	);
	LUT4 #(
		.INIT('ha800)
	) name4835 (
		_w4822_,
		_w4823_,
		_w4825_,
		_w4900_,
		_w4901_
	);
	LUT4 #(
		.INIT('h0057)
	) name4836 (
		_w4822_,
		_w4823_,
		_w4825_,
		_w4900_,
		_w4902_
	);
	LUT4 #(
		.INIT('h07f8)
	) name4837 (
		_w4822_,
		_w4825_,
		_w4823_,
		_w4900_,
		_w4903_
	);
	LUT3 #(
		.INIT('h17)
	) name4838 (
		_w4813_,
		_w4814_,
		_w4815_,
		_w4904_
	);
	LUT2 #(
		.INIT('h6)
	) name4839 (
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT3 #(
		.INIT('h96)
	) name4840 (
		_w4892_,
		_w4896_,
		_w4905_,
		_w4906_
	);
	LUT4 #(
		.INIT('he800)
	) name4841 (
		_w4808_,
		_w4812_,
		_w4827_,
		_w4906_,
		_w4907_
	);
	LUT4 #(
		.INIT('h0017)
	) name4842 (
		_w4808_,
		_w4812_,
		_w4827_,
		_w4906_,
		_w4908_
	);
	LUT4 #(
		.INIT('h31ce)
	) name4843 (
		_w4808_,
		_w4828_,
		_w4829_,
		_w4906_,
		_w4909_
	);
	LUT2 #(
		.INIT('h6)
	) name4844 (
		_w4891_,
		_w4909_,
		_w4910_
	);
	LUT4 #(
		.INIT('hb200)
	) name4845 (
		_w4739_,
		_w4740_,
		_w4804_,
		_w4910_,
		_w4911_
	);
	LUT3 #(
		.INIT('he8)
	) name4846 (
		_w4807_,
		_w4831_,
		_w4851_,
		_w4912_
	);
	LUT3 #(
		.INIT('h45)
	) name4847 (
		_w4794_,
		_w4795_,
		_w4803_,
		_w4913_
	);
	LUT3 #(
		.INIT('h32)
	) name4848 (
		_w4846_,
		_w4848_,
		_w4849_,
		_w4914_
	);
	LUT3 #(
		.INIT('h17)
	) name4849 (
		_w4816_,
		_w4820_,
		_w4826_,
		_w4915_
	);
	LUT3 #(
		.INIT('he8)
	) name4850 (
		_w4809_,
		_w4810_,
		_w4811_,
		_w4916_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		_w4915_,
		_w4916_,
		_w4917_
	);
	LUT2 #(
		.INIT('h8)
	) name4852 (
		_w4915_,
		_w4916_,
		_w4918_
	);
	LUT2 #(
		.INIT('h6)
	) name4853 (
		_w4915_,
		_w4916_,
		_w4919_
	);
	LUT3 #(
		.INIT('h23)
	) name4854 (
		_w4842_,
		_w4843_,
		_w4845_,
		_w4920_
	);
	LUT4 #(
		.INIT('h153f)
	) name4855 (
		\a[18] ,
		\a[19] ,
		\a[49] ,
		\a[50] ,
		_w4921_
	);
	LUT2 #(
		.INIT('h8)
	) name4856 (
		\a[19] ,
		\a[50] ,
		_w4922_
	);
	LUT4 #(
		.INIT('h8000)
	) name4857 (
		\a[18] ,
		\a[19] ,
		\a[49] ,
		\a[50] ,
		_w4923_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4858 (
		\a[18] ,
		\a[19] ,
		\a[49] ,
		\a[50] ,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name4859 (
		\a[30] ,
		\a[38] ,
		_w4925_
	);
	LUT4 #(
		.INIT('h153f)
	) name4860 (
		\a[31] ,
		\a[32] ,
		\a[36] ,
		\a[37] ,
		_w4926_
	);
	LUT4 #(
		.INIT('h8000)
	) name4861 (
		\a[31] ,
		\a[32] ,
		\a[36] ,
		\a[37] ,
		_w4927_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4862 (
		\a[31] ,
		\a[32] ,
		\a[36] ,
		\a[37] ,
		_w4928_
	);
	LUT4 #(
		.INIT('h0660)
	) name4863 (
		_w4759_,
		_w4924_,
		_w4925_,
		_w4928_,
		_w4929_
	);
	LUT4 #(
		.INIT('h9009)
	) name4864 (
		_w4759_,
		_w4924_,
		_w4925_,
		_w4928_,
		_w4930_
	);
	LUT4 #(
		.INIT('h6996)
	) name4865 (
		_w4759_,
		_w4924_,
		_w4925_,
		_w4928_,
		_w4931_
	);
	LUT2 #(
		.INIT('h8)
	) name4866 (
		\a[12] ,
		\a[56] ,
		_w4932_
	);
	LUT4 #(
		.INIT('h153f)
	) name4867 (
		\a[13] ,
		\a[17] ,
		\a[51] ,
		\a[55] ,
		_w4933_
	);
	LUT4 #(
		.INIT('h8000)
	) name4868 (
		\a[13] ,
		\a[17] ,
		\a[51] ,
		\a[55] ,
		_w4934_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4869 (
		\a[13] ,
		\a[17] ,
		\a[51] ,
		\a[55] ,
		_w4935_
	);
	LUT2 #(
		.INIT('h6)
	) name4870 (
		_w4932_,
		_w4935_,
		_w4936_
	);
	LUT2 #(
		.INIT('h8)
	) name4871 (
		\a[14] ,
		\a[54] ,
		_w4937_
	);
	LUT4 #(
		.INIT('h153f)
	) name4872 (
		\a[15] ,
		\a[16] ,
		\a[52] ,
		\a[53] ,
		_w4938_
	);
	LUT4 #(
		.INIT('h8000)
	) name4873 (
		\a[15] ,
		\a[16] ,
		\a[52] ,
		\a[53] ,
		_w4939_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4874 (
		\a[15] ,
		\a[16] ,
		\a[52] ,
		\a[53] ,
		_w4940_
	);
	LUT2 #(
		.INIT('h8)
	) name4875 (
		\a[20] ,
		\a[48] ,
		_w4941_
	);
	LUT4 #(
		.INIT('h153f)
	) name4876 (
		\a[22] ,
		\a[23] ,
		\a[45] ,
		\a[46] ,
		_w4942_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		\a[23] ,
		\a[46] ,
		_w4943_
	);
	LUT4 #(
		.INIT('h8000)
	) name4878 (
		\a[22] ,
		\a[23] ,
		\a[45] ,
		\a[46] ,
		_w4944_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4879 (
		\a[22] ,
		\a[23] ,
		\a[45] ,
		\a[46] ,
		_w4945_
	);
	LUT4 #(
		.INIT('h0660)
	) name4880 (
		_w4937_,
		_w4940_,
		_w4941_,
		_w4945_,
		_w4946_
	);
	LUT4 #(
		.INIT('h9009)
	) name4881 (
		_w4937_,
		_w4940_,
		_w4941_,
		_w4945_,
		_w4947_
	);
	LUT4 #(
		.INIT('h6996)
	) name4882 (
		_w4937_,
		_w4940_,
		_w4941_,
		_w4945_,
		_w4948_
	);
	LUT4 #(
		.INIT('h153f)
	) name4883 (
		\a[25] ,
		\a[26] ,
		\a[42] ,
		\a[43] ,
		_w4949_
	);
	LUT4 #(
		.INIT('h8000)
	) name4884 (
		\a[25] ,
		\a[26] ,
		\a[42] ,
		\a[43] ,
		_w4950_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4885 (
		\a[25] ,
		\a[26] ,
		\a[42] ,
		\a[43] ,
		_w4951_
	);
	LUT2 #(
		.INIT('h6)
	) name4886 (
		_w4779_,
		_w4951_,
		_w4952_
	);
	LUT4 #(
		.INIT('h0660)
	) name4887 (
		_w4931_,
		_w4936_,
		_w4948_,
		_w4952_,
		_w4953_
	);
	LUT4 #(
		.INIT('h9009)
	) name4888 (
		_w4931_,
		_w4936_,
		_w4948_,
		_w4952_,
		_w4954_
	);
	LUT4 #(
		.INIT('h6996)
	) name4889 (
		_w4931_,
		_w4936_,
		_w4948_,
		_w4952_,
		_w4955_
	);
	LUT4 #(
		.INIT('h153f)
	) name4890 (
		\a[10] ,
		\a[11] ,
		\a[57] ,
		\a[58] ,
		_w4956_
	);
	LUT2 #(
		.INIT('h8)
	) name4891 (
		\a[11] ,
		\a[58] ,
		_w4957_
	);
	LUT4 #(
		.INIT('h8000)
	) name4892 (
		\a[10] ,
		\a[11] ,
		\a[57] ,
		\a[58] ,
		_w4958_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4893 (
		\a[10] ,
		\a[11] ,
		\a[57] ,
		\a[58] ,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name4894 (
		\a[27] ,
		\a[41] ,
		_w4960_
	);
	LUT4 #(
		.INIT('h153f)
	) name4895 (
		\a[28] ,
		\a[29] ,
		\a[39] ,
		\a[40] ,
		_w4961_
	);
	LUT4 #(
		.INIT('h8000)
	) name4896 (
		\a[28] ,
		\a[29] ,
		\a[39] ,
		\a[40] ,
		_w4962_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4897 (
		\a[28] ,
		\a[29] ,
		\a[39] ,
		\a[40] ,
		_w4963_
	);
	LUT4 #(
		.INIT('h0660)
	) name4898 (
		_w4775_,
		_w4959_,
		_w4960_,
		_w4963_,
		_w4964_
	);
	LUT4 #(
		.INIT('h9009)
	) name4899 (
		_w4775_,
		_w4959_,
		_w4960_,
		_w4963_,
		_w4965_
	);
	LUT4 #(
		.INIT('h6996)
	) name4900 (
		_w4775_,
		_w4959_,
		_w4960_,
		_w4963_,
		_w4966_
	);
	LUT2 #(
		.INIT('h8)
	) name4901 (
		\a[21] ,
		\a[47] ,
		_w4967_
	);
	LUT4 #(
		.INIT('h153f)
	) name4902 (
		\a[5] ,
		\a[6] ,
		\a[62] ,
		\a[63] ,
		_w4968_
	);
	LUT2 #(
		.INIT('h8)
	) name4903 (
		\a[6] ,
		\a[63] ,
		_w4969_
	);
	LUT4 #(
		.INIT('h8000)
	) name4904 (
		\a[5] ,
		\a[6] ,
		\a[62] ,
		\a[63] ,
		_w4970_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4905 (
		\a[5] ,
		\a[6] ,
		\a[62] ,
		\a[63] ,
		_w4971_
	);
	LUT2 #(
		.INIT('h6)
	) name4906 (
		_w4967_,
		_w4971_,
		_w4972_
	);
	LUT2 #(
		.INIT('h6)
	) name4907 (
		_w4966_,
		_w4972_,
		_w4973_
	);
	LUT2 #(
		.INIT('h6)
	) name4908 (
		_w4955_,
		_w4973_,
		_w4974_
	);
	LUT3 #(
		.INIT('h90)
	) name4909 (
		_w4919_,
		_w4920_,
		_w4974_,
		_w4975_
	);
	LUT3 #(
		.INIT('h06)
	) name4910 (
		_w4919_,
		_w4920_,
		_w4974_,
		_w4976_
	);
	LUT3 #(
		.INIT('h69)
	) name4911 (
		_w4919_,
		_w4920_,
		_w4974_,
		_w4977_
	);
	LUT2 #(
		.INIT('h6)
	) name4912 (
		_w4914_,
		_w4977_,
		_w4978_
	);
	LUT3 #(
		.INIT('h69)
	) name4913 (
		_w4912_,
		_w4913_,
		_w4978_,
		_w4979_
	);
	LUT4 #(
		.INIT('h004d)
	) name4914 (
		_w4739_,
		_w4740_,
		_w4804_,
		_w4910_,
		_w4980_
	);
	LUT3 #(
		.INIT('h04)
	) name4915 (
		_w4911_,
		_w4979_,
		_w4980_,
		_w4981_
	);
	LUT4 #(
		.INIT('h4db2)
	) name4916 (
		_w4739_,
		_w4740_,
		_w4804_,
		_w4910_,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name4917 (
		_w4979_,
		_w4982_,
		_w4983_
	);
	LUT3 #(
		.INIT('hc9)
	) name4918 (
		_w4911_,
		_w4979_,
		_w4980_,
		_w4984_
	);
	LUT3 #(
		.INIT('h01)
	) name4919 (
		_w4866_,
		_w4981_,
		_w4983_,
		_w4985_
	);
	LUT3 #(
		.INIT('h56)
	) name4920 (
		_w4866_,
		_w4981_,
		_w4983_,
		_w4986_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4921 (
		_w4735_,
		_w4856_,
		_w4858_,
		_w4986_,
		_w4987_
	);
	LUT4 #(
		.INIT('h8f00)
	) name4922 (
		_w4601_,
		_w4603_,
		_w4865_,
		_w4987_,
		_w4988_
	);
	LUT3 #(
		.INIT('h0d)
	) name4923 (
		_w4735_,
		_w4856_,
		_w4858_,
		_w4989_
	);
	LUT4 #(
		.INIT('h8f00)
	) name4924 (
		_w4601_,
		_w4603_,
		_w4865_,
		_w4989_,
		_w4990_
	);
	LUT3 #(
		.INIT('h32)
	) name4925 (
		_w4986_,
		_w4988_,
		_w4990_,
		_w4991_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name4926 (
		_w4854_,
		_w4857_,
		_w4866_,
		_w4984_,
		_w4992_
	);
	LUT3 #(
		.INIT('hd0)
	) name4927 (
		_w4735_,
		_w4856_,
		_w4992_,
		_w4993_
	);
	LUT4 #(
		.INIT('h8f00)
	) name4928 (
		_w4601_,
		_w4603_,
		_w4865_,
		_w4993_,
		_w4994_
	);
	LUT3 #(
		.INIT('h51)
	) name4929 (
		_w4911_,
		_w4979_,
		_w4980_,
		_w4995_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4930 (
		_w4802_,
		_w4867_,
		_w4888_,
		_w4889_,
		_w4996_
	);
	LUT3 #(
		.INIT('h32)
	) name4931 (
		_w4953_,
		_w4954_,
		_w4973_,
		_w4997_
	);
	LUT3 #(
		.INIT('h31)
	) name4932 (
		_w4876_,
		_w4885_,
		_w4886_,
		_w4998_
	);
	LUT3 #(
		.INIT('h32)
	) name4933 (
		_w4932_,
		_w4933_,
		_w4934_,
		_w4999_
	);
	LUT3 #(
		.INIT('h0d)
	) name4934 (
		_w4779_,
		_w4949_,
		_w4950_,
		_w5000_
	);
	LUT3 #(
		.INIT('h0d)
	) name4935 (
		_w4960_,
		_w4961_,
		_w4962_,
		_w5001_
	);
	LUT3 #(
		.INIT('h69)
	) name4936 (
		_w4999_,
		_w5000_,
		_w5001_,
		_w5002_
	);
	LUT3 #(
		.INIT('h71)
	) name4937 (
		_w4881_,
		_w4882_,
		_w4883_,
		_w5003_
	);
	LUT3 #(
		.INIT('h8e)
	) name4938 (
		_w4869_,
		_w4870_,
		_w4871_,
		_w5004_
	);
	LUT3 #(
		.INIT('h69)
	) name4939 (
		_w5002_,
		_w5003_,
		_w5004_,
		_w5005_
	);
	LUT4 #(
		.INIT('hb200)
	) name4940 (
		_w4876_,
		_w4880_,
		_w4884_,
		_w5005_,
		_w5006_
	);
	LUT4 #(
		.INIT('h004d)
	) name4941 (
		_w4876_,
		_w4880_,
		_w4884_,
		_w5005_,
		_w5007_
	);
	LUT4 #(
		.INIT('h31ce)
	) name4942 (
		_w4876_,
		_w4885_,
		_w4886_,
		_w5005_,
		_w5008_
	);
	LUT2 #(
		.INIT('h6)
	) name4943 (
		_w4997_,
		_w5008_,
		_w5009_
	);
	LUT3 #(
		.INIT('h32)
	) name4944 (
		_w4929_,
		_w4930_,
		_w4936_,
		_w5010_
	);
	LUT3 #(
		.INIT('h32)
	) name4945 (
		_w4946_,
		_w4947_,
		_w4952_,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name4946 (
		_w5010_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h8)
	) name4947 (
		_w5010_,
		_w5011_,
		_w5013_
	);
	LUT2 #(
		.INIT('h6)
	) name4948 (
		_w5010_,
		_w5011_,
		_w5014_
	);
	LUT3 #(
		.INIT('h54)
	) name4949 (
		_w4901_,
		_w4902_,
		_w4904_,
		_w5015_
	);
	LUT3 #(
		.INIT('h0d)
	) name4950 (
		_w4967_,
		_w4968_,
		_w4970_,
		_w5016_
	);
	LUT3 #(
		.INIT('h0d)
	) name4951 (
		_w4775_,
		_w4956_,
		_w4958_,
		_w5017_
	);
	LUT3 #(
		.INIT('h0d)
	) name4952 (
		_w4941_,
		_w4942_,
		_w4944_,
		_w5018_
	);
	LUT3 #(
		.INIT('h96)
	) name4953 (
		_w5016_,
		_w5017_,
		_w5018_,
		_w5019_
	);
	LUT3 #(
		.INIT('h0d)
	) name4954 (
		_w4925_,
		_w4926_,
		_w4927_,
		_w5020_
	);
	LUT3 #(
		.INIT('h0d)
	) name4955 (
		_w4759_,
		_w4921_,
		_w4923_,
		_w5021_
	);
	LUT3 #(
		.INIT('h0d)
	) name4956 (
		_w4937_,
		_w4938_,
		_w4939_,
		_w5022_
	);
	LUT3 #(
		.INIT('h96)
	) name4957 (
		_w5020_,
		_w5021_,
		_w5022_,
		_w5023_
	);
	LUT3 #(
		.INIT('h32)
	) name4958 (
		_w4964_,
		_w4965_,
		_w4972_,
		_w5024_
	);
	LUT3 #(
		.INIT('h96)
	) name4959 (
		_w5019_,
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT3 #(
		.INIT('h60)
	) name4960 (
		_w5014_,
		_w5015_,
		_w5025_,
		_w5026_
	);
	LUT3 #(
		.INIT('h96)
	) name4961 (
		_w5014_,
		_w5015_,
		_w5025_,
		_w5027_
	);
	LUT4 #(
		.INIT('h8e00)
	) name4962 (
		_w4915_,
		_w4916_,
		_w4920_,
		_w5027_,
		_w5028_
	);
	LUT4 #(
		.INIT('hba45)
	) name4963 (
		_w4917_,
		_w4918_,
		_w4920_,
		_w5027_,
		_w5029_
	);
	LUT3 #(
		.INIT('h96)
	) name4964 (
		_w4996_,
		_w5009_,
		_w5029_,
		_w5030_
	);
	LUT4 #(
		.INIT('h004d)
	) name4965 (
		_w4912_,
		_w4913_,
		_w4978_,
		_w5030_,
		_w5031_
	);
	LUT4 #(
		.INIT('hb200)
	) name4966 (
		_w4912_,
		_w4913_,
		_w4978_,
		_w5030_,
		_w5032_
	);
	LUT3 #(
		.INIT('h0e)
	) name4967 (
		_w4891_,
		_w4907_,
		_w4908_,
		_w5033_
	);
	LUT3 #(
		.INIT('h0e)
	) name4968 (
		_w4914_,
		_w4975_,
		_w4976_,
		_w5034_
	);
	LUT3 #(
		.INIT('he8)
	) name4969 (
		_w4892_,
		_w4896_,
		_w4905_,
		_w5035_
	);
	LUT3 #(
		.INIT('hb2)
	) name4970 (
		_w4893_,
		_w4894_,
		_w4895_,
		_w5036_
	);
	LUT4 #(
		.INIT('h153f)
	) name4971 (
		\a[9] ,
		\a[10] ,
		\a[59] ,
		\a[60] ,
		_w5037_
	);
	LUT4 #(
		.INIT('h8000)
	) name4972 (
		\a[9] ,
		\a[10] ,
		\a[59] ,
		\a[60] ,
		_w5038_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4973 (
		\a[9] ,
		\a[10] ,
		\a[59] ,
		\a[60] ,
		_w5039_
	);
	LUT4 #(
		.INIT('h153f)
	) name4974 (
		\a[24] ,
		\a[25] ,
		\a[44] ,
		\a[45] ,
		_w5040_
	);
	LUT2 #(
		.INIT('h8)
	) name4975 (
		\a[25] ,
		\a[45] ,
		_w5041_
	);
	LUT4 #(
		.INIT('h8000)
	) name4976 (
		\a[24] ,
		\a[25] ,
		\a[44] ,
		\a[45] ,
		_w5042_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4977 (
		\a[24] ,
		\a[25] ,
		\a[44] ,
		\a[45] ,
		_w5043_
	);
	LUT4 #(
		.INIT('h1248)
	) name4978 (
		_w4897_,
		_w4943_,
		_w5039_,
		_w5043_,
		_w5044_
	);
	LUT4 #(
		.INIT('h8421)
	) name4979 (
		_w4897_,
		_w4943_,
		_w5039_,
		_w5043_,
		_w5045_
	);
	LUT4 #(
		.INIT('h6996)
	) name4980 (
		_w4897_,
		_w4943_,
		_w5039_,
		_w5043_,
		_w5046_
	);
	LUT4 #(
		.INIT('h153f)
	) name4981 (
		\a[26] ,
		\a[27] ,
		\a[42] ,
		\a[43] ,
		_w5047_
	);
	LUT4 #(
		.INIT('h8000)
	) name4982 (
		\a[26] ,
		\a[27] ,
		\a[42] ,
		\a[43] ,
		_w5048_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4983 (
		\a[26] ,
		\a[27] ,
		\a[42] ,
		\a[43] ,
		_w5049_
	);
	LUT2 #(
		.INIT('h6)
	) name4984 (
		_w4969_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h6)
	) name4985 (
		_w5046_,
		_w5050_,
		_w5051_
	);
	LUT4 #(
		.INIT('h153f)
	) name4986 (
		\a[7] ,
		\a[8] ,
		\a[60] ,
		\a[61] ,
		_w5052_
	);
	LUT4 #(
		.INIT('h000d)
	) name4987 (
		_w4762_,
		_w4763_,
		_w4764_,
		_w4898_,
		_w5053_
	);
	LUT4 #(
		.INIT('h153f)
	) name4988 (
		\a[12] ,
		\a[13] ,
		\a[56] ,
		\a[57] ,
		_w5054_
	);
	LUT4 #(
		.INIT('h8000)
	) name4989 (
		\a[12] ,
		\a[13] ,
		\a[56] ,
		\a[57] ,
		_w5055_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4990 (
		\a[12] ,
		\a[13] ,
		\a[56] ,
		\a[57] ,
		_w5056_
	);
	LUT2 #(
		.INIT('h6)
	) name4991 (
		_w4957_,
		_w5056_,
		_w5057_
	);
	LUT2 #(
		.INIT('h8)
	) name4992 (
		\a[14] ,
		\a[55] ,
		_w5058_
	);
	LUT4 #(
		.INIT('h153f)
	) name4993 (
		\a[21] ,
		\a[22] ,
		\a[47] ,
		\a[48] ,
		_w5059_
	);
	LUT2 #(
		.INIT('h8)
	) name4994 (
		\a[22] ,
		\a[48] ,
		_w5060_
	);
	LUT4 #(
		.INIT('h8000)
	) name4995 (
		\a[21] ,
		\a[22] ,
		\a[47] ,
		\a[48] ,
		_w5061_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name4996 (
		\a[21] ,
		\a[22] ,
		\a[47] ,
		\a[48] ,
		_w5062_
	);
	LUT2 #(
		.INIT('h6)
	) name4997 (
		_w5058_,
		_w5062_,
		_w5063_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name4998 (
		_w5052_,
		_w5053_,
		_w5057_,
		_w5063_,
		_w5064_
	);
	LUT3 #(
		.INIT('h96)
	) name4999 (
		_w5036_,
		_w5051_,
		_w5064_,
		_w5065_
	);
	LUT3 #(
		.INIT('hd4)
	) name5000 (
		_w4872_,
		_w4873_,
		_w4874_,
		_w5066_
	);
	LUT4 #(
		.INIT('h153f)
	) name5001 (
		\a[17] ,
		\a[18] ,
		\a[51] ,
		\a[52] ,
		_w5067_
	);
	LUT4 #(
		.INIT('h8000)
	) name5002 (
		\a[17] ,
		\a[18] ,
		\a[51] ,
		\a[52] ,
		_w5068_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5003 (
		\a[17] ,
		\a[18] ,
		\a[51] ,
		\a[52] ,
		_w5069_
	);
	LUT2 #(
		.INIT('h8)
	) name5004 (
		\a[28] ,
		\a[41] ,
		_w5070_
	);
	LUT4 #(
		.INIT('h153f)
	) name5005 (
		\a[29] ,
		\a[30] ,
		\a[39] ,
		\a[40] ,
		_w5071_
	);
	LUT4 #(
		.INIT('h8000)
	) name5006 (
		\a[29] ,
		\a[30] ,
		\a[39] ,
		\a[40] ,
		_w5072_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5007 (
		\a[29] ,
		\a[30] ,
		\a[39] ,
		\a[40] ,
		_w5073_
	);
	LUT4 #(
		.INIT('h0660)
	) name5008 (
		_w4922_,
		_w5069_,
		_w5070_,
		_w5073_,
		_w5074_
	);
	LUT4 #(
		.INIT('h6996)
	) name5009 (
		_w4922_,
		_w5069_,
		_w5070_,
		_w5073_,
		_w5075_
	);
	LUT4 #(
		.INIT('h1700)
	) name5010 (
		_w4877_,
		_w4878_,
		_w4879_,
		_w5075_,
		_w5076_
	);
	LUT4 #(
		.INIT('he817)
	) name5011 (
		_w4877_,
		_w4878_,
		_w4879_,
		_w5075_,
		_w5077_
	);
	LUT2 #(
		.INIT('h8)
	) name5012 (
		\a[31] ,
		\a[38] ,
		_w5078_
	);
	LUT4 #(
		.INIT('h153f)
	) name5013 (
		\a[32] ,
		\a[33] ,
		\a[36] ,
		\a[37] ,
		_w5079_
	);
	LUT4 #(
		.INIT('h8000)
	) name5014 (
		\a[32] ,
		\a[33] ,
		\a[36] ,
		\a[37] ,
		_w5080_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5015 (
		\a[32] ,
		\a[33] ,
		\a[36] ,
		\a[37] ,
		_w5081_
	);
	LUT4 #(
		.INIT('h9a30)
	) name5016 (
		\a[7] ,
		\a[34] ,
		\a[35] ,
		\a[62] ,
		_w5082_
	);
	LUT3 #(
		.INIT('h60)
	) name5017 (
		_w5078_,
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT3 #(
		.INIT('h09)
	) name5018 (
		_w5078_,
		_w5081_,
		_w5082_,
		_w5084_
	);
	LUT3 #(
		.INIT('h96)
	) name5019 (
		_w5078_,
		_w5081_,
		_w5082_,
		_w5085_
	);
	LUT2 #(
		.INIT('h8)
	) name5020 (
		\a[15] ,
		\a[54] ,
		_w5086_
	);
	LUT4 #(
		.INIT('h153f)
	) name5021 (
		\a[16] ,
		\a[20] ,
		\a[49] ,
		\a[53] ,
		_w5087_
	);
	LUT4 #(
		.INIT('h8000)
	) name5022 (
		\a[16] ,
		\a[20] ,
		\a[49] ,
		\a[53] ,
		_w5088_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5023 (
		\a[16] ,
		\a[20] ,
		\a[49] ,
		\a[53] ,
		_w5089_
	);
	LUT2 #(
		.INIT('h6)
	) name5024 (
		_w5086_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h6)
	) name5025 (
		_w5085_,
		_w5090_,
		_w5091_
	);
	LUT2 #(
		.INIT('h8)
	) name5026 (
		_w5077_,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h1)
	) name5027 (
		_w5077_,
		_w5091_,
		_w5093_
	);
	LUT2 #(
		.INIT('h6)
	) name5028 (
		_w5077_,
		_w5091_,
		_w5094_
	);
	LUT2 #(
		.INIT('h6)
	) name5029 (
		_w5066_,
		_w5094_,
		_w5095_
	);
	LUT3 #(
		.INIT('h96)
	) name5030 (
		_w5035_,
		_w5065_,
		_w5095_,
		_w5096_
	);
	LUT3 #(
		.INIT('h96)
	) name5031 (
		_w5033_,
		_w5034_,
		_w5096_,
		_w5097_
	);
	LUT3 #(
		.INIT('he1)
	) name5032 (
		_w5031_,
		_w5032_,
		_w5097_,
		_w5098_
	);
	LUT2 #(
		.INIT('h4)
	) name5033 (
		_w4995_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h2)
	) name5034 (
		_w4995_,
		_w5098_,
		_w5100_
	);
	LUT2 #(
		.INIT('h9)
	) name5035 (
		_w4995_,
		_w5098_,
		_w5101_
	);
	LUT3 #(
		.INIT('h1e)
	) name5036 (
		_w4985_,
		_w4994_,
		_w5101_,
		_w5102_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5037 (
		_w4866_,
		_w4981_,
		_w4983_,
		_w5099_,
		_w5103_
	);
	LUT3 #(
		.INIT('h54)
	) name5038 (
		_w5031_,
		_w5032_,
		_w5097_,
		_w5104_
	);
	LUT3 #(
		.INIT('he8)
	) name5039 (
		_w4996_,
		_w5009_,
		_w5029_,
		_w5105_
	);
	LUT3 #(
		.INIT('h31)
	) name5040 (
		_w5066_,
		_w5092_,
		_w5093_,
		_w5106_
	);
	LUT3 #(
		.INIT('h0d)
	) name5041 (
		_w4969_,
		_w5047_,
		_w5048_,
		_w5107_
	);
	LUT3 #(
		.INIT('h0d)
	) name5042 (
		_w5070_,
		_w5071_,
		_w5072_,
		_w5108_
	);
	LUT3 #(
		.INIT('h0d)
	) name5043 (
		_w4943_,
		_w5040_,
		_w5042_,
		_w5109_
	);
	LUT3 #(
		.INIT('h96)
	) name5044 (
		_w5107_,
		_w5108_,
		_w5109_,
		_w5110_
	);
	LUT3 #(
		.INIT('h13)
	) name5045 (
		\a[7] ,
		\a[34] ,
		\a[62] ,
		_w5111_
	);
	LUT2 #(
		.INIT('h8)
	) name5046 (
		\a[8] ,
		\a[62] ,
		_w5112_
	);
	LUT3 #(
		.INIT('h80)
	) name5047 (
		\a[8] ,
		\a[35] ,
		\a[62] ,
		_w5113_
	);
	LUT2 #(
		.INIT('h4)
	) name5048 (
		_w5111_,
		_w5113_,
		_w5114_
	);
	LUT4 #(
		.INIT('he0c0)
	) name5049 (
		\a[7] ,
		\a[34] ,
		\a[35] ,
		\a[62] ,
		_w5115_
	);
	LUT2 #(
		.INIT('h1)
	) name5050 (
		_w5112_,
		_w5115_,
		_w5116_
	);
	LUT3 #(
		.INIT('hd2)
	) name5051 (
		\a[35] ,
		_w5111_,
		_w5112_,
		_w5117_
	);
	LUT3 #(
		.INIT('h0d)
	) name5052 (
		_w5078_,
		_w5079_,
		_w5080_,
		_w5118_
	);
	LUT2 #(
		.INIT('h6)
	) name5053 (
		_w5117_,
		_w5118_,
		_w5119_
	);
	LUT4 #(
		.INIT('he11e)
	) name5054 (
		_w5074_,
		_w5076_,
		_w5110_,
		_w5119_,
		_w5120_
	);
	LUT4 #(
		.INIT('hf110)
	) name5055 (
		_w5052_,
		_w5053_,
		_w5057_,
		_w5063_,
		_w5121_
	);
	LUT3 #(
		.INIT('h32)
	) name5056 (
		_w5044_,
		_w5045_,
		_w5050_,
		_w5122_
	);
	LUT3 #(
		.INIT('h32)
	) name5057 (
		_w5083_,
		_w5084_,
		_w5090_,
		_w5123_
	);
	LUT3 #(
		.INIT('h96)
	) name5058 (
		_w5121_,
		_w5122_,
		_w5123_,
		_w5124_
	);
	LUT3 #(
		.INIT('h69)
	) name5059 (
		_w5106_,
		_w5120_,
		_w5124_,
		_w5125_
	);
	LUT3 #(
		.INIT('h0e)
	) name5060 (
		_w4997_,
		_w5006_,
		_w5007_,
		_w5126_
	);
	LUT3 #(
		.INIT('h71)
	) name5061 (
		_w5019_,
		_w5023_,
		_w5024_,
		_w5127_
	);
	LUT2 #(
		.INIT('h8)
	) name5062 (
		\a[28] ,
		\a[42] ,
		_w5128_
	);
	LUT4 #(
		.INIT('h153f)
	) name5063 (
		\a[7] ,
		\a[23] ,
		\a[47] ,
		\a[63] ,
		_w5129_
	);
	LUT4 #(
		.INIT('h8000)
	) name5064 (
		\a[7] ,
		\a[23] ,
		\a[47] ,
		\a[63] ,
		_w5130_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5065 (
		\a[7] ,
		\a[23] ,
		\a[47] ,
		\a[63] ,
		_w5131_
	);
	LUT2 #(
		.INIT('h8)
	) name5066 (
		\a[29] ,
		\a[41] ,
		_w5132_
	);
	LUT4 #(
		.INIT('h153f)
	) name5067 (
		\a[30] ,
		\a[31] ,
		\a[39] ,
		\a[40] ,
		_w5133_
	);
	LUT4 #(
		.INIT('h8000)
	) name5068 (
		\a[30] ,
		\a[31] ,
		\a[39] ,
		\a[40] ,
		_w5134_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5069 (
		\a[30] ,
		\a[31] ,
		\a[39] ,
		\a[40] ,
		_w5135_
	);
	LUT4 #(
		.INIT('h0660)
	) name5070 (
		_w5128_,
		_w5131_,
		_w5132_,
		_w5135_,
		_w5136_
	);
	LUT4 #(
		.INIT('h6996)
	) name5071 (
		_w5128_,
		_w5131_,
		_w5132_,
		_w5135_,
		_w5137_
	);
	LUT4 #(
		.INIT('h1700)
	) name5072 (
		_w5020_,
		_w5021_,
		_w5022_,
		_w5137_,
		_w5138_
	);
	LUT4 #(
		.INIT('he817)
	) name5073 (
		_w5020_,
		_w5021_,
		_w5022_,
		_w5137_,
		_w5139_
	);
	LUT4 #(
		.INIT('h153f)
	) name5074 (
		\a[14] ,
		\a[15] ,
		\a[55] ,
		\a[56] ,
		_w5140_
	);
	LUT4 #(
		.INIT('h8000)
	) name5075 (
		\a[14] ,
		\a[15] ,
		\a[55] ,
		\a[56] ,
		_w5141_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5076 (
		\a[14] ,
		\a[15] ,
		\a[55] ,
		\a[56] ,
		_w5142_
	);
	LUT4 #(
		.INIT('h153f)
	) name5077 (
		\a[26] ,
		\a[27] ,
		\a[43] ,
		\a[44] ,
		_w5143_
	);
	LUT2 #(
		.INIT('h8)
	) name5078 (
		\a[27] ,
		\a[44] ,
		_w5144_
	);
	LUT4 #(
		.INIT('h8000)
	) name5079 (
		\a[26] ,
		\a[27] ,
		\a[43] ,
		\a[44] ,
		_w5145_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5080 (
		\a[26] ,
		\a[27] ,
		\a[43] ,
		\a[44] ,
		_w5146_
	);
	LUT4 #(
		.INIT('h1428)
	) name5081 (
		_w5041_,
		_w5060_,
		_w5142_,
		_w5146_,
		_w5147_
	);
	LUT4 #(
		.INIT('h8241)
	) name5082 (
		_w5041_,
		_w5060_,
		_w5142_,
		_w5146_,
		_w5148_
	);
	LUT4 #(
		.INIT('h6996)
	) name5083 (
		_w5041_,
		_w5060_,
		_w5142_,
		_w5146_,
		_w5149_
	);
	LUT2 #(
		.INIT('h8)
	) name5084 (
		\a[21] ,
		\a[49] ,
		_w5150_
	);
	LUT4 #(
		.INIT('h153f)
	) name5085 (
		\a[19] ,
		\a[20] ,
		\a[50] ,
		\a[51] ,
		_w5151_
	);
	LUT4 #(
		.INIT('h8000)
	) name5086 (
		\a[19] ,
		\a[20] ,
		\a[50] ,
		\a[51] ,
		_w5152_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5087 (
		\a[19] ,
		\a[20] ,
		\a[50] ,
		\a[51] ,
		_w5153_
	);
	LUT2 #(
		.INIT('h6)
	) name5088 (
		_w5150_,
		_w5153_,
		_w5154_
	);
	LUT2 #(
		.INIT('h6)
	) name5089 (
		_w5149_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h8)
	) name5090 (
		_w5139_,
		_w5155_,
		_w5156_
	);
	LUT2 #(
		.INIT('h1)
	) name5091 (
		_w5139_,
		_w5155_,
		_w5157_
	);
	LUT2 #(
		.INIT('h6)
	) name5092 (
		_w5139_,
		_w5155_,
		_w5158_
	);
	LUT2 #(
		.INIT('h8)
	) name5093 (
		_w5127_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h1)
	) name5094 (
		_w5127_,
		_w5158_,
		_w5160_
	);
	LUT2 #(
		.INIT('h6)
	) name5095 (
		_w5127_,
		_w5158_,
		_w5161_
	);
	LUT3 #(
		.INIT('hd4)
	) name5096 (
		_w5002_,
		_w5003_,
		_w5004_,
		_w5162_
	);
	LUT3 #(
		.INIT('h32)
	) name5097 (
		_w5086_,
		_w5087_,
		_w5088_,
		_w5163_
	);
	LUT3 #(
		.INIT('h0d)
	) name5098 (
		_w4922_,
		_w5067_,
		_w5068_,
		_w5164_
	);
	LUT2 #(
		.INIT('h8)
	) name5099 (
		\a[32] ,
		\a[38] ,
		_w5165_
	);
	LUT4 #(
		.INIT('h153f)
	) name5100 (
		\a[33] ,
		\a[34] ,
		\a[36] ,
		\a[37] ,
		_w5166_
	);
	LUT4 #(
		.INIT('h8000)
	) name5101 (
		\a[33] ,
		\a[34] ,
		\a[36] ,
		\a[37] ,
		_w5167_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5102 (
		\a[33] ,
		\a[34] ,
		\a[36] ,
		\a[37] ,
		_w5168_
	);
	LUT2 #(
		.INIT('h6)
	) name5103 (
		_w5165_,
		_w5168_,
		_w5169_
	);
	LUT3 #(
		.INIT('h96)
	) name5104 (
		_w5163_,
		_w5164_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h8)
	) name5105 (
		\a[9] ,
		\a[61] ,
		_w5171_
	);
	LUT4 #(
		.INIT('h153f)
	) name5106 (
		\a[10] ,
		\a[11] ,
		\a[59] ,
		\a[60] ,
		_w5172_
	);
	LUT2 #(
		.INIT('h8)
	) name5107 (
		\a[11] ,
		\a[60] ,
		_w5173_
	);
	LUT4 #(
		.INIT('h8000)
	) name5108 (
		\a[10] ,
		\a[11] ,
		\a[59] ,
		\a[60] ,
		_w5174_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5109 (
		\a[10] ,
		\a[11] ,
		\a[59] ,
		\a[60] ,
		_w5175_
	);
	LUT4 #(
		.INIT('h153f)
	) name5110 (
		\a[16] ,
		\a[17] ,
		\a[53] ,
		\a[54] ,
		_w5176_
	);
	LUT4 #(
		.INIT('h8000)
	) name5111 (
		\a[16] ,
		\a[17] ,
		\a[53] ,
		\a[54] ,
		_w5177_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5112 (
		\a[16] ,
		\a[17] ,
		\a[53] ,
		\a[54] ,
		_w5178_
	);
	LUT4 #(
		.INIT('h1428)
	) name5113 (
		_w3784_,
		_w5171_,
		_w5175_,
		_w5178_,
		_w5179_
	);
	LUT4 #(
		.INIT('h8241)
	) name5114 (
		_w3784_,
		_w5171_,
		_w5175_,
		_w5178_,
		_w5180_
	);
	LUT4 #(
		.INIT('h6996)
	) name5115 (
		_w3784_,
		_w5171_,
		_w5175_,
		_w5178_,
		_w5181_
	);
	LUT2 #(
		.INIT('h8)
	) name5116 (
		\a[12] ,
		\a[58] ,
		_w5182_
	);
	LUT4 #(
		.INIT('h153f)
	) name5117 (
		\a[13] ,
		\a[24] ,
		\a[46] ,
		\a[57] ,
		_w5183_
	);
	LUT4 #(
		.INIT('h8000)
	) name5118 (
		\a[13] ,
		\a[24] ,
		\a[46] ,
		\a[57] ,
		_w5184_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5119 (
		\a[13] ,
		\a[24] ,
		\a[46] ,
		\a[57] ,
		_w5185_
	);
	LUT2 #(
		.INIT('h6)
	) name5120 (
		_w5182_,
		_w5185_,
		_w5186_
	);
	LUT2 #(
		.INIT('h6)
	) name5121 (
		_w5181_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h4)
	) name5122 (
		_w5170_,
		_w5187_,
		_w5188_
	);
	LUT2 #(
		.INIT('h8)
	) name5123 (
		_w5170_,
		_w5187_,
		_w5189_
	);
	LUT4 #(
		.INIT('h00d4)
	) name5124 (
		_w5002_,
		_w5003_,
		_w5004_,
		_w5170_,
		_w5190_
	);
	LUT4 #(
		.INIT('h606b)
	) name5125 (
		_w5162_,
		_w5170_,
		_w5187_,
		_w5190_,
		_w5191_
	);
	LUT4 #(
		.INIT('h00b2)
	) name5126 (
		_w4997_,
		_w4998_,
		_w5005_,
		_w5191_,
		_w5192_
	);
	LUT4 #(
		.INIT('hed61)
	) name5127 (
		_w5126_,
		_w5161_,
		_w5191_,
		_w5192_,
		_w5193_
	);
	LUT3 #(
		.INIT('h96)
	) name5128 (
		_w5105_,
		_w5125_,
		_w5193_,
		_w5194_
	);
	LUT3 #(
		.INIT('h17)
	) name5129 (
		_w5035_,
		_w5065_,
		_w5095_,
		_w5195_
	);
	LUT3 #(
		.INIT('h17)
	) name5130 (
		_w5036_,
		_w5051_,
		_w5064_,
		_w5196_
	);
	LUT3 #(
		.INIT('h54)
	) name5131 (
		_w5012_,
		_w5013_,
		_w5015_,
		_w5197_
	);
	LUT3 #(
		.INIT('h0d)
	) name5132 (
		_w4957_,
		_w5054_,
		_w5055_,
		_w5198_
	);
	LUT3 #(
		.INIT('h0d)
	) name5133 (
		_w4897_,
		_w5037_,
		_w5038_,
		_w5199_
	);
	LUT3 #(
		.INIT('h0d)
	) name5134 (
		_w5058_,
		_w5059_,
		_w5061_,
		_w5200_
	);
	LUT3 #(
		.INIT('h96)
	) name5135 (
		_w5198_,
		_w5199_,
		_w5200_,
		_w5201_
	);
	LUT3 #(
		.INIT('h17)
	) name5136 (
		_w5016_,
		_w5017_,
		_w5018_,
		_w5202_
	);
	LUT3 #(
		.INIT('h2b)
	) name5137 (
		_w4999_,
		_w5000_,
		_w5001_,
		_w5203_
	);
	LUT3 #(
		.INIT('h69)
	) name5138 (
		_w5201_,
		_w5202_,
		_w5203_,
		_w5204_
	);
	LUT4 #(
		.INIT('he800)
	) name5139 (
		_w5010_,
		_w5011_,
		_w5015_,
		_w5204_,
		_w5205_
	);
	LUT4 #(
		.INIT('h0017)
	) name5140 (
		_w5010_,
		_w5011_,
		_w5015_,
		_w5204_,
		_w5206_
	);
	LUT4 #(
		.INIT('hab54)
	) name5141 (
		_w5012_,
		_w5013_,
		_w5015_,
		_w5204_,
		_w5207_
	);
	LUT2 #(
		.INIT('h9)
	) name5142 (
		_w5196_,
		_w5207_,
		_w5208_
	);
	LUT3 #(
		.INIT('h01)
	) name5143 (
		_w5026_,
		_w5028_,
		_w5208_,
		_w5209_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5144 (
		_w5026_,
		_w5028_,
		_w5195_,
		_w5208_,
		_w5210_
	);
	LUT4 #(
		.INIT('he800)
	) name5145 (
		_w5033_,
		_w5034_,
		_w5096_,
		_w5210_,
		_w5211_
	);
	LUT4 #(
		.INIT('h0017)
	) name5146 (
		_w5033_,
		_w5034_,
		_w5096_,
		_w5210_,
		_w5212_
	);
	LUT4 #(
		.INIT('h17e8)
	) name5147 (
		_w5033_,
		_w5034_,
		_w5096_,
		_w5210_,
		_w5213_
	);
	LUT2 #(
		.INIT('h2)
	) name5148 (
		_w5194_,
		_w5213_,
		_w5214_
	);
	LUT3 #(
		.INIT('h01)
	) name5149 (
		_w5194_,
		_w5211_,
		_w5212_,
		_w5215_
	);
	LUT3 #(
		.INIT('h56)
	) name5150 (
		_w5194_,
		_w5211_,
		_w5212_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name5151 (
		_w5104_,
		_w5216_,
		_w5217_
	);
	LUT3 #(
		.INIT('h02)
	) name5152 (
		_w5104_,
		_w5214_,
		_w5215_,
		_w5218_
	);
	LUT3 #(
		.INIT('ha9)
	) name5153 (
		_w5104_,
		_w5214_,
		_w5215_,
		_w5219_
	);
	LUT4 #(
		.INIT('hdc23)
	) name5154 (
		_w4994_,
		_w5100_,
		_w5103_,
		_w5219_,
		_w5220_
	);
	LUT3 #(
		.INIT('h32)
	) name5155 (
		_w5194_,
		_w5211_,
		_w5212_,
		_w5221_
	);
	LUT4 #(
		.INIT('he800)
	) name5156 (
		_w4996_,
		_w5009_,
		_w5029_,
		_w5125_,
		_w5222_
	);
	LUT4 #(
		.INIT('h17e8)
	) name5157 (
		_w4996_,
		_w5009_,
		_w5029_,
		_w5125_,
		_w5223_
	);
	LUT2 #(
		.INIT('h4)
	) name5158 (
		_w5193_,
		_w5223_,
		_w5224_
	);
	LUT4 #(
		.INIT('hb200)
	) name5159 (
		_w4997_,
		_w4998_,
		_w5005_,
		_w5191_,
		_w5225_
	);
	LUT2 #(
		.INIT('h4)
	) name5160 (
		_w5160_,
		_w5191_,
		_w5226_
	);
	LUT4 #(
		.INIT('h00b2)
	) name5161 (
		_w4997_,
		_w4998_,
		_w5005_,
		_w5160_,
		_w5227_
	);
	LUT4 #(
		.INIT('h2223)
	) name5162 (
		_w5159_,
		_w5225_,
		_w5226_,
		_w5227_,
		_w5228_
	);
	LUT3 #(
		.INIT('h54)
	) name5163 (
		_w5114_,
		_w5116_,
		_w5118_,
		_w5229_
	);
	LUT3 #(
		.INIT('h4d)
	) name5164 (
		_w5163_,
		_w5164_,
		_w5169_,
		_w5230_
	);
	LUT3 #(
		.INIT('h17)
	) name5165 (
		_w5107_,
		_w5108_,
		_w5109_,
		_w5231_
	);
	LUT3 #(
		.INIT('h96)
	) name5166 (
		_w5229_,
		_w5230_,
		_w5231_,
		_w5232_
	);
	LUT4 #(
		.INIT('h0eef)
	) name5167 (
		_w5074_,
		_w5076_,
		_w5110_,
		_w5119_,
		_w5233_
	);
	LUT2 #(
		.INIT('h1)
	) name5168 (
		_w5232_,
		_w5233_,
		_w5234_
	);
	LUT2 #(
		.INIT('h8)
	) name5169 (
		_w5232_,
		_w5233_,
		_w5235_
	);
	LUT2 #(
		.INIT('h6)
	) name5170 (
		_w5232_,
		_w5233_,
		_w5236_
	);
	LUT4 #(
		.INIT('h001b)
	) name5171 (
		_w5162_,
		_w5188_,
		_w5189_,
		_w5190_,
		_w5237_
	);
	LUT2 #(
		.INIT('h9)
	) name5172 (
		_w5236_,
		_w5237_,
		_w5238_
	);
	LUT3 #(
		.INIT('h2b)
	) name5173 (
		_w5106_,
		_w5120_,
		_w5124_,
		_w5239_
	);
	LUT2 #(
		.INIT('h2)
	) name5174 (
		_w5238_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h9)
	) name5175 (
		_w5238_,
		_w5239_,
		_w5241_
	);
	LUT2 #(
		.INIT('h9)
	) name5176 (
		_w5228_,
		_w5241_,
		_w5242_
	);
	LUT4 #(
		.INIT('h0017)
	) name5177 (
		_w4996_,
		_w5009_,
		_w5029_,
		_w5125_,
		_w5243_
	);
	LUT3 #(
		.INIT('h0d)
	) name5178 (
		_w5193_,
		_w5222_,
		_w5243_,
		_w5244_
	);
	LUT4 #(
		.INIT('h0efe)
	) name5179 (
		_w5222_,
		_w5224_,
		_w5242_,
		_w5244_,
		_w5245_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5180 (
		_w5026_,
		_w5028_,
		_w5195_,
		_w5208_,
		_w5246_
	);
	LUT4 #(
		.INIT('hef0e)
	) name5181 (
		_w5026_,
		_w5028_,
		_w5195_,
		_w5208_,
		_w5247_
	);
	LUT3 #(
		.INIT('h31)
	) name5182 (
		_w5127_,
		_w5156_,
		_w5157_,
		_w5248_
	);
	LUT3 #(
		.INIT('h17)
	) name5183 (
		_w5198_,
		_w5199_,
		_w5200_,
		_w5249_
	);
	LUT3 #(
		.INIT('h32)
	) name5184 (
		_w5179_,
		_w5180_,
		_w5186_,
		_w5250_
	);
	LUT3 #(
		.INIT('h32)
	) name5185 (
		_w5147_,
		_w5148_,
		_w5154_,
		_w5251_
	);
	LUT3 #(
		.INIT('h96)
	) name5186 (
		_w5249_,
		_w5250_,
		_w5251_,
		_w5252_
	);
	LUT3 #(
		.INIT('h0d)
	) name5187 (
		_w5182_,
		_w5183_,
		_w5184_,
		_w5253_
	);
	LUT3 #(
		.INIT('h0d)
	) name5188 (
		_w5171_,
		_w5172_,
		_w5174_,
		_w5254_
	);
	LUT3 #(
		.INIT('h0d)
	) name5189 (
		_w5041_,
		_w5143_,
		_w5145_,
		_w5255_
	);
	LUT3 #(
		.INIT('h96)
	) name5190 (
		_w5253_,
		_w5254_,
		_w5255_,
		_w5256_
	);
	LUT3 #(
		.INIT('h32)
	) name5191 (
		_w5128_,
		_w5129_,
		_w5130_,
		_w5257_
	);
	LUT3 #(
		.INIT('h0d)
	) name5192 (
		_w5132_,
		_w5133_,
		_w5134_,
		_w5258_
	);
	LUT3 #(
		.INIT('h0d)
	) name5193 (
		_w5060_,
		_w5140_,
		_w5141_,
		_w5259_
	);
	LUT3 #(
		.INIT('h96)
	) name5194 (
		_w5257_,
		_w5258_,
		_w5259_,
		_w5260_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5195 (
		_w5136_,
		_w5138_,
		_w5256_,
		_w5260_,
		_w5261_
	);
	LUT3 #(
		.INIT('h69)
	) name5196 (
		_w5248_,
		_w5252_,
		_w5261_,
		_w5262_
	);
	LUT3 #(
		.INIT('h32)
	) name5197 (
		_w5196_,
		_w5205_,
		_w5206_,
		_w5263_
	);
	LUT3 #(
		.INIT('hd4)
	) name5198 (
		_w5201_,
		_w5202_,
		_w5203_,
		_w5264_
	);
	LUT3 #(
		.INIT('h0d)
	) name5199 (
		_w3784_,
		_w5176_,
		_w5177_,
		_w5265_
	);
	LUT3 #(
		.INIT('h0d)
	) name5200 (
		_w5165_,
		_w5166_,
		_w5167_,
		_w5266_
	);
	LUT4 #(
		.INIT('h153f)
	) name5201 (
		\a[8] ,
		\a[10] ,
		\a[61] ,
		\a[63] ,
		_w5267_
	);
	LUT4 #(
		.INIT('h8000)
	) name5202 (
		\a[8] ,
		\a[10] ,
		\a[61] ,
		\a[63] ,
		_w5268_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5203 (
		\a[8] ,
		\a[10] ,
		\a[61] ,
		\a[63] ,
		_w5269_
	);
	LUT2 #(
		.INIT('h6)
	) name5204 (
		_w5173_,
		_w5269_,
		_w5270_
	);
	LUT3 #(
		.INIT('h69)
	) name5205 (
		_w5265_,
		_w5266_,
		_w5270_,
		_w5271_
	);
	LUT2 #(
		.INIT('h8)
	) name5206 (
		\a[21] ,
		\a[50] ,
		_w5272_
	);
	LUT4 #(
		.INIT('h153f)
	) name5207 (
		\a[19] ,
		\a[20] ,
		\a[51] ,
		\a[52] ,
		_w5273_
	);
	LUT4 #(
		.INIT('h8000)
	) name5208 (
		\a[19] ,
		\a[20] ,
		\a[51] ,
		\a[52] ,
		_w5274_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5209 (
		\a[19] ,
		\a[20] ,
		\a[51] ,
		\a[52] ,
		_w5275_
	);
	LUT2 #(
		.INIT('h8)
	) name5210 (
		\a[22] ,
		\a[49] ,
		_w5276_
	);
	LUT3 #(
		.INIT('h13)
	) name5211 (
		\a[9] ,
		\a[36] ,
		\a[62] ,
		_w5277_
	);
	LUT3 #(
		.INIT('h80)
	) name5212 (
		\a[9] ,
		\a[36] ,
		\a[62] ,
		_w5278_
	);
	LUT3 #(
		.INIT('h6c)
	) name5213 (
		\a[9] ,
		\a[36] ,
		\a[62] ,
		_w5279_
	);
	LUT4 #(
		.INIT('h0660)
	) name5214 (
		_w5272_,
		_w5275_,
		_w5276_,
		_w5279_,
		_w5280_
	);
	LUT4 #(
		.INIT('h9009)
	) name5215 (
		_w5272_,
		_w5275_,
		_w5276_,
		_w5279_,
		_w5281_
	);
	LUT4 #(
		.INIT('h6996)
	) name5216 (
		_w5272_,
		_w5275_,
		_w5276_,
		_w5279_,
		_w5282_
	);
	LUT2 #(
		.INIT('h8)
	) name5217 (
		\a[33] ,
		\a[38] ,
		_w5283_
	);
	LUT4 #(
		.INIT('h153f)
	) name5218 (
		\a[34] ,
		\a[35] ,
		\a[36] ,
		\a[37] ,
		_w5284_
	);
	LUT4 #(
		.INIT('h8000)
	) name5219 (
		\a[34] ,
		\a[35] ,
		\a[36] ,
		\a[37] ,
		_w5285_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5220 (
		\a[34] ,
		\a[35] ,
		\a[36] ,
		\a[37] ,
		_w5286_
	);
	LUT2 #(
		.INIT('h6)
	) name5221 (
		_w5283_,
		_w5286_,
		_w5287_
	);
	LUT2 #(
		.INIT('h6)
	) name5222 (
		_w5282_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h4)
	) name5223 (
		_w5271_,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('h8)
	) name5224 (
		_w5271_,
		_w5288_,
		_w5290_
	);
	LUT4 #(
		.INIT('h00d4)
	) name5225 (
		_w5201_,
		_w5202_,
		_w5203_,
		_w5271_,
		_w5291_
	);
	LUT4 #(
		.INIT('h606b)
	) name5226 (
		_w5264_,
		_w5271_,
		_w5288_,
		_w5291_,
		_w5292_
	);
	LUT4 #(
		.INIT('hd400)
	) name5227 (
		_w5196_,
		_w5197_,
		_w5204_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h8)
	) name5228 (
		\a[13] ,
		\a[59] ,
		_w5294_
	);
	LUT4 #(
		.INIT('h8000)
	) name5229 (
		\a[12] ,
		\a[13] ,
		\a[58] ,
		\a[59] ,
		_w5295_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5230 (
		\a[12] ,
		\a[13] ,
		\a[58] ,
		\a[59] ,
		_w5296_
	);
	LUT4 #(
		.INIT('hf20d)
	) name5231 (
		_w5150_,
		_w5151_,
		_w5152_,
		_w5296_,
		_w5297_
	);
	LUT2 #(
		.INIT('h8)
	) name5232 (
		\a[14] ,
		\a[57] ,
		_w5298_
	);
	LUT4 #(
		.INIT('h153f)
	) name5233 (
		\a[15] ,
		\a[16] ,
		\a[55] ,
		\a[56] ,
		_w5299_
	);
	LUT4 #(
		.INIT('h8000)
	) name5234 (
		\a[15] ,
		\a[16] ,
		\a[55] ,
		\a[56] ,
		_w5300_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5235 (
		\a[15] ,
		\a[16] ,
		\a[55] ,
		\a[56] ,
		_w5301_
	);
	LUT2 #(
		.INIT('h8)
	) name5236 (
		\a[24] ,
		\a[47] ,
		_w5302_
	);
	LUT4 #(
		.INIT('h153f)
	) name5237 (
		\a[25] ,
		\a[26] ,
		\a[45] ,
		\a[46] ,
		_w5303_
	);
	LUT2 #(
		.INIT('h8)
	) name5238 (
		\a[26] ,
		\a[46] ,
		_w5304_
	);
	LUT4 #(
		.INIT('h8000)
	) name5239 (
		\a[25] ,
		\a[26] ,
		\a[45] ,
		\a[46] ,
		_w5305_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5240 (
		\a[25] ,
		\a[26] ,
		\a[45] ,
		\a[46] ,
		_w5306_
	);
	LUT4 #(
		.INIT('h0660)
	) name5241 (
		_w5298_,
		_w5301_,
		_w5302_,
		_w5306_,
		_w5307_
	);
	LUT4 #(
		.INIT('h9009)
	) name5242 (
		_w5298_,
		_w5301_,
		_w5302_,
		_w5306_,
		_w5308_
	);
	LUT4 #(
		.INIT('h6996)
	) name5243 (
		_w5298_,
		_w5301_,
		_w5302_,
		_w5306_,
		_w5309_
	);
	LUT4 #(
		.INIT('h153f)
	) name5244 (
		\a[28] ,
		\a[29] ,
		\a[42] ,
		\a[43] ,
		_w5310_
	);
	LUT2 #(
		.INIT('h8)
	) name5245 (
		\a[29] ,
		\a[43] ,
		_w5311_
	);
	LUT4 #(
		.INIT('h8000)
	) name5246 (
		\a[28] ,
		\a[29] ,
		\a[42] ,
		\a[43] ,
		_w5312_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5247 (
		\a[28] ,
		\a[29] ,
		\a[42] ,
		\a[43] ,
		_w5313_
	);
	LUT2 #(
		.INIT('h8)
	) name5248 (
		\a[30] ,
		\a[41] ,
		_w5314_
	);
	LUT4 #(
		.INIT('h153f)
	) name5249 (
		\a[31] ,
		\a[32] ,
		\a[39] ,
		\a[40] ,
		_w5315_
	);
	LUT2 #(
		.INIT('h8)
	) name5250 (
		\a[32] ,
		\a[40] ,
		_w5316_
	);
	LUT4 #(
		.INIT('h8000)
	) name5251 (
		\a[31] ,
		\a[32] ,
		\a[39] ,
		\a[40] ,
		_w5317_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5252 (
		\a[31] ,
		\a[32] ,
		\a[39] ,
		\a[40] ,
		_w5318_
	);
	LUT4 #(
		.INIT('h0660)
	) name5253 (
		_w5144_,
		_w5313_,
		_w5314_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('h9009)
	) name5254 (
		_w5144_,
		_w5313_,
		_w5314_,
		_w5318_,
		_w5320_
	);
	LUT4 #(
		.INIT('h6996)
	) name5255 (
		_w5144_,
		_w5313_,
		_w5314_,
		_w5318_,
		_w5321_
	);
	LUT2 #(
		.INIT('h8)
	) name5256 (
		\a[23] ,
		\a[48] ,
		_w5322_
	);
	LUT4 #(
		.INIT('h153f)
	) name5257 (
		\a[17] ,
		\a[18] ,
		\a[53] ,
		\a[54] ,
		_w5323_
	);
	LUT4 #(
		.INIT('h8000)
	) name5258 (
		\a[17] ,
		\a[18] ,
		\a[53] ,
		\a[54] ,
		_w5324_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5259 (
		\a[17] ,
		\a[18] ,
		\a[53] ,
		\a[54] ,
		_w5325_
	);
	LUT2 #(
		.INIT('h6)
	) name5260 (
		_w5322_,
		_w5325_,
		_w5326_
	);
	LUT4 #(
		.INIT('h0990)
	) name5261 (
		_w5297_,
		_w5309_,
		_w5321_,
		_w5326_,
		_w5327_
	);
	LUT4 #(
		.INIT('h9669)
	) name5262 (
		_w5297_,
		_w5309_,
		_w5321_,
		_w5326_,
		_w5328_
	);
	LUT4 #(
		.INIT('he800)
	) name5263 (
		_w5121_,
		_w5122_,
		_w5123_,
		_w5328_,
		_w5329_
	);
	LUT4 #(
		.INIT('h17e8)
	) name5264 (
		_w5121_,
		_w5122_,
		_w5123_,
		_w5328_,
		_w5330_
	);
	LUT4 #(
		.INIT('h0032)
	) name5265 (
		_w5196_,
		_w5205_,
		_w5206_,
		_w5292_,
		_w5331_
	);
	LUT4 #(
		.INIT('hf949)
	) name5266 (
		_w5263_,
		_w5292_,
		_w5330_,
		_w5331_,
		_w5332_
	);
	LUT3 #(
		.INIT('h69)
	) name5267 (
		_w5247_,
		_w5262_,
		_w5332_,
		_w5333_
	);
	LUT3 #(
		.INIT('h28)
	) name5268 (
		_w5221_,
		_w5245_,
		_w5333_,
		_w5334_
	);
	LUT3 #(
		.INIT('h41)
	) name5269 (
		_w5221_,
		_w5245_,
		_w5333_,
		_w5335_
	);
	LUT3 #(
		.INIT('h96)
	) name5270 (
		_w5221_,
		_w5245_,
		_w5333_,
		_w5336_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5271 (
		_w4866_,
		_w4981_,
		_w4983_,
		_w5218_,
		_w5337_
	);
	LUT2 #(
		.INIT('h4)
	) name5272 (
		_w5099_,
		_w5337_,
		_w5338_
	);
	LUT3 #(
		.INIT('h31)
	) name5273 (
		_w5100_,
		_w5217_,
		_w5218_,
		_w5339_
	);
	LUT4 #(
		.INIT('h40cc)
	) name5274 (
		_w4994_,
		_w5336_,
		_w5338_,
		_w5339_,
		_w5340_
	);
	LUT4 #(
		.INIT('h0031)
	) name5275 (
		_w5100_,
		_w5217_,
		_w5218_,
		_w5336_,
		_w5341_
	);
	LUT3 #(
		.INIT('hb0)
	) name5276 (
		_w4994_,
		_w5338_,
		_w5341_,
		_w5342_
	);
	LUT2 #(
		.INIT('he)
	) name5277 (
		_w5340_,
		_w5342_,
		_w5343_
	);
	LUT4 #(
		.INIT('h0031)
	) name5278 (
		_w5100_,
		_w5217_,
		_w5218_,
		_w5334_,
		_w5344_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5279 (
		_w5026_,
		_w5028_,
		_w5208_,
		_w5262_,
		_w5345_
	);
	LUT2 #(
		.INIT('h4)
	) name5280 (
		_w5246_,
		_w5345_,
		_w5346_
	);
	LUT4 #(
		.INIT('he100)
	) name5281 (
		_w5209_,
		_w5246_,
		_w5262_,
		_w5332_,
		_w5347_
	);
	LUT3 #(
		.INIT('h51)
	) name5282 (
		_w5293_,
		_w5330_,
		_w5331_,
		_w5348_
	);
	LUT4 #(
		.INIT('hef0e)
	) name5283 (
		_w5136_,
		_w5138_,
		_w5256_,
		_w5260_,
		_w5349_
	);
	LUT3 #(
		.INIT('h2b)
	) name5284 (
		_w5257_,
		_w5258_,
		_w5259_,
		_w5350_
	);
	LUT4 #(
		.INIT('h153f)
	) name5285 (
		\a[30] ,
		\a[31] ,
		\a[41] ,
		\a[42] ,
		_w5351_
	);
	LUT2 #(
		.INIT('h8)
	) name5286 (
		\a[31] ,
		\a[42] ,
		_w5352_
	);
	LUT4 #(
		.INIT('h8000)
	) name5287 (
		\a[30] ,
		\a[31] ,
		\a[41] ,
		\a[42] ,
		_w5353_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5288 (
		\a[30] ,
		\a[31] ,
		\a[41] ,
		\a[42] ,
		_w5354_
	);
	LUT2 #(
		.INIT('h6)
	) name5289 (
		_w5311_,
		_w5354_,
		_w5355_
	);
	LUT4 #(
		.INIT('h7100)
	) name5290 (
		_w5265_,
		_w5266_,
		_w5270_,
		_w5355_,
		_w5356_
	);
	LUT4 #(
		.INIT('h008e)
	) name5291 (
		_w5265_,
		_w5266_,
		_w5270_,
		_w5355_,
		_w5357_
	);
	LUT3 #(
		.INIT('ha9)
	) name5292 (
		_w5350_,
		_w5356_,
		_w5357_,
		_w5358_
	);
	LUT2 #(
		.INIT('h6)
	) name5293 (
		_w5349_,
		_w5358_,
		_w5359_
	);
	LUT4 #(
		.INIT('h001b)
	) name5294 (
		_w5264_,
		_w5289_,
		_w5290_,
		_w5291_,
		_w5360_
	);
	LUT2 #(
		.INIT('h9)
	) name5295 (
		_w5359_,
		_w5360_,
		_w5361_
	);
	LUT3 #(
		.INIT('h2b)
	) name5296 (
		_w5248_,
		_w5252_,
		_w5261_,
		_w5362_
	);
	LUT2 #(
		.INIT('h2)
	) name5297 (
		_w5361_,
		_w5362_,
		_w5363_
	);
	LUT2 #(
		.INIT('h9)
	) name5298 (
		_w5361_,
		_w5362_,
		_w5364_
	);
	LUT2 #(
		.INIT('h9)
	) name5299 (
		_w5348_,
		_w5364_,
		_w5365_
	);
	LUT4 #(
		.INIT('h0bb0)
	) name5300 (
		_w5246_,
		_w5345_,
		_w5348_,
		_w5364_,
		_w5366_
	);
	LUT2 #(
		.INIT('h4)
	) name5301 (
		_w5347_,
		_w5366_,
		_w5367_
	);
	LUT4 #(
		.INIT('h0eef)
	) name5302 (
		_w5209_,
		_w5246_,
		_w5262_,
		_w5332_,
		_w5368_
	);
	LUT2 #(
		.INIT('h2)
	) name5303 (
		_w5365_,
		_w5368_,
		_w5369_
	);
	LUT3 #(
		.INIT('h1e)
	) name5304 (
		_w5346_,
		_w5347_,
		_w5365_,
		_w5370_
	);
	LUT3 #(
		.INIT('h23)
	) name5305 (
		_w5228_,
		_w5240_,
		_w5241_,
		_w5371_
	);
	LUT3 #(
		.INIT('h17)
	) name5306 (
		_w5253_,
		_w5254_,
		_w5255_,
		_w5372_
	);
	LUT3 #(
		.INIT('h32)
	) name5307 (
		_w5319_,
		_w5320_,
		_w5326_,
		_w5373_
	);
	LUT3 #(
		.INIT('h32)
	) name5308 (
		_w5280_,
		_w5281_,
		_w5287_,
		_w5374_
	);
	LUT3 #(
		.INIT('h96)
	) name5309 (
		_w5372_,
		_w5373_,
		_w5374_,
		_w5375_
	);
	LUT3 #(
		.INIT('h0d)
	) name5310 (
		_w5297_,
		_w5307_,
		_w5308_,
		_w5376_
	);
	LUT3 #(
		.INIT('h0d)
	) name5311 (
		_w5322_,
		_w5323_,
		_w5324_,
		_w5377_
	);
	LUT3 #(
		.INIT('h0d)
	) name5312 (
		_w5144_,
		_w5310_,
		_w5312_,
		_w5378_
	);
	LUT3 #(
		.INIT('h0d)
	) name5313 (
		_w5314_,
		_w5315_,
		_w5317_,
		_w5379_
	);
	LUT3 #(
		.INIT('h96)
	) name5314 (
		_w5377_,
		_w5378_,
		_w5379_,
		_w5380_
	);
	LUT3 #(
		.INIT('h0d)
	) name5315 (
		_w5276_,
		_w5277_,
		_w5278_,
		_w5381_
	);
	LUT3 #(
		.INIT('h32)
	) name5316 (
		_w5283_,
		_w5284_,
		_w5285_,
		_w5382_
	);
	LUT3 #(
		.INIT('h0d)
	) name5317 (
		_w5272_,
		_w5273_,
		_w5274_,
		_w5383_
	);
	LUT3 #(
		.INIT('h69)
	) name5318 (
		_w5381_,
		_w5382_,
		_w5383_,
		_w5384_
	);
	LUT3 #(
		.INIT('h96)
	) name5319 (
		_w5376_,
		_w5380_,
		_w5384_,
		_w5385_
	);
	LUT4 #(
		.INIT('he11e)
	) name5320 (
		_w5327_,
		_w5329_,
		_w5375_,
		_w5385_,
		_w5386_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5321 (
		_w5228_,
		_w5238_,
		_w5239_,
		_w5386_,
		_w5387_
	);
	LUT3 #(
		.INIT('h32)
	) name5322 (
		_w5234_,
		_w5235_,
		_w5237_,
		_w5388_
	);
	LUT3 #(
		.INIT('h71)
	) name5323 (
		_w5229_,
		_w5230_,
		_w5231_,
		_w5389_
	);
	LUT4 #(
		.INIT('h153f)
	) name5324 (
		\a[14] ,
		\a[15] ,
		\a[57] ,
		\a[58] ,
		_w5390_
	);
	LUT4 #(
		.INIT('h8000)
	) name5325 (
		\a[14] ,
		\a[15] ,
		\a[57] ,
		\a[58] ,
		_w5391_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5326 (
		\a[14] ,
		\a[15] ,
		\a[57] ,
		\a[58] ,
		_w5392_
	);
	LUT4 #(
		.INIT('h153f)
	) name5327 (
		\a[27] ,
		\a[28] ,
		\a[44] ,
		\a[45] ,
		_w5393_
	);
	LUT2 #(
		.INIT('h8)
	) name5328 (
		\a[28] ,
		\a[45] ,
		_w5394_
	);
	LUT4 #(
		.INIT('h8000)
	) name5329 (
		\a[27] ,
		\a[28] ,
		\a[44] ,
		\a[45] ,
		_w5395_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5330 (
		\a[27] ,
		\a[28] ,
		\a[44] ,
		\a[45] ,
		_w5396_
	);
	LUT4 #(
		.INIT('h1248)
	) name5331 (
		_w5294_,
		_w5304_,
		_w5392_,
		_w5396_,
		_w5397_
	);
	LUT4 #(
		.INIT('h8421)
	) name5332 (
		_w5294_,
		_w5304_,
		_w5392_,
		_w5396_,
		_w5398_
	);
	LUT4 #(
		.INIT('h6996)
	) name5333 (
		_w5294_,
		_w5304_,
		_w5392_,
		_w5396_,
		_w5399_
	);
	LUT2 #(
		.INIT('h8)
	) name5334 (
		\a[19] ,
		\a[53] ,
		_w5400_
	);
	LUT4 #(
		.INIT('h153f)
	) name5335 (
		\a[33] ,
		\a[34] ,
		\a[38] ,
		\a[39] ,
		_w5401_
	);
	LUT2 #(
		.INIT('h8)
	) name5336 (
		\a[34] ,
		\a[39] ,
		_w5402_
	);
	LUT4 #(
		.INIT('h8000)
	) name5337 (
		\a[33] ,
		\a[34] ,
		\a[38] ,
		\a[39] ,
		_w5403_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5338 (
		\a[33] ,
		\a[34] ,
		\a[38] ,
		\a[39] ,
		_w5404_
	);
	LUT2 #(
		.INIT('h6)
	) name5339 (
		_w5400_,
		_w5404_,
		_w5405_
	);
	LUT2 #(
		.INIT('h6)
	) name5340 (
		_w5399_,
		_w5405_,
		_w5406_
	);
	LUT3 #(
		.INIT('h0d)
	) name5341 (
		_w5302_,
		_w5303_,
		_w5305_,
		_w5407_
	);
	LUT3 #(
		.INIT('h0d)
	) name5342 (
		_w5298_,
		_w5299_,
		_w5300_,
		_w5408_
	);
	LUT3 #(
		.INIT('h0d)
	) name5343 (
		_w5173_,
		_w5267_,
		_w5268_,
		_w5409_
	);
	LUT3 #(
		.INIT('h96)
	) name5344 (
		_w5407_,
		_w5408_,
		_w5409_,
		_w5410_
	);
	LUT4 #(
		.INIT('h7100)
	) name5345 (
		_w5229_,
		_w5230_,
		_w5231_,
		_w5410_,
		_w5411_
	);
	LUT4 #(
		.INIT('hde16)
	) name5346 (
		_w5389_,
		_w5406_,
		_w5410_,
		_w5411_,
		_w5412_
	);
	LUT4 #(
		.INIT('h008e)
	) name5347 (
		_w5232_,
		_w5233_,
		_w5237_,
		_w5412_,
		_w5413_
	);
	LUT3 #(
		.INIT('he8)
	) name5348 (
		_w5249_,
		_w5250_,
		_w5251_,
		_w5414_
	);
	LUT4 #(
		.INIT('h153f)
	) name5349 (
		\a[12] ,
		\a[13] ,
		\a[58] ,
		\a[59] ,
		_w5415_
	);
	LUT4 #(
		.INIT('h000d)
	) name5350 (
		_w5150_,
		_w5151_,
		_w5152_,
		_w5295_,
		_w5416_
	);
	LUT2 #(
		.INIT('h8)
	) name5351 (
		\a[12] ,
		\a[60] ,
		_w5417_
	);
	LUT4 #(
		.INIT('h153f)
	) name5352 (
		\a[24] ,
		\a[25] ,
		\a[47] ,
		\a[48] ,
		_w5418_
	);
	LUT2 #(
		.INIT('h8)
	) name5353 (
		\a[25] ,
		\a[48] ,
		_w5419_
	);
	LUT4 #(
		.INIT('h8000)
	) name5354 (
		\a[24] ,
		\a[25] ,
		\a[47] ,
		\a[48] ,
		_w5420_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5355 (
		\a[24] ,
		\a[25] ,
		\a[47] ,
		\a[48] ,
		_w5421_
	);
	LUT2 #(
		.INIT('h6)
	) name5356 (
		_w5417_,
		_w5421_,
		_w5422_
	);
	LUT2 #(
		.INIT('h8)
	) name5357 (
		\a[9] ,
		\a[63] ,
		_w5423_
	);
	LUT4 #(
		.INIT('h153f)
	) name5358 (
		\a[10] ,
		\a[11] ,
		\a[61] ,
		\a[62] ,
		_w5424_
	);
	LUT4 #(
		.INIT('h8000)
	) name5359 (
		\a[10] ,
		\a[11] ,
		\a[61] ,
		\a[62] ,
		_w5425_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5360 (
		\a[10] ,
		\a[11] ,
		\a[61] ,
		\a[62] ,
		_w5426_
	);
	LUT2 #(
		.INIT('h6)
	) name5361 (
		_w5423_,
		_w5426_,
		_w5427_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5362 (
		_w5415_,
		_w5416_,
		_w5422_,
		_w5427_,
		_w5428_
	);
	LUT4 #(
		.INIT('h153f)
	) name5363 (
		\a[16] ,
		\a[23] ,
		\a[49] ,
		\a[56] ,
		_w5429_
	);
	LUT4 #(
		.INIT('h8000)
	) name5364 (
		\a[16] ,
		\a[23] ,
		\a[49] ,
		\a[56] ,
		_w5430_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5365 (
		\a[16] ,
		\a[23] ,
		\a[49] ,
		\a[56] ,
		_w5431_
	);
	LUT2 #(
		.INIT('h8)
	) name5366 (
		\a[35] ,
		\a[37] ,
		_w5432_
	);
	LUT4 #(
		.INIT('h153f)
	) name5367 (
		\a[21] ,
		\a[22] ,
		\a[50] ,
		\a[51] ,
		_w5433_
	);
	LUT2 #(
		.INIT('h8)
	) name5368 (
		\a[22] ,
		\a[51] ,
		_w5434_
	);
	LUT4 #(
		.INIT('h8000)
	) name5369 (
		\a[21] ,
		\a[22] ,
		\a[50] ,
		\a[51] ,
		_w5435_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5370 (
		\a[21] ,
		\a[22] ,
		\a[50] ,
		\a[51] ,
		_w5436_
	);
	LUT4 #(
		.INIT('h0660)
	) name5371 (
		_w5316_,
		_w5431_,
		_w5432_,
		_w5436_,
		_w5437_
	);
	LUT4 #(
		.INIT('h9009)
	) name5372 (
		_w5316_,
		_w5431_,
		_w5432_,
		_w5436_,
		_w5438_
	);
	LUT4 #(
		.INIT('h6996)
	) name5373 (
		_w5316_,
		_w5431_,
		_w5432_,
		_w5436_,
		_w5439_
	);
	LUT2 #(
		.INIT('h8)
	) name5374 (
		\a[17] ,
		\a[55] ,
		_w5440_
	);
	LUT4 #(
		.INIT('h153f)
	) name5375 (
		\a[18] ,
		\a[20] ,
		\a[52] ,
		\a[54] ,
		_w5441_
	);
	LUT2 #(
		.INIT('h8)
	) name5376 (
		\a[20] ,
		\a[54] ,
		_w5442_
	);
	LUT4 #(
		.INIT('h8000)
	) name5377 (
		\a[18] ,
		\a[20] ,
		\a[52] ,
		\a[54] ,
		_w5443_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5378 (
		\a[18] ,
		\a[20] ,
		\a[52] ,
		\a[54] ,
		_w5444_
	);
	LUT2 #(
		.INIT('h6)
	) name5379 (
		_w5440_,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('h6)
	) name5380 (
		_w5439_,
		_w5445_,
		_w5446_
	);
	LUT2 #(
		.INIT('h8)
	) name5381 (
		_w5428_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h1)
	) name5382 (
		_w5428_,
		_w5446_,
		_w5448_
	);
	LUT2 #(
		.INIT('h6)
	) name5383 (
		_w5428_,
		_w5446_,
		_w5449_
	);
	LUT2 #(
		.INIT('h6)
	) name5384 (
		_w5414_,
		_w5449_,
		_w5450_
	);
	LUT4 #(
		.INIT('h7100)
	) name5385 (
		_w5232_,
		_w5233_,
		_w5237_,
		_w5412_,
		_w5451_
	);
	LUT4 #(
		.INIT('hf616)
	) name5386 (
		_w5388_,
		_w5412_,
		_w5450_,
		_w5451_,
		_w5452_
	);
	LUT3 #(
		.INIT('h0d)
	) name5387 (
		_w5238_,
		_w5239_,
		_w5386_,
		_w5453_
	);
	LUT4 #(
		.INIT('h40f0)
	) name5388 (
		_w5228_,
		_w5241_,
		_w5452_,
		_w5453_,
		_w5454_
	);
	LUT4 #(
		.INIT('h40f9)
	) name5389 (
		_w5371_,
		_w5386_,
		_w5452_,
		_w5454_,
		_w5455_
	);
	LUT3 #(
		.INIT('h70)
	) name5390 (
		_w5242_,
		_w5244_,
		_w5333_,
		_w5456_
	);
	LUT4 #(
		.INIT('h0101)
	) name5391 (
		_w5222_,
		_w5224_,
		_w5242_,
		_w5244_,
		_w5457_
	);
	LUT4 #(
		.INIT('h9990)
	) name5392 (
		_w5370_,
		_w5455_,
		_w5456_,
		_w5457_,
		_w5458_
	);
	LUT4 #(
		.INIT('h0006)
	) name5393 (
		_w5370_,
		_w5455_,
		_w5456_,
		_w5457_,
		_w5459_
	);
	LUT4 #(
		.INIT('h6669)
	) name5394 (
		_w5370_,
		_w5455_,
		_w5456_,
		_w5457_,
		_w5460_
	);
	LUT2 #(
		.INIT('h4)
	) name5395 (
		_w5335_,
		_w5460_,
		_w5461_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5396 (
		_w4994_,
		_w5338_,
		_w5344_,
		_w5461_,
		_w5462_
	);
	LUT4 #(
		.INIT('h1033)
	) name5397 (
		_w4994_,
		_w5335_,
		_w5338_,
		_w5344_,
		_w5463_
	);
	LUT3 #(
		.INIT('hcd)
	) name5398 (
		_w5460_,
		_w5462_,
		_w5463_,
		_w5464_
	);
	LUT2 #(
		.INIT('h1)
	) name5399 (
		_w5335_,
		_w5459_,
		_w5465_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5400 (
		_w4994_,
		_w5338_,
		_w5344_,
		_w5465_,
		_w5466_
	);
	LUT3 #(
		.INIT('h54)
	) name5401 (
		_w5367_,
		_w5369_,
		_w5455_,
		_w5467_
	);
	LUT4 #(
		.INIT('h011f)
	) name5402 (
		_w5327_,
		_w5329_,
		_w5375_,
		_w5385_,
		_w5468_
	);
	LUT2 #(
		.INIT('h2)
	) name5403 (
		_w5406_,
		_w5410_,
		_w5469_
	);
	LUT2 #(
		.INIT('h8)
	) name5404 (
		_w5406_,
		_w5410_,
		_w5470_
	);
	LUT4 #(
		.INIT('h0071)
	) name5405 (
		_w5229_,
		_w5230_,
		_w5231_,
		_w5410_,
		_w5471_
	);
	LUT4 #(
		.INIT('h001b)
	) name5406 (
		_w5389_,
		_w5469_,
		_w5470_,
		_w5471_,
		_w5472_
	);
	LUT3 #(
		.INIT('h17)
	) name5407 (
		_w5377_,
		_w5378_,
		_w5379_,
		_w5473_
	);
	LUT4 #(
		.INIT('h153f)
	) name5408 (
		\a[32] ,
		\a[33] ,
		\a[40] ,
		\a[41] ,
		_w5474_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		\a[33] ,
		\a[41] ,
		_w5475_
	);
	LUT4 #(
		.INIT('h8000)
	) name5410 (
		\a[32] ,
		\a[33] ,
		\a[40] ,
		\a[41] ,
		_w5476_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5411 (
		\a[32] ,
		\a[33] ,
		\a[40] ,
		\a[41] ,
		_w5477_
	);
	LUT2 #(
		.INIT('h6)
	) name5412 (
		_w5352_,
		_w5477_,
		_w5478_
	);
	LUT4 #(
		.INIT('h1700)
	) name5413 (
		_w5407_,
		_w5408_,
		_w5409_,
		_w5478_,
		_w5479_
	);
	LUT4 #(
		.INIT('h00e8)
	) name5414 (
		_w5407_,
		_w5408_,
		_w5409_,
		_w5478_,
		_w5480_
	);
	LUT3 #(
		.INIT('ha9)
	) name5415 (
		_w5473_,
		_w5479_,
		_w5480_,
		_w5481_
	);
	LUT3 #(
		.INIT('h2b)
	) name5416 (
		_w5376_,
		_w5380_,
		_w5384_,
		_w5482_
	);
	LUT2 #(
		.INIT('h6)
	) name5417 (
		_w5481_,
		_w5482_,
		_w5483_
	);
	LUT3 #(
		.INIT('h41)
	) name5418 (
		_w5468_,
		_w5472_,
		_w5483_,
		_w5484_
	);
	LUT3 #(
		.INIT('h96)
	) name5419 (
		_w5468_,
		_w5472_,
		_w5483_,
		_w5485_
	);
	LUT4 #(
		.INIT('hae00)
	) name5420 (
		_w5413_,
		_w5450_,
		_w5451_,
		_w5485_,
		_w5486_
	);
	LUT4 #(
		.INIT('h51ae)
	) name5421 (
		_w5413_,
		_w5450_,
		_w5451_,
		_w5485_,
		_w5487_
	);
	LUT3 #(
		.INIT('he0)
	) name5422 (
		_w5387_,
		_w5454_,
		_w5487_,
		_w5488_
	);
	LUT3 #(
		.INIT('h1e)
	) name5423 (
		_w5387_,
		_w5454_,
		_w5487_,
		_w5489_
	);
	LUT3 #(
		.INIT('h31)
	) name5424 (
		_w5414_,
		_w5447_,
		_w5448_,
		_w5490_
	);
	LUT4 #(
		.INIT('hf110)
	) name5425 (
		_w5415_,
		_w5416_,
		_w5422_,
		_w5427_,
		_w5491_
	);
	LUT3 #(
		.INIT('h4d)
	) name5426 (
		_w5381_,
		_w5382_,
		_w5383_,
		_w5492_
	);
	LUT3 #(
		.INIT('h32)
	) name5427 (
		_w5397_,
		_w5398_,
		_w5405_,
		_w5493_
	);
	LUT3 #(
		.INIT('h96)
	) name5428 (
		_w5491_,
		_w5492_,
		_w5493_,
		_w5494_
	);
	LUT3 #(
		.INIT('h32)
	) name5429 (
		_w5437_,
		_w5438_,
		_w5445_,
		_w5495_
	);
	LUT2 #(
		.INIT('h8)
	) name5430 (
		\a[13] ,
		\a[60] ,
		_w5496_
	);
	LUT4 #(
		.INIT('h0dff)
	) name5431 (
		_w5432_,
		_w5433_,
		_w5435_,
		_w5496_,
		_w5497_
	);
	LUT4 #(
		.INIT('h0df2)
	) name5432 (
		_w5432_,
		_w5433_,
		_w5435_,
		_w5496_,
		_w5498_
	);
	LUT3 #(
		.INIT('h0d)
	) name5433 (
		_w5400_,
		_w5401_,
		_w5403_,
		_w5499_
	);
	LUT2 #(
		.INIT('h6)
	) name5434 (
		_w5498_,
		_w5499_,
		_w5500_
	);
	LUT3 #(
		.INIT('h0d)
	) name5435 (
		_w5417_,
		_w5418_,
		_w5420_,
		_w5501_
	);
	LUT3 #(
		.INIT('h0d)
	) name5436 (
		_w5423_,
		_w5424_,
		_w5425_,
		_w5502_
	);
	LUT3 #(
		.INIT('h0d)
	) name5437 (
		_w5440_,
		_w5441_,
		_w5443_,
		_w5503_
	);
	LUT3 #(
		.INIT('h96)
	) name5438 (
		_w5501_,
		_w5502_,
		_w5503_,
		_w5504_
	);
	LUT3 #(
		.INIT('h96)
	) name5439 (
		_w5495_,
		_w5500_,
		_w5504_,
		_w5505_
	);
	LUT3 #(
		.INIT('h69)
	) name5440 (
		_w5490_,
		_w5494_,
		_w5505_,
		_w5506_
	);
	LUT3 #(
		.INIT('h0d)
	) name5441 (
		_w5361_,
		_w5362_,
		_w5506_,
		_w5507_
	);
	LUT3 #(
		.INIT('hb0)
	) name5442 (
		_w5348_,
		_w5364_,
		_w5507_,
		_w5508_
	);
	LUT3 #(
		.INIT('h0d)
	) name5443 (
		_w5304_,
		_w5393_,
		_w5395_,
		_w5509_
	);
	LUT3 #(
		.INIT('h0d)
	) name5444 (
		_w5294_,
		_w5390_,
		_w5391_,
		_w5510_
	);
	LUT3 #(
		.INIT('h0d)
	) name5445 (
		_w5311_,
		_w5351_,
		_w5353_,
		_w5511_
	);
	LUT3 #(
		.INIT('h96)
	) name5446 (
		_w5509_,
		_w5510_,
		_w5511_,
		_w5512_
	);
	LUT4 #(
		.INIT('hff31)
	) name5447 (
		_w5350_,
		_w5356_,
		_w5357_,
		_w5512_,
		_w5513_
	);
	LUT4 #(
		.INIT('hce31)
	) name5448 (
		_w5350_,
		_w5356_,
		_w5357_,
		_w5512_,
		_w5514_
	);
	LUT4 #(
		.INIT('h153f)
	) name5449 (
		\a[10] ,
		\a[12] ,
		\a[61] ,
		\a[63] ,
		_w5515_
	);
	LUT4 #(
		.INIT('h8000)
	) name5450 (
		\a[10] ,
		\a[12] ,
		\a[61] ,
		\a[63] ,
		_w5516_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5451 (
		\a[10] ,
		\a[12] ,
		\a[61] ,
		\a[63] ,
		_w5517_
	);
	LUT4 #(
		.INIT('h153f)
	) name5452 (
		\a[29] ,
		\a[30] ,
		\a[43] ,
		\a[44] ,
		_w5518_
	);
	LUT4 #(
		.INIT('h8000)
	) name5453 (
		\a[29] ,
		\a[30] ,
		\a[43] ,
		\a[44] ,
		_w5519_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5454 (
		\a[29] ,
		\a[30] ,
		\a[43] ,
		\a[44] ,
		_w5520_
	);
	LUT4 #(
		.INIT('h1428)
	) name5455 (
		_w5394_,
		_w5419_,
		_w5517_,
		_w5520_,
		_w5521_
	);
	LUT4 #(
		.INIT('h8241)
	) name5456 (
		_w5394_,
		_w5419_,
		_w5517_,
		_w5520_,
		_w5522_
	);
	LUT4 #(
		.INIT('h6996)
	) name5457 (
		_w5394_,
		_w5419_,
		_w5517_,
		_w5520_,
		_w5523_
	);
	LUT4 #(
		.INIT('h153f)
	) name5458 (
		\a[35] ,
		\a[36] ,
		\a[37] ,
		\a[38] ,
		_w5524_
	);
	LUT2 #(
		.INIT('h8)
	) name5459 (
		\a[36] ,
		\a[38] ,
		_w5525_
	);
	LUT4 #(
		.INIT('h8000)
	) name5460 (
		\a[35] ,
		\a[36] ,
		\a[37] ,
		\a[38] ,
		_w5526_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5461 (
		\a[35] ,
		\a[36] ,
		\a[37] ,
		\a[38] ,
		_w5527_
	);
	LUT2 #(
		.INIT('h6)
	) name5462 (
		_w5402_,
		_w5527_,
		_w5528_
	);
	LUT2 #(
		.INIT('h6)
	) name5463 (
		_w5523_,
		_w5528_,
		_w5529_
	);
	LUT2 #(
		.INIT('h6)
	) name5464 (
		_w5514_,
		_w5529_,
		_w5530_
	);
	LUT4 #(
		.INIT('h8e00)
	) name5465 (
		_w5349_,
		_w5358_,
		_w5360_,
		_w5530_,
		_w5531_
	);
	LUT3 #(
		.INIT('he8)
	) name5466 (
		_w5372_,
		_w5373_,
		_w5374_,
		_w5532_
	);
	LUT2 #(
		.INIT('h8)
	) name5467 (
		\a[18] ,
		\a[55] ,
		_w5533_
	);
	LUT4 #(
		.INIT('h153f)
	) name5468 (
		\a[19] ,
		\a[24] ,
		\a[49] ,
		\a[54] ,
		_w5534_
	);
	LUT4 #(
		.INIT('h8000)
	) name5469 (
		\a[19] ,
		\a[24] ,
		\a[49] ,
		\a[54] ,
		_w5535_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5470 (
		\a[19] ,
		\a[24] ,
		\a[49] ,
		\a[54] ,
		_w5536_
	);
	LUT2 #(
		.INIT('h8)
	) name5471 (
		\a[23] ,
		\a[50] ,
		_w5537_
	);
	LUT3 #(
		.INIT('h13)
	) name5472 (
		\a[11] ,
		\a[37] ,
		\a[62] ,
		_w5538_
	);
	LUT3 #(
		.INIT('h80)
	) name5473 (
		\a[11] ,
		\a[37] ,
		\a[62] ,
		_w5539_
	);
	LUT3 #(
		.INIT('h6c)
	) name5474 (
		\a[11] ,
		\a[37] ,
		\a[62] ,
		_w5540_
	);
	LUT4 #(
		.INIT('h0660)
	) name5475 (
		_w5533_,
		_w5536_,
		_w5537_,
		_w5540_,
		_w5541_
	);
	LUT4 #(
		.INIT('h9009)
	) name5476 (
		_w5533_,
		_w5536_,
		_w5537_,
		_w5540_,
		_w5542_
	);
	LUT4 #(
		.INIT('h6996)
	) name5477 (
		_w5533_,
		_w5536_,
		_w5537_,
		_w5540_,
		_w5543_
	);
	LUT4 #(
		.INIT('h153f)
	) name5478 (
		\a[20] ,
		\a[21] ,
		\a[52] ,
		\a[53] ,
		_w5544_
	);
	LUT4 #(
		.INIT('h8000)
	) name5479 (
		\a[20] ,
		\a[21] ,
		\a[52] ,
		\a[53] ,
		_w5545_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5480 (
		\a[20] ,
		\a[21] ,
		\a[52] ,
		\a[53] ,
		_w5546_
	);
	LUT2 #(
		.INIT('h6)
	) name5481 (
		_w5434_,
		_w5546_,
		_w5547_
	);
	LUT2 #(
		.INIT('h6)
	) name5482 (
		_w5543_,
		_w5547_,
		_w5548_
	);
	LUT3 #(
		.INIT('h32)
	) name5483 (
		_w5316_,
		_w5429_,
		_w5430_,
		_w5549_
	);
	LUT2 #(
		.INIT('h8)
	) name5484 (
		\a[17] ,
		\a[56] ,
		_w5550_
	);
	LUT4 #(
		.INIT('h153f)
	) name5485 (
		\a[26] ,
		\a[27] ,
		\a[46] ,
		\a[47] ,
		_w5551_
	);
	LUT4 #(
		.INIT('h8000)
	) name5486 (
		\a[26] ,
		\a[27] ,
		\a[46] ,
		\a[47] ,
		_w5552_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5487 (
		\a[26] ,
		\a[27] ,
		\a[46] ,
		\a[47] ,
		_w5553_
	);
	LUT2 #(
		.INIT('h6)
	) name5488 (
		_w5550_,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h8)
	) name5489 (
		\a[14] ,
		\a[59] ,
		_w5555_
	);
	LUT4 #(
		.INIT('h153f)
	) name5490 (
		\a[15] ,
		\a[16] ,
		\a[57] ,
		\a[58] ,
		_w5556_
	);
	LUT4 #(
		.INIT('h8000)
	) name5491 (
		\a[15] ,
		\a[16] ,
		\a[57] ,
		\a[58] ,
		_w5557_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5492 (
		\a[15] ,
		\a[16] ,
		\a[57] ,
		\a[58] ,
		_w5558_
	);
	LUT2 #(
		.INIT('h6)
	) name5493 (
		_w5555_,
		_w5558_,
		_w5559_
	);
	LUT3 #(
		.INIT('h69)
	) name5494 (
		_w5549_,
		_w5554_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h2)
	) name5495 (
		_w5548_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('h4)
	) name5496 (
		_w5548_,
		_w5560_,
		_w5562_
	);
	LUT2 #(
		.INIT('h9)
	) name5497 (
		_w5548_,
		_w5560_,
		_w5563_
	);
	LUT2 #(
		.INIT('h6)
	) name5498 (
		_w5532_,
		_w5563_,
		_w5564_
	);
	LUT4 #(
		.INIT('h7007)
	) name5499 (
		_w5349_,
		_w5358_,
		_w5514_,
		_w5529_,
		_w5565_
	);
	LUT3 #(
		.INIT('hd0)
	) name5500 (
		_w5359_,
		_w5360_,
		_w5565_,
		_w5566_
	);
	LUT4 #(
		.INIT('h20f0)
	) name5501 (
		_w5359_,
		_w5360_,
		_w5564_,
		_w5565_,
		_w5567_
	);
	LUT4 #(
		.INIT('h6006)
	) name5502 (
		_w5514_,
		_w5529_,
		_w5532_,
		_w5563_,
		_w5568_
	);
	LUT4 #(
		.INIT('h8e00)
	) name5503 (
		_w5349_,
		_w5358_,
		_w5360_,
		_w5568_,
		_w5569_
	);
	LUT4 #(
		.INIT('h00cb)
	) name5504 (
		_w5531_,
		_w5564_,
		_w5566_,
		_w5569_,
		_w5570_
	);
	LUT2 #(
		.INIT('h4)
	) name5505 (
		_w5506_,
		_w5570_,
		_w5571_
	);
	LUT4 #(
		.INIT('hb200)
	) name5506 (
		_w5348_,
		_w5361_,
		_w5362_,
		_w5570_,
		_w5572_
	);
	LUT3 #(
		.INIT('h54)
	) name5507 (
		_w5508_,
		_w5571_,
		_w5572_,
		_w5573_
	);
	LUT3 #(
		.INIT('h23)
	) name5508 (
		_w5348_,
		_w5363_,
		_w5364_,
		_w5574_
	);
	LUT3 #(
		.INIT('hed)
	) name5509 (
		_w5506_,
		_w5570_,
		_w5574_,
		_w5575_
	);
	LUT3 #(
		.INIT('h9a)
	) name5510 (
		_w5489_,
		_w5573_,
		_w5575_,
		_w5576_
	);
	LUT2 #(
		.INIT('h1)
	) name5511 (
		_w5467_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h6)
	) name5512 (
		_w5467_,
		_w5576_,
		_w5578_
	);
	LUT3 #(
		.INIT('he1)
	) name5513 (
		_w5458_,
		_w5466_,
		_w5578_,
		_w5579_
	);
	LUT4 #(
		.INIT('h0222)
	) name5514 (
		_w5458_,
		_w5459_,
		_w5467_,
		_w5576_,
		_w5580_
	);
	LUT4 #(
		.INIT('h0111)
	) name5515 (
		_w5335_,
		_w5459_,
		_w5467_,
		_w5576_,
		_w5581_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5516 (
		_w4994_,
		_w5338_,
		_w5344_,
		_w5581_,
		_w5582_
	);
	LUT3 #(
		.INIT('h01)
	) name5517 (
		_w5387_,
		_w5454_,
		_w5487_,
		_w5583_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5518 (
		_w5488_,
		_w5573_,
		_w5575_,
		_w5583_,
		_w5584_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5519 (
		_w5348_,
		_w5361_,
		_w5362_,
		_w5506_,
		_w5585_
	);
	LUT3 #(
		.INIT('h17)
	) name5520 (
		_w5501_,
		_w5502_,
		_w5503_,
		_w5586_
	);
	LUT4 #(
		.INIT('h000d)
	) name5521 (
		_w5432_,
		_w5433_,
		_w5435_,
		_w5496_,
		_w5587_
	);
	LUT3 #(
		.INIT('h07)
	) name5522 (
		_w5497_,
		_w5499_,
		_w5587_,
		_w5588_
	);
	LUT3 #(
		.INIT('h17)
	) name5523 (
		_w5549_,
		_w5554_,
		_w5559_,
		_w5589_
	);
	LUT3 #(
		.INIT('h96)
	) name5524 (
		_w5586_,
		_w5588_,
		_w5589_,
		_w5590_
	);
	LUT3 #(
		.INIT('h2b)
	) name5525 (
		_w5495_,
		_w5500_,
		_w5504_,
		_w5591_
	);
	LUT3 #(
		.INIT('he8)
	) name5526 (
		_w5491_,
		_w5492_,
		_w5493_,
		_w5592_
	);
	LUT3 #(
		.INIT('h69)
	) name5527 (
		_w5590_,
		_w5591_,
		_w5592_,
		_w5593_
	);
	LUT4 #(
		.INIT('hd400)
	) name5528 (
		_w5490_,
		_w5494_,
		_w5505_,
		_w5593_,
		_w5594_
	);
	LUT4 #(
		.INIT('h002b)
	) name5529 (
		_w5490_,
		_w5494_,
		_w5505_,
		_w5593_,
		_w5595_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name5530 (
		_w5490_,
		_w5494_,
		_w5505_,
		_w5593_,
		_w5596_
	);
	LUT3 #(
		.INIT('he0)
	) name5531 (
		_w5531_,
		_w5567_,
		_w5596_,
		_w5597_
	);
	LUT3 #(
		.INIT('h1e)
	) name5532 (
		_w5531_,
		_w5567_,
		_w5596_,
		_w5598_
	);
	LUT3 #(
		.INIT('h31)
	) name5533 (
		_w5532_,
		_w5561_,
		_w5562_,
		_w5599_
	);
	LUT4 #(
		.INIT('h3100)
	) name5534 (
		_w5350_,
		_w5356_,
		_w5357_,
		_w5512_,
		_w5600_
	);
	LUT3 #(
		.INIT('h0d)
	) name5535 (
		_w5513_,
		_w5529_,
		_w5600_,
		_w5601_
	);
	LUT3 #(
		.INIT('h32)
	) name5536 (
		_w5541_,
		_w5542_,
		_w5547_,
		_w5602_
	);
	LUT3 #(
		.INIT('h0d)
	) name5537 (
		_w5402_,
		_w5524_,
		_w5526_,
		_w5603_
	);
	LUT3 #(
		.INIT('h0d)
	) name5538 (
		_w5352_,
		_w5474_,
		_w5476_,
		_w5604_
	);
	LUT2 #(
		.INIT('h8)
	) name5539 (
		\a[14] ,
		\a[60] ,
		_w5605_
	);
	LUT4 #(
		.INIT('h153f)
	) name5540 (
		\a[15] ,
		\a[16] ,
		\a[58] ,
		\a[59] ,
		_w5606_
	);
	LUT4 #(
		.INIT('h8000)
	) name5541 (
		\a[15] ,
		\a[16] ,
		\a[58] ,
		\a[59] ,
		_w5607_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5542 (
		\a[15] ,
		\a[16] ,
		\a[58] ,
		\a[59] ,
		_w5608_
	);
	LUT2 #(
		.INIT('h6)
	) name5543 (
		_w5605_,
		_w5608_,
		_w5609_
	);
	LUT3 #(
		.INIT('h69)
	) name5544 (
		_w5603_,
		_w5604_,
		_w5609_,
		_w5610_
	);
	LUT2 #(
		.INIT('h4)
	) name5545 (
		_w5602_,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('h2)
	) name5546 (
		_w5602_,
		_w5610_,
		_w5612_
	);
	LUT2 #(
		.INIT('h9)
	) name5547 (
		_w5602_,
		_w5610_,
		_w5613_
	);
	LUT3 #(
		.INIT('h0e)
	) name5548 (
		_w5473_,
		_w5479_,
		_w5480_,
		_w5614_
	);
	LUT2 #(
		.INIT('h6)
	) name5549 (
		_w5613_,
		_w5614_,
		_w5615_
	);
	LUT3 #(
		.INIT('h69)
	) name5550 (
		_w5599_,
		_w5601_,
		_w5615_,
		_w5616_
	);
	LUT3 #(
		.INIT('he0)
	) name5551 (
		_w5484_,
		_w5486_,
		_w5616_,
		_w5617_
	);
	LUT3 #(
		.INIT('h0d)
	) name5552 (
		_w5550_,
		_w5551_,
		_w5552_,
		_w5618_
	);
	LUT3 #(
		.INIT('h0d)
	) name5553 (
		_w5394_,
		_w5518_,
		_w5519_,
		_w5619_
	);
	LUT3 #(
		.INIT('h0d)
	) name5554 (
		_w5555_,
		_w5556_,
		_w5557_,
		_w5620_
	);
	LUT3 #(
		.INIT('h96)
	) name5555 (
		_w5618_,
		_w5619_,
		_w5620_,
		_w5621_
	);
	LUT3 #(
		.INIT('h0d)
	) name5556 (
		_w5533_,
		_w5534_,
		_w5535_,
		_w5622_
	);
	LUT3 #(
		.INIT('h0d)
	) name5557 (
		_w5434_,
		_w5544_,
		_w5545_,
		_w5623_
	);
	LUT3 #(
		.INIT('h0d)
	) name5558 (
		_w5419_,
		_w5515_,
		_w5516_,
		_w5624_
	);
	LUT3 #(
		.INIT('h96)
	) name5559 (
		_w5622_,
		_w5623_,
		_w5624_,
		_w5625_
	);
	LUT3 #(
		.INIT('h32)
	) name5560 (
		_w5521_,
		_w5522_,
		_w5528_,
		_w5626_
	);
	LUT3 #(
		.INIT('h96)
	) name5561 (
		_w5621_,
		_w5625_,
		_w5626_,
		_w5627_
	);
	LUT4 #(
		.INIT('hd400)
	) name5562 (
		_w5472_,
		_w5481_,
		_w5482_,
		_w5627_,
		_w5628_
	);
	LUT3 #(
		.INIT('h07)
	) name5563 (
		_w5481_,
		_w5482_,
		_w5627_,
		_w5629_
	);
	LUT3 #(
		.INIT('hb0)
	) name5564 (
		_w5472_,
		_w5483_,
		_w5629_,
		_w5630_
	);
	LUT3 #(
		.INIT('h17)
	) name5565 (
		_w5509_,
		_w5510_,
		_w5511_,
		_w5631_
	);
	LUT4 #(
		.INIT('h8000)
	) name5566 (
		\a[12] ,
		\a[13] ,
		\a[61] ,
		\a[62] ,
		_w5632_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5567 (
		\a[12] ,
		\a[13] ,
		\a[61] ,
		\a[62] ,
		_w5633_
	);
	LUT4 #(
		.INIT('hf20d)
	) name5568 (
		_w5537_,
		_w5538_,
		_w5539_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h8)
	) name5569 (
		\a[29] ,
		\a[45] ,
		_w5635_
	);
	LUT4 #(
		.INIT('h153f)
	) name5570 (
		\a[17] ,
		\a[30] ,
		\a[44] ,
		\a[57] ,
		_w5636_
	);
	LUT4 #(
		.INIT('h8000)
	) name5571 (
		\a[17] ,
		\a[30] ,
		\a[44] ,
		\a[57] ,
		_w5637_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5572 (
		\a[17] ,
		\a[30] ,
		\a[44] ,
		\a[57] ,
		_w5638_
	);
	LUT2 #(
		.INIT('h6)
	) name5573 (
		_w5635_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('h4)
	) name5574 (
		_w5634_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h2)
	) name5575 (
		_w5634_,
		_w5639_,
		_w5641_
	);
	LUT2 #(
		.INIT('h9)
	) name5576 (
		_w5634_,
		_w5639_,
		_w5642_
	);
	LUT2 #(
		.INIT('h8)
	) name5577 (
		\a[11] ,
		\a[63] ,
		_w5643_
	);
	LUT4 #(
		.INIT('h153f)
	) name5578 (
		\a[31] ,
		\a[32] ,
		\a[42] ,
		\a[43] ,
		_w5644_
	);
	LUT4 #(
		.INIT('h8000)
	) name5579 (
		\a[31] ,
		\a[32] ,
		\a[42] ,
		\a[43] ,
		_w5645_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5580 (
		\a[31] ,
		\a[32] ,
		\a[42] ,
		\a[43] ,
		_w5646_
	);
	LUT4 #(
		.INIT('h153f)
	) name5581 (
		\a[18] ,
		\a[25] ,
		\a[49] ,
		\a[56] ,
		_w5647_
	);
	LUT4 #(
		.INIT('h8000)
	) name5582 (
		\a[18] ,
		\a[25] ,
		\a[49] ,
		\a[56] ,
		_w5648_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5583 (
		\a[18] ,
		\a[25] ,
		\a[49] ,
		\a[56] ,
		_w5649_
	);
	LUT4 #(
		.INIT('h1428)
	) name5584 (
		_w5475_,
		_w5643_,
		_w5646_,
		_w5649_,
		_w5650_
	);
	LUT4 #(
		.INIT('h8241)
	) name5585 (
		_w5475_,
		_w5643_,
		_w5646_,
		_w5649_,
		_w5651_
	);
	LUT4 #(
		.INIT('h6996)
	) name5586 (
		_w5475_,
		_w5643_,
		_w5646_,
		_w5649_,
		_w5652_
	);
	LUT2 #(
		.INIT('h8)
	) name5587 (
		\a[26] ,
		\a[48] ,
		_w5653_
	);
	LUT4 #(
		.INIT('h153f)
	) name5588 (
		\a[27] ,
		\a[28] ,
		\a[46] ,
		\a[47] ,
		_w5654_
	);
	LUT4 #(
		.INIT('h8000)
	) name5589 (
		\a[27] ,
		\a[28] ,
		\a[46] ,
		\a[47] ,
		_w5655_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5590 (
		\a[27] ,
		\a[28] ,
		\a[46] ,
		\a[47] ,
		_w5656_
	);
	LUT2 #(
		.INIT('h6)
	) name5591 (
		_w5653_,
		_w5656_,
		_w5657_
	);
	LUT2 #(
		.INIT('h8)
	) name5592 (
		\a[22] ,
		\a[52] ,
		_w5658_
	);
	LUT4 #(
		.INIT('h153f)
	) name5593 (
		\a[19] ,
		\a[21] ,
		\a[53] ,
		\a[55] ,
		_w5659_
	);
	LUT4 #(
		.INIT('h8000)
	) name5594 (
		\a[19] ,
		\a[21] ,
		\a[53] ,
		\a[55] ,
		_w5660_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5595 (
		\a[19] ,
		\a[21] ,
		\a[53] ,
		\a[55] ,
		_w5661_
	);
	LUT4 #(
		.INIT('h153f)
	) name5596 (
		\a[34] ,
		\a[35] ,
		\a[39] ,
		\a[40] ,
		_w5662_
	);
	LUT4 #(
		.INIT('h8000)
	) name5597 (
		\a[34] ,
		\a[35] ,
		\a[39] ,
		\a[40] ,
		_w5663_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5598 (
		\a[34] ,
		\a[35] ,
		\a[39] ,
		\a[40] ,
		_w5664_
	);
	LUT4 #(
		.INIT('h1428)
	) name5599 (
		_w5442_,
		_w5658_,
		_w5661_,
		_w5664_,
		_w5665_
	);
	LUT4 #(
		.INIT('h8241)
	) name5600 (
		_w5442_,
		_w5658_,
		_w5661_,
		_w5664_,
		_w5666_
	);
	LUT4 #(
		.INIT('h6996)
	) name5601 (
		_w5442_,
		_w5658_,
		_w5661_,
		_w5664_,
		_w5667_
	);
	LUT4 #(
		.INIT('h153f)
	) name5602 (
		\a[23] ,
		\a[24] ,
		\a[50] ,
		\a[51] ,
		_w5668_
	);
	LUT4 #(
		.INIT('h8000)
	) name5603 (
		\a[23] ,
		\a[24] ,
		\a[50] ,
		\a[51] ,
		_w5669_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5604 (
		\a[23] ,
		\a[24] ,
		\a[50] ,
		\a[51] ,
		_w5670_
	);
	LUT2 #(
		.INIT('h6)
	) name5605 (
		_w5525_,
		_w5670_,
		_w5671_
	);
	LUT4 #(
		.INIT('h0660)
	) name5606 (
		_w5652_,
		_w5657_,
		_w5667_,
		_w5671_,
		_w5672_
	);
	LUT4 #(
		.INIT('h9009)
	) name5607 (
		_w5652_,
		_w5657_,
		_w5667_,
		_w5671_,
		_w5673_
	);
	LUT4 #(
		.INIT('h6996)
	) name5608 (
		_w5652_,
		_w5657_,
		_w5667_,
		_w5671_,
		_w5674_
	);
	LUT3 #(
		.INIT('h96)
	) name5609 (
		_w5631_,
		_w5642_,
		_w5674_,
		_w5675_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5610 (
		_w5472_,
		_w5483_,
		_w5629_,
		_w5675_,
		_w5676_
	);
	LUT2 #(
		.INIT('h2)
	) name5611 (
		_w5627_,
		_w5675_,
		_w5677_
	);
	LUT4 #(
		.INIT('hd400)
	) name5612 (
		_w5472_,
		_w5481_,
		_w5482_,
		_w5677_,
		_w5678_
	);
	LUT4 #(
		.INIT('h00e3)
	) name5613 (
		_w5628_,
		_w5630_,
		_w5675_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h1)
	) name5614 (
		_w5484_,
		_w5616_,
		_w5680_
	);
	LUT3 #(
		.INIT('h8c)
	) name5615 (
		_w5486_,
		_w5679_,
		_w5680_,
		_w5681_
	);
	LUT4 #(
		.INIT('he11e)
	) name5616 (
		_w5484_,
		_w5486_,
		_w5616_,
		_w5679_,
		_w5682_
	);
	LUT4 #(
		.INIT('h1e00)
	) name5617 (
		_w5573_,
		_w5585_,
		_w5598_,
		_w5682_,
		_w5683_
	);
	LUT4 #(
		.INIT('h00e1)
	) name5618 (
		_w5573_,
		_w5585_,
		_w5598_,
		_w5682_,
		_w5684_
	);
	LUT4 #(
		.INIT('he11e)
	) name5619 (
		_w5573_,
		_w5585_,
		_w5598_,
		_w5682_,
		_w5685_
	);
	LUT2 #(
		.INIT('h1)
	) name5620 (
		_w5584_,
		_w5685_,
		_w5686_
	);
	LUT3 #(
		.INIT('h02)
	) name5621 (
		_w5584_,
		_w5683_,
		_w5684_,
		_w5687_
	);
	LUT3 #(
		.INIT('h01)
	) name5622 (
		_w5577_,
		_w5686_,
		_w5687_,
		_w5688_
	);
	LUT3 #(
		.INIT('h10)
	) name5623 (
		_w5580_,
		_w5582_,
		_w5688_,
		_w5689_
	);
	LUT3 #(
		.INIT('ha9)
	) name5624 (
		_w5584_,
		_w5683_,
		_w5684_,
		_w5690_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5625 (
		_w5577_,
		_w5580_,
		_w5582_,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('h1)
	) name5626 (
		_w5689_,
		_w5691_,
		_w5692_
	);
	LUT4 #(
		.INIT('heee0)
	) name5627 (
		_w5467_,
		_w5576_,
		_w5584_,
		_w5685_,
		_w5693_
	);
	LUT4 #(
		.INIT('h011f)
	) name5628 (
		_w5573_,
		_w5585_,
		_w5598_,
		_w5682_,
		_w5694_
	);
	LUT4 #(
		.INIT('h0f01)
	) name5629 (
		_w5531_,
		_w5567_,
		_w5594_,
		_w5595_,
		_w5695_
	);
	LUT3 #(
		.INIT('h17)
	) name5630 (
		_w5622_,
		_w5623_,
		_w5624_,
		_w5696_
	);
	LUT3 #(
		.INIT('h8e)
	) name5631 (
		_w5603_,
		_w5604_,
		_w5609_,
		_w5697_
	);
	LUT3 #(
		.INIT('h17)
	) name5632 (
		_w5618_,
		_w5619_,
		_w5620_,
		_w5698_
	);
	LUT3 #(
		.INIT('h69)
	) name5633 (
		_w5696_,
		_w5697_,
		_w5698_,
		_w5699_
	);
	LUT4 #(
		.INIT('h00f6)
	) name5634 (
		_w5631_,
		_w5642_,
		_w5672_,
		_w5673_,
		_w5700_
	);
	LUT3 #(
		.INIT('h0e)
	) name5635 (
		_w5631_,
		_w5640_,
		_w5641_,
		_w5701_
	);
	LUT3 #(
		.INIT('h0d)
	) name5636 (
		_w5442_,
		_w5662_,
		_w5663_,
		_w5702_
	);
	LUT3 #(
		.INIT('h0d)
	) name5637 (
		_w5525_,
		_w5668_,
		_w5669_,
		_w5703_
	);
	LUT3 #(
		.INIT('h0d)
	) name5638 (
		_w5658_,
		_w5659_,
		_w5660_,
		_w5704_
	);
	LUT3 #(
		.INIT('h96)
	) name5639 (
		_w5702_,
		_w5703_,
		_w5704_,
		_w5705_
	);
	LUT3 #(
		.INIT('h0d)
	) name5640 (
		_w5475_,
		_w5647_,
		_w5648_,
		_w5706_
	);
	LUT3 #(
		.INIT('h0d)
	) name5641 (
		_w5643_,
		_w5644_,
		_w5645_,
		_w5707_
	);
	LUT4 #(
		.INIT('h153f)
	) name5642 (
		\a[12] ,
		\a[13] ,
		\a[61] ,
		\a[62] ,
		_w5708_
	);
	LUT4 #(
		.INIT('h000d)
	) name5643 (
		_w5537_,
		_w5538_,
		_w5539_,
		_w5632_,
		_w5709_
	);
	LUT4 #(
		.INIT('h6669)
	) name5644 (
		_w5706_,
		_w5707_,
		_w5708_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h4)
	) name5645 (
		_w5705_,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h2)
	) name5646 (
		_w5705_,
		_w5710_,
		_w5712_
	);
	LUT2 #(
		.INIT('h9)
	) name5647 (
		_w5705_,
		_w5710_,
		_w5713_
	);
	LUT4 #(
		.INIT('h6996)
	) name5648 (
		_w5699_,
		_w5700_,
		_w5701_,
		_w5713_,
		_w5714_
	);
	LUT3 #(
		.INIT('hd4)
	) name5649 (
		_w5590_,
		_w5591_,
		_w5592_,
		_w5715_
	);
	LUT3 #(
		.INIT('h32)
	) name5650 (
		_w5635_,
		_w5636_,
		_w5637_,
		_w5716_
	);
	LUT3 #(
		.INIT('h0d)
	) name5651 (
		_w5653_,
		_w5654_,
		_w5655_,
		_w5717_
	);
	LUT3 #(
		.INIT('h0d)
	) name5652 (
		_w5605_,
		_w5606_,
		_w5607_,
		_w5718_
	);
	LUT3 #(
		.INIT('h69)
	) name5653 (
		_w5716_,
		_w5717_,
		_w5718_,
		_w5719_
	);
	LUT3 #(
		.INIT('h32)
	) name5654 (
		_w5665_,
		_w5666_,
		_w5671_,
		_w5720_
	);
	LUT3 #(
		.INIT('h32)
	) name5655 (
		_w5650_,
		_w5651_,
		_w5657_,
		_w5721_
	);
	LUT3 #(
		.INIT('h69)
	) name5656 (
		_w5719_,
		_w5720_,
		_w5721_,
		_w5722_
	);
	LUT3 #(
		.INIT('h8e)
	) name5657 (
		_w5586_,
		_w5588_,
		_w5589_,
		_w5723_
	);
	LUT2 #(
		.INIT('h8)
	) name5658 (
		\a[14] ,
		\a[61] ,
		_w5724_
	);
	LUT4 #(
		.INIT('h153f)
	) name5659 (
		\a[15] ,
		\a[16] ,
		\a[59] ,
		\a[60] ,
		_w5725_
	);
	LUT4 #(
		.INIT('h8000)
	) name5660 (
		\a[15] ,
		\a[16] ,
		\a[59] ,
		\a[60] ,
		_w5726_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5661 (
		\a[15] ,
		\a[16] ,
		\a[59] ,
		\a[60] ,
		_w5727_
	);
	LUT2 #(
		.INIT('h8)
	) name5662 (
		\a[17] ,
		\a[58] ,
		_w5728_
	);
	LUT4 #(
		.INIT('h153f)
	) name5663 (
		\a[18] ,
		\a[26] ,
		\a[49] ,
		\a[57] ,
		_w5729_
	);
	LUT4 #(
		.INIT('h8000)
	) name5664 (
		\a[18] ,
		\a[26] ,
		\a[49] ,
		\a[57] ,
		_w5730_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5665 (
		\a[18] ,
		\a[26] ,
		\a[49] ,
		\a[57] ,
		_w5731_
	);
	LUT4 #(
		.INIT('h0660)
	) name5666 (
		_w5724_,
		_w5727_,
		_w5728_,
		_w5731_,
		_w5732_
	);
	LUT4 #(
		.INIT('h9009)
	) name5667 (
		_w5724_,
		_w5727_,
		_w5728_,
		_w5731_,
		_w5733_
	);
	LUT4 #(
		.INIT('h6996)
	) name5668 (
		_w5724_,
		_w5727_,
		_w5728_,
		_w5731_,
		_w5734_
	);
	LUT2 #(
		.INIT('h8)
	) name5669 (
		\a[27] ,
		\a[48] ,
		_w5735_
	);
	LUT4 #(
		.INIT('h153f)
	) name5670 (
		\a[28] ,
		\a[29] ,
		\a[46] ,
		\a[47] ,
		_w5736_
	);
	LUT4 #(
		.INIT('h8000)
	) name5671 (
		\a[28] ,
		\a[29] ,
		\a[46] ,
		\a[47] ,
		_w5737_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5672 (
		\a[28] ,
		\a[29] ,
		\a[46] ,
		\a[47] ,
		_w5738_
	);
	LUT2 #(
		.INIT('h6)
	) name5673 (
		_w5735_,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h1)
	) name5674 (
		_w5734_,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name5675 (
		_w5734_,
		_w5739_,
		_w5741_
	);
	LUT2 #(
		.INIT('h6)
	) name5676 (
		_w5734_,
		_w5739_,
		_w5742_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		\a[30] ,
		\a[45] ,
		_w5743_
	);
	LUT4 #(
		.INIT('h153f)
	) name5678 (
		\a[12] ,
		\a[19] ,
		\a[56] ,
		\a[63] ,
		_w5744_
	);
	LUT2 #(
		.INIT('h8)
	) name5679 (
		\a[19] ,
		\a[63] ,
		_w5745_
	);
	LUT4 #(
		.INIT('h8000)
	) name5680 (
		\a[12] ,
		\a[19] ,
		\a[56] ,
		\a[63] ,
		_w5746_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5681 (
		\a[12] ,
		\a[19] ,
		\a[56] ,
		\a[63] ,
		_w5747_
	);
	LUT2 #(
		.INIT('h8)
	) name5682 (
		\a[23] ,
		\a[52] ,
		_w5748_
	);
	LUT4 #(
		.INIT('h153f)
	) name5683 (
		\a[35] ,
		\a[36] ,
		\a[39] ,
		\a[40] ,
		_w5749_
	);
	LUT4 #(
		.INIT('h8000)
	) name5684 (
		\a[35] ,
		\a[36] ,
		\a[39] ,
		\a[40] ,
		_w5750_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5685 (
		\a[35] ,
		\a[36] ,
		\a[39] ,
		\a[40] ,
		_w5751_
	);
	LUT4 #(
		.INIT('h0660)
	) name5686 (
		_w5743_,
		_w5747_,
		_w5748_,
		_w5751_,
		_w5752_
	);
	LUT4 #(
		.INIT('h9009)
	) name5687 (
		_w5743_,
		_w5747_,
		_w5748_,
		_w5751_,
		_w5753_
	);
	LUT4 #(
		.INIT('h6996)
	) name5688 (
		_w5743_,
		_w5747_,
		_w5748_,
		_w5751_,
		_w5754_
	);
	LUT4 #(
		.INIT('h9a30)
	) name5689 (
		\a[13] ,
		\a[37] ,
		\a[38] ,
		\a[62] ,
		_w5755_
	);
	LUT2 #(
		.INIT('h6)
	) name5690 (
		_w5754_,
		_w5755_,
		_w5756_
	);
	LUT3 #(
		.INIT('h69)
	) name5691 (
		_w5723_,
		_w5742_,
		_w5756_,
		_w5757_
	);
	LUT4 #(
		.INIT('h4114)
	) name5692 (
		_w5722_,
		_w5723_,
		_w5742_,
		_w5756_,
		_w5758_
	);
	LUT4 #(
		.INIT('h8228)
	) name5693 (
		_w5722_,
		_w5723_,
		_w5742_,
		_w5756_,
		_w5759_
	);
	LUT3 #(
		.INIT('h69)
	) name5694 (
		_w5715_,
		_w5722_,
		_w5757_,
		_w5760_
	);
	LUT4 #(
		.INIT('h1e00)
	) name5695 (
		_w5594_,
		_w5597_,
		_w5714_,
		_w5760_,
		_w5761_
	);
	LUT4 #(
		.INIT('h4114)
	) name5696 (
		_w5714_,
		_w5715_,
		_w5722_,
		_w5757_,
		_w5762_
	);
	LUT4 #(
		.INIT('h8228)
	) name5697 (
		_w5714_,
		_w5715_,
		_w5722_,
		_w5757_,
		_w5763_
	);
	LUT4 #(
		.INIT('h01ef)
	) name5698 (
		_w5594_,
		_w5597_,
		_w5762_,
		_w5763_,
		_w5764_
	);
	LUT2 #(
		.INIT('h4)
	) name5699 (
		_w5761_,
		_w5764_,
		_w5765_
	);
	LUT3 #(
		.INIT('h2b)
	) name5700 (
		_w5599_,
		_w5601_,
		_w5615_,
		_w5766_
	);
	LUT2 #(
		.INIT('h8)
	) name5701 (
		\a[34] ,
		\a[41] ,
		_w5767_
	);
	LUT4 #(
		.INIT('h153f)
	) name5702 (
		\a[20] ,
		\a[25] ,
		\a[50] ,
		\a[55] ,
		_w5768_
	);
	LUT4 #(
		.INIT('h8000)
	) name5703 (
		\a[20] ,
		\a[25] ,
		\a[50] ,
		\a[55] ,
		_w5769_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5704 (
		\a[20] ,
		\a[25] ,
		\a[50] ,
		\a[55] ,
		_w5770_
	);
	LUT2 #(
		.INIT('h8)
	) name5705 (
		\a[31] ,
		\a[44] ,
		_w5771_
	);
	LUT4 #(
		.INIT('h153f)
	) name5706 (
		\a[32] ,
		\a[33] ,
		\a[42] ,
		\a[43] ,
		_w5772_
	);
	LUT2 #(
		.INIT('h8)
	) name5707 (
		\a[33] ,
		\a[43] ,
		_w5773_
	);
	LUT4 #(
		.INIT('h8000)
	) name5708 (
		\a[32] ,
		\a[33] ,
		\a[42] ,
		\a[43] ,
		_w5774_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5709 (
		\a[32] ,
		\a[33] ,
		\a[42] ,
		\a[43] ,
		_w5775_
	);
	LUT4 #(
		.INIT('h0660)
	) name5710 (
		_w5767_,
		_w5770_,
		_w5771_,
		_w5775_,
		_w5776_
	);
	LUT4 #(
		.INIT('h9009)
	) name5711 (
		_w5767_,
		_w5770_,
		_w5771_,
		_w5775_,
		_w5777_
	);
	LUT4 #(
		.INIT('h6996)
	) name5712 (
		_w5767_,
		_w5770_,
		_w5771_,
		_w5775_,
		_w5778_
	);
	LUT2 #(
		.INIT('h8)
	) name5713 (
		\a[21] ,
		\a[54] ,
		_w5779_
	);
	LUT4 #(
		.INIT('h153f)
	) name5714 (
		\a[22] ,
		\a[24] ,
		\a[51] ,
		\a[53] ,
		_w5780_
	);
	LUT4 #(
		.INIT('h8000)
	) name5715 (
		\a[22] ,
		\a[24] ,
		\a[51] ,
		\a[53] ,
		_w5781_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5716 (
		\a[22] ,
		\a[24] ,
		\a[51] ,
		\a[53] ,
		_w5782_
	);
	LUT2 #(
		.INIT('h6)
	) name5717 (
		_w5779_,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h9)
	) name5718 (
		_w5778_,
		_w5783_,
		_w5784_
	);
	LUT4 #(
		.INIT('h8e00)
	) name5719 (
		_w5621_,
		_w5625_,
		_w5626_,
		_w5784_,
		_w5785_
	);
	LUT3 #(
		.INIT('hb2)
	) name5720 (
		_w5602_,
		_w5610_,
		_w5614_,
		_w5786_
	);
	LUT4 #(
		.INIT('h0071)
	) name5721 (
		_w5621_,
		_w5625_,
		_w5626_,
		_w5784_,
		_w5787_
	);
	LUT3 #(
		.INIT('hc9)
	) name5722 (
		_w5785_,
		_w5786_,
		_w5787_,
		_w5788_
	);
	LUT2 #(
		.INIT('h4)
	) name5723 (
		_w5766_,
		_w5788_,
		_w5789_
	);
	LUT4 #(
		.INIT('he00e)
	) name5724 (
		_w5628_,
		_w5676_,
		_w5766_,
		_w5788_,
		_w5790_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5725 (
		_w5628_,
		_w5676_,
		_w5766_,
		_w5788_,
		_w5791_
	);
	LUT4 #(
		.INIT('he000)
	) name5726 (
		_w5484_,
		_w5486_,
		_w5616_,
		_w5791_,
		_w5792_
	);
	LUT4 #(
		.INIT('h8c00)
	) name5727 (
		_w5486_,
		_w5679_,
		_w5680_,
		_w5791_,
		_w5793_
	);
	LUT3 #(
		.INIT('h1e)
	) name5728 (
		_w5617_,
		_w5681_,
		_w5791_,
		_w5794_
	);
	LUT2 #(
		.INIT('h9)
	) name5729 (
		_w5765_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h1)
	) name5730 (
		_w5694_,
		_w5795_,
		_w5796_
	);
	LUT2 #(
		.INIT('h6)
	) name5731 (
		_w5694_,
		_w5795_,
		_w5797_
	);
	LUT2 #(
		.INIT('h4)
	) name5732 (
		_w5687_,
		_w5797_,
		_w5798_
	);
	LUT4 #(
		.INIT('hef00)
	) name5733 (
		_w5580_,
		_w5582_,
		_w5693_,
		_w5798_,
		_w5799_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name5734 (
		_w5580_,
		_w5582_,
		_w5687_,
		_w5693_,
		_w5800_
	);
	LUT3 #(
		.INIT('hcd)
	) name5735 (
		_w5797_,
		_w5799_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h1)
	) name5736 (
		_w5687_,
		_w5796_,
		_w5802_
	);
	LUT4 #(
		.INIT('hef00)
	) name5737 (
		_w5580_,
		_w5582_,
		_w5693_,
		_w5802_,
		_w5803_
	);
	LUT4 #(
		.INIT('h000b)
	) name5738 (
		_w5761_,
		_w5764_,
		_w5792_,
		_w5793_,
		_w5804_
	);
	LUT4 #(
		.INIT('h0073)
	) name5739 (
		_w5486_,
		_w5679_,
		_w5680_,
		_w5791_,
		_w5805_
	);
	LUT2 #(
		.INIT('h4)
	) name5740 (
		_w5617_,
		_w5805_,
		_w5806_
	);
	LUT4 #(
		.INIT('hd400)
	) name5741 (
		_w5590_,
		_w5591_,
		_w5592_,
		_w5722_,
		_w5807_
	);
	LUT4 #(
		.INIT('h0027)
	) name5742 (
		_w5715_,
		_w5758_,
		_w5759_,
		_w5807_,
		_w5808_
	);
	LUT4 #(
		.INIT('h8ee8)
	) name5743 (
		_w5699_,
		_w5700_,
		_w5701_,
		_w5713_,
		_w5809_
	);
	LUT2 #(
		.INIT('h8)
	) name5744 (
		\a[13] ,
		\a[63] ,
		_w5810_
	);
	LUT4 #(
		.INIT('h153f)
	) name5745 (
		\a[31] ,
		\a[32] ,
		\a[44] ,
		\a[45] ,
		_w5811_
	);
	LUT4 #(
		.INIT('h8000)
	) name5746 (
		\a[31] ,
		\a[32] ,
		\a[44] ,
		\a[45] ,
		_w5812_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5747 (
		\a[31] ,
		\a[32] ,
		\a[44] ,
		\a[45] ,
		_w5813_
	);
	LUT4 #(
		.INIT('h153f)
	) name5748 (
		\a[19] ,
		\a[23] ,
		\a[53] ,
		\a[57] ,
		_w5814_
	);
	LUT4 #(
		.INIT('h8000)
	) name5749 (
		\a[19] ,
		\a[23] ,
		\a[53] ,
		\a[57] ,
		_w5815_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5750 (
		\a[19] ,
		\a[23] ,
		\a[53] ,
		\a[57] ,
		_w5816_
	);
	LUT4 #(
		.INIT('h1428)
	) name5751 (
		_w5773_,
		_w5810_,
		_w5813_,
		_w5816_,
		_w5817_
	);
	LUT4 #(
		.INIT('h8241)
	) name5752 (
		_w5773_,
		_w5810_,
		_w5813_,
		_w5816_,
		_w5818_
	);
	LUT4 #(
		.INIT('h6996)
	) name5753 (
		_w5773_,
		_w5810_,
		_w5813_,
		_w5816_,
		_w5819_
	);
	LUT4 #(
		.INIT('h153f)
	) name5754 (
		\a[21] ,
		\a[22] ,
		\a[54] ,
		\a[55] ,
		_w5820_
	);
	LUT4 #(
		.INIT('h8000)
	) name5755 (
		\a[21] ,
		\a[22] ,
		\a[54] ,
		\a[55] ,
		_w5821_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5756 (
		\a[21] ,
		\a[22] ,
		\a[54] ,
		\a[55] ,
		_w5822_
	);
	LUT2 #(
		.INIT('h6)
	) name5757 (
		_w4837_,
		_w5822_,
		_w5823_
	);
	LUT2 #(
		.INIT('h6)
	) name5758 (
		_w5819_,
		_w5823_,
		_w5824_
	);
	LUT4 #(
		.INIT('h002b)
	) name5759 (
		_w5719_,
		_w5720_,
		_w5721_,
		_w5824_,
		_w5825_
	);
	LUT3 #(
		.INIT('h0e)
	) name5760 (
		_w5701_,
		_w5711_,
		_w5712_,
		_w5826_
	);
	LUT4 #(
		.INIT('hd400)
	) name5761 (
		_w5719_,
		_w5720_,
		_w5721_,
		_w5824_,
		_w5827_
	);
	LUT4 #(
		.INIT('h00b2)
	) name5762 (
		_w5701_,
		_w5705_,
		_w5710_,
		_w5827_,
		_w5828_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name5763 (
		_w5719_,
		_w5720_,
		_w5721_,
		_w5824_,
		_w5829_
	);
	LUT4 #(
		.INIT('h004d)
	) name5764 (
		_w5701_,
		_w5705_,
		_w5710_,
		_w5829_,
		_w5830_
	);
	LUT3 #(
		.INIT('hc9)
	) name5765 (
		_w5825_,
		_w5826_,
		_w5827_,
		_w5831_
	);
	LUT4 #(
		.INIT('h008a)
	) name5766 (
		_w5809_,
		_w5825_,
		_w5828_,
		_w5830_,
		_w5832_
	);
	LUT4 #(
		.INIT('h5510)
	) name5767 (
		_w5809_,
		_w5825_,
		_w5828_,
		_w5830_,
		_w5833_
	);
	LUT4 #(
		.INIT('h5a69)
	) name5768 (
		_w5809_,
		_w5825_,
		_w5826_,
		_w5827_,
		_w5834_
	);
	LUT2 #(
		.INIT('h4)
	) name5769 (
		_w5808_,
		_w5834_,
		_w5835_
	);
	LUT2 #(
		.INIT('h9)
	) name5770 (
		_w5808_,
		_w5834_,
		_w5836_
	);
	LUT3 #(
		.INIT('h82)
	) name5771 (
		_w5714_,
		_w5808_,
		_w5834_,
		_w5837_
	);
	LUT4 #(
		.INIT('h2882)
	) name5772 (
		_w5714_,
		_w5715_,
		_w5722_,
		_w5757_,
		_w5838_
	);
	LUT3 #(
		.INIT('h90)
	) name5773 (
		_w5808_,
		_w5834_,
		_w5838_,
		_w5839_
	);
	LUT3 #(
		.INIT('h82)
	) name5774 (
		_w5760_,
		_w5808_,
		_w5834_,
		_w5840_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name5775 (
		_w5695_,
		_w5837_,
		_w5839_,
		_w5840_,
		_w5841_
	);
	LUT3 #(
		.INIT('h0b)
	) name5776 (
		_w5695_,
		_w5714_,
		_w5836_,
		_w5842_
	);
	LUT3 #(
		.INIT('h8c)
	) name5777 (
		_w5761_,
		_w5841_,
		_w5842_,
		_w5843_
	);
	LUT4 #(
		.INIT('h10f1)
	) name5778 (
		_w5628_,
		_w5676_,
		_w5766_,
		_w5788_,
		_w5844_
	);
	LUT4 #(
		.INIT('h8e00)
	) name5779 (
		_w5586_,
		_w5588_,
		_w5589_,
		_w5756_,
		_w5845_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name5780 (
		_w5734_,
		_w5739_,
		_w5754_,
		_w5755_,
		_w5846_
	);
	LUT4 #(
		.INIT('h008e)
	) name5781 (
		_w5586_,
		_w5588_,
		_w5589_,
		_w5740_,
		_w5847_
	);
	LUT4 #(
		.INIT('hdddc)
	) name5782 (
		_w5741_,
		_w5845_,
		_w5846_,
		_w5847_,
		_w5848_
	);
	LUT4 #(
		.INIT('h1117)
	) name5783 (
		_w5706_,
		_w5707_,
		_w5708_,
		_w5709_,
		_w5849_
	);
	LUT3 #(
		.INIT('h2b)
	) name5784 (
		_w5716_,
		_w5717_,
		_w5718_,
		_w5850_
	);
	LUT3 #(
		.INIT('h17)
	) name5785 (
		_w5702_,
		_w5703_,
		_w5704_,
		_w5851_
	);
	LUT3 #(
		.INIT('h96)
	) name5786 (
		_w5849_,
		_w5850_,
		_w5851_,
		_w5852_
	);
	LUT3 #(
		.INIT('h32)
	) name5787 (
		_w5767_,
		_w5768_,
		_w5769_,
		_w5853_
	);
	LUT3 #(
		.INIT('h0d)
	) name5788 (
		_w5735_,
		_w5736_,
		_w5737_,
		_w5854_
	);
	LUT3 #(
		.INIT('h0d)
	) name5789 (
		_w5743_,
		_w5744_,
		_w5746_,
		_w5855_
	);
	LUT3 #(
		.INIT('h69)
	) name5790 (
		_w5853_,
		_w5854_,
		_w5855_,
		_w5856_
	);
	LUT3 #(
		.INIT('h13)
	) name5791 (
		\a[13] ,
		\a[37] ,
		\a[62] ,
		_w5857_
	);
	LUT4 #(
		.INIT('he0c0)
	) name5792 (
		\a[13] ,
		\a[37] ,
		\a[38] ,
		\a[62] ,
		_w5858_
	);
	LUT2 #(
		.INIT('h8)
	) name5793 (
		\a[14] ,
		\a[62] ,
		_w5859_
	);
	LUT2 #(
		.INIT('h1)
	) name5794 (
		_w5858_,
		_w5859_,
		_w5860_
	);
	LUT3 #(
		.INIT('h80)
	) name5795 (
		\a[14] ,
		\a[38] ,
		\a[62] ,
		_w5861_
	);
	LUT2 #(
		.INIT('h4)
	) name5796 (
		_w5857_,
		_w5861_,
		_w5862_
	);
	LUT3 #(
		.INIT('hd2)
	) name5797 (
		\a[38] ,
		_w5857_,
		_w5859_,
		_w5863_
	);
	LUT3 #(
		.INIT('h0d)
	) name5798 (
		_w5748_,
		_w5749_,
		_w5750_,
		_w5864_
	);
	LUT2 #(
		.INIT('h6)
	) name5799 (
		_w5863_,
		_w5864_,
		_w5865_
	);
	LUT3 #(
		.INIT('h45)
	) name5800 (
		_w5776_,
		_w5777_,
		_w5783_,
		_w5866_
	);
	LUT3 #(
		.INIT('h69)
	) name5801 (
		_w5856_,
		_w5865_,
		_w5866_,
		_w5867_
	);
	LUT3 #(
		.INIT('h96)
	) name5802 (
		_w5848_,
		_w5852_,
		_w5867_,
		_w5868_
	);
	LUT3 #(
		.INIT('h0b)
	) name5803 (
		_w5766_,
		_w5788_,
		_w5868_,
		_w5869_
	);
	LUT3 #(
		.INIT('hb2)
	) name5804 (
		_w5696_,
		_w5697_,
		_w5698_,
		_w5870_
	);
	LUT2 #(
		.INIT('h8)
	) name5805 (
		\a[28] ,
		\a[48] ,
		_w5871_
	);
	LUT4 #(
		.INIT('h153f)
	) name5806 (
		\a[29] ,
		\a[30] ,
		\a[46] ,
		\a[47] ,
		_w5872_
	);
	LUT2 #(
		.INIT('h8)
	) name5807 (
		\a[30] ,
		\a[47] ,
		_w5873_
	);
	LUT4 #(
		.INIT('h8000)
	) name5808 (
		\a[29] ,
		\a[30] ,
		\a[46] ,
		\a[47] ,
		_w5874_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5809 (
		\a[29] ,
		\a[30] ,
		\a[46] ,
		\a[47] ,
		_w5875_
	);
	LUT2 #(
		.INIT('h8)
	) name5810 (
		\a[34] ,
		\a[42] ,
		_w5876_
	);
	LUT4 #(
		.INIT('h153f)
	) name5811 (
		\a[35] ,
		\a[36] ,
		\a[40] ,
		\a[41] ,
		_w5877_
	);
	LUT4 #(
		.INIT('h8000)
	) name5812 (
		\a[35] ,
		\a[36] ,
		\a[40] ,
		\a[41] ,
		_w5878_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5813 (
		\a[35] ,
		\a[36] ,
		\a[40] ,
		\a[41] ,
		_w5879_
	);
	LUT4 #(
		.INIT('h0660)
	) name5814 (
		_w5871_,
		_w5875_,
		_w5876_,
		_w5879_,
		_w5880_
	);
	LUT4 #(
		.INIT('h9009)
	) name5815 (
		_w5871_,
		_w5875_,
		_w5876_,
		_w5879_,
		_w5881_
	);
	LUT4 #(
		.INIT('h6996)
	) name5816 (
		_w5871_,
		_w5875_,
		_w5876_,
		_w5879_,
		_w5882_
	);
	LUT2 #(
		.INIT('h8)
	) name5817 (
		\a[37] ,
		\a[39] ,
		_w5883_
	);
	LUT4 #(
		.INIT('h153f)
	) name5818 (
		\a[24] ,
		\a[25] ,
		\a[51] ,
		\a[52] ,
		_w5884_
	);
	LUT2 #(
		.INIT('h8)
	) name5819 (
		\a[25] ,
		\a[52] ,
		_w5885_
	);
	LUT4 #(
		.INIT('h8000)
	) name5820 (
		\a[24] ,
		\a[25] ,
		\a[51] ,
		\a[52] ,
		_w5886_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5821 (
		\a[24] ,
		\a[25] ,
		\a[51] ,
		\a[52] ,
		_w5887_
	);
	LUT2 #(
		.INIT('h6)
	) name5822 (
		_w5883_,
		_w5887_,
		_w5888_
	);
	LUT2 #(
		.INIT('h6)
	) name5823 (
		_w5882_,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h8)
	) name5824 (
		\a[15] ,
		\a[61] ,
		_w5890_
	);
	LUT4 #(
		.INIT('h153f)
	) name5825 (
		\a[16] ,
		\a[17] ,
		\a[59] ,
		\a[60] ,
		_w5891_
	);
	LUT4 #(
		.INIT('h8000)
	) name5826 (
		\a[16] ,
		\a[17] ,
		\a[59] ,
		\a[60] ,
		_w5892_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5827 (
		\a[16] ,
		\a[17] ,
		\a[59] ,
		\a[60] ,
		_w5893_
	);
	LUT2 #(
		.INIT('h6)
	) name5828 (
		_w5890_,
		_w5893_,
		_w5894_
	);
	LUT3 #(
		.INIT('h0d)
	) name5829 (
		_w5779_,
		_w5780_,
		_w5781_,
		_w5895_
	);
	LUT2 #(
		.INIT('h4)
	) name5830 (
		_w5894_,
		_w5895_,
		_w5896_
	);
	LUT2 #(
		.INIT('h8)
	) name5831 (
		\a[18] ,
		\a[58] ,
		_w5897_
	);
	LUT4 #(
		.INIT('h153f)
	) name5832 (
		\a[26] ,
		\a[27] ,
		\a[49] ,
		\a[50] ,
		_w5898_
	);
	LUT2 #(
		.INIT('h8)
	) name5833 (
		\a[27] ,
		\a[50] ,
		_w5899_
	);
	LUT4 #(
		.INIT('h8000)
	) name5834 (
		\a[26] ,
		\a[27] ,
		\a[49] ,
		\a[50] ,
		_w5900_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5835 (
		\a[26] ,
		\a[27] ,
		\a[49] ,
		\a[50] ,
		_w5901_
	);
	LUT2 #(
		.INIT('h6)
	) name5836 (
		_w5897_,
		_w5901_,
		_w5902_
	);
	LUT3 #(
		.INIT('h69)
	) name5837 (
		_w5894_,
		_w5895_,
		_w5902_,
		_w5903_
	);
	LUT3 #(
		.INIT('hf6)
	) name5838 (
		_w5870_,
		_w5889_,
		_w5903_,
		_w5904_
	);
	LUT4 #(
		.INIT('h0023)
	) name5839 (
		_w5611_,
		_w5612_,
		_w5614_,
		_w5787_,
		_w5905_
	);
	LUT3 #(
		.INIT('h0d)
	) name5840 (
		_w5728_,
		_w5729_,
		_w5730_,
		_w5906_
	);
	LUT3 #(
		.INIT('h0d)
	) name5841 (
		_w5724_,
		_w5725_,
		_w5726_,
		_w5907_
	);
	LUT3 #(
		.INIT('h0d)
	) name5842 (
		_w5771_,
		_w5772_,
		_w5774_,
		_w5908_
	);
	LUT3 #(
		.INIT('h96)
	) name5843 (
		_w5906_,
		_w5907_,
		_w5908_,
		_w5909_
	);
	LUT3 #(
		.INIT('h32)
	) name5844 (
		_w5732_,
		_w5733_,
		_w5739_,
		_w5910_
	);
	LUT3 #(
		.INIT('h32)
	) name5845 (
		_w5752_,
		_w5753_,
		_w5755_,
		_w5911_
	);
	LUT3 #(
		.INIT('h69)
	) name5846 (
		_w5909_,
		_w5910_,
		_w5911_,
		_w5912_
	);
	LUT3 #(
		.INIT('h9f)
	) name5847 (
		_w5870_,
		_w5889_,
		_w5903_,
		_w5913_
	);
	LUT4 #(
		.INIT('h1eff)
	) name5848 (
		_w5785_,
		_w5905_,
		_w5912_,
		_w5913_,
		_w5914_
	);
	LUT3 #(
		.INIT('h96)
	) name5849 (
		_w5870_,
		_w5889_,
		_w5903_,
		_w5915_
	);
	LUT4 #(
		.INIT('hffe1)
	) name5850 (
		_w5785_,
		_w5905_,
		_w5912_,
		_w5915_,
		_w5916_
	);
	LUT3 #(
		.INIT('hd0)
	) name5851 (
		_w5904_,
		_w5914_,
		_w5916_,
		_w5917_
	);
	LUT4 #(
		.INIT('h1e00)
	) name5852 (
		_w5789_,
		_w5790_,
		_w5868_,
		_w5917_,
		_w5918_
	);
	LUT3 #(
		.INIT('h04)
	) name5853 (
		_w5790_,
		_w5869_,
		_w5917_,
		_w5919_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5854 (
		_w5868_,
		_w5904_,
		_w5914_,
		_w5916_,
		_w5920_
	);
	LUT2 #(
		.INIT('h4)
	) name5855 (
		_w5844_,
		_w5920_,
		_w5921_
	);
	LUT3 #(
		.INIT('h01)
	) name5856 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5922_
	);
	LUT4 #(
		.INIT('h0110)
	) name5857 (
		_w5804_,
		_w5806_,
		_w5843_,
		_w5922_,
		_w5923_
	);
	LUT4 #(
		.INIT('he00e)
	) name5858 (
		_w5804_,
		_w5806_,
		_w5843_,
		_w5922_,
		_w5924_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5859 (
		_w5804_,
		_w5806_,
		_w5843_,
		_w5922_,
		_w5925_
	);
	LUT3 #(
		.INIT('h87)
	) name5860 (
		_w5694_,
		_w5795_,
		_w5925_,
		_w5926_
	);
	LUT3 #(
		.INIT('hf0)
	) name5861 (
		_w5694_,
		_w5795_,
		_w5925_,
		_w5927_
	);
	LUT3 #(
		.INIT('he4)
	) name5862 (
		_w5803_,
		_w5926_,
		_w5927_,
		_w5928_
	);
	LUT3 #(
		.INIT('h01)
	) name5863 (
		_w5687_,
		_w5796_,
		_w5923_,
		_w5929_
	);
	LUT4 #(
		.INIT('hef00)
	) name5864 (
		_w5580_,
		_w5582_,
		_w5693_,
		_w5929_,
		_w5930_
	);
	LUT3 #(
		.INIT('h08)
	) name5865 (
		_w5694_,
		_w5795_,
		_w5923_,
		_w5931_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5866 (
		_w5841_,
		_w5918_,
		_w5919_,
		_w5921_,
		_w5932_
	);
	LUT3 #(
		.INIT('h40)
	) name5867 (
		_w5761_,
		_w5841_,
		_w5842_,
		_w5933_
	);
	LUT4 #(
		.INIT('h011f)
	) name5868 (
		_w5789_,
		_w5790_,
		_w5868_,
		_w5917_,
		_w5934_
	);
	LUT4 #(
		.INIT('hf111)
	) name5869 (
		_w5785_,
		_w5905_,
		_w5912_,
		_w5913_,
		_w5935_
	);
	LUT4 #(
		.INIT('hff96)
	) name5870 (
		_w5870_,
		_w5889_,
		_w5903_,
		_w5912_,
		_w5936_
	);
	LUT4 #(
		.INIT('hcd00)
	) name5871 (
		_w5785_,
		_w5904_,
		_w5905_,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h8)
	) name5872 (
		\a[34] ,
		\a[43] ,
		_w5938_
	);
	LUT4 #(
		.INIT('h153f)
	) name5873 (
		\a[22] ,
		\a[26] ,
		\a[51] ,
		\a[55] ,
		_w5939_
	);
	LUT4 #(
		.INIT('h8000)
	) name5874 (
		\a[22] ,
		\a[26] ,
		\a[51] ,
		\a[55] ,
		_w5940_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5875 (
		\a[22] ,
		\a[26] ,
		\a[51] ,
		\a[55] ,
		_w5941_
	);
	LUT4 #(
		.INIT('h153f)
	) name5876 (
		\a[23] ,
		\a[24] ,
		\a[53] ,
		\a[54] ,
		_w5942_
	);
	LUT4 #(
		.INIT('h8000)
	) name5877 (
		\a[23] ,
		\a[24] ,
		\a[53] ,
		\a[54] ,
		_w5943_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5878 (
		\a[23] ,
		\a[24] ,
		\a[53] ,
		\a[54] ,
		_w5944_
	);
	LUT4 #(
		.INIT('h1428)
	) name5879 (
		_w5885_,
		_w5938_,
		_w5941_,
		_w5944_,
		_w5945_
	);
	LUT4 #(
		.INIT('h8241)
	) name5880 (
		_w5885_,
		_w5938_,
		_w5941_,
		_w5944_,
		_w5946_
	);
	LUT4 #(
		.INIT('h6996)
	) name5881 (
		_w5885_,
		_w5938_,
		_w5941_,
		_w5944_,
		_w5947_
	);
	LUT2 #(
		.INIT('h8)
	) name5882 (
		\a[16] ,
		\a[61] ,
		_w5948_
	);
	LUT4 #(
		.INIT('h153f)
	) name5883 (
		\a[32] ,
		\a[33] ,
		\a[44] ,
		\a[45] ,
		_w5949_
	);
	LUT4 #(
		.INIT('h8000)
	) name5884 (
		\a[32] ,
		\a[33] ,
		\a[44] ,
		\a[45] ,
		_w5950_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5885 (
		\a[32] ,
		\a[33] ,
		\a[44] ,
		\a[45] ,
		_w5951_
	);
	LUT2 #(
		.INIT('h6)
	) name5886 (
		_w5948_,
		_w5951_,
		_w5952_
	);
	LUT2 #(
		.INIT('h9)
	) name5887 (
		_w5947_,
		_w5952_,
		_w5953_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5888 (
		_w5909_,
		_w5910_,
		_w5911_,
		_w5953_,
		_w5954_
	);
	LUT3 #(
		.INIT('h17)
	) name5889 (
		_w5856_,
		_w5865_,
		_w5866_,
		_w5955_
	);
	LUT4 #(
		.INIT('h00d4)
	) name5890 (
		_w5909_,
		_w5910_,
		_w5911_,
		_w5953_,
		_w5956_
	);
	LUT3 #(
		.INIT('hc9)
	) name5891 (
		_w5954_,
		_w5955_,
		_w5956_,
		_w5957_
	);
	LUT4 #(
		.INIT('he800)
	) name5892 (
		_w5848_,
		_w5852_,
		_w5867_,
		_w5957_,
		_w5958_
	);
	LUT4 #(
		.INIT('h0017)
	) name5893 (
		_w5848_,
		_w5852_,
		_w5867_,
		_w5957_,
		_w5959_
	);
	LUT4 #(
		.INIT('h17e8)
	) name5894 (
		_w5848_,
		_w5852_,
		_w5867_,
		_w5957_,
		_w5960_
	);
	LUT3 #(
		.INIT('h78)
	) name5895 (
		_w5935_,
		_w5937_,
		_w5960_,
		_w5961_
	);
	LUT3 #(
		.INIT('h17)
	) name5896 (
		_w5906_,
		_w5907_,
		_w5908_,
		_w5962_
	);
	LUT2 #(
		.INIT('h8)
	) name5897 (
		\a[18] ,
		\a[60] ,
		_w5963_
	);
	LUT4 #(
		.INIT('h8000)
	) name5898 (
		\a[17] ,
		\a[18] ,
		\a[59] ,
		\a[60] ,
		_w5964_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5899 (
		\a[17] ,
		\a[18] ,
		\a[59] ,
		\a[60] ,
		_w5965_
	);
	LUT4 #(
		.INIT('hf20d)
	) name5900 (
		_w5883_,
		_w5884_,
		_w5886_,
		_w5965_,
		_w5966_
	);
	LUT4 #(
		.INIT('he800)
	) name5901 (
		_w5906_,
		_w5907_,
		_w5908_,
		_w5966_,
		_w5967_
	);
	LUT4 #(
		.INIT('h0017)
	) name5902 (
		_w5906_,
		_w5907_,
		_w5908_,
		_w5966_,
		_w5968_
	);
	LUT4 #(
		.INIT('h17e8)
	) name5903 (
		_w5906_,
		_w5907_,
		_w5908_,
		_w5966_,
		_w5969_
	);
	LUT3 #(
		.INIT('h2b)
	) name5904 (
		_w5853_,
		_w5854_,
		_w5855_,
		_w5970_
	);
	LUT2 #(
		.INIT('h6)
	) name5905 (
		_w5969_,
		_w5970_,
		_w5971_
	);
	LUT3 #(
		.INIT('h17)
	) name5906 (
		_w5870_,
		_w5889_,
		_w5903_,
		_w5972_
	);
	LUT4 #(
		.INIT('he800)
	) name5907 (
		_w5870_,
		_w5889_,
		_w5903_,
		_w5971_,
		_w5973_
	);
	LUT4 #(
		.INIT('h0017)
	) name5908 (
		_w5870_,
		_w5889_,
		_w5903_,
		_w5971_,
		_w5974_
	);
	LUT3 #(
		.INIT('h0d)
	) name5909 (
		_w4837_,
		_w5820_,
		_w5821_,
		_w5975_
	);
	LUT3 #(
		.INIT('h0d)
	) name5910 (
		_w5871_,
		_w5872_,
		_w5874_,
		_w5976_
	);
	LUT3 #(
		.INIT('h0d)
	) name5911 (
		_w5810_,
		_w5811_,
		_w5812_,
		_w5977_
	);
	LUT3 #(
		.INIT('h96)
	) name5912 (
		_w5975_,
		_w5976_,
		_w5977_,
		_w5978_
	);
	LUT3 #(
		.INIT('h0d)
	) name5913 (
		_w5890_,
		_w5891_,
		_w5892_,
		_w5979_
	);
	LUT3 #(
		.INIT('h0d)
	) name5914 (
		_w5897_,
		_w5898_,
		_w5900_,
		_w5980_
	);
	LUT3 #(
		.INIT('h32)
	) name5915 (
		_w5773_,
		_w5814_,
		_w5815_,
		_w5981_
	);
	LUT3 #(
		.INIT('h96)
	) name5916 (
		_w5979_,
		_w5980_,
		_w5981_,
		_w5982_
	);
	LUT3 #(
		.INIT('h32)
	) name5917 (
		_w5817_,
		_w5818_,
		_w5823_,
		_w5983_
	);
	LUT3 #(
		.INIT('h69)
	) name5918 (
		_w5978_,
		_w5982_,
		_w5983_,
		_w5984_
	);
	LUT4 #(
		.INIT('hf299)
	) name5919 (
		_w5971_,
		_w5972_,
		_w5974_,
		_w5984_,
		_w5985_
	);
	LUT4 #(
		.INIT('hd400)
	) name5920 (
		_w5808_,
		_w5809_,
		_w5831_,
		_w5985_,
		_w5986_
	);
	LUT4 #(
		.INIT('h0032)
	) name5921 (
		_w5808_,
		_w5832_,
		_w5833_,
		_w5985_,
		_w5987_
	);
	LUT3 #(
		.INIT('he8)
	) name5922 (
		_w5849_,
		_w5850_,
		_w5851_,
		_w5988_
	);
	LUT2 #(
		.INIT('h8)
	) name5923 (
		\a[35] ,
		\a[42] ,
		_w5989_
	);
	LUT4 #(
		.INIT('h153f)
	) name5924 (
		\a[36] ,
		\a[37] ,
		\a[40] ,
		\a[41] ,
		_w5990_
	);
	LUT2 #(
		.INIT('h8)
	) name5925 (
		\a[37] ,
		\a[41] ,
		_w5991_
	);
	LUT4 #(
		.INIT('h8000)
	) name5926 (
		\a[36] ,
		\a[37] ,
		\a[40] ,
		\a[41] ,
		_w5992_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5927 (
		\a[36] ,
		\a[37] ,
		\a[40] ,
		\a[41] ,
		_w5993_
	);
	LUT4 #(
		.INIT('h153f)
	) name5928 (
		\a[14] ,
		\a[31] ,
		\a[46] ,
		\a[63] ,
		_w5994_
	);
	LUT2 #(
		.INIT('h8)
	) name5929 (
		\a[31] ,
		\a[63] ,
		_w5995_
	);
	LUT4 #(
		.INIT('h8000)
	) name5930 (
		\a[14] ,
		\a[31] ,
		\a[46] ,
		\a[63] ,
		_w5996_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5931 (
		\a[14] ,
		\a[31] ,
		\a[46] ,
		\a[63] ,
		_w5997_
	);
	LUT4 #(
		.INIT('h1428)
	) name5932 (
		_w5873_,
		_w5989_,
		_w5993_,
		_w5997_,
		_w5998_
	);
	LUT4 #(
		.INIT('h8241)
	) name5933 (
		_w5873_,
		_w5989_,
		_w5993_,
		_w5997_,
		_w5999_
	);
	LUT4 #(
		.INIT('h6996)
	) name5934 (
		_w5873_,
		_w5989_,
		_w5993_,
		_w5997_,
		_w6000_
	);
	LUT4 #(
		.INIT('h9a30)
	) name5935 (
		\a[15] ,
		\a[38] ,
		\a[39] ,
		\a[62] ,
		_w6001_
	);
	LUT2 #(
		.INIT('h6)
	) name5936 (
		_w6000_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h8)
	) name5937 (
		\a[19] ,
		\a[58] ,
		_w6003_
	);
	LUT4 #(
		.INIT('h153f)
	) name5938 (
		\a[20] ,
		\a[21] ,
		\a[56] ,
		\a[57] ,
		_w6004_
	);
	LUT4 #(
		.INIT('h8000)
	) name5939 (
		\a[20] ,
		\a[21] ,
		\a[56] ,
		\a[57] ,
		_w6005_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5940 (
		\a[20] ,
		\a[21] ,
		\a[56] ,
		\a[57] ,
		_w6006_
	);
	LUT2 #(
		.INIT('h6)
	) name5941 (
		_w6003_,
		_w6006_,
		_w6007_
	);
	LUT3 #(
		.INIT('h0d)
	) name5942 (
		_w5876_,
		_w5877_,
		_w5878_,
		_w6008_
	);
	LUT4 #(
		.INIT('h153f)
	) name5943 (
		\a[28] ,
		\a[29] ,
		\a[48] ,
		\a[49] ,
		_w6009_
	);
	LUT4 #(
		.INIT('h8000)
	) name5944 (
		\a[28] ,
		\a[29] ,
		\a[48] ,
		\a[49] ,
		_w6010_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5945 (
		\a[28] ,
		\a[29] ,
		\a[48] ,
		\a[49] ,
		_w6011_
	);
	LUT2 #(
		.INIT('h6)
	) name5946 (
		_w5899_,
		_w6011_,
		_w6012_
	);
	LUT3 #(
		.INIT('h69)
	) name5947 (
		_w6007_,
		_w6008_,
		_w6012_,
		_w6013_
	);
	LUT3 #(
		.INIT('hf6)
	) name5948 (
		_w5988_,
		_w6002_,
		_w6013_,
		_w6014_
	);
	LUT4 #(
		.INIT('h004d)
	) name5949 (
		_w5701_,
		_w5705_,
		_w5710_,
		_w5827_,
		_w6015_
	);
	LUT3 #(
		.INIT('h9f)
	) name5950 (
		_w5988_,
		_w6002_,
		_w6013_,
		_w6016_
	);
	LUT3 #(
		.INIT('h45)
	) name5951 (
		_w5860_,
		_w5862_,
		_w5864_,
		_w6017_
	);
	LUT3 #(
		.INIT('h0d)
	) name5952 (
		_w5894_,
		_w5895_,
		_w5902_,
		_w6018_
	);
	LUT3 #(
		.INIT('hb2)
	) name5953 (
		_w5894_,
		_w5895_,
		_w5902_,
		_w6019_
	);
	LUT2 #(
		.INIT('h1)
	) name5954 (
		_w6017_,
		_w6019_,
		_w6020_
	);
	LUT3 #(
		.INIT('h04)
	) name5955 (
		_w5896_,
		_w6017_,
		_w6018_,
		_w6021_
	);
	LUT3 #(
		.INIT('h32)
	) name5956 (
		_w5880_,
		_w5881_,
		_w5888_,
		_w6022_
	);
	LUT3 #(
		.INIT('he1)
	) name5957 (
		_w6020_,
		_w6021_,
		_w6022_,
		_w6023_
	);
	LUT4 #(
		.INIT('h1fef)
	) name5958 (
		_w5825_,
		_w6015_,
		_w6016_,
		_w6023_,
		_w6024_
	);
	LUT3 #(
		.INIT('h96)
	) name5959 (
		_w5988_,
		_w6002_,
		_w6013_,
		_w6025_
	);
	LUT3 #(
		.INIT('h0e)
	) name5960 (
		_w5825_,
		_w6015_,
		_w6023_,
		_w6026_
	);
	LUT4 #(
		.INIT('hffe1)
	) name5961 (
		_w5825_,
		_w6015_,
		_w6023_,
		_w6025_,
		_w6027_
	);
	LUT3 #(
		.INIT('hd0)
	) name5962 (
		_w6014_,
		_w6024_,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h4)
	) name5963 (
		_w5987_,
		_w6028_,
		_w6029_
	);
	LUT3 #(
		.INIT('h10)
	) name5964 (
		_w5986_,
		_w5987_,
		_w6028_,
		_w6030_
	);
	LUT4 #(
		.INIT('hff1e)
	) name5965 (
		_w5832_,
		_w5835_,
		_w5985_,
		_w6028_,
		_w6031_
	);
	LUT4 #(
		.INIT('h9699)
	) name5966 (
		_w5934_,
		_w5961_,
		_w6030_,
		_w6031_,
		_w6032_
	);
	LUT3 #(
		.INIT('h10)
	) name5967 (
		_w5932_,
		_w5933_,
		_w6032_,
		_w6033_
	);
	LUT3 #(
		.INIT('h0e)
	) name5968 (
		_w5932_,
		_w5933_,
		_w6032_,
		_w6034_
	);
	LUT3 #(
		.INIT('he1)
	) name5969 (
		_w5932_,
		_w5933_,
		_w6032_,
		_w6035_
	);
	LUT4 #(
		.INIT('hfe01)
	) name5970 (
		_w5924_,
		_w5930_,
		_w5931_,
		_w6035_,
		_w6036_
	);
	LUT2 #(
		.INIT('h1)
	) name5971 (
		_w5924_,
		_w6034_,
		_w6037_
	);
	LUT2 #(
		.INIT('h4)
	) name5972 (
		_w5931_,
		_w6037_,
		_w6038_
	);
	LUT4 #(
		.INIT('hb2bb)
	) name5973 (
		_w5934_,
		_w5961_,
		_w6030_,
		_w6031_,
		_w6039_
	);
	LUT4 #(
		.INIT('hcd05)
	) name5974 (
		_w5825_,
		_w6014_,
		_w6015_,
		_w6016_,
		_w6040_
	);
	LUT3 #(
		.INIT('hf8)
	) name5975 (
		_w6014_,
		_w6016_,
		_w6023_,
		_w6041_
	);
	LUT3 #(
		.INIT('h40)
	) name5976 (
		_w6026_,
		_w6040_,
		_w6041_,
		_w6042_
	);
	LUT4 #(
		.INIT('h00fb)
	) name5977 (
		_w5896_,
		_w6017_,
		_w6018_,
		_w6022_,
		_w6043_
	);
	LUT4 #(
		.INIT('h153f)
	) name5978 (
		\a[19] ,
		\a[21] ,
		\a[57] ,
		\a[59] ,
		_w6044_
	);
	LUT4 #(
		.INIT('h8000)
	) name5979 (
		\a[19] ,
		\a[21] ,
		\a[57] ,
		\a[59] ,
		_w6045_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5980 (
		\a[19] ,
		\a[21] ,
		\a[57] ,
		\a[59] ,
		_w6046_
	);
	LUT2 #(
		.INIT('h8)
	) name5981 (
		\a[27] ,
		\a[51] ,
		_w6047_
	);
	LUT4 #(
		.INIT('h153f)
	) name5982 (
		\a[28] ,
		\a[29] ,
		\a[49] ,
		\a[50] ,
		_w6048_
	);
	LUT4 #(
		.INIT('h8000)
	) name5983 (
		\a[28] ,
		\a[29] ,
		\a[49] ,
		\a[50] ,
		_w6049_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5984 (
		\a[28] ,
		\a[29] ,
		\a[49] ,
		\a[50] ,
		_w6050_
	);
	LUT4 #(
		.INIT('h0660)
	) name5985 (
		_w5963_,
		_w6046_,
		_w6047_,
		_w6050_,
		_w6051_
	);
	LUT4 #(
		.INIT('h9009)
	) name5986 (
		_w5963_,
		_w6046_,
		_w6047_,
		_w6050_,
		_w6052_
	);
	LUT4 #(
		.INIT('h6996)
	) name5987 (
		_w5963_,
		_w6046_,
		_w6047_,
		_w6050_,
		_w6053_
	);
	LUT2 #(
		.INIT('h8)
	) name5988 (
		\a[15] ,
		\a[63] ,
		_w6054_
	);
	LUT4 #(
		.INIT('h153f)
	) name5989 (
		\a[16] ,
		\a[17] ,
		\a[61] ,
		\a[62] ,
		_w6055_
	);
	LUT4 #(
		.INIT('h8000)
	) name5990 (
		\a[16] ,
		\a[17] ,
		\a[61] ,
		\a[62] ,
		_w6056_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5991 (
		\a[16] ,
		\a[17] ,
		\a[61] ,
		\a[62] ,
		_w6057_
	);
	LUT2 #(
		.INIT('h6)
	) name5992 (
		_w6054_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h6)
	) name5993 (
		_w6053_,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h8)
	) name5994 (
		\a[20] ,
		\a[58] ,
		_w6060_
	);
	LUT4 #(
		.INIT('h153f)
	) name5995 (
		\a[30] ,
		\a[31] ,
		\a[47] ,
		\a[48] ,
		_w6061_
	);
	LUT2 #(
		.INIT('h8)
	) name5996 (
		\a[31] ,
		\a[48] ,
		_w6062_
	);
	LUT4 #(
		.INIT('h8000)
	) name5997 (
		\a[30] ,
		\a[31] ,
		\a[47] ,
		\a[48] ,
		_w6063_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name5998 (
		\a[30] ,
		\a[31] ,
		\a[47] ,
		\a[48] ,
		_w6064_
	);
	LUT2 #(
		.INIT('h8)
	) name5999 (
		\a[32] ,
		\a[46] ,
		_w6065_
	);
	LUT4 #(
		.INIT('h153f)
	) name6000 (
		\a[33] ,
		\a[34] ,
		\a[44] ,
		\a[45] ,
		_w6066_
	);
	LUT4 #(
		.INIT('h8000)
	) name6001 (
		\a[33] ,
		\a[34] ,
		\a[44] ,
		\a[45] ,
		_w6067_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6002 (
		\a[33] ,
		\a[34] ,
		\a[44] ,
		\a[45] ,
		_w6068_
	);
	LUT4 #(
		.INIT('h0660)
	) name6003 (
		_w6060_,
		_w6064_,
		_w6065_,
		_w6068_,
		_w6069_
	);
	LUT4 #(
		.INIT('h9009)
	) name6004 (
		_w6060_,
		_w6064_,
		_w6065_,
		_w6068_,
		_w6070_
	);
	LUT4 #(
		.INIT('h6996)
	) name6005 (
		_w6060_,
		_w6064_,
		_w6065_,
		_w6068_,
		_w6071_
	);
	LUT2 #(
		.INIT('h8)
	) name6006 (
		\a[25] ,
		\a[53] ,
		_w6072_
	);
	LUT4 #(
		.INIT('h153f)
	) name6007 (
		\a[22] ,
		\a[24] ,
		\a[54] ,
		\a[56] ,
		_w6073_
	);
	LUT4 #(
		.INIT('h8000)
	) name6008 (
		\a[22] ,
		\a[24] ,
		\a[54] ,
		\a[56] ,
		_w6074_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6009 (
		\a[22] ,
		\a[24] ,
		\a[54] ,
		\a[56] ,
		_w6075_
	);
	LUT2 #(
		.INIT('h6)
	) name6010 (
		_w6072_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h6)
	) name6011 (
		_w6071_,
		_w6076_,
		_w6077_
	);
	LUT4 #(
		.INIT('h6996)
	) name6012 (
		_w6053_,
		_w6058_,
		_w6071_,
		_w6076_,
		_w6078_
	);
	LUT3 #(
		.INIT('he1)
	) name6013 (
		_w6020_,
		_w6043_,
		_w6078_,
		_w6079_
	);
	LUT4 #(
		.INIT('hba00)
	) name6014 (
		_w5973_,
		_w5974_,
		_w5984_,
		_w6079_,
		_w6080_
	);
	LUT4 #(
		.INIT('h0045)
	) name6015 (
		_w5973_,
		_w5974_,
		_w5984_,
		_w6079_,
		_w6081_
	);
	LUT4 #(
		.INIT('h45ba)
	) name6016 (
		_w5973_,
		_w5974_,
		_w5984_,
		_w6079_,
		_w6082_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6017 (
		_w6026_,
		_w6040_,
		_w6041_,
		_w6082_,
		_w6083_
	);
	LUT4 #(
		.INIT('h0040)
	) name6018 (
		_w6026_,
		_w6040_,
		_w6041_,
		_w6081_,
		_w6084_
	);
	LUT3 #(
		.INIT('h23)
	) name6019 (
		_w6080_,
		_w6083_,
		_w6084_,
		_w6085_
	);
	LUT4 #(
		.INIT('h8882)
	) name6020 (
		_w5986_,
		_w6042_,
		_w6080_,
		_w6081_,
		_w6086_
	);
	LUT3 #(
		.INIT('h07)
	) name6021 (
		_w6029_,
		_w6085_,
		_w6086_,
		_w6087_
	);
	LUT3 #(
		.INIT('h1e)
	) name6022 (
		_w5986_,
		_w6029_,
		_w6085_,
		_w6088_
	);
	LUT3 #(
		.INIT('h07)
	) name6023 (
		_w5935_,
		_w5937_,
		_w5958_,
		_w6089_
	);
	LUT4 #(
		.INIT('h00f8)
	) name6024 (
		_w5935_,
		_w5937_,
		_w5958_,
		_w5959_,
		_w6090_
	);
	LUT3 #(
		.INIT('hb2)
	) name6025 (
		_w6007_,
		_w6008_,
		_w6012_,
		_w6091_
	);
	LUT3 #(
		.INIT('h32)
	) name6026 (
		_w5998_,
		_w5999_,
		_w6001_,
		_w6092_
	);
	LUT3 #(
		.INIT('h45)
	) name6027 (
		_w5945_,
		_w5946_,
		_w5952_,
		_w6093_
	);
	LUT3 #(
		.INIT('h96)
	) name6028 (
		_w6091_,
		_w6092_,
		_w6093_,
		_w6094_
	);
	LUT3 #(
		.INIT('hd4)
	) name6029 (
		_w5978_,
		_w5982_,
		_w5983_,
		_w6095_
	);
	LUT4 #(
		.INIT('he0c0)
	) name6030 (
		\a[15] ,
		\a[38] ,
		\a[39] ,
		\a[62] ,
		_w6096_
	);
	LUT4 #(
		.INIT('h000d)
	) name6031 (
		_w5989_,
		_w5990_,
		_w5992_,
		_w6096_,
		_w6097_
	);
	LUT4 #(
		.INIT('hf200)
	) name6032 (
		_w5989_,
		_w5990_,
		_w5992_,
		_w6096_,
		_w6098_
	);
	LUT4 #(
		.INIT('h0df2)
	) name6033 (
		_w5989_,
		_w5990_,
		_w5992_,
		_w6096_,
		_w6099_
	);
	LUT3 #(
		.INIT('h0d)
	) name6034 (
		_w5885_,
		_w5942_,
		_w5943_,
		_w6100_
	);
	LUT2 #(
		.INIT('h6)
	) name6035 (
		_w6099_,
		_w6100_,
		_w6101_
	);
	LUT3 #(
		.INIT('h0d)
	) name6036 (
		_w5873_,
		_w5994_,
		_w5996_,
		_w6102_
	);
	LUT3 #(
		.INIT('h0d)
	) name6037 (
		_w5899_,
		_w6009_,
		_w6010_,
		_w6103_
	);
	LUT3 #(
		.INIT('h0d)
	) name6038 (
		_w5948_,
		_w5949_,
		_w5950_,
		_w6104_
	);
	LUT3 #(
		.INIT('h96)
	) name6039 (
		_w6102_,
		_w6103_,
		_w6104_,
		_w6105_
	);
	LUT3 #(
		.INIT('h71)
	) name6040 (
		_w5979_,
		_w5980_,
		_w5981_,
		_w6106_
	);
	LUT3 #(
		.INIT('h96)
	) name6041 (
		_w6101_,
		_w6105_,
		_w6106_,
		_w6107_
	);
	LUT3 #(
		.INIT('h69)
	) name6042 (
		_w6094_,
		_w6095_,
		_w6107_,
		_w6108_
	);
	LUT3 #(
		.INIT('h54)
	) name6043 (
		_w5967_,
		_w5968_,
		_w5970_,
		_w6109_
	);
	LUT3 #(
		.INIT('h32)
	) name6044 (
		_w5938_,
		_w5939_,
		_w5940_,
		_w6110_
	);
	LUT3 #(
		.INIT('h0d)
	) name6045 (
		_w6003_,
		_w6004_,
		_w6005_,
		_w6111_
	);
	LUT4 #(
		.INIT('h153f)
	) name6046 (
		\a[17] ,
		\a[18] ,
		\a[59] ,
		\a[60] ,
		_w6112_
	);
	LUT4 #(
		.INIT('h000d)
	) name6047 (
		_w5883_,
		_w5884_,
		_w5886_,
		_w5964_,
		_w6113_
	);
	LUT4 #(
		.INIT('h9996)
	) name6048 (
		_w6110_,
		_w6111_,
		_w6112_,
		_w6113_,
		_w6114_
	);
	LUT2 #(
		.INIT('h8)
	) name6049 (
		\a[23] ,
		\a[55] ,
		_w6115_
	);
	LUT4 #(
		.INIT('h153f)
	) name6050 (
		\a[35] ,
		\a[36] ,
		\a[42] ,
		\a[43] ,
		_w6116_
	);
	LUT2 #(
		.INIT('h8)
	) name6051 (
		\a[36] ,
		\a[43] ,
		_w6117_
	);
	LUT4 #(
		.INIT('h8000)
	) name6052 (
		\a[35] ,
		\a[36] ,
		\a[42] ,
		\a[43] ,
		_w6118_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6053 (
		\a[35] ,
		\a[36] ,
		\a[42] ,
		\a[43] ,
		_w6119_
	);
	LUT2 #(
		.INIT('h8)
	) name6054 (
		\a[26] ,
		\a[52] ,
		_w6120_
	);
	LUT2 #(
		.INIT('h8)
	) name6055 (
		\a[38] ,
		\a[40] ,
		_w6121_
	);
	LUT4 #(
		.INIT('h153f)
	) name6056 (
		\a[26] ,
		\a[38] ,
		\a[40] ,
		\a[52] ,
		_w6122_
	);
	LUT4 #(
		.INIT('h8000)
	) name6057 (
		\a[26] ,
		\a[38] ,
		\a[40] ,
		\a[52] ,
		_w6123_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6058 (
		\a[26] ,
		\a[38] ,
		\a[40] ,
		\a[52] ,
		_w6124_
	);
	LUT4 #(
		.INIT('h1428)
	) name6059 (
		_w5991_,
		_w6115_,
		_w6119_,
		_w6124_,
		_w6125_
	);
	LUT4 #(
		.INIT('h6996)
	) name6060 (
		_w5991_,
		_w6115_,
		_w6119_,
		_w6124_,
		_w6126_
	);
	LUT4 #(
		.INIT('h1700)
	) name6061 (
		_w5975_,
		_w5976_,
		_w5977_,
		_w6126_,
		_w6127_
	);
	LUT4 #(
		.INIT('he817)
	) name6062 (
		_w5975_,
		_w5976_,
		_w5977_,
		_w6126_,
		_w6128_
	);
	LUT2 #(
		.INIT('h4)
	) name6063 (
		_w6114_,
		_w6128_,
		_w6129_
	);
	LUT2 #(
		.INIT('h8)
	) name6064 (
		_w6114_,
		_w6128_,
		_w6130_
	);
	LUT3 #(
		.INIT('h69)
	) name6065 (
		_w6109_,
		_w6114_,
		_w6128_,
		_w6131_
	);
	LUT3 #(
		.INIT('h54)
	) name6066 (
		_w5954_,
		_w5955_,
		_w5956_,
		_w6132_
	);
	LUT3 #(
		.INIT('h17)
	) name6067 (
		_w5988_,
		_w6002_,
		_w6013_,
		_w6133_
	);
	LUT3 #(
		.INIT('h96)
	) name6068 (
		_w6131_,
		_w6132_,
		_w6133_,
		_w6134_
	);
	LUT3 #(
		.INIT('h9f)
	) name6069 (
		_w6090_,
		_w6108_,
		_w6134_,
		_w6135_
	);
	LUT2 #(
		.INIT('h1)
	) name6070 (
		_w5959_,
		_w6134_,
		_w6136_
	);
	LUT3 #(
		.INIT('h40)
	) name6071 (
		_w6089_,
		_w6108_,
		_w6136_,
		_w6137_
	);
	LUT4 #(
		.INIT('h1441)
	) name6072 (
		_w6108_,
		_w6131_,
		_w6132_,
		_w6133_,
		_w6138_
	);
	LUT2 #(
		.INIT('h4)
	) name6073 (
		_w6090_,
		_w6138_,
		_w6139_
	);
	LUT3 #(
		.INIT('h02)
	) name6074 (
		_w6135_,
		_w6137_,
		_w6139_,
		_w6140_
	);
	LUT3 #(
		.INIT('h14)
	) name6075 (
		_w6039_,
		_w6088_,
		_w6140_,
		_w6141_
	);
	LUT3 #(
		.INIT('h82)
	) name6076 (
		_w6039_,
		_w6088_,
		_w6140_,
		_w6142_
	);
	LUT3 #(
		.INIT('h69)
	) name6077 (
		_w6039_,
		_w6088_,
		_w6140_,
		_w6143_
	);
	LUT4 #(
		.INIT('h23dc)
	) name6078 (
		_w5930_,
		_w6033_,
		_w6038_,
		_w6143_,
		_w6144_
	);
	LUT2 #(
		.INIT('h1)
	) name6079 (
		_w6033_,
		_w6141_,
		_w6145_
	);
	LUT3 #(
		.INIT('h45)
	) name6080 (
		_w5986_,
		_w5987_,
		_w6028_,
		_w6146_
	);
	LUT2 #(
		.INIT('h4)
	) name6081 (
		_w6085_,
		_w6146_,
		_w6147_
	);
	LUT3 #(
		.INIT('h0d)
	) name6082 (
		_w6087_,
		_w6140_,
		_w6147_,
		_w6148_
	);
	LUT3 #(
		.INIT('h4d)
	) name6083 (
		_w6131_,
		_w6132_,
		_w6133_,
		_w6149_
	);
	LUT3 #(
		.INIT('h0d)
	) name6084 (
		_w6047_,
		_w6048_,
		_w6049_,
		_w6150_
	);
	LUT3 #(
		.INIT('h0d)
	) name6085 (
		_w5963_,
		_w6044_,
		_w6045_,
		_w6151_
	);
	LUT3 #(
		.INIT('h0d)
	) name6086 (
		_w6072_,
		_w6073_,
		_w6074_,
		_w6152_
	);
	LUT3 #(
		.INIT('h96)
	) name6087 (
		_w6150_,
		_w6151_,
		_w6152_,
		_w6153_
	);
	LUT3 #(
		.INIT('h10)
	) name6088 (
		_w6125_,
		_w6127_,
		_w6153_,
		_w6154_
	);
	LUT3 #(
		.INIT('h0e)
	) name6089 (
		_w6125_,
		_w6127_,
		_w6153_,
		_w6155_
	);
	LUT3 #(
		.INIT('he1)
	) name6090 (
		_w6125_,
		_w6127_,
		_w6153_,
		_w6156_
	);
	LUT4 #(
		.INIT('h222b)
	) name6091 (
		_w6110_,
		_w6111_,
		_w6112_,
		_w6113_,
		_w6157_
	);
	LUT2 #(
		.INIT('h8)
	) name6092 (
		\a[16] ,
		\a[63] ,
		_w6158_
	);
	LUT4 #(
		.INIT('h153f)
	) name6093 (
		\a[34] ,
		\a[35] ,
		\a[44] ,
		\a[45] ,
		_w6159_
	);
	LUT4 #(
		.INIT('h8000)
	) name6094 (
		\a[34] ,
		\a[35] ,
		\a[44] ,
		\a[45] ,
		_w6160_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6095 (
		\a[34] ,
		\a[35] ,
		\a[44] ,
		\a[45] ,
		_w6161_
	);
	LUT2 #(
		.INIT('h6)
	) name6096 (
		_w6158_,
		_w6161_,
		_w6162_
	);
	LUT4 #(
		.INIT('h153f)
	) name6097 (
		\a[23] ,
		\a[27] ,
		\a[52] ,
		\a[56] ,
		_w6163_
	);
	LUT2 #(
		.INIT('h8)
	) name6098 (
		\a[27] ,
		\a[56] ,
		_w6164_
	);
	LUT4 #(
		.INIT('h8000)
	) name6099 (
		\a[23] ,
		\a[27] ,
		\a[52] ,
		\a[56] ,
		_w6165_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6100 (
		\a[23] ,
		\a[27] ,
		\a[52] ,
		\a[56] ,
		_w6166_
	);
	LUT2 #(
		.INIT('h6)
	) name6101 (
		_w6117_,
		_w6166_,
		_w6167_
	);
	LUT4 #(
		.INIT('h1428)
	) name6102 (
		_w6117_,
		_w6158_,
		_w6161_,
		_w6166_,
		_w6168_
	);
	LUT4 #(
		.INIT('h8241)
	) name6103 (
		_w6117_,
		_w6158_,
		_w6161_,
		_w6166_,
		_w6169_
	);
	LUT4 #(
		.INIT('h6996)
	) name6104 (
		_w6117_,
		_w6158_,
		_w6161_,
		_w6166_,
		_w6170_
	);
	LUT2 #(
		.INIT('h6)
	) name6105 (
		_w6157_,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('h6)
	) name6106 (
		_w6156_,
		_w6171_,
		_w6172_
	);
	LUT4 #(
		.INIT('hf110)
	) name6107 (
		_w6020_,
		_w6043_,
		_w6059_,
		_w6077_,
		_w6173_
	);
	LUT2 #(
		.INIT('h8)
	) name6108 (
		\a[18] ,
		\a[61] ,
		_w6174_
	);
	LUT4 #(
		.INIT('he800)
	) name6109 (
		_w5991_,
		_w6120_,
		_w6121_,
		_w6174_,
		_w6175_
	);
	LUT4 #(
		.INIT('h153f)
	) name6110 (
		\a[18] ,
		\a[37] ,
		\a[41] ,
		\a[61] ,
		_w6176_
	);
	LUT4 #(
		.INIT('h88fe)
	) name6111 (
		_w6120_,
		_w6121_,
		_w6174_,
		_w6176_,
		_w6177_
	);
	LUT4 #(
		.INIT('hcd32)
	) name6112 (
		_w5991_,
		_w6122_,
		_w6123_,
		_w6174_,
		_w6178_
	);
	LUT3 #(
		.INIT('h0d)
	) name6113 (
		_w6115_,
		_w6116_,
		_w6118_,
		_w6179_
	);
	LUT2 #(
		.INIT('h6)
	) name6114 (
		_w6178_,
		_w6179_,
		_w6180_
	);
	LUT3 #(
		.INIT('h0d)
	) name6115 (
		_w6054_,
		_w6055_,
		_w6056_,
		_w6181_
	);
	LUT3 #(
		.INIT('h0d)
	) name6116 (
		_w6060_,
		_w6061_,
		_w6063_,
		_w6182_
	);
	LUT3 #(
		.INIT('h0d)
	) name6117 (
		_w6065_,
		_w6066_,
		_w6067_,
		_w6183_
	);
	LUT3 #(
		.INIT('h96)
	) name6118 (
		_w6181_,
		_w6182_,
		_w6183_,
		_w6184_
	);
	LUT3 #(
		.INIT('h32)
	) name6119 (
		_w6069_,
		_w6070_,
		_w6076_,
		_w6185_
	);
	LUT3 #(
		.INIT('h96)
	) name6120 (
		_w6180_,
		_w6184_,
		_w6185_,
		_w6186_
	);
	LUT3 #(
		.INIT('h96)
	) name6121 (
		_w6172_,
		_w6173_,
		_w6186_,
		_w6187_
	);
	LUT2 #(
		.INIT('h1)
	) name6122 (
		_w6149_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h8)
	) name6123 (
		_w6149_,
		_w6187_,
		_w6189_
	);
	LUT2 #(
		.INIT('h6)
	) name6124 (
		_w6149_,
		_w6187_,
		_w6190_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6125 (
		_w6026_,
		_w6040_,
		_w6041_,
		_w6080_,
		_w6191_
	);
	LUT3 #(
		.INIT('hc9)
	) name6126 (
		_w6081_,
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT2 #(
		.INIT('h4)
	) name6127 (
		_w5959_,
		_w6108_,
		_w6193_
	);
	LUT2 #(
		.INIT('h4)
	) name6128 (
		_w6089_,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h8)
	) name6129 (
		\a[24] ,
		\a[55] ,
		_w6195_
	);
	LUT4 #(
		.INIT('h153f)
	) name6130 (
		\a[25] ,
		\a[26] ,
		\a[53] ,
		\a[54] ,
		_w6196_
	);
	LUT4 #(
		.INIT('h8000)
	) name6131 (
		\a[25] ,
		\a[26] ,
		\a[53] ,
		\a[54] ,
		_w6197_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6132 (
		\a[25] ,
		\a[26] ,
		\a[53] ,
		\a[54] ,
		_w6198_
	);
	LUT2 #(
		.INIT('h8)
	) name6133 (
		\a[37] ,
		\a[42] ,
		_w6199_
	);
	LUT4 #(
		.INIT('h153f)
	) name6134 (
		\a[38] ,
		\a[39] ,
		\a[40] ,
		\a[41] ,
		_w6200_
	);
	LUT2 #(
		.INIT('h8)
	) name6135 (
		\a[39] ,
		\a[41] ,
		_w6201_
	);
	LUT4 #(
		.INIT('h8000)
	) name6136 (
		\a[38] ,
		\a[39] ,
		\a[40] ,
		\a[41] ,
		_w6202_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6137 (
		\a[38] ,
		\a[39] ,
		\a[40] ,
		\a[41] ,
		_w6203_
	);
	LUT4 #(
		.INIT('h0660)
	) name6138 (
		_w6195_,
		_w6198_,
		_w6199_,
		_w6203_,
		_w6204_
	);
	LUT4 #(
		.INIT('h9009)
	) name6139 (
		_w6195_,
		_w6198_,
		_w6199_,
		_w6203_,
		_w6205_
	);
	LUT4 #(
		.INIT('h6996)
	) name6140 (
		_w6195_,
		_w6198_,
		_w6199_,
		_w6203_,
		_w6206_
	);
	LUT2 #(
		.INIT('h8)
	) name6141 (
		\a[28] ,
		\a[51] ,
		_w6207_
	);
	LUT3 #(
		.INIT('h13)
	) name6142 (
		\a[17] ,
		\a[40] ,
		\a[62] ,
		_w6208_
	);
	LUT2 #(
		.INIT('h8)
	) name6143 (
		\a[40] ,
		\a[62] ,
		_w6209_
	);
	LUT3 #(
		.INIT('h80)
	) name6144 (
		\a[17] ,
		\a[40] ,
		\a[62] ,
		_w6210_
	);
	LUT3 #(
		.INIT('h6c)
	) name6145 (
		\a[17] ,
		\a[40] ,
		\a[62] ,
		_w6211_
	);
	LUT2 #(
		.INIT('h6)
	) name6146 (
		_w6207_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h8)
	) name6147 (
		\a[19] ,
		\a[60] ,
		_w6213_
	);
	LUT4 #(
		.INIT('h153f)
	) name6148 (
		\a[20] ,
		\a[21] ,
		\a[58] ,
		\a[59] ,
		_w6214_
	);
	LUT4 #(
		.INIT('h8000)
	) name6149 (
		\a[20] ,
		\a[21] ,
		\a[58] ,
		\a[59] ,
		_w6215_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6150 (
		\a[20] ,
		\a[21] ,
		\a[58] ,
		\a[59] ,
		_w6216_
	);
	LUT2 #(
		.INIT('h8)
	) name6151 (
		\a[22] ,
		\a[57] ,
		_w6217_
	);
	LUT4 #(
		.INIT('h153f)
	) name6152 (
		\a[29] ,
		\a[30] ,
		\a[49] ,
		\a[50] ,
		_w6218_
	);
	LUT2 #(
		.INIT('h8)
	) name6153 (
		\a[30] ,
		\a[50] ,
		_w6219_
	);
	LUT4 #(
		.INIT('h8000)
	) name6154 (
		\a[29] ,
		\a[30] ,
		\a[49] ,
		\a[50] ,
		_w6220_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6155 (
		\a[29] ,
		\a[30] ,
		\a[49] ,
		\a[50] ,
		_w6221_
	);
	LUT4 #(
		.INIT('h0660)
	) name6156 (
		_w6213_,
		_w6216_,
		_w6217_,
		_w6221_,
		_w6222_
	);
	LUT4 #(
		.INIT('h9009)
	) name6157 (
		_w6213_,
		_w6216_,
		_w6217_,
		_w6221_,
		_w6223_
	);
	LUT4 #(
		.INIT('h6996)
	) name6158 (
		_w6213_,
		_w6216_,
		_w6217_,
		_w6221_,
		_w6224_
	);
	LUT4 #(
		.INIT('h153f)
	) name6159 (
		\a[32] ,
		\a[33] ,
		\a[46] ,
		\a[47] ,
		_w6225_
	);
	LUT2 #(
		.INIT('h8)
	) name6160 (
		\a[33] ,
		\a[47] ,
		_w6226_
	);
	LUT4 #(
		.INIT('h8000)
	) name6161 (
		\a[32] ,
		\a[33] ,
		\a[46] ,
		\a[47] ,
		_w6227_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6162 (
		\a[32] ,
		\a[33] ,
		\a[46] ,
		\a[47] ,
		_w6228_
	);
	LUT2 #(
		.INIT('h6)
	) name6163 (
		_w6062_,
		_w6228_,
		_w6229_
	);
	LUT4 #(
		.INIT('h0660)
	) name6164 (
		_w6206_,
		_w6212_,
		_w6224_,
		_w6229_,
		_w6230_
	);
	LUT4 #(
		.INIT('h6996)
	) name6165 (
		_w6206_,
		_w6212_,
		_w6224_,
		_w6229_,
		_w6231_
	);
	LUT4 #(
		.INIT('h7100)
	) name6166 (
		_w6101_,
		_w6105_,
		_w6106_,
		_w6231_,
		_w6232_
	);
	LUT4 #(
		.INIT('h8e71)
	) name6167 (
		_w6101_,
		_w6105_,
		_w6106_,
		_w6231_,
		_w6233_
	);
	LUT4 #(
		.INIT('h002b)
	) name6168 (
		_w6094_,
		_w6095_,
		_w6107_,
		_w6233_,
		_w6234_
	);
	LUT4 #(
		.INIT('hd400)
	) name6169 (
		_w6094_,
		_w6095_,
		_w6107_,
		_w6233_,
		_w6235_
	);
	LUT3 #(
		.INIT('h17)
	) name6170 (
		_w6102_,
		_w6103_,
		_w6104_,
		_w6236_
	);
	LUT3 #(
		.INIT('h45)
	) name6171 (
		_w6097_,
		_w6098_,
		_w6100_,
		_w6237_
	);
	LUT3 #(
		.INIT('h32)
	) name6172 (
		_w6051_,
		_w6052_,
		_w6058_,
		_w6238_
	);
	LUT3 #(
		.INIT('h96)
	) name6173 (
		_w6236_,
		_w6237_,
		_w6238_,
		_w6239_
	);
	LUT3 #(
		.INIT('h8e)
	) name6174 (
		_w6091_,
		_w6092_,
		_w6093_,
		_w6240_
	);
	LUT2 #(
		.INIT('h1)
	) name6175 (
		_w6239_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h8)
	) name6176 (
		_w6239_,
		_w6240_,
		_w6242_
	);
	LUT2 #(
		.INIT('h6)
	) name6177 (
		_w6239_,
		_w6240_,
		_w6243_
	);
	LUT4 #(
		.INIT('hb200)
	) name6178 (
		_w5962_,
		_w5966_,
		_w5970_,
		_w6114_,
		_w6244_
	);
	LUT4 #(
		.INIT('h0027)
	) name6179 (
		_w6109_,
		_w6129_,
		_w6130_,
		_w6244_,
		_w6245_
	);
	LUT4 #(
		.INIT('he11e)
	) name6180 (
		_w6234_,
		_w6235_,
		_w6243_,
		_w6245_,
		_w6246_
	);
	LUT3 #(
		.INIT('h40)
	) name6181 (
		_w6089_,
		_w6193_,
		_w6246_,
		_w6247_
	);
	LUT2 #(
		.INIT('h2)
	) name6182 (
		_w5959_,
		_w6108_,
		_w6248_
	);
	LUT4 #(
		.INIT('h0007)
	) name6183 (
		_w5935_,
		_w5937_,
		_w5958_,
		_w6108_,
		_w6249_
	);
	LUT3 #(
		.INIT('h02)
	) name6184 (
		_w6134_,
		_w6248_,
		_w6249_,
		_w6250_
	);
	LUT4 #(
		.INIT('h0008)
	) name6185 (
		_w6134_,
		_w6246_,
		_w6248_,
		_w6249_,
		_w6251_
	);
	LUT2 #(
		.INIT('h1)
	) name6186 (
		_w6247_,
		_w6251_,
		_w6252_
	);
	LUT3 #(
		.INIT('h0b)
	) name6187 (
		_w6089_,
		_w6193_,
		_w6246_,
		_w6253_
	);
	LUT4 #(
		.INIT('h0d3d)
	) name6188 (
		_w6135_,
		_w6194_,
		_w6246_,
		_w6250_,
		_w6254_
	);
	LUT2 #(
		.INIT('h9)
	) name6189 (
		_w6192_,
		_w6254_,
		_w6255_
	);
	LUT3 #(
		.INIT('h96)
	) name6190 (
		_w6142_,
		_w6148_,
		_w6255_,
		_w6256_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6191 (
		_w5930_,
		_w6038_,
		_w6145_,
		_w6256_,
		_w6257_
	);
	LUT3 #(
		.INIT('hc3)
	) name6192 (
		_w6142_,
		_w6148_,
		_w6255_,
		_w6258_
	);
	LUT4 #(
		.INIT('hb000)
	) name6193 (
		_w5930_,
		_w6038_,
		_w6145_,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('he)
	) name6194 (
		_w6257_,
		_w6259_,
		_w6260_
	);
	LUT4 #(
		.INIT('h1101)
	) name6195 (
		_w6033_,
		_w6141_,
		_w6148_,
		_w6255_,
		_w6261_
	);
	LUT3 #(
		.INIT('h4c)
	) name6196 (
		_w6135_,
		_w6192_,
		_w6253_,
		_w6262_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name6197 (
		_w6081_,
		_w6188_,
		_w6189_,
		_w6191_,
		_w6263_
	);
	LUT3 #(
		.INIT('he8)
	) name6198 (
		_w6172_,
		_w6173_,
		_w6186_,
		_w6264_
	);
	LUT4 #(
		.INIT('h8000)
	) name6199 (
		\a[18] ,
		\a[19] ,
		\a[61] ,
		\a[62] ,
		_w6265_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6200 (
		\a[18] ,
		\a[19] ,
		\a[61] ,
		\a[62] ,
		_w6266_
	);
	LUT4 #(
		.INIT('hf20d)
	) name6201 (
		_w6207_,
		_w6208_,
		_w6210_,
		_w6266_,
		_w6267_
	);
	LUT4 #(
		.INIT('h153f)
	) name6202 (
		\a[17] ,
		\a[29] ,
		\a[51] ,
		\a[63] ,
		_w6268_
	);
	LUT4 #(
		.INIT('h8000)
	) name6203 (
		\a[17] ,
		\a[29] ,
		\a[51] ,
		\a[63] ,
		_w6269_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6204 (
		\a[17] ,
		\a[29] ,
		\a[51] ,
		\a[63] ,
		_w6270_
	);
	LUT2 #(
		.INIT('h8)
	) name6205 (
		\a[34] ,
		\a[46] ,
		_w6271_
	);
	LUT4 #(
		.INIT('h153f)
	) name6206 (
		\a[35] ,
		\a[36] ,
		\a[44] ,
		\a[45] ,
		_w6272_
	);
	LUT4 #(
		.INIT('h8000)
	) name6207 (
		\a[35] ,
		\a[36] ,
		\a[44] ,
		\a[45] ,
		_w6273_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6208 (
		\a[35] ,
		\a[36] ,
		\a[44] ,
		\a[45] ,
		_w6274_
	);
	LUT4 #(
		.INIT('h0660)
	) name6209 (
		_w6226_,
		_w6270_,
		_w6271_,
		_w6274_,
		_w6275_
	);
	LUT4 #(
		.INIT('h9009)
	) name6210 (
		_w6226_,
		_w6270_,
		_w6271_,
		_w6274_,
		_w6276_
	);
	LUT4 #(
		.INIT('h6996)
	) name6211 (
		_w6226_,
		_w6270_,
		_w6271_,
		_w6274_,
		_w6277_
	);
	LUT2 #(
		.INIT('h9)
	) name6212 (
		_w6267_,
		_w6277_,
		_w6278_
	);
	LUT4 #(
		.INIT('h153f)
	) name6213 (
		\a[21] ,
		\a[22] ,
		\a[58] ,
		\a[59] ,
		_w6279_
	);
	LUT2 #(
		.INIT('h8)
	) name6214 (
		\a[22] ,
		\a[59] ,
		_w6280_
	);
	LUT4 #(
		.INIT('h8000)
	) name6215 (
		\a[21] ,
		\a[22] ,
		\a[58] ,
		\a[59] ,
		_w6281_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6216 (
		\a[21] ,
		\a[22] ,
		\a[58] ,
		\a[59] ,
		_w6282_
	);
	LUT2 #(
		.INIT('h8)
	) name6217 (
		\a[20] ,
		\a[60] ,
		_w6283_
	);
	LUT2 #(
		.INIT('h6)
	) name6218 (
		_w6282_,
		_w6283_,
		_w6284_
	);
	LUT3 #(
		.INIT('h0d)
	) name6219 (
		_w6199_,
		_w6200_,
		_w6202_,
		_w6285_
	);
	LUT4 #(
		.INIT('h153f)
	) name6220 (
		\a[31] ,
		\a[32] ,
		\a[48] ,
		\a[49] ,
		_w6286_
	);
	LUT4 #(
		.INIT('h8000)
	) name6221 (
		\a[31] ,
		\a[32] ,
		\a[48] ,
		\a[49] ,
		_w6287_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6222 (
		\a[31] ,
		\a[32] ,
		\a[48] ,
		\a[49] ,
		_w6288_
	);
	LUT2 #(
		.INIT('h6)
	) name6223 (
		_w6219_,
		_w6288_,
		_w6289_
	);
	LUT3 #(
		.INIT('h69)
	) name6224 (
		_w6284_,
		_w6285_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h8)
	) name6225 (
		\a[23] ,
		\a[57] ,
		_w6291_
	);
	LUT4 #(
		.INIT('h153f)
	) name6226 (
		\a[24] ,
		\a[26] ,
		\a[54] ,
		\a[56] ,
		_w6292_
	);
	LUT2 #(
		.INIT('h8)
	) name6227 (
		\a[26] ,
		\a[56] ,
		_w6293_
	);
	LUT4 #(
		.INIT('h8000)
	) name6228 (
		\a[24] ,
		\a[26] ,
		\a[54] ,
		\a[56] ,
		_w6294_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6229 (
		\a[24] ,
		\a[26] ,
		\a[54] ,
		\a[56] ,
		_w6295_
	);
	LUT2 #(
		.INIT('h8)
	) name6230 (
		\a[25] ,
		\a[55] ,
		_w6296_
	);
	LUT4 #(
		.INIT('h153f)
	) name6231 (
		\a[37] ,
		\a[38] ,
		\a[42] ,
		\a[43] ,
		_w6297_
	);
	LUT4 #(
		.INIT('h8000)
	) name6232 (
		\a[37] ,
		\a[38] ,
		\a[42] ,
		\a[43] ,
		_w6298_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6233 (
		\a[37] ,
		\a[38] ,
		\a[42] ,
		\a[43] ,
		_w6299_
	);
	LUT4 #(
		.INIT('h0660)
	) name6234 (
		_w6291_,
		_w6295_,
		_w6296_,
		_w6299_,
		_w6300_
	);
	LUT4 #(
		.INIT('h9009)
	) name6235 (
		_w6291_,
		_w6295_,
		_w6296_,
		_w6299_,
		_w6301_
	);
	LUT4 #(
		.INIT('h6996)
	) name6236 (
		_w6291_,
		_w6295_,
		_w6296_,
		_w6299_,
		_w6302_
	);
	LUT4 #(
		.INIT('h153f)
	) name6237 (
		\a[27] ,
		\a[28] ,
		\a[52] ,
		\a[53] ,
		_w6303_
	);
	LUT4 #(
		.INIT('h8000)
	) name6238 (
		\a[27] ,
		\a[28] ,
		\a[52] ,
		\a[53] ,
		_w6304_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6239 (
		\a[27] ,
		\a[28] ,
		\a[52] ,
		\a[53] ,
		_w6305_
	);
	LUT2 #(
		.INIT('h6)
	) name6240 (
		_w6201_,
		_w6305_,
		_w6306_
	);
	LUT2 #(
		.INIT('h6)
	) name6241 (
		_w6302_,
		_w6306_,
		_w6307_
	);
	LUT3 #(
		.INIT('h96)
	) name6242 (
		_w6278_,
		_w6290_,
		_w6307_,
		_w6308_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6243 (
		_w6239_,
		_w6240_,
		_w6245_,
		_w6308_,
		_w6309_
	);
	LUT3 #(
		.INIT('h07)
	) name6244 (
		_w6239_,
		_w6240_,
		_w6308_,
		_w6310_
	);
	LUT3 #(
		.INIT('hd0)
	) name6245 (
		_w6243_,
		_w6245_,
		_w6310_,
		_w6311_
	);
	LUT4 #(
		.INIT('h32cd)
	) name6246 (
		_w6241_,
		_w6242_,
		_w6245_,
		_w6308_,
		_w6312_
	);
	LUT2 #(
		.INIT('h9)
	) name6247 (
		_w6264_,
		_w6312_,
		_w6313_
	);
	LUT4 #(
		.INIT('h7007)
	) name6248 (
		_w6149_,
		_w6187_,
		_w6264_,
		_w6312_,
		_w6314_
	);
	LUT4 #(
		.INIT('hfb00)
	) name6249 (
		_w6081_,
		_w6190_,
		_w6191_,
		_w6314_,
		_w6315_
	);
	LUT4 #(
		.INIT('h5445)
	) name6250 (
		_w6234_,
		_w6235_,
		_w6243_,
		_w6245_,
		_w6316_
	);
	LUT3 #(
		.INIT('h0d)
	) name6251 (
		_w6158_,
		_w6159_,
		_w6160_,
		_w6317_
	);
	LUT3 #(
		.INIT('h0d)
	) name6252 (
		_w6195_,
		_w6196_,
		_w6197_,
		_w6318_
	);
	LUT3 #(
		.INIT('h0d)
	) name6253 (
		_w6117_,
		_w6163_,
		_w6165_,
		_w6319_
	);
	LUT3 #(
		.INIT('h96)
	) name6254 (
		_w6317_,
		_w6318_,
		_w6319_,
		_w6320_
	);
	LUT4 #(
		.INIT('h1700)
	) name6255 (
		_w6157_,
		_w6162_,
		_w6167_,
		_w6320_,
		_w6321_
	);
	LUT4 #(
		.INIT('h00e8)
	) name6256 (
		_w6157_,
		_w6162_,
		_w6167_,
		_w6320_,
		_w6322_
	);
	LUT4 #(
		.INIT('hce31)
	) name6257 (
		_w6157_,
		_w6168_,
		_w6169_,
		_w6320_,
		_w6323_
	);
	LUT3 #(
		.INIT('he8)
	) name6258 (
		_w6236_,
		_w6237_,
		_w6238_,
		_w6324_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name6259 (
		_w6230_,
		_w6232_,
		_w6323_,
		_w6324_,
		_w6325_
	);
	LUT4 #(
		.INIT('h1001)
	) name6260 (
		_w6230_,
		_w6232_,
		_w6323_,
		_w6324_,
		_w6326_
	);
	LUT4 #(
		.INIT('he11e)
	) name6261 (
		_w6230_,
		_w6232_,
		_w6323_,
		_w6324_,
		_w6327_
	);
	LUT3 #(
		.INIT('h0d)
	) name6262 (
		_w6217_,
		_w6218_,
		_w6220_,
		_w6328_
	);
	LUT3 #(
		.INIT('h0d)
	) name6263 (
		_w6213_,
		_w6214_,
		_w6215_,
		_w6329_
	);
	LUT3 #(
		.INIT('h0d)
	) name6264 (
		_w6062_,
		_w6225_,
		_w6227_,
		_w6330_
	);
	LUT3 #(
		.INIT('h96)
	) name6265 (
		_w6328_,
		_w6329_,
		_w6330_,
		_w6331_
	);
	LUT3 #(
		.INIT('h32)
	) name6266 (
		_w6204_,
		_w6205_,
		_w6212_,
		_w6332_
	);
	LUT3 #(
		.INIT('h32)
	) name6267 (
		_w6222_,
		_w6223_,
		_w6229_,
		_w6333_
	);
	LUT3 #(
		.INIT('h69)
	) name6268 (
		_w6331_,
		_w6332_,
		_w6333_,
		_w6334_
	);
	LUT2 #(
		.INIT('h6)
	) name6269 (
		_w6327_,
		_w6334_,
		_w6335_
	);
	LUT3 #(
		.INIT('h54)
	) name6270 (
		_w6154_,
		_w6155_,
		_w6171_,
		_w6336_
	);
	LUT3 #(
		.INIT('h17)
	) name6271 (
		_w6150_,
		_w6151_,
		_w6152_,
		_w6337_
	);
	LUT3 #(
		.INIT('h17)
	) name6272 (
		_w6181_,
		_w6182_,
		_w6183_,
		_w6338_
	);
	LUT3 #(
		.INIT('h51)
	) name6273 (
		_w6175_,
		_w6177_,
		_w6179_,
		_w6339_
	);
	LUT3 #(
		.INIT('h96)
	) name6274 (
		_w6337_,
		_w6338_,
		_w6339_,
		_w6340_
	);
	LUT3 #(
		.INIT('h71)
	) name6275 (
		_w6180_,
		_w6184_,
		_w6185_,
		_w6341_
	);
	LUT3 #(
		.INIT('h69)
	) name6276 (
		_w6336_,
		_w6340_,
		_w6341_,
		_w6342_
	);
	LUT3 #(
		.INIT('h96)
	) name6277 (
		_w6316_,
		_w6335_,
		_w6342_,
		_w6343_
	);
	LUT4 #(
		.INIT('hf10e)
	) name6278 (
		_w6263_,
		_w6313_,
		_w6315_,
		_w6343_,
		_w6344_
	);
	LUT3 #(
		.INIT('h02)
	) name6279 (
		_w6252_,
		_w6262_,
		_w6344_,
		_w6345_
	);
	LUT3 #(
		.INIT('hd0)
	) name6280 (
		_w6252_,
		_w6262_,
		_w6344_,
		_w6346_
	);
	LUT3 #(
		.INIT('h2d)
	) name6281 (
		_w6252_,
		_w6262_,
		_w6344_,
		_w6347_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6282 (
		_w6142_,
		_w6148_,
		_w6255_,
		_w6347_,
		_w6348_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6283 (
		_w5930_,
		_w6038_,
		_w6261_,
		_w6348_,
		_w6349_
	);
	LUT3 #(
		.INIT('h4d)
	) name6284 (
		_w6142_,
		_w6148_,
		_w6255_,
		_w6350_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6285 (
		_w5930_,
		_w6038_,
		_w6261_,
		_w6350_,
		_w6351_
	);
	LUT3 #(
		.INIT('h32)
	) name6286 (
		_w6347_,
		_w6349_,
		_w6351_,
		_w6352_
	);
	LUT4 #(
		.INIT('h004d)
	) name6287 (
		_w6142_,
		_w6148_,
		_w6255_,
		_w6345_,
		_w6353_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6288 (
		_w5930_,
		_w6038_,
		_w6261_,
		_w6353_,
		_w6354_
	);
	LUT4 #(
		.INIT('he0ee)
	) name6289 (
		_w6263_,
		_w6313_,
		_w6315_,
		_w6343_,
		_w6355_
	);
	LUT3 #(
		.INIT('he8)
	) name6290 (
		_w6316_,
		_w6335_,
		_w6342_,
		_w6356_
	);
	LUT3 #(
		.INIT('h32)
	) name6291 (
		_w6325_,
		_w6326_,
		_w6334_,
		_w6357_
	);
	LUT3 #(
		.INIT('h8e)
	) name6292 (
		_w6337_,
		_w6338_,
		_w6339_,
		_w6358_
	);
	LUT4 #(
		.INIT('h153f)
	) name6293 (
		\a[23] ,
		\a[25] ,
		\a[56] ,
		\a[58] ,
		_w6359_
	);
	LUT2 #(
		.INIT('h8)
	) name6294 (
		\a[25] ,
		\a[58] ,
		_w6360_
	);
	LUT4 #(
		.INIT('h8000)
	) name6295 (
		\a[23] ,
		\a[25] ,
		\a[56] ,
		\a[58] ,
		_w6361_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6296 (
		\a[23] ,
		\a[25] ,
		\a[56] ,
		\a[58] ,
		_w6362_
	);
	LUT4 #(
		.INIT('h9a30)
	) name6297 (
		\a[19] ,
		\a[40] ,
		\a[41] ,
		\a[62] ,
		_w6363_
	);
	LUT3 #(
		.INIT('h60)
	) name6298 (
		_w6280_,
		_w6362_,
		_w6363_,
		_w6364_
	);
	LUT3 #(
		.INIT('h09)
	) name6299 (
		_w6280_,
		_w6362_,
		_w6363_,
		_w6365_
	);
	LUT3 #(
		.INIT('h96)
	) name6300 (
		_w6280_,
		_w6362_,
		_w6363_,
		_w6366_
	);
	LUT4 #(
		.INIT('h153f)
	) name6301 (
		\a[33] ,
		\a[34] ,
		\a[47] ,
		\a[48] ,
		_w6367_
	);
	LUT4 #(
		.INIT('h8000)
	) name6302 (
		\a[33] ,
		\a[34] ,
		\a[47] ,
		\a[48] ,
		_w6368_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6303 (
		\a[33] ,
		\a[34] ,
		\a[47] ,
		\a[48] ,
		_w6369_
	);
	LUT2 #(
		.INIT('h6)
	) name6304 (
		_w4607_,
		_w6369_,
		_w6370_
	);
	LUT2 #(
		.INIT('h6)
	) name6305 (
		_w6366_,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h8)
	) name6306 (
		\a[18] ,
		\a[63] ,
		_w6372_
	);
	LUT4 #(
		.INIT('h153f)
	) name6307 (
		\a[20] ,
		\a[21] ,
		\a[60] ,
		\a[61] ,
		_w6373_
	);
	LUT4 #(
		.INIT('h8000)
	) name6308 (
		\a[20] ,
		\a[21] ,
		\a[60] ,
		\a[61] ,
		_w6374_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6309 (
		\a[20] ,
		\a[21] ,
		\a[60] ,
		\a[61] ,
		_w6375_
	);
	LUT2 #(
		.INIT('h8)
	) name6310 (
		\a[35] ,
		\a[46] ,
		_w6376_
	);
	LUT4 #(
		.INIT('h153f)
	) name6311 (
		\a[36] ,
		\a[37] ,
		\a[44] ,
		\a[45] ,
		_w6377_
	);
	LUT4 #(
		.INIT('h8000)
	) name6312 (
		\a[36] ,
		\a[37] ,
		\a[44] ,
		\a[45] ,
		_w6378_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6313 (
		\a[36] ,
		\a[37] ,
		\a[44] ,
		\a[45] ,
		_w6379_
	);
	LUT4 #(
		.INIT('h0660)
	) name6314 (
		_w6372_,
		_w6375_,
		_w6376_,
		_w6379_,
		_w6380_
	);
	LUT4 #(
		.INIT('h9009)
	) name6315 (
		_w6372_,
		_w6375_,
		_w6376_,
		_w6379_,
		_w6381_
	);
	LUT4 #(
		.INIT('h6996)
	) name6316 (
		_w6372_,
		_w6375_,
		_w6376_,
		_w6379_,
		_w6382_
	);
	LUT2 #(
		.INIT('h8)
	) name6317 (
		\a[26] ,
		\a[55] ,
		_w6383_
	);
	LUT4 #(
		.INIT('h153f)
	) name6318 (
		\a[28] ,
		\a[29] ,
		\a[52] ,
		\a[53] ,
		_w6384_
	);
	LUT4 #(
		.INIT('h8000)
	) name6319 (
		\a[28] ,
		\a[29] ,
		\a[52] ,
		\a[53] ,
		_w6385_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6320 (
		\a[28] ,
		\a[29] ,
		\a[52] ,
		\a[53] ,
		_w6386_
	);
	LUT2 #(
		.INIT('h6)
	) name6321 (
		_w6383_,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h6)
	) name6322 (
		_w6382_,
		_w6387_,
		_w6388_
	);
	LUT3 #(
		.INIT('h96)
	) name6323 (
		_w6358_,
		_w6371_,
		_w6388_,
		_w6389_
	);
	LUT4 #(
		.INIT('hb200)
	) name6324 (
		_w6336_,
		_w6340_,
		_w6341_,
		_w6389_,
		_w6390_
	);
	LUT4 #(
		.INIT('h004d)
	) name6325 (
		_w6336_,
		_w6340_,
		_w6341_,
		_w6389_,
		_w6391_
	);
	LUT4 #(
		.INIT('h4db2)
	) name6326 (
		_w6336_,
		_w6340_,
		_w6341_,
		_w6389_,
		_w6392_
	);
	LUT2 #(
		.INIT('h9)
	) name6327 (
		_w6357_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h2)
	) name6328 (
		_w6356_,
		_w6393_,
		_w6394_
	);
	LUT2 #(
		.INIT('h4)
	) name6329 (
		_w6356_,
		_w6393_,
		_w6395_
	);
	LUT2 #(
		.INIT('h9)
	) name6330 (
		_w6356_,
		_w6393_,
		_w6396_
	);
	LUT3 #(
		.INIT('he8)
	) name6331 (
		_w6278_,
		_w6290_,
		_w6307_,
		_w6397_
	);
	LUT3 #(
		.INIT('h0d)
	) name6332 (
		_w6219_,
		_w6286_,
		_w6287_,
		_w6398_
	);
	LUT3 #(
		.INIT('h0d)
	) name6333 (
		_w6226_,
		_w6268_,
		_w6269_,
		_w6399_
	);
	LUT3 #(
		.INIT('h23)
	) name6334 (
		_w6279_,
		_w6281_,
		_w6283_,
		_w6400_
	);
	LUT3 #(
		.INIT('h96)
	) name6335 (
		_w6398_,
		_w6399_,
		_w6400_,
		_w6401_
	);
	LUT3 #(
		.INIT('h0d)
	) name6336 (
		_w6267_,
		_w6275_,
		_w6276_,
		_w6402_
	);
	LUT4 #(
		.INIT('h153f)
	) name6337 (
		\a[18] ,
		\a[19] ,
		\a[61] ,
		\a[62] ,
		_w6403_
	);
	LUT4 #(
		.INIT('h000d)
	) name6338 (
		_w6207_,
		_w6208_,
		_w6210_,
		_w6265_,
		_w6404_
	);
	LUT3 #(
		.INIT('h0d)
	) name6339 (
		_w6271_,
		_w6272_,
		_w6273_,
		_w6405_
	);
	LUT2 #(
		.INIT('h8)
	) name6340 (
		\a[30] ,
		\a[51] ,
		_w6406_
	);
	LUT4 #(
		.INIT('h153f)
	) name6341 (
		\a[31] ,
		\a[32] ,
		\a[49] ,
		\a[50] ,
		_w6407_
	);
	LUT2 #(
		.INIT('h8)
	) name6342 (
		\a[32] ,
		\a[50] ,
		_w6408_
	);
	LUT4 #(
		.INIT('h8000)
	) name6343 (
		\a[31] ,
		\a[32] ,
		\a[49] ,
		\a[50] ,
		_w6409_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6344 (
		\a[31] ,
		\a[32] ,
		\a[49] ,
		\a[50] ,
		_w6410_
	);
	LUT2 #(
		.INIT('h6)
	) name6345 (
		_w6406_,
		_w6410_,
		_w6411_
	);
	LUT4 #(
		.INIT('he11e)
	) name6346 (
		_w6403_,
		_w6404_,
		_w6405_,
		_w6411_,
		_w6412_
	);
	LUT3 #(
		.INIT('h69)
	) name6347 (
		_w6401_,
		_w6402_,
		_w6412_,
		_w6413_
	);
	LUT3 #(
		.INIT('h0d)
	) name6348 (
		_w6296_,
		_w6297_,
		_w6298_,
		_w6414_
	);
	LUT3 #(
		.INIT('h0d)
	) name6349 (
		_w6201_,
		_w6303_,
		_w6304_,
		_w6415_
	);
	LUT3 #(
		.INIT('h0d)
	) name6350 (
		_w6291_,
		_w6292_,
		_w6294_,
		_w6416_
	);
	LUT3 #(
		.INIT('h96)
	) name6351 (
		_w6414_,
		_w6415_,
		_w6416_,
		_w6417_
	);
	LUT3 #(
		.INIT('hb2)
	) name6352 (
		_w6284_,
		_w6285_,
		_w6289_,
		_w6418_
	);
	LUT3 #(
		.INIT('h32)
	) name6353 (
		_w6300_,
		_w6301_,
		_w6306_,
		_w6419_
	);
	LUT3 #(
		.INIT('h69)
	) name6354 (
		_w6417_,
		_w6418_,
		_w6419_,
		_w6420_
	);
	LUT3 #(
		.INIT('h60)
	) name6355 (
		_w6397_,
		_w6413_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h1)
	) name6356 (
		_w6264_,
		_w6309_,
		_w6422_
	);
	LUT3 #(
		.INIT('h54)
	) name6357 (
		_w6321_,
		_w6322_,
		_w6324_,
		_w6423_
	);
	LUT3 #(
		.INIT('h17)
	) name6358 (
		_w6317_,
		_w6318_,
		_w6319_,
		_w6424_
	);
	LUT2 #(
		.INIT('h8)
	) name6359 (
		\a[27] ,
		\a[54] ,
		_w6425_
	);
	LUT4 #(
		.INIT('h153f)
	) name6360 (
		\a[38] ,
		\a[39] ,
		\a[42] ,
		\a[43] ,
		_w6426_
	);
	LUT4 #(
		.INIT('h8000)
	) name6361 (
		\a[38] ,
		\a[39] ,
		\a[42] ,
		\a[43] ,
		_w6427_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6362 (
		\a[38] ,
		\a[39] ,
		\a[42] ,
		\a[43] ,
		_w6428_
	);
	LUT2 #(
		.INIT('h6)
	) name6363 (
		_w6425_,
		_w6428_,
		_w6429_
	);
	LUT4 #(
		.INIT('h1700)
	) name6364 (
		_w6328_,
		_w6329_,
		_w6330_,
		_w6429_,
		_w6430_
	);
	LUT4 #(
		.INIT('h00e8)
	) name6365 (
		_w6328_,
		_w6329_,
		_w6330_,
		_w6429_,
		_w6431_
	);
	LUT3 #(
		.INIT('ha9)
	) name6366 (
		_w6424_,
		_w6430_,
		_w6431_,
		_w6432_
	);
	LUT3 #(
		.INIT('hd4)
	) name6367 (
		_w6331_,
		_w6332_,
		_w6333_,
		_w6433_
	);
	LUT3 #(
		.INIT('h96)
	) name6368 (
		_w6423_,
		_w6432_,
		_w6433_,
		_w6434_
	);
	LUT4 #(
		.INIT('h0e00)
	) name6369 (
		_w6264_,
		_w6309_,
		_w6311_,
		_w6434_,
		_w6435_
	);
	LUT3 #(
		.INIT('h09)
	) name6370 (
		_w6397_,
		_w6413_,
		_w6420_,
		_w6436_
	);
	LUT4 #(
		.INIT('h0096)
	) name6371 (
		_w6423_,
		_w6432_,
		_w6433_,
		_w6436_,
		_w6437_
	);
	LUT4 #(
		.INIT('h002f)
	) name6372 (
		_w6243_,
		_w6245_,
		_w6310_,
		_w6436_,
		_w6438_
	);
	LUT4 #(
		.INIT('h010f)
	) name6373 (
		_w6264_,
		_w6309_,
		_w6437_,
		_w6438_,
		_w6439_
	);
	LUT3 #(
		.INIT('h01)
	) name6374 (
		_w6421_,
		_w6435_,
		_w6439_,
		_w6440_
	);
	LUT3 #(
		.INIT('h96)
	) name6375 (
		_w6397_,
		_w6413_,
		_w6420_,
		_w6441_
	);
	LUT3 #(
		.INIT('h04)
	) name6376 (
		_w6311_,
		_w6434_,
		_w6441_,
		_w6442_
	);
	LUT4 #(
		.INIT('h0069)
	) name6377 (
		_w6423_,
		_w6432_,
		_w6433_,
		_w6441_,
		_w6443_
	);
	LUT4 #(
		.INIT('hf100)
	) name6378 (
		_w6264_,
		_w6309_,
		_w6311_,
		_w6443_,
		_w6444_
	);
	LUT3 #(
		.INIT('h0b)
	) name6379 (
		_w6422_,
		_w6442_,
		_w6444_,
		_w6445_
	);
	LUT3 #(
		.INIT('h9a)
	) name6380 (
		_w6396_,
		_w6440_,
		_w6445_,
		_w6446_
	);
	LUT2 #(
		.INIT('h4)
	) name6381 (
		_w6355_,
		_w6446_,
		_w6447_
	);
	LUT2 #(
		.INIT('h2)
	) name6382 (
		_w6355_,
		_w6446_,
		_w6448_
	);
	LUT2 #(
		.INIT('h9)
	) name6383 (
		_w6355_,
		_w6446_,
		_w6449_
	);
	LUT3 #(
		.INIT('h1e)
	) name6384 (
		_w6346_,
		_w6354_,
		_w6449_,
		_w6450_
	);
	LUT2 #(
		.INIT('h1)
	) name6385 (
		_w6346_,
		_w6447_,
		_w6451_
	);
	LUT4 #(
		.INIT('h2322)
	) name6386 (
		_w6394_,
		_w6395_,
		_w6440_,
		_w6445_,
		_w6452_
	);
	LUT3 #(
		.INIT('he8)
	) name6387 (
		_w6397_,
		_w6413_,
		_w6420_,
		_w6453_
	);
	LUT3 #(
		.INIT('h0e)
	) name6388 (
		_w6424_,
		_w6430_,
		_w6431_,
		_w6454_
	);
	LUT4 #(
		.INIT('h153f)
	) name6389 (
		\a[33] ,
		\a[34] ,
		\a[48] ,
		\a[49] ,
		_w6455_
	);
	LUT4 #(
		.INIT('h8000)
	) name6390 (
		\a[33] ,
		\a[34] ,
		\a[48] ,
		\a[49] ,
		_w6456_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6391 (
		\a[33] ,
		\a[34] ,
		\a[48] ,
		\a[49] ,
		_w6457_
	);
	LUT2 #(
		.INIT('h8)
	) name6392 (
		\a[20] ,
		\a[62] ,
		_w6458_
	);
	LUT4 #(
		.INIT('h153f)
	) name6393 (
		\a[21] ,
		\a[31] ,
		\a[51] ,
		\a[61] ,
		_w6459_
	);
	LUT4 #(
		.INIT('h8000)
	) name6394 (
		\a[21] ,
		\a[31] ,
		\a[51] ,
		\a[61] ,
		_w6460_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6395 (
		\a[21] ,
		\a[31] ,
		\a[51] ,
		\a[61] ,
		_w6461_
	);
	LUT4 #(
		.INIT('h0660)
	) name6396 (
		_w6408_,
		_w6457_,
		_w6458_,
		_w6461_,
		_w6462_
	);
	LUT4 #(
		.INIT('h9009)
	) name6397 (
		_w6408_,
		_w6457_,
		_w6458_,
		_w6461_,
		_w6463_
	);
	LUT4 #(
		.INIT('h6996)
	) name6398 (
		_w6408_,
		_w6457_,
		_w6458_,
		_w6461_,
		_w6464_
	);
	LUT2 #(
		.INIT('h8)
	) name6399 (
		\a[22] ,
		\a[60] ,
		_w6465_
	);
	LUT4 #(
		.INIT('h153f)
	) name6400 (
		\a[23] ,
		\a[24] ,
		\a[58] ,
		\a[59] ,
		_w6466_
	);
	LUT4 #(
		.INIT('h8000)
	) name6401 (
		\a[23] ,
		\a[24] ,
		\a[58] ,
		\a[59] ,
		_w6467_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6402 (
		\a[23] ,
		\a[24] ,
		\a[58] ,
		\a[59] ,
		_w6468_
	);
	LUT2 #(
		.INIT('h6)
	) name6403 (
		_w6465_,
		_w6468_,
		_w6469_
	);
	LUT2 #(
		.INIT('h6)
	) name6404 (
		_w6464_,
		_w6469_,
		_w6470_
	);
	LUT4 #(
		.INIT('h153f)
	) name6405 (
		\a[38] ,
		\a[39] ,
		\a[43] ,
		\a[44] ,
		_w6471_
	);
	LUT4 #(
		.INIT('h8000)
	) name6406 (
		\a[38] ,
		\a[39] ,
		\a[43] ,
		\a[44] ,
		_w6472_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6407 (
		\a[38] ,
		\a[39] ,
		\a[43] ,
		\a[44] ,
		_w6473_
	);
	LUT2 #(
		.INIT('h8)
	) name6408 (
		\a[40] ,
		\a[42] ,
		_w6474_
	);
	LUT4 #(
		.INIT('h153f)
	) name6409 (
		\a[29] ,
		\a[30] ,
		\a[52] ,
		\a[53] ,
		_w6475_
	);
	LUT4 #(
		.INIT('h8000)
	) name6410 (
		\a[29] ,
		\a[30] ,
		\a[52] ,
		\a[53] ,
		_w6476_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6411 (
		\a[29] ,
		\a[30] ,
		\a[52] ,
		\a[53] ,
		_w6477_
	);
	LUT4 #(
		.INIT('h0660)
	) name6412 (
		_w6293_,
		_w6473_,
		_w6474_,
		_w6477_,
		_w6478_
	);
	LUT4 #(
		.INIT('h9009)
	) name6413 (
		_w6293_,
		_w6473_,
		_w6474_,
		_w6477_,
		_w6479_
	);
	LUT4 #(
		.INIT('h6996)
	) name6414 (
		_w6293_,
		_w6473_,
		_w6474_,
		_w6477_,
		_w6480_
	);
	LUT2 #(
		.INIT('h8)
	) name6415 (
		\a[35] ,
		\a[47] ,
		_w6481_
	);
	LUT4 #(
		.INIT('h153f)
	) name6416 (
		\a[36] ,
		\a[37] ,
		\a[45] ,
		\a[46] ,
		_w6482_
	);
	LUT4 #(
		.INIT('h8000)
	) name6417 (
		\a[36] ,
		\a[37] ,
		\a[45] ,
		\a[46] ,
		_w6483_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6418 (
		\a[36] ,
		\a[37] ,
		\a[45] ,
		\a[46] ,
		_w6484_
	);
	LUT2 #(
		.INIT('h6)
	) name6419 (
		_w6481_,
		_w6484_,
		_w6485_
	);
	LUT2 #(
		.INIT('h6)
	) name6420 (
		_w6480_,
		_w6485_,
		_w6486_
	);
	LUT4 #(
		.INIT('h9009)
	) name6421 (
		_w6464_,
		_w6469_,
		_w6480_,
		_w6485_,
		_w6487_
	);
	LUT3 #(
		.INIT('h96)
	) name6422 (
		_w6454_,
		_w6470_,
		_w6486_,
		_w6488_
	);
	LUT4 #(
		.INIT('he800)
	) name6423 (
		_w6423_,
		_w6432_,
		_w6433_,
		_w6488_,
		_w6489_
	);
	LUT4 #(
		.INIT('h0017)
	) name6424 (
		_w6423_,
		_w6432_,
		_w6433_,
		_w6488_,
		_w6490_
	);
	LUT3 #(
		.INIT('ha9)
	) name6425 (
		_w6453_,
		_w6489_,
		_w6490_,
		_w6491_
	);
	LUT4 #(
		.INIT('hcd00)
	) name6426 (
		_w6421_,
		_w6435_,
		_w6439_,
		_w6491_,
		_w6492_
	);
	LUT4 #(
		.INIT('h0032)
	) name6427 (
		_w6421_,
		_w6435_,
		_w6439_,
		_w6491_,
		_w6493_
	);
	LUT4 #(
		.INIT('h32cd)
	) name6428 (
		_w6421_,
		_w6435_,
		_w6439_,
		_w6491_,
		_w6494_
	);
	LUT2 #(
		.INIT('h1)
	) name6429 (
		_w6357_,
		_w6390_,
		_w6495_
	);
	LUT3 #(
		.INIT('h17)
	) name6430 (
		_w6414_,
		_w6415_,
		_w6416_,
		_w6496_
	);
	LUT4 #(
		.INIT('h153f)
	) name6431 (
		\a[25] ,
		\a[27] ,
		\a[55] ,
		\a[57] ,
		_w6497_
	);
	LUT4 #(
		.INIT('h8000)
	) name6432 (
		\a[25] ,
		\a[27] ,
		\a[55] ,
		\a[57] ,
		_w6498_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6433 (
		\a[25] ,
		\a[27] ,
		\a[55] ,
		\a[57] ,
		_w6499_
	);
	LUT2 #(
		.INIT('h6)
	) name6434 (
		_w3231_,
		_w6499_,
		_w6500_
	);
	LUT4 #(
		.INIT('h1700)
	) name6435 (
		_w6398_,
		_w6399_,
		_w6400_,
		_w6500_,
		_w6501_
	);
	LUT4 #(
		.INIT('h00e8)
	) name6436 (
		_w6398_,
		_w6399_,
		_w6400_,
		_w6500_,
		_w6502_
	);
	LUT3 #(
		.INIT('ha9)
	) name6437 (
		_w6496_,
		_w6501_,
		_w6502_,
		_w6503_
	);
	LUT3 #(
		.INIT('hd4)
	) name6438 (
		_w6417_,
		_w6418_,
		_w6419_,
		_w6504_
	);
	LUT3 #(
		.INIT('hd4)
	) name6439 (
		_w6401_,
		_w6402_,
		_w6412_,
		_w6505_
	);
	LUT3 #(
		.INIT('h96)
	) name6440 (
		_w6503_,
		_w6504_,
		_w6505_,
		_w6506_
	);
	LUT4 #(
		.INIT('h00f1)
	) name6441 (
		_w6357_,
		_w6390_,
		_w6391_,
		_w6506_,
		_w6507_
	);
	LUT3 #(
		.INIT('h17)
	) name6442 (
		_w6358_,
		_w6371_,
		_w6388_,
		_w6508_
	);
	LUT3 #(
		.INIT('h0d)
	) name6443 (
		_w4607_,
		_w6367_,
		_w6368_,
		_w6509_
	);
	LUT3 #(
		.INIT('h0d)
	) name6444 (
		_w6406_,
		_w6407_,
		_w6409_,
		_w6510_
	);
	LUT3 #(
		.INIT('h0d)
	) name6445 (
		_w6383_,
		_w6384_,
		_w6385_,
		_w6511_
	);
	LUT3 #(
		.INIT('h96)
	) name6446 (
		_w6509_,
		_w6510_,
		_w6511_,
		_w6512_
	);
	LUT3 #(
		.INIT('h0d)
	) name6447 (
		_w6280_,
		_w6359_,
		_w6361_,
		_w6513_
	);
	LUT3 #(
		.INIT('h0d)
	) name6448 (
		_w6372_,
		_w6373_,
		_w6374_,
		_w6514_
	);
	LUT3 #(
		.INIT('h0d)
	) name6449 (
		_w6376_,
		_w6377_,
		_w6378_,
		_w6515_
	);
	LUT3 #(
		.INIT('h96)
	) name6450 (
		_w6513_,
		_w6514_,
		_w6515_,
		_w6516_
	);
	LUT3 #(
		.INIT('h32)
	) name6451 (
		_w6380_,
		_w6381_,
		_w6387_,
		_w6517_
	);
	LUT3 #(
		.INIT('h96)
	) name6452 (
		_w6512_,
		_w6516_,
		_w6517_,
		_w6518_
	);
	LUT3 #(
		.INIT('h32)
	) name6453 (
		_w6364_,
		_w6365_,
		_w6370_,
		_w6519_
	);
	LUT4 #(
		.INIT('h1f01)
	) name6454 (
		_w6403_,
		_w6404_,
		_w6405_,
		_w6411_,
		_w6520_
	);
	LUT3 #(
		.INIT('h13)
	) name6455 (
		\a[19] ,
		\a[40] ,
		\a[62] ,
		_w6521_
	);
	LUT3 #(
		.INIT('h80)
	) name6456 (
		\a[19] ,
		\a[41] ,
		\a[63] ,
		_w6522_
	);
	LUT2 #(
		.INIT('h4)
	) name6457 (
		_w6521_,
		_w6522_,
		_w6523_
	);
	LUT4 #(
		.INIT('he0c0)
	) name6458 (
		\a[19] ,
		\a[40] ,
		\a[41] ,
		\a[62] ,
		_w6524_
	);
	LUT2 #(
		.INIT('h1)
	) name6459 (
		_w5745_,
		_w6524_,
		_w6525_
	);
	LUT3 #(
		.INIT('hc6)
	) name6460 (
		\a[41] ,
		_w5745_,
		_w6521_,
		_w6526_
	);
	LUT3 #(
		.INIT('h0d)
	) name6461 (
		_w6425_,
		_w6426_,
		_w6427_,
		_w6527_
	);
	LUT2 #(
		.INIT('h6)
	) name6462 (
		_w6526_,
		_w6527_,
		_w6528_
	);
	LUT3 #(
		.INIT('h69)
	) name6463 (
		_w6519_,
		_w6520_,
		_w6528_,
		_w6529_
	);
	LUT3 #(
		.INIT('h69)
	) name6464 (
		_w6508_,
		_w6518_,
		_w6529_,
		_w6530_
	);
	LUT4 #(
		.INIT('h0e00)
	) name6465 (
		_w6357_,
		_w6390_,
		_w6391_,
		_w6506_,
		_w6531_
	);
	LUT3 #(
		.INIT('h04)
	) name6466 (
		_w6507_,
		_w6530_,
		_w6531_,
		_w6532_
	);
	LUT3 #(
		.INIT('h04)
	) name6467 (
		_w6391_,
		_w6506_,
		_w6530_,
		_w6533_
	);
	LUT4 #(
		.INIT('h4114)
	) name6468 (
		_w6506_,
		_w6508_,
		_w6518_,
		_w6529_,
		_w6534_
	);
	LUT4 #(
		.INIT('hf100)
	) name6469 (
		_w6357_,
		_w6390_,
		_w6391_,
		_w6534_,
		_w6535_
	);
	LUT3 #(
		.INIT('h0b)
	) name6470 (
		_w6495_,
		_w6533_,
		_w6535_,
		_w6536_
	);
	LUT3 #(
		.INIT('h45)
	) name6471 (
		_w6494_,
		_w6532_,
		_w6536_,
		_w6537_
	);
	LUT4 #(
		.INIT('h0100)
	) name6472 (
		_w6492_,
		_w6493_,
		_w6532_,
		_w6536_,
		_w6538_
	);
	LUT4 #(
		.INIT('h1e11)
	) name6473 (
		_w6492_,
		_w6493_,
		_w6532_,
		_w6536_,
		_w6539_
	);
	LUT2 #(
		.INIT('h1)
	) name6474 (
		_w6452_,
		_w6539_,
		_w6540_
	);
	LUT3 #(
		.INIT('h02)
	) name6475 (
		_w6452_,
		_w6537_,
		_w6538_,
		_w6541_
	);
	LUT3 #(
		.INIT('h01)
	) name6476 (
		_w6448_,
		_w6540_,
		_w6541_,
		_w6542_
	);
	LUT3 #(
		.INIT('hb0)
	) name6477 (
		_w6354_,
		_w6451_,
		_w6542_,
		_w6543_
	);
	LUT3 #(
		.INIT('ha9)
	) name6478 (
		_w6452_,
		_w6537_,
		_w6538_,
		_w6544_
	);
	LUT2 #(
		.INIT('h2)
	) name6479 (
		_w6448_,
		_w6544_,
		_w6545_
	);
	LUT4 #(
		.INIT('h00fb)
	) name6480 (
		_w6354_,
		_w6451_,
		_w6544_,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('h4)
	) name6481 (
		_w6543_,
		_w6546_,
		_w6547_
	);
	LUT4 #(
		.INIT('h5455)
	) name6482 (
		_w6492_,
		_w6493_,
		_w6532_,
		_w6536_,
		_w6548_
	);
	LUT4 #(
		.INIT('hf110)
	) name6483 (
		_w6391_,
		_w6495_,
		_w6506_,
		_w6530_,
		_w6549_
	);
	LUT3 #(
		.INIT('h2b)
	) name6484 (
		_w6508_,
		_w6518_,
		_w6529_,
		_w6550_
	);
	LUT3 #(
		.INIT('he8)
	) name6485 (
		_w6503_,
		_w6504_,
		_w6505_,
		_w6551_
	);
	LUT3 #(
		.INIT('h0e)
	) name6486 (
		_w6496_,
		_w6501_,
		_w6502_,
		_w6552_
	);
	LUT2 #(
		.INIT('h8)
	) name6487 (
		\a[29] ,
		\a[54] ,
		_w6553_
	);
	LUT4 #(
		.INIT('h153f)
	) name6488 (
		\a[39] ,
		\a[40] ,
		\a[43] ,
		\a[44] ,
		_w6554_
	);
	LUT4 #(
		.INIT('h8000)
	) name6489 (
		\a[39] ,
		\a[40] ,
		\a[43] ,
		\a[44] ,
		_w6555_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6490 (
		\a[39] ,
		\a[40] ,
		\a[43] ,
		\a[44] ,
		_w6556_
	);
	LUT4 #(
		.INIT('h9a30)
	) name6491 (
		\a[21] ,
		\a[41] ,
		\a[42] ,
		\a[62] ,
		_w6557_
	);
	LUT3 #(
		.INIT('h60)
	) name6492 (
		_w6553_,
		_w6556_,
		_w6557_,
		_w6558_
	);
	LUT3 #(
		.INIT('h09)
	) name6493 (
		_w6553_,
		_w6556_,
		_w6557_,
		_w6559_
	);
	LUT3 #(
		.INIT('h96)
	) name6494 (
		_w6553_,
		_w6556_,
		_w6557_,
		_w6560_
	);
	LUT2 #(
		.INIT('h8)
	) name6495 (
		\a[33] ,
		\a[50] ,
		_w6561_
	);
	LUT4 #(
		.INIT('h153f)
	) name6496 (
		\a[34] ,
		\a[35] ,
		\a[48] ,
		\a[49] ,
		_w6562_
	);
	LUT4 #(
		.INIT('h8000)
	) name6497 (
		\a[34] ,
		\a[35] ,
		\a[48] ,
		\a[49] ,
		_w6563_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6498 (
		\a[34] ,
		\a[35] ,
		\a[48] ,
		\a[49] ,
		_w6564_
	);
	LUT2 #(
		.INIT('h6)
	) name6499 (
		_w6561_,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h6)
	) name6500 (
		_w6560_,
		_w6565_,
		_w6566_
	);
	LUT4 #(
		.INIT('h153f)
	) name6501 (
		\a[26] ,
		\a[32] ,
		\a[51] ,
		\a[57] ,
		_w6567_
	);
	LUT4 #(
		.INIT('h8000)
	) name6502 (
		\a[26] ,
		\a[32] ,
		\a[51] ,
		\a[57] ,
		_w6568_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6503 (
		\a[26] ,
		\a[32] ,
		\a[51] ,
		\a[57] ,
		_w6569_
	);
	LUT2 #(
		.INIT('h8)
	) name6504 (
		\a[36] ,
		\a[47] ,
		_w6570_
	);
	LUT4 #(
		.INIT('h153f)
	) name6505 (
		\a[37] ,
		\a[38] ,
		\a[45] ,
		\a[46] ,
		_w6571_
	);
	LUT4 #(
		.INIT('h8000)
	) name6506 (
		\a[37] ,
		\a[38] ,
		\a[45] ,
		\a[46] ,
		_w6572_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6507 (
		\a[37] ,
		\a[38] ,
		\a[45] ,
		\a[46] ,
		_w6573_
	);
	LUT4 #(
		.INIT('h0660)
	) name6508 (
		_w6360_,
		_w6569_,
		_w6570_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h9009)
	) name6509 (
		_w6360_,
		_w6569_,
		_w6570_,
		_w6573_,
		_w6575_
	);
	LUT4 #(
		.INIT('h6996)
	) name6510 (
		_w6360_,
		_w6569_,
		_w6570_,
		_w6573_,
		_w6576_
	);
	LUT4 #(
		.INIT('h153f)
	) name6511 (
		\a[20] ,
		\a[22] ,
		\a[61] ,
		\a[63] ,
		_w6577_
	);
	LUT4 #(
		.INIT('h8000)
	) name6512 (
		\a[20] ,
		\a[22] ,
		\a[61] ,
		\a[63] ,
		_w6578_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6513 (
		\a[20] ,
		\a[22] ,
		\a[61] ,
		\a[63] ,
		_w6579_
	);
	LUT2 #(
		.INIT('h6)
	) name6514 (
		_w6164_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h6)
	) name6515 (
		_w6576_,
		_w6580_,
		_w6581_
	);
	LUT4 #(
		.INIT('h9009)
	) name6516 (
		_w6560_,
		_w6565_,
		_w6576_,
		_w6580_,
		_w6582_
	);
	LUT3 #(
		.INIT('h96)
	) name6517 (
		_w6552_,
		_w6566_,
		_w6581_,
		_w6583_
	);
	LUT2 #(
		.INIT('h8)
	) name6518 (
		_w6551_,
		_w6583_,
		_w6584_
	);
	LUT2 #(
		.INIT('h1)
	) name6519 (
		_w6551_,
		_w6583_,
		_w6585_
	);
	LUT2 #(
		.INIT('h6)
	) name6520 (
		_w6551_,
		_w6583_,
		_w6586_
	);
	LUT2 #(
		.INIT('h9)
	) name6521 (
		_w6550_,
		_w6586_,
		_w6587_
	);
	LUT3 #(
		.INIT('h31)
	) name6522 (
		_w6453_,
		_w6489_,
		_w6490_,
		_w6588_
	);
	LUT3 #(
		.INIT('h17)
	) name6523 (
		_w6509_,
		_w6510_,
		_w6511_,
		_w6589_
	);
	LUT3 #(
		.INIT('h17)
	) name6524 (
		_w6513_,
		_w6514_,
		_w6515_,
		_w6590_
	);
	LUT3 #(
		.INIT('h32)
	) name6525 (
		_w6462_,
		_w6463_,
		_w6469_,
		_w6591_
	);
	LUT3 #(
		.INIT('h96)
	) name6526 (
		_w6589_,
		_w6590_,
		_w6591_,
		_w6592_
	);
	LUT3 #(
		.INIT('h23)
	) name6527 (
		_w6523_,
		_w6525_,
		_w6527_,
		_w6593_
	);
	LUT4 #(
		.INIT('h8000)
	) name6528 (
		\a[23] ,
		\a[24] ,
		\a[59] ,
		\a[60] ,
		_w6594_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6529 (
		\a[23] ,
		\a[24] ,
		\a[59] ,
		\a[60] ,
		_w6595_
	);
	LUT4 #(
		.INIT('hf20d)
	) name6530 (
		_w6474_,
		_w6475_,
		_w6476_,
		_w6595_,
		_w6596_
	);
	LUT2 #(
		.INIT('h8)
	) name6531 (
		\a[31] ,
		\a[52] ,
		_w6597_
	);
	LUT4 #(
		.INIT('h153f)
	) name6532 (
		\a[28] ,
		\a[30] ,
		\a[53] ,
		\a[55] ,
		_w6598_
	);
	LUT4 #(
		.INIT('h8000)
	) name6533 (
		\a[28] ,
		\a[30] ,
		\a[53] ,
		\a[55] ,
		_w6599_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6534 (
		\a[28] ,
		\a[30] ,
		\a[53] ,
		\a[55] ,
		_w6600_
	);
	LUT2 #(
		.INIT('h6)
	) name6535 (
		_w6597_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h4)
	) name6536 (
		_w6596_,
		_w6601_,
		_w6602_
	);
	LUT2 #(
		.INIT('h2)
	) name6537 (
		_w6596_,
		_w6601_,
		_w6603_
	);
	LUT2 #(
		.INIT('h9)
	) name6538 (
		_w6596_,
		_w6601_,
		_w6604_
	);
	LUT2 #(
		.INIT('h6)
	) name6539 (
		_w6593_,
		_w6604_,
		_w6605_
	);
	LUT3 #(
		.INIT('h8e)
	) name6540 (
		_w6519_,
		_w6520_,
		_w6528_,
		_w6606_
	);
	LUT3 #(
		.INIT('h96)
	) name6541 (
		_w6592_,
		_w6605_,
		_w6606_,
		_w6607_
	);
	LUT3 #(
		.INIT('h0d)
	) name6542 (
		_w6465_,
		_w6466_,
		_w6467_,
		_w6608_
	);
	LUT3 #(
		.INIT('h0d)
	) name6543 (
		_w6481_,
		_w6482_,
		_w6483_,
		_w6609_
	);
	LUT3 #(
		.INIT('h0d)
	) name6544 (
		_w6293_,
		_w6471_,
		_w6472_,
		_w6610_
	);
	LUT3 #(
		.INIT('h96)
	) name6545 (
		_w6608_,
		_w6609_,
		_w6610_,
		_w6611_
	);
	LUT3 #(
		.INIT('h32)
	) name6546 (
		_w6458_,
		_w6459_,
		_w6460_,
		_w6612_
	);
	LUT3 #(
		.INIT('h0d)
	) name6547 (
		_w6408_,
		_w6455_,
		_w6456_,
		_w6613_
	);
	LUT3 #(
		.INIT('h0d)
	) name6548 (
		_w3231_,
		_w6497_,
		_w6498_,
		_w6614_
	);
	LUT3 #(
		.INIT('h69)
	) name6549 (
		_w6612_,
		_w6613_,
		_w6614_,
		_w6615_
	);
	LUT3 #(
		.INIT('h32)
	) name6550 (
		_w6478_,
		_w6479_,
		_w6485_,
		_w6616_
	);
	LUT3 #(
		.INIT('h96)
	) name6551 (
		_w6611_,
		_w6615_,
		_w6616_,
		_w6617_
	);
	LUT4 #(
		.INIT('h00f1)
	) name6552 (
		_w6424_,
		_w6430_,
		_w6431_,
		_w6470_,
		_w6618_
	);
	LUT4 #(
		.INIT('h00f1)
	) name6553 (
		_w6424_,
		_w6430_,
		_w6431_,
		_w6486_,
		_w6619_
	);
	LUT3 #(
		.INIT('h01)
	) name6554 (
		_w6487_,
		_w6618_,
		_w6619_,
		_w6620_
	);
	LUT3 #(
		.INIT('h71)
	) name6555 (
		_w6512_,
		_w6516_,
		_w6517_,
		_w6621_
	);
	LUT4 #(
		.INIT('he800)
	) name6556 (
		_w6454_,
		_w6470_,
		_w6486_,
		_w6621_,
		_w6622_
	);
	LUT3 #(
		.INIT('h96)
	) name6557 (
		_w6617_,
		_w6620_,
		_w6621_,
		_w6623_
	);
	LUT3 #(
		.INIT('h96)
	) name6558 (
		_w6588_,
		_w6607_,
		_w6623_,
		_w6624_
	);
	LUT3 #(
		.INIT('h69)
	) name6559 (
		_w6549_,
		_w6587_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h4)
	) name6560 (
		_w6548_,
		_w6625_,
		_w6626_
	);
	LUT2 #(
		.INIT('h2)
	) name6561 (
		_w6548_,
		_w6625_,
		_w6627_
	);
	LUT2 #(
		.INIT('h9)
	) name6562 (
		_w6548_,
		_w6625_,
		_w6628_
	);
	LUT3 #(
		.INIT('h01)
	) name6563 (
		_w6346_,
		_w6447_,
		_w6541_,
		_w6629_
	);
	LUT3 #(
		.INIT('h31)
	) name6564 (
		_w6448_,
		_w6540_,
		_w6541_,
		_w6630_
	);
	LUT4 #(
		.INIT('h63cc)
	) name6565 (
		_w6354_,
		_w6628_,
		_w6629_,
		_w6630_,
		_w6631_
	);
	LUT4 #(
		.INIT('h0031)
	) name6566 (
		_w6448_,
		_w6540_,
		_w6541_,
		_w6627_,
		_w6632_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6567 (
		_w6487_,
		_w6618_,
		_w6619_,
		_w6621_,
		_w6633_
	);
	LUT3 #(
		.INIT('h0e)
	) name6568 (
		_w6617_,
		_w6622_,
		_w6633_,
		_w6634_
	);
	LUT4 #(
		.INIT('h002b)
	) name6569 (
		_w6550_,
		_w6551_,
		_w6583_,
		_w6634_,
		_w6635_
	);
	LUT4 #(
		.INIT('he0c0)
	) name6570 (
		\a[21] ,
		\a[41] ,
		\a[42] ,
		\a[62] ,
		_w6636_
	);
	LUT4 #(
		.INIT('h000d)
	) name6571 (
		_w6553_,
		_w6554_,
		_w6555_,
		_w6636_,
		_w6637_
	);
	LUT4 #(
		.INIT('hf200)
	) name6572 (
		_w6553_,
		_w6554_,
		_w6555_,
		_w6636_,
		_w6638_
	);
	LUT4 #(
		.INIT('h0df2)
	) name6573 (
		_w6553_,
		_w6554_,
		_w6555_,
		_w6636_,
		_w6639_
	);
	LUT3 #(
		.INIT('h0d)
	) name6574 (
		_w6597_,
		_w6598_,
		_w6599_,
		_w6640_
	);
	LUT2 #(
		.INIT('h6)
	) name6575 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT3 #(
		.INIT('h32)
	) name6576 (
		_w6574_,
		_w6575_,
		_w6580_,
		_w6642_
	);
	LUT3 #(
		.INIT('h32)
	) name6577 (
		_w6558_,
		_w6559_,
		_w6565_,
		_w6643_
	);
	LUT3 #(
		.INIT('h69)
	) name6578 (
		_w6641_,
		_w6642_,
		_w6643_,
		_w6644_
	);
	LUT4 #(
		.INIT('h00f1)
	) name6579 (
		_w6496_,
		_w6501_,
		_w6502_,
		_w6566_,
		_w6645_
	);
	LUT4 #(
		.INIT('h00f1)
	) name6580 (
		_w6496_,
		_w6501_,
		_w6502_,
		_w6581_,
		_w6646_
	);
	LUT3 #(
		.INIT('h01)
	) name6581 (
		_w6582_,
		_w6645_,
		_w6646_,
		_w6647_
	);
	LUT3 #(
		.INIT('h71)
	) name6582 (
		_w6611_,
		_w6615_,
		_w6616_,
		_w6648_
	);
	LUT4 #(
		.INIT('he800)
	) name6583 (
		_w6552_,
		_w6566_,
		_w6581_,
		_w6648_,
		_w6649_
	);
	LUT3 #(
		.INIT('h96)
	) name6584 (
		_w6644_,
		_w6647_,
		_w6648_,
		_w6650_
	);
	LUT2 #(
		.INIT('h4)
	) name6585 (
		_w6634_,
		_w6650_,
		_w6651_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6586 (
		_w6550_,
		_w6551_,
		_w6583_,
		_w6650_,
		_w6652_
	);
	LUT3 #(
		.INIT('h54)
	) name6587 (
		_w6635_,
		_w6651_,
		_w6652_,
		_w6653_
	);
	LUT3 #(
		.INIT('h32)
	) name6588 (
		_w6550_,
		_w6584_,
		_w6585_,
		_w6654_
	);
	LUT3 #(
		.INIT('hed)
	) name6589 (
		_w6634_,
		_w6650_,
		_w6654_,
		_w6655_
	);
	LUT4 #(
		.INIT('hce00)
	) name6590 (
		_w6453_,
		_w6489_,
		_w6490_,
		_w6607_,
		_w6656_
	);
	LUT4 #(
		.INIT('h0031)
	) name6591 (
		_w6453_,
		_w6489_,
		_w6490_,
		_w6607_,
		_w6657_
	);
	LUT3 #(
		.INIT('he8)
	) name6592 (
		_w6592_,
		_w6605_,
		_w6606_,
		_w6658_
	);
	LUT3 #(
		.INIT('h0e)
	) name6593 (
		_w6593_,
		_w6602_,
		_w6603_,
		_w6659_
	);
	LUT4 #(
		.INIT('h153f)
	) name6594 (
		\a[23] ,
		\a[24] ,
		\a[59] ,
		\a[60] ,
		_w6660_
	);
	LUT4 #(
		.INIT('h000d)
	) name6595 (
		_w6474_,
		_w6475_,
		_w6476_,
		_w6594_,
		_w6661_
	);
	LUT3 #(
		.INIT('h0d)
	) name6596 (
		_w6164_,
		_w6577_,
		_w6578_,
		_w6662_
	);
	LUT2 #(
		.INIT('h8)
	) name6597 (
		\a[26] ,
		\a[58] ,
		_w6663_
	);
	LUT4 #(
		.INIT('h153f)
	) name6598 (
		\a[31] ,
		\a[32] ,
		\a[52] ,
		\a[53] ,
		_w6664_
	);
	LUT2 #(
		.INIT('h8)
	) name6599 (
		\a[32] ,
		\a[53] ,
		_w6665_
	);
	LUT4 #(
		.INIT('h8000)
	) name6600 (
		\a[31] ,
		\a[32] ,
		\a[52] ,
		\a[53] ,
		_w6666_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6601 (
		\a[31] ,
		\a[32] ,
		\a[52] ,
		\a[53] ,
		_w6667_
	);
	LUT2 #(
		.INIT('h6)
	) name6602 (
		_w6663_,
		_w6667_,
		_w6668_
	);
	LUT4 #(
		.INIT('he11e)
	) name6603 (
		_w6660_,
		_w6661_,
		_w6662_,
		_w6668_,
		_w6669_
	);
	LUT4 #(
		.INIT('h004d)
	) name6604 (
		_w6593_,
		_w6596_,
		_w6601_,
		_w6669_,
		_w6670_
	);
	LUT4 #(
		.INIT('hb200)
	) name6605 (
		_w6593_,
		_w6596_,
		_w6601_,
		_w6669_,
		_w6671_
	);
	LUT4 #(
		.INIT('hf10e)
	) name6606 (
		_w6593_,
		_w6602_,
		_w6603_,
		_w6669_,
		_w6672_
	);
	LUT3 #(
		.INIT('he8)
	) name6607 (
		_w6589_,
		_w6590_,
		_w6591_,
		_w6673_
	);
	LUT3 #(
		.INIT('h0d)
	) name6608 (
		_w6561_,
		_w6562_,
		_w6563_,
		_w6674_
	);
	LUT3 #(
		.INIT('h0d)
	) name6609 (
		_w6570_,
		_w6571_,
		_w6572_,
		_w6675_
	);
	LUT3 #(
		.INIT('h0d)
	) name6610 (
		_w6360_,
		_w6567_,
		_w6568_,
		_w6676_
	);
	LUT3 #(
		.INIT('h96)
	) name6611 (
		_w6674_,
		_w6675_,
		_w6676_,
		_w6677_
	);
	LUT3 #(
		.INIT('h17)
	) name6612 (
		_w6608_,
		_w6609_,
		_w6610_,
		_w6678_
	);
	LUT3 #(
		.INIT('h2b)
	) name6613 (
		_w6612_,
		_w6613_,
		_w6614_,
		_w6679_
	);
	LUT2 #(
		.INIT('h8)
	) name6614 (
		\a[21] ,
		\a[63] ,
		_w6680_
	);
	LUT4 #(
		.INIT('h153f)
	) name6615 (
		\a[22] ,
		\a[23] ,
		\a[61] ,
		\a[62] ,
		_w6681_
	);
	LUT4 #(
		.INIT('h8000)
	) name6616 (
		\a[22] ,
		\a[23] ,
		\a[61] ,
		\a[62] ,
		_w6682_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6617 (
		\a[22] ,
		\a[23] ,
		\a[61] ,
		\a[62] ,
		_w6683_
	);
	LUT2 #(
		.INIT('h8)
	) name6618 (
		\a[33] ,
		\a[51] ,
		_w6684_
	);
	LUT4 #(
		.INIT('h153f)
	) name6619 (
		\a[24] ,
		\a[25] ,
		\a[59] ,
		\a[60] ,
		_w6685_
	);
	LUT2 #(
		.INIT('h8)
	) name6620 (
		\a[25] ,
		\a[60] ,
		_w6686_
	);
	LUT4 #(
		.INIT('h8000)
	) name6621 (
		\a[24] ,
		\a[25] ,
		\a[59] ,
		\a[60] ,
		_w6687_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6622 (
		\a[24] ,
		\a[25] ,
		\a[59] ,
		\a[60] ,
		_w6688_
	);
	LUT4 #(
		.INIT('h0660)
	) name6623 (
		_w6680_,
		_w6683_,
		_w6684_,
		_w6688_,
		_w6689_
	);
	LUT4 #(
		.INIT('h9009)
	) name6624 (
		_w6680_,
		_w6683_,
		_w6684_,
		_w6688_,
		_w6690_
	);
	LUT4 #(
		.INIT('h6996)
	) name6625 (
		_w6680_,
		_w6683_,
		_w6684_,
		_w6688_,
		_w6691_
	);
	LUT2 #(
		.INIT('h8)
	) name6626 (
		\a[34] ,
		\a[50] ,
		_w6692_
	);
	LUT4 #(
		.INIT('h153f)
	) name6627 (
		\a[35] ,
		\a[36] ,
		\a[48] ,
		\a[49] ,
		_w6693_
	);
	LUT2 #(
		.INIT('h8)
	) name6628 (
		\a[36] ,
		\a[49] ,
		_w6694_
	);
	LUT4 #(
		.INIT('h8000)
	) name6629 (
		\a[35] ,
		\a[36] ,
		\a[48] ,
		\a[49] ,
		_w6695_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6630 (
		\a[35] ,
		\a[36] ,
		\a[48] ,
		\a[49] ,
		_w6696_
	);
	LUT2 #(
		.INIT('h6)
	) name6631 (
		_w6692_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h8)
	) name6632 (
		\a[39] ,
		\a[45] ,
		_w6698_
	);
	LUT4 #(
		.INIT('h153f)
	) name6633 (
		\a[40] ,
		\a[41] ,
		\a[43] ,
		\a[44] ,
		_w6699_
	);
	LUT4 #(
		.INIT('h8000)
	) name6634 (
		\a[40] ,
		\a[41] ,
		\a[43] ,
		\a[44] ,
		_w6700_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6635 (
		\a[40] ,
		\a[41] ,
		\a[43] ,
		\a[44] ,
		_w6701_
	);
	LUT2 #(
		.INIT('h8)
	) name6636 (
		\a[28] ,
		\a[56] ,
		_w6702_
	);
	LUT4 #(
		.INIT('h153f)
	) name6637 (
		\a[29] ,
		\a[38] ,
		\a[46] ,
		\a[55] ,
		_w6703_
	);
	LUT4 #(
		.INIT('h8000)
	) name6638 (
		\a[29] ,
		\a[38] ,
		\a[46] ,
		\a[55] ,
		_w6704_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6639 (
		\a[29] ,
		\a[38] ,
		\a[46] ,
		\a[55] ,
		_w6705_
	);
	LUT4 #(
		.INIT('h0660)
	) name6640 (
		_w6698_,
		_w6701_,
		_w6702_,
		_w6705_,
		_w6706_
	);
	LUT4 #(
		.INIT('h9009)
	) name6641 (
		_w6698_,
		_w6701_,
		_w6702_,
		_w6705_,
		_w6707_
	);
	LUT4 #(
		.INIT('h6996)
	) name6642 (
		_w6698_,
		_w6701_,
		_w6702_,
		_w6705_,
		_w6708_
	);
	LUT2 #(
		.INIT('h8)
	) name6643 (
		\a[37] ,
		\a[47] ,
		_w6709_
	);
	LUT4 #(
		.INIT('h153f)
	) name6644 (
		\a[27] ,
		\a[30] ,
		\a[54] ,
		\a[57] ,
		_w6710_
	);
	LUT4 #(
		.INIT('h8000)
	) name6645 (
		\a[27] ,
		\a[30] ,
		\a[54] ,
		\a[57] ,
		_w6711_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6646 (
		\a[27] ,
		\a[30] ,
		\a[54] ,
		\a[57] ,
		_w6712_
	);
	LUT2 #(
		.INIT('h6)
	) name6647 (
		_w6709_,
		_w6712_,
		_w6713_
	);
	LUT4 #(
		.INIT('h0660)
	) name6648 (
		_w6691_,
		_w6697_,
		_w6708_,
		_w6713_,
		_w6714_
	);
	LUT4 #(
		.INIT('h6996)
	) name6649 (
		_w6691_,
		_w6697_,
		_w6708_,
		_w6713_,
		_w6715_
	);
	LUT4 #(
		.INIT('h6900)
	) name6650 (
		_w6677_,
		_w6678_,
		_w6679_,
		_w6715_,
		_w6716_
	);
	LUT4 #(
		.INIT('h9669)
	) name6651 (
		_w6677_,
		_w6678_,
		_w6679_,
		_w6715_,
		_w6717_
	);
	LUT4 #(
		.INIT('h6996)
	) name6652 (
		_w6658_,
		_w6672_,
		_w6673_,
		_w6717_,
		_w6718_
	);
	LUT4 #(
		.INIT('hd400)
	) name6653 (
		_w6588_,
		_w6607_,
		_w6623_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h1)
	) name6654 (
		_w6623_,
		_w6718_,
		_w6720_
	);
	LUT4 #(
		.INIT('h44fd)
	) name6655 (
		_w6588_,
		_w6607_,
		_w6718_,
		_w6720_,
		_w6721_
	);
	LUT4 #(
		.INIT('hf10e)
	) name6656 (
		_w6623_,
		_w6656_,
		_w6657_,
		_w6718_,
		_w6722_
	);
	LUT3 #(
		.INIT('hb4)
	) name6657 (
		_w6653_,
		_w6655_,
		_w6722_,
		_w6723_
	);
	LUT3 #(
		.INIT('h8e)
	) name6658 (
		_w6549_,
		_w6587_,
		_w6624_,
		_w6724_
	);
	LUT2 #(
		.INIT('h8)
	) name6659 (
		_w6723_,
		_w6724_,
		_w6725_
	);
	LUT2 #(
		.INIT('h1)
	) name6660 (
		_w6723_,
		_w6724_,
		_w6726_
	);
	LUT2 #(
		.INIT('h6)
	) name6661 (
		_w6723_,
		_w6724_,
		_w6727_
	);
	LUT4 #(
		.INIT('h0bb0)
	) name6662 (
		_w6548_,
		_w6625_,
		_w6723_,
		_w6724_,
		_w6728_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6663 (
		_w6354_,
		_w6629_,
		_w6632_,
		_w6728_,
		_w6729_
	);
	LUT4 #(
		.INIT('h1033)
	) name6664 (
		_w6354_,
		_w6626_,
		_w6629_,
		_w6632_,
		_w6730_
	);
	LUT3 #(
		.INIT('hcd)
	) name6665 (
		_w6727_,
		_w6729_,
		_w6730_,
		_w6731_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name6666 (
		_w6548_,
		_w6625_,
		_w6723_,
		_w6724_,
		_w6732_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6667 (
		_w6354_,
		_w6629_,
		_w6632_,
		_w6732_,
		_w6733_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name6668 (
		_w6653_,
		_w6655_,
		_w6719_,
		_w6721_,
		_w6734_
	);
	LUT4 #(
		.INIT('hd400)
	) name6669 (
		_w6550_,
		_w6551_,
		_w6583_,
		_w6634_,
		_w6735_
	);
	LUT4 #(
		.INIT('h00ab)
	) name6670 (
		_w6635_,
		_w6651_,
		_w6652_,
		_w6735_,
		_w6736_
	);
	LUT2 #(
		.INIT('h8)
	) name6671 (
		\a[35] ,
		\a[50] ,
		_w6737_
	);
	LUT4 #(
		.INIT('h153f)
	) name6672 (
		\a[22] ,
		\a[28] ,
		\a[57] ,
		\a[63] ,
		_w6738_
	);
	LUT4 #(
		.INIT('h8000)
	) name6673 (
		\a[22] ,
		\a[28] ,
		\a[57] ,
		\a[63] ,
		_w6739_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6674 (
		\a[22] ,
		\a[28] ,
		\a[57] ,
		\a[63] ,
		_w6740_
	);
	LUT4 #(
		.INIT('h153f)
	) name6675 (
		\a[33] ,
		\a[34] ,
		\a[51] ,
		\a[52] ,
		_w6741_
	);
	LUT4 #(
		.INIT('h8000)
	) name6676 (
		\a[33] ,
		\a[34] ,
		\a[51] ,
		\a[52] ,
		_w6742_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6677 (
		\a[33] ,
		\a[34] ,
		\a[51] ,
		\a[52] ,
		_w6743_
	);
	LUT4 #(
		.INIT('h1428)
	) name6678 (
		_w6665_,
		_w6737_,
		_w6740_,
		_w6743_,
		_w6744_
	);
	LUT4 #(
		.INIT('h8241)
	) name6679 (
		_w6665_,
		_w6737_,
		_w6740_,
		_w6743_,
		_w6745_
	);
	LUT4 #(
		.INIT('h6996)
	) name6680 (
		_w6665_,
		_w6737_,
		_w6740_,
		_w6743_,
		_w6746_
	);
	LUT2 #(
		.INIT('h8)
	) name6681 (
		\a[39] ,
		\a[46] ,
		_w6747_
	);
	LUT4 #(
		.INIT('h153f)
	) name6682 (
		\a[40] ,
		\a[41] ,
		\a[44] ,
		\a[45] ,
		_w6748_
	);
	LUT2 #(
		.INIT('h8)
	) name6683 (
		\a[41] ,
		\a[45] ,
		_w6749_
	);
	LUT4 #(
		.INIT('h8000)
	) name6684 (
		\a[40] ,
		\a[41] ,
		\a[44] ,
		\a[45] ,
		_w6750_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6685 (
		\a[40] ,
		\a[41] ,
		\a[44] ,
		\a[45] ,
		_w6751_
	);
	LUT2 #(
		.INIT('h6)
	) name6686 (
		_w6747_,
		_w6751_,
		_w6752_
	);
	LUT4 #(
		.INIT('h153f)
	) name6687 (
		\a[37] ,
		\a[38] ,
		\a[47] ,
		\a[48] ,
		_w6753_
	);
	LUT2 #(
		.INIT('h8)
	) name6688 (
		\a[38] ,
		\a[48] ,
		_w6754_
	);
	LUT4 #(
		.INIT('h8000)
	) name6689 (
		\a[37] ,
		\a[38] ,
		\a[47] ,
		\a[48] ,
		_w6755_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6690 (
		\a[37] ,
		\a[38] ,
		\a[47] ,
		\a[48] ,
		_w6756_
	);
	LUT4 #(
		.INIT('h9a30)
	) name6691 (
		\a[23] ,
		\a[42] ,
		\a[43] ,
		\a[62] ,
		_w6757_
	);
	LUT3 #(
		.INIT('h60)
	) name6692 (
		_w6694_,
		_w6756_,
		_w6757_,
		_w6758_
	);
	LUT3 #(
		.INIT('h09)
	) name6693 (
		_w6694_,
		_w6756_,
		_w6757_,
		_w6759_
	);
	LUT3 #(
		.INIT('h96)
	) name6694 (
		_w6694_,
		_w6756_,
		_w6757_,
		_w6760_
	);
	LUT2 #(
		.INIT('h8)
	) name6695 (
		\a[29] ,
		\a[56] ,
		_w6761_
	);
	LUT4 #(
		.INIT('h153f)
	) name6696 (
		\a[30] ,
		\a[31] ,
		\a[54] ,
		\a[55] ,
		_w6762_
	);
	LUT4 #(
		.INIT('h8000)
	) name6697 (
		\a[30] ,
		\a[31] ,
		\a[54] ,
		\a[55] ,
		_w6763_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6698 (
		\a[30] ,
		\a[31] ,
		\a[54] ,
		\a[55] ,
		_w6764_
	);
	LUT2 #(
		.INIT('h6)
	) name6699 (
		_w6761_,
		_w6764_,
		_w6765_
	);
	LUT4 #(
		.INIT('h0660)
	) name6700 (
		_w6746_,
		_w6752_,
		_w6760_,
		_w6765_,
		_w6766_
	);
	LUT4 #(
		.INIT('h6996)
	) name6701 (
		_w6746_,
		_w6752_,
		_w6760_,
		_w6765_,
		_w6767_
	);
	LUT4 #(
		.INIT('hd400)
	) name6702 (
		_w6641_,
		_w6642_,
		_w6643_,
		_w6767_,
		_w6768_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name6703 (
		_w6641_,
		_w6642_,
		_w6643_,
		_w6767_,
		_w6769_
	);
	LUT3 #(
		.INIT('h0d)
	) name6704 (
		_w6692_,
		_w6693_,
		_w6695_,
		_w6770_
	);
	LUT3 #(
		.INIT('h0d)
	) name6705 (
		_w6680_,
		_w6681_,
		_w6682_,
		_w6771_
	);
	LUT3 #(
		.INIT('h0d)
	) name6706 (
		_w6684_,
		_w6685_,
		_w6687_,
		_w6772_
	);
	LUT3 #(
		.INIT('h96)
	) name6707 (
		_w6770_,
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT3 #(
		.INIT('h32)
	) name6708 (
		_w6706_,
		_w6707_,
		_w6713_,
		_w6774_
	);
	LUT3 #(
		.INIT('h32)
	) name6709 (
		_w6689_,
		_w6690_,
		_w6697_,
		_w6775_
	);
	LUT3 #(
		.INIT('h69)
	) name6710 (
		_w6773_,
		_w6774_,
		_w6775_,
		_w6776_
	);
	LUT3 #(
		.INIT('hd4)
	) name6711 (
		_w6677_,
		_w6678_,
		_w6679_,
		_w6777_
	);
	LUT2 #(
		.INIT('h8)
	) name6712 (
		\a[24] ,
		\a[61] ,
		_w6778_
	);
	LUT4 #(
		.INIT('h0dff)
	) name6713 (
		_w6698_,
		_w6699_,
		_w6700_,
		_w6778_,
		_w6779_
	);
	LUT4 #(
		.INIT('h000d)
	) name6714 (
		_w6698_,
		_w6699_,
		_w6700_,
		_w6778_,
		_w6780_
	);
	LUT4 #(
		.INIT('h0df2)
	) name6715 (
		_w6698_,
		_w6699_,
		_w6700_,
		_w6778_,
		_w6781_
	);
	LUT3 #(
		.INIT('h32)
	) name6716 (
		_w6702_,
		_w6703_,
		_w6704_,
		_w6782_
	);
	LUT2 #(
		.INIT('h6)
	) name6717 (
		_w6781_,
		_w6782_,
		_w6783_
	);
	LUT3 #(
		.INIT('h0d)
	) name6718 (
		_w6663_,
		_w6664_,
		_w6666_,
		_w6784_
	);
	LUT3 #(
		.INIT('h0d)
	) name6719 (
		_w6709_,
		_w6710_,
		_w6711_,
		_w6785_
	);
	LUT4 #(
		.INIT('h153f)
	) name6720 (
		\a[26] ,
		\a[27] ,
		\a[58] ,
		\a[59] ,
		_w6786_
	);
	LUT4 #(
		.INIT('h8000)
	) name6721 (
		\a[26] ,
		\a[27] ,
		\a[58] ,
		\a[59] ,
		_w6787_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6722 (
		\a[26] ,
		\a[27] ,
		\a[58] ,
		\a[59] ,
		_w6788_
	);
	LUT2 #(
		.INIT('h6)
	) name6723 (
		_w6686_,
		_w6788_,
		_w6789_
	);
	LUT3 #(
		.INIT('h69)
	) name6724 (
		_w6784_,
		_w6785_,
		_w6789_,
		_w6790_
	);
	LUT2 #(
		.INIT('h2)
	) name6725 (
		_w6783_,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h4)
	) name6726 (
		_w6783_,
		_w6790_,
		_w6792_
	);
	LUT2 #(
		.INIT('h9)
	) name6727 (
		_w6783_,
		_w6790_,
		_w6793_
	);
	LUT4 #(
		.INIT('h6996)
	) name6728 (
		_w6769_,
		_w6776_,
		_w6777_,
		_w6793_,
		_w6794_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6729 (
		_w6582_,
		_w6645_,
		_w6646_,
		_w6648_,
		_w6795_
	);
	LUT3 #(
		.INIT('h0e)
	) name6730 (
		_w6644_,
		_w6649_,
		_w6795_,
		_w6796_
	);
	LUT3 #(
		.INIT('h17)
	) name6731 (
		_w6674_,
		_w6675_,
		_w6676_,
		_w6797_
	);
	LUT3 #(
		.INIT('h45)
	) name6732 (
		_w6637_,
		_w6638_,
		_w6640_,
		_w6798_
	);
	LUT4 #(
		.INIT('h1f01)
	) name6733 (
		_w6660_,
		_w6661_,
		_w6662_,
		_w6668_,
		_w6799_
	);
	LUT3 #(
		.INIT('h96)
	) name6734 (
		_w6797_,
		_w6798_,
		_w6799_,
		_w6800_
	);
	LUT3 #(
		.INIT('h54)
	) name6735 (
		_w6670_,
		_w6671_,
		_w6673_,
		_w6801_
	);
	LUT4 #(
		.INIT('h0017)
	) name6736 (
		_w6659_,
		_w6669_,
		_w6673_,
		_w6800_,
		_w6802_
	);
	LUT4 #(
		.INIT('he800)
	) name6737 (
		_w6659_,
		_w6669_,
		_w6673_,
		_w6800_,
		_w6803_
	);
	LUT4 #(
		.INIT('hab54)
	) name6738 (
		_w6670_,
		_w6671_,
		_w6673_,
		_w6800_,
		_w6804_
	);
	LUT2 #(
		.INIT('h1)
	) name6739 (
		_w6714_,
		_w6716_,
		_w6805_
	);
	LUT2 #(
		.INIT('h6)
	) name6740 (
		_w6804_,
		_w6805_,
		_w6806_
	);
	LUT4 #(
		.INIT('h41d7)
	) name6741 (
		_w6658_,
		_w6672_,
		_w6673_,
		_w6717_,
		_w6807_
	);
	LUT3 #(
		.INIT('h69)
	) name6742 (
		_w6796_,
		_w6806_,
		_w6807_,
		_w6808_
	);
	LUT2 #(
		.INIT('h1)
	) name6743 (
		_w6735_,
		_w6794_,
		_w6809_
	);
	LUT4 #(
		.INIT('h001e)
	) name6744 (
		_w6653_,
		_w6735_,
		_w6794_,
		_w6808_,
		_w6810_
	);
	LUT3 #(
		.INIT('h40)
	) name6745 (
		_w6653_,
		_w6808_,
		_w6809_,
		_w6811_
	);
	LUT4 #(
		.INIT('hd77d)
	) name6746 (
		_w6794_,
		_w6796_,
		_w6806_,
		_w6807_,
		_w6812_
	);
	LUT2 #(
		.INIT('h1)
	) name6747 (
		_w6736_,
		_w6812_,
		_w6813_
	);
	LUT4 #(
		.INIT('h0001)
	) name6748 (
		_w6734_,
		_w6810_,
		_w6811_,
		_w6813_,
		_w6814_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6749 (
		_w6734_,
		_w6810_,
		_w6811_,
		_w6813_,
		_w6815_
	);
	LUT4 #(
		.INIT('h5556)
	) name6750 (
		_w6734_,
		_w6810_,
		_w6811_,
		_w6813_,
		_w6816_
	);
	LUT3 #(
		.INIT('he1)
	) name6751 (
		_w6726_,
		_w6733_,
		_w6816_,
		_w6817_
	);
	LUT3 #(
		.INIT('h04)
	) name6752 (
		_w6725_,
		_w6726_,
		_w6814_,
		_w6818_
	);
	LUT3 #(
		.INIT('h01)
	) name6753 (
		_w6626_,
		_w6725_,
		_w6814_,
		_w6819_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6754 (
		_w6354_,
		_w6629_,
		_w6632_,
		_w6819_,
		_w6820_
	);
	LUT4 #(
		.INIT('h1f01)
	) name6755 (
		_w6653_,
		_w6735_,
		_w6794_,
		_w6808_,
		_w6821_
	);
	LUT3 #(
		.INIT('h8e)
	) name6756 (
		_w6784_,
		_w6785_,
		_w6789_,
		_w6822_
	);
	LUT3 #(
		.INIT('h45)
	) name6757 (
		_w6744_,
		_w6745_,
		_w6752_,
		_w6823_
	);
	LUT3 #(
		.INIT('h32)
	) name6758 (
		_w6758_,
		_w6759_,
		_w6765_,
		_w6824_
	);
	LUT3 #(
		.INIT('h96)
	) name6759 (
		_w6822_,
		_w6823_,
		_w6824_,
		_w6825_
	);
	LUT3 #(
		.INIT('he8)
	) name6760 (
		_w6797_,
		_w6798_,
		_w6799_,
		_w6826_
	);
	LUT3 #(
		.INIT('h0d)
	) name6761 (
		_w6747_,
		_w6748_,
		_w6750_,
		_w6827_
	);
	LUT3 #(
		.INIT('h0d)
	) name6762 (
		_w6761_,
		_w6762_,
		_w6763_,
		_w6828_
	);
	LUT3 #(
		.INIT('h0d)
	) name6763 (
		_w6694_,
		_w6753_,
		_w6755_,
		_w6829_
	);
	LUT3 #(
		.INIT('h96)
	) name6764 (
		_w6827_,
		_w6828_,
		_w6829_,
		_w6830_
	);
	LUT3 #(
		.INIT('h32)
	) name6765 (
		_w6737_,
		_w6738_,
		_w6739_,
		_w6831_
	);
	LUT3 #(
		.INIT('h0d)
	) name6766 (
		_w6665_,
		_w6741_,
		_w6742_,
		_w6832_
	);
	LUT3 #(
		.INIT('h0d)
	) name6767 (
		_w6686_,
		_w6786_,
		_w6787_,
		_w6833_
	);
	LUT3 #(
		.INIT('h96)
	) name6768 (
		_w6831_,
		_w6832_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h4)
	) name6769 (
		_w6830_,
		_w6834_,
		_w6835_
	);
	LUT2 #(
		.INIT('h2)
	) name6770 (
		_w6830_,
		_w6834_,
		_w6836_
	);
	LUT2 #(
		.INIT('h9)
	) name6771 (
		_w6830_,
		_w6834_,
		_w6837_
	);
	LUT3 #(
		.INIT('h41)
	) name6772 (
		_w6825_,
		_w6826_,
		_w6837_,
		_w6838_
	);
	LUT2 #(
		.INIT('h8)
	) name6773 (
		\a[26] ,
		\a[60] ,
		_w6839_
	);
	LUT4 #(
		.INIT('h153f)
	) name6774 (
		\a[27] ,
		\a[28] ,
		\a[58] ,
		\a[59] ,
		_w6840_
	);
	LUT2 #(
		.INIT('h8)
	) name6775 (
		\a[28] ,
		\a[59] ,
		_w6841_
	);
	LUT4 #(
		.INIT('h8000)
	) name6776 (
		\a[27] ,
		\a[28] ,
		\a[58] ,
		\a[59] ,
		_w6842_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6777 (
		\a[27] ,
		\a[28] ,
		\a[58] ,
		\a[59] ,
		_w6843_
	);
	LUT4 #(
		.INIT('h153f)
	) name6778 (
		\a[32] ,
		\a[42] ,
		\a[44] ,
		\a[54] ,
		_w6844_
	);
	LUT4 #(
		.INIT('h8000)
	) name6779 (
		\a[32] ,
		\a[42] ,
		\a[44] ,
		\a[54] ,
		_w6845_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6780 (
		\a[32] ,
		\a[42] ,
		\a[44] ,
		\a[54] ,
		_w6846_
	);
	LUT4 #(
		.INIT('h1428)
	) name6781 (
		_w6749_,
		_w6839_,
		_w6843_,
		_w6846_,
		_w6847_
	);
	LUT4 #(
		.INIT('h8241)
	) name6782 (
		_w6749_,
		_w6839_,
		_w6843_,
		_w6846_,
		_w6848_
	);
	LUT4 #(
		.INIT('h6996)
	) name6783 (
		_w6749_,
		_w6839_,
		_w6843_,
		_w6846_,
		_w6849_
	);
	LUT2 #(
		.INIT('h8)
	) name6784 (
		\a[30] ,
		\a[56] ,
		_w6850_
	);
	LUT4 #(
		.INIT('h153f)
	) name6785 (
		\a[39] ,
		\a[40] ,
		\a[46] ,
		\a[47] ,
		_w6851_
	);
	LUT2 #(
		.INIT('h8)
	) name6786 (
		\a[40] ,
		\a[47] ,
		_w6852_
	);
	LUT4 #(
		.INIT('h8000)
	) name6787 (
		\a[39] ,
		\a[40] ,
		\a[46] ,
		\a[47] ,
		_w6853_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6788 (
		\a[39] ,
		\a[40] ,
		\a[46] ,
		\a[47] ,
		_w6854_
	);
	LUT2 #(
		.INIT('h6)
	) name6789 (
		_w6850_,
		_w6854_,
		_w6855_
	);
	LUT2 #(
		.INIT('h8)
	) name6790 (
		\a[23] ,
		\a[63] ,
		_w6856_
	);
	LUT4 #(
		.INIT('h153f)
	) name6791 (
		\a[36] ,
		\a[37] ,
		\a[49] ,
		\a[50] ,
		_w6857_
	);
	LUT2 #(
		.INIT('h8)
	) name6792 (
		\a[37] ,
		\a[50] ,
		_w6858_
	);
	LUT4 #(
		.INIT('h8000)
	) name6793 (
		\a[36] ,
		\a[37] ,
		\a[49] ,
		\a[50] ,
		_w6859_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6794 (
		\a[36] ,
		\a[37] ,
		\a[49] ,
		\a[50] ,
		_w6860_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		\a[33] ,
		\a[53] ,
		_w6861_
	);
	LUT4 #(
		.INIT('h153f)
	) name6796 (
		\a[34] ,
		\a[35] ,
		\a[51] ,
		\a[52] ,
		_w6862_
	);
	LUT2 #(
		.INIT('h8)
	) name6797 (
		\a[35] ,
		\a[52] ,
		_w6863_
	);
	LUT4 #(
		.INIT('h8000)
	) name6798 (
		\a[34] ,
		\a[35] ,
		\a[51] ,
		\a[52] ,
		_w6864_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6799 (
		\a[34] ,
		\a[35] ,
		\a[51] ,
		\a[52] ,
		_w6865_
	);
	LUT4 #(
		.INIT('h0660)
	) name6800 (
		_w6856_,
		_w6860_,
		_w6861_,
		_w6865_,
		_w6866_
	);
	LUT4 #(
		.INIT('h9009)
	) name6801 (
		_w6856_,
		_w6860_,
		_w6861_,
		_w6865_,
		_w6867_
	);
	LUT4 #(
		.INIT('h6996)
	) name6802 (
		_w6856_,
		_w6860_,
		_w6861_,
		_w6865_,
		_w6868_
	);
	LUT4 #(
		.INIT('h153f)
	) name6803 (
		\a[29] ,
		\a[31] ,
		\a[55] ,
		\a[57] ,
		_w6869_
	);
	LUT2 #(
		.INIT('h8)
	) name6804 (
		\a[31] ,
		\a[57] ,
		_w6870_
	);
	LUT4 #(
		.INIT('h8000)
	) name6805 (
		\a[29] ,
		\a[31] ,
		\a[55] ,
		\a[57] ,
		_w6871_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6806 (
		\a[29] ,
		\a[31] ,
		\a[55] ,
		\a[57] ,
		_w6872_
	);
	LUT2 #(
		.INIT('h6)
	) name6807 (
		_w6754_,
		_w6872_,
		_w6873_
	);
	LUT4 #(
		.INIT('h0660)
	) name6808 (
		_w6849_,
		_w6855_,
		_w6868_,
		_w6873_,
		_w6874_
	);
	LUT4 #(
		.INIT('h6996)
	) name6809 (
		_w6849_,
		_w6855_,
		_w6868_,
		_w6873_,
		_w6875_
	);
	LUT4 #(
		.INIT('hd400)
	) name6810 (
		_w6773_,
		_w6774_,
		_w6775_,
		_w6875_,
		_w6876_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name6811 (
		_w6773_,
		_w6774_,
		_w6775_,
		_w6875_,
		_w6877_
	);
	LUT4 #(
		.INIT('h6996)
	) name6812 (
		_w6825_,
		_w6826_,
		_w6837_,
		_w6877_,
		_w6878_
	);
	LUT4 #(
		.INIT('h00d4)
	) name6813 (
		_w6796_,
		_w6806_,
		_w6807_,
		_w6878_,
		_w6879_
	);
	LUT4 #(
		.INIT('h8ee8)
	) name6814 (
		_w6769_,
		_w6776_,
		_w6777_,
		_w6793_,
		_w6880_
	);
	LUT3 #(
		.INIT('h45)
	) name6815 (
		_w6802_,
		_w6803_,
		_w6805_,
		_w6881_
	);
	LUT4 #(
		.INIT('h0071)
	) name6816 (
		_w6800_,
		_w6801_,
		_w6805_,
		_w6880_,
		_w6882_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6817 (
		_w6800_,
		_w6801_,
		_w6805_,
		_w6880_,
		_w6883_
	);
	LUT4 #(
		.INIT('hba45)
	) name6818 (
		_w6802_,
		_w6803_,
		_w6805_,
		_w6880_,
		_w6884_
	);
	LUT4 #(
		.INIT('h153f)
	) name6819 (
		\a[24] ,
		\a[25] ,
		\a[61] ,
		\a[62] ,
		_w6885_
	);
	LUT4 #(
		.INIT('h8000)
	) name6820 (
		\a[24] ,
		\a[25] ,
		\a[61] ,
		\a[62] ,
		_w6886_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6821 (
		\a[24] ,
		\a[25] ,
		\a[61] ,
		\a[62] ,
		_w6887_
	);
	LUT4 #(
		.INIT('he0c0)
	) name6822 (
		\a[23] ,
		\a[42] ,
		\a[43] ,
		\a[62] ,
		_w6888_
	);
	LUT2 #(
		.INIT('h6)
	) name6823 (
		_w6887_,
		_w6888_,
		_w6889_
	);
	LUT4 #(
		.INIT('h008a)
	) name6824 (
		_w6779_,
		_w6780_,
		_w6782_,
		_w6889_,
		_w6890_
	);
	LUT4 #(
		.INIT('h7500)
	) name6825 (
		_w6779_,
		_w6780_,
		_w6782_,
		_w6889_,
		_w6891_
	);
	LUT4 #(
		.INIT('hf20d)
	) name6826 (
		_w6779_,
		_w6782_,
		_w6780_,
		_w6889_,
		_w6892_
	);
	LUT3 #(
		.INIT('h17)
	) name6827 (
		_w6770_,
		_w6771_,
		_w6772_,
		_w6893_
	);
	LUT2 #(
		.INIT('h6)
	) name6828 (
		_w6892_,
		_w6893_,
		_w6894_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6829 (
		_w6777_,
		_w6783_,
		_w6790_,
		_w6894_,
		_w6895_
	);
	LUT4 #(
		.INIT('hd00d)
	) name6830 (
		_w6783_,
		_w6790_,
		_w6892_,
		_w6893_,
		_w6896_
	);
	LUT3 #(
		.INIT('h70)
	) name6831 (
		_w6777_,
		_w6793_,
		_w6896_,
		_w6897_
	);
	LUT4 #(
		.INIT('h31ce)
	) name6832 (
		_w6777_,
		_w6791_,
		_w6792_,
		_w6894_,
		_w6898_
	);
	LUT2 #(
		.INIT('h1)
	) name6833 (
		_w6766_,
		_w6768_,
		_w6899_
	);
	LUT2 #(
		.INIT('h6)
	) name6834 (
		_w6898_,
		_w6899_,
		_w6900_
	);
	LUT2 #(
		.INIT('h9)
	) name6835 (
		_w6884_,
		_w6900_,
		_w6901_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6836 (
		_w6796_,
		_w6806_,
		_w6807_,
		_w6878_,
		_w6902_
	);
	LUT3 #(
		.INIT('hc9)
	) name6837 (
		_w6879_,
		_w6901_,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h2)
	) name6838 (
		_w6821_,
		_w6903_,
		_w6904_
	);
	LUT2 #(
		.INIT('h9)
	) name6839 (
		_w6821_,
		_w6903_,
		_w6905_
	);
	LUT4 #(
		.INIT('hfe01)
	) name6840 (
		_w6815_,
		_w6818_,
		_w6820_,
		_w6905_,
		_w6906_
	);
	LUT2 #(
		.INIT('h1)
	) name6841 (
		_w6815_,
		_w6904_,
		_w6907_
	);
	LUT3 #(
		.INIT('h54)
	) name6842 (
		_w6879_,
		_w6901_,
		_w6902_,
		_w6908_
	);
	LUT3 #(
		.INIT('h17)
	) name6843 (
		_w6827_,
		_w6828_,
		_w6829_,
		_w6909_
	);
	LUT3 #(
		.INIT('h32)
	) name6844 (
		_w6866_,
		_w6867_,
		_w6873_,
		_w6910_
	);
	LUT3 #(
		.INIT('h32)
	) name6845 (
		_w6847_,
		_w6848_,
		_w6855_,
		_w6911_
	);
	LUT3 #(
		.INIT('h96)
	) name6846 (
		_w6909_,
		_w6910_,
		_w6911_,
		_w6912_
	);
	LUT3 #(
		.INIT('he0)
	) name6847 (
		_w6874_,
		_w6876_,
		_w6912_,
		_w6913_
	);
	LUT3 #(
		.INIT('h1e)
	) name6848 (
		_w6874_,
		_w6876_,
		_w6912_,
		_w6914_
	);
	LUT4 #(
		.INIT('h2300)
	) name6849 (
		_w6895_,
		_w6897_,
		_w6899_,
		_w6914_,
		_w6915_
	);
	LUT4 #(
		.INIT('hdc23)
	) name6850 (
		_w6895_,
		_w6897_,
		_w6899_,
		_w6914_,
		_w6916_
	);
	LUT4 #(
		.INIT('h0071)
	) name6851 (
		_w6880_,
		_w6881_,
		_w6900_,
		_w6916_,
		_w6917_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6852 (
		_w6880_,
		_w6881_,
		_w6900_,
		_w6916_,
		_w6918_
	);
	LUT4 #(
		.INIT('hba45)
	) name6853 (
		_w6882_,
		_w6883_,
		_w6900_,
		_w6916_,
		_w6919_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6854 (
		_w6825_,
		_w6826_,
		_w6837_,
		_w6877_,
		_w6920_
	);
	LUT4 #(
		.INIT('h153f)
	) name6855 (
		\a[31] ,
		\a[33] ,
		\a[54] ,
		\a[56] ,
		_w6921_
	);
	LUT4 #(
		.INIT('h8000)
	) name6856 (
		\a[31] ,
		\a[33] ,
		\a[54] ,
		\a[56] ,
		_w6922_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6857 (
		\a[31] ,
		\a[33] ,
		\a[54] ,
		\a[56] ,
		_w6923_
	);
	LUT4 #(
		.INIT('h9a30)
	) name6858 (
		\a[25] ,
		\a[43] ,
		\a[44] ,
		\a[62] ,
		_w6924_
	);
	LUT3 #(
		.INIT('h60)
	) name6859 (
		_w6852_,
		_w6923_,
		_w6924_,
		_w6925_
	);
	LUT3 #(
		.INIT('h96)
	) name6860 (
		_w6852_,
		_w6923_,
		_w6924_,
		_w6926_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6861 (
		_w6831_,
		_w6832_,
		_w6833_,
		_w6926_,
		_w6927_
	);
	LUT4 #(
		.INIT('hd42b)
	) name6862 (
		_w6831_,
		_w6832_,
		_w6833_,
		_w6926_,
		_w6928_
	);
	LUT2 #(
		.INIT('h8)
	) name6863 (
		\a[24] ,
		\a[63] ,
		_w6929_
	);
	LUT4 #(
		.INIT('h153f)
	) name6864 (
		\a[26] ,
		\a[27] ,
		\a[60] ,
		\a[61] ,
		_w6930_
	);
	LUT4 #(
		.INIT('h8000)
	) name6865 (
		\a[26] ,
		\a[27] ,
		\a[60] ,
		\a[61] ,
		_w6931_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6866 (
		\a[26] ,
		\a[27] ,
		\a[60] ,
		\a[61] ,
		_w6932_
	);
	LUT4 #(
		.INIT('h153f)
	) name6867 (
		\a[38] ,
		\a[39] ,
		\a[48] ,
		\a[49] ,
		_w6933_
	);
	LUT4 #(
		.INIT('h8000)
	) name6868 (
		\a[38] ,
		\a[39] ,
		\a[48] ,
		\a[49] ,
		_w6934_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6869 (
		\a[38] ,
		\a[39] ,
		\a[48] ,
		\a[49] ,
		_w6935_
	);
	LUT4 #(
		.INIT('h1428)
	) name6870 (
		_w6858_,
		_w6929_,
		_w6932_,
		_w6935_,
		_w6936_
	);
	LUT4 #(
		.INIT('h8241)
	) name6871 (
		_w6858_,
		_w6929_,
		_w6932_,
		_w6935_,
		_w6937_
	);
	LUT4 #(
		.INIT('h6996)
	) name6872 (
		_w6858_,
		_w6929_,
		_w6932_,
		_w6935_,
		_w6938_
	);
	LUT2 #(
		.INIT('h8)
	) name6873 (
		\a[32] ,
		\a[55] ,
		_w6939_
	);
	LUT4 #(
		.INIT('h153f)
	) name6874 (
		\a[41] ,
		\a[42] ,
		\a[45] ,
		\a[46] ,
		_w6940_
	);
	LUT4 #(
		.INIT('h8000)
	) name6875 (
		\a[41] ,
		\a[42] ,
		\a[45] ,
		\a[46] ,
		_w6941_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6876 (
		\a[41] ,
		\a[42] ,
		\a[45] ,
		\a[46] ,
		_w6942_
	);
	LUT2 #(
		.INIT('h6)
	) name6877 (
		_w6939_,
		_w6942_,
		_w6943_
	);
	LUT2 #(
		.INIT('h6)
	) name6878 (
		_w6938_,
		_w6943_,
		_w6944_
	);
	LUT3 #(
		.INIT('h23)
	) name6879 (
		_w6885_,
		_w6886_,
		_w6888_,
		_w6945_
	);
	LUT4 #(
		.INIT('h153f)
	) name6880 (
		\a[30] ,
		\a[34] ,
		\a[53] ,
		\a[57] ,
		_w6946_
	);
	LUT4 #(
		.INIT('h8000)
	) name6881 (
		\a[30] ,
		\a[34] ,
		\a[53] ,
		\a[57] ,
		_w6947_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6882 (
		\a[30] ,
		\a[34] ,
		\a[53] ,
		\a[57] ,
		_w6948_
	);
	LUT2 #(
		.INIT('h6)
	) name6883 (
		_w6841_,
		_w6948_,
		_w6949_
	);
	LUT4 #(
		.INIT('h153f)
	) name6884 (
		\a[29] ,
		\a[36] ,
		\a[51] ,
		\a[58] ,
		_w6950_
	);
	LUT4 #(
		.INIT('h8000)
	) name6885 (
		\a[29] ,
		\a[36] ,
		\a[51] ,
		\a[58] ,
		_w6951_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6886 (
		\a[29] ,
		\a[36] ,
		\a[51] ,
		\a[58] ,
		_w6952_
	);
	LUT2 #(
		.INIT('h6)
	) name6887 (
		_w6863_,
		_w6952_,
		_w6953_
	);
	LUT3 #(
		.INIT('h69)
	) name6888 (
		_w6945_,
		_w6949_,
		_w6953_,
		_w6954_
	);
	LUT3 #(
		.INIT('h96)
	) name6889 (
		_w6928_,
		_w6944_,
		_w6954_,
		_w6955_
	);
	LUT4 #(
		.INIT('hbe00)
	) name6890 (
		_w6825_,
		_w6826_,
		_w6837_,
		_w6955_,
		_w6956_
	);
	LUT4 #(
		.INIT('hbe28)
	) name6891 (
		_w6825_,
		_w6826_,
		_w6837_,
		_w6877_,
		_w6957_
	);
	LUT2 #(
		.INIT('h1)
	) name6892 (
		_w6955_,
		_w6957_,
		_w6958_
	);
	LUT3 #(
		.INIT('he1)
	) name6893 (
		_w6838_,
		_w6920_,
		_w6955_,
		_w6959_
	);
	LUT3 #(
		.INIT('h31)
	) name6894 (
		_w6826_,
		_w6835_,
		_w6836_,
		_w6960_
	);
	LUT3 #(
		.INIT('h71)
	) name6895 (
		_w6822_,
		_w6823_,
		_w6824_,
		_w6961_
	);
	LUT4 #(
		.INIT('h004d)
	) name6896 (
		_w6826_,
		_w6830_,
		_w6834_,
		_w6961_,
		_w6962_
	);
	LUT4 #(
		.INIT('hb200)
	) name6897 (
		_w6826_,
		_w6830_,
		_w6834_,
		_w6961_,
		_w6963_
	);
	LUT4 #(
		.INIT('h31ce)
	) name6898 (
		_w6826_,
		_w6835_,
		_w6836_,
		_w6961_,
		_w6964_
	);
	LUT3 #(
		.INIT('h54)
	) name6899 (
		_w6890_,
		_w6891_,
		_w6893_,
		_w6965_
	);
	LUT3 #(
		.INIT('h32)
	) name6900 (
		_w6749_,
		_w6844_,
		_w6845_,
		_w6966_
	);
	LUT3 #(
		.INIT('h0d)
	) name6901 (
		_w6850_,
		_w6851_,
		_w6853_,
		_w6967_
	);
	LUT3 #(
		.INIT('h0d)
	) name6902 (
		_w6754_,
		_w6869_,
		_w6871_,
		_w6968_
	);
	LUT3 #(
		.INIT('h69)
	) name6903 (
		_w6966_,
		_w6967_,
		_w6968_,
		_w6969_
	);
	LUT3 #(
		.INIT('h0d)
	) name6904 (
		_w6861_,
		_w6862_,
		_w6864_,
		_w6970_
	);
	LUT3 #(
		.INIT('h0d)
	) name6905 (
		_w6839_,
		_w6840_,
		_w6842_,
		_w6971_
	);
	LUT3 #(
		.INIT('h0d)
	) name6906 (
		_w6856_,
		_w6857_,
		_w6859_,
		_w6972_
	);
	LUT3 #(
		.INIT('h96)
	) name6907 (
		_w6970_,
		_w6971_,
		_w6972_,
		_w6973_
	);
	LUT2 #(
		.INIT('h8)
	) name6908 (
		_w6969_,
		_w6973_,
		_w6974_
	);
	LUT2 #(
		.INIT('h1)
	) name6909 (
		_w6969_,
		_w6973_,
		_w6975_
	);
	LUT2 #(
		.INIT('h6)
	) name6910 (
		_w6969_,
		_w6973_,
		_w6976_
	);
	LUT2 #(
		.INIT('h6)
	) name6911 (
		_w6965_,
		_w6976_,
		_w6977_
	);
	LUT2 #(
		.INIT('h6)
	) name6912 (
		_w6964_,
		_w6977_,
		_w6978_
	);
	LUT2 #(
		.INIT('h6)
	) name6913 (
		_w6959_,
		_w6978_,
		_w6979_
	);
	LUT2 #(
		.INIT('h6)
	) name6914 (
		_w6919_,
		_w6979_,
		_w6980_
	);
	LUT2 #(
		.INIT('h1)
	) name6915 (
		_w6908_,
		_w6980_,
		_w6981_
	);
	LUT2 #(
		.INIT('h8)
	) name6916 (
		_w6908_,
		_w6980_,
		_w6982_
	);
	LUT2 #(
		.INIT('h6)
	) name6917 (
		_w6908_,
		_w6980_,
		_w6983_
	);
	LUT3 #(
		.INIT('hb0)
	) name6918 (
		_w6821_,
		_w6903_,
		_w6983_,
		_w6984_
	);
	LUT4 #(
		.INIT('hef00)
	) name6919 (
		_w6818_,
		_w6820_,
		_w6907_,
		_w6984_,
		_w6985_
	);
	LUT3 #(
		.INIT('h04)
	) name6920 (
		_w6821_,
		_w6903_,
		_w6983_,
		_w6986_
	);
	LUT3 #(
		.INIT('h01)
	) name6921 (
		_w6815_,
		_w6904_,
		_w6983_,
		_w6987_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name6922 (
		_w6818_,
		_w6820_,
		_w6986_,
		_w6987_,
		_w6988_
	);
	LUT2 #(
		.INIT('hb)
	) name6923 (
		_w6985_,
		_w6988_,
		_w6989_
	);
	LUT3 #(
		.INIT('h0b)
	) name6924 (
		_w6821_,
		_w6903_,
		_w6982_,
		_w6990_
	);
	LUT4 #(
		.INIT('hef00)
	) name6925 (
		_w6818_,
		_w6820_,
		_w6907_,
		_w6990_,
		_w6991_
	);
	LUT3 #(
		.INIT('h54)
	) name6926 (
		_w6917_,
		_w6918_,
		_w6979_,
		_w6992_
	);
	LUT4 #(
		.INIT('hb00b)
	) name6927 (
		_w6920_,
		_w6956_,
		_w6964_,
		_w6977_,
		_w6993_
	);
	LUT3 #(
		.INIT('h17)
	) name6928 (
		_w6970_,
		_w6971_,
		_w6972_,
		_w6994_
	);
	LUT3 #(
		.INIT('hd4)
	) name6929 (
		_w6945_,
		_w6949_,
		_w6953_,
		_w6995_
	);
	LUT3 #(
		.INIT('h32)
	) name6930 (
		_w6936_,
		_w6937_,
		_w6943_,
		_w6996_
	);
	LUT3 #(
		.INIT('h96)
	) name6931 (
		_w6994_,
		_w6995_,
		_w6996_,
		_w6997_
	);
	LUT3 #(
		.INIT('he8)
	) name6932 (
		_w6928_,
		_w6944_,
		_w6954_,
		_w6998_
	);
	LUT2 #(
		.INIT('h8)
	) name6933 (
		_w6997_,
		_w6998_,
		_w6999_
	);
	LUT2 #(
		.INIT('h6)
	) name6934 (
		_w6997_,
		_w6998_,
		_w7000_
	);
	LUT4 #(
		.INIT('hd400)
	) name6935 (
		_w6960_,
		_w6961_,
		_w6977_,
		_w7000_,
		_w7001_
	);
	LUT4 #(
		.INIT('hab54)
	) name6936 (
		_w6962_,
		_w6963_,
		_w6977_,
		_w7000_,
		_w7002_
	);
	LUT3 #(
		.INIT('h10)
	) name6937 (
		_w6958_,
		_w6993_,
		_w7002_,
		_w7003_
	);
	LUT3 #(
		.INIT('h0e)
	) name6938 (
		_w6958_,
		_w6993_,
		_w7002_,
		_w7004_
	);
	LUT3 #(
		.INIT('he1)
	) name6939 (
		_w6958_,
		_w6993_,
		_w7002_,
		_w7005_
	);
	LUT2 #(
		.INIT('h8)
	) name6940 (
		\a[29] ,
		\a[59] ,
		_w7006_
	);
	LUT4 #(
		.INIT('h153f)
	) name6941 (
		\a[38] ,
		\a[39] ,
		\a[49] ,
		\a[50] ,
		_w7007_
	);
	LUT4 #(
		.INIT('h8000)
	) name6942 (
		\a[38] ,
		\a[39] ,
		\a[49] ,
		\a[50] ,
		_w7008_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6943 (
		\a[38] ,
		\a[39] ,
		\a[49] ,
		\a[50] ,
		_w7009_
	);
	LUT2 #(
		.INIT('h8)
	) name6944 (
		\a[40] ,
		\a[48] ,
		_w7010_
	);
	LUT4 #(
		.INIT('h153f)
	) name6945 (
		\a[30] ,
		\a[32] ,
		\a[56] ,
		\a[58] ,
		_w7011_
	);
	LUT4 #(
		.INIT('h8000)
	) name6946 (
		\a[30] ,
		\a[32] ,
		\a[56] ,
		\a[58] ,
		_w7012_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6947 (
		\a[30] ,
		\a[32] ,
		\a[56] ,
		\a[58] ,
		_w7013_
	);
	LUT4 #(
		.INIT('h0660)
	) name6948 (
		_w7006_,
		_w7009_,
		_w7010_,
		_w7013_,
		_w7014_
	);
	LUT4 #(
		.INIT('h6996)
	) name6949 (
		_w7006_,
		_w7009_,
		_w7010_,
		_w7013_,
		_w7015_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6950 (
		_w6966_,
		_w6967_,
		_w6968_,
		_w7015_,
		_w7016_
	);
	LUT4 #(
		.INIT('hd42b)
	) name6951 (
		_w6966_,
		_w6967_,
		_w6968_,
		_w7015_,
		_w7017_
	);
	LUT3 #(
		.INIT('h13)
	) name6952 (
		\a[25] ,
		\a[43] ,
		\a[62] ,
		_w7018_
	);
	LUT2 #(
		.INIT('h8)
	) name6953 (
		\a[25] ,
		\a[63] ,
		_w7019_
	);
	LUT3 #(
		.INIT('h80)
	) name6954 (
		\a[25] ,
		\a[44] ,
		\a[63] ,
		_w7020_
	);
	LUT2 #(
		.INIT('h4)
	) name6955 (
		_w7018_,
		_w7020_,
		_w7021_
	);
	LUT4 #(
		.INIT('he0c0)
	) name6956 (
		\a[25] ,
		\a[43] ,
		\a[44] ,
		\a[62] ,
		_w7022_
	);
	LUT2 #(
		.INIT('h1)
	) name6957 (
		_w7019_,
		_w7022_,
		_w7023_
	);
	LUT3 #(
		.INIT('hd2)
	) name6958 (
		\a[44] ,
		_w7018_,
		_w7019_,
		_w7024_
	);
	LUT3 #(
		.INIT('h0d)
	) name6959 (
		_w6939_,
		_w6940_,
		_w6941_,
		_w7025_
	);
	LUT2 #(
		.INIT('h6)
	) name6960 (
		_w7024_,
		_w7025_,
		_w7026_
	);
	LUT2 #(
		.INIT('h8)
	) name6961 (
		\a[26] ,
		\a[62] ,
		_w7027_
	);
	LUT4 #(
		.INIT('h153f)
	) name6962 (
		\a[27] ,
		\a[28] ,
		\a[60] ,
		\a[61] ,
		_w7028_
	);
	LUT4 #(
		.INIT('h8000)
	) name6963 (
		\a[27] ,
		\a[28] ,
		\a[60] ,
		\a[61] ,
		_w7029_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6964 (
		\a[27] ,
		\a[28] ,
		\a[60] ,
		\a[61] ,
		_w7030_
	);
	LUT4 #(
		.INIT('h153f)
	) name6965 (
		\a[41] ,
		\a[42] ,
		\a[46] ,
		\a[47] ,
		_w7031_
	);
	LUT4 #(
		.INIT('h8000)
	) name6966 (
		\a[41] ,
		\a[42] ,
		\a[46] ,
		\a[47] ,
		_w7032_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6967 (
		\a[41] ,
		\a[42] ,
		\a[46] ,
		\a[47] ,
		_w7033_
	);
	LUT4 #(
		.INIT('h1428)
	) name6968 (
		_w6870_,
		_w7027_,
		_w7030_,
		_w7033_,
		_w7034_
	);
	LUT4 #(
		.INIT('h8241)
	) name6969 (
		_w6870_,
		_w7027_,
		_w7030_,
		_w7033_,
		_w7035_
	);
	LUT4 #(
		.INIT('h6996)
	) name6970 (
		_w6870_,
		_w7027_,
		_w7030_,
		_w7033_,
		_w7036_
	);
	LUT2 #(
		.INIT('h8)
	) name6971 (
		\a[35] ,
		\a[53] ,
		_w7037_
	);
	LUT4 #(
		.INIT('h153f)
	) name6972 (
		\a[36] ,
		\a[37] ,
		\a[51] ,
		\a[52] ,
		_w7038_
	);
	LUT4 #(
		.INIT('h8000)
	) name6973 (
		\a[36] ,
		\a[37] ,
		\a[51] ,
		\a[52] ,
		_w7039_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6974 (
		\a[36] ,
		\a[37] ,
		\a[51] ,
		\a[52] ,
		_w7040_
	);
	LUT2 #(
		.INIT('h6)
	) name6975 (
		_w7037_,
		_w7040_,
		_w7041_
	);
	LUT2 #(
		.INIT('h6)
	) name6976 (
		_w7036_,
		_w7041_,
		_w7042_
	);
	LUT3 #(
		.INIT('h69)
	) name6977 (
		_w7017_,
		_w7026_,
		_w7042_,
		_w7043_
	);
	LUT3 #(
		.INIT('h32)
	) name6978 (
		_w6965_,
		_w6974_,
		_w6975_,
		_w7044_
	);
	LUT3 #(
		.INIT('he8)
	) name6979 (
		_w6909_,
		_w6910_,
		_w6911_,
		_w7045_
	);
	LUT4 #(
		.INIT('h00d4)
	) name6980 (
		_w6965_,
		_w6969_,
		_w6973_,
		_w7045_,
		_w7046_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6981 (
		_w6965_,
		_w6969_,
		_w6973_,
		_w7045_,
		_w7047_
	);
	LUT4 #(
		.INIT('hcd32)
	) name6982 (
		_w6965_,
		_w6974_,
		_w6975_,
		_w7045_,
		_w7048_
	);
	LUT3 #(
		.INIT('h32)
	) name6983 (
		_w6841_,
		_w6946_,
		_w6947_,
		_w7049_
	);
	LUT3 #(
		.INIT('h0d)
	) name6984 (
		_w6929_,
		_w6930_,
		_w6931_,
		_w7050_
	);
	LUT3 #(
		.INIT('h0d)
	) name6985 (
		_w6858_,
		_w6933_,
		_w6934_,
		_w7051_
	);
	LUT3 #(
		.INIT('h69)
	) name6986 (
		_w7049_,
		_w7050_,
		_w7051_,
		_w7052_
	);
	LUT3 #(
		.INIT('h32)
	) name6987 (
		_w6863_,
		_w6950_,
		_w6951_,
		_w7053_
	);
	LUT3 #(
		.INIT('h0d)
	) name6988 (
		_w6852_,
		_w6921_,
		_w6922_,
		_w7054_
	);
	LUT2 #(
		.INIT('h8)
	) name6989 (
		\a[43] ,
		\a[45] ,
		_w7055_
	);
	LUT4 #(
		.INIT('h153f)
	) name6990 (
		\a[33] ,
		\a[34] ,
		\a[54] ,
		\a[55] ,
		_w7056_
	);
	LUT2 #(
		.INIT('h8)
	) name6991 (
		\a[34] ,
		\a[55] ,
		_w7057_
	);
	LUT4 #(
		.INIT('h8000)
	) name6992 (
		\a[33] ,
		\a[34] ,
		\a[54] ,
		\a[55] ,
		_w7058_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name6993 (
		\a[33] ,
		\a[34] ,
		\a[54] ,
		\a[55] ,
		_w7059_
	);
	LUT2 #(
		.INIT('h6)
	) name6994 (
		_w7055_,
		_w7059_,
		_w7060_
	);
	LUT3 #(
		.INIT('h69)
	) name6995 (
		_w7053_,
		_w7054_,
		_w7060_,
		_w7061_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6996 (
		_w6925_,
		_w6927_,
		_w7052_,
		_w7061_,
		_w7062_
	);
	LUT2 #(
		.INIT('h6)
	) name6997 (
		_w7048_,
		_w7062_,
		_w7063_
	);
	LUT4 #(
		.INIT('h001f)
	) name6998 (
		_w6874_,
		_w6876_,
		_w6912_,
		_w7043_,
		_w7064_
	);
	LUT4 #(
		.INIT('h1e00)
	) name6999 (
		_w6913_,
		_w6915_,
		_w7043_,
		_w7063_,
		_w7065_
	);
	LUT3 #(
		.INIT('h90)
	) name7000 (
		_w7048_,
		_w7062_,
		_w7064_,
		_w7066_
	);
	LUT3 #(
		.INIT('h82)
	) name7001 (
		_w7043_,
		_w7048_,
		_w7062_,
		_w7067_
	);
	LUT4 #(
		.INIT('h01cf)
	) name7002 (
		_w6913_,
		_w6915_,
		_w7066_,
		_w7067_,
		_w7068_
	);
	LUT3 #(
		.INIT('h9a)
	) name7003 (
		_w7005_,
		_w7065_,
		_w7068_,
		_w7069_
	);
	LUT2 #(
		.INIT('h6)
	) name7004 (
		_w6992_,
		_w7069_,
		_w7070_
	);
	LUT3 #(
		.INIT('he1)
	) name7005 (
		_w6981_,
		_w6991_,
		_w7070_,
		_w7071_
	);
	LUT3 #(
		.INIT('h0d)
	) name7006 (
		_w7037_,
		_w7038_,
		_w7039_,
		_w7072_
	);
	LUT3 #(
		.INIT('h0d)
	) name7007 (
		_w7027_,
		_w7028_,
		_w7029_,
		_w7073_
	);
	LUT3 #(
		.INIT('h0d)
	) name7008 (
		_w7010_,
		_w7011_,
		_w7012_,
		_w7074_
	);
	LUT3 #(
		.INIT('h96)
	) name7009 (
		_w7072_,
		_w7073_,
		_w7074_,
		_w7075_
	);
	LUT4 #(
		.INIT('h8000)
	) name7010 (
		\a[28] ,
		\a[29] ,
		\a[60] ,
		\a[61] ,
		_w7076_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7011 (
		\a[28] ,
		\a[29] ,
		\a[60] ,
		\a[61] ,
		_w7077_
	);
	LUT4 #(
		.INIT('hf20d)
	) name7012 (
		_w7055_,
		_w7056_,
		_w7058_,
		_w7077_,
		_w7078_
	);
	LUT4 #(
		.INIT('h153f)
	) name7013 (
		\a[42] ,
		\a[43] ,
		\a[46] ,
		\a[47] ,
		_w7079_
	);
	LUT4 #(
		.INIT('h8000)
	) name7014 (
		\a[42] ,
		\a[43] ,
		\a[46] ,
		\a[47] ,
		_w7080_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7015 (
		\a[42] ,
		\a[43] ,
		\a[46] ,
		\a[47] ,
		_w7081_
	);
	LUT4 #(
		.INIT('h9a30)
	) name7016 (
		\a[27] ,
		\a[44] ,
		\a[45] ,
		\a[62] ,
		_w7082_
	);
	LUT3 #(
		.INIT('h60)
	) name7017 (
		_w7057_,
		_w7081_,
		_w7082_,
		_w7083_
	);
	LUT3 #(
		.INIT('h09)
	) name7018 (
		_w7057_,
		_w7081_,
		_w7082_,
		_w7084_
	);
	LUT3 #(
		.INIT('h96)
	) name7019 (
		_w7057_,
		_w7081_,
		_w7082_,
		_w7085_
	);
	LUT2 #(
		.INIT('h9)
	) name7020 (
		_w7078_,
		_w7085_,
		_w7086_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		\a[41] ,
		\a[48] ,
		_w7087_
	);
	LUT4 #(
		.INIT('h153f)
	) name7022 (
		\a[33] ,
		\a[35] ,
		\a[54] ,
		\a[56] ,
		_w7088_
	);
	LUT2 #(
		.INIT('h8)
	) name7023 (
		\a[35] ,
		\a[56] ,
		_w7089_
	);
	LUT4 #(
		.INIT('h8000)
	) name7024 (
		\a[33] ,
		\a[35] ,
		\a[54] ,
		\a[56] ,
		_w7090_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7025 (
		\a[33] ,
		\a[35] ,
		\a[54] ,
		\a[56] ,
		_w7091_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		\a[36] ,
		\a[53] ,
		_w7092_
	);
	LUT4 #(
		.INIT('h153f)
	) name7027 (
		\a[37] ,
		\a[38] ,
		\a[51] ,
		\a[52] ,
		_w7093_
	);
	LUT4 #(
		.INIT('h8000)
	) name7028 (
		\a[37] ,
		\a[38] ,
		\a[51] ,
		\a[52] ,
		_w7094_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7029 (
		\a[37] ,
		\a[38] ,
		\a[51] ,
		\a[52] ,
		_w7095_
	);
	LUT4 #(
		.INIT('h0660)
	) name7030 (
		_w7087_,
		_w7091_,
		_w7092_,
		_w7095_,
		_w7096_
	);
	LUT4 #(
		.INIT('h9009)
	) name7031 (
		_w7087_,
		_w7091_,
		_w7092_,
		_w7095_,
		_w7097_
	);
	LUT4 #(
		.INIT('h6996)
	) name7032 (
		_w7087_,
		_w7091_,
		_w7092_,
		_w7095_,
		_w7098_
	);
	LUT2 #(
		.INIT('h8)
	) name7033 (
		\a[30] ,
		\a[59] ,
		_w7099_
	);
	LUT4 #(
		.INIT('h153f)
	) name7034 (
		\a[31] ,
		\a[32] ,
		\a[57] ,
		\a[58] ,
		_w7100_
	);
	LUT4 #(
		.INIT('h8000)
	) name7035 (
		\a[31] ,
		\a[32] ,
		\a[57] ,
		\a[58] ,
		_w7101_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7036 (
		\a[31] ,
		\a[32] ,
		\a[57] ,
		\a[58] ,
		_w7102_
	);
	LUT2 #(
		.INIT('h6)
	) name7037 (
		_w7099_,
		_w7102_,
		_w7103_
	);
	LUT2 #(
		.INIT('h6)
	) name7038 (
		_w7098_,
		_w7103_,
		_w7104_
	);
	LUT3 #(
		.INIT('h69)
	) name7039 (
		_w7075_,
		_w7086_,
		_w7104_,
		_w7105_
	);
	LUT3 #(
		.INIT('he0)
	) name7040 (
		_w6999_,
		_w7001_,
		_w7105_,
		_w7106_
	);
	LUT3 #(
		.INIT('h2b)
	) name7041 (
		_w7049_,
		_w7050_,
		_w7051_,
		_w7107_
	);
	LUT3 #(
		.INIT('h23)
	) name7042 (
		_w7021_,
		_w7023_,
		_w7025_,
		_w7108_
	);
	LUT3 #(
		.INIT('hb2)
	) name7043 (
		_w7053_,
		_w7054_,
		_w7060_,
		_w7109_
	);
	LUT3 #(
		.INIT('h96)
	) name7044 (
		_w7107_,
		_w7108_,
		_w7109_,
		_w7110_
	);
	LUT3 #(
		.INIT('he8)
	) name7045 (
		_w6994_,
		_w6995_,
		_w6996_,
		_w7111_
	);
	LUT4 #(
		.INIT('h10f1)
	) name7046 (
		_w6925_,
		_w6927_,
		_w7052_,
		_w7061_,
		_w7112_
	);
	LUT3 #(
		.INIT('h96)
	) name7047 (
		_w7110_,
		_w7111_,
		_w7112_,
		_w7113_
	);
	LUT3 #(
		.INIT('h07)
	) name7048 (
		_w6997_,
		_w6998_,
		_w7105_,
		_w7114_
	);
	LUT4 #(
		.INIT('h001e)
	) name7049 (
		_w6999_,
		_w7001_,
		_w7105_,
		_w7113_,
		_w7115_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name7050 (
		_w6999_,
		_w7001_,
		_w7105_,
		_w7113_,
		_w7116_
	);
	LUT3 #(
		.INIT('h32)
	) name7051 (
		_w7034_,
		_w7035_,
		_w7041_,
		_w7117_
	);
	LUT3 #(
		.INIT('h0d)
	) name7052 (
		_w6870_,
		_w7031_,
		_w7032_,
		_w7118_
	);
	LUT3 #(
		.INIT('h0d)
	) name7053 (
		_w7006_,
		_w7007_,
		_w7008_,
		_w7119_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		\a[26] ,
		\a[63] ,
		_w7120_
	);
	LUT4 #(
		.INIT('h153f)
	) name7055 (
		\a[39] ,
		\a[40] ,
		\a[49] ,
		\a[50] ,
		_w7121_
	);
	LUT4 #(
		.INIT('h8000)
	) name7056 (
		\a[39] ,
		\a[40] ,
		\a[49] ,
		\a[50] ,
		_w7122_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7057 (
		\a[39] ,
		\a[40] ,
		\a[49] ,
		\a[50] ,
		_w7123_
	);
	LUT2 #(
		.INIT('h6)
	) name7058 (
		_w7120_,
		_w7123_,
		_w7124_
	);
	LUT3 #(
		.INIT('h69)
	) name7059 (
		_w7118_,
		_w7119_,
		_w7124_,
		_w7125_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name7060 (
		_w7014_,
		_w7016_,
		_w7117_,
		_w7125_,
		_w7126_
	);
	LUT3 #(
		.INIT('hb2)
	) name7061 (
		_w7017_,
		_w7026_,
		_w7042_,
		_w7127_
	);
	LUT2 #(
		.INIT('h8)
	) name7062 (
		_w7126_,
		_w7127_,
		_w7128_
	);
	LUT2 #(
		.INIT('h6)
	) name7063 (
		_w7126_,
		_w7127_,
		_w7129_
	);
	LUT4 #(
		.INIT('he800)
	) name7064 (
		_w7044_,
		_w7045_,
		_w7062_,
		_w7129_,
		_w7130_
	);
	LUT4 #(
		.INIT('hab54)
	) name7065 (
		_w7046_,
		_w7047_,
		_w7062_,
		_w7129_,
		_w7131_
	);
	LUT4 #(
		.INIT('he000)
	) name7066 (
		_w6913_,
		_w6915_,
		_w7043_,
		_w7131_,
		_w7132_
	);
	LUT4 #(
		.INIT('h1680)
	) name7067 (
		_w7044_,
		_w7045_,
		_w7062_,
		_w7129_,
		_w7133_
	);
	LUT3 #(
		.INIT('hb0)
	) name7068 (
		_w6915_,
		_w7064_,
		_w7133_,
		_w7134_
	);
	LUT2 #(
		.INIT('h1)
	) name7069 (
		_w7132_,
		_w7134_,
		_w7135_
	);
	LUT4 #(
		.INIT('h001f)
	) name7070 (
		_w6913_,
		_w6915_,
		_w7043_,
		_w7131_,
		_w7136_
	);
	LUT4 #(
		.INIT('h0203)
	) name7071 (
		_w7065_,
		_w7132_,
		_w7134_,
		_w7136_,
		_w7137_
	);
	LUT4 #(
		.INIT('h2322)
	) name7072 (
		_w7003_,
		_w7004_,
		_w7065_,
		_w7068_,
		_w7138_
	);
	LUT3 #(
		.INIT('h60)
	) name7073 (
		_w7116_,
		_w7137_,
		_w7138_,
		_w7139_
	);
	LUT3 #(
		.INIT('h09)
	) name7074 (
		_w7116_,
		_w7137_,
		_w7138_,
		_w7140_
	);
	LUT3 #(
		.INIT('h96)
	) name7075 (
		_w7116_,
		_w7137_,
		_w7138_,
		_w7141_
	);
	LUT4 #(
		.INIT('h0777)
	) name7076 (
		_w6908_,
		_w6980_,
		_w6992_,
		_w7069_,
		_w7142_
	);
	LUT3 #(
		.INIT('hb0)
	) name7077 (
		_w6821_,
		_w6903_,
		_w7142_,
		_w7143_
	);
	LUT4 #(
		.INIT('hef00)
	) name7078 (
		_w6818_,
		_w6820_,
		_w6907_,
		_w7143_,
		_w7144_
	);
	LUT4 #(
		.INIT('hfee0)
	) name7079 (
		_w6908_,
		_w6980_,
		_w6992_,
		_w7069_,
		_w7145_
	);
	LUT3 #(
		.INIT('h9a)
	) name7080 (
		_w7141_,
		_w7144_,
		_w7145_,
		_w7146_
	);
	LUT2 #(
		.INIT('h4)
	) name7081 (
		_w7140_,
		_w7145_,
		_w7147_
	);
	LUT3 #(
		.INIT('h8c)
	) name7082 (
		_w7065_,
		_w7116_,
		_w7136_,
		_w7148_
	);
	LUT2 #(
		.INIT('h2)
	) name7083 (
		_w7135_,
		_w7148_,
		_w7149_
	);
	LUT3 #(
		.INIT('h8e)
	) name7084 (
		_w7110_,
		_w7111_,
		_w7112_,
		_w7150_
	);
	LUT4 #(
		.INIT('he0c0)
	) name7085 (
		\a[27] ,
		\a[44] ,
		\a[45] ,
		\a[62] ,
		_w7151_
	);
	LUT3 #(
		.INIT('h0d)
	) name7086 (
		_w7057_,
		_w7079_,
		_w7080_,
		_w7152_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7087 (
		_w7057_,
		_w7079_,
		_w7080_,
		_w7151_,
		_w7153_
	);
	LUT3 #(
		.INIT('h0d)
	) name7088 (
		_w7087_,
		_w7088_,
		_w7090_,
		_w7154_
	);
	LUT2 #(
		.INIT('h6)
	) name7089 (
		_w7153_,
		_w7154_,
		_w7155_
	);
	LUT3 #(
		.INIT('h0d)
	) name7090 (
		_w7078_,
		_w7083_,
		_w7084_,
		_w7156_
	);
	LUT3 #(
		.INIT('h32)
	) name7091 (
		_w7096_,
		_w7097_,
		_w7103_,
		_w7157_
	);
	LUT3 #(
		.INIT('h69)
	) name7092 (
		_w7155_,
		_w7156_,
		_w7157_,
		_w7158_
	);
	LUT3 #(
		.INIT('hd4)
	) name7093 (
		_w7075_,
		_w7086_,
		_w7104_,
		_w7159_
	);
	LUT2 #(
		.INIT('h8)
	) name7094 (
		_w7158_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h1)
	) name7095 (
		_w7158_,
		_w7159_,
		_w7161_
	);
	LUT2 #(
		.INIT('h6)
	) name7096 (
		_w7158_,
		_w7159_,
		_w7162_
	);
	LUT2 #(
		.INIT('h6)
	) name7097 (
		_w7150_,
		_w7162_,
		_w7163_
	);
	LUT4 #(
		.INIT('h001f)
	) name7098 (
		_w6999_,
		_w7001_,
		_w7105_,
		_w7163_,
		_w7164_
	);
	LUT2 #(
		.INIT('h4)
	) name7099 (
		_w7115_,
		_w7164_,
		_w7165_
	);
	LUT3 #(
		.INIT('h28)
	) name7100 (
		_w7105_,
		_w7150_,
		_w7162_,
		_w7166_
	);
	LUT3 #(
		.INIT('he0)
	) name7101 (
		_w6999_,
		_w7001_,
		_w7166_,
		_w7167_
	);
	LUT3 #(
		.INIT('h14)
	) name7102 (
		_w7113_,
		_w7150_,
		_w7162_,
		_w7168_
	);
	LUT3 #(
		.INIT('hb0)
	) name7103 (
		_w7001_,
		_w7114_,
		_w7168_,
		_w7169_
	);
	LUT2 #(
		.INIT('h1)
	) name7104 (
		_w7167_,
		_w7169_,
		_w7170_
	);
	LUT3 #(
		.INIT('he8)
	) name7105 (
		_w7107_,
		_w7108_,
		_w7109_,
		_w7171_
	);
	LUT3 #(
		.INIT('h0d)
	) name7106 (
		_w7092_,
		_w7093_,
		_w7094_,
		_w7172_
	);
	LUT3 #(
		.INIT('h0d)
	) name7107 (
		_w7099_,
		_w7100_,
		_w7101_,
		_w7173_
	);
	LUT3 #(
		.INIT('h0d)
	) name7108 (
		_w7120_,
		_w7121_,
		_w7122_,
		_w7174_
	);
	LUT3 #(
		.INIT('h96)
	) name7109 (
		_w7172_,
		_w7173_,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('h8)
	) name7110 (
		\a[35] ,
		\a[55] ,
		_w7176_
	);
	LUT4 #(
		.INIT('h153f)
	) name7111 (
		\a[33] ,
		\a[34] ,
		\a[56] ,
		\a[57] ,
		_w7177_
	);
	LUT4 #(
		.INIT('h8000)
	) name7112 (
		\a[33] ,
		\a[34] ,
		\a[56] ,
		\a[57] ,
		_w7178_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7113 (
		\a[33] ,
		\a[34] ,
		\a[56] ,
		\a[57] ,
		_w7179_
	);
	LUT2 #(
		.INIT('h8)
	) name7114 (
		\a[36] ,
		\a[54] ,
		_w7180_
	);
	LUT4 #(
		.INIT('h153f)
	) name7115 (
		\a[37] ,
		\a[38] ,
		\a[52] ,
		\a[53] ,
		_w7181_
	);
	LUT4 #(
		.INIT('h8000)
	) name7116 (
		\a[37] ,
		\a[38] ,
		\a[52] ,
		\a[53] ,
		_w7182_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7117 (
		\a[37] ,
		\a[38] ,
		\a[52] ,
		\a[53] ,
		_w7183_
	);
	LUT4 #(
		.INIT('h0660)
	) name7118 (
		_w7176_,
		_w7179_,
		_w7180_,
		_w7183_,
		_w7184_
	);
	LUT4 #(
		.INIT('h9009)
	) name7119 (
		_w7176_,
		_w7179_,
		_w7180_,
		_w7183_,
		_w7185_
	);
	LUT4 #(
		.INIT('h6996)
	) name7120 (
		_w7176_,
		_w7179_,
		_w7180_,
		_w7183_,
		_w7186_
	);
	LUT2 #(
		.INIT('h8)
	) name7121 (
		\a[42] ,
		\a[48] ,
		_w7187_
	);
	LUT4 #(
		.INIT('h153f)
	) name7122 (
		\a[43] ,
		\a[44] ,
		\a[46] ,
		\a[47] ,
		_w7188_
	);
	LUT4 #(
		.INIT('h8000)
	) name7123 (
		\a[43] ,
		\a[44] ,
		\a[46] ,
		\a[47] ,
		_w7189_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7124 (
		\a[43] ,
		\a[44] ,
		\a[46] ,
		\a[47] ,
		_w7190_
	);
	LUT2 #(
		.INIT('h6)
	) name7125 (
		_w7187_,
		_w7190_,
		_w7191_
	);
	LUT2 #(
		.INIT('h6)
	) name7126 (
		_w7186_,
		_w7191_,
		_w7192_
	);
	LUT2 #(
		.INIT('h8)
	) name7127 (
		_w7175_,
		_w7192_,
		_w7193_
	);
	LUT2 #(
		.INIT('h4)
	) name7128 (
		_w7175_,
		_w7192_,
		_w7194_
	);
	LUT3 #(
		.INIT('h69)
	) name7129 (
		_w7171_,
		_w7175_,
		_w7192_,
		_w7195_
	);
	LUT3 #(
		.INIT('he0)
	) name7130 (
		_w7128_,
		_w7130_,
		_w7195_,
		_w7196_
	);
	LUT4 #(
		.INIT('h1f01)
	) name7131 (
		_w7014_,
		_w7016_,
		_w7117_,
		_w7125_,
		_w7197_
	);
	LUT2 #(
		.INIT('h8)
	) name7132 (
		\a[39] ,
		\a[51] ,
		_w7198_
	);
	LUT4 #(
		.INIT('h153f)
	) name7133 (
		\a[40] ,
		\a[41] ,
		\a[49] ,
		\a[50] ,
		_w7199_
	);
	LUT4 #(
		.INIT('h8000)
	) name7134 (
		\a[40] ,
		\a[41] ,
		\a[49] ,
		\a[50] ,
		_w7200_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7135 (
		\a[40] ,
		\a[41] ,
		\a[49] ,
		\a[50] ,
		_w7201_
	);
	LUT2 #(
		.INIT('h6)
	) name7136 (
		_w7198_,
		_w7201_,
		_w7202_
	);
	LUT4 #(
		.INIT('h00e8)
	) name7137 (
		_w7072_,
		_w7073_,
		_w7074_,
		_w7202_,
		_w7203_
	);
	LUT4 #(
		.INIT('h1700)
	) name7138 (
		_w7072_,
		_w7073_,
		_w7074_,
		_w7202_,
		_w7204_
	);
	LUT3 #(
		.INIT('h8e)
	) name7139 (
		_w7118_,
		_w7119_,
		_w7124_,
		_w7205_
	);
	LUT4 #(
		.INIT('h153f)
	) name7140 (
		\a[28] ,
		\a[29] ,
		\a[60] ,
		\a[61] ,
		_w7206_
	);
	LUT4 #(
		.INIT('h000d)
	) name7141 (
		_w7055_,
		_w7056_,
		_w7058_,
		_w7076_,
		_w7207_
	);
	LUT4 #(
		.INIT('h153f)
	) name7142 (
		\a[31] ,
		\a[32] ,
		\a[58] ,
		\a[59] ,
		_w7208_
	);
	LUT4 #(
		.INIT('h8000)
	) name7143 (
		\a[31] ,
		\a[32] ,
		\a[58] ,
		\a[59] ,
		_w7209_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7144 (
		\a[31] ,
		\a[32] ,
		\a[58] ,
		\a[59] ,
		_w7210_
	);
	LUT2 #(
		.INIT('h8)
	) name7145 (
		\a[30] ,
		\a[60] ,
		_w7211_
	);
	LUT2 #(
		.INIT('h6)
	) name7146 (
		_w7210_,
		_w7211_,
		_w7212_
	);
	LUT2 #(
		.INIT('h8)
	) name7147 (
		\a[27] ,
		\a[63] ,
		_w7213_
	);
	LUT4 #(
		.INIT('h153f)
	) name7148 (
		\a[28] ,
		\a[29] ,
		\a[61] ,
		\a[62] ,
		_w7214_
	);
	LUT4 #(
		.INIT('h8000)
	) name7149 (
		\a[28] ,
		\a[29] ,
		\a[61] ,
		\a[62] ,
		_w7215_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7150 (
		\a[28] ,
		\a[29] ,
		\a[61] ,
		\a[62] ,
		_w7216_
	);
	LUT2 #(
		.INIT('h6)
	) name7151 (
		_w7213_,
		_w7216_,
		_w7217_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name7152 (
		_w7206_,
		_w7207_,
		_w7212_,
		_w7217_,
		_w7218_
	);
	LUT4 #(
		.INIT('h1e00)
	) name7153 (
		_w7203_,
		_w7204_,
		_w7205_,
		_w7218_,
		_w7219_
	);
	LUT4 #(
		.INIT('h00e1)
	) name7154 (
		_w7203_,
		_w7204_,
		_w7205_,
		_w7218_,
		_w7220_
	);
	LUT4 #(
		.INIT('he11e)
	) name7155 (
		_w7203_,
		_w7204_,
		_w7205_,
		_w7218_,
		_w7221_
	);
	LUT2 #(
		.INIT('h9)
	) name7156 (
		_w7197_,
		_w7221_,
		_w7222_
	);
	LUT2 #(
		.INIT('h1)
	) name7157 (
		_w7128_,
		_w7195_,
		_w7223_
	);
	LUT3 #(
		.INIT('h8c)
	) name7158 (
		_w7130_,
		_w7222_,
		_w7223_,
		_w7224_
	);
	LUT4 #(
		.INIT('h1e00)
	) name7159 (
		_w7128_,
		_w7130_,
		_w7195_,
		_w7222_,
		_w7225_
	);
	LUT4 #(
		.INIT('he11e)
	) name7160 (
		_w7128_,
		_w7130_,
		_w7195_,
		_w7222_,
		_w7226_
	);
	LUT3 #(
		.INIT('hb4)
	) name7161 (
		_w7165_,
		_w7170_,
		_w7226_,
		_w7227_
	);
	LUT2 #(
		.INIT('h2)
	) name7162 (
		_w7149_,
		_w7227_,
		_w7228_
	);
	LUT2 #(
		.INIT('h9)
	) name7163 (
		_w7149_,
		_w7227_,
		_w7229_
	);
	LUT4 #(
		.INIT('h45ba)
	) name7164 (
		_w7139_,
		_w7144_,
		_w7147_,
		_w7229_,
		_w7230_
	);
	LUT3 #(
		.INIT('h45)
	) name7165 (
		_w7139_,
		_w7149_,
		_w7227_,
		_w7231_
	);
	LUT3 #(
		.INIT('h45)
	) name7166 (
		_w7203_,
		_w7204_,
		_w7205_,
		_w7232_
	);
	LUT3 #(
		.INIT('h0d)
	) name7167 (
		_w7180_,
		_w7181_,
		_w7182_,
		_w7233_
	);
	LUT3 #(
		.INIT('h0d)
	) name7168 (
		_w7213_,
		_w7214_,
		_w7215_,
		_w7234_
	);
	LUT3 #(
		.INIT('h23)
	) name7169 (
		_w7208_,
		_w7209_,
		_w7211_,
		_w7235_
	);
	LUT3 #(
		.INIT('h96)
	) name7170 (
		_w7233_,
		_w7234_,
		_w7235_,
		_w7236_
	);
	LUT2 #(
		.INIT('h8)
	) name7171 (
		\a[28] ,
		\a[63] ,
		_w7237_
	);
	LUT4 #(
		.INIT('h153f)
	) name7172 (
		\a[40] ,
		\a[41] ,
		\a[50] ,
		\a[51] ,
		_w7238_
	);
	LUT4 #(
		.INIT('h8000)
	) name7173 (
		\a[40] ,
		\a[41] ,
		\a[50] ,
		\a[51] ,
		_w7239_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7174 (
		\a[40] ,
		\a[41] ,
		\a[50] ,
		\a[51] ,
		_w7240_
	);
	LUT4 #(
		.INIT('h153f)
	) name7175 (
		\a[43] ,
		\a[44] ,
		\a[47] ,
		\a[48] ,
		_w7241_
	);
	LUT4 #(
		.INIT('h8000)
	) name7176 (
		\a[43] ,
		\a[44] ,
		\a[47] ,
		\a[48] ,
		_w7242_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7177 (
		\a[43] ,
		\a[44] ,
		\a[47] ,
		\a[48] ,
		_w7243_
	);
	LUT4 #(
		.INIT('h1428)
	) name7178 (
		_w7089_,
		_w7237_,
		_w7240_,
		_w7243_,
		_w7244_
	);
	LUT4 #(
		.INIT('h8241)
	) name7179 (
		_w7089_,
		_w7237_,
		_w7240_,
		_w7243_,
		_w7245_
	);
	LUT4 #(
		.INIT('h6996)
	) name7180 (
		_w7089_,
		_w7237_,
		_w7240_,
		_w7243_,
		_w7246_
	);
	LUT4 #(
		.INIT('h9a30)
	) name7181 (
		\a[29] ,
		\a[45] ,
		\a[46] ,
		\a[62] ,
		_w7247_
	);
	LUT2 #(
		.INIT('h6)
	) name7182 (
		_w7246_,
		_w7247_,
		_w7248_
	);
	LUT2 #(
		.INIT('h2)
	) name7183 (
		_w7236_,
		_w7248_,
		_w7249_
	);
	LUT3 #(
		.INIT('h69)
	) name7184 (
		_w7232_,
		_w7236_,
		_w7248_,
		_w7250_
	);
	LUT4 #(
		.INIT('h17ff)
	) name7185 (
		_w7150_,
		_w7158_,
		_w7159_,
		_w7250_,
		_w7251_
	);
	LUT4 #(
		.INIT('h0017)
	) name7186 (
		_w7150_,
		_w7158_,
		_w7159_,
		_w7250_,
		_w7252_
	);
	LUT4 #(
		.INIT('h31ce)
	) name7187 (
		_w7150_,
		_w7160_,
		_w7161_,
		_w7250_,
		_w7253_
	);
	LUT2 #(
		.INIT('h8)
	) name7188 (
		\a[37] ,
		\a[54] ,
		_w7254_
	);
	LUT4 #(
		.INIT('h153f)
	) name7189 (
		\a[38] ,
		\a[39] ,
		\a[52] ,
		\a[53] ,
		_w7255_
	);
	LUT2 #(
		.INIT('h8)
	) name7190 (
		\a[39] ,
		\a[53] ,
		_w7256_
	);
	LUT4 #(
		.INIT('h8000)
	) name7191 (
		\a[38] ,
		\a[39] ,
		\a[52] ,
		\a[53] ,
		_w7257_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7192 (
		\a[38] ,
		\a[39] ,
		\a[52] ,
		\a[53] ,
		_w7258_
	);
	LUT2 #(
		.INIT('h6)
	) name7193 (
		_w7254_,
		_w7258_,
		_w7259_
	);
	LUT3 #(
		.INIT('h0d)
	) name7194 (
		_w7198_,
		_w7199_,
		_w7200_,
		_w7260_
	);
	LUT2 #(
		.INIT('h8)
	) name7195 (
		\a[31] ,
		\a[60] ,
		_w7261_
	);
	LUT4 #(
		.INIT('h153f)
	) name7196 (
		\a[32] ,
		\a[33] ,
		\a[58] ,
		\a[59] ,
		_w7262_
	);
	LUT4 #(
		.INIT('h8000)
	) name7197 (
		\a[32] ,
		\a[33] ,
		\a[58] ,
		\a[59] ,
		_w7263_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7198 (
		\a[32] ,
		\a[33] ,
		\a[58] ,
		\a[59] ,
		_w7264_
	);
	LUT2 #(
		.INIT('h6)
	) name7199 (
		_w7261_,
		_w7264_,
		_w7265_
	);
	LUT3 #(
		.INIT('h96)
	) name7200 (
		_w7259_,
		_w7260_,
		_w7265_,
		_w7266_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7201 (
		_w7155_,
		_w7156_,
		_w7157_,
		_w7266_,
		_w7267_
	);
	LUT3 #(
		.INIT('h17)
	) name7202 (
		_w7172_,
		_w7173_,
		_w7174_,
		_w7268_
	);
	LUT2 #(
		.INIT('h8)
	) name7203 (
		\a[42] ,
		\a[49] ,
		_w7269_
	);
	LUT4 #(
		.INIT('h153f)
	) name7204 (
		\a[34] ,
		\a[36] ,
		\a[55] ,
		\a[57] ,
		_w7270_
	);
	LUT4 #(
		.INIT('h8000)
	) name7205 (
		\a[34] ,
		\a[36] ,
		\a[55] ,
		\a[57] ,
		_w7271_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7206 (
		\a[34] ,
		\a[36] ,
		\a[55] ,
		\a[57] ,
		_w7272_
	);
	LUT2 #(
		.INIT('h6)
	) name7207 (
		_w7269_,
		_w7272_,
		_w7273_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7208 (
		_w7151_,
		_w7152_,
		_w7154_,
		_w7273_,
		_w7274_
	);
	LUT4 #(
		.INIT('h00d4)
	) name7209 (
		_w7151_,
		_w7152_,
		_w7154_,
		_w7273_,
		_w7275_
	);
	LUT3 #(
		.INIT('ha9)
	) name7210 (
		_w7268_,
		_w7274_,
		_w7275_,
		_w7276_
	);
	LUT4 #(
		.INIT('h00d4)
	) name7211 (
		_w7155_,
		_w7156_,
		_w7157_,
		_w7266_,
		_w7277_
	);
	LUT3 #(
		.INIT('hc9)
	) name7212 (
		_w7267_,
		_w7276_,
		_w7277_,
		_w7278_
	);
	LUT2 #(
		.INIT('h6)
	) name7213 (
		_w7253_,
		_w7278_,
		_w7279_
	);
	LUT3 #(
		.INIT('h0d)
	) name7214 (
		_w7197_,
		_w7219_,
		_w7220_,
		_w7280_
	);
	LUT4 #(
		.INIT('h00e8)
	) name7215 (
		_w7107_,
		_w7108_,
		_w7109_,
		_w7175_,
		_w7281_
	);
	LUT4 #(
		.INIT('h0027)
	) name7216 (
		_w7171_,
		_w7193_,
		_w7194_,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('h8)
	) name7217 (
		\a[30] ,
		\a[61] ,
		_w7283_
	);
	LUT4 #(
		.INIT('h0dff)
	) name7218 (
		_w7187_,
		_w7188_,
		_w7189_,
		_w7283_,
		_w7284_
	);
	LUT4 #(
		.INIT('h000d)
	) name7219 (
		_w7187_,
		_w7188_,
		_w7189_,
		_w7283_,
		_w7285_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7220 (
		_w7187_,
		_w7188_,
		_w7189_,
		_w7283_,
		_w7286_
	);
	LUT3 #(
		.INIT('h0d)
	) name7221 (
		_w7176_,
		_w7177_,
		_w7178_,
		_w7287_
	);
	LUT2 #(
		.INIT('h6)
	) name7222 (
		_w7286_,
		_w7287_,
		_w7288_
	);
	LUT4 #(
		.INIT('hf110)
	) name7223 (
		_w7206_,
		_w7207_,
		_w7212_,
		_w7217_,
		_w7289_
	);
	LUT3 #(
		.INIT('h32)
	) name7224 (
		_w7184_,
		_w7185_,
		_w7191_,
		_w7290_
	);
	LUT3 #(
		.INIT('h69)
	) name7225 (
		_w7288_,
		_w7289_,
		_w7290_,
		_w7291_
	);
	LUT3 #(
		.INIT('h69)
	) name7226 (
		_w7280_,
		_w7282_,
		_w7291_,
		_w7292_
	);
	LUT4 #(
		.INIT('h0e01)
	) name7227 (
		_w7196_,
		_w7224_,
		_w7279_,
		_w7292_,
		_w7293_
	);
	LUT3 #(
		.INIT('h01)
	) name7228 (
		_w7167_,
		_w7169_,
		_w7226_,
		_w7294_
	);
	LUT4 #(
		.INIT('h00dc)
	) name7229 (
		_w7001_,
		_w7113_,
		_w7114_,
		_w7163_,
		_w7295_
	);
	LUT2 #(
		.INIT('h4)
	) name7230 (
		_w7106_,
		_w7295_,
		_w7296_
	);
	LUT4 #(
		.INIT('h10e0)
	) name7231 (
		_w7196_,
		_w7225_,
		_w7279_,
		_w7292_,
		_w7297_
	);
	LUT4 #(
		.INIT('h0001)
	) name7232 (
		_w7293_,
		_w7294_,
		_w7296_,
		_w7297_,
		_w7298_
	);
	LUT4 #(
		.INIT('he11e)
	) name7233 (
		_w7196_,
		_w7225_,
		_w7279_,
		_w7292_,
		_w7299_
	);
	LUT3 #(
		.INIT('h0e)
	) name7234 (
		_w7294_,
		_w7296_,
		_w7299_,
		_w7300_
	);
	LUT4 #(
		.INIT('h0356)
	) name7235 (
		_w7293_,
		_w7294_,
		_w7296_,
		_w7297_,
		_w7301_
	);
	LUT3 #(
		.INIT('hd0)
	) name7236 (
		_w7149_,
		_w7227_,
		_w7301_,
		_w7302_
	);
	LUT4 #(
		.INIT('h4f00)
	) name7237 (
		_w7144_,
		_w7147_,
		_w7231_,
		_w7302_,
		_w7303_
	);
	LUT4 #(
		.INIT('h040f)
	) name7238 (
		_w7144_,
		_w7147_,
		_w7228_,
		_w7231_,
		_w7304_
	);
	LUT3 #(
		.INIT('h32)
	) name7239 (
		_w7301_,
		_w7303_,
		_w7304_,
		_w7305_
	);
	LUT3 #(
		.INIT('h02)
	) name7240 (
		_w7149_,
		_w7227_,
		_w7298_,
		_w7306_
	);
	LUT4 #(
		.INIT('h0045)
	) name7241 (
		_w7139_,
		_w7149_,
		_w7227_,
		_w7298_,
		_w7307_
	);
	LUT4 #(
		.INIT('h040f)
	) name7242 (
		_w7144_,
		_w7147_,
		_w7306_,
		_w7307_,
		_w7308_
	);
	LUT3 #(
		.INIT('h0e)
	) name7243 (
		_w7268_,
		_w7274_,
		_w7275_,
		_w7309_
	);
	LUT3 #(
		.INIT('h0d)
	) name7244 (
		_w7254_,
		_w7255_,
		_w7257_,
		_w7310_
	);
	LUT3 #(
		.INIT('h0d)
	) name7245 (
		_w7261_,
		_w7262_,
		_w7263_,
		_w7311_
	);
	LUT3 #(
		.INIT('h0d)
	) name7246 (
		_w7237_,
		_w7238_,
		_w7239_,
		_w7312_
	);
	LUT3 #(
		.INIT('h96)
	) name7247 (
		_w7310_,
		_w7311_,
		_w7312_,
		_w7313_
	);
	LUT3 #(
		.INIT('h0d)
	) name7248 (
		_w7089_,
		_w7241_,
		_w7242_,
		_w7314_
	);
	LUT3 #(
		.INIT('h0d)
	) name7249 (
		_w7269_,
		_w7270_,
		_w7271_,
		_w7315_
	);
	LUT2 #(
		.INIT('h8)
	) name7250 (
		\a[32] ,
		\a[60] ,
		_w7316_
	);
	LUT4 #(
		.INIT('h153f)
	) name7251 (
		\a[37] ,
		\a[38] ,
		\a[54] ,
		\a[55] ,
		_w7317_
	);
	LUT4 #(
		.INIT('h8000)
	) name7252 (
		\a[37] ,
		\a[38] ,
		\a[54] ,
		\a[55] ,
		_w7318_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7253 (
		\a[37] ,
		\a[38] ,
		\a[54] ,
		\a[55] ,
		_w7319_
	);
	LUT2 #(
		.INIT('h6)
	) name7254 (
		_w7316_,
		_w7319_,
		_w7320_
	);
	LUT3 #(
		.INIT('h69)
	) name7255 (
		_w7314_,
		_w7315_,
		_w7320_,
		_w7321_
	);
	LUT2 #(
		.INIT('h1)
	) name7256 (
		_w7313_,
		_w7321_,
		_w7322_
	);
	LUT2 #(
		.INIT('h6)
	) name7257 (
		_w7313_,
		_w7321_,
		_w7323_
	);
	LUT2 #(
		.INIT('h6)
	) name7258 (
		_w7309_,
		_w7323_,
		_w7324_
	);
	LUT4 #(
		.INIT('hba00)
	) name7259 (
		_w7203_,
		_w7204_,
		_w7205_,
		_w7236_,
		_w7325_
	);
	LUT4 #(
		.INIT('h00ba)
	) name7260 (
		_w7203_,
		_w7204_,
		_w7205_,
		_w7248_,
		_w7326_
	);
	LUT3 #(
		.INIT('h01)
	) name7261 (
		_w7249_,
		_w7325_,
		_w7326_,
		_w7327_
	);
	LUT3 #(
		.INIT('h17)
	) name7262 (
		_w7233_,
		_w7234_,
		_w7235_,
		_w7328_
	);
	LUT3 #(
		.INIT('h4d)
	) name7263 (
		_w7259_,
		_w7260_,
		_w7265_,
		_w7329_
	);
	LUT3 #(
		.INIT('h32)
	) name7264 (
		_w7244_,
		_w7245_,
		_w7247_,
		_w7330_
	);
	LUT3 #(
		.INIT('h69)
	) name7265 (
		_w7328_,
		_w7329_,
		_w7330_,
		_w7331_
	);
	LUT4 #(
		.INIT('hfe01)
	) name7266 (
		_w7249_,
		_w7325_,
		_w7326_,
		_w7331_,
		_w7332_
	);
	LUT2 #(
		.INIT('h6)
	) name7267 (
		_w7324_,
		_w7332_,
		_w7333_
	);
	LUT4 #(
		.INIT('h00ce)
	) name7268 (
		_w7251_,
		_w7252_,
		_w7278_,
		_w7333_,
		_w7334_
	);
	LUT3 #(
		.INIT('hb2)
	) name7269 (
		_w7280_,
		_w7282_,
		_w7291_,
		_w7335_
	);
	LUT3 #(
		.INIT('h54)
	) name7270 (
		_w7267_,
		_w7276_,
		_w7277_,
		_w7336_
	);
	LUT3 #(
		.INIT('hd4)
	) name7271 (
		_w7288_,
		_w7289_,
		_w7290_,
		_w7337_
	);
	LUT4 #(
		.INIT('he0c0)
	) name7272 (
		\a[29] ,
		\a[45] ,
		\a[46] ,
		\a[62] ,
		_w7338_
	);
	LUT4 #(
		.INIT('h153f)
	) name7273 (
		\a[30] ,
		\a[31] ,
		\a[61] ,
		\a[62] ,
		_w7339_
	);
	LUT4 #(
		.INIT('h8000)
	) name7274 (
		\a[30] ,
		\a[31] ,
		\a[61] ,
		\a[62] ,
		_w7340_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7275 (
		\a[30] ,
		\a[31] ,
		\a[61] ,
		\a[62] ,
		_w7341_
	);
	LUT4 #(
		.INIT('h153f)
	) name7276 (
		\a[40] ,
		\a[41] ,
		\a[51] ,
		\a[52] ,
		_w7342_
	);
	LUT4 #(
		.INIT('h8000)
	) name7277 (
		\a[40] ,
		\a[41] ,
		\a[51] ,
		\a[52] ,
		_w7343_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7278 (
		\a[40] ,
		\a[41] ,
		\a[51] ,
		\a[52] ,
		_w7344_
	);
	LUT4 #(
		.INIT('h1428)
	) name7279 (
		_w7256_,
		_w7338_,
		_w7341_,
		_w7344_,
		_w7345_
	);
	LUT4 #(
		.INIT('h8241)
	) name7280 (
		_w7256_,
		_w7338_,
		_w7341_,
		_w7344_,
		_w7346_
	);
	LUT4 #(
		.INIT('h6996)
	) name7281 (
		_w7256_,
		_w7338_,
		_w7341_,
		_w7344_,
		_w7347_
	);
	LUT4 #(
		.INIT('hf807)
	) name7282 (
		_w7284_,
		_w7287_,
		_w7285_,
		_w7347_,
		_w7348_
	);
	LUT2 #(
		.INIT('h8)
	) name7283 (
		\a[43] ,
		\a[49] ,
		_w7349_
	);
	LUT4 #(
		.INIT('h153f)
	) name7284 (
		\a[44] ,
		\a[45] ,
		\a[47] ,
		\a[48] ,
		_w7350_
	);
	LUT4 #(
		.INIT('h8000)
	) name7285 (
		\a[44] ,
		\a[45] ,
		\a[47] ,
		\a[48] ,
		_w7351_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7286 (
		\a[44] ,
		\a[45] ,
		\a[47] ,
		\a[48] ,
		_w7352_
	);
	LUT2 #(
		.INIT('h8)
	) name7287 (
		\a[34] ,
		\a[58] ,
		_w7353_
	);
	LUT4 #(
		.INIT('h153f)
	) name7288 (
		\a[35] ,
		\a[42] ,
		\a[50] ,
		\a[57] ,
		_w7354_
	);
	LUT4 #(
		.INIT('h8000)
	) name7289 (
		\a[35] ,
		\a[42] ,
		\a[50] ,
		\a[57] ,
		_w7355_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7290 (
		\a[35] ,
		\a[42] ,
		\a[50] ,
		\a[57] ,
		_w7356_
	);
	LUT4 #(
		.INIT('h0660)
	) name7291 (
		_w7349_,
		_w7352_,
		_w7353_,
		_w7356_,
		_w7357_
	);
	LUT4 #(
		.INIT('h9009)
	) name7292 (
		_w7349_,
		_w7352_,
		_w7353_,
		_w7356_,
		_w7358_
	);
	LUT4 #(
		.INIT('h6996)
	) name7293 (
		_w7349_,
		_w7352_,
		_w7353_,
		_w7356_,
		_w7359_
	);
	LUT2 #(
		.INIT('h8)
	) name7294 (
		\a[36] ,
		\a[56] ,
		_w7360_
	);
	LUT4 #(
		.INIT('h153f)
	) name7295 (
		\a[29] ,
		\a[33] ,
		\a[59] ,
		\a[63] ,
		_w7361_
	);
	LUT4 #(
		.INIT('h8000)
	) name7296 (
		\a[29] ,
		\a[33] ,
		\a[59] ,
		\a[63] ,
		_w7362_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7297 (
		\a[29] ,
		\a[33] ,
		\a[59] ,
		\a[63] ,
		_w7363_
	);
	LUT2 #(
		.INIT('h6)
	) name7298 (
		_w7360_,
		_w7363_,
		_w7364_
	);
	LUT2 #(
		.INIT('h6)
	) name7299 (
		_w7359_,
		_w7364_,
		_w7365_
	);
	LUT2 #(
		.INIT('h1)
	) name7300 (
		_w7348_,
		_w7365_,
		_w7366_
	);
	LUT2 #(
		.INIT('h8)
	) name7301 (
		_w7348_,
		_w7365_,
		_w7367_
	);
	LUT2 #(
		.INIT('h6)
	) name7302 (
		_w7348_,
		_w7365_,
		_w7368_
	);
	LUT2 #(
		.INIT('h6)
	) name7303 (
		_w7337_,
		_w7368_,
		_w7369_
	);
	LUT2 #(
		.INIT('h8)
	) name7304 (
		_w7336_,
		_w7369_,
		_w7370_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w7336_,
		_w7369_,
		_w7371_
	);
	LUT2 #(
		.INIT('h6)
	) name7306 (
		_w7336_,
		_w7369_,
		_w7372_
	);
	LUT2 #(
		.INIT('h6)
	) name7307 (
		_w7335_,
		_w7372_,
		_w7373_
	);
	LUT4 #(
		.INIT('h3100)
	) name7308 (
		_w7251_,
		_w7252_,
		_w7278_,
		_w7333_,
		_w7374_
	);
	LUT3 #(
		.INIT('hc9)
	) name7309 (
		_w7334_,
		_w7373_,
		_w7374_,
		_w7375_
	);
	LUT4 #(
		.INIT('h011f)
	) name7310 (
		_w7196_,
		_w7225_,
		_w7279_,
		_w7292_,
		_w7376_
	);
	LUT2 #(
		.INIT('h4)
	) name7311 (
		_w7375_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h2)
	) name7312 (
		_w7375_,
		_w7376_,
		_w7378_
	);
	LUT2 #(
		.INIT('h9)
	) name7313 (
		_w7375_,
		_w7376_,
		_w7379_
	);
	LUT3 #(
		.INIT('hb4)
	) name7314 (
		_w7300_,
		_w7308_,
		_w7379_,
		_w7380_
	);
	LUT2 #(
		.INIT('h1)
	) name7315 (
		_w7300_,
		_w7377_,
		_w7381_
	);
	LUT3 #(
		.INIT('h54)
	) name7316 (
		_w7334_,
		_w7373_,
		_w7374_,
		_w7382_
	);
	LUT3 #(
		.INIT('h31)
	) name7317 (
		_w7335_,
		_w7370_,
		_w7371_,
		_w7383_
	);
	LUT3 #(
		.INIT('h17)
	) name7318 (
		_w7310_,
		_w7311_,
		_w7312_,
		_w7384_
	);
	LUT3 #(
		.INIT('h8e)
	) name7319 (
		_w7314_,
		_w7315_,
		_w7320_,
		_w7385_
	);
	LUT3 #(
		.INIT('h32)
	) name7320 (
		_w7357_,
		_w7358_,
		_w7364_,
		_w7386_
	);
	LUT3 #(
		.INIT('h69)
	) name7321 (
		_w7384_,
		_w7385_,
		_w7386_,
		_w7387_
	);
	LUT2 #(
		.INIT('h8)
	) name7322 (
		_w7313_,
		_w7321_,
		_w7388_
	);
	LUT3 #(
		.INIT('h0e)
	) name7323 (
		_w7309_,
		_w7322_,
		_w7388_,
		_w7389_
	);
	LUT4 #(
		.INIT('hf01e)
	) name7324 (
		_w7309_,
		_w7322_,
		_w7387_,
		_w7388_,
		_w7390_
	);
	LUT4 #(
		.INIT('h00a8)
	) name7325 (
		_w7284_,
		_w7285_,
		_w7287_,
		_w7345_,
		_w7391_
	);
	LUT3 #(
		.INIT('h32)
	) name7326 (
		_w7353_,
		_w7354_,
		_w7355_,
		_w7392_
	);
	LUT3 #(
		.INIT('h0d)
	) name7327 (
		_w7349_,
		_w7350_,
		_w7351_,
		_w7393_
	);
	LUT3 #(
		.INIT('h0d)
	) name7328 (
		_w7256_,
		_w7342_,
		_w7343_,
		_w7394_
	);
	LUT3 #(
		.INIT('h69)
	) name7329 (
		_w7392_,
		_w7393_,
		_w7394_,
		_w7395_
	);
	LUT3 #(
		.INIT('h32)
	) name7330 (
		_w7360_,
		_w7361_,
		_w7362_,
		_w7396_
	);
	LUT3 #(
		.INIT('h0d)
	) name7331 (
		_w7316_,
		_w7317_,
		_w7318_,
		_w7397_
	);
	LUT3 #(
		.INIT('h0d)
	) name7332 (
		_w7338_,
		_w7339_,
		_w7340_,
		_w7398_
	);
	LUT3 #(
		.INIT('h69)
	) name7333 (
		_w7396_,
		_w7397_,
		_w7398_,
		_w7399_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name7334 (
		_w7346_,
		_w7391_,
		_w7395_,
		_w7399_,
		_w7400_
	);
	LUT2 #(
		.INIT('h6)
	) name7335 (
		_w7390_,
		_w7400_,
		_w7401_
	);
	LUT4 #(
		.INIT('he800)
	) name7336 (
		_w7335_,
		_w7336_,
		_w7369_,
		_w7401_,
		_w7402_
	);
	LUT4 #(
		.INIT('h7007)
	) name7337 (
		_w7336_,
		_w7369_,
		_w7390_,
		_w7400_,
		_w7403_
	);
	LUT3 #(
		.INIT('h70)
	) name7338 (
		_w7335_,
		_w7372_,
		_w7403_,
		_w7404_
	);
	LUT4 #(
		.INIT('hf660)
	) name7339 (
		_w7309_,
		_w7323_,
		_w7327_,
		_w7331_,
		_w7405_
	);
	LUT2 #(
		.INIT('h8)
	) name7340 (
		\a[30] ,
		\a[63] ,
		_w7406_
	);
	LUT4 #(
		.INIT('h153f)
	) name7341 (
		\a[32] ,
		\a[33] ,
		\a[60] ,
		\a[61] ,
		_w7407_
	);
	LUT4 #(
		.INIT('h8000)
	) name7342 (
		\a[32] ,
		\a[33] ,
		\a[60] ,
		\a[61] ,
		_w7408_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7343 (
		\a[32] ,
		\a[33] ,
		\a[60] ,
		\a[61] ,
		_w7409_
	);
	LUT2 #(
		.INIT('h8)
	) name7344 (
		\a[35] ,
		\a[58] ,
		_w7410_
	);
	LUT4 #(
		.INIT('h153f)
	) name7345 (
		\a[36] ,
		\a[39] ,
		\a[54] ,
		\a[57] ,
		_w7411_
	);
	LUT4 #(
		.INIT('h8000)
	) name7346 (
		\a[36] ,
		\a[39] ,
		\a[54] ,
		\a[57] ,
		_w7412_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7347 (
		\a[36] ,
		\a[39] ,
		\a[54] ,
		\a[57] ,
		_w7413_
	);
	LUT4 #(
		.INIT('h0660)
	) name7348 (
		_w7406_,
		_w7409_,
		_w7410_,
		_w7413_,
		_w7414_
	);
	LUT4 #(
		.INIT('h9009)
	) name7349 (
		_w7406_,
		_w7409_,
		_w7410_,
		_w7413_,
		_w7415_
	);
	LUT4 #(
		.INIT('h6996)
	) name7350 (
		_w7406_,
		_w7409_,
		_w7410_,
		_w7413_,
		_w7416_
	);
	LUT2 #(
		.INIT('h8)
	) name7351 (
		\a[34] ,
		\a[59] ,
		_w7417_
	);
	LUT4 #(
		.INIT('h153f)
	) name7352 (
		\a[40] ,
		\a[41] ,
		\a[52] ,
		\a[53] ,
		_w7418_
	);
	LUT4 #(
		.INIT('h8000)
	) name7353 (
		\a[40] ,
		\a[41] ,
		\a[52] ,
		\a[53] ,
		_w7419_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7354 (
		\a[40] ,
		\a[41] ,
		\a[52] ,
		\a[53] ,
		_w7420_
	);
	LUT2 #(
		.INIT('h6)
	) name7355 (
		_w7417_,
		_w7420_,
		_w7421_
	);
	LUT2 #(
		.INIT('h8)
	) name7356 (
		\a[37] ,
		\a[56] ,
		_w7422_
	);
	LUT4 #(
		.INIT('h153f)
	) name7357 (
		\a[38] ,
		\a[45] ,
		\a[48] ,
		\a[55] ,
		_w7423_
	);
	LUT4 #(
		.INIT('h8000)
	) name7358 (
		\a[38] ,
		\a[45] ,
		\a[48] ,
		\a[55] ,
		_w7424_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7359 (
		\a[38] ,
		\a[45] ,
		\a[48] ,
		\a[55] ,
		_w7425_
	);
	LUT2 #(
		.INIT('h8)
	) name7360 (
		\a[42] ,
		\a[51] ,
		_w7426_
	);
	LUT4 #(
		.INIT('h153f)
	) name7361 (
		\a[43] ,
		\a[44] ,
		\a[49] ,
		\a[50] ,
		_w7427_
	);
	LUT4 #(
		.INIT('h8000)
	) name7362 (
		\a[43] ,
		\a[44] ,
		\a[49] ,
		\a[50] ,
		_w7428_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7363 (
		\a[43] ,
		\a[44] ,
		\a[49] ,
		\a[50] ,
		_w7429_
	);
	LUT4 #(
		.INIT('h0660)
	) name7364 (
		_w7422_,
		_w7425_,
		_w7426_,
		_w7429_,
		_w7430_
	);
	LUT4 #(
		.INIT('h9009)
	) name7365 (
		_w7422_,
		_w7425_,
		_w7426_,
		_w7429_,
		_w7431_
	);
	LUT4 #(
		.INIT('h6996)
	) name7366 (
		_w7422_,
		_w7425_,
		_w7426_,
		_w7429_,
		_w7432_
	);
	LUT4 #(
		.INIT('h9a30)
	) name7367 (
		\a[31] ,
		\a[46] ,
		\a[47] ,
		\a[62] ,
		_w7433_
	);
	LUT4 #(
		.INIT('h0660)
	) name7368 (
		_w7416_,
		_w7421_,
		_w7432_,
		_w7433_,
		_w7434_
	);
	LUT4 #(
		.INIT('h6996)
	) name7369 (
		_w7416_,
		_w7421_,
		_w7432_,
		_w7433_,
		_w7435_
	);
	LUT4 #(
		.INIT('hb200)
	) name7370 (
		_w7328_,
		_w7329_,
		_w7330_,
		_w7435_,
		_w7436_
	);
	LUT4 #(
		.INIT('h4db2)
	) name7371 (
		_w7328_,
		_w7329_,
		_w7330_,
		_w7435_,
		_w7437_
	);
	LUT4 #(
		.INIT('he800)
	) name7372 (
		_w7337_,
		_w7348_,
		_w7365_,
		_w7437_,
		_w7438_
	);
	LUT4 #(
		.INIT('h0017)
	) name7373 (
		_w7337_,
		_w7348_,
		_w7365_,
		_w7437_,
		_w7439_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7374 (
		_w7337_,
		_w7366_,
		_w7367_,
		_w7437_,
		_w7440_
	);
	LUT2 #(
		.INIT('h6)
	) name7375 (
		_w7405_,
		_w7440_,
		_w7441_
	);
	LUT3 #(
		.INIT('h10)
	) name7376 (
		_w7402_,
		_w7404_,
		_w7441_,
		_w7442_
	);
	LUT3 #(
		.INIT('h41)
	) name7377 (
		_w7401_,
		_w7405_,
		_w7440_,
		_w7443_
	);
	LUT3 #(
		.INIT('h82)
	) name7378 (
		_w7401_,
		_w7405_,
		_w7440_,
		_w7444_
	);
	LUT3 #(
		.INIT('h27)
	) name7379 (
		_w7383_,
		_w7443_,
		_w7444_,
		_w7445_
	);
	LUT3 #(
		.INIT('h20)
	) name7380 (
		_w7382_,
		_w7442_,
		_w7445_,
		_w7446_
	);
	LUT3 #(
		.INIT('h45)
	) name7381 (
		_w7382_,
		_w7442_,
		_w7445_,
		_w7447_
	);
	LUT3 #(
		.INIT('h9a)
	) name7382 (
		_w7382_,
		_w7442_,
		_w7445_,
		_w7448_
	);
	LUT4 #(
		.INIT('h13ec)
	) name7383 (
		_w7308_,
		_w7378_,
		_w7381_,
		_w7448_,
		_w7449_
	);
	LUT2 #(
		.INIT('h1)
	) name7384 (
		_w7378_,
		_w7446_,
		_w7450_
	);
	LUT3 #(
		.INIT('h90)
	) name7385 (
		_w7309_,
		_w7323_,
		_w7331_,
		_w7451_
	);
	LUT3 #(
		.INIT('h60)
	) name7386 (
		_w7309_,
		_w7323_,
		_w7331_,
		_w7452_
	);
	LUT3 #(
		.INIT('h27)
	) name7387 (
		_w7327_,
		_w7451_,
		_w7452_,
		_w7453_
	);
	LUT3 #(
		.INIT('h07)
	) name7388 (
		_w7324_,
		_w7327_,
		_w7438_,
		_w7454_
	);
	LUT3 #(
		.INIT('h2b)
	) name7389 (
		_w7396_,
		_w7397_,
		_w7398_,
		_w7455_
	);
	LUT3 #(
		.INIT('h2b)
	) name7390 (
		_w7392_,
		_w7393_,
		_w7394_,
		_w7456_
	);
	LUT3 #(
		.INIT('h32)
	) name7391 (
		_w7414_,
		_w7415_,
		_w7421_,
		_w7457_
	);
	LUT3 #(
		.INIT('h96)
	) name7392 (
		_w7455_,
		_w7456_,
		_w7457_,
		_w7458_
	);
	LUT4 #(
		.INIT('h011f)
	) name7393 (
		_w7346_,
		_w7391_,
		_w7395_,
		_w7399_,
		_w7459_
	);
	LUT2 #(
		.INIT('h8)
	) name7394 (
		_w7458_,
		_w7459_,
		_w7460_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name7395 (
		_w7434_,
		_w7436_,
		_w7458_,
		_w7459_,
		_w7461_
	);
	LUT4 #(
		.INIT('he11e)
	) name7396 (
		_w7434_,
		_w7436_,
		_w7458_,
		_w7459_,
		_w7462_
	);
	LUT4 #(
		.INIT('h00ea)
	) name7397 (
		_w7439_,
		_w7453_,
		_w7454_,
		_w7462_,
		_w7463_
	);
	LUT2 #(
		.INIT('h4)
	) name7398 (
		_w7439_,
		_w7462_,
		_w7464_
	);
	LUT3 #(
		.INIT('h70)
	) name7399 (
		_w7453_,
		_w7454_,
		_w7464_,
		_w7465_
	);
	LUT3 #(
		.INIT('hb2)
	) name7400 (
		_w7384_,
		_w7385_,
		_w7386_,
		_w7466_
	);
	LUT2 #(
		.INIT('h8)
	) name7401 (
		\a[36] ,
		\a[58] ,
		_w7467_
	);
	LUT4 #(
		.INIT('h153f)
	) name7402 (
		\a[43] ,
		\a[44] ,
		\a[50] ,
		\a[51] ,
		_w7468_
	);
	LUT4 #(
		.INIT('h8000)
	) name7403 (
		\a[43] ,
		\a[44] ,
		\a[50] ,
		\a[51] ,
		_w7469_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7404 (
		\a[43] ,
		\a[44] ,
		\a[50] ,
		\a[51] ,
		_w7470_
	);
	LUT2 #(
		.INIT('h8)
	) name7405 (
		\a[40] ,
		\a[54] ,
		_w7471_
	);
	LUT4 #(
		.INIT('h153f)
	) name7406 (
		\a[41] ,
		\a[42] ,
		\a[52] ,
		\a[53] ,
		_w7472_
	);
	LUT2 #(
		.INIT('h8)
	) name7407 (
		\a[42] ,
		\a[53] ,
		_w7473_
	);
	LUT4 #(
		.INIT('h8000)
	) name7408 (
		\a[41] ,
		\a[42] ,
		\a[52] ,
		\a[53] ,
		_w7474_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7409 (
		\a[41] ,
		\a[42] ,
		\a[52] ,
		\a[53] ,
		_w7475_
	);
	LUT4 #(
		.INIT('h0660)
	) name7410 (
		_w7467_,
		_w7470_,
		_w7471_,
		_w7475_,
		_w7476_
	);
	LUT4 #(
		.INIT('h9009)
	) name7411 (
		_w7467_,
		_w7470_,
		_w7471_,
		_w7475_,
		_w7477_
	);
	LUT4 #(
		.INIT('h6996)
	) name7412 (
		_w7467_,
		_w7470_,
		_w7471_,
		_w7475_,
		_w7478_
	);
	LUT2 #(
		.INIT('h8)
	) name7413 (
		\a[45] ,
		\a[49] ,
		_w7479_
	);
	LUT4 #(
		.INIT('h153f)
	) name7414 (
		\a[38] ,
		\a[46] ,
		\a[48] ,
		\a[56] ,
		_w7480_
	);
	LUT4 #(
		.INIT('h8000)
	) name7415 (
		\a[38] ,
		\a[46] ,
		\a[48] ,
		\a[56] ,
		_w7481_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7416 (
		\a[38] ,
		\a[46] ,
		\a[48] ,
		\a[56] ,
		_w7482_
	);
	LUT2 #(
		.INIT('h6)
	) name7417 (
		_w7479_,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h6)
	) name7418 (
		_w7478_,
		_w7483_,
		_w7484_
	);
	LUT4 #(
		.INIT('h153f)
	) name7419 (
		\a[33] ,
		\a[35] ,
		\a[59] ,
		\a[61] ,
		_w7485_
	);
	LUT4 #(
		.INIT('h8000)
	) name7420 (
		\a[33] ,
		\a[35] ,
		\a[59] ,
		\a[61] ,
		_w7486_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7421 (
		\a[33] ,
		\a[35] ,
		\a[59] ,
		\a[61] ,
		_w7487_
	);
	LUT2 #(
		.INIT('h6)
	) name7422 (
		_w4382_,
		_w7487_,
		_w7488_
	);
	LUT3 #(
		.INIT('h0d)
	) name7423 (
		_w7426_,
		_w7427_,
		_w7428_,
		_w7489_
	);
	LUT2 #(
		.INIT('h8)
	) name7424 (
		\a[37] ,
		\a[57] ,
		_w7490_
	);
	LUT4 #(
		.INIT('h153f)
	) name7425 (
		\a[34] ,
		\a[39] ,
		\a[55] ,
		\a[60] ,
		_w7491_
	);
	LUT4 #(
		.INIT('h8000)
	) name7426 (
		\a[34] ,
		\a[39] ,
		\a[55] ,
		\a[60] ,
		_w7492_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7427 (
		\a[34] ,
		\a[39] ,
		\a[55] ,
		\a[60] ,
		_w7493_
	);
	LUT2 #(
		.INIT('h6)
	) name7428 (
		_w7490_,
		_w7493_,
		_w7494_
	);
	LUT3 #(
		.INIT('h69)
	) name7429 (
		_w7488_,
		_w7489_,
		_w7494_,
		_w7495_
	);
	LUT3 #(
		.INIT('h13)
	) name7430 (
		\a[31] ,
		\a[46] ,
		\a[62] ,
		_w7496_
	);
	LUT3 #(
		.INIT('h80)
	) name7431 (
		\a[31] ,
		\a[47] ,
		\a[63] ,
		_w7497_
	);
	LUT2 #(
		.INIT('h4)
	) name7432 (
		_w7496_,
		_w7497_,
		_w7498_
	);
	LUT4 #(
		.INIT('he0c0)
	) name7433 (
		\a[31] ,
		\a[46] ,
		\a[47] ,
		\a[62] ,
		_w7499_
	);
	LUT2 #(
		.INIT('h1)
	) name7434 (
		_w5995_,
		_w7499_,
		_w7500_
	);
	LUT3 #(
		.INIT('hc6)
	) name7435 (
		\a[47] ,
		_w5995_,
		_w7496_,
		_w7501_
	);
	LUT3 #(
		.INIT('h0d)
	) name7436 (
		_w7422_,
		_w7423_,
		_w7424_,
		_w7502_
	);
	LUT2 #(
		.INIT('h6)
	) name7437 (
		_w7501_,
		_w7502_,
		_w7503_
	);
	LUT3 #(
		.INIT('h32)
	) name7438 (
		_w7430_,
		_w7431_,
		_w7433_,
		_w7504_
	);
	LUT3 #(
		.INIT('h0d)
	) name7439 (
		_w7410_,
		_w7411_,
		_w7412_,
		_w7505_
	);
	LUT3 #(
		.INIT('h0d)
	) name7440 (
		_w7406_,
		_w7407_,
		_w7408_,
		_w7506_
	);
	LUT3 #(
		.INIT('h0d)
	) name7441 (
		_w7417_,
		_w7418_,
		_w7419_,
		_w7507_
	);
	LUT3 #(
		.INIT('h96)
	) name7442 (
		_w7505_,
		_w7506_,
		_w7507_,
		_w7508_
	);
	LUT3 #(
		.INIT('h96)
	) name7443 (
		_w7503_,
		_w7504_,
		_w7508_,
		_w7509_
	);
	LUT4 #(
		.INIT('h9600)
	) name7444 (
		_w7466_,
		_w7484_,
		_w7495_,
		_w7509_,
		_w7510_
	);
	LUT4 #(
		.INIT('h1700)
	) name7445 (
		_w7387_,
		_w7389_,
		_w7400_,
		_w7510_,
		_w7511_
	);
	LUT4 #(
		.INIT('h0096)
	) name7446 (
		_w7466_,
		_w7484_,
		_w7495_,
		_w7509_,
		_w7512_
	);
	LUT4 #(
		.INIT('he800)
	) name7447 (
		_w7387_,
		_w7389_,
		_w7400_,
		_w7512_,
		_w7513_
	);
	LUT4 #(
		.INIT('h6900)
	) name7448 (
		_w7466_,
		_w7484_,
		_w7495_,
		_w7509_,
		_w7514_
	);
	LUT4 #(
		.INIT('he800)
	) name7449 (
		_w7387_,
		_w7389_,
		_w7400_,
		_w7514_,
		_w7515_
	);
	LUT4 #(
		.INIT('h0069)
	) name7450 (
		_w7466_,
		_w7484_,
		_w7495_,
		_w7509_,
		_w7516_
	);
	LUT4 #(
		.INIT('h1700)
	) name7451 (
		_w7387_,
		_w7389_,
		_w7400_,
		_w7516_,
		_w7517_
	);
	LUT4 #(
		.INIT('h0001)
	) name7452 (
		_w7511_,
		_w7513_,
		_w7515_,
		_w7517_,
		_w7518_
	);
	LUT3 #(
		.INIT('he1)
	) name7453 (
		_w7463_,
		_w7465_,
		_w7518_,
		_w7519_
	);
	LUT3 #(
		.INIT('h45)
	) name7454 (
		_w7402_,
		_w7404_,
		_w7441_,
		_w7520_
	);
	LUT2 #(
		.INIT('h4)
	) name7455 (
		_w7519_,
		_w7520_,
		_w7521_
	);
	LUT2 #(
		.INIT('h2)
	) name7456 (
		_w7519_,
		_w7520_,
		_w7522_
	);
	LUT2 #(
		.INIT('h9)
	) name7457 (
		_w7519_,
		_w7520_,
		_w7523_
	);
	LUT2 #(
		.INIT('h9)
	) name7458 (
		_w7447_,
		_w7523_,
		_w7524_
	);
	LUT4 #(
		.INIT('h8f00)
	) name7459 (
		_w7308_,
		_w7381_,
		_w7450_,
		_w7524_,
		_w7525_
	);
	LUT2 #(
		.INIT('hc)
	) name7460 (
		_w7447_,
		_w7523_,
		_w7526_
	);
	LUT4 #(
		.INIT('h7000)
	) name7461 (
		_w7308_,
		_w7381_,
		_w7450_,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('he)
	) name7462 (
		_w7525_,
		_w7527_,
		_w7528_
	);
	LUT4 #(
		.INIT('he800)
	) name7463 (
		_w7387_,
		_w7389_,
		_w7400_,
		_w7509_,
		_w7529_
	);
	LUT3 #(
		.INIT('h17)
	) name7464 (
		_w7466_,
		_w7484_,
		_w7495_,
		_w7530_
	);
	LUT3 #(
		.INIT('h23)
	) name7465 (
		_w7498_,
		_w7500_,
		_w7502_,
		_w7531_
	);
	LUT2 #(
		.INIT('h8)
	) name7466 (
		\a[36] ,
		\a[60] ,
		_w7532_
	);
	LUT4 #(
		.INIT('h8000)
	) name7467 (
		\a[35] ,
		\a[36] ,
		\a[59] ,
		\a[60] ,
		_w7533_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7468 (
		\a[35] ,
		\a[36] ,
		\a[59] ,
		\a[60] ,
		_w7534_
	);
	LUT4 #(
		.INIT('hcd32)
	) name7469 (
		_w7479_,
		_w7480_,
		_w7481_,
		_w7534_,
		_w7535_
	);
	LUT4 #(
		.INIT('h00dc)
	) name7470 (
		_w7498_,
		_w7500_,
		_w7502_,
		_w7535_,
		_w7536_
	);
	LUT4 #(
		.INIT('h2300)
	) name7471 (
		_w7498_,
		_w7500_,
		_w7502_,
		_w7535_,
		_w7537_
	);
	LUT4 #(
		.INIT('hdc23)
	) name7472 (
		_w7498_,
		_w7500_,
		_w7502_,
		_w7535_,
		_w7538_
	);
	LUT3 #(
		.INIT('h17)
	) name7473 (
		_w7505_,
		_w7506_,
		_w7507_,
		_w7539_
	);
	LUT2 #(
		.INIT('h6)
	) name7474 (
		_w7538_,
		_w7539_,
		_w7540_
	);
	LUT3 #(
		.INIT('h4d)
	) name7475 (
		_w7503_,
		_w7504_,
		_w7508_,
		_w7541_
	);
	LUT2 #(
		.INIT('h6)
	) name7476 (
		_w7540_,
		_w7541_,
		_w7542_
	);
	LUT2 #(
		.INIT('h9)
	) name7477 (
		_w7530_,
		_w7542_,
		_w7543_
	);
	LUT4 #(
		.INIT('h0001)
	) name7478 (
		_w7511_,
		_w7513_,
		_w7529_,
		_w7543_,
		_w7544_
	);
	LUT4 #(
		.INIT('hfe00)
	) name7479 (
		_w7511_,
		_w7513_,
		_w7529_,
		_w7543_,
		_w7545_
	);
	LUT4 #(
		.INIT('h01fe)
	) name7480 (
		_w7511_,
		_w7513_,
		_w7529_,
		_w7543_,
		_w7546_
	);
	LUT4 #(
		.INIT('h011f)
	) name7481 (
		_w7434_,
		_w7436_,
		_w7458_,
		_w7459_,
		_w7547_
	);
	LUT3 #(
		.INIT('h32)
	) name7482 (
		_w7490_,
		_w7491_,
		_w7492_,
		_w7548_
	);
	LUT3 #(
		.INIT('h0d)
	) name7483 (
		_w4382_,
		_w7485_,
		_w7486_,
		_w7549_
	);
	LUT3 #(
		.INIT('h0d)
	) name7484 (
		_w7471_,
		_w7472_,
		_w7474_,
		_w7550_
	);
	LUT3 #(
		.INIT('h69)
	) name7485 (
		_w7548_,
		_w7549_,
		_w7550_,
		_w7551_
	);
	LUT3 #(
		.INIT('h32)
	) name7486 (
		_w7476_,
		_w7477_,
		_w7483_,
		_w7552_
	);
	LUT3 #(
		.INIT('hb2)
	) name7487 (
		_w7488_,
		_w7489_,
		_w7494_,
		_w7553_
	);
	LUT3 #(
		.INIT('h69)
	) name7488 (
		_w7551_,
		_w7552_,
		_w7553_,
		_w7554_
	);
	LUT2 #(
		.INIT('h4)
	) name7489 (
		_w7547_,
		_w7554_,
		_w7555_
	);
	LUT3 #(
		.INIT('h07)
	) name7490 (
		_w7458_,
		_w7459_,
		_w7554_,
		_w7556_
	);
	LUT2 #(
		.INIT('h4)
	) name7491 (
		_w7461_,
		_w7556_,
		_w7557_
	);
	LUT3 #(
		.INIT('he8)
	) name7492 (
		_w7455_,
		_w7456_,
		_w7457_,
		_w7558_
	);
	LUT2 #(
		.INIT('h8)
	) name7493 (
		\a[39] ,
		\a[56] ,
		_w7559_
	);
	LUT4 #(
		.INIT('h153f)
	) name7494 (
		\a[45] ,
		\a[46] ,
		\a[49] ,
		\a[50] ,
		_w7560_
	);
	LUT4 #(
		.INIT('h8000)
	) name7495 (
		\a[45] ,
		\a[46] ,
		\a[49] ,
		\a[50] ,
		_w7561_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7496 (
		\a[45] ,
		\a[46] ,
		\a[49] ,
		\a[50] ,
		_w7562_
	);
	LUT4 #(
		.INIT('h9a30)
	) name7497 (
		\a[33] ,
		\a[47] ,
		\a[48] ,
		\a[62] ,
		_w7563_
	);
	LUT3 #(
		.INIT('h60)
	) name7498 (
		_w7559_,
		_w7562_,
		_w7563_,
		_w7564_
	);
	LUT3 #(
		.INIT('h09)
	) name7499 (
		_w7559_,
		_w7562_,
		_w7563_,
		_w7565_
	);
	LUT3 #(
		.INIT('h96)
	) name7500 (
		_w7559_,
		_w7562_,
		_w7563_,
		_w7566_
	);
	LUT4 #(
		.INIT('h153f)
	) name7501 (
		\a[43] ,
		\a[44] ,
		\a[51] ,
		\a[52] ,
		_w7567_
	);
	LUT2 #(
		.INIT('h8)
	) name7502 (
		\a[44] ,
		\a[52] ,
		_w7568_
	);
	LUT4 #(
		.INIT('h8000)
	) name7503 (
		\a[43] ,
		\a[44] ,
		\a[51] ,
		\a[52] ,
		_w7569_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7504 (
		\a[43] ,
		\a[44] ,
		\a[51] ,
		\a[52] ,
		_w7570_
	);
	LUT2 #(
		.INIT('h6)
	) name7505 (
		_w7473_,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h6)
	) name7506 (
		_w7566_,
		_w7571_,
		_w7572_
	);
	LUT2 #(
		.INIT('h8)
	) name7507 (
		\a[37] ,
		\a[58] ,
		_w7573_
	);
	LUT4 #(
		.INIT('h153f)
	) name7508 (
		\a[38] ,
		\a[40] ,
		\a[55] ,
		\a[57] ,
		_w7574_
	);
	LUT2 #(
		.INIT('h8)
	) name7509 (
		\a[40] ,
		\a[57] ,
		_w7575_
	);
	LUT4 #(
		.INIT('h8000)
	) name7510 (
		\a[38] ,
		\a[40] ,
		\a[55] ,
		\a[57] ,
		_w7576_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7511 (
		\a[38] ,
		\a[40] ,
		\a[55] ,
		\a[57] ,
		_w7577_
	);
	LUT2 #(
		.INIT('h6)
	) name7512 (
		_w7573_,
		_w7577_,
		_w7578_
	);
	LUT3 #(
		.INIT('h0d)
	) name7513 (
		_w7467_,
		_w7468_,
		_w7469_,
		_w7579_
	);
	LUT2 #(
		.INIT('h8)
	) name7514 (
		\a[41] ,
		\a[54] ,
		_w7580_
	);
	LUT4 #(
		.INIT('h153f)
	) name7515 (
		\a[32] ,
		\a[34] ,
		\a[61] ,
		\a[63] ,
		_w7581_
	);
	LUT4 #(
		.INIT('h8000)
	) name7516 (
		\a[32] ,
		\a[34] ,
		\a[61] ,
		\a[63] ,
		_w7582_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7517 (
		\a[32] ,
		\a[34] ,
		\a[61] ,
		\a[63] ,
		_w7583_
	);
	LUT2 #(
		.INIT('h6)
	) name7518 (
		_w7580_,
		_w7583_,
		_w7584_
	);
	LUT3 #(
		.INIT('h96)
	) name7519 (
		_w7578_,
		_w7579_,
		_w7584_,
		_w7585_
	);
	LUT3 #(
		.INIT('h69)
	) name7520 (
		_w7558_,
		_w7572_,
		_w7585_,
		_w7586_
	);
	LUT3 #(
		.INIT('hb0)
	) name7521 (
		_w7461_,
		_w7556_,
		_w7586_,
		_w7587_
	);
	LUT3 #(
		.INIT('h04)
	) name7522 (
		_w7461_,
		_w7556_,
		_w7586_,
		_w7588_
	);
	LUT4 #(
		.INIT('h8228)
	) name7523 (
		_w7554_,
		_w7558_,
		_w7572_,
		_w7585_,
		_w7589_
	);
	LUT2 #(
		.INIT('h4)
	) name7524 (
		_w7547_,
		_w7589_,
		_w7590_
	);
	LUT4 #(
		.INIT('h000b)
	) name7525 (
		_w7555_,
		_w7587_,
		_w7588_,
		_w7590_,
		_w7591_
	);
	LUT2 #(
		.INIT('h1)
	) name7526 (
		_w7546_,
		_w7591_,
		_w7592_
	);
	LUT3 #(
		.INIT('h54)
	) name7527 (
		_w7463_,
		_w7465_,
		_w7518_,
		_w7593_
	);
	LUT2 #(
		.INIT('h8)
	) name7528 (
		_w7546_,
		_w7591_,
		_w7594_
	);
	LUT3 #(
		.INIT('h04)
	) name7529 (
		_w7592_,
		_w7593_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('h6)
	) name7530 (
		_w7546_,
		_w7591_,
		_w7596_
	);
	LUT3 #(
		.INIT('h96)
	) name7531 (
		_w7546_,
		_w7591_,
		_w7593_,
		_w7597_
	);
	LUT4 #(
		.INIT('h0070)
	) name7532 (
		_w7308_,
		_w7381_,
		_w7450_,
		_w7522_,
		_w7598_
	);
	LUT3 #(
		.INIT('h31)
	) name7533 (
		_w7447_,
		_w7521_,
		_w7522_,
		_w7599_
	);
	LUT3 #(
		.INIT('h9a)
	) name7534 (
		_w7597_,
		_w7598_,
		_w7599_,
		_w7600_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name7535 (
		_w7519_,
		_w7520_,
		_w7593_,
		_w7596_,
		_w7601_
	);
	LUT3 #(
		.INIT('hd0)
	) name7536 (
		_w7447_,
		_w7522_,
		_w7601_,
		_w7602_
	);
	LUT4 #(
		.INIT('he0c0)
	) name7537 (
		\a[33] ,
		\a[47] ,
		\a[48] ,
		\a[62] ,
		_w7603_
	);
	LUT3 #(
		.INIT('h0d)
	) name7538 (
		_w7559_,
		_w7560_,
		_w7561_,
		_w7604_
	);
	LUT4 #(
		.INIT('h000d)
	) name7539 (
		_w7559_,
		_w7560_,
		_w7561_,
		_w7603_,
		_w7605_
	);
	LUT4 #(
		.INIT('hf200)
	) name7540 (
		_w7559_,
		_w7560_,
		_w7561_,
		_w7603_,
		_w7606_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7541 (
		_w7559_,
		_w7560_,
		_w7561_,
		_w7603_,
		_w7607_
	);
	LUT3 #(
		.INIT('h0d)
	) name7542 (
		_w7473_,
		_w7567_,
		_w7569_,
		_w7608_
	);
	LUT2 #(
		.INIT('h6)
	) name7543 (
		_w7607_,
		_w7608_,
		_w7609_
	);
	LUT3 #(
		.INIT('h32)
	) name7544 (
		_w7564_,
		_w7565_,
		_w7571_,
		_w7610_
	);
	LUT3 #(
		.INIT('h4d)
	) name7545 (
		_w7578_,
		_w7579_,
		_w7584_,
		_w7611_
	);
	LUT3 #(
		.INIT('h96)
	) name7546 (
		_w7609_,
		_w7610_,
		_w7611_,
		_w7612_
	);
	LUT4 #(
		.INIT('hd400)
	) name7547 (
		_w7530_,
		_w7540_,
		_w7541_,
		_w7612_,
		_w7613_
	);
	LUT3 #(
		.INIT('h07)
	) name7548 (
		_w7540_,
		_w7541_,
		_w7612_,
		_w7614_
	);
	LUT3 #(
		.INIT('hb0)
	) name7549 (
		_w7530_,
		_w7542_,
		_w7614_,
		_w7615_
	);
	LUT2 #(
		.INIT('h8)
	) name7550 (
		\a[41] ,
		\a[55] ,
		_w7616_
	);
	LUT4 #(
		.INIT('h153f)
	) name7551 (
		\a[42] ,
		\a[43] ,
		\a[53] ,
		\a[54] ,
		_w7617_
	);
	LUT2 #(
		.INIT('h8)
	) name7552 (
		\a[43] ,
		\a[54] ,
		_w7618_
	);
	LUT4 #(
		.INIT('h8000)
	) name7553 (
		\a[42] ,
		\a[43] ,
		\a[53] ,
		\a[54] ,
		_w7619_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7554 (
		\a[42] ,
		\a[43] ,
		\a[53] ,
		\a[54] ,
		_w7620_
	);
	LUT2 #(
		.INIT('h8)
	) name7555 (
		\a[33] ,
		\a[63] ,
		_w7621_
	);
	LUT4 #(
		.INIT('h153f)
	) name7556 (
		\a[34] ,
		\a[35] ,
		\a[61] ,
		\a[62] ,
		_w7622_
	);
	LUT4 #(
		.INIT('h8000)
	) name7557 (
		\a[34] ,
		\a[35] ,
		\a[61] ,
		\a[62] ,
		_w7623_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7558 (
		\a[34] ,
		\a[35] ,
		\a[61] ,
		\a[62] ,
		_w7624_
	);
	LUT4 #(
		.INIT('h0660)
	) name7559 (
		_w7616_,
		_w7620_,
		_w7621_,
		_w7624_,
		_w7625_
	);
	LUT4 #(
		.INIT('h6996)
	) name7560 (
		_w7616_,
		_w7620_,
		_w7621_,
		_w7624_,
		_w7626_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7561 (
		_w7548_,
		_w7549_,
		_w7550_,
		_w7626_,
		_w7627_
	);
	LUT4 #(
		.INIT('hd42b)
	) name7562 (
		_w7548_,
		_w7549_,
		_w7550_,
		_w7626_,
		_w7628_
	);
	LUT3 #(
		.INIT('h0d)
	) name7563 (
		_w7573_,
		_w7574_,
		_w7576_,
		_w7629_
	);
	LUT3 #(
		.INIT('h0d)
	) name7564 (
		_w7580_,
		_w7581_,
		_w7582_,
		_w7630_
	);
	LUT3 #(
		.INIT('h01)
	) name7565 (
		_w7479_,
		_w7481_,
		_w7533_,
		_w7631_
	);
	LUT4 #(
		.INIT('h153f)
	) name7566 (
		\a[35] ,
		\a[36] ,
		\a[59] ,
		\a[60] ,
		_w7632_
	);
	LUT3 #(
		.INIT('h0d)
	) name7567 (
		_w7480_,
		_w7533_,
		_w7632_,
		_w7633_
	);
	LUT4 #(
		.INIT('h6966)
	) name7568 (
		_w7629_,
		_w7630_,
		_w7631_,
		_w7633_,
		_w7634_
	);
	LUT3 #(
		.INIT('h54)
	) name7569 (
		_w7536_,
		_w7537_,
		_w7539_,
		_w7635_
	);
	LUT4 #(
		.INIT('h0017)
	) name7570 (
		_w7531_,
		_w7535_,
		_w7539_,
		_w7634_,
		_w7636_
	);
	LUT4 #(
		.INIT('he800)
	) name7571 (
		_w7531_,
		_w7535_,
		_w7539_,
		_w7634_,
		_w7637_
	);
	LUT4 #(
		.INIT('hab54)
	) name7572 (
		_w7536_,
		_w7537_,
		_w7539_,
		_w7634_,
		_w7638_
	);
	LUT2 #(
		.INIT('h6)
	) name7573 (
		_w7628_,
		_w7638_,
		_w7639_
	);
	LUT4 #(
		.INIT('h4f00)
	) name7574 (
		_w7530_,
		_w7542_,
		_w7614_,
		_w7639_,
		_w7640_
	);
	LUT3 #(
		.INIT('h82)
	) name7575 (
		_w7612_,
		_w7628_,
		_w7638_,
		_w7641_
	);
	LUT4 #(
		.INIT('hd400)
	) name7576 (
		_w7530_,
		_w7540_,
		_w7541_,
		_w7641_,
		_w7642_
	);
	LUT4 #(
		.INIT('h00e3)
	) name7577 (
		_w7613_,
		_w7615_,
		_w7639_,
		_w7642_,
		_w7643_
	);
	LUT4 #(
		.INIT('h4114)
	) name7578 (
		_w7554_,
		_w7558_,
		_w7572_,
		_w7585_,
		_w7644_
	);
	LUT4 #(
		.INIT('h00fe)
	) name7579 (
		_w7460_,
		_w7461_,
		_w7586_,
		_w7644_,
		_w7645_
	);
	LUT4 #(
		.INIT('h153f)
	) name7580 (
		\a[37] ,
		\a[40] ,
		\a[56] ,
		\a[59] ,
		_w7646_
	);
	LUT2 #(
		.INIT('h8)
	) name7581 (
		\a[40] ,
		\a[59] ,
		_w7647_
	);
	LUT4 #(
		.INIT('h8000)
	) name7582 (
		\a[37] ,
		\a[40] ,
		\a[56] ,
		\a[59] ,
		_w7648_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7583 (
		\a[37] ,
		\a[40] ,
		\a[56] ,
		\a[59] ,
		_w7649_
	);
	LUT4 #(
		.INIT('h153f)
	) name7584 (
		\a[38] ,
		\a[39] ,
		\a[57] ,
		\a[58] ,
		_w7650_
	);
	LUT4 #(
		.INIT('h8000)
	) name7585 (
		\a[38] ,
		\a[39] ,
		\a[57] ,
		\a[58] ,
		_w7651_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7586 (
		\a[38] ,
		\a[39] ,
		\a[57] ,
		\a[58] ,
		_w7652_
	);
	LUT4 #(
		.INIT('h1248)
	) name7587 (
		_w7532_,
		_w7568_,
		_w7649_,
		_w7652_,
		_w7653_
	);
	LUT4 #(
		.INIT('h8421)
	) name7588 (
		_w7532_,
		_w7568_,
		_w7649_,
		_w7652_,
		_w7654_
	);
	LUT4 #(
		.INIT('h6996)
	) name7589 (
		_w7532_,
		_w7568_,
		_w7649_,
		_w7652_,
		_w7655_
	);
	LUT2 #(
		.INIT('h8)
	) name7590 (
		\a[45] ,
		\a[51] ,
		_w7656_
	);
	LUT4 #(
		.INIT('h153f)
	) name7591 (
		\a[46] ,
		\a[47] ,
		\a[49] ,
		\a[50] ,
		_w7657_
	);
	LUT4 #(
		.INIT('h8000)
	) name7592 (
		\a[46] ,
		\a[47] ,
		\a[49] ,
		\a[50] ,
		_w7658_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7593 (
		\a[46] ,
		\a[47] ,
		\a[49] ,
		\a[50] ,
		_w7659_
	);
	LUT2 #(
		.INIT('h6)
	) name7594 (
		_w7656_,
		_w7659_,
		_w7660_
	);
	LUT2 #(
		.INIT('h6)
	) name7595 (
		_w7655_,
		_w7660_,
		_w7661_
	);
	LUT4 #(
		.INIT('hd400)
	) name7596 (
		_w7551_,
		_w7552_,
		_w7553_,
		_w7661_,
		_w7662_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name7597 (
		_w7551_,
		_w7552_,
		_w7553_,
		_w7661_,
		_w7663_
	);
	LUT4 #(
		.INIT('h0017)
	) name7598 (
		_w7455_,
		_w7456_,
		_w7457_,
		_w7572_,
		_w7664_
	);
	LUT4 #(
		.INIT('he800)
	) name7599 (
		_w7455_,
		_w7456_,
		_w7457_,
		_w7572_,
		_w7665_
	);
	LUT4 #(
		.INIT('h8e00)
	) name7600 (
		_w7558_,
		_w7572_,
		_w7585_,
		_w7663_,
		_w7666_
	);
	LUT4 #(
		.INIT('hc3c9)
	) name7601 (
		_w7585_,
		_w7663_,
		_w7664_,
		_w7665_,
		_w7667_
	);
	LUT3 #(
		.INIT('hb0)
	) name7602 (
		_w7461_,
		_w7556_,
		_w7667_,
		_w7668_
	);
	LUT2 #(
		.INIT('h8)
	) name7603 (
		_w7645_,
		_w7668_,
		_w7669_
	);
	LUT3 #(
		.INIT('h04)
	) name7604 (
		_w7461_,
		_w7556_,
		_w7667_,
		_w7670_
	);
	LUT3 #(
		.INIT('h0e)
	) name7605 (
		_w7645_,
		_w7667_,
		_w7670_,
		_w7671_
	);
	LUT3 #(
		.INIT('hb4)
	) name7606 (
		_w7557_,
		_w7645_,
		_w7667_,
		_w7672_
	);
	LUT2 #(
		.INIT('h6)
	) name7607 (
		_w7643_,
		_w7672_,
		_w7673_
	);
	LUT3 #(
		.INIT('h54)
	) name7608 (
		_w7544_,
		_w7545_,
		_w7591_,
		_w7674_
	);
	LUT2 #(
		.INIT('h1)
	) name7609 (
		_w7673_,
		_w7674_,
		_w7675_
	);
	LUT2 #(
		.INIT('h8)
	) name7610 (
		_w7673_,
		_w7674_,
		_w7676_
	);
	LUT2 #(
		.INIT('h6)
	) name7611 (
		_w7673_,
		_w7674_,
		_w7677_
	);
	LUT4 #(
		.INIT('h45ba)
	) name7612 (
		_w7595_,
		_w7598_,
		_w7602_,
		_w7677_,
		_w7678_
	);
	LUT2 #(
		.INIT('h1)
	) name7613 (
		_w7595_,
		_w7676_,
		_w7679_
	);
	LUT2 #(
		.INIT('h8)
	) name7614 (
		\a[37] ,
		\a[60] ,
		_w7680_
	);
	LUT4 #(
		.INIT('h153f)
	) name7615 (
		\a[38] ,
		\a[39] ,
		\a[58] ,
		\a[59] ,
		_w7681_
	);
	LUT4 #(
		.INIT('h8000)
	) name7616 (
		\a[38] ,
		\a[39] ,
		\a[58] ,
		\a[59] ,
		_w7682_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7617 (
		\a[38] ,
		\a[39] ,
		\a[58] ,
		\a[59] ,
		_w7683_
	);
	LUT2 #(
		.INIT('h8)
	) name7618 (
		\a[41] ,
		\a[56] ,
		_w7684_
	);
	LUT4 #(
		.INIT('h153f)
	) name7619 (
		\a[34] ,
		\a[42] ,
		\a[55] ,
		\a[63] ,
		_w7685_
	);
	LUT4 #(
		.INIT('h8000)
	) name7620 (
		\a[34] ,
		\a[42] ,
		\a[55] ,
		\a[63] ,
		_w7686_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7621 (
		\a[34] ,
		\a[42] ,
		\a[55] ,
		\a[63] ,
		_w7687_
	);
	LUT4 #(
		.INIT('h0660)
	) name7622 (
		_w7680_,
		_w7683_,
		_w7684_,
		_w7687_,
		_w7688_
	);
	LUT4 #(
		.INIT('h9009)
	) name7623 (
		_w7680_,
		_w7683_,
		_w7684_,
		_w7687_,
		_w7689_
	);
	LUT4 #(
		.INIT('h6996)
	) name7624 (
		_w7680_,
		_w7683_,
		_w7684_,
		_w7687_,
		_w7690_
	);
	LUT4 #(
		.INIT('h153f)
	) name7625 (
		\a[44] ,
		\a[45] ,
		\a[52] ,
		\a[53] ,
		_w7691_
	);
	LUT2 #(
		.INIT('h8)
	) name7626 (
		\a[45] ,
		\a[53] ,
		_w7692_
	);
	LUT4 #(
		.INIT('h8000)
	) name7627 (
		\a[44] ,
		\a[45] ,
		\a[52] ,
		\a[53] ,
		_w7693_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7628 (
		\a[44] ,
		\a[45] ,
		\a[52] ,
		\a[53] ,
		_w7694_
	);
	LUT2 #(
		.INIT('h6)
	) name7629 (
		_w7618_,
		_w7694_,
		_w7695_
	);
	LUT2 #(
		.INIT('h6)
	) name7630 (
		_w7690_,
		_w7695_,
		_w7696_
	);
	LUT4 #(
		.INIT('h4d00)
	) name7631 (
		_w7609_,
		_w7610_,
		_w7611_,
		_w7696_,
		_w7697_
	);
	LUT4 #(
		.INIT('h00b2)
	) name7632 (
		_w7609_,
		_w7610_,
		_w7611_,
		_w7696_,
		_w7698_
	);
	LUT4 #(
		.INIT('hb24d)
	) name7633 (
		_w7609_,
		_w7610_,
		_w7611_,
		_w7696_,
		_w7699_
	);
	LUT4 #(
		.INIT('hcd32)
	) name7634 (
		_w7628_,
		_w7636_,
		_w7637_,
		_w7699_,
		_w7700_
	);
	LUT3 #(
		.INIT('h32)
	) name7635 (
		_w7653_,
		_w7654_,
		_w7660_,
		_w7701_
	);
	LUT2 #(
		.INIT('h8)
	) name7636 (
		\a[36] ,
		\a[61] ,
		_w7702_
	);
	LUT4 #(
		.INIT('h0dff)
	) name7637 (
		_w7656_,
		_w7657_,
		_w7658_,
		_w7702_,
		_w7703_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7638 (
		_w7656_,
		_w7657_,
		_w7658_,
		_w7702_,
		_w7704_
	);
	LUT3 #(
		.INIT('h0d)
	) name7639 (
		_w7568_,
		_w7650_,
		_w7651_,
		_w7705_
	);
	LUT2 #(
		.INIT('h6)
	) name7640 (
		_w7704_,
		_w7705_,
		_w7706_
	);
	LUT4 #(
		.INIT('h1711)
	) name7641 (
		_w7629_,
		_w7630_,
		_w7631_,
		_w7633_,
		_w7707_
	);
	LUT3 #(
		.INIT('h69)
	) name7642 (
		_w7701_,
		_w7706_,
		_w7707_,
		_w7708_
	);
	LUT4 #(
		.INIT('h153f)
	) name7643 (
		\a[46] ,
		\a[47] ,
		\a[50] ,
		\a[51] ,
		_w7709_
	);
	LUT4 #(
		.INIT('h8000)
	) name7644 (
		\a[46] ,
		\a[47] ,
		\a[50] ,
		\a[51] ,
		_w7710_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7645 (
		\a[46] ,
		\a[47] ,
		\a[50] ,
		\a[51] ,
		_w7711_
	);
	LUT4 #(
		.INIT('h9a30)
	) name7646 (
		\a[35] ,
		\a[48] ,
		\a[49] ,
		\a[62] ,
		_w7712_
	);
	LUT3 #(
		.INIT('h60)
	) name7647 (
		_w7575_,
		_w7711_,
		_w7712_,
		_w7713_
	);
	LUT3 #(
		.INIT('h96)
	) name7648 (
		_w7575_,
		_w7711_,
		_w7712_,
		_w7714_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7649 (
		_w7603_,
		_w7604_,
		_w7608_,
		_w7714_,
		_w7715_
	);
	LUT4 #(
		.INIT('hba45)
	) name7650 (
		_w7605_,
		_w7606_,
		_w7608_,
		_w7714_,
		_w7716_
	);
	LUT3 #(
		.INIT('h0d)
	) name7651 (
		_w7532_,
		_w7646_,
		_w7648_,
		_w7717_
	);
	LUT3 #(
		.INIT('h0d)
	) name7652 (
		_w7621_,
		_w7622_,
		_w7623_,
		_w7718_
	);
	LUT3 #(
		.INIT('h0d)
	) name7653 (
		_w7616_,
		_w7617_,
		_w7619_,
		_w7719_
	);
	LUT3 #(
		.INIT('h96)
	) name7654 (
		_w7717_,
		_w7718_,
		_w7719_,
		_w7720_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name7655 (
		_w7625_,
		_w7627_,
		_w7716_,
		_w7720_,
		_w7721_
	);
	LUT2 #(
		.INIT('h8)
	) name7656 (
		_w7708_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h1)
	) name7657 (
		_w7708_,
		_w7721_,
		_w7723_
	);
	LUT2 #(
		.INIT('h6)
	) name7658 (
		_w7708_,
		_w7721_,
		_w7724_
	);
	LUT3 #(
		.INIT('he0)
	) name7659 (
		_w7662_,
		_w7666_,
		_w7724_,
		_w7725_
	);
	LUT3 #(
		.INIT('h1e)
	) name7660 (
		_w7662_,
		_w7666_,
		_w7724_,
		_w7726_
	);
	LUT4 #(
		.INIT('he11e)
	) name7661 (
		_w7613_,
		_w7640_,
		_w7700_,
		_w7726_,
		_w7727_
	);
	LUT4 #(
		.INIT('hec00)
	) name7662 (
		_w7643_,
		_w7669_,
		_w7671_,
		_w7727_,
		_w7728_
	);
	LUT4 #(
		.INIT('h0013)
	) name7663 (
		_w7643_,
		_w7669_,
		_w7671_,
		_w7727_,
		_w7729_
	);
	LUT4 #(
		.INIT('h13ec)
	) name7664 (
		_w7643_,
		_w7669_,
		_w7671_,
		_w7727_,
		_w7730_
	);
	LUT3 #(
		.INIT('he0)
	) name7665 (
		_w7673_,
		_w7674_,
		_w7730_,
		_w7731_
	);
	LUT4 #(
		.INIT('h4f00)
	) name7666 (
		_w7598_,
		_w7602_,
		_w7679_,
		_w7731_,
		_w7732_
	);
	LUT4 #(
		.INIT('h040f)
	) name7667 (
		_w7598_,
		_w7602_,
		_w7675_,
		_w7679_,
		_w7733_
	);
	LUT3 #(
		.INIT('h32)
	) name7668 (
		_w7730_,
		_w7732_,
		_w7733_,
		_w7734_
	);
	LUT3 #(
		.INIT('h07)
	) name7669 (
		_w7673_,
		_w7674_,
		_w7728_,
		_w7735_
	);
	LUT3 #(
		.INIT('h01)
	) name7670 (
		_w7673_,
		_w7674_,
		_w7728_,
		_w7736_
	);
	LUT2 #(
		.INIT('h4)
	) name7671 (
		_w7595_,
		_w7735_,
		_w7737_
	);
	LUT4 #(
		.INIT('h040f)
	) name7672 (
		_w7598_,
		_w7602_,
		_w7736_,
		_w7737_,
		_w7738_
	);
	LUT4 #(
		.INIT('h011f)
	) name7673 (
		_w7613_,
		_w7640_,
		_w7700_,
		_w7726_,
		_w7739_
	);
	LUT4 #(
		.INIT('h0f01)
	) name7674 (
		_w7662_,
		_w7666_,
		_w7722_,
		_w7723_,
		_w7740_
	);
	LUT4 #(
		.INIT('he0fe)
	) name7675 (
		_w7625_,
		_w7627_,
		_w7716_,
		_w7720_,
		_w7741_
	);
	LUT4 #(
		.INIT('h153f)
	) name7676 (
		\a[43] ,
		\a[44] ,
		\a[54] ,
		\a[55] ,
		_w7742_
	);
	LUT4 #(
		.INIT('h8000)
	) name7677 (
		\a[43] ,
		\a[44] ,
		\a[54] ,
		\a[55] ,
		_w7743_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7678 (
		\a[43] ,
		\a[44] ,
		\a[54] ,
		\a[55] ,
		_w7744_
	);
	LUT2 #(
		.INIT('h8)
	) name7679 (
		\a[35] ,
		\a[63] ,
		_w7745_
	);
	LUT2 #(
		.INIT('h6)
	) name7680 (
		_w7744_,
		_w7745_,
		_w7746_
	);
	LUT3 #(
		.INIT('h0d)
	) name7681 (
		_w7575_,
		_w7709_,
		_w7710_,
		_w7747_
	);
	LUT2 #(
		.INIT('h8)
	) name7682 (
		\a[38] ,
		\a[60] ,
		_w7748_
	);
	LUT4 #(
		.INIT('h153f)
	) name7683 (
		\a[41] ,
		\a[42] ,
		\a[56] ,
		\a[57] ,
		_w7749_
	);
	LUT4 #(
		.INIT('h8000)
	) name7684 (
		\a[41] ,
		\a[42] ,
		\a[56] ,
		\a[57] ,
		_w7750_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7685 (
		\a[41] ,
		\a[42] ,
		\a[56] ,
		\a[57] ,
		_w7751_
	);
	LUT2 #(
		.INIT('h6)
	) name7686 (
		_w7748_,
		_w7751_,
		_w7752_
	);
	LUT3 #(
		.INIT('h69)
	) name7687 (
		_w7746_,
		_w7747_,
		_w7752_,
		_w7753_
	);
	LUT4 #(
		.INIT('hb200)
	) name7688 (
		_w7701_,
		_w7706_,
		_w7707_,
		_w7753_,
		_w7754_
	);
	LUT4 #(
		.INIT('h004d)
	) name7689 (
		_w7701_,
		_w7706_,
		_w7707_,
		_w7753_,
		_w7755_
	);
	LUT4 #(
		.INIT('h4db2)
	) name7690 (
		_w7701_,
		_w7706_,
		_w7707_,
		_w7753_,
		_w7756_
	);
	LUT2 #(
		.INIT('h6)
	) name7691 (
		_w7741_,
		_w7756_,
		_w7757_
	);
	LUT4 #(
		.INIT('h0017)
	) name7692 (
		_w7628_,
		_w7634_,
		_w7635_,
		_w7697_,
		_w7758_
	);
	LUT3 #(
		.INIT('h17)
	) name7693 (
		_w7717_,
		_w7718_,
		_w7719_,
		_w7759_
	);
	LUT4 #(
		.INIT('h000d)
	) name7694 (
		_w7656_,
		_w7657_,
		_w7658_,
		_w7702_,
		_w7760_
	);
	LUT3 #(
		.INIT('h07)
	) name7695 (
		_w7703_,
		_w7705_,
		_w7760_,
		_w7761_
	);
	LUT3 #(
		.INIT('h32)
	) name7696 (
		_w7688_,
		_w7689_,
		_w7695_,
		_w7762_
	);
	LUT3 #(
		.INIT('h96)
	) name7697 (
		_w7759_,
		_w7761_,
		_w7762_,
		_w7763_
	);
	LUT3 #(
		.INIT('h32)
	) name7698 (
		_w7684_,
		_w7685_,
		_w7686_,
		_w7764_
	);
	LUT3 #(
		.INIT('h0d)
	) name7699 (
		_w7680_,
		_w7681_,
		_w7682_,
		_w7765_
	);
	LUT3 #(
		.INIT('h0d)
	) name7700 (
		_w7618_,
		_w7691_,
		_w7693_,
		_w7766_
	);
	LUT3 #(
		.INIT('h69)
	) name7701 (
		_w7764_,
		_w7765_,
		_w7766_,
		_w7767_
	);
	LUT4 #(
		.INIT('h153f)
	) name7702 (
		\a[36] ,
		\a[37] ,
		\a[61] ,
		\a[62] ,
		_w7768_
	);
	LUT4 #(
		.INIT('h8000)
	) name7703 (
		\a[36] ,
		\a[37] ,
		\a[61] ,
		\a[62] ,
		_w7769_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7704 (
		\a[36] ,
		\a[37] ,
		\a[61] ,
		\a[62] ,
		_w7770_
	);
	LUT4 #(
		.INIT('he0c0)
	) name7705 (
		\a[35] ,
		\a[48] ,
		\a[49] ,
		\a[62] ,
		_w7771_
	);
	LUT2 #(
		.INIT('h8)
	) name7706 (
		_w7770_,
		_w7771_,
		_w7772_
	);
	LUT2 #(
		.INIT('h6)
	) name7707 (
		_w7770_,
		_w7771_,
		_w7773_
	);
	LUT4 #(
		.INIT('h153f)
	) name7708 (
		\a[39] ,
		\a[40] ,
		\a[58] ,
		\a[59] ,
		_w7774_
	);
	LUT4 #(
		.INIT('h8000)
	) name7709 (
		\a[39] ,
		\a[40] ,
		\a[58] ,
		\a[59] ,
		_w7775_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7710 (
		\a[39] ,
		\a[40] ,
		\a[58] ,
		\a[59] ,
		_w7776_
	);
	LUT2 #(
		.INIT('h8)
	) name7711 (
		\a[46] ,
		\a[52] ,
		_w7777_
	);
	LUT4 #(
		.INIT('h153f)
	) name7712 (
		\a[47] ,
		\a[48] ,
		\a[50] ,
		\a[51] ,
		_w7778_
	);
	LUT2 #(
		.INIT('h8)
	) name7713 (
		\a[48] ,
		\a[51] ,
		_w7779_
	);
	LUT4 #(
		.INIT('h8000)
	) name7714 (
		\a[47] ,
		\a[48] ,
		\a[50] ,
		\a[51] ,
		_w7780_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7715 (
		\a[47] ,
		\a[48] ,
		\a[50] ,
		\a[51] ,
		_w7781_
	);
	LUT4 #(
		.INIT('h0660)
	) name7716 (
		_w7692_,
		_w7776_,
		_w7777_,
		_w7781_,
		_w7782_
	);
	LUT4 #(
		.INIT('h9009)
	) name7717 (
		_w7692_,
		_w7776_,
		_w7777_,
		_w7781_,
		_w7783_
	);
	LUT4 #(
		.INIT('h6996)
	) name7718 (
		_w7692_,
		_w7776_,
		_w7777_,
		_w7781_,
		_w7784_
	);
	LUT2 #(
		.INIT('h6)
	) name7719 (
		_w7773_,
		_w7784_,
		_w7785_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name7720 (
		_w7713_,
		_w7715_,
		_w7767_,
		_w7785_,
		_w7786_
	);
	LUT2 #(
		.INIT('h8)
	) name7721 (
		_w7763_,
		_w7786_,
		_w7787_
	);
	LUT2 #(
		.INIT('h1)
	) name7722 (
		_w7763_,
		_w7786_,
		_w7788_
	);
	LUT2 #(
		.INIT('h6)
	) name7723 (
		_w7763_,
		_w7786_,
		_w7789_
	);
	LUT3 #(
		.INIT('he1)
	) name7724 (
		_w7698_,
		_w7758_,
		_w7789_,
		_w7790_
	);
	LUT4 #(
		.INIT('h7007)
	) name7725 (
		_w7708_,
		_w7721_,
		_w7741_,
		_w7756_,
		_w7791_
	);
	LUT4 #(
		.INIT('h1f00)
	) name7726 (
		_w7662_,
		_w7666_,
		_w7724_,
		_w7791_,
		_w7792_
	);
	LUT4 #(
		.INIT('hf04b)
	) name7727 (
		_w7740_,
		_w7757_,
		_w7790_,
		_w7792_,
		_w7793_
	);
	LUT2 #(
		.INIT('h2)
	) name7728 (
		_w7739_,
		_w7793_,
		_w7794_
	);
	LUT2 #(
		.INIT('h4)
	) name7729 (
		_w7739_,
		_w7793_,
		_w7795_
	);
	LUT2 #(
		.INIT('h9)
	) name7730 (
		_w7739_,
		_w7793_,
		_w7796_
	);
	LUT3 #(
		.INIT('hb4)
	) name7731 (
		_w7729_,
		_w7738_,
		_w7796_,
		_w7797_
	);
	LUT2 #(
		.INIT('h1)
	) name7732 (
		_w7729_,
		_w7794_,
		_w7798_
	);
	LUT4 #(
		.INIT('h011f)
	) name7733 (
		_w7722_,
		_w7725_,
		_w7757_,
		_w7790_,
		_w7799_
	);
	LUT3 #(
		.INIT('he8)
	) name7734 (
		_w7759_,
		_w7761_,
		_w7762_,
		_w7800_
	);
	LUT2 #(
		.INIT('h8)
	) name7735 (
		\a[45] ,
		\a[54] ,
		_w7801_
	);
	LUT4 #(
		.INIT('h153f)
	) name7736 (
		\a[46] ,
		\a[47] ,
		\a[52] ,
		\a[53] ,
		_w7802_
	);
	LUT2 #(
		.INIT('h8)
	) name7737 (
		\a[47] ,
		\a[53] ,
		_w7803_
	);
	LUT4 #(
		.INIT('h8000)
	) name7738 (
		\a[46] ,
		\a[47] ,
		\a[52] ,
		\a[53] ,
		_w7804_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7739 (
		\a[46] ,
		\a[47] ,
		\a[52] ,
		\a[53] ,
		_w7805_
	);
	LUT4 #(
		.INIT('h153f)
	) name7740 (
		\a[41] ,
		\a[44] ,
		\a[55] ,
		\a[58] ,
		_w7806_
	);
	LUT4 #(
		.INIT('h8000)
	) name7741 (
		\a[41] ,
		\a[44] ,
		\a[55] ,
		\a[58] ,
		_w7807_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7742 (
		\a[41] ,
		\a[44] ,
		\a[55] ,
		\a[58] ,
		_w7808_
	);
	LUT4 #(
		.INIT('h1428)
	) name7743 (
		_w7647_,
		_w7801_,
		_w7805_,
		_w7808_,
		_w7809_
	);
	LUT4 #(
		.INIT('h8241)
	) name7744 (
		_w7647_,
		_w7801_,
		_w7805_,
		_w7808_,
		_w7810_
	);
	LUT4 #(
		.INIT('h6996)
	) name7745 (
		_w7647_,
		_w7801_,
		_w7805_,
		_w7808_,
		_w7811_
	);
	LUT4 #(
		.INIT('h153f)
	) name7746 (
		\a[42] ,
		\a[43] ,
		\a[56] ,
		\a[57] ,
		_w7812_
	);
	LUT2 #(
		.INIT('h8)
	) name7747 (
		\a[43] ,
		\a[57] ,
		_w7813_
	);
	LUT4 #(
		.INIT('h8000)
	) name7748 (
		\a[42] ,
		\a[43] ,
		\a[56] ,
		\a[57] ,
		_w7814_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7749 (
		\a[42] ,
		\a[43] ,
		\a[56] ,
		\a[57] ,
		_w7815_
	);
	LUT2 #(
		.INIT('h6)
	) name7750 (
		_w7779_,
		_w7815_,
		_w7816_
	);
	LUT2 #(
		.INIT('h6)
	) name7751 (
		_w7811_,
		_w7816_,
		_w7817_
	);
	LUT4 #(
		.INIT('h0017)
	) name7752 (
		_w7759_,
		_w7761_,
		_w7762_,
		_w7817_,
		_w7818_
	);
	LUT4 #(
		.INIT('he800)
	) name7753 (
		_w7759_,
		_w7761_,
		_w7762_,
		_w7817_,
		_w7819_
	);
	LUT4 #(
		.INIT('h17e8)
	) name7754 (
		_w7759_,
		_w7761_,
		_w7762_,
		_w7817_,
		_w7820_
	);
	LUT4 #(
		.INIT('hef0e)
	) name7755 (
		_w7713_,
		_w7715_,
		_w7767_,
		_w7785_,
		_w7821_
	);
	LUT2 #(
		.INIT('h6)
	) name7756 (
		_w7820_,
		_w7821_,
		_w7822_
	);
	LUT3 #(
		.INIT('h0e)
	) name7757 (
		_w7698_,
		_w7758_,
		_w7787_,
		_w7823_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7758 (
		_w7698_,
		_w7758_,
		_w7787_,
		_w7788_,
		_w7824_
	);
	LUT3 #(
		.INIT('h0e)
	) name7759 (
		_w7741_,
		_w7754_,
		_w7755_,
		_w7825_
	);
	LUT3 #(
		.INIT('hb2)
	) name7760 (
		_w7746_,
		_w7747_,
		_w7752_,
		_w7826_
	);
	LUT4 #(
		.INIT('h9a30)
	) name7761 (
		\a[37] ,
		\a[49] ,
		\a[50] ,
		\a[62] ,
		_w7827_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7762 (
		_w7764_,
		_w7765_,
		_w7766_,
		_w7827_,
		_w7828_
	);
	LUT4 #(
		.INIT('h00d4)
	) name7763 (
		_w7764_,
		_w7765_,
		_w7766_,
		_w7827_,
		_w7829_
	);
	LUT4 #(
		.INIT('hd42b)
	) name7764 (
		_w7764_,
		_w7765_,
		_w7766_,
		_w7827_,
		_w7830_
	);
	LUT2 #(
		.INIT('h6)
	) name7765 (
		_w7826_,
		_w7830_,
		_w7831_
	);
	LUT3 #(
		.INIT('h0d)
	) name7766 (
		_w7777_,
		_w7778_,
		_w7780_,
		_w7832_
	);
	LUT3 #(
		.INIT('h0d)
	) name7767 (
		_w7692_,
		_w7774_,
		_w7775_,
		_w7833_
	);
	LUT3 #(
		.INIT('h23)
	) name7768 (
		_w7742_,
		_w7743_,
		_w7745_,
		_w7834_
	);
	LUT3 #(
		.INIT('h96)
	) name7769 (
		_w7832_,
		_w7833_,
		_w7834_,
		_w7835_
	);
	LUT3 #(
		.INIT('h0e)
	) name7770 (
		_w7773_,
		_w7782_,
		_w7783_,
		_w7836_
	);
	LUT2 #(
		.INIT('h4)
	) name7771 (
		_w7835_,
		_w7836_,
		_w7837_
	);
	LUT2 #(
		.INIT('h2)
	) name7772 (
		_w7835_,
		_w7836_,
		_w7838_
	);
	LUT2 #(
		.INIT('h9)
	) name7773 (
		_w7835_,
		_w7836_,
		_w7839_
	);
	LUT3 #(
		.INIT('h23)
	) name7774 (
		_w7768_,
		_w7769_,
		_w7771_,
		_w7840_
	);
	LUT3 #(
		.INIT('h0d)
	) name7775 (
		_w7748_,
		_w7749_,
		_w7750_,
		_w7841_
	);
	LUT2 #(
		.INIT('h1)
	) name7776 (
		_w7840_,
		_w7841_,
		_w7842_
	);
	LUT2 #(
		.INIT('h8)
	) name7777 (
		\a[36] ,
		\a[63] ,
		_w7843_
	);
	LUT4 #(
		.INIT('h153f)
	) name7778 (
		\a[38] ,
		\a[39] ,
		\a[60] ,
		\a[61] ,
		_w7844_
	);
	LUT4 #(
		.INIT('h8000)
	) name7779 (
		\a[38] ,
		\a[39] ,
		\a[60] ,
		\a[61] ,
		_w7845_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7780 (
		\a[38] ,
		\a[39] ,
		\a[60] ,
		\a[61] ,
		_w7846_
	);
	LUT2 #(
		.INIT('h6)
	) name7781 (
		_w7843_,
		_w7846_,
		_w7847_
	);
	LUT4 #(
		.INIT('h000d)
	) name7782 (
		_w7748_,
		_w7749_,
		_w7750_,
		_w7769_,
		_w7848_
	);
	LUT2 #(
		.INIT('h4)
	) name7783 (
		_w7772_,
		_w7848_,
		_w7849_
	);
	LUT3 #(
		.INIT('h36)
	) name7784 (
		_w7842_,
		_w7847_,
		_w7849_,
		_w7850_
	);
	LUT3 #(
		.INIT('h82)
	) name7785 (
		_w7831_,
		_w7839_,
		_w7850_,
		_w7851_
	);
	LUT3 #(
		.INIT('h14)
	) name7786 (
		_w7831_,
		_w7839_,
		_w7850_,
		_w7852_
	);
	LUT3 #(
		.INIT('h69)
	) name7787 (
		_w7831_,
		_w7839_,
		_w7850_,
		_w7853_
	);
	LUT2 #(
		.INIT('h6)
	) name7788 (
		_w7825_,
		_w7853_,
		_w7854_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name7789 (
		_w7763_,
		_w7786_,
		_w7820_,
		_w7821_,
		_w7855_
	);
	LUT4 #(
		.INIT('hf100)
	) name7790 (
		_w7698_,
		_w7758_,
		_w7787_,
		_w7855_,
		_w7856_
	);
	LUT4 #(
		.INIT('hf01e)
	) name7791 (
		_w7822_,
		_w7824_,
		_w7854_,
		_w7856_,
		_w7857_
	);
	LUT2 #(
		.INIT('h9)
	) name7792 (
		_w7799_,
		_w7857_,
		_w7858_
	);
	LUT4 #(
		.INIT('h13ec)
	) name7793 (
		_w7738_,
		_w7795_,
		_w7798_,
		_w7858_,
		_w7859_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7794 (
		_w7739_,
		_w7793_,
		_w7799_,
		_w7857_,
		_w7860_
	);
	LUT4 #(
		.INIT('hcd04)
	) name7795 (
		_w7788_,
		_w7822_,
		_w7823_,
		_w7854_,
		_w7861_
	);
	LUT4 #(
		.INIT('h153f)
	) name7796 (
		\a[48] ,
		\a[49] ,
		\a[51] ,
		\a[52] ,
		_w7862_
	);
	LUT4 #(
		.INIT('h8000)
	) name7797 (
		\a[48] ,
		\a[49] ,
		\a[51] ,
		\a[52] ,
		_w7863_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7798 (
		\a[48] ,
		\a[49] ,
		\a[51] ,
		\a[52] ,
		_w7864_
	);
	LUT2 #(
		.INIT('h6)
	) name7799 (
		_w7803_,
		_w7864_,
		_w7865_
	);
	LUT4 #(
		.INIT('h1700)
	) name7800 (
		_w7832_,
		_w7833_,
		_w7834_,
		_w7865_,
		_w7866_
	);
	LUT4 #(
		.INIT('h00e8)
	) name7801 (
		_w7832_,
		_w7833_,
		_w7834_,
		_w7865_,
		_w7867_
	);
	LUT4 #(
		.INIT('he817)
	) name7802 (
		_w7832_,
		_w7833_,
		_w7834_,
		_w7865_,
		_w7868_
	);
	LUT3 #(
		.INIT('h0e)
	) name7803 (
		_w7840_,
		_w7841_,
		_w7847_,
		_w7869_
	);
	LUT3 #(
		.INIT('hc9)
	) name7804 (
		_w7849_,
		_w7868_,
		_w7869_,
		_w7870_
	);
	LUT4 #(
		.INIT('h0023)
	) name7805 (
		_w7818_,
		_w7819_,
		_w7821_,
		_w7870_,
		_w7871_
	);
	LUT4 #(
		.INIT('he800)
	) name7806 (
		_w7800_,
		_w7817_,
		_w7821_,
		_w7870_,
		_w7872_
	);
	LUT4 #(
		.INIT('h17e8)
	) name7807 (
		_w7800_,
		_w7817_,
		_w7821_,
		_w7870_,
		_w7873_
	);
	LUT3 #(
		.INIT('h0d)
	) name7808 (
		_w7843_,
		_w7844_,
		_w7845_,
		_w7874_
	);
	LUT3 #(
		.INIT('h0d)
	) name7809 (
		_w7801_,
		_w7802_,
		_w7804_,
		_w7875_
	);
	LUT3 #(
		.INIT('h32)
	) name7810 (
		_w7647_,
		_w7806_,
		_w7807_,
		_w7876_
	);
	LUT3 #(
		.INIT('h96)
	) name7811 (
		_w7874_,
		_w7875_,
		_w7876_,
		_w7877_
	);
	LUT3 #(
		.INIT('h32)
	) name7812 (
		_w7809_,
		_w7810_,
		_w7816_,
		_w7878_
	);
	LUT3 #(
		.INIT('h13)
	) name7813 (
		\a[37] ,
		\a[49] ,
		\a[62] ,
		_w7879_
	);
	LUT2 #(
		.INIT('h8)
	) name7814 (
		\a[37] ,
		\a[63] ,
		_w7880_
	);
	LUT3 #(
		.INIT('h80)
	) name7815 (
		\a[37] ,
		\a[50] ,
		\a[63] ,
		_w7881_
	);
	LUT2 #(
		.INIT('h4)
	) name7816 (
		_w7879_,
		_w7881_,
		_w7882_
	);
	LUT4 #(
		.INIT('he0c0)
	) name7817 (
		\a[37] ,
		\a[49] ,
		\a[50] ,
		\a[62] ,
		_w7883_
	);
	LUT2 #(
		.INIT('h1)
	) name7818 (
		_w7880_,
		_w7883_,
		_w7884_
	);
	LUT3 #(
		.INIT('hd2)
	) name7819 (
		\a[50] ,
		_w7879_,
		_w7880_,
		_w7885_
	);
	LUT3 #(
		.INIT('h0d)
	) name7820 (
		_w7779_,
		_w7812_,
		_w7814_,
		_w7886_
	);
	LUT2 #(
		.INIT('h6)
	) name7821 (
		_w7885_,
		_w7886_,
		_w7887_
	);
	LUT3 #(
		.INIT('h69)
	) name7822 (
		_w7877_,
		_w7878_,
		_w7887_,
		_w7888_
	);
	LUT2 #(
		.INIT('h6)
	) name7823 (
		_w7873_,
		_w7888_,
		_w7889_
	);
	LUT2 #(
		.INIT('h8)
	) name7824 (
		\a[38] ,
		\a[62] ,
		_w7890_
	);
	LUT4 #(
		.INIT('h153f)
	) name7825 (
		\a[39] ,
		\a[40] ,
		\a[60] ,
		\a[61] ,
		_w7891_
	);
	LUT4 #(
		.INIT('h8000)
	) name7826 (
		\a[39] ,
		\a[40] ,
		\a[60] ,
		\a[61] ,
		_w7892_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7827 (
		\a[39] ,
		\a[40] ,
		\a[60] ,
		\a[61] ,
		_w7893_
	);
	LUT4 #(
		.INIT('h153f)
	) name7828 (
		\a[44] ,
		\a[45] ,
		\a[55] ,
		\a[56] ,
		_w7894_
	);
	LUT4 #(
		.INIT('h8000)
	) name7829 (
		\a[44] ,
		\a[45] ,
		\a[55] ,
		\a[56] ,
		_w7895_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7830 (
		\a[44] ,
		\a[45] ,
		\a[55] ,
		\a[56] ,
		_w7896_
	);
	LUT4 #(
		.INIT('h1428)
	) name7831 (
		_w7813_,
		_w7890_,
		_w7893_,
		_w7896_,
		_w7897_
	);
	LUT4 #(
		.INIT('h8241)
	) name7832 (
		_w7813_,
		_w7890_,
		_w7893_,
		_w7896_,
		_w7898_
	);
	LUT4 #(
		.INIT('h6996)
	) name7833 (
		_w7813_,
		_w7890_,
		_w7893_,
		_w7896_,
		_w7899_
	);
	LUT2 #(
		.INIT('h8)
	) name7834 (
		\a[46] ,
		\a[54] ,
		_w7900_
	);
	LUT4 #(
		.INIT('h153f)
	) name7835 (
		\a[41] ,
		\a[42] ,
		\a[58] ,
		\a[59] ,
		_w7901_
	);
	LUT2 #(
		.INIT('h8)
	) name7836 (
		\a[42] ,
		\a[59] ,
		_w7902_
	);
	LUT4 #(
		.INIT('h8000)
	) name7837 (
		\a[41] ,
		\a[42] ,
		\a[58] ,
		\a[59] ,
		_w7903_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7838 (
		\a[41] ,
		\a[42] ,
		\a[58] ,
		\a[59] ,
		_w7904_
	);
	LUT2 #(
		.INIT('h6)
	) name7839 (
		_w7900_,
		_w7904_,
		_w7905_
	);
	LUT2 #(
		.INIT('h6)
	) name7840 (
		_w7899_,
		_w7905_,
		_w7906_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7841 (
		_w7826_,
		_w7828_,
		_w7829_,
		_w7906_,
		_w7907_
	);
	LUT4 #(
		.INIT('h0e00)
	) name7842 (
		_w7826_,
		_w7828_,
		_w7829_,
		_w7906_,
		_w7908_
	);
	LUT4 #(
		.INIT('hf10e)
	) name7843 (
		_w7826_,
		_w7828_,
		_w7829_,
		_w7906_,
		_w7909_
	);
	LUT4 #(
		.INIT('hdc23)
	) name7844 (
		_w7837_,
		_w7838_,
		_w7850_,
		_w7909_,
		_w7910_
	);
	LUT4 #(
		.INIT('hec00)
	) name7845 (
		_w7825_,
		_w7851_,
		_w7853_,
		_w7910_,
		_w7911_
	);
	LUT4 #(
		.INIT('h0031)
	) name7846 (
		_w7825_,
		_w7851_,
		_w7852_,
		_w7910_,
		_w7912_
	);
	LUT4 #(
		.INIT('h31ce)
	) name7847 (
		_w7825_,
		_w7851_,
		_w7852_,
		_w7910_,
		_w7913_
	);
	LUT2 #(
		.INIT('h9)
	) name7848 (
		_w7889_,
		_w7913_,
		_w7914_
	);
	LUT2 #(
		.INIT('h4)
	) name7849 (
		_w7861_,
		_w7914_,
		_w7915_
	);
	LUT4 #(
		.INIT('h2dd2)
	) name7850 (
		_w7799_,
		_w7857_,
		_w7861_,
		_w7914_,
		_w7916_
	);
	LUT4 #(
		.INIT('h8f00)
	) name7851 (
		_w7738_,
		_w7798_,
		_w7860_,
		_w7916_,
		_w7917_
	);
	LUT4 #(
		.INIT('hf00f)
	) name7852 (
		_w7799_,
		_w7857_,
		_w7861_,
		_w7914_,
		_w7918_
	);
	LUT4 #(
		.INIT('h7000)
	) name7853 (
		_w7738_,
		_w7798_,
		_w7860_,
		_w7918_,
		_w7919_
	);
	LUT2 #(
		.INIT('he)
	) name7854 (
		_w7917_,
		_w7919_,
		_w7920_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name7855 (
		_w7799_,
		_w7857_,
		_w7861_,
		_w7914_,
		_w7921_
	);
	LUT2 #(
		.INIT('h4)
	) name7856 (
		_w7795_,
		_w7921_,
		_w7922_
	);
	LUT4 #(
		.INIT('h2202)
	) name7857 (
		_w7799_,
		_w7857_,
		_w7861_,
		_w7914_,
		_w7923_
	);
	LUT3 #(
		.INIT('h0e)
	) name7858 (
		_w7889_,
		_w7911_,
		_w7912_,
		_w7924_
	);
	LUT4 #(
		.INIT('h0c0d)
	) name7859 (
		_w7849_,
		_w7866_,
		_w7867_,
		_w7869_,
		_w7925_
	);
	LUT2 #(
		.INIT('h8)
	) name7860 (
		\a[38] ,
		\a[63] ,
		_w7926_
	);
	LUT4 #(
		.INIT('h153f)
	) name7861 (
		\a[46] ,
		\a[47] ,
		\a[54] ,
		\a[55] ,
		_w7927_
	);
	LUT4 #(
		.INIT('h8000)
	) name7862 (
		\a[46] ,
		\a[47] ,
		\a[54] ,
		\a[55] ,
		_w7928_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7863 (
		\a[46] ,
		\a[47] ,
		\a[54] ,
		\a[55] ,
		_w7929_
	);
	LUT4 #(
		.INIT('h153f)
	) name7864 (
		\a[43] ,
		\a[45] ,
		\a[56] ,
		\a[58] ,
		_w7930_
	);
	LUT4 #(
		.INIT('h8000)
	) name7865 (
		\a[43] ,
		\a[45] ,
		\a[56] ,
		\a[58] ,
		_w7931_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7866 (
		\a[43] ,
		\a[45] ,
		\a[56] ,
		\a[58] ,
		_w7932_
	);
	LUT4 #(
		.INIT('h1428)
	) name7867 (
		_w7902_,
		_w7926_,
		_w7929_,
		_w7932_,
		_w7933_
	);
	LUT4 #(
		.INIT('h8241)
	) name7868 (
		_w7902_,
		_w7926_,
		_w7929_,
		_w7932_,
		_w7934_
	);
	LUT4 #(
		.INIT('h6996)
	) name7869 (
		_w7902_,
		_w7926_,
		_w7929_,
		_w7932_,
		_w7935_
	);
	LUT2 #(
		.INIT('h8)
	) name7870 (
		\a[48] ,
		\a[53] ,
		_w7936_
	);
	LUT4 #(
		.INIT('h153f)
	) name7871 (
		\a[44] ,
		\a[49] ,
		\a[52] ,
		\a[57] ,
		_w7937_
	);
	LUT4 #(
		.INIT('h8000)
	) name7872 (
		\a[44] ,
		\a[49] ,
		\a[52] ,
		\a[57] ,
		_w7938_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7873 (
		\a[44] ,
		\a[49] ,
		\a[52] ,
		\a[57] ,
		_w7939_
	);
	LUT2 #(
		.INIT('h6)
	) name7874 (
		_w7936_,
		_w7939_,
		_w7940_
	);
	LUT2 #(
		.INIT('h6)
	) name7875 (
		_w7935_,
		_w7940_,
		_w7941_
	);
	LUT3 #(
		.INIT('h23)
	) name7876 (
		_w7882_,
		_w7884_,
		_w7886_,
		_w7942_
	);
	LUT3 #(
		.INIT('h0d)
	) name7877 (
		_w7803_,
		_w7862_,
		_w7863_,
		_w7943_
	);
	LUT4 #(
		.INIT('h8000)
	) name7878 (
		\a[40] ,
		\a[41] ,
		\a[60] ,
		\a[61] ,
		_w7944_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7879 (
		\a[40] ,
		\a[41] ,
		\a[60] ,
		\a[61] ,
		_w7945_
	);
	LUT4 #(
		.INIT('h9a30)
	) name7880 (
		\a[39] ,
		\a[50] ,
		\a[51] ,
		\a[62] ,
		_w7946_
	);
	LUT3 #(
		.INIT('h6f)
	) name7881 (
		_w7943_,
		_w7945_,
		_w7946_,
		_w7947_
	);
	LUT3 #(
		.INIT('hf9)
	) name7882 (
		_w7943_,
		_w7945_,
		_w7946_,
		_w7948_
	);
	LUT3 #(
		.INIT('h69)
	) name7883 (
		_w7943_,
		_w7945_,
		_w7946_,
		_w7949_
	);
	LUT2 #(
		.INIT('h6)
	) name7884 (
		_w7942_,
		_w7949_,
		_w7950_
	);
	LUT3 #(
		.INIT('h96)
	) name7885 (
		_w7925_,
		_w7941_,
		_w7950_,
		_w7951_
	);
	LUT4 #(
		.INIT('h23ff)
	) name7886 (
		_w7871_,
		_w7872_,
		_w7888_,
		_w7951_,
		_w7952_
	);
	LUT4 #(
		.INIT('h0023)
	) name7887 (
		_w7871_,
		_w7872_,
		_w7888_,
		_w7951_,
		_w7953_
	);
	LUT4 #(
		.INIT('h23dc)
	) name7888 (
		_w7871_,
		_w7872_,
		_w7888_,
		_w7951_,
		_w7954_
	);
	LUT3 #(
		.INIT('h0d)
	) name7889 (
		_w7900_,
		_w7901_,
		_w7903_,
		_w7955_
	);
	LUT3 #(
		.INIT('h0d)
	) name7890 (
		_w7890_,
		_w7891_,
		_w7892_,
		_w7956_
	);
	LUT3 #(
		.INIT('h0d)
	) name7891 (
		_w7813_,
		_w7894_,
		_w7895_,
		_w7957_
	);
	LUT3 #(
		.INIT('h96)
	) name7892 (
		_w7955_,
		_w7956_,
		_w7957_,
		_w7958_
	);
	LUT3 #(
		.INIT('h71)
	) name7893 (
		_w7874_,
		_w7875_,
		_w7876_,
		_w7959_
	);
	LUT3 #(
		.INIT('h32)
	) name7894 (
		_w7897_,
		_w7898_,
		_w7905_,
		_w7960_
	);
	LUT3 #(
		.INIT('h14)
	) name7895 (
		_w7958_,
		_w7959_,
		_w7960_,
		_w7961_
	);
	LUT4 #(
		.INIT('h00b2)
	) name7896 (
		_w7835_,
		_w7836_,
		_w7850_,
		_w7908_,
		_w7962_
	);
	LUT3 #(
		.INIT('h8e)
	) name7897 (
		_w7877_,
		_w7878_,
		_w7887_,
		_w7963_
	);
	LUT2 #(
		.INIT('h4)
	) name7898 (
		_w7907_,
		_w7963_,
		_w7964_
	);
	LUT2 #(
		.INIT('h4)
	) name7899 (
		_w7962_,
		_w7964_,
		_w7965_
	);
	LUT3 #(
		.INIT('h45)
	) name7900 (
		_w7961_,
		_w7962_,
		_w7964_,
		_w7966_
	);
	LUT3 #(
		.INIT('h82)
	) name7901 (
		_w7958_,
		_w7959_,
		_w7960_,
		_w7967_
	);
	LUT2 #(
		.INIT('h2)
	) name7902 (
		_w7963_,
		_w7967_,
		_w7968_
	);
	LUT2 #(
		.INIT('h1)
	) name7903 (
		_w7907_,
		_w7967_,
		_w7969_
	);
	LUT3 #(
		.INIT('h23)
	) name7904 (
		_w7962_,
		_w7968_,
		_w7969_,
		_w7970_
	);
	LUT3 #(
		.INIT('h69)
	) name7905 (
		_w7958_,
		_w7959_,
		_w7960_,
		_w7971_
	);
	LUT4 #(
		.INIT('hffe1)
	) name7906 (
		_w7907_,
		_w7962_,
		_w7963_,
		_w7971_,
		_w7972_
	);
	LUT3 #(
		.INIT('hd0)
	) name7907 (
		_w7966_,
		_w7970_,
		_w7972_,
		_w7973_
	);
	LUT4 #(
		.INIT('h5100)
	) name7908 (
		_w7954_,
		_w7966_,
		_w7970_,
		_w7972_,
		_w7974_
	);
	LUT4 #(
		.INIT('h08aa)
	) name7909 (
		_w7952_,
		_w7966_,
		_w7970_,
		_w7972_,
		_w7975_
	);
	LUT4 #(
		.INIT('ha208)
	) name7910 (
		_w7924_,
		_w7952_,
		_w7953_,
		_w7973_,
		_w7976_
	);
	LUT4 #(
		.INIT('h0451)
	) name7911 (
		_w7924_,
		_w7952_,
		_w7953_,
		_w7973_,
		_w7977_
	);
	LUT4 #(
		.INIT('h595a)
	) name7912 (
		_w7924_,
		_w7953_,
		_w7974_,
		_w7975_,
		_w7978_
	);
	LUT3 #(
		.INIT('h10)
	) name7913 (
		_w7915_,
		_w7923_,
		_w7978_,
		_w7979_
	);
	LUT4 #(
		.INIT('h8f00)
	) name7914 (
		_w7738_,
		_w7798_,
		_w7922_,
		_w7979_,
		_w7980_
	);
	LUT4 #(
		.INIT('hd0fd)
	) name7915 (
		_w7799_,
		_w7857_,
		_w7861_,
		_w7914_,
		_w7981_
	);
	LUT4 #(
		.INIT('h8f00)
	) name7916 (
		_w7738_,
		_w7798_,
		_w7922_,
		_w7981_,
		_w7982_
	);
	LUT3 #(
		.INIT('h32)
	) name7917 (
		_w7978_,
		_w7980_,
		_w7982_,
		_w7983_
	);
	LUT3 #(
		.INIT('h01)
	) name7918 (
		_w7915_,
		_w7923_,
		_w7977_,
		_w7984_
	);
	LUT4 #(
		.INIT('h8f00)
	) name7919 (
		_w7738_,
		_w7798_,
		_w7922_,
		_w7984_,
		_w7985_
	);
	LUT4 #(
		.INIT('h153f)
	) name7920 (
		\a[40] ,
		\a[41] ,
		\a[60] ,
		\a[61] ,
		_w7986_
	);
	LUT4 #(
		.INIT('h000d)
	) name7921 (
		_w7803_,
		_w7862_,
		_w7863_,
		_w7944_,
		_w7987_
	);
	LUT3 #(
		.INIT('h0d)
	) name7922 (
		_w7902_,
		_w7930_,
		_w7931_,
		_w7988_
	);
	LUT2 #(
		.INIT('h8)
	) name7923 (
		\a[39] ,
		\a[63] ,
		_w7989_
	);
	LUT4 #(
		.INIT('h153f)
	) name7924 (
		\a[41] ,
		\a[42] ,
		\a[60] ,
		\a[61] ,
		_w7990_
	);
	LUT2 #(
		.INIT('h8)
	) name7925 (
		\a[42] ,
		\a[61] ,
		_w7991_
	);
	LUT4 #(
		.INIT('h8000)
	) name7926 (
		\a[41] ,
		\a[42] ,
		\a[60] ,
		\a[61] ,
		_w7992_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7927 (
		\a[41] ,
		\a[42] ,
		\a[60] ,
		\a[61] ,
		_w7993_
	);
	LUT2 #(
		.INIT('h6)
	) name7928 (
		_w7989_,
		_w7993_,
		_w7994_
	);
	LUT4 #(
		.INIT('he11e)
	) name7929 (
		_w7986_,
		_w7987_,
		_w7988_,
		_w7994_,
		_w7995_
	);
	LUT4 #(
		.INIT('h004f)
	) name7930 (
		_w7942_,
		_w7947_,
		_w7948_,
		_w7995_,
		_w7996_
	);
	LUT4 #(
		.INIT('hb000)
	) name7931 (
		_w7942_,
		_w7947_,
		_w7948_,
		_w7995_,
		_w7997_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name7932 (
		_w7942_,
		_w7947_,
		_w7948_,
		_w7995_,
		_w7998_
	);
	LUT4 #(
		.INIT('h153f)
	) name7933 (
		\a[43] ,
		\a[44] ,
		\a[58] ,
		\a[59] ,
		_w7999_
	);
	LUT4 #(
		.INIT('h8000)
	) name7934 (
		\a[43] ,
		\a[44] ,
		\a[58] ,
		\a[59] ,
		_w8000_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7935 (
		\a[43] ,
		\a[44] ,
		\a[58] ,
		\a[59] ,
		_w8001_
	);
	LUT2 #(
		.INIT('h8)
	) name7936 (
		\a[45] ,
		\a[57] ,
		_w8002_
	);
	LUT4 #(
		.INIT('h153f)
	) name7937 (
		\a[46] ,
		\a[47] ,
		\a[55] ,
		\a[56] ,
		_w8003_
	);
	LUT4 #(
		.INIT('h8000)
	) name7938 (
		\a[46] ,
		\a[47] ,
		\a[55] ,
		\a[56] ,
		_w8004_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7939 (
		\a[46] ,
		\a[47] ,
		\a[55] ,
		\a[56] ,
		_w8005_
	);
	LUT4 #(
		.INIT('h0660)
	) name7940 (
		_w6209_,
		_w8001_,
		_w8002_,
		_w8005_,
		_w8006_
	);
	LUT4 #(
		.INIT('h9009)
	) name7941 (
		_w6209_,
		_w8001_,
		_w8002_,
		_w8005_,
		_w8007_
	);
	LUT4 #(
		.INIT('h6996)
	) name7942 (
		_w6209_,
		_w8001_,
		_w8002_,
		_w8005_,
		_w8008_
	);
	LUT2 #(
		.INIT('h8)
	) name7943 (
		\a[48] ,
		\a[54] ,
		_w8009_
	);
	LUT4 #(
		.INIT('h153f)
	) name7944 (
		\a[49] ,
		\a[50] ,
		\a[52] ,
		\a[53] ,
		_w8010_
	);
	LUT4 #(
		.INIT('h8000)
	) name7945 (
		\a[49] ,
		\a[50] ,
		\a[52] ,
		\a[53] ,
		_w8011_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7946 (
		\a[49] ,
		\a[50] ,
		\a[52] ,
		\a[53] ,
		_w8012_
	);
	LUT2 #(
		.INIT('h6)
	) name7947 (
		_w8009_,
		_w8012_,
		_w8013_
	);
	LUT2 #(
		.INIT('h6)
	) name7948 (
		_w8008_,
		_w8013_,
		_w8014_
	);
	LUT2 #(
		.INIT('h6)
	) name7949 (
		_w7998_,
		_w8014_,
		_w8015_
	);
	LUT4 #(
		.INIT('hae00)
	) name7950 (
		_w7965_,
		_w7966_,
		_w7970_,
		_w8015_,
		_w8016_
	);
	LUT3 #(
		.INIT('h17)
	) name7951 (
		_w7925_,
		_w7941_,
		_w7950_,
		_w8017_
	);
	LUT3 #(
		.INIT('hd4)
	) name7952 (
		_w7958_,
		_w7959_,
		_w7960_,
		_w8018_
	);
	LUT4 #(
		.INIT('he800)
	) name7953 (
		_w7925_,
		_w7941_,
		_w7950_,
		_w8018_,
		_w8019_
	);
	LUT4 #(
		.INIT('he0c0)
	) name7954 (
		\a[39] ,
		\a[50] ,
		\a[51] ,
		\a[62] ,
		_w8020_
	);
	LUT4 #(
		.INIT('h000d)
	) name7955 (
		_w7936_,
		_w7937_,
		_w7938_,
		_w8020_,
		_w8021_
	);
	LUT4 #(
		.INIT('hf200)
	) name7956 (
		_w7936_,
		_w7937_,
		_w7938_,
		_w8020_,
		_w8022_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7957 (
		_w7936_,
		_w7937_,
		_w7938_,
		_w8020_,
		_w8023_
	);
	LUT3 #(
		.INIT('h0d)
	) name7958 (
		_w7926_,
		_w7927_,
		_w7928_,
		_w8024_
	);
	LUT2 #(
		.INIT('h6)
	) name7959 (
		_w8023_,
		_w8024_,
		_w8025_
	);
	LUT3 #(
		.INIT('h17)
	) name7960 (
		_w7955_,
		_w7956_,
		_w7957_,
		_w8026_
	);
	LUT3 #(
		.INIT('h32)
	) name7961 (
		_w7933_,
		_w7934_,
		_w7940_,
		_w8027_
	);
	LUT3 #(
		.INIT('h69)
	) name7962 (
		_w8025_,
		_w8026_,
		_w8027_,
		_w8028_
	);
	LUT4 #(
		.INIT('h0017)
	) name7963 (
		_w7925_,
		_w7941_,
		_w7950_,
		_w8018_,
		_w8029_
	);
	LUT4 #(
		.INIT('hf949)
	) name7964 (
		_w8017_,
		_w8018_,
		_w8028_,
		_w8029_,
		_w8030_
	);
	LUT3 #(
		.INIT('h0b)
	) name7965 (
		_w7962_,
		_w7964_,
		_w8015_,
		_w8031_
	);
	LUT3 #(
		.INIT('hd0)
	) name7966 (
		_w7966_,
		_w7970_,
		_w8031_,
		_w8032_
	);
	LUT4 #(
		.INIT('h20f0)
	) name7967 (
		_w7966_,
		_w7970_,
		_w8030_,
		_w8031_,
		_w8033_
	);
	LUT2 #(
		.INIT('h4)
	) name7968 (
		_w8016_,
		_w8033_,
		_w8034_
	);
	LUT4 #(
		.INIT('h32cd)
	) name7969 (
		_w7961_,
		_w7965_,
		_w7970_,
		_w8015_,
		_w8035_
	);
	LUT2 #(
		.INIT('h1)
	) name7970 (
		_w8030_,
		_w8035_,
		_w8036_
	);
	LUT3 #(
		.INIT('hc9)
	) name7971 (
		_w8016_,
		_w8030_,
		_w8032_,
		_w8037_
	);
	LUT2 #(
		.INIT('h1)
	) name7972 (
		_w7953_,
		_w7975_,
		_w8038_
	);
	LUT2 #(
		.INIT('h1)
	) name7973 (
		_w8037_,
		_w8038_,
		_w8039_
	);
	LUT4 #(
		.INIT('h1011)
	) name7974 (
		_w7953_,
		_w7975_,
		_w8016_,
		_w8033_,
		_w8040_
	);
	LUT3 #(
		.INIT('he1)
	) name7975 (
		_w8034_,
		_w8036_,
		_w8038_,
		_w8041_
	);
	LUT3 #(
		.INIT('h1e)
	) name7976 (
		_w7976_,
		_w7985_,
		_w8041_,
		_w8042_
	);
	LUT3 #(
		.INIT('h45)
	) name7977 (
		_w7976_,
		_w8036_,
		_w8040_,
		_w8043_
	);
	LUT3 #(
		.INIT('h45)
	) name7978 (
		_w8021_,
		_w8022_,
		_w8024_,
		_w8044_
	);
	LUT4 #(
		.INIT('h1f01)
	) name7979 (
		_w7986_,
		_w7987_,
		_w7988_,
		_w7994_,
		_w8045_
	);
	LUT3 #(
		.INIT('h32)
	) name7980 (
		_w8006_,
		_w8007_,
		_w8013_,
		_w8046_
	);
	LUT3 #(
		.INIT('h96)
	) name7981 (
		_w8044_,
		_w8045_,
		_w8046_,
		_w8047_
	);
	LUT3 #(
		.INIT('h54)
	) name7982 (
		_w7996_,
		_w7997_,
		_w8014_,
		_w8048_
	);
	LUT3 #(
		.INIT('hd4)
	) name7983 (
		_w8025_,
		_w8026_,
		_w8027_,
		_w8049_
	);
	LUT4 #(
		.INIT('hab54)
	) name7984 (
		_w7996_,
		_w7997_,
		_w8014_,
		_w8049_,
		_w8050_
	);
	LUT2 #(
		.INIT('h6)
	) name7985 (
		_w8047_,
		_w8050_,
		_w8051_
	);
	LUT2 #(
		.INIT('h8)
	) name7986 (
		\a[40] ,
		\a[63] ,
		_w8052_
	);
	LUT4 #(
		.INIT('h0dff)
	) name7987 (
		_w8009_,
		_w8010_,
		_w8011_,
		_w8052_,
		_w8053_
	);
	LUT4 #(
		.INIT('h000d)
	) name7988 (
		_w8009_,
		_w8010_,
		_w8011_,
		_w8052_,
		_w8054_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7989 (
		_w8009_,
		_w8010_,
		_w8011_,
		_w8052_,
		_w8055_
	);
	LUT3 #(
		.INIT('h0d)
	) name7990 (
		_w8002_,
		_w8003_,
		_w8004_,
		_w8056_
	);
	LUT2 #(
		.INIT('h6)
	) name7991 (
		_w8055_,
		_w8056_,
		_w8057_
	);
	LUT3 #(
		.INIT('h0d)
	) name7992 (
		_w7989_,
		_w7990_,
		_w7992_,
		_w8058_
	);
	LUT3 #(
		.INIT('h0d)
	) name7993 (
		_w6209_,
		_w7999_,
		_w8000_,
		_w8059_
	);
	LUT4 #(
		.INIT('h153f)
	) name7994 (
		\a[44] ,
		\a[45] ,
		\a[58] ,
		\a[59] ,
		_w8060_
	);
	LUT4 #(
		.INIT('h8000)
	) name7995 (
		\a[44] ,
		\a[45] ,
		\a[58] ,
		\a[59] ,
		_w8061_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7996 (
		\a[44] ,
		\a[45] ,
		\a[58] ,
		\a[59] ,
		_w8062_
	);
	LUT2 #(
		.INIT('h6)
	) name7997 (
		_w7991_,
		_w8062_,
		_w8063_
	);
	LUT3 #(
		.INIT('h69)
	) name7998 (
		_w8058_,
		_w8059_,
		_w8063_,
		_w8064_
	);
	LUT2 #(
		.INIT('h8)
	) name7999 (
		\a[43] ,
		\a[60] ,
		_w8065_
	);
	LUT4 #(
		.INIT('h153f)
	) name8000 (
		\a[46] ,
		\a[47] ,
		\a[56] ,
		\a[57] ,
		_w8066_
	);
	LUT4 #(
		.INIT('h8000)
	) name8001 (
		\a[46] ,
		\a[47] ,
		\a[56] ,
		\a[57] ,
		_w8067_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8002 (
		\a[46] ,
		\a[47] ,
		\a[56] ,
		\a[57] ,
		_w8068_
	);
	LUT2 #(
		.INIT('h8)
	) name8003 (
		\a[48] ,
		\a[55] ,
		_w8069_
	);
	LUT4 #(
		.INIT('h153f)
	) name8004 (
		\a[49] ,
		\a[50] ,
		\a[53] ,
		\a[54] ,
		_w8070_
	);
	LUT4 #(
		.INIT('h8000)
	) name8005 (
		\a[49] ,
		\a[50] ,
		\a[53] ,
		\a[54] ,
		_w8071_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8006 (
		\a[49] ,
		\a[50] ,
		\a[53] ,
		\a[54] ,
		_w8072_
	);
	LUT4 #(
		.INIT('h0660)
	) name8007 (
		_w8065_,
		_w8068_,
		_w8069_,
		_w8072_,
		_w8073_
	);
	LUT4 #(
		.INIT('h9009)
	) name8008 (
		_w8065_,
		_w8068_,
		_w8069_,
		_w8072_,
		_w8074_
	);
	LUT4 #(
		.INIT('h6996)
	) name8009 (
		_w8065_,
		_w8068_,
		_w8069_,
		_w8072_,
		_w8075_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8010 (
		\a[41] ,
		\a[51] ,
		\a[52] ,
		\a[62] ,
		_w8076_
	);
	LUT2 #(
		.INIT('h6)
	) name8011 (
		_w8075_,
		_w8076_,
		_w8077_
	);
	LUT3 #(
		.INIT('h96)
	) name8012 (
		_w8057_,
		_w8064_,
		_w8077_,
		_w8078_
	);
	LUT4 #(
		.INIT('hae00)
	) name8013 (
		_w8019_,
		_w8028_,
		_w8029_,
		_w8078_,
		_w8079_
	);
	LUT4 #(
		.INIT('h0051)
	) name8014 (
		_w8019_,
		_w8028_,
		_w8029_,
		_w8078_,
		_w8080_
	);
	LUT4 #(
		.INIT('h51ae)
	) name8015 (
		_w8019_,
		_w8028_,
		_w8029_,
		_w8078_,
		_w8081_
	);
	LUT2 #(
		.INIT('h1)
	) name8016 (
		_w8051_,
		_w8081_,
		_w8082_
	);
	LUT3 #(
		.INIT('h02)
	) name8017 (
		_w8051_,
		_w8079_,
		_w8080_,
		_w8083_
	);
	LUT4 #(
		.INIT('h000e)
	) name8018 (
		_w8016_,
		_w8033_,
		_w8082_,
		_w8083_,
		_w8084_
	);
	LUT3 #(
		.INIT('ha9)
	) name8019 (
		_w8051_,
		_w8079_,
		_w8080_,
		_w8085_
	);
	LUT3 #(
		.INIT('h01)
	) name8020 (
		_w8016_,
		_w8033_,
		_w8085_,
		_w8086_
	);
	LUT4 #(
		.INIT('heee1)
	) name8021 (
		_w8016_,
		_w8033_,
		_w8082_,
		_w8083_,
		_w8087_
	);
	LUT4 #(
		.INIT('hdc23)
	) name8022 (
		_w7985_,
		_w8039_,
		_w8043_,
		_w8087_,
		_w8088_
	);
	LUT4 #(
		.INIT('h000e)
	) name8023 (
		_w8034_,
		_w8036_,
		_w8038_,
		_w8084_,
		_w8089_
	);
	LUT4 #(
		.INIT('h0045)
	) name8024 (
		_w7976_,
		_w8036_,
		_w8040_,
		_w8084_,
		_w8090_
	);
	LUT3 #(
		.INIT('h31)
	) name8025 (
		_w8051_,
		_w8079_,
		_w8080_,
		_w8091_
	);
	LUT3 #(
		.INIT('h0d)
	) name8026 (
		_w8069_,
		_w8070_,
		_w8071_,
		_w8092_
	);
	LUT3 #(
		.INIT('h0d)
	) name8027 (
		_w8065_,
		_w8066_,
		_w8067_,
		_w8093_
	);
	LUT3 #(
		.INIT('h0d)
	) name8028 (
		_w7991_,
		_w8060_,
		_w8061_,
		_w8094_
	);
	LUT3 #(
		.INIT('h96)
	) name8029 (
		_w8092_,
		_w8093_,
		_w8094_,
		_w8095_
	);
	LUT3 #(
		.INIT('h32)
	) name8030 (
		_w8073_,
		_w8074_,
		_w8076_,
		_w8096_
	);
	LUT2 #(
		.INIT('h8)
	) name8031 (
		\a[44] ,
		\a[60] ,
		_w8097_
	);
	LUT4 #(
		.INIT('h153f)
	) name8032 (
		\a[43] ,
		\a[45] ,
		\a[59] ,
		\a[61] ,
		_w8098_
	);
	LUT4 #(
		.INIT('h8000)
	) name8033 (
		\a[43] ,
		\a[45] ,
		\a[59] ,
		\a[61] ,
		_w8099_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8034 (
		\a[43] ,
		\a[45] ,
		\a[59] ,
		\a[61] ,
		_w8100_
	);
	LUT2 #(
		.INIT('h8)
	) name8035 (
		\a[46] ,
		\a[58] ,
		_w8101_
	);
	LUT4 #(
		.INIT('h153f)
	) name8036 (
		\a[47] ,
		\a[48] ,
		\a[56] ,
		\a[57] ,
		_w8102_
	);
	LUT4 #(
		.INIT('h8000)
	) name8037 (
		\a[47] ,
		\a[48] ,
		\a[56] ,
		\a[57] ,
		_w8103_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8038 (
		\a[47] ,
		\a[48] ,
		\a[56] ,
		\a[57] ,
		_w8104_
	);
	LUT4 #(
		.INIT('h0660)
	) name8039 (
		_w8097_,
		_w8100_,
		_w8101_,
		_w8104_,
		_w8105_
	);
	LUT4 #(
		.INIT('h9009)
	) name8040 (
		_w8097_,
		_w8100_,
		_w8101_,
		_w8104_,
		_w8106_
	);
	LUT4 #(
		.INIT('h6996)
	) name8041 (
		_w8097_,
		_w8100_,
		_w8101_,
		_w8104_,
		_w8107_
	);
	LUT2 #(
		.INIT('h8)
	) name8042 (
		\a[49] ,
		\a[55] ,
		_w8108_
	);
	LUT4 #(
		.INIT('h153f)
	) name8043 (
		\a[50] ,
		\a[51] ,
		\a[53] ,
		\a[54] ,
		_w8109_
	);
	LUT4 #(
		.INIT('h8000)
	) name8044 (
		\a[50] ,
		\a[51] ,
		\a[53] ,
		\a[54] ,
		_w8110_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8045 (
		\a[50] ,
		\a[51] ,
		\a[53] ,
		\a[54] ,
		_w8111_
	);
	LUT2 #(
		.INIT('h6)
	) name8046 (
		_w8108_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h6)
	) name8047 (
		_w8107_,
		_w8112_,
		_w8113_
	);
	LUT3 #(
		.INIT('h69)
	) name8048 (
		_w8095_,
		_w8096_,
		_w8113_,
		_w8114_
	);
	LUT4 #(
		.INIT('h0017)
	) name8049 (
		_w8047_,
		_w8048_,
		_w8049_,
		_w8114_,
		_w8115_
	);
	LUT3 #(
		.INIT('he8)
	) name8050 (
		_w8044_,
		_w8045_,
		_w8046_,
		_w8116_
	);
	LUT3 #(
		.INIT('h71)
	) name8051 (
		_w8057_,
		_w8064_,
		_w8077_,
		_w8117_
	);
	LUT2 #(
		.INIT('h1)
	) name8052 (
		_w8116_,
		_w8117_,
		_w8118_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8053 (
		\a[41] ,
		\a[51] ,
		\a[52] ,
		\a[62] ,
		_w8119_
	);
	LUT4 #(
		.INIT('h153f)
	) name8054 (
		\a[41] ,
		\a[42] ,
		\a[62] ,
		\a[63] ,
		_w8120_
	);
	LUT2 #(
		.INIT('h8)
	) name8055 (
		\a[42] ,
		\a[63] ,
		_w8121_
	);
	LUT4 #(
		.INIT('h8000)
	) name8056 (
		\a[41] ,
		\a[42] ,
		\a[62] ,
		\a[63] ,
		_w8122_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8057 (
		\a[41] ,
		\a[42] ,
		\a[62] ,
		\a[63] ,
		_w8123_
	);
	LUT2 #(
		.INIT('h6)
	) name8058 (
		_w8119_,
		_w8123_,
		_w8124_
	);
	LUT4 #(
		.INIT('h00a8)
	) name8059 (
		_w8053_,
		_w8054_,
		_w8056_,
		_w8124_,
		_w8125_
	);
	LUT4 #(
		.INIT('h5700)
	) name8060 (
		_w8053_,
		_w8054_,
		_w8056_,
		_w8124_,
		_w8126_
	);
	LUT4 #(
		.INIT('hf807)
	) name8061 (
		_w8053_,
		_w8056_,
		_w8054_,
		_w8124_,
		_w8127_
	);
	LUT3 #(
		.INIT('h8e)
	) name8062 (
		_w8058_,
		_w8059_,
		_w8063_,
		_w8128_
	);
	LUT2 #(
		.INIT('h6)
	) name8063 (
		_w8127_,
		_w8128_,
		_w8129_
	);
	LUT3 #(
		.INIT('h69)
	) name8064 (
		_w8116_,
		_w8117_,
		_w8129_,
		_w8130_
	);
	LUT4 #(
		.INIT('he800)
	) name8065 (
		_w8047_,
		_w8048_,
		_w8049_,
		_w8114_,
		_w8131_
	);
	LUT3 #(
		.INIT('hc9)
	) name8066 (
		_w8115_,
		_w8130_,
		_w8131_,
		_w8132_
	);
	LUT2 #(
		.INIT('h4)
	) name8067 (
		_w8091_,
		_w8132_,
		_w8133_
	);
	LUT2 #(
		.INIT('h2)
	) name8068 (
		_w8091_,
		_w8132_,
		_w8134_
	);
	LUT2 #(
		.INIT('h9)
	) name8069 (
		_w8091_,
		_w8132_,
		_w8135_
	);
	LUT2 #(
		.INIT('h4)
	) name8070 (
		_w8086_,
		_w8135_,
		_w8136_
	);
	LUT4 #(
		.INIT('h2300)
	) name8071 (
		_w7985_,
		_w8089_,
		_w8090_,
		_w8136_,
		_w8137_
	);
	LUT4 #(
		.INIT('h0203)
	) name8072 (
		_w7985_,
		_w8086_,
		_w8089_,
		_w8090_,
		_w8138_
	);
	LUT3 #(
		.INIT('h32)
	) name8073 (
		_w8135_,
		_w8137_,
		_w8138_,
		_w8139_
	);
	LUT2 #(
		.INIT('h1)
	) name8074 (
		_w8086_,
		_w8134_,
		_w8140_
	);
	LUT4 #(
		.INIT('h2300)
	) name8075 (
		_w7985_,
		_w8089_,
		_w8090_,
		_w8140_,
		_w8141_
	);
	LUT3 #(
		.INIT('h70)
	) name8076 (
		_w8116_,
		_w8117_,
		_w8129_,
		_w8142_
	);
	LUT3 #(
		.INIT('h8e)
	) name8077 (
		_w8116_,
		_w8117_,
		_w8129_,
		_w8143_
	);
	LUT3 #(
		.INIT('hd4)
	) name8078 (
		_w8095_,
		_w8096_,
		_w8113_,
		_w8144_
	);
	LUT2 #(
		.INIT('h8)
	) name8079 (
		\a[49] ,
		\a[56] ,
		_w8145_
	);
	LUT4 #(
		.INIT('h153f)
	) name8080 (
		\a[50] ,
		\a[51] ,
		\a[54] ,
		\a[55] ,
		_w8146_
	);
	LUT4 #(
		.INIT('h8000)
	) name8081 (
		\a[50] ,
		\a[51] ,
		\a[54] ,
		\a[55] ,
		_w8147_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8082 (
		\a[50] ,
		\a[51] ,
		\a[54] ,
		\a[55] ,
		_w8148_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8083 (
		\a[43] ,
		\a[52] ,
		\a[53] ,
		\a[62] ,
		_w8149_
	);
	LUT3 #(
		.INIT('h60)
	) name8084 (
		_w8145_,
		_w8148_,
		_w8149_,
		_w8150_
	);
	LUT3 #(
		.INIT('h96)
	) name8085 (
		_w8145_,
		_w8148_,
		_w8149_,
		_w8151_
	);
	LUT4 #(
		.INIT('h1700)
	) name8086 (
		_w8092_,
		_w8093_,
		_w8094_,
		_w8151_,
		_w8152_
	);
	LUT4 #(
		.INIT('he817)
	) name8087 (
		_w8092_,
		_w8093_,
		_w8094_,
		_w8151_,
		_w8153_
	);
	LUT3 #(
		.INIT('h0d)
	) name8088 (
		_w8119_,
		_w8120_,
		_w8122_,
		_w8154_
	);
	LUT4 #(
		.INIT('h153f)
	) name8089 (
		\a[44] ,
		\a[45] ,
		\a[60] ,
		\a[61] ,
		_w8155_
	);
	LUT4 #(
		.INIT('h8000)
	) name8090 (
		\a[44] ,
		\a[45] ,
		\a[60] ,
		\a[61] ,
		_w8156_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8091 (
		\a[44] ,
		\a[45] ,
		\a[60] ,
		\a[61] ,
		_w8157_
	);
	LUT2 #(
		.INIT('h6)
	) name8092 (
		_w8121_,
		_w8157_,
		_w8158_
	);
	LUT2 #(
		.INIT('h8)
	) name8093 (
		\a[46] ,
		\a[59] ,
		_w8159_
	);
	LUT4 #(
		.INIT('h153f)
	) name8094 (
		\a[47] ,
		\a[48] ,
		\a[57] ,
		\a[58] ,
		_w8160_
	);
	LUT4 #(
		.INIT('h8000)
	) name8095 (
		\a[47] ,
		\a[48] ,
		\a[57] ,
		\a[58] ,
		_w8161_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8096 (
		\a[47] ,
		\a[48] ,
		\a[57] ,
		\a[58] ,
		_w8162_
	);
	LUT2 #(
		.INIT('h6)
	) name8097 (
		_w8159_,
		_w8162_,
		_w8163_
	);
	LUT3 #(
		.INIT('h69)
	) name8098 (
		_w8154_,
		_w8158_,
		_w8163_,
		_w8164_
	);
	LUT2 #(
		.INIT('h1)
	) name8099 (
		_w8153_,
		_w8164_,
		_w8165_
	);
	LUT2 #(
		.INIT('h8)
	) name8100 (
		_w8153_,
		_w8164_,
		_w8166_
	);
	LUT2 #(
		.INIT('h6)
	) name8101 (
		_w8153_,
		_w8164_,
		_w8167_
	);
	LUT2 #(
		.INIT('h8)
	) name8102 (
		_w8144_,
		_w8167_,
		_w8168_
	);
	LUT2 #(
		.INIT('h6)
	) name8103 (
		_w8144_,
		_w8167_,
		_w8169_
	);
	LUT3 #(
		.INIT('h0d)
	) name8104 (
		_w8101_,
		_w8102_,
		_w8103_,
		_w8170_
	);
	LUT3 #(
		.INIT('h0d)
	) name8105 (
		_w8108_,
		_w8109_,
		_w8110_,
		_w8171_
	);
	LUT3 #(
		.INIT('h0d)
	) name8106 (
		_w8097_,
		_w8098_,
		_w8099_,
		_w8172_
	);
	LUT3 #(
		.INIT('h96)
	) name8107 (
		_w8170_,
		_w8171_,
		_w8172_,
		_w8173_
	);
	LUT3 #(
		.INIT('h32)
	) name8108 (
		_w8105_,
		_w8106_,
		_w8112_,
		_w8174_
	);
	LUT2 #(
		.INIT('h2)
	) name8109 (
		_w8173_,
		_w8174_,
		_w8175_
	);
	LUT2 #(
		.INIT('h4)
	) name8110 (
		_w8173_,
		_w8174_,
		_w8176_
	);
	LUT2 #(
		.INIT('h9)
	) name8111 (
		_w8173_,
		_w8174_,
		_w8177_
	);
	LUT3 #(
		.INIT('h45)
	) name8112 (
		_w8125_,
		_w8126_,
		_w8128_,
		_w8178_
	);
	LUT2 #(
		.INIT('h6)
	) name8113 (
		_w8177_,
		_w8178_,
		_w8179_
	);
	LUT3 #(
		.INIT('hed)
	) name8114 (
		_w8143_,
		_w8169_,
		_w8179_,
		_w8180_
	);
	LUT4 #(
		.INIT('h10e0)
	) name8115 (
		_w8118_,
		_w8142_,
		_w8169_,
		_w8179_,
		_w8181_
	);
	LUT2 #(
		.INIT('h2)
	) name8116 (
		_w8180_,
		_w8181_,
		_w8182_
	);
	LUT3 #(
		.INIT('h54)
	) name8117 (
		_w8115_,
		_w8130_,
		_w8131_,
		_w8183_
	);
	LUT2 #(
		.INIT('h9)
	) name8118 (
		_w8182_,
		_w8183_,
		_w8184_
	);
	LUT3 #(
		.INIT('h1e)
	) name8119 (
		_w8133_,
		_w8141_,
		_w8184_,
		_w8185_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8120 (
		_w8091_,
		_w8132_,
		_w8182_,
		_w8183_,
		_w8186_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name8121 (
		_w8116_,
		_w8117_,
		_w8177_,
		_w8178_,
		_w8187_
	);
	LUT2 #(
		.INIT('h4)
	) name8122 (
		_w8142_,
		_w8187_,
		_w8188_
	);
	LUT3 #(
		.INIT('h23)
	) name8123 (
		_w8142_,
		_w8168_,
		_w8187_,
		_w8189_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name8124 (
		_w8144_,
		_w8167_,
		_w8177_,
		_w8178_,
		_w8190_
	);
	LUT4 #(
		.INIT('heee0)
	) name8125 (
		_w8116_,
		_w8117_,
		_w8144_,
		_w8167_,
		_w8191_
	);
	LUT3 #(
		.INIT('h23)
	) name8126 (
		_w8142_,
		_w8190_,
		_w8191_,
		_w8192_
	);
	LUT3 #(
		.INIT('h13)
	) name8127 (
		\a[43] ,
		\a[52] ,
		\a[62] ,
		_w8193_
	);
	LUT2 #(
		.INIT('h8)
	) name8128 (
		\a[43] ,
		\a[63] ,
		_w8194_
	);
	LUT3 #(
		.INIT('h80)
	) name8129 (
		\a[43] ,
		\a[53] ,
		\a[63] ,
		_w8195_
	);
	LUT2 #(
		.INIT('h4)
	) name8130 (
		_w8193_,
		_w8195_,
		_w8196_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8131 (
		\a[43] ,
		\a[52] ,
		\a[53] ,
		\a[62] ,
		_w8197_
	);
	LUT2 #(
		.INIT('h1)
	) name8132 (
		_w8194_,
		_w8197_,
		_w8198_
	);
	LUT3 #(
		.INIT('hd2)
	) name8133 (
		\a[53] ,
		_w8193_,
		_w8194_,
		_w8199_
	);
	LUT3 #(
		.INIT('h0d)
	) name8134 (
		_w8145_,
		_w8146_,
		_w8147_,
		_w8200_
	);
	LUT2 #(
		.INIT('h6)
	) name8135 (
		_w8199_,
		_w8200_,
		_w8201_
	);
	LUT3 #(
		.INIT('hd4)
	) name8136 (
		_w8154_,
		_w8158_,
		_w8163_,
		_w8202_
	);
	LUT4 #(
		.INIT('he11e)
	) name8137 (
		_w8150_,
		_w8152_,
		_w8201_,
		_w8202_,
		_w8203_
	);
	LUT4 #(
		.INIT('h00e8)
	) name8138 (
		_w8144_,
		_w8153_,
		_w8164_,
		_w8203_,
		_w8204_
	);
	LUT4 #(
		.INIT('h1700)
	) name8139 (
		_w8144_,
		_w8153_,
		_w8164_,
		_w8203_,
		_w8205_
	);
	LUT4 #(
		.INIT('hf20d)
	) name8140 (
		_w8144_,
		_w8165_,
		_w8166_,
		_w8203_,
		_w8206_
	);
	LUT2 #(
		.INIT('h8)
	) name8141 (
		\a[47] ,
		\a[59] ,
		_w8207_
	);
	LUT4 #(
		.INIT('h153f)
	) name8142 (
		\a[48] ,
		\a[49] ,
		\a[57] ,
		\a[58] ,
		_w8208_
	);
	LUT4 #(
		.INIT('h8000)
	) name8143 (
		\a[48] ,
		\a[49] ,
		\a[57] ,
		\a[58] ,
		_w8209_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8144 (
		\a[48] ,
		\a[49] ,
		\a[57] ,
		\a[58] ,
		_w8210_
	);
	LUT2 #(
		.INIT('h8)
	) name8145 (
		\a[50] ,
		\a[56] ,
		_w8211_
	);
	LUT4 #(
		.INIT('h153f)
	) name8146 (
		\a[51] ,
		\a[52] ,
		\a[54] ,
		\a[55] ,
		_w8212_
	);
	LUT4 #(
		.INIT('h8000)
	) name8147 (
		\a[51] ,
		\a[52] ,
		\a[54] ,
		\a[55] ,
		_w8213_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8148 (
		\a[51] ,
		\a[52] ,
		\a[54] ,
		\a[55] ,
		_w8214_
	);
	LUT4 #(
		.INIT('h0660)
	) name8149 (
		_w8207_,
		_w8210_,
		_w8211_,
		_w8214_,
		_w8215_
	);
	LUT4 #(
		.INIT('h6996)
	) name8150 (
		_w8207_,
		_w8210_,
		_w8211_,
		_w8214_,
		_w8216_
	);
	LUT4 #(
		.INIT('h1700)
	) name8151 (
		_w8170_,
		_w8171_,
		_w8172_,
		_w8216_,
		_w8217_
	);
	LUT4 #(
		.INIT('he817)
	) name8152 (
		_w8170_,
		_w8171_,
		_w8172_,
		_w8216_,
		_w8218_
	);
	LUT3 #(
		.INIT('h0d)
	) name8153 (
		_w8121_,
		_w8155_,
		_w8156_,
		_w8219_
	);
	LUT3 #(
		.INIT('h0d)
	) name8154 (
		_w8159_,
		_w8160_,
		_w8161_,
		_w8220_
	);
	LUT2 #(
		.INIT('h8)
	) name8155 (
		\a[44] ,
		\a[62] ,
		_w8221_
	);
	LUT4 #(
		.INIT('h153f)
	) name8156 (
		\a[45] ,
		\a[46] ,
		\a[60] ,
		\a[61] ,
		_w8222_
	);
	LUT4 #(
		.INIT('h8000)
	) name8157 (
		\a[45] ,
		\a[46] ,
		\a[60] ,
		\a[61] ,
		_w8223_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8158 (
		\a[45] ,
		\a[46] ,
		\a[60] ,
		\a[61] ,
		_w8224_
	);
	LUT2 #(
		.INIT('h6)
	) name8159 (
		_w8221_,
		_w8224_,
		_w8225_
	);
	LUT3 #(
		.INIT('h69)
	) name8160 (
		_w8219_,
		_w8220_,
		_w8225_,
		_w8226_
	);
	LUT2 #(
		.INIT('h2)
	) name8161 (
		_w8218_,
		_w8226_,
		_w8227_
	);
	LUT2 #(
		.INIT('h9)
	) name8162 (
		_w8218_,
		_w8226_,
		_w8228_
	);
	LUT4 #(
		.INIT('hd400)
	) name8163 (
		_w8173_,
		_w8174_,
		_w8178_,
		_w8228_,
		_w8229_
	);
	LUT4 #(
		.INIT('hab54)
	) name8164 (
		_w8175_,
		_w8176_,
		_w8178_,
		_w8228_,
		_w8230_
	);
	LUT2 #(
		.INIT('h6)
	) name8165 (
		_w8206_,
		_w8230_,
		_w8231_
	);
	LUT4 #(
		.INIT('hae00)
	) name8166 (
		_w8188_,
		_w8189_,
		_w8192_,
		_w8231_,
		_w8232_
	);
	LUT4 #(
		.INIT('h0051)
	) name8167 (
		_w8188_,
		_w8189_,
		_w8192_,
		_w8231_,
		_w8233_
	);
	LUT4 #(
		.INIT('h32cd)
	) name8168 (
		_w8168_,
		_w8188_,
		_w8192_,
		_w8231_,
		_w8234_
	);
	LUT3 #(
		.INIT('h2d)
	) name8169 (
		_w8182_,
		_w8183_,
		_w8234_,
		_w8235_
	);
	LUT3 #(
		.INIT('hf0)
	) name8170 (
		_w8182_,
		_w8183_,
		_w8234_,
		_w8236_
	);
	LUT4 #(
		.INIT('hf4b0)
	) name8171 (
		_w8141_,
		_w8186_,
		_w8235_,
		_w8236_,
		_w8237_
	);
	LUT3 #(
		.INIT('h32)
	) name8172 (
		_w8204_,
		_w8205_,
		_w8230_,
		_w8238_
	);
	LUT3 #(
		.INIT('h23)
	) name8173 (
		_w8196_,
		_w8198_,
		_w8200_,
		_w8239_
	);
	LUT3 #(
		.INIT('h8e)
	) name8174 (
		_w8219_,
		_w8220_,
		_w8225_,
		_w8240_
	);
	LUT4 #(
		.INIT('he00e)
	) name8175 (
		_w8215_,
		_w8217_,
		_w8239_,
		_w8240_,
		_w8241_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name8176 (
		_w8215_,
		_w8217_,
		_w8239_,
		_w8240_,
		_w8242_
	);
	LUT4 #(
		.INIT('hef0e)
	) name8177 (
		_w8150_,
		_w8152_,
		_w8201_,
		_w8202_,
		_w8243_
	);
	LUT4 #(
		.INIT('h8000)
	) name8178 (
		\a[46] ,
		\a[47] ,
		\a[60] ,
		\a[61] ,
		_w8244_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8179 (
		\a[46] ,
		\a[47] ,
		\a[60] ,
		\a[61] ,
		_w8245_
	);
	LUT4 #(
		.INIT('hf20d)
	) name8180 (
		_w8211_,
		_w8212_,
		_w8213_,
		_w8245_,
		_w8246_
	);
	LUT2 #(
		.INIT('h8)
	) name8181 (
		\a[50] ,
		\a[57] ,
		_w8247_
	);
	LUT4 #(
		.INIT('h153f)
	) name8182 (
		\a[51] ,
		\a[52] ,
		\a[55] ,
		\a[56] ,
		_w8248_
	);
	LUT4 #(
		.INIT('h8000)
	) name8183 (
		\a[51] ,
		\a[52] ,
		\a[55] ,
		\a[56] ,
		_w8249_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8184 (
		\a[51] ,
		\a[52] ,
		\a[55] ,
		\a[56] ,
		_w8250_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8185 (
		\a[45] ,
		\a[53] ,
		\a[54] ,
		\a[62] ,
		_w8251_
	);
	LUT3 #(
		.INIT('h60)
	) name8186 (
		_w8247_,
		_w8250_,
		_w8251_,
		_w8252_
	);
	LUT3 #(
		.INIT('h09)
	) name8187 (
		_w8247_,
		_w8250_,
		_w8251_,
		_w8253_
	);
	LUT3 #(
		.INIT('h96)
	) name8188 (
		_w8247_,
		_w8250_,
		_w8251_,
		_w8254_
	);
	LUT2 #(
		.INIT('h9)
	) name8189 (
		_w8246_,
		_w8254_,
		_w8255_
	);
	LUT3 #(
		.INIT('h0d)
	) name8190 (
		_w8221_,
		_w8222_,
		_w8223_,
		_w8256_
	);
	LUT3 #(
		.INIT('h0d)
	) name8191 (
		_w8207_,
		_w8208_,
		_w8209_,
		_w8257_
	);
	LUT2 #(
		.INIT('h8)
	) name8192 (
		\a[48] ,
		\a[59] ,
		_w8258_
	);
	LUT4 #(
		.INIT('h153f)
	) name8193 (
		\a[44] ,
		\a[49] ,
		\a[58] ,
		\a[63] ,
		_w8259_
	);
	LUT2 #(
		.INIT('h8)
	) name8194 (
		\a[49] ,
		\a[63] ,
		_w8260_
	);
	LUT4 #(
		.INIT('h8000)
	) name8195 (
		\a[44] ,
		\a[49] ,
		\a[58] ,
		\a[63] ,
		_w8261_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8196 (
		\a[44] ,
		\a[49] ,
		\a[58] ,
		\a[63] ,
		_w8262_
	);
	LUT2 #(
		.INIT('h6)
	) name8197 (
		_w8258_,
		_w8262_,
		_w8263_
	);
	LUT3 #(
		.INIT('h69)
	) name8198 (
		_w8256_,
		_w8257_,
		_w8263_,
		_w8264_
	);
	LUT2 #(
		.INIT('h2)
	) name8199 (
		_w8255_,
		_w8264_,
		_w8265_
	);
	LUT2 #(
		.INIT('h4)
	) name8200 (
		_w8255_,
		_w8264_,
		_w8266_
	);
	LUT2 #(
		.INIT('h9)
	) name8201 (
		_w8255_,
		_w8264_,
		_w8267_
	);
	LUT2 #(
		.INIT('h6)
	) name8202 (
		_w8243_,
		_w8267_,
		_w8268_
	);
	LUT4 #(
		.INIT('he11e)
	) name8203 (
		_w8227_,
		_w8229_,
		_w8242_,
		_w8268_,
		_w8269_
	);
	LUT2 #(
		.INIT('h1)
	) name8204 (
		_w8238_,
		_w8269_,
		_w8270_
	);
	LUT2 #(
		.INIT('h8)
	) name8205 (
		_w8238_,
		_w8269_,
		_w8271_
	);
	LUT2 #(
		.INIT('h6)
	) name8206 (
		_w8238_,
		_w8269_,
		_w8272_
	);
	LUT3 #(
		.INIT('h0b)
	) name8207 (
		_w8182_,
		_w8183_,
		_w8232_,
		_w8273_
	);
	LUT2 #(
		.INIT('h4)
	) name8208 (
		_w8133_,
		_w8273_,
		_w8274_
	);
	LUT3 #(
		.INIT('h02)
	) name8209 (
		_w8182_,
		_w8183_,
		_w8232_,
		_w8275_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8210 (
		_w8182_,
		_w8183_,
		_w8232_,
		_w8233_,
		_w8276_
	);
	LUT4 #(
		.INIT('h63cc)
	) name8211 (
		_w8141_,
		_w8272_,
		_w8274_,
		_w8276_,
		_w8277_
	);
	LUT2 #(
		.INIT('h1)
	) name8212 (
		_w8233_,
		_w8270_,
		_w8278_
	);
	LUT2 #(
		.INIT('h4)
	) name8213 (
		_w8275_,
		_w8278_,
		_w8279_
	);
	LUT4 #(
		.INIT('h011f)
	) name8214 (
		_w8227_,
		_w8229_,
		_w8242_,
		_w8268_,
		_w8280_
	);
	LUT3 #(
		.INIT('h0d)
	) name8215 (
		_w8246_,
		_w8252_,
		_w8253_,
		_w8281_
	);
	LUT2 #(
		.INIT('h8)
	) name8216 (
		\a[51] ,
		\a[57] ,
		_w8282_
	);
	LUT4 #(
		.INIT('h153f)
	) name8217 (
		\a[52] ,
		\a[53] ,
		\a[55] ,
		\a[56] ,
		_w8283_
	);
	LUT4 #(
		.INIT('h8000)
	) name8218 (
		\a[52] ,
		\a[53] ,
		\a[55] ,
		\a[56] ,
		_w8284_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8219 (
		\a[52] ,
		\a[53] ,
		\a[55] ,
		\a[56] ,
		_w8285_
	);
	LUT2 #(
		.INIT('h6)
	) name8220 (
		_w8282_,
		_w8285_,
		_w8286_
	);
	LUT4 #(
		.INIT('h7100)
	) name8221 (
		_w8256_,
		_w8257_,
		_w8263_,
		_w8286_,
		_w8287_
	);
	LUT4 #(
		.INIT('h008e)
	) name8222 (
		_w8256_,
		_w8257_,
		_w8263_,
		_w8286_,
		_w8288_
	);
	LUT4 #(
		.INIT('h8e71)
	) name8223 (
		_w8256_,
		_w8257_,
		_w8263_,
		_w8286_,
		_w8289_
	);
	LUT2 #(
		.INIT('h6)
	) name8224 (
		_w8281_,
		_w8289_,
		_w8290_
	);
	LUT4 #(
		.INIT('hd00d)
	) name8225 (
		_w8255_,
		_w8264_,
		_w8281_,
		_w8289_,
		_w8291_
	);
	LUT3 #(
		.INIT('h70)
	) name8226 (
		_w8243_,
		_w8267_,
		_w8291_,
		_w8292_
	);
	LUT4 #(
		.INIT('h8e00)
	) name8227 (
		_w8243_,
		_w8255_,
		_w8264_,
		_w8290_,
		_w8293_
	);
	LUT4 #(
		.INIT('h31ce)
	) name8228 (
		_w8243_,
		_w8265_,
		_w8266_,
		_w8290_,
		_w8294_
	);
	LUT3 #(
		.INIT('h13)
	) name8229 (
		\a[45] ,
		\a[53] ,
		\a[62] ,
		_w8295_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8230 (
		\a[45] ,
		\a[53] ,
		\a[54] ,
		\a[62] ,
		_w8296_
	);
	LUT3 #(
		.INIT('h0d)
	) name8231 (
		_w8247_,
		_w8248_,
		_w8249_,
		_w8297_
	);
	LUT4 #(
		.INIT('hf20d)
	) name8232 (
		_w8247_,
		_w8248_,
		_w8249_,
		_w8296_,
		_w8298_
	);
	LUT3 #(
		.INIT('h0d)
	) name8233 (
		_w8258_,
		_w8259_,
		_w8261_,
		_w8299_
	);
	LUT2 #(
		.INIT('h9)
	) name8234 (
		_w8298_,
		_w8299_,
		_w8300_
	);
	LUT3 #(
		.INIT('hd0)
	) name8235 (
		_w8239_,
		_w8240_,
		_w8300_,
		_w8301_
	);
	LUT3 #(
		.INIT('h0b)
	) name8236 (
		_w8239_,
		_w8240_,
		_w8300_,
		_w8302_
	);
	LUT4 #(
		.INIT('h1101)
	) name8237 (
		_w8215_,
		_w8217_,
		_w8239_,
		_w8240_,
		_w8303_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name8238 (
		_w8241_,
		_w8301_,
		_w8302_,
		_w8303_,
		_w8304_
	);
	LUT4 #(
		.INIT('h153f)
	) name8239 (
		\a[46] ,
		\a[47] ,
		\a[60] ,
		\a[61] ,
		_w8305_
	);
	LUT4 #(
		.INIT('h000d)
	) name8240 (
		_w8211_,
		_w8212_,
		_w8213_,
		_w8244_,
		_w8306_
	);
	LUT2 #(
		.INIT('h8)
	) name8241 (
		\a[45] ,
		\a[63] ,
		_w8307_
	);
	LUT4 #(
		.INIT('h153f)
	) name8242 (
		\a[46] ,
		\a[47] ,
		\a[61] ,
		\a[62] ,
		_w8308_
	);
	LUT4 #(
		.INIT('h8000)
	) name8243 (
		\a[46] ,
		\a[47] ,
		\a[61] ,
		\a[62] ,
		_w8309_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8244 (
		\a[46] ,
		\a[47] ,
		\a[61] ,
		\a[62] ,
		_w8310_
	);
	LUT2 #(
		.INIT('h6)
	) name8245 (
		_w8307_,
		_w8310_,
		_w8311_
	);
	LUT2 #(
		.INIT('h8)
	) name8246 (
		\a[48] ,
		\a[60] ,
		_w8312_
	);
	LUT4 #(
		.INIT('h153f)
	) name8247 (
		\a[49] ,
		\a[50] ,
		\a[58] ,
		\a[59] ,
		_w8313_
	);
	LUT4 #(
		.INIT('h8000)
	) name8248 (
		\a[49] ,
		\a[50] ,
		\a[58] ,
		\a[59] ,
		_w8314_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8249 (
		\a[49] ,
		\a[50] ,
		\a[58] ,
		\a[59] ,
		_w8315_
	);
	LUT2 #(
		.INIT('h6)
	) name8250 (
		_w8312_,
		_w8315_,
		_w8316_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name8251 (
		_w8305_,
		_w8306_,
		_w8311_,
		_w8316_,
		_w8317_
	);
	LUT3 #(
		.INIT('h96)
	) name8252 (
		_w8294_,
		_w8304_,
		_w8317_,
		_w8318_
	);
	LUT2 #(
		.INIT('h2)
	) name8253 (
		_w8280_,
		_w8318_,
		_w8319_
	);
	LUT2 #(
		.INIT('h4)
	) name8254 (
		_w8280_,
		_w8318_,
		_w8320_
	);
	LUT2 #(
		.INIT('h9)
	) name8255 (
		_w8280_,
		_w8318_,
		_w8321_
	);
	LUT4 #(
		.INIT('h7007)
	) name8256 (
		_w8238_,
		_w8269_,
		_w8280_,
		_w8318_,
		_w8322_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8257 (
		_w8141_,
		_w8274_,
		_w8279_,
		_w8322_,
		_w8323_
	);
	LUT4 #(
		.INIT('h1033)
	) name8258 (
		_w8141_,
		_w8271_,
		_w8274_,
		_w8279_,
		_w8324_
	);
	LUT3 #(
		.INIT('hcd)
	) name8259 (
		_w8321_,
		_w8323_,
		_w8324_,
		_w8325_
	);
	LUT4 #(
		.INIT('h7077)
	) name8260 (
		_w8238_,
		_w8269_,
		_w8280_,
		_w8318_,
		_w8326_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8261 (
		_w8141_,
		_w8274_,
		_w8279_,
		_w8326_,
		_w8327_
	);
	LUT4 #(
		.INIT('h4554)
	) name8262 (
		_w8292_,
		_w8293_,
		_w8304_,
		_w8317_,
		_w8328_
	);
	LUT4 #(
		.INIT('hf110)
	) name8263 (
		_w8305_,
		_w8306_,
		_w8311_,
		_w8316_,
		_w8329_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8264 (
		\a[47] ,
		\a[54] ,
		\a[55] ,
		\a[62] ,
		_w8330_
	);
	LUT4 #(
		.INIT('hff2b)
	) name8265 (
		_w8296_,
		_w8297_,
		_w8299_,
		_w8330_,
		_w8331_
	);
	LUT3 #(
		.INIT('h80)
	) name8266 (
		\a[47] ,
		\a[54] ,
		\a[62] ,
		_w8332_
	);
	LUT2 #(
		.INIT('h4)
	) name8267 (
		_w8295_,
		_w8332_,
		_w8333_
	);
	LUT4 #(
		.INIT('h88ef)
	) name8268 (
		_w8297_,
		_w8299_,
		_w8330_,
		_w8333_,
		_w8334_
	);
	LUT3 #(
		.INIT('h6a)
	) name8269 (
		_w8329_,
		_w8331_,
		_w8334_,
		_w8335_
	);
	LUT3 #(
		.INIT('h0d)
	) name8270 (
		_w8302_,
		_w8303_,
		_w8317_,
		_w8336_
	);
	LUT4 #(
		.INIT('h4404)
	) name8271 (
		_w8241_,
		_w8301_,
		_w8302_,
		_w8303_,
		_w8337_
	);
	LUT3 #(
		.INIT('h54)
	) name8272 (
		_w8335_,
		_w8336_,
		_w8337_,
		_w8338_
	);
	LUT3 #(
		.INIT('h20)
	) name8273 (
		_w8302_,
		_w8303_,
		_w8335_,
		_w8339_
	);
	LUT4 #(
		.INIT('h2888)
	) name8274 (
		_w8317_,
		_w8329_,
		_w8331_,
		_w8334_,
		_w8340_
	);
	LUT3 #(
		.INIT('hb0)
	) name8275 (
		_w8241_,
		_w8301_,
		_w8340_,
		_w8341_
	);
	LUT2 #(
		.INIT('h1)
	) name8276 (
		_w8339_,
		_w8341_,
		_w8342_
	);
	LUT2 #(
		.INIT('h8)
	) name8277 (
		\a[46] ,
		\a[63] ,
		_w8343_
	);
	LUT4 #(
		.INIT('h0dff)
	) name8278 (
		_w8282_,
		_w8283_,
		_w8284_,
		_w8343_,
		_w8344_
	);
	LUT4 #(
		.INIT('h000d)
	) name8279 (
		_w8282_,
		_w8283_,
		_w8284_,
		_w8343_,
		_w8345_
	);
	LUT4 #(
		.INIT('h0df2)
	) name8280 (
		_w8282_,
		_w8283_,
		_w8284_,
		_w8343_,
		_w8346_
	);
	LUT3 #(
		.INIT('h0d)
	) name8281 (
		_w8312_,
		_w8313_,
		_w8314_,
		_w8347_
	);
	LUT2 #(
		.INIT('h6)
	) name8282 (
		_w8346_,
		_w8347_,
		_w8348_
	);
	LUT3 #(
		.INIT('h0e)
	) name8283 (
		_w8281_,
		_w8287_,
		_w8288_,
		_w8349_
	);
	LUT4 #(
		.INIT('hf100)
	) name8284 (
		_w8281_,
		_w8287_,
		_w8288_,
		_w8348_,
		_w8350_
	);
	LUT4 #(
		.INIT('hff31)
	) name8285 (
		_w8281_,
		_w8287_,
		_w8288_,
		_w8348_,
		_w8351_
	);
	LUT2 #(
		.INIT('h8)
	) name8286 (
		\a[48] ,
		\a[61] ,
		_w8352_
	);
	LUT4 #(
		.INIT('h153f)
	) name8287 (
		\a[49] ,
		\a[50] ,
		\a[59] ,
		\a[60] ,
		_w8353_
	);
	LUT4 #(
		.INIT('h8000)
	) name8288 (
		\a[49] ,
		\a[50] ,
		\a[59] ,
		\a[60] ,
		_w8354_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8289 (
		\a[49] ,
		\a[50] ,
		\a[59] ,
		\a[60] ,
		_w8355_
	);
	LUT2 #(
		.INIT('h6)
	) name8290 (
		_w8352_,
		_w8355_,
		_w8356_
	);
	LUT3 #(
		.INIT('h0d)
	) name8291 (
		_w8307_,
		_w8308_,
		_w8309_,
		_w8357_
	);
	LUT2 #(
		.INIT('h8)
	) name8292 (
		\a[51] ,
		\a[58] ,
		_w8358_
	);
	LUT4 #(
		.INIT('h153f)
	) name8293 (
		\a[52] ,
		\a[53] ,
		\a[56] ,
		\a[57] ,
		_w8359_
	);
	LUT4 #(
		.INIT('h8000)
	) name8294 (
		\a[52] ,
		\a[53] ,
		\a[56] ,
		\a[57] ,
		_w8360_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8295 (
		\a[52] ,
		\a[53] ,
		\a[56] ,
		\a[57] ,
		_w8361_
	);
	LUT2 #(
		.INIT('h6)
	) name8296 (
		_w8358_,
		_w8361_,
		_w8362_
	);
	LUT3 #(
		.INIT('h69)
	) name8297 (
		_w8356_,
		_w8357_,
		_w8362_,
		_w8363_
	);
	LUT3 #(
		.INIT('h40)
	) name8298 (
		_w8350_,
		_w8351_,
		_w8363_,
		_w8364_
	);
	LUT4 #(
		.INIT('h000e)
	) name8299 (
		_w8281_,
		_w8287_,
		_w8288_,
		_w8348_,
		_w8365_
	);
	LUT4 #(
		.INIT('hf0fd)
	) name8300 (
		_w8348_,
		_w8349_,
		_w8363_,
		_w8365_,
		_w8366_
	);
	LUT2 #(
		.INIT('h4)
	) name8301 (
		_w8364_,
		_w8366_,
		_w8367_
	);
	LUT4 #(
		.INIT('h0100)
	) name8302 (
		_w8339_,
		_w8341_,
		_w8364_,
		_w8366_,
		_w8368_
	);
	LUT4 #(
		.INIT('h8a20)
	) name8303 (
		_w8328_,
		_w8338_,
		_w8342_,
		_w8367_,
		_w8369_
	);
	LUT4 #(
		.INIT('h1045)
	) name8304 (
		_w8328_,
		_w8338_,
		_w8342_,
		_w8367_,
		_w8370_
	);
	LUT4 #(
		.INIT('h659a)
	) name8305 (
		_w8328_,
		_w8338_,
		_w8342_,
		_w8367_,
		_w8371_
	);
	LUT3 #(
		.INIT('he1)
	) name8306 (
		_w8319_,
		_w8327_,
		_w8371_,
		_w8372_
	);
	LUT3 #(
		.INIT('h02)
	) name8307 (
		_w8319_,
		_w8320_,
		_w8369_,
		_w8373_
	);
	LUT3 #(
		.INIT('h01)
	) name8308 (
		_w8271_,
		_w8320_,
		_w8369_,
		_w8374_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8309 (
		_w8141_,
		_w8274_,
		_w8279_,
		_w8374_,
		_w8375_
	);
	LUT3 #(
		.INIT('hb2)
	) name8310 (
		_w8356_,
		_w8357_,
		_w8362_,
		_w8376_
	);
	LUT3 #(
		.INIT('h0d)
	) name8311 (
		_w8352_,
		_w8353_,
		_w8354_,
		_w8377_
	);
	LUT3 #(
		.INIT('h0d)
	) name8312 (
		_w8358_,
		_w8359_,
		_w8360_,
		_w8378_
	);
	LUT2 #(
		.INIT('h8)
	) name8313 (
		\a[49] ,
		\a[61] ,
		_w8379_
	);
	LUT4 #(
		.INIT('h153f)
	) name8314 (
		\a[50] ,
		\a[51] ,
		\a[59] ,
		\a[60] ,
		_w8380_
	);
	LUT4 #(
		.INIT('h8000)
	) name8315 (
		\a[50] ,
		\a[51] ,
		\a[59] ,
		\a[60] ,
		_w8381_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8316 (
		\a[50] ,
		\a[51] ,
		\a[59] ,
		\a[60] ,
		_w8382_
	);
	LUT2 #(
		.INIT('h6)
	) name8317 (
		_w8379_,
		_w8382_,
		_w8383_
	);
	LUT3 #(
		.INIT('h69)
	) name8318 (
		_w8377_,
		_w8378_,
		_w8383_,
		_w8384_
	);
	LUT2 #(
		.INIT('h9)
	) name8319 (
		_w8376_,
		_w8384_,
		_w8385_
	);
	LUT3 #(
		.INIT('h70)
	) name8320 (
		_w8329_,
		_w8331_,
		_w8334_,
		_w8386_
	);
	LUT2 #(
		.INIT('h9)
	) name8321 (
		_w8385_,
		_w8386_,
		_w8387_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8322 (
		\a[47] ,
		\a[54] ,
		\a[55] ,
		\a[62] ,
		_w8388_
	);
	LUT4 #(
		.INIT('h153f)
	) name8323 (
		\a[47] ,
		\a[48] ,
		\a[62] ,
		\a[63] ,
		_w8389_
	);
	LUT2 #(
		.INIT('h8)
	) name8324 (
		\a[48] ,
		\a[63] ,
		_w8390_
	);
	LUT4 #(
		.INIT('h8000)
	) name8325 (
		\a[47] ,
		\a[48] ,
		\a[62] ,
		\a[63] ,
		_w8391_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8326 (
		\a[47] ,
		\a[48] ,
		\a[62] ,
		\a[63] ,
		_w8392_
	);
	LUT2 #(
		.INIT('h8)
	) name8327 (
		\a[52] ,
		\a[58] ,
		_w8393_
	);
	LUT4 #(
		.INIT('h153f)
	) name8328 (
		\a[53] ,
		\a[54] ,
		\a[56] ,
		\a[57] ,
		_w8394_
	);
	LUT4 #(
		.INIT('h8000)
	) name8329 (
		\a[53] ,
		\a[54] ,
		\a[56] ,
		\a[57] ,
		_w8395_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8330 (
		\a[53] ,
		\a[54] ,
		\a[56] ,
		\a[57] ,
		_w8396_
	);
	LUT4 #(
		.INIT('h0660)
	) name8331 (
		_w8388_,
		_w8392_,
		_w8393_,
		_w8396_,
		_w8397_
	);
	LUT4 #(
		.INIT('h9009)
	) name8332 (
		_w8388_,
		_w8392_,
		_w8393_,
		_w8396_,
		_w8398_
	);
	LUT4 #(
		.INIT('h6996)
	) name8333 (
		_w8388_,
		_w8392_,
		_w8393_,
		_w8396_,
		_w8399_
	);
	LUT4 #(
		.INIT('hf807)
	) name8334 (
		_w8344_,
		_w8347_,
		_w8345_,
		_w8399_,
		_w8400_
	);
	LUT4 #(
		.INIT('h8cff)
	) name8335 (
		_w8350_,
		_w8351_,
		_w8363_,
		_w8400_,
		_w8401_
	);
	LUT4 #(
		.INIT('h008c)
	) name8336 (
		_w8350_,
		_w8351_,
		_w8363_,
		_w8400_,
		_w8402_
	);
	LUT4 #(
		.INIT('h8c73)
	) name8337 (
		_w8350_,
		_w8351_,
		_w8363_,
		_w8400_,
		_w8403_
	);
	LUT2 #(
		.INIT('h6)
	) name8338 (
		_w8387_,
		_w8403_,
		_w8404_
	);
	LUT4 #(
		.INIT('h008c)
	) name8339 (
		_w8338_,
		_w8342_,
		_w8368_,
		_w8404_,
		_w8405_
	);
	LUT4 #(
		.INIT('h7300)
	) name8340 (
		_w8338_,
		_w8342_,
		_w8368_,
		_w8404_,
		_w8406_
	);
	LUT4 #(
		.INIT('h8c73)
	) name8341 (
		_w8338_,
		_w8342_,
		_w8367_,
		_w8404_,
		_w8407_
	);
	LUT4 #(
		.INIT('hfe01)
	) name8342 (
		_w8370_,
		_w8373_,
		_w8375_,
		_w8407_,
		_w8408_
	);
	LUT2 #(
		.INIT('h1)
	) name8343 (
		_w8370_,
		_w8405_,
		_w8409_
	);
	LUT3 #(
		.INIT('hc4)
	) name8344 (
		_w8387_,
		_w8401_,
		_w8402_,
		_w8410_
	);
	LUT4 #(
		.INIT('h153f)
	) name8345 (
		\a[50] ,
		\a[51] ,
		\a[60] ,
		\a[61] ,
		_w8411_
	);
	LUT4 #(
		.INIT('h8000)
	) name8346 (
		\a[50] ,
		\a[51] ,
		\a[60] ,
		\a[61] ,
		_w8412_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8347 (
		\a[50] ,
		\a[51] ,
		\a[60] ,
		\a[61] ,
		_w8413_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8348 (
		\a[49] ,
		\a[55] ,
		\a[56] ,
		\a[62] ,
		_w8414_
	);
	LUT3 #(
		.INIT('h60)
	) name8349 (
		_w8390_,
		_w8413_,
		_w8414_,
		_w8415_
	);
	LUT3 #(
		.INIT('h09)
	) name8350 (
		_w8390_,
		_w8413_,
		_w8414_,
		_w8416_
	);
	LUT3 #(
		.INIT('h96)
	) name8351 (
		_w8390_,
		_w8413_,
		_w8414_,
		_w8417_
	);
	LUT2 #(
		.INIT('h8)
	) name8352 (
		\a[52] ,
		\a[59] ,
		_w8418_
	);
	LUT4 #(
		.INIT('h153f)
	) name8353 (
		\a[53] ,
		\a[54] ,
		\a[57] ,
		\a[58] ,
		_w8419_
	);
	LUT4 #(
		.INIT('h8000)
	) name8354 (
		\a[53] ,
		\a[54] ,
		\a[57] ,
		\a[58] ,
		_w8420_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8355 (
		\a[53] ,
		\a[54] ,
		\a[57] ,
		\a[58] ,
		_w8421_
	);
	LUT2 #(
		.INIT('h6)
	) name8356 (
		_w8418_,
		_w8421_,
		_w8422_
	);
	LUT2 #(
		.INIT('h6)
	) name8357 (
		_w8417_,
		_w8422_,
		_w8423_
	);
	LUT4 #(
		.INIT('h2b00)
	) name8358 (
		_w8376_,
		_w8384_,
		_w8386_,
		_w8423_,
		_w8424_
	);
	LUT3 #(
		.INIT('h0d)
	) name8359 (
		_w8379_,
		_w8380_,
		_w8381_,
		_w8425_
	);
	LUT3 #(
		.INIT('h0d)
	) name8360 (
		_w8393_,
		_w8394_,
		_w8395_,
		_w8426_
	);
	LUT3 #(
		.INIT('h0d)
	) name8361 (
		_w8388_,
		_w8389_,
		_w8391_,
		_w8427_
	);
	LUT3 #(
		.INIT('h96)
	) name8362 (
		_w8425_,
		_w8426_,
		_w8427_,
		_w8428_
	);
	LUT3 #(
		.INIT('h8e)
	) name8363 (
		_w8377_,
		_w8378_,
		_w8383_,
		_w8429_
	);
	LUT2 #(
		.INIT('h8)
	) name8364 (
		_w8428_,
		_w8429_,
		_w8430_
	);
	LUT4 #(
		.INIT('h00a8)
	) name8365 (
		_w8344_,
		_w8345_,
		_w8347_,
		_w8397_,
		_w8431_
	);
	LUT4 #(
		.INIT('h3c69)
	) name8366 (
		_w8398_,
		_w8428_,
		_w8429_,
		_w8431_,
		_w8432_
	);
	LUT3 #(
		.INIT('h0d)
	) name8367 (
		_w8376_,
		_w8384_,
		_w8423_,
		_w8433_
	);
	LUT3 #(
		.INIT('hd0)
	) name8368 (
		_w8385_,
		_w8386_,
		_w8433_,
		_w8434_
	);
	LUT4 #(
		.INIT('h20f0)
	) name8369 (
		_w8385_,
		_w8386_,
		_w8432_,
		_w8433_,
		_w8435_
	);
	LUT3 #(
		.INIT('hc9)
	) name8370 (
		_w8424_,
		_w8432_,
		_w8434_,
		_w8436_
	);
	LUT2 #(
		.INIT('h4)
	) name8371 (
		_w8410_,
		_w8436_,
		_w8437_
	);
	LUT2 #(
		.INIT('h9)
	) name8372 (
		_w8410_,
		_w8436_,
		_w8438_
	);
	LUT2 #(
		.INIT('h4)
	) name8373 (
		_w8406_,
		_w8438_,
		_w8439_
	);
	LUT4 #(
		.INIT('hef00)
	) name8374 (
		_w8373_,
		_w8375_,
		_w8409_,
		_w8439_,
		_w8440_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name8375 (
		_w8373_,
		_w8375_,
		_w8406_,
		_w8409_,
		_w8441_
	);
	LUT3 #(
		.INIT('hcd)
	) name8376 (
		_w8438_,
		_w8440_,
		_w8441_,
		_w8442_
	);
	LUT2 #(
		.INIT('h1)
	) name8377 (
		_w8406_,
		_w8437_,
		_w8443_
	);
	LUT4 #(
		.INIT('hef00)
	) name8378 (
		_w8373_,
		_w8375_,
		_w8409_,
		_w8443_,
		_w8444_
	);
	LUT4 #(
		.INIT('hfca8)
	) name8379 (
		_w8398_,
		_w8428_,
		_w8429_,
		_w8431_,
		_w8445_
	);
	LUT4 #(
		.INIT('h153f)
	) name8380 (
		\a[51] ,
		\a[52] ,
		\a[60] ,
		\a[61] ,
		_w8446_
	);
	LUT4 #(
		.INIT('h8000)
	) name8381 (
		\a[51] ,
		\a[52] ,
		\a[60] ,
		\a[61] ,
		_w8447_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8382 (
		\a[51] ,
		\a[52] ,
		\a[60] ,
		\a[61] ,
		_w8448_
	);
	LUT2 #(
		.INIT('h6)
	) name8383 (
		_w8260_,
		_w8448_,
		_w8449_
	);
	LUT3 #(
		.INIT('h0d)
	) name8384 (
		_w8390_,
		_w8411_,
		_w8412_,
		_w8450_
	);
	LUT2 #(
		.INIT('h8)
	) name8385 (
		\a[53] ,
		\a[59] ,
		_w8451_
	);
	LUT4 #(
		.INIT('h153f)
	) name8386 (
		\a[54] ,
		\a[55] ,
		\a[57] ,
		\a[58] ,
		_w8452_
	);
	LUT4 #(
		.INIT('h8000)
	) name8387 (
		\a[54] ,
		\a[55] ,
		\a[57] ,
		\a[58] ,
		_w8453_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8388 (
		\a[54] ,
		\a[55] ,
		\a[57] ,
		\a[58] ,
		_w8454_
	);
	LUT2 #(
		.INIT('h6)
	) name8389 (
		_w8451_,
		_w8454_,
		_w8455_
	);
	LUT3 #(
		.INIT('h69)
	) name8390 (
		_w8449_,
		_w8450_,
		_w8455_,
		_w8456_
	);
	LUT3 #(
		.INIT('h32)
	) name8391 (
		_w8415_,
		_w8416_,
		_w8422_,
		_w8457_
	);
	LUT3 #(
		.INIT('h13)
	) name8392 (
		\a[49] ,
		\a[55] ,
		\a[62] ,
		_w8458_
	);
	LUT2 #(
		.INIT('h8)
	) name8393 (
		\a[50] ,
		\a[62] ,
		_w8459_
	);
	LUT3 #(
		.INIT('h80)
	) name8394 (
		\a[50] ,
		\a[56] ,
		\a[62] ,
		_w8460_
	);
	LUT2 #(
		.INIT('h4)
	) name8395 (
		_w8458_,
		_w8460_,
		_w8461_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8396 (
		\a[49] ,
		\a[55] ,
		\a[56] ,
		\a[62] ,
		_w8462_
	);
	LUT2 #(
		.INIT('h1)
	) name8397 (
		_w8459_,
		_w8462_,
		_w8463_
	);
	LUT3 #(
		.INIT('hd2)
	) name8398 (
		\a[56] ,
		_w8458_,
		_w8459_,
		_w8464_
	);
	LUT3 #(
		.INIT('h0d)
	) name8399 (
		_w8418_,
		_w8419_,
		_w8420_,
		_w8465_
	);
	LUT2 #(
		.INIT('h6)
	) name8400 (
		_w8464_,
		_w8465_,
		_w8466_
	);
	LUT3 #(
		.INIT('h17)
	) name8401 (
		_w8425_,
		_w8426_,
		_w8427_,
		_w8467_
	);
	LUT3 #(
		.INIT('h69)
	) name8402 (
		_w8457_,
		_w8466_,
		_w8467_,
		_w8468_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name8403 (
		_w8430_,
		_w8445_,
		_w8456_,
		_w8468_,
		_w8469_
	);
	LUT3 #(
		.INIT('h01)
	) name8404 (
		_w8424_,
		_w8435_,
		_w8469_,
		_w8470_
	);
	LUT3 #(
		.INIT('he0)
	) name8405 (
		_w8424_,
		_w8435_,
		_w8469_,
		_w8471_
	);
	LUT3 #(
		.INIT('h1e)
	) name8406 (
		_w8424_,
		_w8435_,
		_w8469_,
		_w8472_
	);
	LUT3 #(
		.INIT('h2d)
	) name8407 (
		_w8410_,
		_w8436_,
		_w8472_,
		_w8473_
	);
	LUT3 #(
		.INIT('hf0)
	) name8408 (
		_w8410_,
		_w8436_,
		_w8472_,
		_w8474_
	);
	LUT3 #(
		.INIT('he4)
	) name8409 (
		_w8444_,
		_w8473_,
		_w8474_,
		_w8475_
	);
	LUT4 #(
		.INIT('hf110)
	) name8410 (
		_w8430_,
		_w8445_,
		_w8456_,
		_w8468_,
		_w8476_
	);
	LUT3 #(
		.INIT('h4d)
	) name8411 (
		_w8457_,
		_w8466_,
		_w8467_,
		_w8477_
	);
	LUT2 #(
		.INIT('h8)
	) name8412 (
		\a[50] ,
		\a[63] ,
		_w8478_
	);
	LUT4 #(
		.INIT('h153f)
	) name8413 (
		\a[54] ,
		\a[55] ,
		\a[58] ,
		\a[59] ,
		_w8479_
	);
	LUT4 #(
		.INIT('h8000)
	) name8414 (
		\a[54] ,
		\a[55] ,
		\a[58] ,
		\a[59] ,
		_w8480_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8415 (
		\a[54] ,
		\a[55] ,
		\a[58] ,
		\a[59] ,
		_w8481_
	);
	LUT2 #(
		.INIT('h6)
	) name8416 (
		_w8478_,
		_w8481_,
		_w8482_
	);
	LUT3 #(
		.INIT('h0d)
	) name8417 (
		_w8260_,
		_w8446_,
		_w8447_,
		_w8483_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8418 (
		\a[51] ,
		\a[56] ,
		\a[57] ,
		\a[62] ,
		_w8484_
	);
	LUT3 #(
		.INIT('h69)
	) name8419 (
		_w8482_,
		_w8483_,
		_w8484_,
		_w8485_
	);
	LUT4 #(
		.INIT('hb200)
	) name8420 (
		_w8457_,
		_w8466_,
		_w8467_,
		_w8485_,
		_w8486_
	);
	LUT3 #(
		.INIT('h23)
	) name8421 (
		_w8461_,
		_w8463_,
		_w8465_,
		_w8487_
	);
	LUT4 #(
		.INIT('h8000)
	) name8422 (
		\a[52] ,
		\a[53] ,
		\a[60] ,
		\a[61] ,
		_w8488_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8423 (
		\a[52] ,
		\a[53] ,
		\a[60] ,
		\a[61] ,
		_w8489_
	);
	LUT4 #(
		.INIT('hf20d)
	) name8424 (
		_w8451_,
		_w8452_,
		_w8453_,
		_w8489_,
		_w8490_
	);
	LUT4 #(
		.INIT('hdc00)
	) name8425 (
		_w8461_,
		_w8463_,
		_w8465_,
		_w8490_,
		_w8491_
	);
	LUT4 #(
		.INIT('h0023)
	) name8426 (
		_w8461_,
		_w8463_,
		_w8465_,
		_w8490_,
		_w8492_
	);
	LUT4 #(
		.INIT('h23dc)
	) name8427 (
		_w8461_,
		_w8463_,
		_w8465_,
		_w8490_,
		_w8493_
	);
	LUT3 #(
		.INIT('hb2)
	) name8428 (
		_w8449_,
		_w8450_,
		_w8455_,
		_w8494_
	);
	LUT2 #(
		.INIT('h6)
	) name8429 (
		_w8493_,
		_w8494_,
		_w8495_
	);
	LUT4 #(
		.INIT('h004d)
	) name8430 (
		_w8457_,
		_w8466_,
		_w8467_,
		_w8485_,
		_w8496_
	);
	LUT4 #(
		.INIT('hf949)
	) name8431 (
		_w8477_,
		_w8485_,
		_w8495_,
		_w8496_,
		_w8497_
	);
	LUT2 #(
		.INIT('h1)
	) name8432 (
		_w8476_,
		_w8497_,
		_w8498_
	);
	LUT2 #(
		.INIT('h8)
	) name8433 (
		_w8476_,
		_w8497_,
		_w8499_
	);
	LUT2 #(
		.INIT('h6)
	) name8434 (
		_w8476_,
		_w8497_,
		_w8500_
	);
	LUT3 #(
		.INIT('h02)
	) name8435 (
		_w8410_,
		_w8436_,
		_w8471_,
		_w8501_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name8436 (
		_w8410_,
		_w8436_,
		_w8470_,
		_w8471_,
		_w8502_
	);
	LUT4 #(
		.INIT('h20f0)
	) name8437 (
		_w8444_,
		_w8471_,
		_w8500_,
		_w8502_,
		_w8503_
	);
	LUT2 #(
		.INIT('h1)
	) name8438 (
		_w8470_,
		_w8500_,
		_w8504_
	);
	LUT2 #(
		.INIT('h4)
	) name8439 (
		_w8501_,
		_w8504_,
		_w8505_
	);
	LUT3 #(
		.INIT('hd0)
	) name8440 (
		_w8444_,
		_w8471_,
		_w8505_,
		_w8506_
	);
	LUT2 #(
		.INIT('he)
	) name8441 (
		_w8503_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h1)
	) name8442 (
		_w8470_,
		_w8498_,
		_w8508_
	);
	LUT2 #(
		.INIT('h4)
	) name8443 (
		_w8501_,
		_w8508_,
		_w8509_
	);
	LUT3 #(
		.INIT('h51)
	) name8444 (
		_w8486_,
		_w8495_,
		_w8496_,
		_w8510_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8445 (
		\a[51] ,
		\a[56] ,
		\a[57] ,
		\a[62] ,
		_w8511_
	);
	LUT4 #(
		.INIT('h000d)
	) name8446 (
		_w8478_,
		_w8479_,
		_w8480_,
		_w8511_,
		_w8512_
	);
	LUT4 #(
		.INIT('hf200)
	) name8447 (
		_w8478_,
		_w8479_,
		_w8480_,
		_w8511_,
		_w8513_
	);
	LUT4 #(
		.INIT('h0df2)
	) name8448 (
		_w8478_,
		_w8479_,
		_w8480_,
		_w8511_,
		_w8514_
	);
	LUT4 #(
		.INIT('h153f)
	) name8449 (
		\a[52] ,
		\a[53] ,
		\a[60] ,
		\a[61] ,
		_w8515_
	);
	LUT4 #(
		.INIT('h000d)
	) name8450 (
		_w8451_,
		_w8452_,
		_w8453_,
		_w8488_,
		_w8516_
	);
	LUT3 #(
		.INIT('ha9)
	) name8451 (
		_w8514_,
		_w8515_,
		_w8516_,
		_w8517_
	);
	LUT4 #(
		.INIT('hb200)
	) name8452 (
		_w8487_,
		_w8490_,
		_w8494_,
		_w8517_,
		_w8518_
	);
	LUT4 #(
		.INIT('h0023)
	) name8453 (
		_w8491_,
		_w8492_,
		_w8494_,
		_w8517_,
		_w8519_
	);
	LUT2 #(
		.INIT('h8)
	) name8454 (
		\a[51] ,
		\a[63] ,
		_w8520_
	);
	LUT4 #(
		.INIT('h153f)
	) name8455 (
		\a[52] ,
		\a[53] ,
		\a[61] ,
		\a[62] ,
		_w8521_
	);
	LUT4 #(
		.INIT('h8000)
	) name8456 (
		\a[52] ,
		\a[53] ,
		\a[61] ,
		\a[62] ,
		_w8522_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8457 (
		\a[52] ,
		\a[53] ,
		\a[61] ,
		\a[62] ,
		_w8523_
	);
	LUT2 #(
		.INIT('h8)
	) name8458 (
		\a[54] ,
		\a[60] ,
		_w8524_
	);
	LUT4 #(
		.INIT('h153f)
	) name8459 (
		\a[55] ,
		\a[56] ,
		\a[58] ,
		\a[59] ,
		_w8525_
	);
	LUT4 #(
		.INIT('h8000)
	) name8460 (
		\a[55] ,
		\a[56] ,
		\a[58] ,
		\a[59] ,
		_w8526_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8461 (
		\a[55] ,
		\a[56] ,
		\a[58] ,
		\a[59] ,
		_w8527_
	);
	LUT4 #(
		.INIT('h0660)
	) name8462 (
		_w8520_,
		_w8523_,
		_w8524_,
		_w8527_,
		_w8528_
	);
	LUT4 #(
		.INIT('h9009)
	) name8463 (
		_w8520_,
		_w8523_,
		_w8524_,
		_w8527_,
		_w8529_
	);
	LUT4 #(
		.INIT('h6996)
	) name8464 (
		_w8520_,
		_w8523_,
		_w8524_,
		_w8527_,
		_w8530_
	);
	LUT4 #(
		.INIT('h4db2)
	) name8465 (
		_w8482_,
		_w8483_,
		_w8484_,
		_w8530_,
		_w8531_
	);
	LUT3 #(
		.INIT('he1)
	) name8466 (
		_w8518_,
		_w8519_,
		_w8531_,
		_w8532_
	);
	LUT2 #(
		.INIT('h2)
	) name8467 (
		_w8510_,
		_w8532_,
		_w8533_
	);
	LUT2 #(
		.INIT('h9)
	) name8468 (
		_w8510_,
		_w8532_,
		_w8534_
	);
	LUT4 #(
		.INIT('h7007)
	) name8469 (
		_w8476_,
		_w8497_,
		_w8510_,
		_w8532_,
		_w8535_
	);
	LUT4 #(
		.INIT('h2f00)
	) name8470 (
		_w8444_,
		_w8471_,
		_w8509_,
		_w8535_,
		_w8536_
	);
	LUT4 #(
		.INIT('h020f)
	) name8471 (
		_w8444_,
		_w8471_,
		_w8499_,
		_w8509_,
		_w8537_
	);
	LUT3 #(
		.INIT('hcd)
	) name8472 (
		_w8534_,
		_w8536_,
		_w8537_,
		_w8538_
	);
	LUT4 #(
		.INIT('h7077)
	) name8473 (
		_w8476_,
		_w8497_,
		_w8510_,
		_w8532_,
		_w8539_
	);
	LUT4 #(
		.INIT('h2f00)
	) name8474 (
		_w8444_,
		_w8471_,
		_w8509_,
		_w8539_,
		_w8540_
	);
	LUT3 #(
		.INIT('h45)
	) name8475 (
		_w8518_,
		_w8519_,
		_w8531_,
		_w8541_
	);
	LUT2 #(
		.INIT('h8)
	) name8476 (
		\a[52] ,
		\a[63] ,
		_w8542_
	);
	LUT4 #(
		.INIT('h0dff)
	) name8477 (
		_w8524_,
		_w8525_,
		_w8526_,
		_w8542_,
		_w8543_
	);
	LUT4 #(
		.INIT('h000d)
	) name8478 (
		_w8524_,
		_w8525_,
		_w8526_,
		_w8542_,
		_w8544_
	);
	LUT4 #(
		.INIT('h0df2)
	) name8479 (
		_w8524_,
		_w8525_,
		_w8526_,
		_w8542_,
		_w8545_
	);
	LUT3 #(
		.INIT('h0d)
	) name8480 (
		_w8520_,
		_w8521_,
		_w8522_,
		_w8546_
	);
	LUT2 #(
		.INIT('h6)
	) name8481 (
		_w8545_,
		_w8546_,
		_w8547_
	);
	LUT4 #(
		.INIT('h004d)
	) name8482 (
		_w8482_,
		_w8483_,
		_w8484_,
		_w8528_,
		_w8548_
	);
	LUT3 #(
		.INIT('hc8)
	) name8483 (
		_w8529_,
		_w8547_,
		_w8548_,
		_w8549_
	);
	LUT4 #(
		.INIT('h4445)
	) name8484 (
		_w8512_,
		_w8513_,
		_w8515_,
		_w8516_,
		_w8550_
	);
	LUT2 #(
		.INIT('h8)
	) name8485 (
		\a[54] ,
		\a[61] ,
		_w8551_
	);
	LUT4 #(
		.INIT('h153f)
	) name8486 (
		\a[55] ,
		\a[56] ,
		\a[59] ,
		\a[60] ,
		_w8552_
	);
	LUT4 #(
		.INIT('h8000)
	) name8487 (
		\a[55] ,
		\a[56] ,
		\a[59] ,
		\a[60] ,
		_w8553_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8488 (
		\a[55] ,
		\a[56] ,
		\a[59] ,
		\a[60] ,
		_w8554_
	);
	LUT2 #(
		.INIT('h6)
	) name8489 (
		_w8551_,
		_w8554_,
		_w8555_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8490 (
		\a[53] ,
		\a[57] ,
		\a[58] ,
		\a[62] ,
		_w8556_
	);
	LUT3 #(
		.INIT('h60)
	) name8491 (
		_w8551_,
		_w8554_,
		_w8556_,
		_w8557_
	);
	LUT3 #(
		.INIT('h09)
	) name8492 (
		_w8551_,
		_w8554_,
		_w8556_,
		_w8558_
	);
	LUT3 #(
		.INIT('h96)
	) name8493 (
		_w8551_,
		_w8554_,
		_w8556_,
		_w8559_
	);
	LUT2 #(
		.INIT('h6)
	) name8494 (
		_w8550_,
		_w8559_,
		_w8560_
	);
	LUT3 #(
		.INIT('h41)
	) name8495 (
		_w8529_,
		_w8545_,
		_w8546_,
		_w8561_
	);
	LUT2 #(
		.INIT('h4)
	) name8496 (
		_w8548_,
		_w8561_,
		_w8562_
	);
	LUT3 #(
		.INIT('hc9)
	) name8497 (
		_w8549_,
		_w8560_,
		_w8562_,
		_w8563_
	);
	LUT2 #(
		.INIT('h2)
	) name8498 (
		_w8541_,
		_w8563_,
		_w8564_
	);
	LUT2 #(
		.INIT('h9)
	) name8499 (
		_w8541_,
		_w8563_,
		_w8565_
	);
	LUT3 #(
		.INIT('he1)
	) name8500 (
		_w8533_,
		_w8540_,
		_w8565_,
		_w8566_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8501 (
		_w8510_,
		_w8532_,
		_w8541_,
		_w8563_,
		_w8567_
	);
	LUT4 #(
		.INIT('h2022)
	) name8502 (
		_w8510_,
		_w8532_,
		_w8541_,
		_w8563_,
		_w8568_
	);
	LUT2 #(
		.INIT('h4)
	) name8503 (
		_w8499_,
		_w8567_,
		_w8569_
	);
	LUT4 #(
		.INIT('h2f00)
	) name8504 (
		_w8444_,
		_w8471_,
		_w8509_,
		_w8569_,
		_w8570_
	);
	LUT3 #(
		.INIT('h0d)
	) name8505 (
		_w8551_,
		_w8552_,
		_w8553_,
		_w8571_
	);
	LUT4 #(
		.INIT('h153f)
	) name8506 (
		\a[53] ,
		\a[54] ,
		\a[62] ,
		\a[63] ,
		_w8572_
	);
	LUT2 #(
		.INIT('h8)
	) name8507 (
		\a[54] ,
		\a[63] ,
		_w8573_
	);
	LUT4 #(
		.INIT('h8000)
	) name8508 (
		\a[53] ,
		\a[54] ,
		\a[62] ,
		\a[63] ,
		_w8574_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8509 (
		\a[53] ,
		\a[54] ,
		\a[62] ,
		\a[63] ,
		_w8575_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8510 (
		\a[53] ,
		\a[57] ,
		\a[58] ,
		\a[62] ,
		_w8576_
	);
	LUT2 #(
		.INIT('h8)
	) name8511 (
		_w8575_,
		_w8576_,
		_w8577_
	);
	LUT2 #(
		.INIT('h6)
	) name8512 (
		_w8575_,
		_w8576_,
		_w8578_
	);
	LUT2 #(
		.INIT('h8)
	) name8513 (
		\a[55] ,
		\a[61] ,
		_w8579_
	);
	LUT4 #(
		.INIT('h153f)
	) name8514 (
		\a[56] ,
		\a[57] ,
		\a[59] ,
		\a[60] ,
		_w8580_
	);
	LUT4 #(
		.INIT('h8000)
	) name8515 (
		\a[56] ,
		\a[57] ,
		\a[59] ,
		\a[60] ,
		_w8581_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8516 (
		\a[56] ,
		\a[57] ,
		\a[59] ,
		\a[60] ,
		_w8582_
	);
	LUT2 #(
		.INIT('h6)
	) name8517 (
		_w8579_,
		_w8582_,
		_w8583_
	);
	LUT4 #(
		.INIT('h6996)
	) name8518 (
		_w8575_,
		_w8576_,
		_w8579_,
		_w8582_,
		_w8584_
	);
	LUT2 #(
		.INIT('h6)
	) name8519 (
		_w8571_,
		_w8584_,
		_w8585_
	);
	LUT3 #(
		.INIT('h07)
	) name8520 (
		_w8543_,
		_w8546_,
		_w8544_,
		_w8586_
	);
	LUT4 #(
		.INIT('he800)
	) name8521 (
		_w8550_,
		_w8555_,
		_w8556_,
		_w8586_,
		_w8587_
	);
	LUT4 #(
		.INIT('h00a8)
	) name8522 (
		_w8543_,
		_w8544_,
		_w8546_,
		_w8557_,
		_w8588_
	);
	LUT3 #(
		.INIT('h70)
	) name8523 (
		_w8550_,
		_w8559_,
		_w8588_,
		_w8589_
	);
	LUT4 #(
		.INIT('h31ce)
	) name8524 (
		_w8550_,
		_w8557_,
		_w8558_,
		_w8586_,
		_w8590_
	);
	LUT2 #(
		.INIT('h2)
	) name8525 (
		_w8585_,
		_w8590_,
		_w8591_
	);
	LUT4 #(
		.INIT('h080f)
	) name8526 (
		_w8550_,
		_w8559_,
		_w8585_,
		_w8588_,
		_w8592_
	);
	LUT2 #(
		.INIT('h4)
	) name8527 (
		_w8587_,
		_w8592_,
		_w8593_
	);
	LUT3 #(
		.INIT('h56)
	) name8528 (
		_w8585_,
		_w8587_,
		_w8589_,
		_w8594_
	);
	LUT4 #(
		.INIT('h82c3)
	) name8529 (
		_w8548_,
		_w8550_,
		_w8559_,
		_w8561_,
		_w8595_
	);
	LUT2 #(
		.INIT('h1)
	) name8530 (
		_w8549_,
		_w8595_,
		_w8596_
	);
	LUT4 #(
		.INIT('h0045)
	) name8531 (
		_w8549_,
		_w8587_,
		_w8592_,
		_w8595_,
		_w8597_
	);
	LUT2 #(
		.INIT('h4)
	) name8532 (
		_w8591_,
		_w8597_,
		_w8598_
	);
	LUT3 #(
		.INIT('he1)
	) name8533 (
		_w8591_,
		_w8593_,
		_w8596_,
		_w8599_
	);
	LUT4 #(
		.INIT('hfe01)
	) name8534 (
		_w8564_,
		_w8568_,
		_w8570_,
		_w8599_,
		_w8600_
	);
	LUT4 #(
		.INIT('hddd0)
	) name8535 (
		_w8541_,
		_w8563_,
		_w8594_,
		_w8596_,
		_w8601_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8536 (
		\a[55] ,
		\a[58] ,
		\a[59] ,
		\a[62] ,
		_w8602_
	);
	LUT4 #(
		.INIT('hf200)
	) name8537 (
		_w8551_,
		_w8552_,
		_w8553_,
		_w8602_,
		_w8603_
	);
	LUT4 #(
		.INIT('h117f)
	) name8538 (
		_w8578_,
		_w8583_,
		_w8602_,
		_w8603_,
		_w8604_
	);
	LUT4 #(
		.INIT('hffd4)
	) name8539 (
		_w8571_,
		_w8578_,
		_w8583_,
		_w8602_,
		_w8605_
	);
	LUT2 #(
		.INIT('h8)
	) name8540 (
		_w8604_,
		_w8605_,
		_w8606_
	);
	LUT3 #(
		.INIT('h23)
	) name8541 (
		_w8572_,
		_w8574_,
		_w8576_,
		_w8607_
	);
	LUT3 #(
		.INIT('h0d)
	) name8542 (
		_w8579_,
		_w8580_,
		_w8581_,
		_w8608_
	);
	LUT2 #(
		.INIT('h1)
	) name8543 (
		_w8607_,
		_w8608_,
		_w8609_
	);
	LUT4 #(
		.INIT('h153f)
	) name8544 (
		\a[56] ,
		\a[57] ,
		\a[60] ,
		\a[61] ,
		_w8610_
	);
	LUT4 #(
		.INIT('h8000)
	) name8545 (
		\a[56] ,
		\a[57] ,
		\a[60] ,
		\a[61] ,
		_w8611_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8546 (
		\a[56] ,
		\a[57] ,
		\a[60] ,
		\a[61] ,
		_w8612_
	);
	LUT2 #(
		.INIT('h6)
	) name8547 (
		_w8573_,
		_w8612_,
		_w8613_
	);
	LUT4 #(
		.INIT('h0051)
	) name8548 (
		_w8574_,
		_w8579_,
		_w8580_,
		_w8581_,
		_w8614_
	);
	LUT2 #(
		.INIT('h4)
	) name8549 (
		_w8577_,
		_w8614_,
		_w8615_
	);
	LUT3 #(
		.INIT('h36)
	) name8550 (
		_w8609_,
		_w8613_,
		_w8615_,
		_w8616_
	);
	LUT4 #(
		.INIT('he00e)
	) name8551 (
		_w8587_,
		_w8592_,
		_w8606_,
		_w8616_,
		_w8617_
	);
	LUT4 #(
		.INIT('h0110)
	) name8552 (
		_w8587_,
		_w8592_,
		_w8606_,
		_w8616_,
		_w8618_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name8553 (
		_w8587_,
		_w8592_,
		_w8606_,
		_w8616_,
		_w8619_
	);
	LUT3 #(
		.INIT('hb0)
	) name8554 (
		_w8591_,
		_w8597_,
		_w8619_,
		_w8620_
	);
	LUT4 #(
		.INIT('hef00)
	) name8555 (
		_w8568_,
		_w8570_,
		_w8601_,
		_w8620_,
		_w8621_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name8556 (
		_w8568_,
		_w8570_,
		_w8598_,
		_w8601_,
		_w8622_
	);
	LUT3 #(
		.INIT('hcd)
	) name8557 (
		_w8619_,
		_w8621_,
		_w8622_,
		_w8623_
	);
	LUT3 #(
		.INIT('h0b)
	) name8558 (
		_w8591_,
		_w8597_,
		_w8617_,
		_w8624_
	);
	LUT4 #(
		.INIT('hef00)
	) name8559 (
		_w8568_,
		_w8570_,
		_w8601_,
		_w8624_,
		_w8625_
	);
	LUT3 #(
		.INIT('h13)
	) name8560 (
		\a[55] ,
		\a[58] ,
		\a[62] ,
		_w8626_
	);
	LUT2 #(
		.INIT('h8)
	) name8561 (
		\a[55] ,
		\a[63] ,
		_w8627_
	);
	LUT3 #(
		.INIT('h80)
	) name8562 (
		\a[55] ,
		\a[59] ,
		\a[63] ,
		_w8628_
	);
	LUT2 #(
		.INIT('h4)
	) name8563 (
		_w8626_,
		_w8628_,
		_w8629_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8564 (
		\a[55] ,
		\a[58] ,
		\a[59] ,
		\a[62] ,
		_w8630_
	);
	LUT2 #(
		.INIT('h1)
	) name8565 (
		_w8627_,
		_w8630_,
		_w8631_
	);
	LUT3 #(
		.INIT('hd2)
	) name8566 (
		\a[59] ,
		_w8626_,
		_w8627_,
		_w8632_
	);
	LUT3 #(
		.INIT('h0d)
	) name8567 (
		_w8573_,
		_w8610_,
		_w8611_,
		_w8633_
	);
	LUT2 #(
		.INIT('h6)
	) name8568 (
		_w8632_,
		_w8633_,
		_w8634_
	);
	LUT3 #(
		.INIT('h0e)
	) name8569 (
		_w8607_,
		_w8608_,
		_w8613_,
		_w8635_
	);
	LUT2 #(
		.INIT('h8)
	) name8570 (
		\a[56] ,
		\a[62] ,
		_w8636_
	);
	LUT4 #(
		.INIT('h153f)
	) name8571 (
		\a[57] ,
		\a[58] ,
		\a[60] ,
		\a[61] ,
		_w8637_
	);
	LUT4 #(
		.INIT('h8000)
	) name8572 (
		\a[57] ,
		\a[58] ,
		\a[60] ,
		\a[61] ,
		_w8638_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8573 (
		\a[57] ,
		\a[58] ,
		\a[60] ,
		\a[61] ,
		_w8639_
	);
	LUT2 #(
		.INIT('h6)
	) name8574 (
		_w8636_,
		_w8639_,
		_w8640_
	);
	LUT3 #(
		.INIT('hb0)
	) name8575 (
		_w8577_,
		_w8614_,
		_w8640_,
		_w8641_
	);
	LUT4 #(
		.INIT('hf10e)
	) name8576 (
		_w8609_,
		_w8613_,
		_w8615_,
		_w8640_,
		_w8642_
	);
	LUT2 #(
		.INIT('h9)
	) name8577 (
		_w8634_,
		_w8642_,
		_w8643_
	);
	LUT3 #(
		.INIT('ha2)
	) name8578 (
		_w8604_,
		_w8605_,
		_w8616_,
		_w8644_
	);
	LUT2 #(
		.INIT('h4)
	) name8579 (
		_w8643_,
		_w8644_,
		_w8645_
	);
	LUT3 #(
		.INIT('h96)
	) name8580 (
		_w8618_,
		_w8643_,
		_w8644_,
		_w8646_
	);
	LUT3 #(
		.INIT('hc3)
	) name8581 (
		_w8618_,
		_w8643_,
		_w8644_,
		_w8647_
	);
	LUT3 #(
		.INIT('he4)
	) name8582 (
		_w8625_,
		_w8646_,
		_w8647_,
		_w8648_
	);
	LUT3 #(
		.INIT('h51)
	) name8583 (
		_w8617_,
		_w8643_,
		_w8644_,
		_w8649_
	);
	LUT2 #(
		.INIT('h4)
	) name8584 (
		_w8598_,
		_w8649_,
		_w8650_
	);
	LUT4 #(
		.INIT('hef00)
	) name8585 (
		_w8568_,
		_w8570_,
		_w8601_,
		_w8650_,
		_w8651_
	);
	LUT3 #(
		.INIT('ha2)
	) name8586 (
		_w8618_,
		_w8643_,
		_w8644_,
		_w8652_
	);
	LUT3 #(
		.INIT('h23)
	) name8587 (
		_w8629_,
		_w8631_,
		_w8633_,
		_w8653_
	);
	LUT3 #(
		.INIT('h0d)
	) name8588 (
		_w8636_,
		_w8637_,
		_w8638_,
		_w8654_
	);
	LUT2 #(
		.INIT('h8)
	) name8589 (
		\a[58] ,
		\a[63] ,
		_w8655_
	);
	LUT4 #(
		.INIT('h8000)
	) name8590 (
		\a[56] ,
		\a[58] ,
		\a[61] ,
		\a[63] ,
		_w8656_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8591 (
		\a[56] ,
		\a[58] ,
		\a[61] ,
		\a[63] ,
		_w8657_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8592 (
		\a[57] ,
		\a[59] ,
		\a[60] ,
		\a[62] ,
		_w8658_
	);
	LUT3 #(
		.INIT('h6f)
	) name8593 (
		_w8654_,
		_w8657_,
		_w8658_,
		_w8659_
	);
	LUT3 #(
		.INIT('hf9)
	) name8594 (
		_w8654_,
		_w8657_,
		_w8658_,
		_w8660_
	);
	LUT3 #(
		.INIT('h69)
	) name8595 (
		_w8654_,
		_w8657_,
		_w8658_,
		_w8661_
	);
	LUT2 #(
		.INIT('h6)
	) name8596 (
		_w8653_,
		_w8661_,
		_w8662_
	);
	LUT3 #(
		.INIT('h8a)
	) name8597 (
		_w8634_,
		_w8635_,
		_w8641_,
		_w8663_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8598 (
		_w8609_,
		_w8613_,
		_w8615_,
		_w8640_,
		_w8664_
	);
	LUT3 #(
		.INIT('h02)
	) name8599 (
		_w8662_,
		_w8663_,
		_w8664_,
		_w8665_
	);
	LUT3 #(
		.INIT('h54)
	) name8600 (
		_w8662_,
		_w8663_,
		_w8664_,
		_w8666_
	);
	LUT3 #(
		.INIT('ha9)
	) name8601 (
		_w8662_,
		_w8663_,
		_w8664_,
		_w8667_
	);
	LUT4 #(
		.INIT('hfe01)
	) name8602 (
		_w8645_,
		_w8651_,
		_w8652_,
		_w8667_,
		_w8668_
	);
	LUT4 #(
		.INIT('h004d)
	) name8603 (
		_w8618_,
		_w8643_,
		_w8644_,
		_w8666_,
		_w8669_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8604 (
		\a[57] ,
		\a[59] ,
		\a[60] ,
		\a[62] ,
		_w8670_
	);
	LUT4 #(
		.INIT('h153f)
	) name8605 (
		\a[56] ,
		\a[58] ,
		\a[61] ,
		\a[63] ,
		_w8671_
	);
	LUT4 #(
		.INIT('h000d)
	) name8606 (
		_w8636_,
		_w8637_,
		_w8638_,
		_w8656_,
		_w8672_
	);
	LUT2 #(
		.INIT('h8)
	) name8607 (
		\a[57] ,
		\a[63] ,
		_w8673_
	);
	LUT4 #(
		.INIT('h153f)
	) name8608 (
		\a[58] ,
		\a[59] ,
		\a[61] ,
		\a[62] ,
		_w8674_
	);
	LUT4 #(
		.INIT('h8000)
	) name8609 (
		\a[58] ,
		\a[59] ,
		\a[61] ,
		\a[62] ,
		_w8675_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8610 (
		\a[58] ,
		\a[59] ,
		\a[61] ,
		\a[62] ,
		_w8676_
	);
	LUT2 #(
		.INIT('h6)
	) name8611 (
		_w8673_,
		_w8676_,
		_w8677_
	);
	LUT4 #(
		.INIT('h56a9)
	) name8612 (
		_w8670_,
		_w8671_,
		_w8672_,
		_w8677_,
		_w8678_
	);
	LUT4 #(
		.INIT('h004f)
	) name8613 (
		_w8653_,
		_w8659_,
		_w8660_,
		_w8678_,
		_w8679_
	);
	LUT4 #(
		.INIT('hb000)
	) name8614 (
		_w8653_,
		_w8659_,
		_w8660_,
		_w8678_,
		_w8680_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name8615 (
		_w8653_,
		_w8659_,
		_w8660_,
		_w8678_,
		_w8681_
	);
	LUT4 #(
		.INIT('h23dc)
	) name8616 (
		_w8651_,
		_w8665_,
		_w8669_,
		_w8681_,
		_w8682_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8617 (
		_w8662_,
		_w8663_,
		_w8664_,
		_w8680_,
		_w8683_
	);
	LUT4 #(
		.INIT('h33f7)
	) name8618 (
		\a[57] ,
		_w8655_,
		_w8674_,
		_w8675_,
		_w8684_
	);
	LUT4 #(
		.INIT('h0051)
	) name8619 (
		_w8655_,
		_w8673_,
		_w8674_,
		_w8675_,
		_w8685_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8620 (
		\a[59] ,
		\a[60] ,
		\a[61] ,
		\a[62] ,
		_w8686_
	);
	LUT3 #(
		.INIT('h2d)
	) name8621 (
		_w8684_,
		_w8685_,
		_w8686_,
		_w8687_
	);
	LUT4 #(
		.INIT('hab02)
	) name8622 (
		_w8670_,
		_w8671_,
		_w8672_,
		_w8677_,
		_w8688_
	);
	LUT2 #(
		.INIT('h2)
	) name8623 (
		_w8687_,
		_w8688_,
		_w8689_
	);
	LUT2 #(
		.INIT('h4)
	) name8624 (
		_w8687_,
		_w8688_,
		_w8690_
	);
	LUT2 #(
		.INIT('h9)
	) name8625 (
		_w8687_,
		_w8688_,
		_w8691_
	);
	LUT2 #(
		.INIT('h9)
	) name8626 (
		_w8679_,
		_w8691_,
		_w8692_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8627 (
		_w8651_,
		_w8669_,
		_w8683_,
		_w8692_,
		_w8693_
	);
	LUT2 #(
		.INIT('hc)
	) name8628 (
		_w8679_,
		_w8691_,
		_w8694_
	);
	LUT4 #(
		.INIT('hb000)
	) name8629 (
		_w8651_,
		_w8669_,
		_w8683_,
		_w8694_,
		_w8695_
	);
	LUT2 #(
		.INIT('he)
	) name8630 (
		_w8693_,
		_w8695_,
		_w8696_
	);
	LUT2 #(
		.INIT('h1)
	) name8631 (
		_w8680_,
		_w8690_,
		_w8697_
	);
	LUT2 #(
		.INIT('h4)
	) name8632 (
		_w8665_,
		_w8697_,
		_w8698_
	);
	LUT4 #(
		.INIT('h153f)
	) name8633 (
		\a[59] ,
		\a[60] ,
		\a[62] ,
		\a[63] ,
		_w8699_
	);
	LUT4 #(
		.INIT('h8000)
	) name8634 (
		\a[59] ,
		\a[60] ,
		\a[62] ,
		\a[63] ,
		_w8700_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name8635 (
		\a[59] ,
		\a[60] ,
		\a[62] ,
		\a[63] ,
		_w8701_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8636 (
		\a[59] ,
		\a[60] ,
		\a[61] ,
		\a[62] ,
		_w8702_
	);
	LUT2 #(
		.INIT('h6)
	) name8637 (
		_w8701_,
		_w8702_,
		_w8703_
	);
	LUT4 #(
		.INIT('h00ce)
	) name8638 (
		_w8684_,
		_w8685_,
		_w8686_,
		_w8703_,
		_w8704_
	);
	LUT4 #(
		.INIT('h3100)
	) name8639 (
		_w8684_,
		_w8685_,
		_w8686_,
		_w8703_,
		_w8705_
	);
	LUT4 #(
		.INIT('hce31)
	) name8640 (
		_w8684_,
		_w8685_,
		_w8686_,
		_w8703_,
		_w8706_
	);
	LUT3 #(
		.INIT('hd0)
	) name8641 (
		_w8687_,
		_w8688_,
		_w8706_,
		_w8707_
	);
	LUT3 #(
		.INIT('hd0)
	) name8642 (
		_w8679_,
		_w8690_,
		_w8707_,
		_w8708_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8643 (
		_w8651_,
		_w8669_,
		_w8698_,
		_w8708_,
		_w8709_
	);
	LUT3 #(
		.INIT('h31)
	) name8644 (
		_w8679_,
		_w8689_,
		_w8690_,
		_w8710_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8645 (
		_w8651_,
		_w8669_,
		_w8698_,
		_w8710_,
		_w8711_
	);
	LUT3 #(
		.INIT('h32)
	) name8646 (
		_w8706_,
		_w8709_,
		_w8711_,
		_w8712_
	);
	LUT3 #(
		.INIT('h0d)
	) name8647 (
		_w8687_,
		_w8688_,
		_w8704_,
		_w8713_
	);
	LUT3 #(
		.INIT('hd0)
	) name8648 (
		_w8679_,
		_w8690_,
		_w8713_,
		_w8714_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8649 (
		_w8651_,
		_w8669_,
		_w8698_,
		_w8714_,
		_w8715_
	);
	LUT4 #(
		.INIT('h9a30)
	) name8650 (
		\a[60] ,
		\a[61] ,
		\a[62] ,
		\a[63] ,
		_w8716_
	);
	LUT4 #(
		.INIT('h0023)
	) name8651 (
		_w8699_,
		_w8700_,
		_w8702_,
		_w8716_,
		_w8717_
	);
	LUT4 #(
		.INIT('hea00)
	) name8652 (
		_w8700_,
		_w8701_,
		_w8702_,
		_w8716_,
		_w8718_
	);
	LUT4 #(
		.INIT('h15ea)
	) name8653 (
		_w8700_,
		_w8701_,
		_w8702_,
		_w8716_,
		_w8719_
	);
	LUT3 #(
		.INIT('h1e)
	) name8654 (
		_w8705_,
		_w8715_,
		_w8719_,
		_w8720_
	);
	LUT4 #(
		.INIT('h2cc0)
	) name8655 (
		\a[60] ,
		\a[61] ,
		\a[62] ,
		\a[63] ,
		_w8721_
	);
	LUT2 #(
		.INIT('h8)
	) name8656 (
		_w8717_,
		_w8721_,
		_w8722_
	);
	LUT2 #(
		.INIT('h4)
	) name8657 (
		_w8718_,
		_w8721_,
		_w8723_
	);
	LUT2 #(
		.INIT('h4)
	) name8658 (
		_w8705_,
		_w8723_,
		_w8724_
	);
	LUT3 #(
		.INIT('h23)
	) name8659 (
		_w8715_,
		_w8722_,
		_w8724_,
		_w8725_
	);
	LUT2 #(
		.INIT('h1)
	) name8660 (
		_w8705_,
		_w8718_,
		_w8726_
	);
	LUT2 #(
		.INIT('h1)
	) name8661 (
		_w8717_,
		_w8721_,
		_w8727_
	);
	LUT3 #(
		.INIT('hb0)
	) name8662 (
		_w8715_,
		_w8726_,
		_w8727_,
		_w8728_
	);
	LUT2 #(
		.INIT('hd)
	) name8663 (
		_w8725_,
		_w8728_,
		_w8729_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8664 (
		\a[60] ,
		\a[61] ,
		\a[62] ,
		\a[63] ,
		_w8730_
	);
	LUT2 #(
		.INIT('h4)
	) name8665 (
		_w8717_,
		_w8730_,
		_w8731_
	);
	LUT3 #(
		.INIT('hb0)
	) name8666 (
		_w8715_,
		_w8726_,
		_w8731_,
		_w8732_
	);
	LUT4 #(
		.INIT('hecc0)
	) name8667 (
		\a[60] ,
		\a[61] ,
		\a[62] ,
		\a[63] ,
		_w8733_
	);
	LUT2 #(
		.INIT('h4)
	) name8668 (
		_w8717_,
		_w8733_,
		_w8734_
	);
	LUT3 #(
		.INIT('hb0)
	) name8669 (
		\a[61] ,
		\a[62] ,
		\a[63] ,
		_w8735_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8670 (
		_w8715_,
		_w8726_,
		_w8734_,
		_w8735_,
		_w8736_
	);
	LUT2 #(
		.INIT('he)
	) name8671 (
		_w8732_,
		_w8736_,
		_w8737_
	);
	LUT4 #(
		.INIT('h1055)
	) name8672 (
		\a[62] ,
		_w8715_,
		_w8726_,
		_w8734_,
		_w8738_
	);
	LUT2 #(
		.INIT('h2)
	) name8673 (
		\a[63] ,
		_w8738_,
		_w8739_
	);
	assign \asquared[0]  = \a[0] ;
	assign \asquared[1]  = 1'b0;
	assign \asquared[2]  = _w66_ ;
	assign \asquared[3]  = _w68_ ;
	assign \asquared[4]  = _w70_ ;
	assign \asquared[5]  = _w73_ ;
	assign \asquared[6]  = _w83_ ;
	assign \asquared[7]  = _w98_ ;
	assign \asquared[8]  = _w112_ ;
	assign \asquared[9]  = _w131_ ;
	assign \asquared[10]  = _w145_ ;
	assign \asquared[11]  = _w170_ ;
	assign \asquared[12]  = _w197_ ;
	assign \asquared[13]  = _w219_ ;
	assign \asquared[14]  = _w249_ ;
	assign \asquared[15]  = _w278_ ;
	assign \asquared[16]  = _w309_ ;
	assign \asquared[17]  = _w345_ ;
	assign \asquared[18]  = _w389_ ;
	assign \asquared[19]  = _w418_ ;
	assign \asquared[20]  = _w461_ ;
	assign \asquared[21]  = _w506_ ;
	assign \asquared[22]  = _w552_ ;
	assign \asquared[23]  = _w608_ ;
	assign \asquared[24]  = _w661_ ;
	assign \asquared[25]  = _w712_ ;
	assign \asquared[26]  = _w763_ ;
	assign \asquared[27]  = _w820_ ;
	assign \asquared[28]  = _w876_ ;
	assign \asquared[29]  = _w943_ ;
	assign \asquared[30]  = _w1003_ ;
	assign \asquared[31]  = _w1059_ ;
	assign \asquared[32]  = _w1133_ ;
	assign \asquared[33]  = _w1209_ ;
	assign \asquared[34]  = _w1273_ ;
	assign \asquared[35]  = _w1343_ ;
	assign \asquared[36]  = _w1417_ ;
	assign \asquared[37]  = _w1494_ ;
	assign \asquared[38]  = _w1576_ ;
	assign \asquared[39]  = _w1660_ ;
	assign \asquared[40]  = _w1741_ ;
	assign \asquared[41]  = _w1825_ ;
	assign \asquared[42]  = _w1914_ ;
	assign \asquared[43]  = _w2000_ ;
	assign \asquared[44]  = _w2088_ ;
	assign \asquared[45]  = _w2190_ ;
	assign \asquared[46]  = _w2293_ ;
	assign \asquared[47]  = _w2400_ ;
	assign \asquared[48]  = _w2495_ ;
	assign \asquared[49]  = _w2586_ ;
	assign \asquared[50]  = _w2692_ ;
	assign \asquared[51]  = _w2797_ ;
	assign \asquared[52]  = _w2900_ ;
	assign \asquared[53]  = _w3000_ ;
	assign \asquared[54]  = _w3112_ ;
	assign \asquared[55]  = _w3220_ ;
	assign \asquared[56]  = _w3350_ ;
	assign \asquared[57]  = _w3466_ ;
	assign \asquared[58]  = _w3584_ ;
	assign \asquared[59]  = _w3701_ ;
	assign \asquared[60]  = _w3828_ ;
	assign \asquared[61]  = _w3946_ ;
	assign \asquared[62]  = _w4076_ ;
	assign \asquared[63]  = _w4219_ ;
	assign \asquared[64]  = _w4344_ ;
	assign \asquared[65]  = _w4477_ ;
	assign \asquared[66]  = _w4602_ ;
	assign \asquared[67]  = _w4737_ ;
	assign \asquared[68]  = _w4864_ ;
	assign \asquared[69]  = _w4991_ ;
	assign \asquared[70]  = _w5102_ ;
	assign \asquared[71]  = _w5220_ ;
	assign \asquared[72]  = _w5343_ ;
	assign \asquared[73]  = _w5464_ ;
	assign \asquared[74]  = _w5579_ ;
	assign \asquared[75]  = _w5692_ ;
	assign \asquared[76]  = _w5801_ ;
	assign \asquared[77]  = _w5928_ ;
	assign \asquared[78]  = _w6036_ ;
	assign \asquared[79]  = _w6144_ ;
	assign \asquared[80]  = _w6260_ ;
	assign \asquared[81]  = _w6352_ ;
	assign \asquared[82]  = _w6450_ ;
	assign \asquared[83]  = _w6547_ ;
	assign \asquared[84]  = _w6631_ ;
	assign \asquared[85]  = _w6731_ ;
	assign \asquared[86]  = _w6817_ ;
	assign \asquared[87]  = _w6906_ ;
	assign \asquared[88]  = _w6989_ ;
	assign \asquared[89]  = _w7071_ ;
	assign \asquared[90]  = _w7146_ ;
	assign \asquared[91]  = _w7230_ ;
	assign \asquared[92]  = _w7305_ ;
	assign \asquared[93]  = _w7380_ ;
	assign \asquared[94]  = _w7449_ ;
	assign \asquared[95]  = _w7528_ ;
	assign \asquared[96]  = _w7600_ ;
	assign \asquared[97]  = _w7678_ ;
	assign \asquared[98]  = _w7734_ ;
	assign \asquared[99]  = _w7797_ ;
	assign \asquared[100]  = _w7859_ ;
	assign \asquared[101]  = _w7920_ ;
	assign \asquared[102]  = _w7983_ ;
	assign \asquared[103]  = _w8042_ ;
	assign \asquared[104]  = _w8088_ ;
	assign \asquared[105]  = _w8139_ ;
	assign \asquared[106]  = _w8185_ ;
	assign \asquared[107]  = _w8237_ ;
	assign \asquared[108]  = _w8277_ ;
	assign \asquared[109]  = _w8325_ ;
	assign \asquared[110]  = _w8372_ ;
	assign \asquared[111]  = _w8408_ ;
	assign \asquared[112]  = _w8442_ ;
	assign \asquared[113]  = _w8475_ ;
	assign \asquared[114]  = _w8507_ ;
	assign \asquared[115]  = _w8538_ ;
	assign \asquared[116]  = _w8566_ ;
	assign \asquared[117]  = _w8600_ ;
	assign \asquared[118]  = _w8623_ ;
	assign \asquared[119]  = _w8648_ ;
	assign \asquared[120]  = _w8668_ ;
	assign \asquared[121]  = _w8682_ ;
	assign \asquared[122]  = _w8696_ ;
	assign \asquared[123]  = _w8712_ ;
	assign \asquared[124]  = _w8720_ ;
	assign \asquared[125]  = _w8729_ ;
	assign \asquared[126]  = _w8737_ ;
	assign \asquared[127]  = _w8739_ ;
endmodule;