module top( \G0_pad  , \G10_reg/NET0131  , \G11_reg/NET0131  , \G12_reg/NET0131  , \G13_reg/NET0131  , \G147_pad  , \G148_pad  , \G14_reg/NET0131  , \G15_reg/NET0131  , \G16_reg/NET0131  , \G17_reg/NET0131  , \G18_reg/NET0131  , \G198_pad  , \G199_pad  , \G19_reg/NET0131  , \G1_pad  , \G20_reg/NET0131  , \G213_pad  , \G214_pad  , \G21_reg/NET0131  , \G22_reg/NET0131  , \G29_reg/NET0131  , \G2_pad  , \G30_reg/NET0131  , \_al_n0  , \_al_n1  , \g1001/_0_  , \g1006/_0_  , \g1008/_0_  , \g1012/_0_  , \g1020/_0_  , \g1036/_0_  , \g1056/_0_  , \g1068/_0_  , \g1070/_0_  , \g1152/_0_  , \g1298/_0_  , \g1331/_2_  , \g971/_2_  , \g973/_2_  , \g975/_2_  , \g983/_0_  , \g984/_0_  , \g985/_0_  , \g991/_2_  , \g993/_0_  , \g997/_0_  );
  input \G0_pad  ;
  input \G10_reg/NET0131  ;
  input \G11_reg/NET0131  ;
  input \G12_reg/NET0131  ;
  input \G13_reg/NET0131  ;
  input \G147_pad  ;
  input \G148_pad  ;
  input \G14_reg/NET0131  ;
  input \G15_reg/NET0131  ;
  input \G16_reg/NET0131  ;
  input \G17_reg/NET0131  ;
  input \G18_reg/NET0131  ;
  input \G198_pad  ;
  input \G199_pad  ;
  input \G19_reg/NET0131  ;
  input \G1_pad  ;
  input \G20_reg/NET0131  ;
  input \G213_pad  ;
  input \G214_pad  ;
  input \G21_reg/NET0131  ;
  input \G22_reg/NET0131  ;
  input \G29_reg/NET0131  ;
  input \G2_pad  ;
  input \G30_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1001/_0_  ;
  output \g1006/_0_  ;
  output \g1008/_0_  ;
  output \g1012/_0_  ;
  output \g1020/_0_  ;
  output \g1036/_0_  ;
  output \g1056/_0_  ;
  output \g1068/_0_  ;
  output \g1070/_0_  ;
  output \g1152/_0_  ;
  output \g1298/_0_  ;
  output \g1331/_2_  ;
  output \g971/_2_  ;
  output \g973/_2_  ;
  output \g975/_2_  ;
  output \g983/_0_  ;
  output \g984/_0_  ;
  output \g985/_0_  ;
  output \g991/_2_  ;
  output \g993/_0_  ;
  output \g997/_0_  ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 ;
  assign n25 = ~\G14_reg/NET0131  & \G15_reg/NET0131  ;
  assign n26 = \G10_reg/NET0131  & ~\G11_reg/NET0131  ;
  assign n27 = n25 & n26 ;
  assign n28 = ~\G30_reg/NET0131  & ~n27 ;
  assign n29 = \G16_reg/NET0131  & ~n28 ;
  assign n30 = \G17_reg/NET0131  & n29 ;
  assign n32 = \G18_reg/NET0131  & n30 ;
  assign n31 = ~\G18_reg/NET0131  & ~n30 ;
  assign n33 = ~\G0_pad  & ~n31 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = ~\G17_reg/NET0131  & ~\G18_reg/NET0131  ;
  assign n36 = \G16_reg/NET0131  & \G19_reg/NET0131  ;
  assign n37 = n35 & n36 ;
  assign n38 = ~n28 & n37 ;
  assign n39 = ~\G20_reg/NET0131  & ~n38 ;
  assign n40 = \G20_reg/NET0131  & n38 ;
  assign n41 = ~\G0_pad  & ~n40 ;
  assign n42 = ~n39 & n41 ;
  assign n44 = \G12_reg/NET0131  & ~\G13_reg/NET0131  ;
  assign n43 = \G20_reg/NET0131  & ~\G21_reg/NET0131  ;
  assign n45 = ~\G29_reg/NET0131  & n43 ;
  assign n46 = n44 & n45 ;
  assign n47 = \G22_reg/NET0131  & ~n46 ;
  assign n48 = ~\G20_reg/NET0131  & ~\G21_reg/NET0131  ;
  assign n49 = \G29_reg/NET0131  & n48 ;
  assign n50 = n44 & n49 ;
  assign n51 = ~n47 & ~n50 ;
  assign n52 = ~\G0_pad  & ~n51 ;
  assign n53 = ~\G16_reg/NET0131  & n28 ;
  assign n54 = ~\G0_pad  & ~n29 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = \G10_reg/NET0131  & \G11_reg/NET0131  ;
  assign n58 = ~\G14_reg/NET0131  & ~n56 ;
  assign n57 = \G14_reg/NET0131  & n56 ;
  assign n59 = ~\G0_pad  & ~n57 ;
  assign n60 = ~n58 & n59 ;
  assign n63 = \G15_reg/NET0131  & n57 ;
  assign n62 = ~\G15_reg/NET0131  & ~n57 ;
  assign n61 = ~\G14_reg/NET0131  & n26 ;
  assign n64 = ~\G0_pad  & ~n61 ;
  assign n65 = ~n62 & n64 ;
  assign n66 = ~n63 & n65 ;
  assign n67 = \G10_reg/NET0131  & ~n25 ;
  assign n68 = ~\G11_reg/NET0131  & ~n67 ;
  assign n69 = ~\G0_pad  & ~n56 ;
  assign n70 = ~n68 & n69 ;
  assign n71 = \G1_pad  & ~\G30_reg/NET0131  ;
  assign n72 = ~\G1_pad  & \G30_reg/NET0131  ;
  assign n73 = ~n71 & ~n72 ;
  assign n74 = ~\G0_pad  & ~n73 ;
  assign n75 = \G29_reg/NET0131  & ~\G2_pad  ;
  assign n76 = ~\G29_reg/NET0131  & \G2_pad  ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = ~\G0_pad  & ~n77 ;
  assign n79 = ~\G0_pad  & ~\G10_reg/NET0131  ;
  assign n80 = \G12_reg/NET0131  & \G21_reg/NET0131  ;
  assign n81 = ~\G12_reg/NET0131  & ~\G21_reg/NET0131  ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = n40 & ~n82 ;
  assign n84 = ~\G0_pad  & \G13_reg/NET0131  ;
  assign n85 = ~n83 & n84 ;
  assign n86 = ~\G0_pad  & \G12_reg/NET0131  ;
  assign n87 = ~\G13_reg/NET0131  & \G20_reg/NET0131  ;
  assign n88 = \G21_reg/NET0131  & n87 ;
  assign n89 = n86 & n88 ;
  assign n90 = n38 & n89 ;
  assign n91 = ~n85 & ~n90 ;
  assign n92 = ~\G18_reg/NET0131  & ~n51 ;
  assign n95 = \G13_reg/NET0131  & ~\G20_reg/NET0131  ;
  assign n96 = ~\G21_reg/NET0131  & n95 ;
  assign n93 = \G13_reg/NET0131  & \G21_reg/NET0131  ;
  assign n94 = \G199_pad  & n93 ;
  assign n97 = ~\G12_reg/NET0131  & ~n94 ;
  assign n98 = ~n96 & n97 ;
  assign n99 = n51 & ~n98 ;
  assign n100 = ~n92 & ~n99 ;
  assign n101 = \G13_reg/NET0131  & ~\G22_reg/NET0131  ;
  assign n102 = \G12_reg/NET0131  & ~\G199_pad  ;
  assign n103 = n101 & n102 ;
  assign n104 = ~n100 & ~n103 ;
  assign n107 = n81 & n95 ;
  assign n108 = ~n44 & ~n107 ;
  assign n105 = ~\G12_reg/NET0131  & ~n93 ;
  assign n106 = ~\G148_pad  & ~n105 ;
  assign n109 = ~n88 & ~n106 ;
  assign n110 = n108 & n109 ;
  assign n111 = n51 & n110 ;
  assign n112 = ~\G198_pad  & ~n105 ;
  assign n113 = n108 & ~n112 ;
  assign n114 = n51 & n113 ;
  assign n115 = \G13_reg/NET0131  & \G214_pad  ;
  assign n116 = ~n87 & ~n115 ;
  assign n117 = ~n44 & ~n81 ;
  assign n118 = ~n116 & n117 ;
  assign n119 = n51 & n118 ;
  assign n120 = \G21_reg/NET0131  & n41 ;
  assign n121 = ~\G12_reg/NET0131  & \G13_reg/NET0131  ;
  assign n122 = ~\G0_pad  & n43 ;
  assign n123 = ~n121 & n122 ;
  assign n124 = n38 & n123 ;
  assign n125 = ~n120 & ~n124 ;
  assign n127 = ~\G12_reg/NET0131  & n43 ;
  assign n126 = ~\G213_pad  & ~n81 ;
  assign n128 = n101 & ~n126 ;
  assign n129 = ~n127 & n128 ;
  assign n130 = ~n92 & ~n129 ;
  assign n131 = \G21_reg/NET0131  & n40 ;
  assign n132 = n86 & ~n131 ;
  assign n133 = ~\G0_pad  & ~\G12_reg/NET0131  ;
  assign n134 = n131 & n133 ;
  assign n135 = ~n132 & ~n134 ;
  assign n136 = ~\G19_reg/NET0131  & ~n32 ;
  assign n137 = \G17_reg/NET0131  & \G18_reg/NET0131  ;
  assign n138 = \G19_reg/NET0131  & n137 ;
  assign n139 = ~n35 & ~n138 ;
  assign n140 = n29 & ~n139 ;
  assign n141 = ~\G0_pad  & ~n140 ;
  assign n142 = ~n136 & n141 ;
  assign n143 = \G13_reg/NET0131  & ~\G147_pad  ;
  assign n144 = ~n105 & ~n143 ;
  assign n145 = n51 & n144 ;
  assign n146 = ~\G18_reg/NET0131  & \G19_reg/NET0131  ;
  assign n147 = n29 & ~n146 ;
  assign n148 = ~\G17_reg/NET0131  & ~n147 ;
  assign n149 = ~\G0_pad  & ~n30 ;
  assign n150 = ~n148 & n149 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1001/_0_  = n34 ;
  assign \g1006/_0_  = n42 ;
  assign \g1008/_0_  = n52 ;
  assign \g1012/_0_  = n55 ;
  assign \g1020/_0_  = n60 ;
  assign \g1036/_0_  = n66 ;
  assign \g1056/_0_  = n70 ;
  assign \g1068/_0_  = n74 ;
  assign \g1070/_0_  = n78 ;
  assign \g1152/_0_  = n79 ;
  assign \g1298/_0_  = ~n91 ;
  assign \g1331/_2_  = n104 ;
  assign \g971/_2_  = n111 ;
  assign \g973/_2_  = n114 ;
  assign \g975/_2_  = n119 ;
  assign \g983/_0_  = ~n125 ;
  assign \g984/_0_  = ~n130 ;
  assign \g985/_0_  = ~n135 ;
  assign \g991/_2_  = n142 ;
  assign \g993/_0_  = n145 ;
  assign \g997/_0_  = n150 ;
endmodule
