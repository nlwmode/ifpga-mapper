module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	output p_pad ;
	output q_pad ;
	output r_pad ;
	output s_pad ;
	output t_pad ;
	output u_pad ;
	output v_pad ;
	output w_pad ;
	output x_pad ;
	output y_pad ;
	output z_pad ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		e_pad,
		f_pad,
		_w15_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		c_pad,
		f_pad,
		_w16_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		c_pad,
		e_pad,
		_w17_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w16_,
		_w17_,
		_w18_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		d_pad,
		_w15_,
		_w19_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		_w18_,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		a_pad,
		b_pad,
		_w21_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		d_pad,
		e_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		o_pad,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w16_,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w21_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		a_pad,
		_w24_,
		_w26_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		b_pad,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		a_pad,
		b_pad,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w24_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		b_pad,
		_w26_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		j_pad,
		_w21_,
		_w31_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		f_pad,
		n_pad,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		o_pad,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		b_pad,
		m_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		b_pad,
		k_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		a_pad,
		l_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w34_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w35_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		a_pad,
		_w34_,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		l_pad,
		_w21_,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w35_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w39_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		i_pad,
		_w31_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w33_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		_w38_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w42_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		c_pad,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		f_pad,
		o_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		c_pad,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		d_pad,
		e_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		_w47_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		c_pad,
		_w33_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		_w51_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		g_pad,
		o_pad,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		c_pad,
		f_pad,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		d_pad,
		g_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w56_,
		_w57_,
		_w58_
	);
	assign p_pad = _w20_ ;
	assign q_pad = _w20_ ;
	assign r_pad = _w25_ ;
	assign s_pad = _w27_ ;
	assign t_pad = _w29_ ;
	assign u_pad = _w30_ ;
	assign v_pad = _w52_ ;
	assign w_pad = _w24_ ;
	assign x_pad = _w54_ ;
	assign y_pad = _w55_ ;
	assign z_pad = _w58_ ;
endmodule;