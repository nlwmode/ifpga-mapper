module top (\coda0_reg[0]/NET0131 , \coda0_reg[1]/NET0131 , \coda0_reg[2]/NET0131 , \coda1_reg[0]/NET0131 , \coda1_reg[1]/NET0131 , \coda1_reg[2]/NET0131 , \coda2_reg[0]/NET0131 , \coda2_reg[1]/NET0131 , \coda2_reg[2]/NET0131 , \coda3_reg[0]/NET0131 , \coda3_reg[1]/NET0131 , \coda3_reg[2]/NET0131 , \fu1_reg/NET0131 , \fu2_reg/NET0131 , \fu3_reg/NET0131 , \fu4_reg/NET0131 , \grant_o[0]_pad , \grant_o[1]_pad , \grant_o[2]_pad , \grant_o[3]_pad , \grant_reg[0]/NET0131 , \grant_reg[1]/NET0131 , \grant_reg[2]/NET0131 , \grant_reg[3]/NET0131 , \request1_pad , \request2_pad , \request3_pad , \request4_pad , \ru1_reg/NET0131 , \ru2_reg/NET0131 , \ru3_reg/NET0131 , \ru4_reg/NET0131 , \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , \_al_n0 , \_al_n1 , \g1143/_0_ , \g1144/_0_ , \g1145/_0_ , \g1146/_0_ , \g1147/_0_ , \g1148/_0_ , \g1149/_0_ , \g1150/_0_ , \g1151/_0_ , \g1152/_0_ , \g1153/_0_ , \g1154/_0_ , \g1174/_0_ , \g1175/_0_ , \g1176/_0_ , \g1177/_0_ , \g1238/_0_ , \g1239/_0_ , \g1240/_0_ , \g1241/_0_ , \g1242/_0_ , \g1243/_0_ , \g1244/_0_ , \g1245/_0_ , \g1247/_0_ , \g1248/_0_ , \g1249/_0_ , \g1250/_0_ , \g1520/_0_ );
	input \coda0_reg[0]/NET0131  ;
	input \coda0_reg[1]/NET0131  ;
	input \coda0_reg[2]/NET0131  ;
	input \coda1_reg[0]/NET0131  ;
	input \coda1_reg[1]/NET0131  ;
	input \coda1_reg[2]/NET0131  ;
	input \coda2_reg[0]/NET0131  ;
	input \coda2_reg[1]/NET0131  ;
	input \coda2_reg[2]/NET0131  ;
	input \coda3_reg[0]/NET0131  ;
	input \coda3_reg[1]/NET0131  ;
	input \coda3_reg[2]/NET0131  ;
	input \fu1_reg/NET0131  ;
	input \fu2_reg/NET0131  ;
	input \fu3_reg/NET0131  ;
	input \fu4_reg/NET0131  ;
	input \grant_o[0]_pad  ;
	input \grant_o[1]_pad  ;
	input \grant_o[2]_pad  ;
	input \grant_o[3]_pad  ;
	input \grant_reg[0]/NET0131  ;
	input \grant_reg[1]/NET0131  ;
	input \grant_reg[2]/NET0131  ;
	input \grant_reg[3]/NET0131  ;
	input \request1_pad  ;
	input \request2_pad  ;
	input \request3_pad  ;
	input \request4_pad  ;
	input \ru1_reg/NET0131  ;
	input \ru2_reg/NET0131  ;
	input \ru3_reg/NET0131  ;
	input \ru4_reg/NET0131  ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1143/_0_  ;
	output \g1144/_0_  ;
	output \g1145/_0_  ;
	output \g1146/_0_  ;
	output \g1147/_0_  ;
	output \g1148/_0_  ;
	output \g1149/_0_  ;
	output \g1150/_0_  ;
	output \g1151/_0_  ;
	output \g1152/_0_  ;
	output \g1153/_0_  ;
	output \g1154/_0_  ;
	output \g1174/_0_  ;
	output \g1175/_0_  ;
	output \g1176/_0_  ;
	output \g1177/_0_  ;
	output \g1238/_0_  ;
	output \g1239/_0_  ;
	output \g1240/_0_  ;
	output \g1241/_0_  ;
	output \g1242/_0_  ;
	output \g1243/_0_  ;
	output \g1244/_0_  ;
	output \g1245/_0_  ;
	output \g1247/_0_  ;
	output \g1248/_0_  ;
	output \g1249/_0_  ;
	output \g1250/_0_  ;
	output \g1520/_0_  ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\coda0_reg[2]/NET0131 ,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\coda0_reg[2]/NET0131 ,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\ru4_reg/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\coda0_reg[2]/NET0131 ,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w41_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\ru2_reg/NET0131 ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\ru1_reg/NET0131 ,
		_w39_,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w36_,
		_w37_,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\fu1_reg/NET0131 ,
		\fu2_reg/NET0131 ,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\fu3_reg/NET0131 ,
		\fu4_reg/NET0131 ,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\stato_reg[1]/NET0131 ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\coda0_reg[2]/NET0131 ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\coda1_reg[2]/NET0131 ,
		_w53_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\stato_reg[0]/NET0131 ,
		_w54_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w49_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\coda0_reg[0]/NET0131 ,
		_w35_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w41_,
		_w42_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\ru2_reg/NET0131 ,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\coda0_reg[0]/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w61_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\ru1_reg/NET0131 ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w59_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		_w37_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\coda0_reg[0]/NET0131 ,
		_w53_,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\coda1_reg[0]/NET0131 ,
		_w53_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\stato_reg[0]/NET0131 ,
		_w68_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w69_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w67_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\coda0_reg[1]/NET0131 ,
		_w35_,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		\coda0_reg[1]/NET0131 ,
		_w38_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\coda0_reg[1]/NET0131 ,
		_w42_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\ru2_reg/NET0131 ,
		_w41_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\ru1_reg/NET0131 ,
		_w74_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w77_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w73_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		_w37_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\coda0_reg[1]/NET0131 ,
		_w53_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\coda1_reg[1]/NET0131 ,
		_w53_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\stato_reg[0]/NET0131 ,
		_w82_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w81_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\ru1_reg/NET0131 ,
		_w37_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\coda0_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\coda1_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\ru3_reg/NET0131 ,
		_w88_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\fu4_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\coda1_reg[1]/NET0131 ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\coda0_reg[1]/NET0131 ,
		_w92_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\ru3_reg/NET0131 ,
		_w93_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w91_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\ru2_reg/NET0131 ,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\coda0_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\coda1_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\ru2_reg/NET0131 ,
		_w99_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w98_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w87_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\stato_reg[0]/NET0131 ,
		_w35_,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		\stato_reg[0]/NET0131 ,
		_w52_,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\stato_reg[1]/NET0131 ,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w105_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\coda1_reg[1]/NET0131 ,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\stato_reg[0]/NET0131 ,
		_w53_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\coda2_reg[1]/NET0131 ,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\ru1_reg/NET0131 ,
		_w37_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\fu1_reg/NET0131 ,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\coda0_reg[1]/NET0131 ,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w111_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w109_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w104_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\coda1_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\coda2_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w119_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\ru3_reg/NET0131 ,
		_w118_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\coda2_reg[2]/NET0131 ,
		_w92_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		\coda1_reg[2]/NET0131 ,
		_w92_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\ru3_reg/NET0131 ,
		_w122_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w121_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\ru2_reg/NET0131 ,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\coda1_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\coda2_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w129_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\ru2_reg/NET0131 ,
		_w128_,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w127_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w87_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\coda2_reg[2]/NET0131 ,
		_w108_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\coda3_reg[2]/NET0131 ,
		_w110_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		\coda1_reg[2]/NET0131 ,
		_w113_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w135_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w134_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w133_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\coda0_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\coda1_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\ru3_reg/NET0131 ,
		_w140_,
		_w142_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w141_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\coda1_reg[2]/NET0131 ,
		_w92_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\coda0_reg[2]/NET0131 ,
		_w92_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\ru3_reg/NET0131 ,
		_w144_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w143_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\ru2_reg/NET0131 ,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\coda0_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w150_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		\coda1_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\ru2_reg/NET0131 ,
		_w150_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w149_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		_w87_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		\coda1_reg[2]/NET0131 ,
		_w108_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\coda2_reg[2]/NET0131 ,
		_w110_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\coda0_reg[2]/NET0131 ,
		_w113_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w156_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w155_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		\coda0_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w162_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		\coda1_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		\ru3_reg/NET0131 ,
		_w162_,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\coda1_reg[0]/NET0131 ,
		_w92_,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		\coda0_reg[0]/NET0131 ,
		_w92_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\ru3_reg/NET0131 ,
		_w166_,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w167_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w165_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\ru2_reg/NET0131 ,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\coda0_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		\coda1_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\ru2_reg/NET0131 ,
		_w172_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w173_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w171_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		_w87_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\coda1_reg[0]/NET0131 ,
		_w108_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\coda2_reg[0]/NET0131 ,
		_w110_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\coda0_reg[0]/NET0131 ,
		_w113_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w179_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w178_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		_w177_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\coda1_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		\coda2_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w185_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\ru3_reg/NET0131 ,
		_w184_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\coda2_reg[0]/NET0131 ,
		_w92_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		\coda1_reg[0]/NET0131 ,
		_w92_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\ru3_reg/NET0131 ,
		_w188_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w187_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\ru2_reg/NET0131 ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\coda1_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\coda2_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w195_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		\ru2_reg/NET0131 ,
		_w194_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w193_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		_w87_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\coda2_reg[0]/NET0131 ,
		_w108_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\coda3_reg[0]/NET0131 ,
		_w110_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\coda1_reg[0]/NET0131 ,
		_w113_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		_w200_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w199_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		\coda1_reg[1]/NET0131 ,
		\fu1_reg/NET0131 ,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		\coda2_reg[1]/NET0131 ,
		\fu1_reg/NET0131 ,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w112_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\coda2_reg[1]/NET0131 ,
		_w53_,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		\coda3_reg[1]/NET0131 ,
		_w53_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\stato_reg[0]/NET0131 ,
		_w210_,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w211_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\coda1_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		\coda2_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\ru3_reg/NET0131 ,
		_w214_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\coda2_reg[1]/NET0131 ,
		_w92_,
		_w218_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		\coda1_reg[1]/NET0131 ,
		_w92_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\ru3_reg/NET0131 ,
		_w218_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		_w219_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w217_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\ru2_reg/NET0131 ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\coda1_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		\coda2_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w225_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\ru2_reg/NET0131 ,
		_w224_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		_w225_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w223_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		_w87_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w209_,
		_w213_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		_w229_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		\coda2_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		\coda3_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w234_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		\ru3_reg/NET0131 ,
		_w233_,
		_w235_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w234_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\coda3_reg[0]/NET0131 ,
		_w92_,
		_w237_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		\coda2_reg[0]/NET0131 ,
		_w92_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		\ru3_reg/NET0131 ,
		_w237_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w238_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w236_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		_w232_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\coda2_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		\coda3_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w245_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		_w243_,
		_w244_,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w245_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w242_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		_w37_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\coda3_reg[0]/NET0131 ,
		_w108_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		\coda2_reg[0]/NET0131 ,
		_w113_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w249_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		\coda2_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\coda3_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w255_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\ru3_reg/NET0131 ,
		_w254_,
		_w256_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w255_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\coda3_reg[1]/NET0131 ,
		_w92_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name224 (
		\coda2_reg[1]/NET0131 ,
		_w92_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		\ru3_reg/NET0131 ,
		_w258_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w259_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w257_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		_w232_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		\coda2_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		\coda3_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		_w243_,
		_w264_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		_w265_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w263_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		_w37_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\coda2_reg[1]/NET0131 ,
		_w113_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		\coda3_reg[1]/NET0131 ,
		_w108_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w270_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w269_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\coda2_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w274_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		\coda3_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		\ru3_reg/NET0131 ,
		_w274_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\coda3_reg[2]/NET0131 ,
		_w92_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		\coda2_reg[2]/NET0131 ,
		_w92_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\ru3_reg/NET0131 ,
		_w278_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w277_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		_w232_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		\coda2_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\coda3_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w285_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w243_,
		_w284_,
		_w286_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w285_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w283_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		_w37_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		\coda2_reg[2]/NET0131 ,
		_w113_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\coda3_reg[2]/NET0131 ,
		_w108_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		_w289_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name259 (
		\grant_reg[0]/NET0131 ,
		_w107_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\coda0_reg[1]/NET0131 ,
		_w110_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w294_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\grant_reg[1]/NET0131 ,
		_w107_,
		_w299_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		\coda0_reg[1]/NET0131 ,
		_w110_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w300_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w299_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\grant_reg[2]/NET0131 ,
		_w107_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w295_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w304_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\grant_reg[3]/NET0131 ,
		_w107_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name274 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w300_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w308_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\fu1_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w112_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		\ru2_reg/NET0131 ,
		_w37_,
		_w314_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\fu2_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		\ru3_reg/NET0131 ,
		_w37_,
		_w317_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		\fu3_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		\ru4_reg/NET0131 ,
		_w37_,
		_w320_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		\fu4_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\grant_reg[0]/NET0131 ,
		_w37_,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		\grant_o[0]_pad ,
		\stato_reg[0]/NET0131 ,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w323_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\grant_reg[1]/NET0131 ,
		_w37_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		\grant_o[1]_pad ,
		\stato_reg[0]/NET0131 ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w326_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\grant_reg[2]/NET0131 ,
		_w37_,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		\grant_o[2]_pad ,
		\stato_reg[0]/NET0131 ,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w329_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\grant_reg[3]/NET0131 ,
		_w37_,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		\grant_o[3]_pad ,
		\stato_reg[0]/NET0131 ,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w332_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\request1_pad ,
		\stato_reg[0]/NET0131 ,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w112_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		\request2_pad ,
		\stato_reg[0]/NET0131 ,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w314_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		\request3_pad ,
		\stato_reg[0]/NET0131 ,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w317_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		\request4_pad ,
		\stato_reg[0]/NET0131 ,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w320_,
		_w341_,
		_w342_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1143/_0_  = _w58_ ;
	assign \g1144/_0_  = _w72_ ;
	assign \g1145/_0_  = _w86_ ;
	assign \g1146/_0_  = _w117_ ;
	assign \g1147/_0_  = _w139_ ;
	assign \g1148/_0_  = _w161_ ;
	assign \g1149/_0_  = _w183_ ;
	assign \g1150/_0_  = _w205_ ;
	assign \g1151/_0_  = _w231_ ;
	assign \g1152/_0_  = _w253_ ;
	assign \g1153/_0_  = _w273_ ;
	assign \g1154/_0_  = _w293_ ;
	assign \g1174/_0_  = _w298_ ;
	assign \g1175/_0_  = _w303_ ;
	assign \g1176/_0_  = _w307_ ;
	assign \g1177/_0_  = _w311_ ;
	assign \g1238/_0_  = _w313_ ;
	assign \g1239/_0_  = _w316_ ;
	assign \g1240/_0_  = _w319_ ;
	assign \g1241/_0_  = _w322_ ;
	assign \g1242/_0_  = _w325_ ;
	assign \g1243/_0_  = _w328_ ;
	assign \g1244/_0_  = _w331_ ;
	assign \g1245/_0_  = _w334_ ;
	assign \g1247/_0_  = _w336_ ;
	assign \g1248/_0_  = _w338_ ;
	assign \g1249/_0_  = _w340_ ;
	assign \g1250/_0_  = _w342_ ;
	assign \g1520/_0_  = \stato_reg[0]/NET0131 ;
endmodule;