module top (\A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] , \A[1000] , maj);
	input \A[0]  ;
	input \A[1]  ;
	input \A[2]  ;
	input \A[3]  ;
	input \A[4]  ;
	input \A[5]  ;
	input \A[6]  ;
	input \A[7]  ;
	input \A[8]  ;
	input \A[9]  ;
	input \A[10]  ;
	input \A[11]  ;
	input \A[12]  ;
	input \A[13]  ;
	input \A[14]  ;
	input \A[15]  ;
	input \A[16]  ;
	input \A[17]  ;
	input \A[18]  ;
	input \A[19]  ;
	input \A[20]  ;
	input \A[21]  ;
	input \A[22]  ;
	input \A[23]  ;
	input \A[24]  ;
	input \A[25]  ;
	input \A[26]  ;
	input \A[27]  ;
	input \A[28]  ;
	input \A[29]  ;
	input \A[30]  ;
	input \A[31]  ;
	input \A[32]  ;
	input \A[33]  ;
	input \A[34]  ;
	input \A[35]  ;
	input \A[36]  ;
	input \A[37]  ;
	input \A[38]  ;
	input \A[39]  ;
	input \A[40]  ;
	input \A[41]  ;
	input \A[42]  ;
	input \A[43]  ;
	input \A[44]  ;
	input \A[45]  ;
	input \A[46]  ;
	input \A[47]  ;
	input \A[48]  ;
	input \A[49]  ;
	input \A[50]  ;
	input \A[51]  ;
	input \A[52]  ;
	input \A[53]  ;
	input \A[54]  ;
	input \A[55]  ;
	input \A[56]  ;
	input \A[57]  ;
	input \A[58]  ;
	input \A[59]  ;
	input \A[60]  ;
	input \A[61]  ;
	input \A[62]  ;
	input \A[63]  ;
	input \A[64]  ;
	input \A[65]  ;
	input \A[66]  ;
	input \A[67]  ;
	input \A[68]  ;
	input \A[69]  ;
	input \A[70]  ;
	input \A[71]  ;
	input \A[72]  ;
	input \A[73]  ;
	input \A[74]  ;
	input \A[75]  ;
	input \A[76]  ;
	input \A[77]  ;
	input \A[78]  ;
	input \A[79]  ;
	input \A[80]  ;
	input \A[81]  ;
	input \A[82]  ;
	input \A[83]  ;
	input \A[84]  ;
	input \A[85]  ;
	input \A[86]  ;
	input \A[87]  ;
	input \A[88]  ;
	input \A[89]  ;
	input \A[90]  ;
	input \A[91]  ;
	input \A[92]  ;
	input \A[93]  ;
	input \A[94]  ;
	input \A[95]  ;
	input \A[96]  ;
	input \A[97]  ;
	input \A[98]  ;
	input \A[99]  ;
	input \A[100]  ;
	input \A[101]  ;
	input \A[102]  ;
	input \A[103]  ;
	input \A[104]  ;
	input \A[105]  ;
	input \A[106]  ;
	input \A[107]  ;
	input \A[108]  ;
	input \A[109]  ;
	input \A[110]  ;
	input \A[111]  ;
	input \A[112]  ;
	input \A[113]  ;
	input \A[114]  ;
	input \A[115]  ;
	input \A[116]  ;
	input \A[117]  ;
	input \A[118]  ;
	input \A[119]  ;
	input \A[120]  ;
	input \A[121]  ;
	input \A[122]  ;
	input \A[123]  ;
	input \A[124]  ;
	input \A[125]  ;
	input \A[126]  ;
	input \A[127]  ;
	input \A[128]  ;
	input \A[129]  ;
	input \A[130]  ;
	input \A[131]  ;
	input \A[132]  ;
	input \A[133]  ;
	input \A[134]  ;
	input \A[135]  ;
	input \A[136]  ;
	input \A[137]  ;
	input \A[138]  ;
	input \A[139]  ;
	input \A[140]  ;
	input \A[141]  ;
	input \A[142]  ;
	input \A[143]  ;
	input \A[144]  ;
	input \A[145]  ;
	input \A[146]  ;
	input \A[147]  ;
	input \A[148]  ;
	input \A[149]  ;
	input \A[150]  ;
	input \A[151]  ;
	input \A[152]  ;
	input \A[153]  ;
	input \A[154]  ;
	input \A[155]  ;
	input \A[156]  ;
	input \A[157]  ;
	input \A[158]  ;
	input \A[159]  ;
	input \A[160]  ;
	input \A[161]  ;
	input \A[162]  ;
	input \A[163]  ;
	input \A[164]  ;
	input \A[165]  ;
	input \A[166]  ;
	input \A[167]  ;
	input \A[168]  ;
	input \A[169]  ;
	input \A[170]  ;
	input \A[171]  ;
	input \A[172]  ;
	input \A[173]  ;
	input \A[174]  ;
	input \A[175]  ;
	input \A[176]  ;
	input \A[177]  ;
	input \A[178]  ;
	input \A[179]  ;
	input \A[180]  ;
	input \A[181]  ;
	input \A[182]  ;
	input \A[183]  ;
	input \A[184]  ;
	input \A[185]  ;
	input \A[186]  ;
	input \A[187]  ;
	input \A[188]  ;
	input \A[189]  ;
	input \A[190]  ;
	input \A[191]  ;
	input \A[192]  ;
	input \A[193]  ;
	input \A[194]  ;
	input \A[195]  ;
	input \A[196]  ;
	input \A[197]  ;
	input \A[198]  ;
	input \A[199]  ;
	input \A[200]  ;
	input \A[201]  ;
	input \A[202]  ;
	input \A[203]  ;
	input \A[204]  ;
	input \A[205]  ;
	input \A[206]  ;
	input \A[207]  ;
	input \A[208]  ;
	input \A[209]  ;
	input \A[210]  ;
	input \A[211]  ;
	input \A[212]  ;
	input \A[213]  ;
	input \A[214]  ;
	input \A[215]  ;
	input \A[216]  ;
	input \A[217]  ;
	input \A[218]  ;
	input \A[219]  ;
	input \A[220]  ;
	input \A[221]  ;
	input \A[222]  ;
	input \A[223]  ;
	input \A[224]  ;
	input \A[225]  ;
	input \A[226]  ;
	input \A[227]  ;
	input \A[228]  ;
	input \A[229]  ;
	input \A[230]  ;
	input \A[231]  ;
	input \A[232]  ;
	input \A[233]  ;
	input \A[234]  ;
	input \A[235]  ;
	input \A[236]  ;
	input \A[237]  ;
	input \A[238]  ;
	input \A[239]  ;
	input \A[240]  ;
	input \A[241]  ;
	input \A[242]  ;
	input \A[243]  ;
	input \A[244]  ;
	input \A[245]  ;
	input \A[246]  ;
	input \A[247]  ;
	input \A[248]  ;
	input \A[249]  ;
	input \A[250]  ;
	input \A[251]  ;
	input \A[252]  ;
	input \A[253]  ;
	input \A[254]  ;
	input \A[255]  ;
	input \A[256]  ;
	input \A[257]  ;
	input \A[258]  ;
	input \A[259]  ;
	input \A[260]  ;
	input \A[261]  ;
	input \A[262]  ;
	input \A[263]  ;
	input \A[264]  ;
	input \A[265]  ;
	input \A[266]  ;
	input \A[267]  ;
	input \A[268]  ;
	input \A[269]  ;
	input \A[270]  ;
	input \A[271]  ;
	input \A[272]  ;
	input \A[273]  ;
	input \A[274]  ;
	input \A[275]  ;
	input \A[276]  ;
	input \A[277]  ;
	input \A[278]  ;
	input \A[279]  ;
	input \A[280]  ;
	input \A[281]  ;
	input \A[282]  ;
	input \A[283]  ;
	input \A[284]  ;
	input \A[285]  ;
	input \A[286]  ;
	input \A[287]  ;
	input \A[288]  ;
	input \A[289]  ;
	input \A[290]  ;
	input \A[291]  ;
	input \A[292]  ;
	input \A[293]  ;
	input \A[294]  ;
	input \A[295]  ;
	input \A[296]  ;
	input \A[297]  ;
	input \A[298]  ;
	input \A[299]  ;
	input \A[300]  ;
	input \A[301]  ;
	input \A[302]  ;
	input \A[303]  ;
	input \A[304]  ;
	input \A[305]  ;
	input \A[306]  ;
	input \A[307]  ;
	input \A[308]  ;
	input \A[309]  ;
	input \A[310]  ;
	input \A[311]  ;
	input \A[312]  ;
	input \A[313]  ;
	input \A[314]  ;
	input \A[315]  ;
	input \A[316]  ;
	input \A[317]  ;
	input \A[318]  ;
	input \A[319]  ;
	input \A[320]  ;
	input \A[321]  ;
	input \A[322]  ;
	input \A[323]  ;
	input \A[324]  ;
	input \A[325]  ;
	input \A[326]  ;
	input \A[327]  ;
	input \A[328]  ;
	input \A[329]  ;
	input \A[330]  ;
	input \A[331]  ;
	input \A[332]  ;
	input \A[333]  ;
	input \A[334]  ;
	input \A[335]  ;
	input \A[336]  ;
	input \A[337]  ;
	input \A[338]  ;
	input \A[339]  ;
	input \A[340]  ;
	input \A[341]  ;
	input \A[342]  ;
	input \A[343]  ;
	input \A[344]  ;
	input \A[345]  ;
	input \A[346]  ;
	input \A[347]  ;
	input \A[348]  ;
	input \A[349]  ;
	input \A[350]  ;
	input \A[351]  ;
	input \A[352]  ;
	input \A[353]  ;
	input \A[354]  ;
	input \A[355]  ;
	input \A[356]  ;
	input \A[357]  ;
	input \A[358]  ;
	input \A[359]  ;
	input \A[360]  ;
	input \A[361]  ;
	input \A[362]  ;
	input \A[363]  ;
	input \A[364]  ;
	input \A[365]  ;
	input \A[366]  ;
	input \A[367]  ;
	input \A[368]  ;
	input \A[369]  ;
	input \A[370]  ;
	input \A[371]  ;
	input \A[372]  ;
	input \A[373]  ;
	input \A[374]  ;
	input \A[375]  ;
	input \A[376]  ;
	input \A[377]  ;
	input \A[378]  ;
	input \A[379]  ;
	input \A[380]  ;
	input \A[381]  ;
	input \A[382]  ;
	input \A[383]  ;
	input \A[384]  ;
	input \A[385]  ;
	input \A[386]  ;
	input \A[387]  ;
	input \A[388]  ;
	input \A[389]  ;
	input \A[390]  ;
	input \A[391]  ;
	input \A[392]  ;
	input \A[393]  ;
	input \A[394]  ;
	input \A[395]  ;
	input \A[396]  ;
	input \A[397]  ;
	input \A[398]  ;
	input \A[399]  ;
	input \A[400]  ;
	input \A[401]  ;
	input \A[402]  ;
	input \A[403]  ;
	input \A[404]  ;
	input \A[405]  ;
	input \A[406]  ;
	input \A[407]  ;
	input \A[408]  ;
	input \A[409]  ;
	input \A[410]  ;
	input \A[411]  ;
	input \A[412]  ;
	input \A[413]  ;
	input \A[414]  ;
	input \A[415]  ;
	input \A[416]  ;
	input \A[417]  ;
	input \A[418]  ;
	input \A[419]  ;
	input \A[420]  ;
	input \A[421]  ;
	input \A[422]  ;
	input \A[423]  ;
	input \A[424]  ;
	input \A[425]  ;
	input \A[426]  ;
	input \A[427]  ;
	input \A[428]  ;
	input \A[429]  ;
	input \A[430]  ;
	input \A[431]  ;
	input \A[432]  ;
	input \A[433]  ;
	input \A[434]  ;
	input \A[435]  ;
	input \A[436]  ;
	input \A[437]  ;
	input \A[438]  ;
	input \A[439]  ;
	input \A[440]  ;
	input \A[441]  ;
	input \A[442]  ;
	input \A[443]  ;
	input \A[444]  ;
	input \A[445]  ;
	input \A[446]  ;
	input \A[447]  ;
	input \A[448]  ;
	input \A[449]  ;
	input \A[450]  ;
	input \A[451]  ;
	input \A[452]  ;
	input \A[453]  ;
	input \A[454]  ;
	input \A[455]  ;
	input \A[456]  ;
	input \A[457]  ;
	input \A[458]  ;
	input \A[459]  ;
	input \A[460]  ;
	input \A[461]  ;
	input \A[462]  ;
	input \A[463]  ;
	input \A[464]  ;
	input \A[465]  ;
	input \A[466]  ;
	input \A[467]  ;
	input \A[468]  ;
	input \A[469]  ;
	input \A[470]  ;
	input \A[471]  ;
	input \A[472]  ;
	input \A[473]  ;
	input \A[474]  ;
	input \A[475]  ;
	input \A[476]  ;
	input \A[477]  ;
	input \A[478]  ;
	input \A[479]  ;
	input \A[480]  ;
	input \A[481]  ;
	input \A[482]  ;
	input \A[483]  ;
	input \A[484]  ;
	input \A[485]  ;
	input \A[486]  ;
	input \A[487]  ;
	input \A[488]  ;
	input \A[489]  ;
	input \A[490]  ;
	input \A[491]  ;
	input \A[492]  ;
	input \A[493]  ;
	input \A[494]  ;
	input \A[495]  ;
	input \A[496]  ;
	input \A[497]  ;
	input \A[498]  ;
	input \A[499]  ;
	input \A[500]  ;
	input \A[501]  ;
	input \A[502]  ;
	input \A[503]  ;
	input \A[504]  ;
	input \A[505]  ;
	input \A[506]  ;
	input \A[507]  ;
	input \A[508]  ;
	input \A[509]  ;
	input \A[510]  ;
	input \A[511]  ;
	input \A[512]  ;
	input \A[513]  ;
	input \A[514]  ;
	input \A[515]  ;
	input \A[516]  ;
	input \A[517]  ;
	input \A[518]  ;
	input \A[519]  ;
	input \A[520]  ;
	input \A[521]  ;
	input \A[522]  ;
	input \A[523]  ;
	input \A[524]  ;
	input \A[525]  ;
	input \A[526]  ;
	input \A[527]  ;
	input \A[528]  ;
	input \A[529]  ;
	input \A[530]  ;
	input \A[531]  ;
	input \A[532]  ;
	input \A[533]  ;
	input \A[534]  ;
	input \A[535]  ;
	input \A[536]  ;
	input \A[537]  ;
	input \A[538]  ;
	input \A[539]  ;
	input \A[540]  ;
	input \A[541]  ;
	input \A[542]  ;
	input \A[543]  ;
	input \A[544]  ;
	input \A[545]  ;
	input \A[546]  ;
	input \A[547]  ;
	input \A[548]  ;
	input \A[549]  ;
	input \A[550]  ;
	input \A[551]  ;
	input \A[552]  ;
	input \A[553]  ;
	input \A[554]  ;
	input \A[555]  ;
	input \A[556]  ;
	input \A[557]  ;
	input \A[558]  ;
	input \A[559]  ;
	input \A[560]  ;
	input \A[561]  ;
	input \A[562]  ;
	input \A[563]  ;
	input \A[564]  ;
	input \A[565]  ;
	input \A[566]  ;
	input \A[567]  ;
	input \A[568]  ;
	input \A[569]  ;
	input \A[570]  ;
	input \A[571]  ;
	input \A[572]  ;
	input \A[573]  ;
	input \A[574]  ;
	input \A[575]  ;
	input \A[576]  ;
	input \A[577]  ;
	input \A[578]  ;
	input \A[579]  ;
	input \A[580]  ;
	input \A[581]  ;
	input \A[582]  ;
	input \A[583]  ;
	input \A[584]  ;
	input \A[585]  ;
	input \A[586]  ;
	input \A[587]  ;
	input \A[588]  ;
	input \A[589]  ;
	input \A[590]  ;
	input \A[591]  ;
	input \A[592]  ;
	input \A[593]  ;
	input \A[594]  ;
	input \A[595]  ;
	input \A[596]  ;
	input \A[597]  ;
	input \A[598]  ;
	input \A[599]  ;
	input \A[600]  ;
	input \A[601]  ;
	input \A[602]  ;
	input \A[603]  ;
	input \A[604]  ;
	input \A[605]  ;
	input \A[606]  ;
	input \A[607]  ;
	input \A[608]  ;
	input \A[609]  ;
	input \A[610]  ;
	input \A[611]  ;
	input \A[612]  ;
	input \A[613]  ;
	input \A[614]  ;
	input \A[615]  ;
	input \A[616]  ;
	input \A[617]  ;
	input \A[618]  ;
	input \A[619]  ;
	input \A[620]  ;
	input \A[621]  ;
	input \A[622]  ;
	input \A[623]  ;
	input \A[624]  ;
	input \A[625]  ;
	input \A[626]  ;
	input \A[627]  ;
	input \A[628]  ;
	input \A[629]  ;
	input \A[630]  ;
	input \A[631]  ;
	input \A[632]  ;
	input \A[633]  ;
	input \A[634]  ;
	input \A[635]  ;
	input \A[636]  ;
	input \A[637]  ;
	input \A[638]  ;
	input \A[639]  ;
	input \A[640]  ;
	input \A[641]  ;
	input \A[642]  ;
	input \A[643]  ;
	input \A[644]  ;
	input \A[645]  ;
	input \A[646]  ;
	input \A[647]  ;
	input \A[648]  ;
	input \A[649]  ;
	input \A[650]  ;
	input \A[651]  ;
	input \A[652]  ;
	input \A[653]  ;
	input \A[654]  ;
	input \A[655]  ;
	input \A[656]  ;
	input \A[657]  ;
	input \A[658]  ;
	input \A[659]  ;
	input \A[660]  ;
	input \A[661]  ;
	input \A[662]  ;
	input \A[663]  ;
	input \A[664]  ;
	input \A[665]  ;
	input \A[666]  ;
	input \A[667]  ;
	input \A[668]  ;
	input \A[669]  ;
	input \A[670]  ;
	input \A[671]  ;
	input \A[672]  ;
	input \A[673]  ;
	input \A[674]  ;
	input \A[675]  ;
	input \A[676]  ;
	input \A[677]  ;
	input \A[678]  ;
	input \A[679]  ;
	input \A[680]  ;
	input \A[681]  ;
	input \A[682]  ;
	input \A[683]  ;
	input \A[684]  ;
	input \A[685]  ;
	input \A[686]  ;
	input \A[687]  ;
	input \A[688]  ;
	input \A[689]  ;
	input \A[690]  ;
	input \A[691]  ;
	input \A[692]  ;
	input \A[693]  ;
	input \A[694]  ;
	input \A[695]  ;
	input \A[696]  ;
	input \A[697]  ;
	input \A[698]  ;
	input \A[699]  ;
	input \A[700]  ;
	input \A[701]  ;
	input \A[702]  ;
	input \A[703]  ;
	input \A[704]  ;
	input \A[705]  ;
	input \A[706]  ;
	input \A[707]  ;
	input \A[708]  ;
	input \A[709]  ;
	input \A[710]  ;
	input \A[711]  ;
	input \A[712]  ;
	input \A[713]  ;
	input \A[714]  ;
	input \A[715]  ;
	input \A[716]  ;
	input \A[717]  ;
	input \A[718]  ;
	input \A[719]  ;
	input \A[720]  ;
	input \A[721]  ;
	input \A[722]  ;
	input \A[723]  ;
	input \A[724]  ;
	input \A[725]  ;
	input \A[726]  ;
	input \A[727]  ;
	input \A[728]  ;
	input \A[729]  ;
	input \A[730]  ;
	input \A[731]  ;
	input \A[732]  ;
	input \A[733]  ;
	input \A[734]  ;
	input \A[735]  ;
	input \A[736]  ;
	input \A[737]  ;
	input \A[738]  ;
	input \A[739]  ;
	input \A[740]  ;
	input \A[741]  ;
	input \A[742]  ;
	input \A[743]  ;
	input \A[744]  ;
	input \A[745]  ;
	input \A[746]  ;
	input \A[747]  ;
	input \A[748]  ;
	input \A[749]  ;
	input \A[750]  ;
	input \A[751]  ;
	input \A[752]  ;
	input \A[753]  ;
	input \A[754]  ;
	input \A[755]  ;
	input \A[756]  ;
	input \A[757]  ;
	input \A[758]  ;
	input \A[759]  ;
	input \A[760]  ;
	input \A[761]  ;
	input \A[762]  ;
	input \A[763]  ;
	input \A[764]  ;
	input \A[765]  ;
	input \A[766]  ;
	input \A[767]  ;
	input \A[768]  ;
	input \A[769]  ;
	input \A[770]  ;
	input \A[771]  ;
	input \A[772]  ;
	input \A[773]  ;
	input \A[774]  ;
	input \A[775]  ;
	input \A[776]  ;
	input \A[777]  ;
	input \A[778]  ;
	input \A[779]  ;
	input \A[780]  ;
	input \A[781]  ;
	input \A[782]  ;
	input \A[783]  ;
	input \A[784]  ;
	input \A[785]  ;
	input \A[786]  ;
	input \A[787]  ;
	input \A[788]  ;
	input \A[789]  ;
	input \A[790]  ;
	input \A[791]  ;
	input \A[792]  ;
	input \A[793]  ;
	input \A[794]  ;
	input \A[795]  ;
	input \A[796]  ;
	input \A[797]  ;
	input \A[798]  ;
	input \A[799]  ;
	input \A[800]  ;
	input \A[801]  ;
	input \A[802]  ;
	input \A[803]  ;
	input \A[804]  ;
	input \A[805]  ;
	input \A[806]  ;
	input \A[807]  ;
	input \A[808]  ;
	input \A[809]  ;
	input \A[810]  ;
	input \A[811]  ;
	input \A[812]  ;
	input \A[813]  ;
	input \A[814]  ;
	input \A[815]  ;
	input \A[816]  ;
	input \A[817]  ;
	input \A[818]  ;
	input \A[819]  ;
	input \A[820]  ;
	input \A[821]  ;
	input \A[822]  ;
	input \A[823]  ;
	input \A[824]  ;
	input \A[825]  ;
	input \A[826]  ;
	input \A[827]  ;
	input \A[828]  ;
	input \A[829]  ;
	input \A[830]  ;
	input \A[831]  ;
	input \A[832]  ;
	input \A[833]  ;
	input \A[834]  ;
	input \A[835]  ;
	input \A[836]  ;
	input \A[837]  ;
	input \A[838]  ;
	input \A[839]  ;
	input \A[840]  ;
	input \A[841]  ;
	input \A[842]  ;
	input \A[843]  ;
	input \A[844]  ;
	input \A[845]  ;
	input \A[846]  ;
	input \A[847]  ;
	input \A[848]  ;
	input \A[849]  ;
	input \A[850]  ;
	input \A[851]  ;
	input \A[852]  ;
	input \A[853]  ;
	input \A[854]  ;
	input \A[855]  ;
	input \A[856]  ;
	input \A[857]  ;
	input \A[858]  ;
	input \A[859]  ;
	input \A[860]  ;
	input \A[861]  ;
	input \A[862]  ;
	input \A[863]  ;
	input \A[864]  ;
	input \A[865]  ;
	input \A[866]  ;
	input \A[867]  ;
	input \A[868]  ;
	input \A[869]  ;
	input \A[870]  ;
	input \A[871]  ;
	input \A[872]  ;
	input \A[873]  ;
	input \A[874]  ;
	input \A[875]  ;
	input \A[876]  ;
	input \A[877]  ;
	input \A[878]  ;
	input \A[879]  ;
	input \A[880]  ;
	input \A[881]  ;
	input \A[882]  ;
	input \A[883]  ;
	input \A[884]  ;
	input \A[885]  ;
	input \A[886]  ;
	input \A[887]  ;
	input \A[888]  ;
	input \A[889]  ;
	input \A[890]  ;
	input \A[891]  ;
	input \A[892]  ;
	input \A[893]  ;
	input \A[894]  ;
	input \A[895]  ;
	input \A[896]  ;
	input \A[897]  ;
	input \A[898]  ;
	input \A[899]  ;
	input \A[900]  ;
	input \A[901]  ;
	input \A[902]  ;
	input \A[903]  ;
	input \A[904]  ;
	input \A[905]  ;
	input \A[906]  ;
	input \A[907]  ;
	input \A[908]  ;
	input \A[909]  ;
	input \A[910]  ;
	input \A[911]  ;
	input \A[912]  ;
	input \A[913]  ;
	input \A[914]  ;
	input \A[915]  ;
	input \A[916]  ;
	input \A[917]  ;
	input \A[918]  ;
	input \A[919]  ;
	input \A[920]  ;
	input \A[921]  ;
	input \A[922]  ;
	input \A[923]  ;
	input \A[924]  ;
	input \A[925]  ;
	input \A[926]  ;
	input \A[927]  ;
	input \A[928]  ;
	input \A[929]  ;
	input \A[930]  ;
	input \A[931]  ;
	input \A[932]  ;
	input \A[933]  ;
	input \A[934]  ;
	input \A[935]  ;
	input \A[936]  ;
	input \A[937]  ;
	input \A[938]  ;
	input \A[939]  ;
	input \A[940]  ;
	input \A[941]  ;
	input \A[942]  ;
	input \A[943]  ;
	input \A[944]  ;
	input \A[945]  ;
	input \A[946]  ;
	input \A[947]  ;
	input \A[948]  ;
	input \A[949]  ;
	input \A[950]  ;
	input \A[951]  ;
	input \A[952]  ;
	input \A[953]  ;
	input \A[954]  ;
	input \A[955]  ;
	input \A[956]  ;
	input \A[957]  ;
	input \A[958]  ;
	input \A[959]  ;
	input \A[960]  ;
	input \A[961]  ;
	input \A[962]  ;
	input \A[963]  ;
	input \A[964]  ;
	input \A[965]  ;
	input \A[966]  ;
	input \A[967]  ;
	input \A[968]  ;
	input \A[969]  ;
	input \A[970]  ;
	input \A[971]  ;
	input \A[972]  ;
	input \A[973]  ;
	input \A[974]  ;
	input \A[975]  ;
	input \A[976]  ;
	input \A[977]  ;
	input \A[978]  ;
	input \A[979]  ;
	input \A[980]  ;
	input \A[981]  ;
	input \A[982]  ;
	input \A[983]  ;
	input \A[984]  ;
	input \A[985]  ;
	input \A[986]  ;
	input \A[987]  ;
	input \A[988]  ;
	input \A[989]  ;
	input \A[990]  ;
	input \A[991]  ;
	input \A[992]  ;
	input \A[993]  ;
	input \A[994]  ;
	input \A[995]  ;
	input \A[996]  ;
	input \A[997]  ;
	input \A[998]  ;
	input \A[999]  ;
	input \A[1000]  ;
	output maj ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	LUT3 #(
		.INIT('h17)
	) name0 (
		\A[67] ,
		\A[68] ,
		\A[69] ,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\A[70] ,
		\A[71] ,
		_w1004_
	);
	LUT3 #(
		.INIT('h96)
	) name2 (
		\A[67] ,
		\A[68] ,
		\A[69] ,
		_w1005_
	);
	LUT3 #(
		.INIT('h96)
	) name3 (
		\A[70] ,
		\A[71] ,
		\A[72] ,
		_w1006_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		_w1004_,
		_w1005_,
		_w1006_,
		_w1007_
	);
	LUT3 #(
		.INIT('h17)
	) name5 (
		\A[70] ,
		\A[71] ,
		\A[72] ,
		_w1008_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name6 (
		\A[70] ,
		\A[71] ,
		\A[72] ,
		_w1005_,
		_w1009_
	);
	LUT2 #(
		.INIT('h9)
	) name7 (
		_w1003_,
		_w1009_,
		_w1010_
	);
	LUT3 #(
		.INIT('h96)
	) name8 (
		\A[73] ,
		\A[74] ,
		\A[75] ,
		_w1011_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\A[76] ,
		\A[77] ,
		_w1012_
	);
	LUT3 #(
		.INIT('h96)
	) name10 (
		\A[76] ,
		\A[77] ,
		\A[78] ,
		_w1013_
	);
	LUT3 #(
		.INIT('h17)
	) name11 (
		\A[76] ,
		\A[77] ,
		\A[78] ,
		_w1014_
	);
	LUT3 #(
		.INIT('h17)
	) name12 (
		\A[73] ,
		\A[74] ,
		\A[75] ,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w1014_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h6)
	) name14 (
		_w1014_,
		_w1015_,
		_w1017_
	);
	LUT4 #(
		.INIT('h8008)
	) name15 (
		_w1011_,
		_w1013_,
		_w1014_,
		_w1015_,
		_w1018_
	);
	LUT4 #(
		.INIT('h0770)
	) name16 (
		_w1011_,
		_w1013_,
		_w1014_,
		_w1015_,
		_w1019_
	);
	LUT4 #(
		.INIT('h0660)
	) name17 (
		_w1005_,
		_w1006_,
		_w1011_,
		_w1013_,
		_w1020_
	);
	LUT3 #(
		.INIT('h01)
	) name18 (
		_w1019_,
		_w1020_,
		_w1018_,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w1017_,
		_w1020_,
		_w1022_
	);
	LUT4 #(
		.INIT('h4000)
	) name20 (
		_w1003_,
		_w1004_,
		_w1005_,
		_w1006_,
		_w1023_
	);
	LUT3 #(
		.INIT('h08)
	) name21 (
		_w1017_,
		_w1020_,
		_w1023_,
		_w1024_
	);
	LUT4 #(
		.INIT('h80a0)
	) name22 (
		_w1011_,
		_w1012_,
		_w1013_,
		_w1015_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w1016_,
		_w1025_,
		_w1026_
	);
	LUT4 #(
		.INIT('h00f2)
	) name24 (
		_w1010_,
		_w1021_,
		_w1024_,
		_w1026_,
		_w1027_
	);
	LUT4 #(
		.INIT('h4055)
	) name25 (
		_w1003_,
		_w1005_,
		_w1006_,
		_w1008_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w1007_,
		_w1028_,
		_w1029_
	);
	LUT4 #(
		.INIT('h0d00)
	) name27 (
		_w1010_,
		_w1021_,
		_w1024_,
		_w1026_,
		_w1030_
	);
	LUT3 #(
		.INIT('h54)
	) name28 (
		_w1027_,
		_w1029_,
		_w1030_,
		_w1031_
	);
	LUT3 #(
		.INIT('h96)
	) name29 (
		\A[61] ,
		\A[62] ,
		\A[63] ,
		_w1032_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\A[64] ,
		\A[65] ,
		_w1033_
	);
	LUT3 #(
		.INIT('h96)
	) name31 (
		\A[64] ,
		\A[65] ,
		\A[66] ,
		_w1034_
	);
	LUT3 #(
		.INIT('h96)
	) name32 (
		\A[55] ,
		\A[56] ,
		\A[57] ,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\A[58] ,
		\A[59] ,
		_w1036_
	);
	LUT3 #(
		.INIT('h96)
	) name34 (
		\A[58] ,
		\A[59] ,
		\A[60] ,
		_w1037_
	);
	LUT4 #(
		.INIT('h0660)
	) name35 (
		_w1032_,
		_w1034_,
		_w1035_,
		_w1037_,
		_w1038_
	);
	LUT3 #(
		.INIT('h17)
	) name36 (
		\A[61] ,
		\A[62] ,
		\A[63] ,
		_w1039_
	);
	LUT3 #(
		.INIT('h17)
	) name37 (
		\A[64] ,
		\A[65] ,
		\A[66] ,
		_w1040_
	);
	LUT3 #(
		.INIT('h80)
	) name38 (
		_w1032_,
		_w1033_,
		_w1034_,
		_w1041_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name39 (
		\A[64] ,
		\A[65] ,
		\A[66] ,
		_w1032_,
		_w1042_
	);
	LUT2 #(
		.INIT('h9)
	) name40 (
		_w1039_,
		_w1042_,
		_w1043_
	);
	LUT3 #(
		.INIT('h14)
	) name41 (
		_w1038_,
		_w1039_,
		_w1042_,
		_w1044_
	);
	LUT3 #(
		.INIT('h17)
	) name42 (
		\A[55] ,
		\A[56] ,
		\A[57] ,
		_w1045_
	);
	LUT3 #(
		.INIT('h80)
	) name43 (
		_w1035_,
		_w1036_,
		_w1037_,
		_w1046_
	);
	LUT3 #(
		.INIT('h17)
	) name44 (
		\A[58] ,
		\A[59] ,
		\A[60] ,
		_w1047_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name45 (
		\A[58] ,
		\A[59] ,
		\A[60] ,
		_w1035_,
		_w1048_
	);
	LUT2 #(
		.INIT('h9)
	) name46 (
		_w1045_,
		_w1048_,
		_w1049_
	);
	LUT3 #(
		.INIT('h82)
	) name47 (
		_w1038_,
		_w1039_,
		_w1042_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w1039_,
		_w1040_,
		_w1051_
	);
	LUT4 #(
		.INIT('h0080)
	) name49 (
		_w1035_,
		_w1036_,
		_w1037_,
		_w1045_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w1051_,
		_w1052_,
		_w1053_
	);
	LUT4 #(
		.INIT('h171f)
	) name51 (
		_w1038_,
		_w1043_,
		_w1049_,
		_w1053_,
		_w1054_
	);
	LUT4 #(
		.INIT('h080f)
	) name52 (
		_w1032_,
		_w1034_,
		_w1039_,
		_w1040_,
		_w1055_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w1041_,
		_w1055_,
		_w1056_
	);
	LUT4 #(
		.INIT('h080f)
	) name54 (
		_w1035_,
		_w1037_,
		_w1045_,
		_w1047_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w1046_,
		_w1057_,
		_w1058_
	);
	LUT3 #(
		.INIT('he8)
	) name56 (
		_w1054_,
		_w1056_,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w1031_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w1031_,
		_w1059_,
		_w1061_
	);
	LUT3 #(
		.INIT('h69)
	) name59 (
		_w1054_,
		_w1056_,
		_w1058_,
		_w1062_
	);
	LUT4 #(
		.INIT('hf20d)
	) name60 (
		_w1010_,
		_w1021_,
		_w1024_,
		_w1026_,
		_w1063_
	);
	LUT2 #(
		.INIT('h9)
	) name61 (
		_w1029_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('h6996)
	) name62 (
		_w1005_,
		_w1006_,
		_w1011_,
		_w1013_,
		_w1065_
	);
	LUT4 #(
		.INIT('h6996)
	) name63 (
		_w1032_,
		_w1034_,
		_w1035_,
		_w1037_,
		_w1066_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w1065_,
		_w1066_,
		_w1067_
	);
	LUT4 #(
		.INIT('h89a9)
	) name65 (
		_w1010_,
		_w1021_,
		_w1022_,
		_w1023_,
		_w1068_
	);
	LUT4 #(
		.INIT('hc989)
	) name66 (
		_w1044_,
		_w1049_,
		_w1050_,
		_w1053_,
		_w1069_
	);
	LUT3 #(
		.INIT('he8)
	) name67 (
		_w1067_,
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT3 #(
		.INIT('he8)
	) name68 (
		_w1062_,
		_w1064_,
		_w1070_,
		_w1071_
	);
	LUT3 #(
		.INIT('h54)
	) name69 (
		_w1060_,
		_w1061_,
		_w1071_,
		_w1072_
	);
	LUT3 #(
		.INIT('h17)
	) name70 (
		\A[43] ,
		\A[44] ,
		\A[45] ,
		_w1073_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\A[46] ,
		\A[47] ,
		_w1074_
	);
	LUT3 #(
		.INIT('h96)
	) name72 (
		\A[43] ,
		\A[44] ,
		\A[45] ,
		_w1075_
	);
	LUT3 #(
		.INIT('h96)
	) name73 (
		\A[46] ,
		\A[47] ,
		\A[48] ,
		_w1076_
	);
	LUT3 #(
		.INIT('h80)
	) name74 (
		_w1074_,
		_w1075_,
		_w1076_,
		_w1077_
	);
	LUT3 #(
		.INIT('h17)
	) name75 (
		\A[46] ,
		\A[47] ,
		\A[48] ,
		_w1078_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name76 (
		\A[46] ,
		\A[47] ,
		\A[48] ,
		_w1075_,
		_w1079_
	);
	LUT2 #(
		.INIT('h9)
	) name77 (
		_w1073_,
		_w1079_,
		_w1080_
	);
	LUT3 #(
		.INIT('h96)
	) name78 (
		\A[49] ,
		\A[50] ,
		\A[51] ,
		_w1081_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\A[52] ,
		\A[53] ,
		_w1082_
	);
	LUT3 #(
		.INIT('h96)
	) name80 (
		\A[52] ,
		\A[53] ,
		\A[54] ,
		_w1083_
	);
	LUT3 #(
		.INIT('h17)
	) name81 (
		\A[52] ,
		\A[53] ,
		\A[54] ,
		_w1084_
	);
	LUT3 #(
		.INIT('h17)
	) name82 (
		\A[49] ,
		\A[50] ,
		\A[51] ,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w1084_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h6)
	) name84 (
		_w1084_,
		_w1085_,
		_w1087_
	);
	LUT4 #(
		.INIT('h8008)
	) name85 (
		_w1081_,
		_w1083_,
		_w1084_,
		_w1085_,
		_w1088_
	);
	LUT4 #(
		.INIT('h0770)
	) name86 (
		_w1081_,
		_w1083_,
		_w1084_,
		_w1085_,
		_w1089_
	);
	LUT4 #(
		.INIT('h0660)
	) name87 (
		_w1075_,
		_w1076_,
		_w1081_,
		_w1083_,
		_w1090_
	);
	LUT3 #(
		.INIT('h01)
	) name88 (
		_w1089_,
		_w1090_,
		_w1088_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w1087_,
		_w1090_,
		_w1092_
	);
	LUT4 #(
		.INIT('h4000)
	) name90 (
		_w1073_,
		_w1074_,
		_w1075_,
		_w1076_,
		_w1093_
	);
	LUT3 #(
		.INIT('h08)
	) name91 (
		_w1087_,
		_w1090_,
		_w1093_,
		_w1094_
	);
	LUT3 #(
		.INIT('h0d)
	) name92 (
		_w1080_,
		_w1091_,
		_w1094_,
		_w1095_
	);
	LUT4 #(
		.INIT('h80a0)
	) name93 (
		_w1081_,
		_w1082_,
		_w1083_,
		_w1085_,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w1086_,
		_w1096_,
		_w1097_
	);
	LUT4 #(
		.INIT('h00f2)
	) name95 (
		_w1080_,
		_w1091_,
		_w1094_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h4055)
	) name96 (
		_w1073_,
		_w1075_,
		_w1076_,
		_w1078_,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w1077_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('h0d00)
	) name98 (
		_w1080_,
		_w1091_,
		_w1094_,
		_w1097_,
		_w1101_
	);
	LUT3 #(
		.INIT('h96)
	) name99 (
		\A[37] ,
		\A[38] ,
		\A[39] ,
		_w1102_
	);
	LUT3 #(
		.INIT('h96)
	) name100 (
		\A[40] ,
		\A[41] ,
		\A[42] ,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT3 #(
		.INIT('h96)
	) name102 (
		\A[31] ,
		\A[32] ,
		\A[33] ,
		_w1105_
	);
	LUT3 #(
		.INIT('h96)
	) name103 (
		\A[34] ,
		\A[35] ,
		\A[36] ,
		_w1106_
	);
	LUT4 #(
		.INIT('h0660)
	) name104 (
		_w1102_,
		_w1103_,
		_w1105_,
		_w1106_,
		_w1107_
	);
	LUT3 #(
		.INIT('h17)
	) name105 (
		\A[40] ,
		\A[41] ,
		\A[42] ,
		_w1108_
	);
	LUT3 #(
		.INIT('h17)
	) name106 (
		\A[37] ,
		\A[38] ,
		\A[39] ,
		_w1109_
	);
	LUT2 #(
		.INIT('h6)
	) name107 (
		_w1108_,
		_w1109_,
		_w1110_
	);
	LUT3 #(
		.INIT('h17)
	) name108 (
		\A[34] ,
		\A[35] ,
		\A[36] ,
		_w1111_
	);
	LUT3 #(
		.INIT('h17)
	) name109 (
		\A[31] ,
		\A[32] ,
		\A[33] ,
		_w1112_
	);
	LUT4 #(
		.INIT('h7887)
	) name110 (
		_w1105_,
		_w1106_,
		_w1111_,
		_w1112_,
		_w1113_
	);
	LUT4 #(
		.INIT('hc0de)
	) name111 (
		_w1104_,
		_w1107_,
		_w1110_,
		_w1113_,
		_w1114_
	);
	LUT4 #(
		.INIT('h088f)
	) name112 (
		_w1102_,
		_w1103_,
		_w1108_,
		_w1109_,
		_w1115_
	);
	LUT4 #(
		.INIT('h088f)
	) name113 (
		_w1105_,
		_w1106_,
		_w1111_,
		_w1112_,
		_w1116_
	);
	LUT3 #(
		.INIT('he8)
	) name114 (
		_w1114_,
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT4 #(
		.INIT('h1700)
	) name115 (
		_w1095_,
		_w1097_,
		_w1100_,
		_w1117_,
		_w1118_
	);
	LUT4 #(
		.INIT('h00e8)
	) name116 (
		_w1095_,
		_w1097_,
		_w1100_,
		_w1117_,
		_w1119_
	);
	LUT4 #(
		.INIT('hf20d)
	) name117 (
		_w1080_,
		_w1091_,
		_w1094_,
		_w1097_,
		_w1120_
	);
	LUT3 #(
		.INIT('h69)
	) name118 (
		_w1114_,
		_w1115_,
		_w1116_,
		_w1121_
	);
	LUT3 #(
		.INIT('h09)
	) name119 (
		_w1100_,
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT3 #(
		.INIT('h60)
	) name120 (
		_w1100_,
		_w1120_,
		_w1121_,
		_w1123_
	);
	LUT4 #(
		.INIT('h6996)
	) name121 (
		_w1075_,
		_w1076_,
		_w1081_,
		_w1083_,
		_w1124_
	);
	LUT4 #(
		.INIT('h6996)
	) name122 (
		_w1102_,
		_w1103_,
		_w1105_,
		_w1106_,
		_w1125_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT4 #(
		.INIT('h89a9)
	) name124 (
		_w1080_,
		_w1091_,
		_w1092_,
		_w1093_,
		_w1127_
	);
	LUT4 #(
		.INIT('he11e)
	) name125 (
		_w1104_,
		_w1107_,
		_w1110_,
		_w1113_,
		_w1128_
	);
	LUT3 #(
		.INIT('h71)
	) name126 (
		_w1126_,
		_w1127_,
		_w1128_,
		_w1129_
	);
	LUT4 #(
		.INIT('h4445)
	) name127 (
		_w1119_,
		_w1122_,
		_w1123_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w1118_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		_w1072_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w1072_,
		_w1131_,
		_w1133_
	);
	LUT2 #(
		.INIT('h6)
	) name131 (
		_w1031_,
		_w1059_,
		_w1134_
	);
	LUT4 #(
		.INIT('h54ab)
	) name132 (
		_w1098_,
		_w1100_,
		_w1101_,
		_w1117_,
		_w1135_
	);
	LUT4 #(
		.INIT('h54ab)
	) name133 (
		_w1122_,
		_w1123_,
		_w1129_,
		_w1135_,
		_w1136_
	);
	LUT3 #(
		.INIT('h09)
	) name134 (
		_w1071_,
		_w1134_,
		_w1136_,
		_w1137_
	);
	LUT3 #(
		.INIT('h60)
	) name135 (
		_w1071_,
		_w1134_,
		_w1136_,
		_w1138_
	);
	LUT3 #(
		.INIT('h96)
	) name136 (
		_w1062_,
		_w1064_,
		_w1070_,
		_w1139_
	);
	LUT3 #(
		.INIT('h96)
	) name137 (
		_w1100_,
		_w1120_,
		_w1121_,
		_w1140_
	);
	LUT2 #(
		.INIT('h9)
	) name138 (
		_w1129_,
		_w1140_,
		_w1141_
	);
	LUT4 #(
		.INIT('h0660)
	) name139 (
		_w1065_,
		_w1066_,
		_w1124_,
		_w1125_,
		_w1142_
	);
	LUT4 #(
		.INIT('h9600)
	) name140 (
		_w1067_,
		_w1068_,
		_w1069_,
		_w1142_,
		_w1143_
	);
	LUT4 #(
		.INIT('h0069)
	) name141 (
		_w1067_,
		_w1068_,
		_w1069_,
		_w1142_,
		_w1144_
	);
	LUT3 #(
		.INIT('h69)
	) name142 (
		_w1126_,
		_w1127_,
		_w1128_,
		_w1145_
	);
	LUT3 #(
		.INIT('h45)
	) name143 (
		_w1143_,
		_w1144_,
		_w1145_,
		_w1146_
	);
	LUT3 #(
		.INIT('h71)
	) name144 (
		_w1139_,
		_w1141_,
		_w1146_,
		_w1147_
	);
	LUT3 #(
		.INIT('h45)
	) name145 (
		_w1137_,
		_w1138_,
		_w1147_,
		_w1148_
	);
	LUT3 #(
		.INIT('h17)
	) name146 (
		\A[3] ,
		\A[4] ,
		\A[5] ,
		_w1149_
	);
	LUT3 #(
		.INIT('h17)
	) name147 (
		\A[0] ,
		\A[1] ,
		\A[2] ,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w1149_,
		_w1150_,
		_w1151_
	);
	LUT3 #(
		.INIT('h96)
	) name149 (
		\A[0] ,
		\A[1] ,
		\A[2] ,
		_w1152_
	);
	LUT4 #(
		.INIT('h6996)
	) name150 (
		\A[0] ,
		\A[1] ,
		\A[2] ,
		\A[6] ,
		_w1153_
	);
	LUT3 #(
		.INIT('h96)
	) name151 (
		\A[3] ,
		\A[4] ,
		\A[5] ,
		_w1154_
	);
	LUT3 #(
		.INIT('h17)
	) name152 (
		\A[6] ,
		_w1152_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w1149_,
		_w1150_,
		_w1156_
	);
	LUT2 #(
		.INIT('h6)
	) name154 (
		_w1149_,
		_w1150_,
		_w1157_
	);
	LUT3 #(
		.INIT('h54)
	) name155 (
		_w1151_,
		_w1155_,
		_w1156_,
		_w1158_
	);
	LUT3 #(
		.INIT('h96)
	) name156 (
		\A[997] ,
		\A[998] ,
		\A[999] ,
		_w1159_
	);
	LUT3 #(
		.INIT('h60)
	) name157 (
		_w1153_,
		_w1154_,
		_w1159_,
		_w1160_
	);
	LUT3 #(
		.INIT('h17)
	) name158 (
		\A[997] ,
		\A[998] ,
		\A[999] ,
		_w1161_
	);
	LUT4 #(
		.INIT('h90f9)
	) name159 (
		_w1155_,
		_w1157_,
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w1158_,
		_w1162_,
		_w1163_
	);
	LUT3 #(
		.INIT('h96)
	) name161 (
		_w1153_,
		_w1154_,
		_w1159_,
		_w1164_
	);
	LUT3 #(
		.INIT('h96)
	) name162 (
		\A[991] ,
		\A[992] ,
		\A[993] ,
		_w1165_
	);
	LUT3 #(
		.INIT('h96)
	) name163 (
		\A[994] ,
		\A[995] ,
		\A[996] ,
		_w1166_
	);
	LUT2 #(
		.INIT('h6)
	) name164 (
		_w1165_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w1164_,
		_w1167_,
		_w1168_
	);
	LUT4 #(
		.INIT('h6996)
	) name166 (
		_w1155_,
		_w1157_,
		_w1160_,
		_w1161_,
		_w1169_
	);
	LUT3 #(
		.INIT('h17)
	) name167 (
		\A[994] ,
		\A[995] ,
		\A[996] ,
		_w1170_
	);
	LUT3 #(
		.INIT('h17)
	) name168 (
		\A[991] ,
		\A[992] ,
		\A[993] ,
		_w1171_
	);
	LUT4 #(
		.INIT('h7887)
	) name169 (
		_w1165_,
		_w1166_,
		_w1170_,
		_w1171_,
		_w1172_
	);
	LUT3 #(
		.INIT('h8e)
	) name170 (
		_w1168_,
		_w1169_,
		_w1172_,
		_w1173_
	);
	LUT4 #(
		.INIT('h088f)
	) name171 (
		_w1165_,
		_w1166_,
		_w1170_,
		_w1171_,
		_w1174_
	);
	LUT4 #(
		.INIT('h8e00)
	) name172 (
		_w1168_,
		_w1169_,
		_w1172_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w1163_,
		_w1175_,
		_w1176_
	);
	LUT3 #(
		.INIT('h96)
	) name174 (
		\A[19] ,
		\A[20] ,
		\A[21] ,
		_w1177_
	);
	LUT3 #(
		.INIT('h96)
	) name175 (
		\A[22] ,
		\A[23] ,
		\A[24] ,
		_w1178_
	);
	LUT3 #(
		.INIT('h96)
	) name176 (
		\A[25] ,
		\A[26] ,
		\A[27] ,
		_w1179_
	);
	LUT3 #(
		.INIT('h96)
	) name177 (
		\A[28] ,
		\A[29] ,
		\A[30] ,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w1179_,
		_w1180_,
		_w1181_
	);
	LUT4 #(
		.INIT('h0660)
	) name179 (
		_w1177_,
		_w1178_,
		_w1179_,
		_w1180_,
		_w1182_
	);
	LUT3 #(
		.INIT('h17)
	) name180 (
		\A[28] ,
		\A[29] ,
		\A[30] ,
		_w1183_
	);
	LUT3 #(
		.INIT('h17)
	) name181 (
		\A[25] ,
		\A[26] ,
		\A[27] ,
		_w1184_
	);
	LUT2 #(
		.INIT('h6)
	) name182 (
		_w1183_,
		_w1184_,
		_w1185_
	);
	LUT3 #(
		.INIT('h17)
	) name183 (
		\A[22] ,
		\A[23] ,
		\A[24] ,
		_w1186_
	);
	LUT3 #(
		.INIT('h17)
	) name184 (
		\A[19] ,
		\A[20] ,
		\A[21] ,
		_w1187_
	);
	LUT4 #(
		.INIT('h7887)
	) name185 (
		_w1177_,
		_w1178_,
		_w1186_,
		_w1187_,
		_w1188_
	);
	LUT4 #(
		.INIT('hc0de)
	) name186 (
		_w1181_,
		_w1182_,
		_w1185_,
		_w1188_,
		_w1189_
	);
	LUT4 #(
		.INIT('hf770)
	) name187 (
		_w1179_,
		_w1180_,
		_w1183_,
		_w1184_,
		_w1190_
	);
	LUT4 #(
		.INIT('h088f)
	) name188 (
		_w1177_,
		_w1178_,
		_w1186_,
		_w1187_,
		_w1191_
	);
	LUT3 #(
		.INIT('hb2)
	) name189 (
		_w1189_,
		_w1190_,
		_w1191_,
		_w1192_
	);
	LUT3 #(
		.INIT('h96)
	) name190 (
		\A[7] ,
		\A[8] ,
		\A[9] ,
		_w1193_
	);
	LUT3 #(
		.INIT('h96)
	) name191 (
		\A[10] ,
		\A[11] ,
		\A[12] ,
		_w1194_
	);
	LUT3 #(
		.INIT('h96)
	) name192 (
		\A[13] ,
		\A[14] ,
		\A[15] ,
		_w1195_
	);
	LUT3 #(
		.INIT('h96)
	) name193 (
		\A[16] ,
		\A[17] ,
		\A[18] ,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w1195_,
		_w1196_,
		_w1197_
	);
	LUT4 #(
		.INIT('h0660)
	) name195 (
		_w1193_,
		_w1194_,
		_w1195_,
		_w1196_,
		_w1198_
	);
	LUT3 #(
		.INIT('h17)
	) name196 (
		\A[16] ,
		\A[17] ,
		\A[18] ,
		_w1199_
	);
	LUT3 #(
		.INIT('h17)
	) name197 (
		\A[13] ,
		\A[14] ,
		\A[15] ,
		_w1200_
	);
	LUT2 #(
		.INIT('h6)
	) name198 (
		_w1199_,
		_w1200_,
		_w1201_
	);
	LUT3 #(
		.INIT('h17)
	) name199 (
		\A[10] ,
		\A[11] ,
		\A[12] ,
		_w1202_
	);
	LUT3 #(
		.INIT('h17)
	) name200 (
		\A[7] ,
		\A[8] ,
		\A[9] ,
		_w1203_
	);
	LUT4 #(
		.INIT('h7887)
	) name201 (
		_w1193_,
		_w1194_,
		_w1202_,
		_w1203_,
		_w1204_
	);
	LUT4 #(
		.INIT('hc0de)
	) name202 (
		_w1197_,
		_w1198_,
		_w1201_,
		_w1204_,
		_w1205_
	);
	LUT4 #(
		.INIT('hf770)
	) name203 (
		_w1195_,
		_w1196_,
		_w1199_,
		_w1200_,
		_w1206_
	);
	LUT4 #(
		.INIT('h088f)
	) name204 (
		_w1193_,
		_w1194_,
		_w1202_,
		_w1203_,
		_w1207_
	);
	LUT3 #(
		.INIT('hb2)
	) name205 (
		_w1205_,
		_w1206_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w1192_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w1192_,
		_w1208_,
		_w1210_
	);
	LUT3 #(
		.INIT('h96)
	) name208 (
		_w1205_,
		_w1206_,
		_w1207_,
		_w1211_
	);
	LUT3 #(
		.INIT('h96)
	) name209 (
		_w1189_,
		_w1190_,
		_w1191_,
		_w1212_
	);
	LUT4 #(
		.INIT('h6996)
	) name210 (
		_w1177_,
		_w1178_,
		_w1179_,
		_w1180_,
		_w1213_
	);
	LUT4 #(
		.INIT('h6996)
	) name211 (
		_w1193_,
		_w1194_,
		_w1195_,
		_w1196_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w1213_,
		_w1214_,
		_w1215_
	);
	LUT4 #(
		.INIT('he11e)
	) name213 (
		_w1181_,
		_w1182_,
		_w1185_,
		_w1188_,
		_w1216_
	);
	LUT4 #(
		.INIT('he11e)
	) name214 (
		_w1197_,
		_w1198_,
		_w1201_,
		_w1204_,
		_w1217_
	);
	LUT3 #(
		.INIT('hd4)
	) name215 (
		_w1215_,
		_w1216_,
		_w1217_,
		_w1218_
	);
	LUT3 #(
		.INIT('he8)
	) name216 (
		_w1211_,
		_w1212_,
		_w1218_,
		_w1219_
	);
	LUT4 #(
		.INIT('h80a8)
	) name217 (
		_w1176_,
		_w1192_,
		_w1208_,
		_w1219_,
		_w1220_
	);
	LUT4 #(
		.INIT('h1501)
	) name218 (
		_w1176_,
		_w1192_,
		_w1208_,
		_w1219_,
		_w1221_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		_w1158_,
		_w1162_,
		_w1222_
	);
	LUT4 #(
		.INIT('h9581)
	) name220 (
		_w1163_,
		_w1173_,
		_w1174_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h6)
	) name221 (
		_w1192_,
		_w1208_,
		_w1224_
	);
	LUT2 #(
		.INIT('h9)
	) name222 (
		_w1219_,
		_w1224_,
		_w1225_
	);
	LUT3 #(
		.INIT('h48)
	) name223 (
		_w1219_,
		_w1223_,
		_w1224_,
		_w1226_
	);
	LUT3 #(
		.INIT('h21)
	) name224 (
		_w1219_,
		_w1223_,
		_w1224_,
		_w1227_
	);
	LUT3 #(
		.INIT('h96)
	) name225 (
		_w1158_,
		_w1162_,
		_w1174_,
		_w1228_
	);
	LUT2 #(
		.INIT('h6)
	) name226 (
		_w1173_,
		_w1228_,
		_w1229_
	);
	LUT3 #(
		.INIT('h69)
	) name227 (
		_w1211_,
		_w1212_,
		_w1218_,
		_w1230_
	);
	LUT4 #(
		.INIT('h0660)
	) name228 (
		_w1164_,
		_w1167_,
		_w1213_,
		_w1214_,
		_w1231_
	);
	LUT4 #(
		.INIT('h9600)
	) name229 (
		_w1215_,
		_w1216_,
		_w1217_,
		_w1231_,
		_w1232_
	);
	LUT4 #(
		.INIT('h0069)
	) name230 (
		_w1215_,
		_w1216_,
		_w1217_,
		_w1231_,
		_w1233_
	);
	LUT3 #(
		.INIT('h96)
	) name231 (
		_w1168_,
		_w1169_,
		_w1172_,
		_w1234_
	);
	LUT3 #(
		.INIT('h54)
	) name232 (
		_w1232_,
		_w1233_,
		_w1234_,
		_w1235_
	);
	LUT3 #(
		.INIT('hb2)
	) name233 (
		_w1229_,
		_w1230_,
		_w1235_,
		_w1236_
	);
	LUT4 #(
		.INIT('h1051)
	) name234 (
		_w1221_,
		_w1223_,
		_w1225_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w1220_,
		_w1237_,
		_w1238_
	);
	LUT4 #(
		.INIT('h4d00)
	) name236 (
		_w1072_,
		_w1131_,
		_w1148_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('h00b2)
	) name237 (
		_w1072_,
		_w1131_,
		_w1148_,
		_w1238_,
		_w1240_
	);
	LUT4 #(
		.INIT('hba45)
	) name238 (
		_w1132_,
		_w1133_,
		_w1148_,
		_w1238_,
		_w1241_
	);
	LUT2 #(
		.INIT('h9)
	) name239 (
		_w1072_,
		_w1131_,
		_w1242_
	);
	LUT4 #(
		.INIT('h6665)
	) name240 (
		_w1176_,
		_w1209_,
		_w1210_,
		_w1219_,
		_w1243_
	);
	LUT4 #(
		.INIT('h45ba)
	) name241 (
		_w1226_,
		_w1227_,
		_w1236_,
		_w1243_,
		_w1244_
	);
	LUT3 #(
		.INIT('h06)
	) name242 (
		_w1148_,
		_w1242_,
		_w1244_,
		_w1245_
	);
	LUT3 #(
		.INIT('h90)
	) name243 (
		_w1148_,
		_w1242_,
		_w1244_,
		_w1246_
	);
	LUT3 #(
		.INIT('h96)
	) name244 (
		_w1071_,
		_w1134_,
		_w1136_,
		_w1247_
	);
	LUT3 #(
		.INIT('h96)
	) name245 (
		_w1219_,
		_w1223_,
		_w1224_,
		_w1248_
	);
	LUT2 #(
		.INIT('h6)
	) name246 (
		_w1236_,
		_w1248_,
		_w1249_
	);
	LUT3 #(
		.INIT('h09)
	) name247 (
		_w1147_,
		_w1247_,
		_w1249_,
		_w1250_
	);
	LUT3 #(
		.INIT('h60)
	) name248 (
		_w1147_,
		_w1247_,
		_w1249_,
		_w1251_
	);
	LUT3 #(
		.INIT('h96)
	) name249 (
		_w1229_,
		_w1230_,
		_w1235_,
		_w1252_
	);
	LUT4 #(
		.INIT('h0096)
	) name250 (
		_w1139_,
		_w1141_,
		_w1146_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('h6900)
	) name251 (
		_w1139_,
		_w1141_,
		_w1146_,
		_w1252_,
		_w1254_
	);
	LUT4 #(
		.INIT('h6996)
	) name252 (
		_w1164_,
		_w1167_,
		_w1213_,
		_w1214_,
		_w1255_
	);
	LUT4 #(
		.INIT('h6996)
	) name253 (
		_w1065_,
		_w1066_,
		_w1124_,
		_w1125_,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT4 #(
		.INIT('h6996)
	) name255 (
		_w1067_,
		_w1068_,
		_w1069_,
		_w1142_,
		_w1258_
	);
	LUT4 #(
		.INIT('h6996)
	) name256 (
		_w1215_,
		_w1216_,
		_w1217_,
		_w1231_,
		_w1259_
	);
	LUT2 #(
		.INIT('h9)
	) name257 (
		_w1234_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h21b7)
	) name258 (
		_w1145_,
		_w1257_,
		_w1258_,
		_w1260_,
		_w1261_
	);
	LUT3 #(
		.INIT('h45)
	) name259 (
		_w1253_,
		_w1254_,
		_w1261_,
		_w1262_
	);
	LUT3 #(
		.INIT('h45)
	) name260 (
		_w1250_,
		_w1251_,
		_w1262_,
		_w1263_
	);
	LUT4 #(
		.INIT('h6665)
	) name261 (
		_w1241_,
		_w1245_,
		_w1246_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\A[946] ,
		\A[947] ,
		_w1265_
	);
	LUT3 #(
		.INIT('h96)
	) name263 (
		\A[943] ,
		\A[944] ,
		\A[945] ,
		_w1266_
	);
	LUT3 #(
		.INIT('h96)
	) name264 (
		\A[946] ,
		\A[947] ,
		\A[948] ,
		_w1267_
	);
	LUT3 #(
		.INIT('h80)
	) name265 (
		_w1265_,
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT3 #(
		.INIT('h17)
	) name266 (
		\A[943] ,
		\A[944] ,
		\A[945] ,
		_w1269_
	);
	LUT3 #(
		.INIT('h17)
	) name267 (
		\A[946] ,
		\A[947] ,
		\A[948] ,
		_w1270_
	);
	LUT4 #(
		.INIT('h080f)
	) name268 (
		_w1266_,
		_w1267_,
		_w1269_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w1268_,
		_w1271_,
		_w1272_
	);
	LUT3 #(
		.INIT('h17)
	) name270 (
		\A[952] ,
		\A[953] ,
		\A[954] ,
		_w1273_
	);
	LUT3 #(
		.INIT('h17)
	) name271 (
		\A[949] ,
		\A[950] ,
		\A[951] ,
		_w1274_
	);
	LUT3 #(
		.INIT('h96)
	) name272 (
		\A[949] ,
		\A[950] ,
		\A[951] ,
		_w1275_
	);
	LUT3 #(
		.INIT('h96)
	) name273 (
		\A[952] ,
		\A[953] ,
		\A[954] ,
		_w1276_
	);
	LUT4 #(
		.INIT('h7111)
	) name274 (
		_w1273_,
		_w1274_,
		_w1275_,
		_w1276_,
		_w1277_
	);
	LUT4 #(
		.INIT('h0660)
	) name275 (
		_w1266_,
		_w1267_,
		_w1275_,
		_w1276_,
		_w1278_
	);
	LUT4 #(
		.INIT('h0080)
	) name276 (
		_w1265_,
		_w1266_,
		_w1267_,
		_w1269_,
		_w1279_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		_w1278_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('h6999)
	) name278 (
		_w1273_,
		_w1274_,
		_w1275_,
		_w1276_,
		_w1281_
	);
	LUT3 #(
		.INIT('h02)
	) name279 (
		_w1278_,
		_w1279_,
		_w1281_,
		_w1282_
	);
	LUT3 #(
		.INIT('hd0)
	) name280 (
		_w1278_,
		_w1279_,
		_w1281_,
		_w1283_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name281 (
		\A[946] ,
		\A[947] ,
		\A[948] ,
		_w1266_,
		_w1284_
	);
	LUT2 #(
		.INIT('h9)
	) name282 (
		_w1269_,
		_w1284_,
		_w1285_
	);
	LUT4 #(
		.INIT('h8a08)
	) name283 (
		_w1277_,
		_w1280_,
		_w1281_,
		_w1285_,
		_w1286_
	);
	LUT4 #(
		.INIT('h1051)
	) name284 (
		_w1277_,
		_w1280_,
		_w1281_,
		_w1285_,
		_w1287_
	);
	LUT4 #(
		.INIT('h6566)
	) name285 (
		_w1277_,
		_w1282_,
		_w1283_,
		_w1285_,
		_w1288_
	);
	LUT2 #(
		.INIT('h6)
	) name286 (
		_w1272_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\A[958] ,
		\A[959] ,
		_w1290_
	);
	LUT3 #(
		.INIT('h96)
	) name288 (
		\A[955] ,
		\A[956] ,
		\A[957] ,
		_w1291_
	);
	LUT3 #(
		.INIT('h96)
	) name289 (
		\A[958] ,
		\A[959] ,
		\A[960] ,
		_w1292_
	);
	LUT3 #(
		.INIT('h80)
	) name290 (
		_w1290_,
		_w1291_,
		_w1292_,
		_w1293_
	);
	LUT3 #(
		.INIT('h17)
	) name291 (
		\A[955] ,
		\A[956] ,
		\A[957] ,
		_w1294_
	);
	LUT3 #(
		.INIT('h17)
	) name292 (
		\A[958] ,
		\A[959] ,
		\A[960] ,
		_w1295_
	);
	LUT4 #(
		.INIT('h080f)
	) name293 (
		_w1291_,
		_w1292_,
		_w1294_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w1293_,
		_w1296_,
		_w1297_
	);
	LUT3 #(
		.INIT('h17)
	) name295 (
		\A[964] ,
		\A[965] ,
		\A[966] ,
		_w1298_
	);
	LUT3 #(
		.INIT('h17)
	) name296 (
		\A[961] ,
		\A[962] ,
		\A[963] ,
		_w1299_
	);
	LUT3 #(
		.INIT('h96)
	) name297 (
		\A[961] ,
		\A[962] ,
		\A[963] ,
		_w1300_
	);
	LUT3 #(
		.INIT('h96)
	) name298 (
		\A[964] ,
		\A[965] ,
		\A[966] ,
		_w1301_
	);
	LUT4 #(
		.INIT('h7111)
	) name299 (
		_w1298_,
		_w1299_,
		_w1300_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('h0660)
	) name300 (
		_w1291_,
		_w1292_,
		_w1300_,
		_w1301_,
		_w1303_
	);
	LUT4 #(
		.INIT('h0080)
	) name301 (
		_w1290_,
		_w1291_,
		_w1292_,
		_w1294_,
		_w1304_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		_w1303_,
		_w1304_,
		_w1305_
	);
	LUT4 #(
		.INIT('h6999)
	) name303 (
		_w1298_,
		_w1299_,
		_w1300_,
		_w1301_,
		_w1306_
	);
	LUT3 #(
		.INIT('h02)
	) name304 (
		_w1303_,
		_w1304_,
		_w1306_,
		_w1307_
	);
	LUT3 #(
		.INIT('hd0)
	) name305 (
		_w1303_,
		_w1304_,
		_w1306_,
		_w1308_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name306 (
		\A[958] ,
		\A[959] ,
		\A[960] ,
		_w1291_,
		_w1309_
	);
	LUT2 #(
		.INIT('h9)
	) name307 (
		_w1294_,
		_w1309_,
		_w1310_
	);
	LUT4 #(
		.INIT('h8a08)
	) name308 (
		_w1302_,
		_w1305_,
		_w1306_,
		_w1310_,
		_w1311_
	);
	LUT4 #(
		.INIT('h1051)
	) name309 (
		_w1302_,
		_w1305_,
		_w1306_,
		_w1310_,
		_w1312_
	);
	LUT4 #(
		.INIT('h6566)
	) name310 (
		_w1302_,
		_w1307_,
		_w1308_,
		_w1310_,
		_w1313_
	);
	LUT2 #(
		.INIT('h6)
	) name311 (
		_w1297_,
		_w1313_,
		_w1314_
	);
	LUT4 #(
		.INIT('h9009)
	) name312 (
		_w1272_,
		_w1288_,
		_w1297_,
		_w1313_,
		_w1315_
	);
	LUT4 #(
		.INIT('h0660)
	) name313 (
		_w1272_,
		_w1288_,
		_w1297_,
		_w1313_,
		_w1316_
	);
	LUT4 #(
		.INIT('h6996)
	) name314 (
		_w1291_,
		_w1292_,
		_w1300_,
		_w1301_,
		_w1317_
	);
	LUT4 #(
		.INIT('h6996)
	) name315 (
		_w1266_,
		_w1267_,
		_w1275_,
		_w1276_,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT3 #(
		.INIT('h2d)
	) name317 (
		_w1303_,
		_w1304_,
		_w1306_,
		_w1320_
	);
	LUT3 #(
		.INIT('h48)
	) name318 (
		_w1310_,
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT3 #(
		.INIT('h21)
	) name319 (
		_w1310_,
		_w1319_,
		_w1320_,
		_w1322_
	);
	LUT3 #(
		.INIT('h2d)
	) name320 (
		_w1278_,
		_w1279_,
		_w1281_,
		_w1323_
	);
	LUT2 #(
		.INIT('h6)
	) name321 (
		_w1285_,
		_w1323_,
		_w1324_
	);
	LUT3 #(
		.INIT('h45)
	) name322 (
		_w1321_,
		_w1322_,
		_w1324_,
		_w1325_
	);
	LUT3 #(
		.INIT('h54)
	) name323 (
		_w1315_,
		_w1316_,
		_w1325_,
		_w1326_
	);
	LUT3 #(
		.INIT('h32)
	) name324 (
		_w1297_,
		_w1311_,
		_w1312_,
		_w1327_
	);
	LUT4 #(
		.INIT('h0017)
	) name325 (
		_w1289_,
		_w1314_,
		_w1325_,
		_w1327_,
		_w1328_
	);
	LUT4 #(
		.INIT('he800)
	) name326 (
		_w1289_,
		_w1314_,
		_w1325_,
		_w1327_,
		_w1329_
	);
	LUT3 #(
		.INIT('h32)
	) name327 (
		_w1272_,
		_w1286_,
		_w1287_,
		_w1330_
	);
	LUT3 #(
		.INIT('h96)
	) name328 (
		\A[979] ,
		\A[980] ,
		\A[981] ,
		_w1331_
	);
	LUT3 #(
		.INIT('h96)
	) name329 (
		\A[982] ,
		\A[983] ,
		\A[984] ,
		_w1332_
	);
	LUT3 #(
		.INIT('h96)
	) name330 (
		\A[985] ,
		\A[986] ,
		\A[987] ,
		_w1333_
	);
	LUT3 #(
		.INIT('h96)
	) name331 (
		\A[988] ,
		\A[989] ,
		\A[990] ,
		_w1334_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT4 #(
		.INIT('h0660)
	) name333 (
		_w1331_,
		_w1332_,
		_w1333_,
		_w1334_,
		_w1336_
	);
	LUT3 #(
		.INIT('h17)
	) name334 (
		\A[988] ,
		\A[989] ,
		\A[990] ,
		_w1337_
	);
	LUT3 #(
		.INIT('h17)
	) name335 (
		\A[985] ,
		\A[986] ,
		\A[987] ,
		_w1338_
	);
	LUT2 #(
		.INIT('h6)
	) name336 (
		_w1337_,
		_w1338_,
		_w1339_
	);
	LUT3 #(
		.INIT('h17)
	) name337 (
		\A[982] ,
		\A[983] ,
		\A[984] ,
		_w1340_
	);
	LUT3 #(
		.INIT('h17)
	) name338 (
		\A[979] ,
		\A[980] ,
		\A[981] ,
		_w1341_
	);
	LUT4 #(
		.INIT('h7887)
	) name339 (
		_w1331_,
		_w1332_,
		_w1340_,
		_w1341_,
		_w1342_
	);
	LUT4 #(
		.INIT('hc0de)
	) name340 (
		_w1335_,
		_w1336_,
		_w1339_,
		_w1342_,
		_w1343_
	);
	LUT4 #(
		.INIT('hf770)
	) name341 (
		_w1333_,
		_w1334_,
		_w1337_,
		_w1338_,
		_w1344_
	);
	LUT4 #(
		.INIT('h088f)
	) name342 (
		_w1331_,
		_w1332_,
		_w1340_,
		_w1341_,
		_w1345_
	);
	LUT3 #(
		.INIT('hb2)
	) name343 (
		_w1343_,
		_w1344_,
		_w1345_,
		_w1346_
	);
	LUT3 #(
		.INIT('h96)
	) name344 (
		\A[967] ,
		\A[968] ,
		\A[969] ,
		_w1347_
	);
	LUT3 #(
		.INIT('h96)
	) name345 (
		\A[970] ,
		\A[971] ,
		\A[972] ,
		_w1348_
	);
	LUT3 #(
		.INIT('h96)
	) name346 (
		\A[973] ,
		\A[974] ,
		\A[975] ,
		_w1349_
	);
	LUT3 #(
		.INIT('h96)
	) name347 (
		\A[976] ,
		\A[977] ,
		\A[978] ,
		_w1350_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		_w1349_,
		_w1350_,
		_w1351_
	);
	LUT4 #(
		.INIT('h0660)
	) name349 (
		_w1347_,
		_w1348_,
		_w1349_,
		_w1350_,
		_w1352_
	);
	LUT3 #(
		.INIT('h17)
	) name350 (
		\A[976] ,
		\A[977] ,
		\A[978] ,
		_w1353_
	);
	LUT3 #(
		.INIT('h17)
	) name351 (
		\A[973] ,
		\A[974] ,
		\A[975] ,
		_w1354_
	);
	LUT2 #(
		.INIT('h6)
	) name352 (
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT3 #(
		.INIT('h17)
	) name353 (
		\A[970] ,
		\A[971] ,
		\A[972] ,
		_w1356_
	);
	LUT3 #(
		.INIT('h17)
	) name354 (
		\A[967] ,
		\A[968] ,
		\A[969] ,
		_w1357_
	);
	LUT4 #(
		.INIT('h7887)
	) name355 (
		_w1347_,
		_w1348_,
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('hc0de)
	) name356 (
		_w1351_,
		_w1352_,
		_w1355_,
		_w1358_,
		_w1359_
	);
	LUT4 #(
		.INIT('hf770)
	) name357 (
		_w1349_,
		_w1350_,
		_w1353_,
		_w1354_,
		_w1360_
	);
	LUT4 #(
		.INIT('h088f)
	) name358 (
		_w1347_,
		_w1348_,
		_w1356_,
		_w1357_,
		_w1361_
	);
	LUT3 #(
		.INIT('hb2)
	) name359 (
		_w1359_,
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		_w1346_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w1346_,
		_w1362_,
		_w1364_
	);
	LUT3 #(
		.INIT('h96)
	) name362 (
		_w1359_,
		_w1360_,
		_w1361_,
		_w1365_
	);
	LUT3 #(
		.INIT('h96)
	) name363 (
		_w1343_,
		_w1344_,
		_w1345_,
		_w1366_
	);
	LUT4 #(
		.INIT('h6996)
	) name364 (
		_w1331_,
		_w1332_,
		_w1333_,
		_w1334_,
		_w1367_
	);
	LUT4 #(
		.INIT('h6996)
	) name365 (
		_w1347_,
		_w1348_,
		_w1349_,
		_w1350_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		_w1367_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('he11e)
	) name367 (
		_w1335_,
		_w1336_,
		_w1339_,
		_w1342_,
		_w1370_
	);
	LUT4 #(
		.INIT('he11e)
	) name368 (
		_w1351_,
		_w1352_,
		_w1355_,
		_w1358_,
		_w1371_
	);
	LUT3 #(
		.INIT('hd4)
	) name369 (
		_w1369_,
		_w1370_,
		_w1371_,
		_w1372_
	);
	LUT3 #(
		.INIT('he8)
	) name370 (
		_w1365_,
		_w1366_,
		_w1372_,
		_w1373_
	);
	LUT3 #(
		.INIT('h54)
	) name371 (
		_w1363_,
		_w1364_,
		_w1373_,
		_w1374_
	);
	LUT4 #(
		.INIT('h0017)
	) name372 (
		_w1326_,
		_w1327_,
		_w1330_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('he800)
	) name373 (
		_w1326_,
		_w1327_,
		_w1330_,
		_w1374_,
		_w1376_
	);
	LUT4 #(
		.INIT('hab54)
	) name374 (
		_w1315_,
		_w1316_,
		_w1325_,
		_w1327_,
		_w1377_
	);
	LUT2 #(
		.INIT('h6)
	) name375 (
		_w1346_,
		_w1362_,
		_w1378_
	);
	LUT2 #(
		.INIT('h9)
	) name376 (
		_w1373_,
		_w1378_,
		_w1379_
	);
	LUT4 #(
		.INIT('h6996)
	) name377 (
		_w1272_,
		_w1288_,
		_w1297_,
		_w1313_,
		_w1380_
	);
	LUT3 #(
		.INIT('h69)
	) name378 (
		_w1365_,
		_w1366_,
		_w1372_,
		_w1381_
	);
	LUT4 #(
		.INIT('h0660)
	) name379 (
		_w1317_,
		_w1318_,
		_w1367_,
		_w1368_,
		_w1382_
	);
	LUT4 #(
		.INIT('h9600)
	) name380 (
		_w1369_,
		_w1370_,
		_w1371_,
		_w1382_,
		_w1383_
	);
	LUT4 #(
		.INIT('h0069)
	) name381 (
		_w1369_,
		_w1370_,
		_w1371_,
		_w1382_,
		_w1384_
	);
	LUT3 #(
		.INIT('h96)
	) name382 (
		_w1310_,
		_w1319_,
		_w1320_,
		_w1385_
	);
	LUT4 #(
		.INIT('h3231)
	) name383 (
		_w1324_,
		_w1383_,
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT4 #(
		.INIT('h6f06)
	) name384 (
		_w1325_,
		_w1380_,
		_w1381_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h6f06)
	) name385 (
		_w1330_,
		_w1377_,
		_w1379_,
		_w1387_,
		_w1388_
	);
	LUT3 #(
		.INIT('h54)
	) name386 (
		_w1375_,
		_w1376_,
		_w1388_,
		_w1389_
	);
	LUT4 #(
		.INIT('hab54)
	) name387 (
		_w1328_,
		_w1329_,
		_w1330_,
		_w1374_,
		_w1390_
	);
	LUT2 #(
		.INIT('h9)
	) name388 (
		_w1388_,
		_w1390_,
		_w1391_
	);
	LUT3 #(
		.INIT('h69)
	) name389 (
		_w1148_,
		_w1242_,
		_w1244_,
		_w1392_
	);
	LUT3 #(
		.INIT('h96)
	) name390 (
		_w1147_,
		_w1247_,
		_w1249_,
		_w1393_
	);
	LUT4 #(
		.INIT('h6996)
	) name391 (
		_w1330_,
		_w1377_,
		_w1379_,
		_w1387_,
		_w1394_
	);
	LUT4 #(
		.INIT('h6996)
	) name392 (
		_w1325_,
		_w1380_,
		_w1381_,
		_w1386_,
		_w1395_
	);
	LUT4 #(
		.INIT('h9669)
	) name393 (
		_w1139_,
		_w1141_,
		_w1146_,
		_w1252_,
		_w1396_
	);
	LUT4 #(
		.INIT('h6996)
	) name394 (
		_w1317_,
		_w1318_,
		_w1367_,
		_w1368_,
		_w1397_
	);
	LUT3 #(
		.INIT('h60)
	) name395 (
		_w1255_,
		_w1256_,
		_w1397_,
		_w1398_
	);
	LUT4 #(
		.INIT('h9669)
	) name396 (
		_w1145_,
		_w1257_,
		_w1258_,
		_w1260_,
		_w1399_
	);
	LUT4 #(
		.INIT('h6996)
	) name397 (
		_w1369_,
		_w1370_,
		_w1371_,
		_w1382_,
		_w1400_
	);
	LUT3 #(
		.INIT('h96)
	) name398 (
		_w1324_,
		_w1385_,
		_w1400_,
		_w1401_
	);
	LUT3 #(
		.INIT('h4d)
	) name399 (
		_w1398_,
		_w1399_,
		_w1401_,
		_w1402_
	);
	LUT4 #(
		.INIT('h84ed)
	) name400 (
		_w1261_,
		_w1395_,
		_w1396_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('hf660)
	) name401 (
		_w1262_,
		_w1393_,
		_w1394_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('hed84)
	) name402 (
		_w1263_,
		_w1391_,
		_w1392_,
		_w1404_,
		_w1405_
	);
	LUT3 #(
		.INIT('h4d)
	) name403 (
		_w1264_,
		_w1389_,
		_w1405_,
		_w1406_
	);
	LUT4 #(
		.INIT('h4445)
	) name404 (
		_w1239_,
		_w1245_,
		_w1246_,
		_w1263_,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w1240_,
		_w1407_,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w1406_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		\A[874] ,
		\A[875] ,
		_w1410_
	);
	LUT3 #(
		.INIT('h96)
	) name408 (
		\A[871] ,
		\A[872] ,
		\A[873] ,
		_w1411_
	);
	LUT3 #(
		.INIT('h96)
	) name409 (
		\A[874] ,
		\A[875] ,
		\A[876] ,
		_w1412_
	);
	LUT3 #(
		.INIT('h80)
	) name410 (
		_w1410_,
		_w1411_,
		_w1412_,
		_w1413_
	);
	LUT3 #(
		.INIT('h17)
	) name411 (
		\A[871] ,
		\A[872] ,
		\A[873] ,
		_w1414_
	);
	LUT3 #(
		.INIT('h17)
	) name412 (
		\A[874] ,
		\A[875] ,
		\A[876] ,
		_w1415_
	);
	LUT4 #(
		.INIT('h080f)
	) name413 (
		_w1411_,
		_w1412_,
		_w1414_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w1413_,
		_w1416_,
		_w1417_
	);
	LUT3 #(
		.INIT('h17)
	) name415 (
		\A[880] ,
		\A[881] ,
		\A[882] ,
		_w1418_
	);
	LUT3 #(
		.INIT('h17)
	) name416 (
		\A[877] ,
		\A[878] ,
		\A[879] ,
		_w1419_
	);
	LUT3 #(
		.INIT('h96)
	) name417 (
		\A[877] ,
		\A[878] ,
		\A[879] ,
		_w1420_
	);
	LUT3 #(
		.INIT('h96)
	) name418 (
		\A[880] ,
		\A[881] ,
		\A[882] ,
		_w1421_
	);
	LUT4 #(
		.INIT('h7111)
	) name419 (
		_w1418_,
		_w1419_,
		_w1420_,
		_w1421_,
		_w1422_
	);
	LUT4 #(
		.INIT('h0660)
	) name420 (
		_w1411_,
		_w1412_,
		_w1420_,
		_w1421_,
		_w1423_
	);
	LUT4 #(
		.INIT('h0080)
	) name421 (
		_w1410_,
		_w1411_,
		_w1412_,
		_w1414_,
		_w1424_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT4 #(
		.INIT('h6999)
	) name423 (
		_w1418_,
		_w1419_,
		_w1420_,
		_w1421_,
		_w1426_
	);
	LUT3 #(
		.INIT('h02)
	) name424 (
		_w1423_,
		_w1424_,
		_w1426_,
		_w1427_
	);
	LUT3 #(
		.INIT('hd0)
	) name425 (
		_w1423_,
		_w1424_,
		_w1426_,
		_w1428_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name426 (
		\A[874] ,
		\A[875] ,
		\A[876] ,
		_w1411_,
		_w1429_
	);
	LUT2 #(
		.INIT('h9)
	) name427 (
		_w1414_,
		_w1429_,
		_w1430_
	);
	LUT4 #(
		.INIT('h8a08)
	) name428 (
		_w1422_,
		_w1425_,
		_w1426_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('h1051)
	) name429 (
		_w1422_,
		_w1425_,
		_w1426_,
		_w1430_,
		_w1432_
	);
	LUT4 #(
		.INIT('h6566)
	) name430 (
		_w1422_,
		_w1427_,
		_w1428_,
		_w1430_,
		_w1433_
	);
	LUT2 #(
		.INIT('h6)
	) name431 (
		_w1417_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		\A[886] ,
		\A[887] ,
		_w1435_
	);
	LUT3 #(
		.INIT('h96)
	) name433 (
		\A[883] ,
		\A[884] ,
		\A[885] ,
		_w1436_
	);
	LUT3 #(
		.INIT('h96)
	) name434 (
		\A[886] ,
		\A[887] ,
		\A[888] ,
		_w1437_
	);
	LUT3 #(
		.INIT('h80)
	) name435 (
		_w1435_,
		_w1436_,
		_w1437_,
		_w1438_
	);
	LUT3 #(
		.INIT('h17)
	) name436 (
		\A[883] ,
		\A[884] ,
		\A[885] ,
		_w1439_
	);
	LUT3 #(
		.INIT('h17)
	) name437 (
		\A[886] ,
		\A[887] ,
		\A[888] ,
		_w1440_
	);
	LUT4 #(
		.INIT('h080f)
	) name438 (
		_w1436_,
		_w1437_,
		_w1439_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w1438_,
		_w1441_,
		_w1442_
	);
	LUT3 #(
		.INIT('h17)
	) name440 (
		\A[892] ,
		\A[893] ,
		\A[894] ,
		_w1443_
	);
	LUT3 #(
		.INIT('h17)
	) name441 (
		\A[889] ,
		\A[890] ,
		\A[891] ,
		_w1444_
	);
	LUT3 #(
		.INIT('h96)
	) name442 (
		\A[889] ,
		\A[890] ,
		\A[891] ,
		_w1445_
	);
	LUT3 #(
		.INIT('h96)
	) name443 (
		\A[892] ,
		\A[893] ,
		\A[894] ,
		_w1446_
	);
	LUT4 #(
		.INIT('h7111)
	) name444 (
		_w1443_,
		_w1444_,
		_w1445_,
		_w1446_,
		_w1447_
	);
	LUT4 #(
		.INIT('h0660)
	) name445 (
		_w1436_,
		_w1437_,
		_w1445_,
		_w1446_,
		_w1448_
	);
	LUT4 #(
		.INIT('h0080)
	) name446 (
		_w1435_,
		_w1436_,
		_w1437_,
		_w1439_,
		_w1449_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		_w1448_,
		_w1449_,
		_w1450_
	);
	LUT4 #(
		.INIT('h6999)
	) name448 (
		_w1443_,
		_w1444_,
		_w1445_,
		_w1446_,
		_w1451_
	);
	LUT3 #(
		.INIT('h02)
	) name449 (
		_w1448_,
		_w1449_,
		_w1451_,
		_w1452_
	);
	LUT3 #(
		.INIT('hd0)
	) name450 (
		_w1448_,
		_w1449_,
		_w1451_,
		_w1453_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name451 (
		\A[886] ,
		\A[887] ,
		\A[888] ,
		_w1436_,
		_w1454_
	);
	LUT2 #(
		.INIT('h9)
	) name452 (
		_w1439_,
		_w1454_,
		_w1455_
	);
	LUT4 #(
		.INIT('h8a08)
	) name453 (
		_w1447_,
		_w1450_,
		_w1451_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h1051)
	) name454 (
		_w1447_,
		_w1450_,
		_w1451_,
		_w1455_,
		_w1457_
	);
	LUT4 #(
		.INIT('h6566)
	) name455 (
		_w1447_,
		_w1452_,
		_w1453_,
		_w1455_,
		_w1458_
	);
	LUT2 #(
		.INIT('h6)
	) name456 (
		_w1442_,
		_w1458_,
		_w1459_
	);
	LUT4 #(
		.INIT('h9009)
	) name457 (
		_w1417_,
		_w1433_,
		_w1442_,
		_w1458_,
		_w1460_
	);
	LUT4 #(
		.INIT('h0660)
	) name458 (
		_w1417_,
		_w1433_,
		_w1442_,
		_w1458_,
		_w1461_
	);
	LUT4 #(
		.INIT('h6996)
	) name459 (
		_w1436_,
		_w1437_,
		_w1445_,
		_w1446_,
		_w1462_
	);
	LUT4 #(
		.INIT('h6996)
	) name460 (
		_w1411_,
		_w1412_,
		_w1420_,
		_w1421_,
		_w1463_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT3 #(
		.INIT('h2d)
	) name462 (
		_w1448_,
		_w1449_,
		_w1451_,
		_w1465_
	);
	LUT3 #(
		.INIT('h48)
	) name463 (
		_w1455_,
		_w1464_,
		_w1465_,
		_w1466_
	);
	LUT3 #(
		.INIT('h21)
	) name464 (
		_w1455_,
		_w1464_,
		_w1465_,
		_w1467_
	);
	LUT3 #(
		.INIT('h2d)
	) name465 (
		_w1423_,
		_w1424_,
		_w1426_,
		_w1468_
	);
	LUT2 #(
		.INIT('h6)
	) name466 (
		_w1430_,
		_w1468_,
		_w1469_
	);
	LUT3 #(
		.INIT('h45)
	) name467 (
		_w1466_,
		_w1467_,
		_w1469_,
		_w1470_
	);
	LUT3 #(
		.INIT('h32)
	) name468 (
		_w1442_,
		_w1456_,
		_w1457_,
		_w1471_
	);
	LUT4 #(
		.INIT('h0017)
	) name469 (
		_w1434_,
		_w1459_,
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT4 #(
		.INIT('he800)
	) name470 (
		_w1434_,
		_w1459_,
		_w1470_,
		_w1471_,
		_w1473_
	);
	LUT3 #(
		.INIT('h32)
	) name471 (
		_w1417_,
		_w1431_,
		_w1432_,
		_w1474_
	);
	LUT3 #(
		.INIT('h54)
	) name472 (
		_w1472_,
		_w1473_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('hab54)
	) name473 (
		_w1460_,
		_w1461_,
		_w1470_,
		_w1471_,
		_w1476_
	);
	LUT2 #(
		.INIT('h9)
	) name474 (
		_w1474_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		\A[850] ,
		\A[851] ,
		_w1478_
	);
	LUT3 #(
		.INIT('h96)
	) name476 (
		\A[847] ,
		\A[848] ,
		\A[849] ,
		_w1479_
	);
	LUT3 #(
		.INIT('h96)
	) name477 (
		\A[850] ,
		\A[851] ,
		\A[852] ,
		_w1480_
	);
	LUT3 #(
		.INIT('h80)
	) name478 (
		_w1478_,
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT3 #(
		.INIT('h17)
	) name479 (
		\A[847] ,
		\A[848] ,
		\A[849] ,
		_w1482_
	);
	LUT3 #(
		.INIT('h17)
	) name480 (
		\A[850] ,
		\A[851] ,
		\A[852] ,
		_w1483_
	);
	LUT4 #(
		.INIT('h080f)
	) name481 (
		_w1479_,
		_w1480_,
		_w1482_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w1481_,
		_w1484_,
		_w1485_
	);
	LUT3 #(
		.INIT('h17)
	) name483 (
		\A[856] ,
		\A[857] ,
		\A[858] ,
		_w1486_
	);
	LUT3 #(
		.INIT('h17)
	) name484 (
		\A[853] ,
		\A[854] ,
		\A[855] ,
		_w1487_
	);
	LUT3 #(
		.INIT('h96)
	) name485 (
		\A[853] ,
		\A[854] ,
		\A[855] ,
		_w1488_
	);
	LUT3 #(
		.INIT('h96)
	) name486 (
		\A[856] ,
		\A[857] ,
		\A[858] ,
		_w1489_
	);
	LUT4 #(
		.INIT('h7111)
	) name487 (
		_w1486_,
		_w1487_,
		_w1488_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('h0660)
	) name488 (
		_w1479_,
		_w1480_,
		_w1488_,
		_w1489_,
		_w1491_
	);
	LUT4 #(
		.INIT('h0080)
	) name489 (
		_w1478_,
		_w1479_,
		_w1480_,
		_w1482_,
		_w1492_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		_w1491_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('h6999)
	) name491 (
		_w1486_,
		_w1487_,
		_w1488_,
		_w1489_,
		_w1494_
	);
	LUT3 #(
		.INIT('h02)
	) name492 (
		_w1491_,
		_w1492_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('hd0)
	) name493 (
		_w1491_,
		_w1492_,
		_w1494_,
		_w1496_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name494 (
		\A[850] ,
		\A[851] ,
		\A[852] ,
		_w1479_,
		_w1497_
	);
	LUT2 #(
		.INIT('h9)
	) name495 (
		_w1482_,
		_w1497_,
		_w1498_
	);
	LUT4 #(
		.INIT('h8a08)
	) name496 (
		_w1490_,
		_w1493_,
		_w1494_,
		_w1498_,
		_w1499_
	);
	LUT4 #(
		.INIT('h1051)
	) name497 (
		_w1490_,
		_w1493_,
		_w1494_,
		_w1498_,
		_w1500_
	);
	LUT4 #(
		.INIT('h6566)
	) name498 (
		_w1490_,
		_w1495_,
		_w1496_,
		_w1498_,
		_w1501_
	);
	LUT2 #(
		.INIT('h6)
	) name499 (
		_w1485_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\A[862] ,
		\A[863] ,
		_w1503_
	);
	LUT3 #(
		.INIT('h96)
	) name501 (
		\A[859] ,
		\A[860] ,
		\A[861] ,
		_w1504_
	);
	LUT3 #(
		.INIT('h96)
	) name502 (
		\A[862] ,
		\A[863] ,
		\A[864] ,
		_w1505_
	);
	LUT3 #(
		.INIT('h80)
	) name503 (
		_w1503_,
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT3 #(
		.INIT('h17)
	) name504 (
		\A[859] ,
		\A[860] ,
		\A[861] ,
		_w1507_
	);
	LUT3 #(
		.INIT('h17)
	) name505 (
		\A[862] ,
		\A[863] ,
		\A[864] ,
		_w1508_
	);
	LUT4 #(
		.INIT('h080f)
	) name506 (
		_w1504_,
		_w1505_,
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w1506_,
		_w1509_,
		_w1510_
	);
	LUT3 #(
		.INIT('h17)
	) name508 (
		\A[868] ,
		\A[869] ,
		\A[870] ,
		_w1511_
	);
	LUT3 #(
		.INIT('h17)
	) name509 (
		\A[865] ,
		\A[866] ,
		\A[867] ,
		_w1512_
	);
	LUT3 #(
		.INIT('h96)
	) name510 (
		\A[865] ,
		\A[866] ,
		\A[867] ,
		_w1513_
	);
	LUT3 #(
		.INIT('h96)
	) name511 (
		\A[868] ,
		\A[869] ,
		\A[870] ,
		_w1514_
	);
	LUT4 #(
		.INIT('h7111)
	) name512 (
		_w1511_,
		_w1512_,
		_w1513_,
		_w1514_,
		_w1515_
	);
	LUT4 #(
		.INIT('h0660)
	) name513 (
		_w1504_,
		_w1505_,
		_w1513_,
		_w1514_,
		_w1516_
	);
	LUT4 #(
		.INIT('h0080)
	) name514 (
		_w1503_,
		_w1504_,
		_w1505_,
		_w1507_,
		_w1517_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		_w1516_,
		_w1517_,
		_w1518_
	);
	LUT4 #(
		.INIT('h6999)
	) name516 (
		_w1511_,
		_w1512_,
		_w1513_,
		_w1514_,
		_w1519_
	);
	LUT3 #(
		.INIT('h02)
	) name517 (
		_w1516_,
		_w1517_,
		_w1519_,
		_w1520_
	);
	LUT3 #(
		.INIT('hd0)
	) name518 (
		_w1516_,
		_w1517_,
		_w1519_,
		_w1521_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name519 (
		\A[862] ,
		\A[863] ,
		\A[864] ,
		_w1504_,
		_w1522_
	);
	LUT2 #(
		.INIT('h9)
	) name520 (
		_w1507_,
		_w1522_,
		_w1523_
	);
	LUT4 #(
		.INIT('h8a08)
	) name521 (
		_w1515_,
		_w1518_,
		_w1519_,
		_w1523_,
		_w1524_
	);
	LUT4 #(
		.INIT('h1051)
	) name522 (
		_w1515_,
		_w1518_,
		_w1519_,
		_w1523_,
		_w1525_
	);
	LUT4 #(
		.INIT('h6566)
	) name523 (
		_w1515_,
		_w1520_,
		_w1521_,
		_w1523_,
		_w1526_
	);
	LUT2 #(
		.INIT('h6)
	) name524 (
		_w1510_,
		_w1526_,
		_w1527_
	);
	LUT4 #(
		.INIT('h9009)
	) name525 (
		_w1485_,
		_w1501_,
		_w1510_,
		_w1526_,
		_w1528_
	);
	LUT4 #(
		.INIT('h0660)
	) name526 (
		_w1485_,
		_w1501_,
		_w1510_,
		_w1526_,
		_w1529_
	);
	LUT4 #(
		.INIT('h6996)
	) name527 (
		_w1504_,
		_w1505_,
		_w1513_,
		_w1514_,
		_w1530_
	);
	LUT4 #(
		.INIT('h6996)
	) name528 (
		_w1479_,
		_w1480_,
		_w1488_,
		_w1489_,
		_w1531_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT3 #(
		.INIT('h2d)
	) name530 (
		_w1516_,
		_w1517_,
		_w1519_,
		_w1533_
	);
	LUT3 #(
		.INIT('h48)
	) name531 (
		_w1523_,
		_w1532_,
		_w1533_,
		_w1534_
	);
	LUT3 #(
		.INIT('h21)
	) name532 (
		_w1523_,
		_w1532_,
		_w1533_,
		_w1535_
	);
	LUT3 #(
		.INIT('h2d)
	) name533 (
		_w1491_,
		_w1492_,
		_w1494_,
		_w1536_
	);
	LUT2 #(
		.INIT('h6)
	) name534 (
		_w1498_,
		_w1536_,
		_w1537_
	);
	LUT3 #(
		.INIT('h45)
	) name535 (
		_w1534_,
		_w1535_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('h32)
	) name536 (
		_w1510_,
		_w1524_,
		_w1525_,
		_w1539_
	);
	LUT4 #(
		.INIT('h0017)
	) name537 (
		_w1502_,
		_w1527_,
		_w1538_,
		_w1539_,
		_w1540_
	);
	LUT4 #(
		.INIT('he800)
	) name538 (
		_w1502_,
		_w1527_,
		_w1538_,
		_w1539_,
		_w1541_
	);
	LUT4 #(
		.INIT('hab54)
	) name539 (
		_w1528_,
		_w1529_,
		_w1538_,
		_w1539_,
		_w1542_
	);
	LUT3 #(
		.INIT('h32)
	) name540 (
		_w1485_,
		_w1499_,
		_w1500_,
		_w1543_
	);
	LUT2 #(
		.INIT('h9)
	) name541 (
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT4 #(
		.INIT('h0660)
	) name542 (
		_w1474_,
		_w1476_,
		_w1542_,
		_w1543_,
		_w1545_
	);
	LUT4 #(
		.INIT('h9009)
	) name543 (
		_w1474_,
		_w1476_,
		_w1542_,
		_w1543_,
		_w1546_
	);
	LUT4 #(
		.INIT('h6996)
	) name544 (
		_w1485_,
		_w1501_,
		_w1510_,
		_w1526_,
		_w1547_
	);
	LUT4 #(
		.INIT('h6996)
	) name545 (
		_w1417_,
		_w1433_,
		_w1442_,
		_w1458_,
		_w1548_
	);
	LUT4 #(
		.INIT('h1428)
	) name546 (
		_w1470_,
		_w1538_,
		_w1547_,
		_w1548_,
		_w1549_
	);
	LUT4 #(
		.INIT('h8241)
	) name547 (
		_w1470_,
		_w1538_,
		_w1547_,
		_w1548_,
		_w1550_
	);
	LUT4 #(
		.INIT('h0660)
	) name548 (
		_w1462_,
		_w1463_,
		_w1530_,
		_w1531_,
		_w1551_
	);
	LUT3 #(
		.INIT('h96)
	) name549 (
		_w1455_,
		_w1464_,
		_w1465_,
		_w1552_
	);
	LUT3 #(
		.INIT('h48)
	) name550 (
		_w1469_,
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT3 #(
		.INIT('h21)
	) name551 (
		_w1469_,
		_w1551_,
		_w1552_,
		_w1554_
	);
	LUT3 #(
		.INIT('h96)
	) name552 (
		_w1523_,
		_w1532_,
		_w1533_,
		_w1555_
	);
	LUT2 #(
		.INIT('h9)
	) name553 (
		_w1537_,
		_w1555_,
		_w1556_
	);
	LUT3 #(
		.INIT('h54)
	) name554 (
		_w1553_,
		_w1554_,
		_w1556_,
		_w1557_
	);
	LUT3 #(
		.INIT('h45)
	) name555 (
		_w1549_,
		_w1550_,
		_w1557_,
		_w1558_
	);
	LUT4 #(
		.INIT('h022a)
	) name556 (
		_w1475_,
		_w1477_,
		_w1544_,
		_w1558_,
		_w1559_
	);
	LUT4 #(
		.INIT('h5440)
	) name557 (
		_w1475_,
		_w1477_,
		_w1544_,
		_w1558_,
		_w1560_
	);
	LUT4 #(
		.INIT('h6665)
	) name558 (
		_w1475_,
		_w1545_,
		_w1546_,
		_w1558_,
		_w1561_
	);
	LUT3 #(
		.INIT('h54)
	) name559 (
		_w1540_,
		_w1541_,
		_w1543_,
		_w1562_
	);
	LUT2 #(
		.INIT('h6)
	) name560 (
		_w1561_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		\A[922] ,
		\A[923] ,
		_w1564_
	);
	LUT3 #(
		.INIT('h96)
	) name562 (
		\A[919] ,
		\A[920] ,
		\A[921] ,
		_w1565_
	);
	LUT3 #(
		.INIT('h96)
	) name563 (
		\A[922] ,
		\A[923] ,
		\A[924] ,
		_w1566_
	);
	LUT3 #(
		.INIT('h80)
	) name564 (
		_w1564_,
		_w1565_,
		_w1566_,
		_w1567_
	);
	LUT3 #(
		.INIT('h17)
	) name565 (
		\A[919] ,
		\A[920] ,
		\A[921] ,
		_w1568_
	);
	LUT3 #(
		.INIT('h17)
	) name566 (
		\A[922] ,
		\A[923] ,
		\A[924] ,
		_w1569_
	);
	LUT4 #(
		.INIT('h080f)
	) name567 (
		_w1565_,
		_w1566_,
		_w1568_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w1567_,
		_w1570_,
		_w1571_
	);
	LUT3 #(
		.INIT('h17)
	) name569 (
		\A[928] ,
		\A[929] ,
		\A[930] ,
		_w1572_
	);
	LUT3 #(
		.INIT('h17)
	) name570 (
		\A[925] ,
		\A[926] ,
		\A[927] ,
		_w1573_
	);
	LUT3 #(
		.INIT('h96)
	) name571 (
		\A[925] ,
		\A[926] ,
		\A[927] ,
		_w1574_
	);
	LUT3 #(
		.INIT('h96)
	) name572 (
		\A[928] ,
		\A[929] ,
		\A[930] ,
		_w1575_
	);
	LUT4 #(
		.INIT('h7111)
	) name573 (
		_w1572_,
		_w1573_,
		_w1574_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h0660)
	) name574 (
		_w1565_,
		_w1566_,
		_w1574_,
		_w1575_,
		_w1577_
	);
	LUT4 #(
		.INIT('h0080)
	) name575 (
		_w1564_,
		_w1565_,
		_w1566_,
		_w1568_,
		_w1578_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT4 #(
		.INIT('h6999)
	) name577 (
		_w1572_,
		_w1573_,
		_w1574_,
		_w1575_,
		_w1580_
	);
	LUT3 #(
		.INIT('h02)
	) name578 (
		_w1577_,
		_w1578_,
		_w1580_,
		_w1581_
	);
	LUT3 #(
		.INIT('hd0)
	) name579 (
		_w1577_,
		_w1578_,
		_w1580_,
		_w1582_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name580 (
		\A[922] ,
		\A[923] ,
		\A[924] ,
		_w1565_,
		_w1583_
	);
	LUT2 #(
		.INIT('h9)
	) name581 (
		_w1568_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('h8a08)
	) name582 (
		_w1576_,
		_w1579_,
		_w1580_,
		_w1584_,
		_w1585_
	);
	LUT4 #(
		.INIT('h1051)
	) name583 (
		_w1576_,
		_w1579_,
		_w1580_,
		_w1584_,
		_w1586_
	);
	LUT4 #(
		.INIT('h6566)
	) name584 (
		_w1576_,
		_w1581_,
		_w1582_,
		_w1584_,
		_w1587_
	);
	LUT2 #(
		.INIT('h6)
	) name585 (
		_w1571_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		\A[934] ,
		\A[935] ,
		_w1589_
	);
	LUT3 #(
		.INIT('h96)
	) name587 (
		\A[931] ,
		\A[932] ,
		\A[933] ,
		_w1590_
	);
	LUT3 #(
		.INIT('h96)
	) name588 (
		\A[934] ,
		\A[935] ,
		\A[936] ,
		_w1591_
	);
	LUT3 #(
		.INIT('h80)
	) name589 (
		_w1589_,
		_w1590_,
		_w1591_,
		_w1592_
	);
	LUT3 #(
		.INIT('h17)
	) name590 (
		\A[931] ,
		\A[932] ,
		\A[933] ,
		_w1593_
	);
	LUT3 #(
		.INIT('h17)
	) name591 (
		\A[934] ,
		\A[935] ,
		\A[936] ,
		_w1594_
	);
	LUT4 #(
		.INIT('h080f)
	) name592 (
		_w1590_,
		_w1591_,
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w1592_,
		_w1595_,
		_w1596_
	);
	LUT3 #(
		.INIT('h17)
	) name594 (
		\A[940] ,
		\A[941] ,
		\A[942] ,
		_w1597_
	);
	LUT3 #(
		.INIT('h17)
	) name595 (
		\A[937] ,
		\A[938] ,
		\A[939] ,
		_w1598_
	);
	LUT3 #(
		.INIT('h96)
	) name596 (
		\A[937] ,
		\A[938] ,
		\A[939] ,
		_w1599_
	);
	LUT3 #(
		.INIT('h96)
	) name597 (
		\A[940] ,
		\A[941] ,
		\A[942] ,
		_w1600_
	);
	LUT4 #(
		.INIT('h7111)
	) name598 (
		_w1597_,
		_w1598_,
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT4 #(
		.INIT('h0660)
	) name599 (
		_w1590_,
		_w1591_,
		_w1599_,
		_w1600_,
		_w1602_
	);
	LUT4 #(
		.INIT('h0080)
	) name600 (
		_w1589_,
		_w1590_,
		_w1591_,
		_w1593_,
		_w1603_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		_w1602_,
		_w1603_,
		_w1604_
	);
	LUT4 #(
		.INIT('h6999)
	) name602 (
		_w1597_,
		_w1598_,
		_w1599_,
		_w1600_,
		_w1605_
	);
	LUT3 #(
		.INIT('h02)
	) name603 (
		_w1602_,
		_w1603_,
		_w1605_,
		_w1606_
	);
	LUT3 #(
		.INIT('hd0)
	) name604 (
		_w1602_,
		_w1603_,
		_w1605_,
		_w1607_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name605 (
		\A[934] ,
		\A[935] ,
		\A[936] ,
		_w1590_,
		_w1608_
	);
	LUT2 #(
		.INIT('h9)
	) name606 (
		_w1593_,
		_w1608_,
		_w1609_
	);
	LUT4 #(
		.INIT('h8a08)
	) name607 (
		_w1601_,
		_w1604_,
		_w1605_,
		_w1609_,
		_w1610_
	);
	LUT4 #(
		.INIT('h1051)
	) name608 (
		_w1601_,
		_w1604_,
		_w1605_,
		_w1609_,
		_w1611_
	);
	LUT4 #(
		.INIT('h6566)
	) name609 (
		_w1601_,
		_w1606_,
		_w1607_,
		_w1609_,
		_w1612_
	);
	LUT2 #(
		.INIT('h6)
	) name610 (
		_w1596_,
		_w1612_,
		_w1613_
	);
	LUT4 #(
		.INIT('h9009)
	) name611 (
		_w1571_,
		_w1587_,
		_w1596_,
		_w1612_,
		_w1614_
	);
	LUT4 #(
		.INIT('h0660)
	) name612 (
		_w1571_,
		_w1587_,
		_w1596_,
		_w1612_,
		_w1615_
	);
	LUT4 #(
		.INIT('h6996)
	) name613 (
		_w1590_,
		_w1591_,
		_w1599_,
		_w1600_,
		_w1616_
	);
	LUT4 #(
		.INIT('h6996)
	) name614 (
		_w1565_,
		_w1566_,
		_w1574_,
		_w1575_,
		_w1617_
	);
	LUT2 #(
		.INIT('h8)
	) name615 (
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT3 #(
		.INIT('h2d)
	) name616 (
		_w1602_,
		_w1603_,
		_w1605_,
		_w1619_
	);
	LUT3 #(
		.INIT('h48)
	) name617 (
		_w1609_,
		_w1618_,
		_w1619_,
		_w1620_
	);
	LUT3 #(
		.INIT('h21)
	) name618 (
		_w1609_,
		_w1618_,
		_w1619_,
		_w1621_
	);
	LUT3 #(
		.INIT('h2d)
	) name619 (
		_w1577_,
		_w1578_,
		_w1580_,
		_w1622_
	);
	LUT2 #(
		.INIT('h6)
	) name620 (
		_w1584_,
		_w1622_,
		_w1623_
	);
	LUT3 #(
		.INIT('h45)
	) name621 (
		_w1620_,
		_w1621_,
		_w1623_,
		_w1624_
	);
	LUT3 #(
		.INIT('h32)
	) name622 (
		_w1596_,
		_w1610_,
		_w1611_,
		_w1625_
	);
	LUT4 #(
		.INIT('h0017)
	) name623 (
		_w1588_,
		_w1613_,
		_w1624_,
		_w1625_,
		_w1626_
	);
	LUT4 #(
		.INIT('he800)
	) name624 (
		_w1588_,
		_w1613_,
		_w1624_,
		_w1625_,
		_w1627_
	);
	LUT3 #(
		.INIT('h32)
	) name625 (
		_w1571_,
		_w1585_,
		_w1586_,
		_w1628_
	);
	LUT3 #(
		.INIT('h54)
	) name626 (
		_w1626_,
		_w1627_,
		_w1628_,
		_w1629_
	);
	LUT4 #(
		.INIT('hab54)
	) name627 (
		_w1614_,
		_w1615_,
		_w1624_,
		_w1625_,
		_w1630_
	);
	LUT2 #(
		.INIT('h9)
	) name628 (
		_w1628_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		\A[898] ,
		\A[899] ,
		_w1632_
	);
	LUT3 #(
		.INIT('h96)
	) name630 (
		\A[895] ,
		\A[896] ,
		\A[897] ,
		_w1633_
	);
	LUT3 #(
		.INIT('h96)
	) name631 (
		\A[898] ,
		\A[899] ,
		\A[900] ,
		_w1634_
	);
	LUT3 #(
		.INIT('h80)
	) name632 (
		_w1632_,
		_w1633_,
		_w1634_,
		_w1635_
	);
	LUT3 #(
		.INIT('h17)
	) name633 (
		\A[895] ,
		\A[896] ,
		\A[897] ,
		_w1636_
	);
	LUT3 #(
		.INIT('h17)
	) name634 (
		\A[898] ,
		\A[899] ,
		\A[900] ,
		_w1637_
	);
	LUT4 #(
		.INIT('h080f)
	) name635 (
		_w1633_,
		_w1634_,
		_w1636_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w1635_,
		_w1638_,
		_w1639_
	);
	LUT3 #(
		.INIT('h17)
	) name637 (
		\A[904] ,
		\A[905] ,
		\A[906] ,
		_w1640_
	);
	LUT3 #(
		.INIT('h17)
	) name638 (
		\A[901] ,
		\A[902] ,
		\A[903] ,
		_w1641_
	);
	LUT3 #(
		.INIT('h96)
	) name639 (
		\A[901] ,
		\A[902] ,
		\A[903] ,
		_w1642_
	);
	LUT3 #(
		.INIT('h96)
	) name640 (
		\A[904] ,
		\A[905] ,
		\A[906] ,
		_w1643_
	);
	LUT4 #(
		.INIT('h7111)
	) name641 (
		_w1640_,
		_w1641_,
		_w1642_,
		_w1643_,
		_w1644_
	);
	LUT4 #(
		.INIT('h0660)
	) name642 (
		_w1633_,
		_w1634_,
		_w1642_,
		_w1643_,
		_w1645_
	);
	LUT4 #(
		.INIT('h0080)
	) name643 (
		_w1632_,
		_w1633_,
		_w1634_,
		_w1636_,
		_w1646_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		_w1645_,
		_w1646_,
		_w1647_
	);
	LUT4 #(
		.INIT('h6999)
	) name645 (
		_w1640_,
		_w1641_,
		_w1642_,
		_w1643_,
		_w1648_
	);
	LUT3 #(
		.INIT('h02)
	) name646 (
		_w1645_,
		_w1646_,
		_w1648_,
		_w1649_
	);
	LUT3 #(
		.INIT('hd0)
	) name647 (
		_w1645_,
		_w1646_,
		_w1648_,
		_w1650_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name648 (
		\A[898] ,
		\A[899] ,
		\A[900] ,
		_w1633_,
		_w1651_
	);
	LUT2 #(
		.INIT('h9)
	) name649 (
		_w1636_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h8a08)
	) name650 (
		_w1644_,
		_w1647_,
		_w1648_,
		_w1652_,
		_w1653_
	);
	LUT4 #(
		.INIT('h1051)
	) name651 (
		_w1644_,
		_w1647_,
		_w1648_,
		_w1652_,
		_w1654_
	);
	LUT4 #(
		.INIT('h6566)
	) name652 (
		_w1644_,
		_w1649_,
		_w1650_,
		_w1652_,
		_w1655_
	);
	LUT2 #(
		.INIT('h6)
	) name653 (
		_w1639_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h8)
	) name654 (
		\A[910] ,
		\A[911] ,
		_w1657_
	);
	LUT3 #(
		.INIT('h96)
	) name655 (
		\A[907] ,
		\A[908] ,
		\A[909] ,
		_w1658_
	);
	LUT3 #(
		.INIT('h96)
	) name656 (
		\A[910] ,
		\A[911] ,
		\A[912] ,
		_w1659_
	);
	LUT3 #(
		.INIT('h80)
	) name657 (
		_w1657_,
		_w1658_,
		_w1659_,
		_w1660_
	);
	LUT3 #(
		.INIT('h17)
	) name658 (
		\A[907] ,
		\A[908] ,
		\A[909] ,
		_w1661_
	);
	LUT3 #(
		.INIT('h17)
	) name659 (
		\A[910] ,
		\A[911] ,
		\A[912] ,
		_w1662_
	);
	LUT4 #(
		.INIT('h080f)
	) name660 (
		_w1658_,
		_w1659_,
		_w1661_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w1660_,
		_w1663_,
		_w1664_
	);
	LUT3 #(
		.INIT('h17)
	) name662 (
		\A[916] ,
		\A[917] ,
		\A[918] ,
		_w1665_
	);
	LUT3 #(
		.INIT('h17)
	) name663 (
		\A[913] ,
		\A[914] ,
		\A[915] ,
		_w1666_
	);
	LUT3 #(
		.INIT('h96)
	) name664 (
		\A[913] ,
		\A[914] ,
		\A[915] ,
		_w1667_
	);
	LUT3 #(
		.INIT('h96)
	) name665 (
		\A[916] ,
		\A[917] ,
		\A[918] ,
		_w1668_
	);
	LUT4 #(
		.INIT('h7111)
	) name666 (
		_w1665_,
		_w1666_,
		_w1667_,
		_w1668_,
		_w1669_
	);
	LUT4 #(
		.INIT('h0660)
	) name667 (
		_w1658_,
		_w1659_,
		_w1667_,
		_w1668_,
		_w1670_
	);
	LUT4 #(
		.INIT('h0080)
	) name668 (
		_w1657_,
		_w1658_,
		_w1659_,
		_w1661_,
		_w1671_
	);
	LUT2 #(
		.INIT('h2)
	) name669 (
		_w1670_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('h6999)
	) name670 (
		_w1665_,
		_w1666_,
		_w1667_,
		_w1668_,
		_w1673_
	);
	LUT3 #(
		.INIT('h02)
	) name671 (
		_w1670_,
		_w1671_,
		_w1673_,
		_w1674_
	);
	LUT3 #(
		.INIT('hd0)
	) name672 (
		_w1670_,
		_w1671_,
		_w1673_,
		_w1675_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name673 (
		\A[910] ,
		\A[911] ,
		\A[912] ,
		_w1658_,
		_w1676_
	);
	LUT2 #(
		.INIT('h9)
	) name674 (
		_w1661_,
		_w1676_,
		_w1677_
	);
	LUT4 #(
		.INIT('h8a08)
	) name675 (
		_w1669_,
		_w1672_,
		_w1673_,
		_w1677_,
		_w1678_
	);
	LUT4 #(
		.INIT('h1051)
	) name676 (
		_w1669_,
		_w1672_,
		_w1673_,
		_w1677_,
		_w1679_
	);
	LUT4 #(
		.INIT('h6566)
	) name677 (
		_w1669_,
		_w1674_,
		_w1675_,
		_w1677_,
		_w1680_
	);
	LUT2 #(
		.INIT('h6)
	) name678 (
		_w1664_,
		_w1680_,
		_w1681_
	);
	LUT4 #(
		.INIT('h9009)
	) name679 (
		_w1639_,
		_w1655_,
		_w1664_,
		_w1680_,
		_w1682_
	);
	LUT4 #(
		.INIT('h0660)
	) name680 (
		_w1639_,
		_w1655_,
		_w1664_,
		_w1680_,
		_w1683_
	);
	LUT4 #(
		.INIT('h6996)
	) name681 (
		_w1658_,
		_w1659_,
		_w1667_,
		_w1668_,
		_w1684_
	);
	LUT4 #(
		.INIT('h6996)
	) name682 (
		_w1633_,
		_w1634_,
		_w1642_,
		_w1643_,
		_w1685_
	);
	LUT2 #(
		.INIT('h8)
	) name683 (
		_w1684_,
		_w1685_,
		_w1686_
	);
	LUT3 #(
		.INIT('h2d)
	) name684 (
		_w1670_,
		_w1671_,
		_w1673_,
		_w1687_
	);
	LUT3 #(
		.INIT('h48)
	) name685 (
		_w1677_,
		_w1686_,
		_w1687_,
		_w1688_
	);
	LUT3 #(
		.INIT('h21)
	) name686 (
		_w1677_,
		_w1686_,
		_w1687_,
		_w1689_
	);
	LUT3 #(
		.INIT('h2d)
	) name687 (
		_w1645_,
		_w1646_,
		_w1648_,
		_w1690_
	);
	LUT2 #(
		.INIT('h6)
	) name688 (
		_w1652_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h45)
	) name689 (
		_w1688_,
		_w1689_,
		_w1691_,
		_w1692_
	);
	LUT3 #(
		.INIT('h32)
	) name690 (
		_w1664_,
		_w1678_,
		_w1679_,
		_w1693_
	);
	LUT4 #(
		.INIT('h0017)
	) name691 (
		_w1656_,
		_w1681_,
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT4 #(
		.INIT('he800)
	) name692 (
		_w1656_,
		_w1681_,
		_w1692_,
		_w1693_,
		_w1695_
	);
	LUT4 #(
		.INIT('hab54)
	) name693 (
		_w1682_,
		_w1683_,
		_w1692_,
		_w1693_,
		_w1696_
	);
	LUT3 #(
		.INIT('h32)
	) name694 (
		_w1639_,
		_w1653_,
		_w1654_,
		_w1697_
	);
	LUT2 #(
		.INIT('h9)
	) name695 (
		_w1696_,
		_w1697_,
		_w1698_
	);
	LUT4 #(
		.INIT('h0660)
	) name696 (
		_w1628_,
		_w1630_,
		_w1696_,
		_w1697_,
		_w1699_
	);
	LUT4 #(
		.INIT('h9009)
	) name697 (
		_w1628_,
		_w1630_,
		_w1696_,
		_w1697_,
		_w1700_
	);
	LUT4 #(
		.INIT('h6996)
	) name698 (
		_w1639_,
		_w1655_,
		_w1664_,
		_w1680_,
		_w1701_
	);
	LUT4 #(
		.INIT('h6996)
	) name699 (
		_w1571_,
		_w1587_,
		_w1596_,
		_w1612_,
		_w1702_
	);
	LUT4 #(
		.INIT('h1428)
	) name700 (
		_w1624_,
		_w1692_,
		_w1701_,
		_w1702_,
		_w1703_
	);
	LUT4 #(
		.INIT('h8241)
	) name701 (
		_w1624_,
		_w1692_,
		_w1701_,
		_w1702_,
		_w1704_
	);
	LUT4 #(
		.INIT('h0660)
	) name702 (
		_w1616_,
		_w1617_,
		_w1684_,
		_w1685_,
		_w1705_
	);
	LUT3 #(
		.INIT('h96)
	) name703 (
		_w1609_,
		_w1618_,
		_w1619_,
		_w1706_
	);
	LUT3 #(
		.INIT('h48)
	) name704 (
		_w1623_,
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT3 #(
		.INIT('h21)
	) name705 (
		_w1623_,
		_w1705_,
		_w1706_,
		_w1708_
	);
	LUT3 #(
		.INIT('h96)
	) name706 (
		_w1677_,
		_w1686_,
		_w1687_,
		_w1709_
	);
	LUT2 #(
		.INIT('h9)
	) name707 (
		_w1691_,
		_w1709_,
		_w1710_
	);
	LUT3 #(
		.INIT('h54)
	) name708 (
		_w1707_,
		_w1708_,
		_w1710_,
		_w1711_
	);
	LUT3 #(
		.INIT('h45)
	) name709 (
		_w1703_,
		_w1704_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h022a)
	) name710 (
		_w1629_,
		_w1631_,
		_w1698_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('h5440)
	) name711 (
		_w1629_,
		_w1631_,
		_w1698_,
		_w1712_,
		_w1714_
	);
	LUT4 #(
		.INIT('h6665)
	) name712 (
		_w1629_,
		_w1699_,
		_w1700_,
		_w1712_,
		_w1715_
	);
	LUT3 #(
		.INIT('h54)
	) name713 (
		_w1694_,
		_w1695_,
		_w1697_,
		_w1716_
	);
	LUT2 #(
		.INIT('h6)
	) name714 (
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('h9009)
	) name715 (
		_w1561_,
		_w1562_,
		_w1715_,
		_w1716_,
		_w1718_
	);
	LUT4 #(
		.INIT('h0660)
	) name716 (
		_w1561_,
		_w1562_,
		_w1715_,
		_w1716_,
		_w1719_
	);
	LUT4 #(
		.INIT('h6996)
	) name717 (
		_w1628_,
		_w1630_,
		_w1696_,
		_w1697_,
		_w1720_
	);
	LUT4 #(
		.INIT('h6996)
	) name718 (
		_w1474_,
		_w1476_,
		_w1542_,
		_w1543_,
		_w1721_
	);
	LUT4 #(
		.INIT('h1428)
	) name719 (
		_w1558_,
		_w1712_,
		_w1720_,
		_w1721_,
		_w1722_
	);
	LUT4 #(
		.INIT('h8241)
	) name720 (
		_w1558_,
		_w1712_,
		_w1720_,
		_w1721_,
		_w1723_
	);
	LUT4 #(
		.INIT('h6996)
	) name721 (
		_w1470_,
		_w1538_,
		_w1547_,
		_w1548_,
		_w1724_
	);
	LUT4 #(
		.INIT('h6996)
	) name722 (
		_w1624_,
		_w1692_,
		_w1701_,
		_w1702_,
		_w1725_
	);
	LUT4 #(
		.INIT('h1248)
	) name723 (
		_w1557_,
		_w1711_,
		_w1724_,
		_w1725_,
		_w1726_
	);
	LUT4 #(
		.INIT('h8421)
	) name724 (
		_w1557_,
		_w1711_,
		_w1724_,
		_w1725_,
		_w1727_
	);
	LUT4 #(
		.INIT('h6996)
	) name725 (
		_w1616_,
		_w1617_,
		_w1684_,
		_w1685_,
		_w1728_
	);
	LUT4 #(
		.INIT('h6996)
	) name726 (
		_w1462_,
		_w1463_,
		_w1530_,
		_w1531_,
		_w1729_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		_w1728_,
		_w1729_,
		_w1730_
	);
	LUT3 #(
		.INIT('h96)
	) name728 (
		_w1623_,
		_w1705_,
		_w1706_,
		_w1731_
	);
	LUT3 #(
		.INIT('h84)
	) name729 (
		_w1710_,
		_w1730_,
		_w1731_,
		_w1732_
	);
	LUT3 #(
		.INIT('h12)
	) name730 (
		_w1710_,
		_w1730_,
		_w1731_,
		_w1733_
	);
	LUT3 #(
		.INIT('h96)
	) name731 (
		_w1469_,
		_w1551_,
		_w1552_,
		_w1734_
	);
	LUT2 #(
		.INIT('h9)
	) name732 (
		_w1556_,
		_w1734_,
		_w1735_
	);
	LUT3 #(
		.INIT('h45)
	) name733 (
		_w1732_,
		_w1733_,
		_w1735_,
		_w1736_
	);
	LUT3 #(
		.INIT('h45)
	) name734 (
		_w1726_,
		_w1727_,
		_w1736_,
		_w1737_
	);
	LUT3 #(
		.INIT('h45)
	) name735 (
		_w1722_,
		_w1723_,
		_w1737_,
		_w1738_
	);
	LUT3 #(
		.INIT('h45)
	) name736 (
		_w1713_,
		_w1714_,
		_w1716_,
		_w1739_
	);
	LUT4 #(
		.INIT('h00e8)
	) name737 (
		_w1563_,
		_w1717_,
		_w1738_,
		_w1739_,
		_w1740_
	);
	LUT4 #(
		.INIT('h1700)
	) name738 (
		_w1563_,
		_w1717_,
		_w1738_,
		_w1739_,
		_w1741_
	);
	LUT3 #(
		.INIT('h45)
	) name739 (
		_w1559_,
		_w1560_,
		_w1562_,
		_w1742_
	);
	LUT3 #(
		.INIT('h54)
	) name740 (
		_w1740_,
		_w1741_,
		_w1742_,
		_w1743_
	);
	LUT3 #(
		.INIT('h09)
	) name741 (
		_w1406_,
		_w1408_,
		_w1743_,
		_w1744_
	);
	LUT3 #(
		.INIT('h69)
	) name742 (
		_w1264_,
		_w1389_,
		_w1405_,
		_w1745_
	);
	LUT4 #(
		.INIT('h54ab)
	) name743 (
		_w1718_,
		_w1719_,
		_w1738_,
		_w1739_,
		_w1746_
	);
	LUT2 #(
		.INIT('h6)
	) name744 (
		_w1742_,
		_w1746_,
		_w1747_
	);
	LUT4 #(
		.INIT('h6996)
	) name745 (
		_w1561_,
		_w1562_,
		_w1715_,
		_w1716_,
		_w1748_
	);
	LUT2 #(
		.INIT('h9)
	) name746 (
		_w1738_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('h6996)
	) name747 (
		_w1263_,
		_w1391_,
		_w1392_,
		_w1404_,
		_w1750_
	);
	LUT4 #(
		.INIT('h9669)
	) name748 (
		_w1262_,
		_w1393_,
		_w1394_,
		_w1403_,
		_w1751_
	);
	LUT4 #(
		.INIT('h6996)
	) name749 (
		_w1558_,
		_w1712_,
		_w1720_,
		_w1721_,
		_w1752_
	);
	LUT2 #(
		.INIT('h6)
	) name750 (
		_w1737_,
		_w1752_,
		_w1753_
	);
	LUT4 #(
		.INIT('h6996)
	) name751 (
		_w1557_,
		_w1711_,
		_w1724_,
		_w1725_,
		_w1754_
	);
	LUT2 #(
		.INIT('h9)
	) name752 (
		_w1736_,
		_w1754_,
		_w1755_
	);
	LUT4 #(
		.INIT('h6996)
	) name753 (
		_w1261_,
		_w1395_,
		_w1396_,
		_w1402_,
		_w1756_
	);
	LUT2 #(
		.INIT('h6)
	) name754 (
		_w1728_,
		_w1729_,
		_w1757_
	);
	LUT3 #(
		.INIT('h96)
	) name755 (
		_w1255_,
		_w1256_,
		_w1397_,
		_w1758_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		_w1757_,
		_w1758_,
		_w1759_
	);
	LUT4 #(
		.INIT('h6900)
	) name757 (
		_w1398_,
		_w1399_,
		_w1401_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('h0096)
	) name758 (
		_w1398_,
		_w1399_,
		_w1401_,
		_w1759_,
		_w1761_
	);
	LUT3 #(
		.INIT('h69)
	) name759 (
		_w1710_,
		_w1730_,
		_w1731_,
		_w1762_
	);
	LUT2 #(
		.INIT('h9)
	) name760 (
		_w1735_,
		_w1762_,
		_w1763_
	);
	LUT3 #(
		.INIT('h54)
	) name761 (
		_w1760_,
		_w1761_,
		_w1763_,
		_w1764_
	);
	LUT3 #(
		.INIT('h8e)
	) name762 (
		_w1755_,
		_w1756_,
		_w1764_,
		_w1765_
	);
	LUT3 #(
		.INIT('hd4)
	) name763 (
		_w1751_,
		_w1753_,
		_w1765_,
		_w1766_
	);
	LUT3 #(
		.INIT('hb2)
	) name764 (
		_w1749_,
		_w1750_,
		_w1766_,
		_w1767_
	);
	LUT3 #(
		.INIT('he8)
	) name765 (
		_w1745_,
		_w1747_,
		_w1767_,
		_w1768_
	);
	LUT3 #(
		.INIT('h20)
	) name766 (
		_w1409_,
		_w1744_,
		_w1768_,
		_w1769_
	);
	LUT3 #(
		.INIT('h17)
	) name767 (
		\A[403] ,
		\A[404] ,
		\A[405] ,
		_w1770_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		\A[406] ,
		\A[407] ,
		_w1771_
	);
	LUT3 #(
		.INIT('h96)
	) name769 (
		\A[403] ,
		\A[404] ,
		\A[405] ,
		_w1772_
	);
	LUT3 #(
		.INIT('h96)
	) name770 (
		\A[406] ,
		\A[407] ,
		\A[408] ,
		_w1773_
	);
	LUT3 #(
		.INIT('h80)
	) name771 (
		_w1771_,
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT3 #(
		.INIT('h17)
	) name772 (
		\A[406] ,
		\A[407] ,
		\A[408] ,
		_w1775_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name773 (
		\A[406] ,
		\A[407] ,
		\A[408] ,
		_w1772_,
		_w1776_
	);
	LUT2 #(
		.INIT('h9)
	) name774 (
		_w1770_,
		_w1776_,
		_w1777_
	);
	LUT3 #(
		.INIT('h96)
	) name775 (
		\A[409] ,
		\A[410] ,
		\A[411] ,
		_w1778_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		\A[412] ,
		\A[413] ,
		_w1779_
	);
	LUT3 #(
		.INIT('h96)
	) name777 (
		\A[412] ,
		\A[413] ,
		\A[414] ,
		_w1780_
	);
	LUT3 #(
		.INIT('h17)
	) name778 (
		\A[412] ,
		\A[413] ,
		\A[414] ,
		_w1781_
	);
	LUT3 #(
		.INIT('h17)
	) name779 (
		\A[409] ,
		\A[410] ,
		\A[411] ,
		_w1782_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w1781_,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h6)
	) name781 (
		_w1781_,
		_w1782_,
		_w1784_
	);
	LUT4 #(
		.INIT('h8008)
	) name782 (
		_w1778_,
		_w1780_,
		_w1781_,
		_w1782_,
		_w1785_
	);
	LUT4 #(
		.INIT('h0770)
	) name783 (
		_w1778_,
		_w1780_,
		_w1781_,
		_w1782_,
		_w1786_
	);
	LUT4 #(
		.INIT('h0660)
	) name784 (
		_w1772_,
		_w1773_,
		_w1778_,
		_w1780_,
		_w1787_
	);
	LUT3 #(
		.INIT('h01)
	) name785 (
		_w1786_,
		_w1787_,
		_w1785_,
		_w1788_
	);
	LUT2 #(
		.INIT('h8)
	) name786 (
		_w1784_,
		_w1787_,
		_w1789_
	);
	LUT4 #(
		.INIT('h4000)
	) name787 (
		_w1770_,
		_w1771_,
		_w1772_,
		_w1773_,
		_w1790_
	);
	LUT3 #(
		.INIT('h08)
	) name788 (
		_w1784_,
		_w1787_,
		_w1790_,
		_w1791_
	);
	LUT4 #(
		.INIT('h80a0)
	) name789 (
		_w1778_,
		_w1779_,
		_w1780_,
		_w1782_,
		_w1792_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w1783_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h00f2)
	) name791 (
		_w1777_,
		_w1788_,
		_w1791_,
		_w1793_,
		_w1794_
	);
	LUT4 #(
		.INIT('h4055)
	) name792 (
		_w1770_,
		_w1772_,
		_w1773_,
		_w1775_,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w1774_,
		_w1795_,
		_w1796_
	);
	LUT4 #(
		.INIT('h0d00)
	) name794 (
		_w1777_,
		_w1788_,
		_w1791_,
		_w1793_,
		_w1797_
	);
	LUT3 #(
		.INIT('h54)
	) name795 (
		_w1794_,
		_w1796_,
		_w1797_,
		_w1798_
	);
	LUT3 #(
		.INIT('h96)
	) name796 (
		\A[397] ,
		\A[398] ,
		\A[399] ,
		_w1799_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		\A[400] ,
		\A[401] ,
		_w1800_
	);
	LUT3 #(
		.INIT('h96)
	) name798 (
		\A[400] ,
		\A[401] ,
		\A[402] ,
		_w1801_
	);
	LUT3 #(
		.INIT('h96)
	) name799 (
		\A[391] ,
		\A[392] ,
		\A[393] ,
		_w1802_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		\A[394] ,
		\A[395] ,
		_w1803_
	);
	LUT3 #(
		.INIT('h96)
	) name801 (
		\A[394] ,
		\A[395] ,
		\A[396] ,
		_w1804_
	);
	LUT4 #(
		.INIT('h0660)
	) name802 (
		_w1799_,
		_w1801_,
		_w1802_,
		_w1804_,
		_w1805_
	);
	LUT3 #(
		.INIT('h17)
	) name803 (
		\A[397] ,
		\A[398] ,
		\A[399] ,
		_w1806_
	);
	LUT3 #(
		.INIT('h17)
	) name804 (
		\A[400] ,
		\A[401] ,
		\A[402] ,
		_w1807_
	);
	LUT3 #(
		.INIT('h80)
	) name805 (
		_w1799_,
		_w1800_,
		_w1801_,
		_w1808_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name806 (
		\A[400] ,
		\A[401] ,
		\A[402] ,
		_w1799_,
		_w1809_
	);
	LUT2 #(
		.INIT('h9)
	) name807 (
		_w1806_,
		_w1809_,
		_w1810_
	);
	LUT3 #(
		.INIT('h14)
	) name808 (
		_w1805_,
		_w1806_,
		_w1809_,
		_w1811_
	);
	LUT3 #(
		.INIT('h17)
	) name809 (
		\A[391] ,
		\A[392] ,
		\A[393] ,
		_w1812_
	);
	LUT3 #(
		.INIT('h80)
	) name810 (
		_w1802_,
		_w1803_,
		_w1804_,
		_w1813_
	);
	LUT3 #(
		.INIT('h17)
	) name811 (
		\A[394] ,
		\A[395] ,
		\A[396] ,
		_w1814_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name812 (
		\A[394] ,
		\A[395] ,
		\A[396] ,
		_w1802_,
		_w1815_
	);
	LUT2 #(
		.INIT('h9)
	) name813 (
		_w1812_,
		_w1815_,
		_w1816_
	);
	LUT3 #(
		.INIT('h82)
	) name814 (
		_w1805_,
		_w1806_,
		_w1809_,
		_w1817_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w1806_,
		_w1807_,
		_w1818_
	);
	LUT4 #(
		.INIT('h0080)
	) name816 (
		_w1802_,
		_w1803_,
		_w1804_,
		_w1812_,
		_w1819_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w1818_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('h171f)
	) name818 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h080f)
	) name819 (
		_w1799_,
		_w1801_,
		_w1806_,
		_w1807_,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w1808_,
		_w1822_,
		_w1823_
	);
	LUT4 #(
		.INIT('h080f)
	) name821 (
		_w1802_,
		_w1804_,
		_w1812_,
		_w1814_,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w1813_,
		_w1824_,
		_w1825_
	);
	LUT3 #(
		.INIT('he8)
	) name823 (
		_w1821_,
		_w1823_,
		_w1825_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w1798_,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		_w1798_,
		_w1826_,
		_w1828_
	);
	LUT3 #(
		.INIT('h69)
	) name826 (
		_w1821_,
		_w1823_,
		_w1825_,
		_w1829_
	);
	LUT4 #(
		.INIT('hf20d)
	) name827 (
		_w1777_,
		_w1788_,
		_w1791_,
		_w1793_,
		_w1830_
	);
	LUT2 #(
		.INIT('h9)
	) name828 (
		_w1796_,
		_w1830_,
		_w1831_
	);
	LUT4 #(
		.INIT('h6996)
	) name829 (
		_w1772_,
		_w1773_,
		_w1778_,
		_w1780_,
		_w1832_
	);
	LUT4 #(
		.INIT('h6996)
	) name830 (
		_w1799_,
		_w1801_,
		_w1802_,
		_w1804_,
		_w1833_
	);
	LUT2 #(
		.INIT('h8)
	) name831 (
		_w1832_,
		_w1833_,
		_w1834_
	);
	LUT4 #(
		.INIT('h89a9)
	) name832 (
		_w1777_,
		_w1788_,
		_w1789_,
		_w1790_,
		_w1835_
	);
	LUT4 #(
		.INIT('hc989)
	) name833 (
		_w1811_,
		_w1816_,
		_w1817_,
		_w1820_,
		_w1836_
	);
	LUT3 #(
		.INIT('he8)
	) name834 (
		_w1834_,
		_w1835_,
		_w1836_,
		_w1837_
	);
	LUT3 #(
		.INIT('he8)
	) name835 (
		_w1829_,
		_w1831_,
		_w1837_,
		_w1838_
	);
	LUT3 #(
		.INIT('h45)
	) name836 (
		_w1827_,
		_w1828_,
		_w1838_,
		_w1839_
	);
	LUT3 #(
		.INIT('h96)
	) name837 (
		\A[385] ,
		\A[386] ,
		\A[387] ,
		_w1840_
	);
	LUT3 #(
		.INIT('h96)
	) name838 (
		\A[388] ,
		\A[389] ,
		\A[390] ,
		_w1841_
	);
	LUT2 #(
		.INIT('h8)
	) name839 (
		_w1840_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('h96)
	) name840 (
		\A[379] ,
		\A[380] ,
		\A[381] ,
		_w1843_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		\A[382] ,
		\A[383] ,
		_w1844_
	);
	LUT3 #(
		.INIT('h96)
	) name842 (
		\A[382] ,
		\A[383] ,
		\A[384] ,
		_w1845_
	);
	LUT4 #(
		.INIT('h0660)
	) name843 (
		_w1840_,
		_w1841_,
		_w1843_,
		_w1845_,
		_w1846_
	);
	LUT3 #(
		.INIT('h17)
	) name844 (
		\A[388] ,
		\A[389] ,
		\A[390] ,
		_w1847_
	);
	LUT3 #(
		.INIT('h17)
	) name845 (
		\A[385] ,
		\A[386] ,
		\A[387] ,
		_w1848_
	);
	LUT2 #(
		.INIT('h6)
	) name846 (
		_w1847_,
		_w1848_,
		_w1849_
	);
	LUT3 #(
		.INIT('h17)
	) name847 (
		\A[379] ,
		\A[380] ,
		\A[381] ,
		_w1850_
	);
	LUT3 #(
		.INIT('h17)
	) name848 (
		\A[382] ,
		\A[383] ,
		\A[384] ,
		_w1851_
	);
	LUT3 #(
		.INIT('h80)
	) name849 (
		_w1843_,
		_w1844_,
		_w1845_,
		_w1852_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name850 (
		\A[382] ,
		\A[383] ,
		\A[384] ,
		_w1843_,
		_w1853_
	);
	LUT2 #(
		.INIT('h9)
	) name851 (
		_w1850_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('h0770)
	) name852 (
		_w1846_,
		_w1849_,
		_w1850_,
		_w1853_,
		_w1855_
	);
	LUT4 #(
		.INIT('h8008)
	) name853 (
		_w1840_,
		_w1841_,
		_w1847_,
		_w1848_,
		_w1856_
	);
	LUT4 #(
		.INIT('h0770)
	) name854 (
		_w1840_,
		_w1841_,
		_w1847_,
		_w1848_,
		_w1857_
	);
	LUT3 #(
		.INIT('h01)
	) name855 (
		_w1846_,
		_w1857_,
		_w1856_,
		_w1858_
	);
	LUT4 #(
		.INIT('h088f)
	) name856 (
		_w1840_,
		_w1841_,
		_w1847_,
		_w1848_,
		_w1859_
	);
	LUT4 #(
		.INIT('h080f)
	) name857 (
		_w1843_,
		_w1845_,
		_w1850_,
		_w1851_,
		_w1860_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		_w1852_,
		_w1860_,
		_w1861_
	);
	LUT4 #(
		.INIT('h10f1)
	) name859 (
		_w1855_,
		_w1858_,
		_w1859_,
		_w1861_,
		_w1862_
	);
	LUT4 #(
		.INIT('he11e)
	) name860 (
		_w1855_,
		_w1858_,
		_w1859_,
		_w1861_,
		_w1863_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		\A[370] ,
		\A[371] ,
		_w1864_
	);
	LUT3 #(
		.INIT('h96)
	) name862 (
		\A[367] ,
		\A[368] ,
		\A[369] ,
		_w1865_
	);
	LUT3 #(
		.INIT('h96)
	) name863 (
		\A[370] ,
		\A[371] ,
		\A[372] ,
		_w1866_
	);
	LUT3 #(
		.INIT('h80)
	) name864 (
		_w1864_,
		_w1865_,
		_w1866_,
		_w1867_
	);
	LUT3 #(
		.INIT('h17)
	) name865 (
		\A[367] ,
		\A[368] ,
		\A[369] ,
		_w1868_
	);
	LUT3 #(
		.INIT('h17)
	) name866 (
		\A[370] ,
		\A[371] ,
		\A[372] ,
		_w1869_
	);
	LUT4 #(
		.INIT('h080f)
	) name867 (
		_w1865_,
		_w1866_,
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1867_,
		_w1870_,
		_w1871_
	);
	LUT3 #(
		.INIT('h96)
	) name869 (
		\A[373] ,
		\A[374] ,
		\A[375] ,
		_w1872_
	);
	LUT3 #(
		.INIT('h96)
	) name870 (
		\A[376] ,
		\A[377] ,
		\A[378] ,
		_w1873_
	);
	LUT2 #(
		.INIT('h8)
	) name871 (
		_w1872_,
		_w1873_,
		_w1874_
	);
	LUT4 #(
		.INIT('h0660)
	) name872 (
		_w1865_,
		_w1866_,
		_w1872_,
		_w1873_,
		_w1875_
	);
	LUT3 #(
		.INIT('h17)
	) name873 (
		\A[376] ,
		\A[377] ,
		\A[378] ,
		_w1876_
	);
	LUT3 #(
		.INIT('h17)
	) name874 (
		\A[373] ,
		\A[374] ,
		\A[375] ,
		_w1877_
	);
	LUT2 #(
		.INIT('h6)
	) name875 (
		_w1876_,
		_w1877_,
		_w1878_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name876 (
		\A[370] ,
		\A[371] ,
		\A[372] ,
		_w1865_,
		_w1879_
	);
	LUT2 #(
		.INIT('h9)
	) name877 (
		_w1868_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('h152a)
	) name878 (
		_w1868_,
		_w1875_,
		_w1878_,
		_w1879_,
		_w1881_
	);
	LUT4 #(
		.INIT('h8008)
	) name879 (
		_w1872_,
		_w1873_,
		_w1876_,
		_w1877_,
		_w1882_
	);
	LUT4 #(
		.INIT('h0770)
	) name880 (
		_w1872_,
		_w1873_,
		_w1876_,
		_w1877_,
		_w1883_
	);
	LUT3 #(
		.INIT('h01)
	) name881 (
		_w1875_,
		_w1883_,
		_w1882_,
		_w1884_
	);
	LUT4 #(
		.INIT('h088f)
	) name882 (
		_w1872_,
		_w1873_,
		_w1876_,
		_w1877_,
		_w1885_
	);
	LUT4 #(
		.INIT('ha956)
	) name883 (
		_w1871_,
		_w1881_,
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		_w1863_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w1863_,
		_w1886_,
		_w1888_
	);
	LUT4 #(
		.INIT('h6996)
	) name886 (
		_w1840_,
		_w1841_,
		_w1843_,
		_w1845_,
		_w1889_
	);
	LUT4 #(
		.INIT('h6996)
	) name887 (
		_w1865_,
		_w1866_,
		_w1872_,
		_w1873_,
		_w1890_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		_w1889_,
		_w1890_,
		_w1891_
	);
	LUT3 #(
		.INIT('h1e)
	) name889 (
		_w1842_,
		_w1846_,
		_w1849_,
		_w1892_
	);
	LUT3 #(
		.INIT('h48)
	) name890 (
		_w1854_,
		_w1891_,
		_w1892_,
		_w1893_
	);
	LUT3 #(
		.INIT('h21)
	) name891 (
		_w1854_,
		_w1891_,
		_w1892_,
		_w1894_
	);
	LUT3 #(
		.INIT('h1e)
	) name892 (
		_w1874_,
		_w1875_,
		_w1878_,
		_w1895_
	);
	LUT2 #(
		.INIT('h9)
	) name893 (
		_w1880_,
		_w1895_,
		_w1896_
	);
	LUT3 #(
		.INIT('h54)
	) name894 (
		_w1893_,
		_w1894_,
		_w1896_,
		_w1897_
	);
	LUT4 #(
		.INIT('h80a8)
	) name895 (
		_w1862_,
		_w1863_,
		_w1886_,
		_w1897_,
		_w1898_
	);
	LUT4 #(
		.INIT('h1501)
	) name896 (
		_w1862_,
		_w1863_,
		_w1886_,
		_w1897_,
		_w1899_
	);
	LUT4 #(
		.INIT('h5701)
	) name897 (
		_w1871_,
		_w1881_,
		_w1884_,
		_w1885_,
		_w1900_
	);
	LUT3 #(
		.INIT('h45)
	) name898 (
		_w1898_,
		_w1899_,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w1839_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		_w1839_,
		_w1901_,
		_w1903_
	);
	LUT2 #(
		.INIT('h6)
	) name901 (
		_w1798_,
		_w1826_,
		_w1904_
	);
	LUT4 #(
		.INIT('h6665)
	) name902 (
		_w1862_,
		_w1887_,
		_w1888_,
		_w1897_,
		_w1905_
	);
	LUT4 #(
		.INIT('h1248)
	) name903 (
		_w1838_,
		_w1900_,
		_w1904_,
		_w1905_,
		_w1906_
	);
	LUT4 #(
		.INIT('h8421)
	) name904 (
		_w1838_,
		_w1900_,
		_w1904_,
		_w1905_,
		_w1907_
	);
	LUT3 #(
		.INIT('h96)
	) name905 (
		_w1829_,
		_w1831_,
		_w1837_,
		_w1908_
	);
	LUT2 #(
		.INIT('h6)
	) name906 (
		_w1863_,
		_w1886_,
		_w1909_
	);
	LUT2 #(
		.INIT('h9)
	) name907 (
		_w1897_,
		_w1909_,
		_w1910_
	);
	LUT4 #(
		.INIT('h0660)
	) name908 (
		_w1832_,
		_w1833_,
		_w1889_,
		_w1890_,
		_w1911_
	);
	LUT4 #(
		.INIT('h9600)
	) name909 (
		_w1834_,
		_w1835_,
		_w1836_,
		_w1911_,
		_w1912_
	);
	LUT4 #(
		.INIT('h0069)
	) name910 (
		_w1834_,
		_w1835_,
		_w1836_,
		_w1911_,
		_w1913_
	);
	LUT3 #(
		.INIT('h96)
	) name911 (
		_w1854_,
		_w1891_,
		_w1892_,
		_w1914_
	);
	LUT2 #(
		.INIT('h9)
	) name912 (
		_w1896_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('h45)
	) name913 (
		_w1912_,
		_w1913_,
		_w1915_,
		_w1916_
	);
	LUT3 #(
		.INIT('h71)
	) name914 (
		_w1908_,
		_w1910_,
		_w1916_,
		_w1917_
	);
	LUT3 #(
		.INIT('h54)
	) name915 (
		_w1906_,
		_w1907_,
		_w1917_,
		_w1918_
	);
	LUT3 #(
		.INIT('h54)
	) name916 (
		_w1902_,
		_w1903_,
		_w1918_,
		_w1919_
	);
	LUT3 #(
		.INIT('h96)
	) name917 (
		\A[445] ,
		\A[446] ,
		\A[447] ,
		_w1920_
	);
	LUT2 #(
		.INIT('h8)
	) name918 (
		\A[448] ,
		\A[449] ,
		_w1921_
	);
	LUT3 #(
		.INIT('h96)
	) name919 (
		\A[448] ,
		\A[449] ,
		\A[450] ,
		_w1922_
	);
	LUT3 #(
		.INIT('h96)
	) name920 (
		\A[439] ,
		\A[440] ,
		\A[441] ,
		_w1923_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		\A[442] ,
		\A[443] ,
		_w1924_
	);
	LUT3 #(
		.INIT('h96)
	) name922 (
		\A[442] ,
		\A[443] ,
		\A[444] ,
		_w1925_
	);
	LUT4 #(
		.INIT('h0660)
	) name923 (
		_w1920_,
		_w1922_,
		_w1923_,
		_w1925_,
		_w1926_
	);
	LUT3 #(
		.INIT('h17)
	) name924 (
		\A[445] ,
		\A[446] ,
		\A[447] ,
		_w1927_
	);
	LUT3 #(
		.INIT('h17)
	) name925 (
		\A[448] ,
		\A[449] ,
		\A[450] ,
		_w1928_
	);
	LUT3 #(
		.INIT('h80)
	) name926 (
		_w1920_,
		_w1921_,
		_w1922_,
		_w1929_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name927 (
		\A[448] ,
		\A[449] ,
		\A[450] ,
		_w1920_,
		_w1930_
	);
	LUT2 #(
		.INIT('h9)
	) name928 (
		_w1927_,
		_w1930_,
		_w1931_
	);
	LUT3 #(
		.INIT('h14)
	) name929 (
		_w1926_,
		_w1927_,
		_w1930_,
		_w1932_
	);
	LUT3 #(
		.INIT('h17)
	) name930 (
		\A[439] ,
		\A[440] ,
		\A[441] ,
		_w1933_
	);
	LUT3 #(
		.INIT('h80)
	) name931 (
		_w1923_,
		_w1924_,
		_w1925_,
		_w1934_
	);
	LUT3 #(
		.INIT('h17)
	) name932 (
		\A[442] ,
		\A[443] ,
		\A[444] ,
		_w1935_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name933 (
		\A[442] ,
		\A[443] ,
		\A[444] ,
		_w1923_,
		_w1936_
	);
	LUT2 #(
		.INIT('h9)
	) name934 (
		_w1933_,
		_w1936_,
		_w1937_
	);
	LUT3 #(
		.INIT('h82)
	) name935 (
		_w1926_,
		_w1927_,
		_w1930_,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1927_,
		_w1928_,
		_w1939_
	);
	LUT4 #(
		.INIT('h0080)
	) name937 (
		_w1923_,
		_w1924_,
		_w1925_,
		_w1933_,
		_w1940_
	);
	LUT2 #(
		.INIT('h1)
	) name938 (
		_w1939_,
		_w1940_,
		_w1941_
	);
	LUT4 #(
		.INIT('h171f)
	) name939 (
		_w1926_,
		_w1931_,
		_w1937_,
		_w1941_,
		_w1942_
	);
	LUT4 #(
		.INIT('h080f)
	) name940 (
		_w1920_,
		_w1922_,
		_w1927_,
		_w1928_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name941 (
		_w1929_,
		_w1943_,
		_w1944_
	);
	LUT4 #(
		.INIT('h080f)
	) name942 (
		_w1923_,
		_w1925_,
		_w1933_,
		_w1935_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		_w1934_,
		_w1945_,
		_w1946_
	);
	LUT3 #(
		.INIT('h96)
	) name944 (
		\A[451] ,
		\A[452] ,
		\A[453] ,
		_w1947_
	);
	LUT3 #(
		.INIT('h96)
	) name945 (
		\A[454] ,
		\A[455] ,
		\A[456] ,
		_w1948_
	);
	LUT3 #(
		.INIT('h17)
	) name946 (
		\A[454] ,
		\A[455] ,
		\A[456] ,
		_w1949_
	);
	LUT3 #(
		.INIT('h17)
	) name947 (
		\A[451] ,
		\A[452] ,
		\A[453] ,
		_w1950_
	);
	LUT4 #(
		.INIT('h7887)
	) name948 (
		_w1947_,
		_w1948_,
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT3 #(
		.INIT('h96)
	) name949 (
		\A[457] ,
		\A[458] ,
		\A[459] ,
		_w1952_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		\A[460] ,
		\A[461] ,
		_w1953_
	);
	LUT3 #(
		.INIT('h96)
	) name951 (
		\A[460] ,
		\A[461] ,
		\A[462] ,
		_w1954_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		_w1952_,
		_w1954_,
		_w1955_
	);
	LUT3 #(
		.INIT('h17)
	) name953 (
		\A[460] ,
		\A[461] ,
		\A[462] ,
		_w1956_
	);
	LUT3 #(
		.INIT('h17)
	) name954 (
		\A[457] ,
		\A[458] ,
		\A[459] ,
		_w1957_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w1956_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h6)
	) name956 (
		_w1956_,
		_w1957_,
		_w1959_
	);
	LUT4 #(
		.INIT('h0660)
	) name957 (
		_w1947_,
		_w1948_,
		_w1952_,
		_w1954_,
		_w1960_
	);
	LUT4 #(
		.INIT('h5514)
	) name958 (
		_w1951_,
		_w1955_,
		_w1959_,
		_w1960_,
		_w1961_
	);
	LUT4 #(
		.INIT('h0008)
	) name959 (
		_w1947_,
		_w1948_,
		_w1949_,
		_w1950_,
		_w1962_
	);
	LUT3 #(
		.INIT('h08)
	) name960 (
		_w1959_,
		_w1960_,
		_w1962_,
		_w1963_
	);
	LUT4 #(
		.INIT('h80a0)
	) name961 (
		_w1952_,
		_w1953_,
		_w1954_,
		_w1957_,
		_w1964_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w1958_,
		_w1964_,
		_w1965_
	);
	LUT4 #(
		.INIT('h088f)
	) name963 (
		_w1947_,
		_w1948_,
		_w1949_,
		_w1950_,
		_w1966_
	);
	LUT4 #(
		.INIT('hef0e)
	) name964 (
		_w1961_,
		_w1963_,
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h1700)
	) name965 (
		_w1942_,
		_w1944_,
		_w1946_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('h00e8)
	) name966 (
		_w1942_,
		_w1944_,
		_w1946_,
		_w1967_,
		_w1969_
	);
	LUT3 #(
		.INIT('h69)
	) name967 (
		_w1942_,
		_w1944_,
		_w1946_,
		_w1970_
	);
	LUT4 #(
		.INIT('he11e)
	) name968 (
		_w1961_,
		_w1963_,
		_w1965_,
		_w1966_,
		_w1971_
	);
	LUT4 #(
		.INIT('h0069)
	) name969 (
		_w1942_,
		_w1944_,
		_w1946_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h9600)
	) name970 (
		_w1942_,
		_w1944_,
		_w1946_,
		_w1971_,
		_w1973_
	);
	LUT4 #(
		.INIT('h6996)
	) name971 (
		_w1947_,
		_w1948_,
		_w1952_,
		_w1954_,
		_w1974_
	);
	LUT4 #(
		.INIT('h6996)
	) name972 (
		_w1920_,
		_w1922_,
		_w1923_,
		_w1925_,
		_w1975_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		_w1974_,
		_w1975_,
		_w1976_
	);
	LUT4 #(
		.INIT('ha082)
	) name974 (
		_w1951_,
		_w1955_,
		_w1959_,
		_w1960_,
		_w1977_
	);
	LUT4 #(
		.INIT('h0f02)
	) name975 (
		_w1961_,
		_w1963_,
		_w1976_,
		_w1977_,
		_w1978_
	);
	LUT4 #(
		.INIT('hc989)
	) name976 (
		_w1932_,
		_w1937_,
		_w1938_,
		_w1941_,
		_w1979_
	);
	LUT4 #(
		.INIT('h00d0)
	) name977 (
		_w1961_,
		_w1963_,
		_w1976_,
		_w1977_,
		_w1980_
	);
	LUT3 #(
		.INIT('h54)
	) name978 (
		_w1978_,
		_w1979_,
		_w1980_,
		_w1981_
	);
	LUT4 #(
		.INIT('h4504)
	) name979 (
		_w1969_,
		_w1970_,
		_w1971_,
		_w1981_,
		_w1982_
	);
	LUT3 #(
		.INIT('h17)
	) name980 (
		\A[427] ,
		\A[428] ,
		\A[429] ,
		_w1983_
	);
	LUT2 #(
		.INIT('h8)
	) name981 (
		\A[430] ,
		\A[431] ,
		_w1984_
	);
	LUT3 #(
		.INIT('h96)
	) name982 (
		\A[427] ,
		\A[428] ,
		\A[429] ,
		_w1985_
	);
	LUT3 #(
		.INIT('h96)
	) name983 (
		\A[430] ,
		\A[431] ,
		\A[432] ,
		_w1986_
	);
	LUT3 #(
		.INIT('h80)
	) name984 (
		_w1984_,
		_w1985_,
		_w1986_,
		_w1987_
	);
	LUT3 #(
		.INIT('h17)
	) name985 (
		\A[430] ,
		\A[431] ,
		\A[432] ,
		_w1988_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name986 (
		\A[430] ,
		\A[431] ,
		\A[432] ,
		_w1985_,
		_w1989_
	);
	LUT2 #(
		.INIT('h9)
	) name987 (
		_w1983_,
		_w1989_,
		_w1990_
	);
	LUT3 #(
		.INIT('h96)
	) name988 (
		\A[433] ,
		\A[434] ,
		\A[435] ,
		_w1991_
	);
	LUT2 #(
		.INIT('h8)
	) name989 (
		\A[436] ,
		\A[437] ,
		_w1992_
	);
	LUT3 #(
		.INIT('h96)
	) name990 (
		\A[436] ,
		\A[437] ,
		\A[438] ,
		_w1993_
	);
	LUT3 #(
		.INIT('h17)
	) name991 (
		\A[436] ,
		\A[437] ,
		\A[438] ,
		_w1994_
	);
	LUT3 #(
		.INIT('h17)
	) name992 (
		\A[433] ,
		\A[434] ,
		\A[435] ,
		_w1995_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h6)
	) name994 (
		_w1994_,
		_w1995_,
		_w1997_
	);
	LUT4 #(
		.INIT('h8008)
	) name995 (
		_w1991_,
		_w1993_,
		_w1994_,
		_w1995_,
		_w1998_
	);
	LUT4 #(
		.INIT('h0770)
	) name996 (
		_w1991_,
		_w1993_,
		_w1994_,
		_w1995_,
		_w1999_
	);
	LUT4 #(
		.INIT('h0660)
	) name997 (
		_w1985_,
		_w1986_,
		_w1991_,
		_w1993_,
		_w2000_
	);
	LUT3 #(
		.INIT('h01)
	) name998 (
		_w1999_,
		_w2000_,
		_w1998_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name999 (
		_w1997_,
		_w2000_,
		_w2002_
	);
	LUT4 #(
		.INIT('h4000)
	) name1000 (
		_w1983_,
		_w1984_,
		_w1985_,
		_w1986_,
		_w2003_
	);
	LUT3 #(
		.INIT('h08)
	) name1001 (
		_w1997_,
		_w2000_,
		_w2003_,
		_w2004_
	);
	LUT3 #(
		.INIT('h0d)
	) name1002 (
		_w1990_,
		_w2001_,
		_w2004_,
		_w2005_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1003 (
		_w1991_,
		_w1992_,
		_w1993_,
		_w1995_,
		_w2006_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w1996_,
		_w2006_,
		_w2007_
	);
	LUT4 #(
		.INIT('h00f2)
	) name1005 (
		_w1990_,
		_w2001_,
		_w2004_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('h4055)
	) name1006 (
		_w1983_,
		_w1985_,
		_w1986_,
		_w1988_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		_w1987_,
		_w2009_,
		_w2010_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1008 (
		_w1990_,
		_w2001_,
		_w2004_,
		_w2007_,
		_w2011_
	);
	LUT3 #(
		.INIT('h96)
	) name1009 (
		\A[421] ,
		\A[422] ,
		\A[423] ,
		_w2012_
	);
	LUT3 #(
		.INIT('h96)
	) name1010 (
		\A[424] ,
		\A[425] ,
		\A[426] ,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1011 (
		_w2012_,
		_w2013_,
		_w2014_
	);
	LUT3 #(
		.INIT('h96)
	) name1012 (
		\A[415] ,
		\A[416] ,
		\A[417] ,
		_w2015_
	);
	LUT3 #(
		.INIT('h96)
	) name1013 (
		\A[418] ,
		\A[419] ,
		\A[420] ,
		_w2016_
	);
	LUT4 #(
		.INIT('h0660)
	) name1014 (
		_w2012_,
		_w2013_,
		_w2015_,
		_w2016_,
		_w2017_
	);
	LUT3 #(
		.INIT('h17)
	) name1015 (
		\A[424] ,
		\A[425] ,
		\A[426] ,
		_w2018_
	);
	LUT3 #(
		.INIT('h17)
	) name1016 (
		\A[421] ,
		\A[422] ,
		\A[423] ,
		_w2019_
	);
	LUT2 #(
		.INIT('h6)
	) name1017 (
		_w2018_,
		_w2019_,
		_w2020_
	);
	LUT3 #(
		.INIT('h17)
	) name1018 (
		\A[418] ,
		\A[419] ,
		\A[420] ,
		_w2021_
	);
	LUT3 #(
		.INIT('h17)
	) name1019 (
		\A[415] ,
		\A[416] ,
		\A[417] ,
		_w2022_
	);
	LUT4 #(
		.INIT('h7887)
	) name1020 (
		_w2015_,
		_w2016_,
		_w2021_,
		_w2022_,
		_w2023_
	);
	LUT4 #(
		.INIT('hc0de)
	) name1021 (
		_w2014_,
		_w2017_,
		_w2020_,
		_w2023_,
		_w2024_
	);
	LUT4 #(
		.INIT('h088f)
	) name1022 (
		_w2012_,
		_w2013_,
		_w2018_,
		_w2019_,
		_w2025_
	);
	LUT4 #(
		.INIT('h088f)
	) name1023 (
		_w2015_,
		_w2016_,
		_w2021_,
		_w2022_,
		_w2026_
	);
	LUT3 #(
		.INIT('he8)
	) name1024 (
		_w2024_,
		_w2025_,
		_w2026_,
		_w2027_
	);
	LUT4 #(
		.INIT('h1700)
	) name1025 (
		_w2005_,
		_w2007_,
		_w2010_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1026 (
		_w2005_,
		_w2007_,
		_w2010_,
		_w2027_,
		_w2029_
	);
	LUT4 #(
		.INIT('hf20d)
	) name1027 (
		_w1990_,
		_w2001_,
		_w2004_,
		_w2007_,
		_w2030_
	);
	LUT3 #(
		.INIT('h69)
	) name1028 (
		_w2024_,
		_w2025_,
		_w2026_,
		_w2031_
	);
	LUT3 #(
		.INIT('h09)
	) name1029 (
		_w2010_,
		_w2030_,
		_w2031_,
		_w2032_
	);
	LUT3 #(
		.INIT('h60)
	) name1030 (
		_w2010_,
		_w2030_,
		_w2031_,
		_w2033_
	);
	LUT4 #(
		.INIT('h6996)
	) name1031 (
		_w1985_,
		_w1986_,
		_w1991_,
		_w1993_,
		_w2034_
	);
	LUT4 #(
		.INIT('h6996)
	) name1032 (
		_w2012_,
		_w2013_,
		_w2015_,
		_w2016_,
		_w2035_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		_w2034_,
		_w2035_,
		_w2036_
	);
	LUT4 #(
		.INIT('h89a9)
	) name1034 (
		_w1990_,
		_w2001_,
		_w2002_,
		_w2003_,
		_w2037_
	);
	LUT4 #(
		.INIT('he11e)
	) name1035 (
		_w2014_,
		_w2017_,
		_w2020_,
		_w2023_,
		_w2038_
	);
	LUT3 #(
		.INIT('h71)
	) name1036 (
		_w2036_,
		_w2037_,
		_w2038_,
		_w2039_
	);
	LUT4 #(
		.INIT('h4445)
	) name1037 (
		_w2029_,
		_w2032_,
		_w2033_,
		_w2039_,
		_w2040_
	);
	LUT4 #(
		.INIT('heee0)
	) name1038 (
		_w1968_,
		_w1982_,
		_w2028_,
		_w2040_,
		_w2041_
	);
	LUT4 #(
		.INIT('h0001)
	) name1039 (
		_w1968_,
		_w1982_,
		_w2028_,
		_w2040_,
		_w2042_
	);
	LUT4 #(
		.INIT('he817)
	) name1040 (
		_w1942_,
		_w1944_,
		_w1946_,
		_w1967_,
		_w2043_
	);
	LUT4 #(
		.INIT('h45ba)
	) name1041 (
		_w1972_,
		_w1973_,
		_w1981_,
		_w2043_,
		_w2044_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1042 (
		_w2008_,
		_w2010_,
		_w2011_,
		_w2027_,
		_w2045_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1043 (
		_w2032_,
		_w2033_,
		_w2039_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		_w2044_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		_w2044_,
		_w2046_,
		_w2048_
	);
	LUT3 #(
		.INIT('h96)
	) name1046 (
		_w2010_,
		_w2030_,
		_w2031_,
		_w2049_
	);
	LUT4 #(
		.INIT('h6996)
	) name1047 (
		_w1942_,
		_w1944_,
		_w1946_,
		_w1971_,
		_w2050_
	);
	LUT4 #(
		.INIT('h4182)
	) name1048 (
		_w1981_,
		_w2039_,
		_w2049_,
		_w2050_,
		_w2051_
	);
	LUT4 #(
		.INIT('h2814)
	) name1049 (
		_w1981_,
		_w2039_,
		_w2049_,
		_w2050_,
		_w2052_
	);
	LUT4 #(
		.INIT('h0660)
	) name1050 (
		_w1974_,
		_w1975_,
		_w2034_,
		_w2035_,
		_w2053_
	);
	LUT4 #(
		.INIT('hf02d)
	) name1051 (
		_w1961_,
		_w1963_,
		_w1976_,
		_w1977_,
		_w2054_
	);
	LUT3 #(
		.INIT('h48)
	) name1052 (
		_w1979_,
		_w2053_,
		_w2054_,
		_w2055_
	);
	LUT3 #(
		.INIT('h21)
	) name1053 (
		_w1979_,
		_w2053_,
		_w2054_,
		_w2056_
	);
	LUT3 #(
		.INIT('h69)
	) name1054 (
		_w2036_,
		_w2037_,
		_w2038_,
		_w2057_
	);
	LUT3 #(
		.INIT('h45)
	) name1055 (
		_w2055_,
		_w2056_,
		_w2057_,
		_w2058_
	);
	LUT3 #(
		.INIT('h54)
	) name1056 (
		_w2051_,
		_w2052_,
		_w2058_,
		_w2059_
	);
	LUT4 #(
		.INIT('h4054)
	) name1057 (
		_w2042_,
		_w2044_,
		_w2046_,
		_w2059_,
		_w2060_
	);
	LUT2 #(
		.INIT('h1)
	) name1058 (
		_w2041_,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		_w1919_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		_w1919_,
		_w2061_,
		_w2063_
	);
	LUT4 #(
		.INIT('h111e)
	) name1061 (
		_w1968_,
		_w1982_,
		_w2028_,
		_w2040_,
		_w2064_
	);
	LUT4 #(
		.INIT('h45ba)
	) name1062 (
		_w2047_,
		_w2048_,
		_w2059_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h6)
	) name1063 (
		_w1839_,
		_w1901_,
		_w2066_
	);
	LUT3 #(
		.INIT('h48)
	) name1064 (
		_w1918_,
		_w2065_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('h21)
	) name1065 (
		_w1918_,
		_w2065_,
		_w2066_,
		_w2068_
	);
	LUT4 #(
		.INIT('h6996)
	) name1066 (
		_w1838_,
		_w1900_,
		_w1904_,
		_w1905_,
		_w2069_
	);
	LUT2 #(
		.INIT('h6)
	) name1067 (
		_w2044_,
		_w2046_,
		_w2070_
	);
	LUT4 #(
		.INIT('h1248)
	) name1068 (
		_w1917_,
		_w2059_,
		_w2069_,
		_w2070_,
		_w2071_
	);
	LUT4 #(
		.INIT('h8421)
	) name1069 (
		_w1917_,
		_w2059_,
		_w2069_,
		_w2070_,
		_w2072_
	);
	LUT3 #(
		.INIT('h69)
	) name1070 (
		_w1908_,
		_w1910_,
		_w1916_,
		_w2073_
	);
	LUT4 #(
		.INIT('h9669)
	) name1071 (
		_w1981_,
		_w2039_,
		_w2049_,
		_w2050_,
		_w2074_
	);
	LUT2 #(
		.INIT('h9)
	) name1072 (
		_w2058_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('h6996)
	) name1073 (
		_w1974_,
		_w1975_,
		_w2034_,
		_w2035_,
		_w2076_
	);
	LUT4 #(
		.INIT('h6996)
	) name1074 (
		_w1832_,
		_w1833_,
		_w1889_,
		_w1890_,
		_w2077_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT3 #(
		.INIT('h96)
	) name1076 (
		_w1979_,
		_w2053_,
		_w2054_,
		_w2079_
	);
	LUT3 #(
		.INIT('h48)
	) name1077 (
		_w2057_,
		_w2078_,
		_w2079_,
		_w2080_
	);
	LUT3 #(
		.INIT('h21)
	) name1078 (
		_w2057_,
		_w2078_,
		_w2079_,
		_w2081_
	);
	LUT4 #(
		.INIT('h6996)
	) name1079 (
		_w1834_,
		_w1835_,
		_w1836_,
		_w1911_,
		_w2082_
	);
	LUT2 #(
		.INIT('h9)
	) name1080 (
		_w1915_,
		_w2082_,
		_w2083_
	);
	LUT3 #(
		.INIT('h54)
	) name1081 (
		_w2080_,
		_w2081_,
		_w2083_,
		_w2084_
	);
	LUT3 #(
		.INIT('h8e)
	) name1082 (
		_w2073_,
		_w2075_,
		_w2084_,
		_w2085_
	);
	LUT3 #(
		.INIT('h54)
	) name1083 (
		_w2071_,
		_w2072_,
		_w2085_,
		_w2086_
	);
	LUT3 #(
		.INIT('h54)
	) name1084 (
		_w2067_,
		_w2068_,
		_w2086_,
		_w2087_
	);
	LUT3 #(
		.INIT('h45)
	) name1085 (
		_w2062_,
		_w2063_,
		_w2087_,
		_w2088_
	);
	LUT3 #(
		.INIT('h17)
	) name1086 (
		\A[355] ,
		\A[356] ,
		\A[357] ,
		_w2089_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		\A[358] ,
		\A[359] ,
		_w2090_
	);
	LUT3 #(
		.INIT('h96)
	) name1088 (
		\A[355] ,
		\A[356] ,
		\A[357] ,
		_w2091_
	);
	LUT3 #(
		.INIT('h96)
	) name1089 (
		\A[358] ,
		\A[359] ,
		\A[360] ,
		_w2092_
	);
	LUT3 #(
		.INIT('h80)
	) name1090 (
		_w2090_,
		_w2091_,
		_w2092_,
		_w2093_
	);
	LUT3 #(
		.INIT('h17)
	) name1091 (
		\A[358] ,
		\A[359] ,
		\A[360] ,
		_w2094_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1092 (
		\A[358] ,
		\A[359] ,
		\A[360] ,
		_w2091_,
		_w2095_
	);
	LUT2 #(
		.INIT('h9)
	) name1093 (
		_w2089_,
		_w2095_,
		_w2096_
	);
	LUT3 #(
		.INIT('h96)
	) name1094 (
		\A[361] ,
		\A[362] ,
		\A[363] ,
		_w2097_
	);
	LUT2 #(
		.INIT('h8)
	) name1095 (
		\A[364] ,
		\A[365] ,
		_w2098_
	);
	LUT3 #(
		.INIT('h96)
	) name1096 (
		\A[364] ,
		\A[365] ,
		\A[366] ,
		_w2099_
	);
	LUT3 #(
		.INIT('h17)
	) name1097 (
		\A[364] ,
		\A[365] ,
		\A[366] ,
		_w2100_
	);
	LUT3 #(
		.INIT('h17)
	) name1098 (
		\A[361] ,
		\A[362] ,
		\A[363] ,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h6)
	) name1100 (
		_w2100_,
		_w2101_,
		_w2103_
	);
	LUT4 #(
		.INIT('h8008)
	) name1101 (
		_w2097_,
		_w2099_,
		_w2100_,
		_w2101_,
		_w2104_
	);
	LUT4 #(
		.INIT('h0770)
	) name1102 (
		_w2097_,
		_w2099_,
		_w2100_,
		_w2101_,
		_w2105_
	);
	LUT4 #(
		.INIT('h0660)
	) name1103 (
		_w2091_,
		_w2092_,
		_w2097_,
		_w2099_,
		_w2106_
	);
	LUT3 #(
		.INIT('h01)
	) name1104 (
		_w2105_,
		_w2106_,
		_w2104_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		_w2103_,
		_w2106_,
		_w2108_
	);
	LUT4 #(
		.INIT('h4000)
	) name1106 (
		_w2089_,
		_w2090_,
		_w2091_,
		_w2092_,
		_w2109_
	);
	LUT3 #(
		.INIT('h08)
	) name1107 (
		_w2103_,
		_w2106_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1108 (
		_w2097_,
		_w2098_,
		_w2099_,
		_w2101_,
		_w2111_
	);
	LUT2 #(
		.INIT('h1)
	) name1109 (
		_w2102_,
		_w2111_,
		_w2112_
	);
	LUT4 #(
		.INIT('h00f2)
	) name1110 (
		_w2096_,
		_w2107_,
		_w2110_,
		_w2112_,
		_w2113_
	);
	LUT4 #(
		.INIT('h4055)
	) name1111 (
		_w2089_,
		_w2091_,
		_w2092_,
		_w2094_,
		_w2114_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w2093_,
		_w2114_,
		_w2115_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1113 (
		_w2096_,
		_w2107_,
		_w2110_,
		_w2112_,
		_w2116_
	);
	LUT3 #(
		.INIT('h54)
	) name1114 (
		_w2113_,
		_w2115_,
		_w2116_,
		_w2117_
	);
	LUT3 #(
		.INIT('h96)
	) name1115 (
		\A[349] ,
		\A[350] ,
		\A[351] ,
		_w2118_
	);
	LUT2 #(
		.INIT('h8)
	) name1116 (
		\A[352] ,
		\A[353] ,
		_w2119_
	);
	LUT3 #(
		.INIT('h96)
	) name1117 (
		\A[352] ,
		\A[353] ,
		\A[354] ,
		_w2120_
	);
	LUT3 #(
		.INIT('h96)
	) name1118 (
		\A[343] ,
		\A[344] ,
		\A[345] ,
		_w2121_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		\A[346] ,
		\A[347] ,
		_w2122_
	);
	LUT3 #(
		.INIT('h96)
	) name1120 (
		\A[346] ,
		\A[347] ,
		\A[348] ,
		_w2123_
	);
	LUT4 #(
		.INIT('h0660)
	) name1121 (
		_w2118_,
		_w2120_,
		_w2121_,
		_w2123_,
		_w2124_
	);
	LUT3 #(
		.INIT('h17)
	) name1122 (
		\A[349] ,
		\A[350] ,
		\A[351] ,
		_w2125_
	);
	LUT3 #(
		.INIT('h17)
	) name1123 (
		\A[352] ,
		\A[353] ,
		\A[354] ,
		_w2126_
	);
	LUT3 #(
		.INIT('h80)
	) name1124 (
		_w2118_,
		_w2119_,
		_w2120_,
		_w2127_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1125 (
		\A[352] ,
		\A[353] ,
		\A[354] ,
		_w2118_,
		_w2128_
	);
	LUT2 #(
		.INIT('h9)
	) name1126 (
		_w2125_,
		_w2128_,
		_w2129_
	);
	LUT3 #(
		.INIT('h14)
	) name1127 (
		_w2124_,
		_w2125_,
		_w2128_,
		_w2130_
	);
	LUT3 #(
		.INIT('h17)
	) name1128 (
		\A[343] ,
		\A[344] ,
		\A[345] ,
		_w2131_
	);
	LUT3 #(
		.INIT('h80)
	) name1129 (
		_w2121_,
		_w2122_,
		_w2123_,
		_w2132_
	);
	LUT3 #(
		.INIT('h17)
	) name1130 (
		\A[346] ,
		\A[347] ,
		\A[348] ,
		_w2133_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1131 (
		\A[346] ,
		\A[347] ,
		\A[348] ,
		_w2121_,
		_w2134_
	);
	LUT2 #(
		.INIT('h9)
	) name1132 (
		_w2131_,
		_w2134_,
		_w2135_
	);
	LUT3 #(
		.INIT('h82)
	) name1133 (
		_w2124_,
		_w2125_,
		_w2128_,
		_w2136_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		_w2125_,
		_w2126_,
		_w2137_
	);
	LUT4 #(
		.INIT('h0080)
	) name1135 (
		_w2121_,
		_w2122_,
		_w2123_,
		_w2131_,
		_w2138_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		_w2137_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('h171f)
	) name1137 (
		_w2124_,
		_w2129_,
		_w2135_,
		_w2139_,
		_w2140_
	);
	LUT4 #(
		.INIT('h080f)
	) name1138 (
		_w2118_,
		_w2120_,
		_w2125_,
		_w2126_,
		_w2141_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		_w2127_,
		_w2141_,
		_w2142_
	);
	LUT4 #(
		.INIT('h080f)
	) name1140 (
		_w2121_,
		_w2123_,
		_w2131_,
		_w2133_,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w2132_,
		_w2143_,
		_w2144_
	);
	LUT3 #(
		.INIT('he8)
	) name1142 (
		_w2140_,
		_w2142_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w2117_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		_w2117_,
		_w2145_,
		_w2147_
	);
	LUT3 #(
		.INIT('h69)
	) name1145 (
		_w2140_,
		_w2142_,
		_w2144_,
		_w2148_
	);
	LUT4 #(
		.INIT('hf20d)
	) name1146 (
		_w2096_,
		_w2107_,
		_w2110_,
		_w2112_,
		_w2149_
	);
	LUT2 #(
		.INIT('h9)
	) name1147 (
		_w2115_,
		_w2149_,
		_w2150_
	);
	LUT4 #(
		.INIT('h6996)
	) name1148 (
		_w2091_,
		_w2092_,
		_w2097_,
		_w2099_,
		_w2151_
	);
	LUT4 #(
		.INIT('h6996)
	) name1149 (
		_w2118_,
		_w2120_,
		_w2121_,
		_w2123_,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT4 #(
		.INIT('h89a9)
	) name1151 (
		_w2096_,
		_w2107_,
		_w2108_,
		_w2109_,
		_w2154_
	);
	LUT4 #(
		.INIT('hc989)
	) name1152 (
		_w2130_,
		_w2135_,
		_w2136_,
		_w2139_,
		_w2155_
	);
	LUT3 #(
		.INIT('he8)
	) name1153 (
		_w2153_,
		_w2154_,
		_w2155_,
		_w2156_
	);
	LUT3 #(
		.INIT('he8)
	) name1154 (
		_w2148_,
		_w2150_,
		_w2156_,
		_w2157_
	);
	LUT3 #(
		.INIT('h45)
	) name1155 (
		_w2146_,
		_w2147_,
		_w2157_,
		_w2158_
	);
	LUT3 #(
		.INIT('h17)
	) name1156 (
		\A[331] ,
		\A[332] ,
		\A[333] ,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1157 (
		\A[334] ,
		\A[335] ,
		_w2160_
	);
	LUT3 #(
		.INIT('h96)
	) name1158 (
		\A[331] ,
		\A[332] ,
		\A[333] ,
		_w2161_
	);
	LUT3 #(
		.INIT('h96)
	) name1159 (
		\A[334] ,
		\A[335] ,
		\A[336] ,
		_w2162_
	);
	LUT3 #(
		.INIT('h80)
	) name1160 (
		_w2160_,
		_w2161_,
		_w2162_,
		_w2163_
	);
	LUT3 #(
		.INIT('h17)
	) name1161 (
		\A[334] ,
		\A[335] ,
		\A[336] ,
		_w2164_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1162 (
		\A[334] ,
		\A[335] ,
		\A[336] ,
		_w2161_,
		_w2165_
	);
	LUT2 #(
		.INIT('h9)
	) name1163 (
		_w2159_,
		_w2165_,
		_w2166_
	);
	LUT3 #(
		.INIT('h96)
	) name1164 (
		\A[337] ,
		\A[338] ,
		\A[339] ,
		_w2167_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		\A[340] ,
		\A[341] ,
		_w2168_
	);
	LUT3 #(
		.INIT('h96)
	) name1166 (
		\A[340] ,
		\A[341] ,
		\A[342] ,
		_w2169_
	);
	LUT3 #(
		.INIT('h17)
	) name1167 (
		\A[340] ,
		\A[341] ,
		\A[342] ,
		_w2170_
	);
	LUT3 #(
		.INIT('h17)
	) name1168 (
		\A[337] ,
		\A[338] ,
		\A[339] ,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w2170_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h6)
	) name1170 (
		_w2170_,
		_w2171_,
		_w2173_
	);
	LUT4 #(
		.INIT('h8008)
	) name1171 (
		_w2167_,
		_w2169_,
		_w2170_,
		_w2171_,
		_w2174_
	);
	LUT4 #(
		.INIT('h0770)
	) name1172 (
		_w2167_,
		_w2169_,
		_w2170_,
		_w2171_,
		_w2175_
	);
	LUT4 #(
		.INIT('h0660)
	) name1173 (
		_w2161_,
		_w2162_,
		_w2167_,
		_w2169_,
		_w2176_
	);
	LUT3 #(
		.INIT('h01)
	) name1174 (
		_w2175_,
		_w2176_,
		_w2174_,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		_w2173_,
		_w2176_,
		_w2178_
	);
	LUT4 #(
		.INIT('h4000)
	) name1176 (
		_w2159_,
		_w2160_,
		_w2161_,
		_w2162_,
		_w2179_
	);
	LUT3 #(
		.INIT('h08)
	) name1177 (
		_w2173_,
		_w2176_,
		_w2179_,
		_w2180_
	);
	LUT3 #(
		.INIT('h0d)
	) name1178 (
		_w2166_,
		_w2177_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1179 (
		_w2167_,
		_w2168_,
		_w2169_,
		_w2171_,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w2172_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h00f2)
	) name1181 (
		_w2166_,
		_w2177_,
		_w2180_,
		_w2183_,
		_w2184_
	);
	LUT4 #(
		.INIT('h4055)
	) name1182 (
		_w2159_,
		_w2161_,
		_w2162_,
		_w2164_,
		_w2185_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w2163_,
		_w2185_,
		_w2186_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1184 (
		_w2166_,
		_w2177_,
		_w2180_,
		_w2183_,
		_w2187_
	);
	LUT3 #(
		.INIT('h96)
	) name1185 (
		\A[325] ,
		\A[326] ,
		\A[327] ,
		_w2188_
	);
	LUT3 #(
		.INIT('h96)
	) name1186 (
		\A[328] ,
		\A[329] ,
		\A[330] ,
		_w2189_
	);
	LUT2 #(
		.INIT('h8)
	) name1187 (
		_w2188_,
		_w2189_,
		_w2190_
	);
	LUT3 #(
		.INIT('h96)
	) name1188 (
		\A[319] ,
		\A[320] ,
		\A[321] ,
		_w2191_
	);
	LUT3 #(
		.INIT('h96)
	) name1189 (
		\A[322] ,
		\A[323] ,
		\A[324] ,
		_w2192_
	);
	LUT4 #(
		.INIT('h0660)
	) name1190 (
		_w2188_,
		_w2189_,
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT3 #(
		.INIT('h17)
	) name1191 (
		\A[328] ,
		\A[329] ,
		\A[330] ,
		_w2194_
	);
	LUT3 #(
		.INIT('h17)
	) name1192 (
		\A[325] ,
		\A[326] ,
		\A[327] ,
		_w2195_
	);
	LUT2 #(
		.INIT('h6)
	) name1193 (
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT3 #(
		.INIT('h17)
	) name1194 (
		\A[322] ,
		\A[323] ,
		\A[324] ,
		_w2197_
	);
	LUT3 #(
		.INIT('h17)
	) name1195 (
		\A[319] ,
		\A[320] ,
		\A[321] ,
		_w2198_
	);
	LUT4 #(
		.INIT('h7887)
	) name1196 (
		_w2191_,
		_w2192_,
		_w2197_,
		_w2198_,
		_w2199_
	);
	LUT4 #(
		.INIT('hc0de)
	) name1197 (
		_w2190_,
		_w2193_,
		_w2196_,
		_w2199_,
		_w2200_
	);
	LUT4 #(
		.INIT('h088f)
	) name1198 (
		_w2188_,
		_w2189_,
		_w2194_,
		_w2195_,
		_w2201_
	);
	LUT4 #(
		.INIT('h088f)
	) name1199 (
		_w2191_,
		_w2192_,
		_w2197_,
		_w2198_,
		_w2202_
	);
	LUT3 #(
		.INIT('he8)
	) name1200 (
		_w2200_,
		_w2201_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h1700)
	) name1201 (
		_w2181_,
		_w2183_,
		_w2186_,
		_w2203_,
		_w2204_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1202 (
		_w2181_,
		_w2183_,
		_w2186_,
		_w2203_,
		_w2205_
	);
	LUT4 #(
		.INIT('hf20d)
	) name1203 (
		_w2166_,
		_w2177_,
		_w2180_,
		_w2183_,
		_w2206_
	);
	LUT3 #(
		.INIT('h69)
	) name1204 (
		_w2200_,
		_w2201_,
		_w2202_,
		_w2207_
	);
	LUT3 #(
		.INIT('h09)
	) name1205 (
		_w2186_,
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT3 #(
		.INIT('h60)
	) name1206 (
		_w2186_,
		_w2206_,
		_w2207_,
		_w2209_
	);
	LUT4 #(
		.INIT('h6996)
	) name1207 (
		_w2161_,
		_w2162_,
		_w2167_,
		_w2169_,
		_w2210_
	);
	LUT4 #(
		.INIT('h6996)
	) name1208 (
		_w2188_,
		_w2189_,
		_w2191_,
		_w2192_,
		_w2211_
	);
	LUT2 #(
		.INIT('h8)
	) name1209 (
		_w2210_,
		_w2211_,
		_w2212_
	);
	LUT4 #(
		.INIT('h89a9)
	) name1210 (
		_w2166_,
		_w2177_,
		_w2178_,
		_w2179_,
		_w2213_
	);
	LUT4 #(
		.INIT('he11e)
	) name1211 (
		_w2190_,
		_w2193_,
		_w2196_,
		_w2199_,
		_w2214_
	);
	LUT3 #(
		.INIT('h71)
	) name1212 (
		_w2212_,
		_w2213_,
		_w2214_,
		_w2215_
	);
	LUT4 #(
		.INIT('h4445)
	) name1213 (
		_w2205_,
		_w2208_,
		_w2209_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w2204_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h1)
	) name1215 (
		_w2158_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		_w2158_,
		_w2217_,
		_w2219_
	);
	LUT2 #(
		.INIT('h6)
	) name1217 (
		_w2117_,
		_w2145_,
		_w2220_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1218 (
		_w2184_,
		_w2186_,
		_w2187_,
		_w2203_,
		_w2221_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1219 (
		_w2208_,
		_w2209_,
		_w2215_,
		_w2221_,
		_w2222_
	);
	LUT3 #(
		.INIT('h09)
	) name1220 (
		_w2157_,
		_w2220_,
		_w2222_,
		_w2223_
	);
	LUT3 #(
		.INIT('h60)
	) name1221 (
		_w2157_,
		_w2220_,
		_w2222_,
		_w2224_
	);
	LUT3 #(
		.INIT('h96)
	) name1222 (
		_w2148_,
		_w2150_,
		_w2156_,
		_w2225_
	);
	LUT3 #(
		.INIT('h96)
	) name1223 (
		_w2186_,
		_w2206_,
		_w2207_,
		_w2226_
	);
	LUT2 #(
		.INIT('h9)
	) name1224 (
		_w2215_,
		_w2226_,
		_w2227_
	);
	LUT4 #(
		.INIT('h0660)
	) name1225 (
		_w2151_,
		_w2152_,
		_w2210_,
		_w2211_,
		_w2228_
	);
	LUT4 #(
		.INIT('h9600)
	) name1226 (
		_w2153_,
		_w2154_,
		_w2155_,
		_w2228_,
		_w2229_
	);
	LUT4 #(
		.INIT('h0069)
	) name1227 (
		_w2153_,
		_w2154_,
		_w2155_,
		_w2228_,
		_w2230_
	);
	LUT3 #(
		.INIT('h69)
	) name1228 (
		_w2212_,
		_w2213_,
		_w2214_,
		_w2231_
	);
	LUT3 #(
		.INIT('h45)
	) name1229 (
		_w2229_,
		_w2230_,
		_w2231_,
		_w2232_
	);
	LUT3 #(
		.INIT('h71)
	) name1230 (
		_w2225_,
		_w2227_,
		_w2232_,
		_w2233_
	);
	LUT3 #(
		.INIT('h45)
	) name1231 (
		_w2223_,
		_w2224_,
		_w2233_,
		_w2234_
	);
	LUT3 #(
		.INIT('h96)
	) name1232 (
		\A[301] ,
		\A[302] ,
		\A[303] ,
		_w2235_
	);
	LUT3 #(
		.INIT('h96)
	) name1233 (
		\A[304] ,
		\A[305] ,
		\A[306] ,
		_w2236_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		_w2235_,
		_w2236_,
		_w2237_
	);
	LUT3 #(
		.INIT('h96)
	) name1235 (
		\A[295] ,
		\A[296] ,
		\A[297] ,
		_w2238_
	);
	LUT3 #(
		.INIT('h96)
	) name1236 (
		\A[298] ,
		\A[299] ,
		\A[300] ,
		_w2239_
	);
	LUT4 #(
		.INIT('h0660)
	) name1237 (
		_w2235_,
		_w2236_,
		_w2238_,
		_w2239_,
		_w2240_
	);
	LUT3 #(
		.INIT('h17)
	) name1238 (
		\A[304] ,
		\A[305] ,
		\A[306] ,
		_w2241_
	);
	LUT3 #(
		.INIT('h17)
	) name1239 (
		\A[301] ,
		\A[302] ,
		\A[303] ,
		_w2242_
	);
	LUT2 #(
		.INIT('h6)
	) name1240 (
		_w2241_,
		_w2242_,
		_w2243_
	);
	LUT3 #(
		.INIT('h17)
	) name1241 (
		\A[298] ,
		\A[299] ,
		\A[300] ,
		_w2244_
	);
	LUT3 #(
		.INIT('h17)
	) name1242 (
		\A[295] ,
		\A[296] ,
		\A[297] ,
		_w2245_
	);
	LUT4 #(
		.INIT('h7887)
	) name1243 (
		_w2238_,
		_w2239_,
		_w2244_,
		_w2245_,
		_w2246_
	);
	LUT4 #(
		.INIT('hc0de)
	) name1244 (
		_w2237_,
		_w2240_,
		_w2243_,
		_w2246_,
		_w2247_
	);
	LUT4 #(
		.INIT('h088f)
	) name1245 (
		_w2235_,
		_w2236_,
		_w2241_,
		_w2242_,
		_w2248_
	);
	LUT4 #(
		.INIT('h088f)
	) name1246 (
		_w2238_,
		_w2239_,
		_w2244_,
		_w2245_,
		_w2249_
	);
	LUT3 #(
		.INIT('he8)
	) name1247 (
		_w2247_,
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT3 #(
		.INIT('h69)
	) name1248 (
		_w2247_,
		_w2248_,
		_w2249_,
		_w2251_
	);
	LUT3 #(
		.INIT('h96)
	) name1249 (
		\A[313] ,
		\A[314] ,
		\A[315] ,
		_w2252_
	);
	LUT3 #(
		.INIT('h96)
	) name1250 (
		\A[316] ,
		\A[317] ,
		\A[318] ,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT3 #(
		.INIT('h96)
	) name1252 (
		\A[307] ,
		\A[308] ,
		\A[309] ,
		_w2255_
	);
	LUT3 #(
		.INIT('h96)
	) name1253 (
		\A[310] ,
		\A[311] ,
		\A[312] ,
		_w2256_
	);
	LUT4 #(
		.INIT('h0660)
	) name1254 (
		_w2252_,
		_w2253_,
		_w2255_,
		_w2256_,
		_w2257_
	);
	LUT3 #(
		.INIT('h17)
	) name1255 (
		\A[316] ,
		\A[317] ,
		\A[318] ,
		_w2258_
	);
	LUT3 #(
		.INIT('h17)
	) name1256 (
		\A[313] ,
		\A[314] ,
		\A[315] ,
		_w2259_
	);
	LUT2 #(
		.INIT('h6)
	) name1257 (
		_w2258_,
		_w2259_,
		_w2260_
	);
	LUT3 #(
		.INIT('h17)
	) name1258 (
		\A[310] ,
		\A[311] ,
		\A[312] ,
		_w2261_
	);
	LUT3 #(
		.INIT('h17)
	) name1259 (
		\A[307] ,
		\A[308] ,
		\A[309] ,
		_w2262_
	);
	LUT4 #(
		.INIT('h7887)
	) name1260 (
		_w2255_,
		_w2256_,
		_w2261_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('hc0de)
	) name1261 (
		_w2254_,
		_w2257_,
		_w2260_,
		_w2263_,
		_w2264_
	);
	LUT4 #(
		.INIT('h088f)
	) name1262 (
		_w2252_,
		_w2253_,
		_w2258_,
		_w2259_,
		_w2265_
	);
	LUT4 #(
		.INIT('h088f)
	) name1263 (
		_w2255_,
		_w2256_,
		_w2261_,
		_w2262_,
		_w2266_
	);
	LUT3 #(
		.INIT('h69)
	) name1264 (
		_w2264_,
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('h6996)
	) name1265 (
		_w2252_,
		_w2253_,
		_w2255_,
		_w2256_,
		_w2268_
	);
	LUT4 #(
		.INIT('h6996)
	) name1266 (
		_w2235_,
		_w2236_,
		_w2238_,
		_w2239_,
		_w2269_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		_w2268_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('he11e)
	) name1268 (
		_w2254_,
		_w2257_,
		_w2260_,
		_w2263_,
		_w2271_
	);
	LUT4 #(
		.INIT('he11e)
	) name1269 (
		_w2237_,
		_w2240_,
		_w2243_,
		_w2246_,
		_w2272_
	);
	LUT3 #(
		.INIT('hd4)
	) name1270 (
		_w2270_,
		_w2271_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h022a)
	) name1271 (
		_w2250_,
		_w2251_,
		_w2267_,
		_w2273_,
		_w2274_
	);
	LUT4 #(
		.INIT('h5440)
	) name1272 (
		_w2250_,
		_w2251_,
		_w2267_,
		_w2273_,
		_w2275_
	);
	LUT3 #(
		.INIT('he8)
	) name1273 (
		_w2264_,
		_w2265_,
		_w2266_,
		_w2276_
	);
	LUT3 #(
		.INIT('h45)
	) name1274 (
		_w2274_,
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT3 #(
		.INIT('h96)
	) name1275 (
		\A[277] ,
		\A[278] ,
		\A[279] ,
		_w2278_
	);
	LUT3 #(
		.INIT('h96)
	) name1276 (
		\A[280] ,
		\A[281] ,
		\A[282] ,
		_w2279_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT3 #(
		.INIT('h96)
	) name1278 (
		\A[271] ,
		\A[272] ,
		\A[273] ,
		_w2281_
	);
	LUT3 #(
		.INIT('h96)
	) name1279 (
		\A[274] ,
		\A[275] ,
		\A[276] ,
		_w2282_
	);
	LUT4 #(
		.INIT('h0660)
	) name1280 (
		_w2278_,
		_w2279_,
		_w2281_,
		_w2282_,
		_w2283_
	);
	LUT3 #(
		.INIT('h17)
	) name1281 (
		\A[280] ,
		\A[281] ,
		\A[282] ,
		_w2284_
	);
	LUT3 #(
		.INIT('h17)
	) name1282 (
		\A[277] ,
		\A[278] ,
		\A[279] ,
		_w2285_
	);
	LUT2 #(
		.INIT('h6)
	) name1283 (
		_w2284_,
		_w2285_,
		_w2286_
	);
	LUT3 #(
		.INIT('h17)
	) name1284 (
		\A[274] ,
		\A[275] ,
		\A[276] ,
		_w2287_
	);
	LUT3 #(
		.INIT('h17)
	) name1285 (
		\A[271] ,
		\A[272] ,
		\A[273] ,
		_w2288_
	);
	LUT4 #(
		.INIT('h7887)
	) name1286 (
		_w2281_,
		_w2282_,
		_w2287_,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('hc0de)
	) name1287 (
		_w2280_,
		_w2283_,
		_w2286_,
		_w2289_,
		_w2290_
	);
	LUT4 #(
		.INIT('h088f)
	) name1288 (
		_w2278_,
		_w2279_,
		_w2284_,
		_w2285_,
		_w2291_
	);
	LUT4 #(
		.INIT('h088f)
	) name1289 (
		_w2281_,
		_w2282_,
		_w2287_,
		_w2288_,
		_w2292_
	);
	LUT3 #(
		.INIT('he8)
	) name1290 (
		_w2290_,
		_w2291_,
		_w2292_,
		_w2293_
	);
	LUT3 #(
		.INIT('h69)
	) name1291 (
		_w2290_,
		_w2291_,
		_w2292_,
		_w2294_
	);
	LUT3 #(
		.INIT('h96)
	) name1292 (
		\A[289] ,
		\A[290] ,
		\A[291] ,
		_w2295_
	);
	LUT3 #(
		.INIT('h96)
	) name1293 (
		\A[292] ,
		\A[293] ,
		\A[294] ,
		_w2296_
	);
	LUT2 #(
		.INIT('h8)
	) name1294 (
		_w2295_,
		_w2296_,
		_w2297_
	);
	LUT3 #(
		.INIT('h96)
	) name1295 (
		\A[283] ,
		\A[284] ,
		\A[285] ,
		_w2298_
	);
	LUT3 #(
		.INIT('h96)
	) name1296 (
		\A[286] ,
		\A[287] ,
		\A[288] ,
		_w2299_
	);
	LUT4 #(
		.INIT('h0660)
	) name1297 (
		_w2295_,
		_w2296_,
		_w2298_,
		_w2299_,
		_w2300_
	);
	LUT3 #(
		.INIT('h17)
	) name1298 (
		\A[292] ,
		\A[293] ,
		\A[294] ,
		_w2301_
	);
	LUT3 #(
		.INIT('h17)
	) name1299 (
		\A[289] ,
		\A[290] ,
		\A[291] ,
		_w2302_
	);
	LUT2 #(
		.INIT('h6)
	) name1300 (
		_w2301_,
		_w2302_,
		_w2303_
	);
	LUT3 #(
		.INIT('h17)
	) name1301 (
		\A[286] ,
		\A[287] ,
		\A[288] ,
		_w2304_
	);
	LUT3 #(
		.INIT('h17)
	) name1302 (
		\A[283] ,
		\A[284] ,
		\A[285] ,
		_w2305_
	);
	LUT4 #(
		.INIT('h7887)
	) name1303 (
		_w2298_,
		_w2299_,
		_w2304_,
		_w2305_,
		_w2306_
	);
	LUT4 #(
		.INIT('hc0de)
	) name1304 (
		_w2297_,
		_w2300_,
		_w2303_,
		_w2306_,
		_w2307_
	);
	LUT4 #(
		.INIT('h088f)
	) name1305 (
		_w2295_,
		_w2296_,
		_w2301_,
		_w2302_,
		_w2308_
	);
	LUT4 #(
		.INIT('h088f)
	) name1306 (
		_w2298_,
		_w2299_,
		_w2304_,
		_w2305_,
		_w2309_
	);
	LUT3 #(
		.INIT('h69)
	) name1307 (
		_w2307_,
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('h6996)
	) name1308 (
		_w2295_,
		_w2296_,
		_w2298_,
		_w2299_,
		_w2311_
	);
	LUT4 #(
		.INIT('h6996)
	) name1309 (
		_w2278_,
		_w2279_,
		_w2281_,
		_w2282_,
		_w2312_
	);
	LUT2 #(
		.INIT('h8)
	) name1310 (
		_w2311_,
		_w2312_,
		_w2313_
	);
	LUT4 #(
		.INIT('he11e)
	) name1311 (
		_w2297_,
		_w2300_,
		_w2303_,
		_w2306_,
		_w2314_
	);
	LUT4 #(
		.INIT('he11e)
	) name1312 (
		_w2280_,
		_w2283_,
		_w2286_,
		_w2289_,
		_w2315_
	);
	LUT3 #(
		.INIT('hd4)
	) name1313 (
		_w2313_,
		_w2314_,
		_w2315_,
		_w2316_
	);
	LUT4 #(
		.INIT('h022a)
	) name1314 (
		_w2293_,
		_w2294_,
		_w2310_,
		_w2316_,
		_w2317_
	);
	LUT4 #(
		.INIT('h5440)
	) name1315 (
		_w2293_,
		_w2294_,
		_w2310_,
		_w2316_,
		_w2318_
	);
	LUT3 #(
		.INIT('he8)
	) name1316 (
		_w2307_,
		_w2308_,
		_w2309_,
		_w2319_
	);
	LUT3 #(
		.INIT('h45)
	) name1317 (
		_w2317_,
		_w2318_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h1)
	) name1318 (
		_w2277_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('h8)
	) name1319 (
		_w2277_,
		_w2320_,
		_w2322_
	);
	LUT4 #(
		.INIT('ha995)
	) name1320 (
		_w2250_,
		_w2251_,
		_w2267_,
		_w2273_,
		_w2323_
	);
	LUT4 #(
		.INIT('ha995)
	) name1321 (
		_w2293_,
		_w2294_,
		_w2310_,
		_w2316_,
		_w2324_
	);
	LUT4 #(
		.INIT('h8421)
	) name1322 (
		_w2276_,
		_w2319_,
		_w2323_,
		_w2324_,
		_w2325_
	);
	LUT4 #(
		.INIT('h1248)
	) name1323 (
		_w2276_,
		_w2319_,
		_w2323_,
		_w2324_,
		_w2326_
	);
	LUT3 #(
		.INIT('h69)
	) name1324 (
		_w2294_,
		_w2310_,
		_w2316_,
		_w2327_
	);
	LUT3 #(
		.INIT('h69)
	) name1325 (
		_w2251_,
		_w2267_,
		_w2273_,
		_w2328_
	);
	LUT4 #(
		.INIT('h0660)
	) name1326 (
		_w2268_,
		_w2269_,
		_w2311_,
		_w2312_,
		_w2329_
	);
	LUT4 #(
		.INIT('h9600)
	) name1327 (
		_w2270_,
		_w2271_,
		_w2272_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('h0069)
	) name1328 (
		_w2270_,
		_w2271_,
		_w2272_,
		_w2329_,
		_w2331_
	);
	LUT3 #(
		.INIT('h96)
	) name1329 (
		_w2313_,
		_w2314_,
		_w2315_,
		_w2332_
	);
	LUT3 #(
		.INIT('h45)
	) name1330 (
		_w2330_,
		_w2331_,
		_w2332_,
		_w2333_
	);
	LUT3 #(
		.INIT('h8e)
	) name1331 (
		_w2327_,
		_w2328_,
		_w2333_,
		_w2334_
	);
	LUT3 #(
		.INIT('h54)
	) name1332 (
		_w2325_,
		_w2326_,
		_w2334_,
		_w2335_
	);
	LUT3 #(
		.INIT('h45)
	) name1333 (
		_w2321_,
		_w2322_,
		_w2335_,
		_w2336_
	);
	LUT4 #(
		.INIT('h0071)
	) name1334 (
		_w2158_,
		_w2217_,
		_w2234_,
		_w2336_,
		_w2337_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1335 (
		_w2158_,
		_w2217_,
		_w2234_,
		_w2336_,
		_w2338_
	);
	LUT2 #(
		.INIT('h6)
	) name1336 (
		_w2158_,
		_w2217_,
		_w2339_
	);
	LUT2 #(
		.INIT('h6)
	) name1337 (
		_w2277_,
		_w2320_,
		_w2340_
	);
	LUT2 #(
		.INIT('h9)
	) name1338 (
		_w2335_,
		_w2340_,
		_w2341_
	);
	LUT3 #(
		.INIT('h06)
	) name1339 (
		_w2234_,
		_w2339_,
		_w2341_,
		_w2342_
	);
	LUT3 #(
		.INIT('h90)
	) name1340 (
		_w2234_,
		_w2339_,
		_w2341_,
		_w2343_
	);
	LUT4 #(
		.INIT('h6996)
	) name1341 (
		_w2276_,
		_w2319_,
		_w2323_,
		_w2324_,
		_w2344_
	);
	LUT2 #(
		.INIT('h9)
	) name1342 (
		_w2334_,
		_w2344_,
		_w2345_
	);
	LUT3 #(
		.INIT('h96)
	) name1343 (
		_w2157_,
		_w2220_,
		_w2222_,
		_w2346_
	);
	LUT3 #(
		.INIT('h21)
	) name1344 (
		_w2233_,
		_w2345_,
		_w2346_,
		_w2347_
	);
	LUT3 #(
		.INIT('h48)
	) name1345 (
		_w2233_,
		_w2345_,
		_w2346_,
		_w2348_
	);
	LUT3 #(
		.INIT('h69)
	) name1346 (
		_w2327_,
		_w2328_,
		_w2333_,
		_w2349_
	);
	LUT4 #(
		.INIT('h0096)
	) name1347 (
		_w2225_,
		_w2227_,
		_w2232_,
		_w2349_,
		_w2350_
	);
	LUT4 #(
		.INIT('h6900)
	) name1348 (
		_w2225_,
		_w2227_,
		_w2232_,
		_w2349_,
		_w2351_
	);
	LUT4 #(
		.INIT('h6996)
	) name1349 (
		_w2151_,
		_w2152_,
		_w2210_,
		_w2211_,
		_w2352_
	);
	LUT4 #(
		.INIT('h6996)
	) name1350 (
		_w2268_,
		_w2269_,
		_w2311_,
		_w2312_,
		_w2353_
	);
	LUT2 #(
		.INIT('h8)
	) name1351 (
		_w2352_,
		_w2353_,
		_w2354_
	);
	LUT4 #(
		.INIT('h6996)
	) name1352 (
		_w2153_,
		_w2154_,
		_w2155_,
		_w2228_,
		_w2355_
	);
	LUT4 #(
		.INIT('h6996)
	) name1353 (
		_w2270_,
		_w2271_,
		_w2272_,
		_w2329_,
		_w2356_
	);
	LUT2 #(
		.INIT('h9)
	) name1354 (
		_w2332_,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('hb721)
	) name1355 (
		_w2231_,
		_w2354_,
		_w2355_,
		_w2357_,
		_w2358_
	);
	LUT3 #(
		.INIT('h45)
	) name1356 (
		_w2350_,
		_w2351_,
		_w2358_,
		_w2359_
	);
	LUT3 #(
		.INIT('h45)
	) name1357 (
		_w2347_,
		_w2348_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('h4445)
	) name1358 (
		_w2338_,
		_w2342_,
		_w2343_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		_w2337_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		_w2088_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		_w2088_,
		_w2362_,
		_w2364_
	);
	LUT2 #(
		.INIT('h6)
	) name1362 (
		_w1919_,
		_w2061_,
		_w2365_
	);
	LUT4 #(
		.INIT('hba45)
	) name1363 (
		_w2218_,
		_w2219_,
		_w2234_,
		_w2336_,
		_w2366_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1364 (
		_w2342_,
		_w2343_,
		_w2360_,
		_w2366_,
		_w2367_
	);
	LUT3 #(
		.INIT('h09)
	) name1365 (
		_w2087_,
		_w2365_,
		_w2367_,
		_w2368_
	);
	LUT3 #(
		.INIT('h60)
	) name1366 (
		_w2087_,
		_w2365_,
		_w2367_,
		_w2369_
	);
	LUT3 #(
		.INIT('h69)
	) name1367 (
		_w2234_,
		_w2339_,
		_w2341_,
		_w2370_
	);
	LUT3 #(
		.INIT('h96)
	) name1368 (
		_w1918_,
		_w2065_,
		_w2066_,
		_w2371_
	);
	LUT4 #(
		.INIT('h2814)
	) name1369 (
		_w2086_,
		_w2360_,
		_w2370_,
		_w2371_,
		_w2372_
	);
	LUT4 #(
		.INIT('h4182)
	) name1370 (
		_w2086_,
		_w2360_,
		_w2370_,
		_w2371_,
		_w2373_
	);
	LUT4 #(
		.INIT('h6996)
	) name1371 (
		_w1917_,
		_w2059_,
		_w2069_,
		_w2070_,
		_w2374_
	);
	LUT3 #(
		.INIT('h96)
	) name1372 (
		_w2233_,
		_w2345_,
		_w2346_,
		_w2375_
	);
	LUT4 #(
		.INIT('h8421)
	) name1373 (
		_w2085_,
		_w2359_,
		_w2374_,
		_w2375_,
		_w2376_
	);
	LUT4 #(
		.INIT('h1248)
	) name1374 (
		_w2085_,
		_w2359_,
		_w2374_,
		_w2375_,
		_w2377_
	);
	LUT4 #(
		.INIT('h9669)
	) name1375 (
		_w2225_,
		_w2227_,
		_w2232_,
		_w2349_,
		_w2378_
	);
	LUT2 #(
		.INIT('h9)
	) name1376 (
		_w2358_,
		_w2378_,
		_w2379_
	);
	LUT3 #(
		.INIT('h69)
	) name1377 (
		_w2073_,
		_w2075_,
		_w2084_,
		_w2380_
	);
	LUT4 #(
		.INIT('h0660)
	) name1378 (
		_w2076_,
		_w2077_,
		_w2352_,
		_w2353_,
		_w2381_
	);
	LUT3 #(
		.INIT('h96)
	) name1379 (
		_w2057_,
		_w2078_,
		_w2079_,
		_w2382_
	);
	LUT4 #(
		.INIT('h9669)
	) name1380 (
		_w2231_,
		_w2354_,
		_w2355_,
		_w2357_,
		_w2383_
	);
	LUT4 #(
		.INIT('h127b)
	) name1381 (
		_w2083_,
		_w2381_,
		_w2382_,
		_w2383_,
		_w2384_
	);
	LUT3 #(
		.INIT('h8e)
	) name1382 (
		_w2379_,
		_w2380_,
		_w2384_,
		_w2385_
	);
	LUT3 #(
		.INIT('h54)
	) name1383 (
		_w2376_,
		_w2377_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('h54)
	) name1384 (
		_w2372_,
		_w2373_,
		_w2386_,
		_w2387_
	);
	LUT3 #(
		.INIT('h54)
	) name1385 (
		_w2368_,
		_w2369_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h45)
	) name1386 (
		_w2363_,
		_w2364_,
		_w2388_,
		_w2389_
	);
	LUT3 #(
		.INIT('h17)
	) name1387 (
		\A[211] ,
		\A[212] ,
		\A[213] ,
		_w2390_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		\A[214] ,
		\A[215] ,
		_w2391_
	);
	LUT3 #(
		.INIT('h96)
	) name1389 (
		\A[211] ,
		\A[212] ,
		\A[213] ,
		_w2392_
	);
	LUT3 #(
		.INIT('h96)
	) name1390 (
		\A[214] ,
		\A[215] ,
		\A[216] ,
		_w2393_
	);
	LUT3 #(
		.INIT('h80)
	) name1391 (
		_w2391_,
		_w2392_,
		_w2393_,
		_w2394_
	);
	LUT3 #(
		.INIT('h17)
	) name1392 (
		\A[214] ,
		\A[215] ,
		\A[216] ,
		_w2395_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1393 (
		\A[214] ,
		\A[215] ,
		\A[216] ,
		_w2392_,
		_w2396_
	);
	LUT2 #(
		.INIT('h9)
	) name1394 (
		_w2390_,
		_w2396_,
		_w2397_
	);
	LUT3 #(
		.INIT('h96)
	) name1395 (
		\A[217] ,
		\A[218] ,
		\A[219] ,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name1396 (
		\A[220] ,
		\A[221] ,
		_w2399_
	);
	LUT3 #(
		.INIT('h96)
	) name1397 (
		\A[220] ,
		\A[221] ,
		\A[222] ,
		_w2400_
	);
	LUT3 #(
		.INIT('h17)
	) name1398 (
		\A[220] ,
		\A[221] ,
		\A[222] ,
		_w2401_
	);
	LUT3 #(
		.INIT('h17)
	) name1399 (
		\A[217] ,
		\A[218] ,
		\A[219] ,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name1400 (
		_w2401_,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h6)
	) name1401 (
		_w2401_,
		_w2402_,
		_w2404_
	);
	LUT4 #(
		.INIT('h8008)
	) name1402 (
		_w2398_,
		_w2400_,
		_w2401_,
		_w2402_,
		_w2405_
	);
	LUT4 #(
		.INIT('h0770)
	) name1403 (
		_w2398_,
		_w2400_,
		_w2401_,
		_w2402_,
		_w2406_
	);
	LUT4 #(
		.INIT('h0660)
	) name1404 (
		_w2392_,
		_w2393_,
		_w2398_,
		_w2400_,
		_w2407_
	);
	LUT3 #(
		.INIT('h01)
	) name1405 (
		_w2406_,
		_w2407_,
		_w2405_,
		_w2408_
	);
	LUT2 #(
		.INIT('h8)
	) name1406 (
		_w2404_,
		_w2407_,
		_w2409_
	);
	LUT4 #(
		.INIT('h4000)
	) name1407 (
		_w2390_,
		_w2391_,
		_w2392_,
		_w2393_,
		_w2410_
	);
	LUT3 #(
		.INIT('h08)
	) name1408 (
		_w2404_,
		_w2407_,
		_w2410_,
		_w2411_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1409 (
		_w2398_,
		_w2399_,
		_w2400_,
		_w2402_,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		_w2403_,
		_w2412_,
		_w2413_
	);
	LUT4 #(
		.INIT('h00f2)
	) name1411 (
		_w2397_,
		_w2408_,
		_w2411_,
		_w2413_,
		_w2414_
	);
	LUT4 #(
		.INIT('h4055)
	) name1412 (
		_w2390_,
		_w2392_,
		_w2393_,
		_w2395_,
		_w2415_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w2394_,
		_w2415_,
		_w2416_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1414 (
		_w2397_,
		_w2408_,
		_w2411_,
		_w2413_,
		_w2417_
	);
	LUT3 #(
		.INIT('h54)
	) name1415 (
		_w2414_,
		_w2416_,
		_w2417_,
		_w2418_
	);
	LUT3 #(
		.INIT('h96)
	) name1416 (
		\A[205] ,
		\A[206] ,
		\A[207] ,
		_w2419_
	);
	LUT2 #(
		.INIT('h8)
	) name1417 (
		\A[208] ,
		\A[209] ,
		_w2420_
	);
	LUT3 #(
		.INIT('h96)
	) name1418 (
		\A[208] ,
		\A[209] ,
		\A[210] ,
		_w2421_
	);
	LUT3 #(
		.INIT('h96)
	) name1419 (
		\A[199] ,
		\A[200] ,
		\A[201] ,
		_w2422_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		\A[202] ,
		\A[203] ,
		_w2423_
	);
	LUT3 #(
		.INIT('h96)
	) name1421 (
		\A[202] ,
		\A[203] ,
		\A[204] ,
		_w2424_
	);
	LUT4 #(
		.INIT('h0660)
	) name1422 (
		_w2419_,
		_w2421_,
		_w2422_,
		_w2424_,
		_w2425_
	);
	LUT3 #(
		.INIT('h17)
	) name1423 (
		\A[205] ,
		\A[206] ,
		\A[207] ,
		_w2426_
	);
	LUT3 #(
		.INIT('h17)
	) name1424 (
		\A[208] ,
		\A[209] ,
		\A[210] ,
		_w2427_
	);
	LUT3 #(
		.INIT('h80)
	) name1425 (
		_w2419_,
		_w2420_,
		_w2421_,
		_w2428_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1426 (
		\A[208] ,
		\A[209] ,
		\A[210] ,
		_w2419_,
		_w2429_
	);
	LUT2 #(
		.INIT('h9)
	) name1427 (
		_w2426_,
		_w2429_,
		_w2430_
	);
	LUT3 #(
		.INIT('h14)
	) name1428 (
		_w2425_,
		_w2426_,
		_w2429_,
		_w2431_
	);
	LUT3 #(
		.INIT('h17)
	) name1429 (
		\A[199] ,
		\A[200] ,
		\A[201] ,
		_w2432_
	);
	LUT3 #(
		.INIT('h80)
	) name1430 (
		_w2422_,
		_w2423_,
		_w2424_,
		_w2433_
	);
	LUT3 #(
		.INIT('h17)
	) name1431 (
		\A[202] ,
		\A[203] ,
		\A[204] ,
		_w2434_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1432 (
		\A[202] ,
		\A[203] ,
		\A[204] ,
		_w2422_,
		_w2435_
	);
	LUT2 #(
		.INIT('h9)
	) name1433 (
		_w2432_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('h82)
	) name1434 (
		_w2425_,
		_w2426_,
		_w2429_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w2426_,
		_w2427_,
		_w2438_
	);
	LUT4 #(
		.INIT('h0080)
	) name1436 (
		_w2422_,
		_w2423_,
		_w2424_,
		_w2432_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT4 #(
		.INIT('h171f)
	) name1438 (
		_w2425_,
		_w2430_,
		_w2436_,
		_w2440_,
		_w2441_
	);
	LUT4 #(
		.INIT('h080f)
	) name1439 (
		_w2419_,
		_w2421_,
		_w2426_,
		_w2427_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		_w2428_,
		_w2442_,
		_w2443_
	);
	LUT4 #(
		.INIT('h080f)
	) name1441 (
		_w2422_,
		_w2424_,
		_w2432_,
		_w2434_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		_w2433_,
		_w2444_,
		_w2445_
	);
	LUT3 #(
		.INIT('he8)
	) name1443 (
		_w2441_,
		_w2443_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h1)
	) name1444 (
		_w2418_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		_w2418_,
		_w2446_,
		_w2448_
	);
	LUT3 #(
		.INIT('h69)
	) name1446 (
		_w2441_,
		_w2443_,
		_w2445_,
		_w2449_
	);
	LUT4 #(
		.INIT('hf20d)
	) name1447 (
		_w2397_,
		_w2408_,
		_w2411_,
		_w2413_,
		_w2450_
	);
	LUT2 #(
		.INIT('h9)
	) name1448 (
		_w2416_,
		_w2450_,
		_w2451_
	);
	LUT4 #(
		.INIT('h6996)
	) name1449 (
		_w2392_,
		_w2393_,
		_w2398_,
		_w2400_,
		_w2452_
	);
	LUT4 #(
		.INIT('h6996)
	) name1450 (
		_w2419_,
		_w2421_,
		_w2422_,
		_w2424_,
		_w2453_
	);
	LUT2 #(
		.INIT('h8)
	) name1451 (
		_w2452_,
		_w2453_,
		_w2454_
	);
	LUT4 #(
		.INIT('h89a9)
	) name1452 (
		_w2397_,
		_w2408_,
		_w2409_,
		_w2410_,
		_w2455_
	);
	LUT4 #(
		.INIT('hc989)
	) name1453 (
		_w2431_,
		_w2436_,
		_w2437_,
		_w2440_,
		_w2456_
	);
	LUT3 #(
		.INIT('he8)
	) name1454 (
		_w2454_,
		_w2455_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('he8)
	) name1455 (
		_w2449_,
		_w2451_,
		_w2457_,
		_w2458_
	);
	LUT3 #(
		.INIT('h45)
	) name1456 (
		_w2447_,
		_w2448_,
		_w2458_,
		_w2459_
	);
	LUT3 #(
		.INIT('h96)
	) name1457 (
		\A[193] ,
		\A[194] ,
		\A[195] ,
		_w2460_
	);
	LUT3 #(
		.INIT('h96)
	) name1458 (
		\A[196] ,
		\A[197] ,
		\A[198] ,
		_w2461_
	);
	LUT2 #(
		.INIT('h8)
	) name1459 (
		_w2460_,
		_w2461_,
		_w2462_
	);
	LUT3 #(
		.INIT('h96)
	) name1460 (
		\A[187] ,
		\A[188] ,
		\A[189] ,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		\A[190] ,
		\A[191] ,
		_w2464_
	);
	LUT3 #(
		.INIT('h96)
	) name1462 (
		\A[190] ,
		\A[191] ,
		\A[192] ,
		_w2465_
	);
	LUT4 #(
		.INIT('h0660)
	) name1463 (
		_w2460_,
		_w2461_,
		_w2463_,
		_w2465_,
		_w2466_
	);
	LUT3 #(
		.INIT('h17)
	) name1464 (
		\A[196] ,
		\A[197] ,
		\A[198] ,
		_w2467_
	);
	LUT3 #(
		.INIT('h17)
	) name1465 (
		\A[193] ,
		\A[194] ,
		\A[195] ,
		_w2468_
	);
	LUT2 #(
		.INIT('h6)
	) name1466 (
		_w2467_,
		_w2468_,
		_w2469_
	);
	LUT3 #(
		.INIT('h17)
	) name1467 (
		\A[187] ,
		\A[188] ,
		\A[189] ,
		_w2470_
	);
	LUT3 #(
		.INIT('h17)
	) name1468 (
		\A[190] ,
		\A[191] ,
		\A[192] ,
		_w2471_
	);
	LUT3 #(
		.INIT('h80)
	) name1469 (
		_w2463_,
		_w2464_,
		_w2465_,
		_w2472_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1470 (
		\A[190] ,
		\A[191] ,
		\A[192] ,
		_w2463_,
		_w2473_
	);
	LUT2 #(
		.INIT('h9)
	) name1471 (
		_w2470_,
		_w2473_,
		_w2474_
	);
	LUT4 #(
		.INIT('h0770)
	) name1472 (
		_w2466_,
		_w2469_,
		_w2470_,
		_w2473_,
		_w2475_
	);
	LUT4 #(
		.INIT('h8008)
	) name1473 (
		_w2460_,
		_w2461_,
		_w2467_,
		_w2468_,
		_w2476_
	);
	LUT4 #(
		.INIT('h0770)
	) name1474 (
		_w2460_,
		_w2461_,
		_w2467_,
		_w2468_,
		_w2477_
	);
	LUT3 #(
		.INIT('h01)
	) name1475 (
		_w2466_,
		_w2477_,
		_w2476_,
		_w2478_
	);
	LUT4 #(
		.INIT('h088f)
	) name1476 (
		_w2460_,
		_w2461_,
		_w2467_,
		_w2468_,
		_w2479_
	);
	LUT4 #(
		.INIT('h080f)
	) name1477 (
		_w2463_,
		_w2465_,
		_w2470_,
		_w2471_,
		_w2480_
	);
	LUT2 #(
		.INIT('h1)
	) name1478 (
		_w2472_,
		_w2480_,
		_w2481_
	);
	LUT4 #(
		.INIT('h10f1)
	) name1479 (
		_w2475_,
		_w2478_,
		_w2479_,
		_w2481_,
		_w2482_
	);
	LUT4 #(
		.INIT('he11e)
	) name1480 (
		_w2475_,
		_w2478_,
		_w2479_,
		_w2481_,
		_w2483_
	);
	LUT2 #(
		.INIT('h8)
	) name1481 (
		\A[178] ,
		\A[179] ,
		_w2484_
	);
	LUT3 #(
		.INIT('h96)
	) name1482 (
		\A[175] ,
		\A[176] ,
		\A[177] ,
		_w2485_
	);
	LUT3 #(
		.INIT('h96)
	) name1483 (
		\A[178] ,
		\A[179] ,
		\A[180] ,
		_w2486_
	);
	LUT3 #(
		.INIT('h80)
	) name1484 (
		_w2484_,
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT3 #(
		.INIT('h17)
	) name1485 (
		\A[175] ,
		\A[176] ,
		\A[177] ,
		_w2488_
	);
	LUT3 #(
		.INIT('h17)
	) name1486 (
		\A[178] ,
		\A[179] ,
		\A[180] ,
		_w2489_
	);
	LUT4 #(
		.INIT('h080f)
	) name1487 (
		_w2485_,
		_w2486_,
		_w2488_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h1)
	) name1488 (
		_w2487_,
		_w2490_,
		_w2491_
	);
	LUT3 #(
		.INIT('h96)
	) name1489 (
		\A[181] ,
		\A[182] ,
		\A[183] ,
		_w2492_
	);
	LUT3 #(
		.INIT('h96)
	) name1490 (
		\A[184] ,
		\A[185] ,
		\A[186] ,
		_w2493_
	);
	LUT2 #(
		.INIT('h8)
	) name1491 (
		_w2492_,
		_w2493_,
		_w2494_
	);
	LUT4 #(
		.INIT('h0660)
	) name1492 (
		_w2485_,
		_w2486_,
		_w2492_,
		_w2493_,
		_w2495_
	);
	LUT3 #(
		.INIT('h17)
	) name1493 (
		\A[184] ,
		\A[185] ,
		\A[186] ,
		_w2496_
	);
	LUT3 #(
		.INIT('h17)
	) name1494 (
		\A[181] ,
		\A[182] ,
		\A[183] ,
		_w2497_
	);
	LUT2 #(
		.INIT('h6)
	) name1495 (
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1496 (
		\A[178] ,
		\A[179] ,
		\A[180] ,
		_w2485_,
		_w2499_
	);
	LUT2 #(
		.INIT('h9)
	) name1497 (
		_w2488_,
		_w2499_,
		_w2500_
	);
	LUT4 #(
		.INIT('h152a)
	) name1498 (
		_w2488_,
		_w2495_,
		_w2498_,
		_w2499_,
		_w2501_
	);
	LUT4 #(
		.INIT('h8008)
	) name1499 (
		_w2492_,
		_w2493_,
		_w2496_,
		_w2497_,
		_w2502_
	);
	LUT4 #(
		.INIT('h0770)
	) name1500 (
		_w2492_,
		_w2493_,
		_w2496_,
		_w2497_,
		_w2503_
	);
	LUT3 #(
		.INIT('h01)
	) name1501 (
		_w2495_,
		_w2503_,
		_w2502_,
		_w2504_
	);
	LUT4 #(
		.INIT('h088f)
	) name1502 (
		_w2492_,
		_w2493_,
		_w2496_,
		_w2497_,
		_w2505_
	);
	LUT4 #(
		.INIT('ha956)
	) name1503 (
		_w2491_,
		_w2501_,
		_w2504_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h8)
	) name1504 (
		_w2483_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w2483_,
		_w2506_,
		_w2508_
	);
	LUT4 #(
		.INIT('h6996)
	) name1506 (
		_w2460_,
		_w2461_,
		_w2463_,
		_w2465_,
		_w2509_
	);
	LUT4 #(
		.INIT('h6996)
	) name1507 (
		_w2485_,
		_w2486_,
		_w2492_,
		_w2493_,
		_w2510_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		_w2509_,
		_w2510_,
		_w2511_
	);
	LUT3 #(
		.INIT('h1e)
	) name1509 (
		_w2462_,
		_w2466_,
		_w2469_,
		_w2512_
	);
	LUT3 #(
		.INIT('h48)
	) name1510 (
		_w2474_,
		_w2511_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('h21)
	) name1511 (
		_w2474_,
		_w2511_,
		_w2512_,
		_w2514_
	);
	LUT3 #(
		.INIT('h1e)
	) name1512 (
		_w2494_,
		_w2495_,
		_w2498_,
		_w2515_
	);
	LUT2 #(
		.INIT('h9)
	) name1513 (
		_w2500_,
		_w2515_,
		_w2516_
	);
	LUT3 #(
		.INIT('h54)
	) name1514 (
		_w2513_,
		_w2514_,
		_w2516_,
		_w2517_
	);
	LUT4 #(
		.INIT('h80a8)
	) name1515 (
		_w2482_,
		_w2483_,
		_w2506_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('h1501)
	) name1516 (
		_w2482_,
		_w2483_,
		_w2506_,
		_w2517_,
		_w2519_
	);
	LUT4 #(
		.INIT('h5701)
	) name1517 (
		_w2491_,
		_w2501_,
		_w2504_,
		_w2505_,
		_w2520_
	);
	LUT3 #(
		.INIT('h45)
	) name1518 (
		_w2518_,
		_w2519_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h1)
	) name1519 (
		_w2459_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('h8)
	) name1520 (
		_w2459_,
		_w2521_,
		_w2523_
	);
	LUT2 #(
		.INIT('h6)
	) name1521 (
		_w2418_,
		_w2446_,
		_w2524_
	);
	LUT4 #(
		.INIT('h6665)
	) name1522 (
		_w2482_,
		_w2507_,
		_w2508_,
		_w2517_,
		_w2525_
	);
	LUT4 #(
		.INIT('h1248)
	) name1523 (
		_w2458_,
		_w2520_,
		_w2524_,
		_w2525_,
		_w2526_
	);
	LUT4 #(
		.INIT('h8421)
	) name1524 (
		_w2458_,
		_w2520_,
		_w2524_,
		_w2525_,
		_w2527_
	);
	LUT3 #(
		.INIT('h96)
	) name1525 (
		_w2449_,
		_w2451_,
		_w2457_,
		_w2528_
	);
	LUT2 #(
		.INIT('h6)
	) name1526 (
		_w2483_,
		_w2506_,
		_w2529_
	);
	LUT2 #(
		.INIT('h9)
	) name1527 (
		_w2517_,
		_w2529_,
		_w2530_
	);
	LUT4 #(
		.INIT('h0660)
	) name1528 (
		_w2452_,
		_w2453_,
		_w2509_,
		_w2510_,
		_w2531_
	);
	LUT4 #(
		.INIT('h9600)
	) name1529 (
		_w2454_,
		_w2455_,
		_w2456_,
		_w2531_,
		_w2532_
	);
	LUT4 #(
		.INIT('h0069)
	) name1530 (
		_w2454_,
		_w2455_,
		_w2456_,
		_w2531_,
		_w2533_
	);
	LUT3 #(
		.INIT('h96)
	) name1531 (
		_w2474_,
		_w2511_,
		_w2512_,
		_w2534_
	);
	LUT2 #(
		.INIT('h9)
	) name1532 (
		_w2516_,
		_w2534_,
		_w2535_
	);
	LUT3 #(
		.INIT('h45)
	) name1533 (
		_w2532_,
		_w2533_,
		_w2535_,
		_w2536_
	);
	LUT3 #(
		.INIT('h71)
	) name1534 (
		_w2528_,
		_w2530_,
		_w2536_,
		_w2537_
	);
	LUT3 #(
		.INIT('h54)
	) name1535 (
		_w2526_,
		_w2527_,
		_w2537_,
		_w2538_
	);
	LUT3 #(
		.INIT('h54)
	) name1536 (
		_w2522_,
		_w2523_,
		_w2538_,
		_w2539_
	);
	LUT3 #(
		.INIT('h17)
	) name1537 (
		\A[259] ,
		\A[260] ,
		\A[261] ,
		_w2540_
	);
	LUT2 #(
		.INIT('h8)
	) name1538 (
		\A[262] ,
		\A[263] ,
		_w2541_
	);
	LUT3 #(
		.INIT('h96)
	) name1539 (
		\A[259] ,
		\A[260] ,
		\A[261] ,
		_w2542_
	);
	LUT3 #(
		.INIT('h96)
	) name1540 (
		\A[262] ,
		\A[263] ,
		\A[264] ,
		_w2543_
	);
	LUT3 #(
		.INIT('h80)
	) name1541 (
		_w2541_,
		_w2542_,
		_w2543_,
		_w2544_
	);
	LUT3 #(
		.INIT('h17)
	) name1542 (
		\A[262] ,
		\A[263] ,
		\A[264] ,
		_w2545_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1543 (
		\A[262] ,
		\A[263] ,
		\A[264] ,
		_w2542_,
		_w2546_
	);
	LUT2 #(
		.INIT('h9)
	) name1544 (
		_w2540_,
		_w2546_,
		_w2547_
	);
	LUT3 #(
		.INIT('h96)
	) name1545 (
		\A[265] ,
		\A[266] ,
		\A[267] ,
		_w2548_
	);
	LUT2 #(
		.INIT('h8)
	) name1546 (
		\A[268] ,
		\A[269] ,
		_w2549_
	);
	LUT3 #(
		.INIT('h96)
	) name1547 (
		\A[268] ,
		\A[269] ,
		\A[270] ,
		_w2550_
	);
	LUT3 #(
		.INIT('h17)
	) name1548 (
		\A[268] ,
		\A[269] ,
		\A[270] ,
		_w2551_
	);
	LUT3 #(
		.INIT('h17)
	) name1549 (
		\A[265] ,
		\A[266] ,
		\A[267] ,
		_w2552_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		_w2551_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h6)
	) name1551 (
		_w2551_,
		_w2552_,
		_w2554_
	);
	LUT4 #(
		.INIT('h8008)
	) name1552 (
		_w2548_,
		_w2550_,
		_w2551_,
		_w2552_,
		_w2555_
	);
	LUT4 #(
		.INIT('h0770)
	) name1553 (
		_w2548_,
		_w2550_,
		_w2551_,
		_w2552_,
		_w2556_
	);
	LUT4 #(
		.INIT('h0660)
	) name1554 (
		_w2542_,
		_w2543_,
		_w2548_,
		_w2550_,
		_w2557_
	);
	LUT3 #(
		.INIT('h01)
	) name1555 (
		_w2556_,
		_w2557_,
		_w2555_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name1556 (
		_w2554_,
		_w2557_,
		_w2559_
	);
	LUT4 #(
		.INIT('h4000)
	) name1557 (
		_w2540_,
		_w2541_,
		_w2542_,
		_w2543_,
		_w2560_
	);
	LUT3 #(
		.INIT('h08)
	) name1558 (
		_w2554_,
		_w2557_,
		_w2560_,
		_w2561_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1559 (
		_w2548_,
		_w2549_,
		_w2550_,
		_w2552_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w2553_,
		_w2562_,
		_w2563_
	);
	LUT4 #(
		.INIT('h00f2)
	) name1561 (
		_w2547_,
		_w2558_,
		_w2561_,
		_w2563_,
		_w2564_
	);
	LUT4 #(
		.INIT('h4055)
	) name1562 (
		_w2540_,
		_w2542_,
		_w2543_,
		_w2545_,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name1563 (
		_w2544_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1564 (
		_w2547_,
		_w2558_,
		_w2561_,
		_w2563_,
		_w2567_
	);
	LUT3 #(
		.INIT('h54)
	) name1565 (
		_w2564_,
		_w2566_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('h96)
	) name1566 (
		\A[253] ,
		\A[254] ,
		\A[255] ,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name1567 (
		\A[256] ,
		\A[257] ,
		_w2570_
	);
	LUT3 #(
		.INIT('h96)
	) name1568 (
		\A[256] ,
		\A[257] ,
		\A[258] ,
		_w2571_
	);
	LUT3 #(
		.INIT('h96)
	) name1569 (
		\A[247] ,
		\A[248] ,
		\A[249] ,
		_w2572_
	);
	LUT2 #(
		.INIT('h8)
	) name1570 (
		\A[250] ,
		\A[251] ,
		_w2573_
	);
	LUT3 #(
		.INIT('h96)
	) name1571 (
		\A[250] ,
		\A[251] ,
		\A[252] ,
		_w2574_
	);
	LUT4 #(
		.INIT('h0660)
	) name1572 (
		_w2569_,
		_w2571_,
		_w2572_,
		_w2574_,
		_w2575_
	);
	LUT3 #(
		.INIT('h17)
	) name1573 (
		\A[253] ,
		\A[254] ,
		\A[255] ,
		_w2576_
	);
	LUT3 #(
		.INIT('h17)
	) name1574 (
		\A[256] ,
		\A[257] ,
		\A[258] ,
		_w2577_
	);
	LUT3 #(
		.INIT('h80)
	) name1575 (
		_w2569_,
		_w2570_,
		_w2571_,
		_w2578_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1576 (
		\A[256] ,
		\A[257] ,
		\A[258] ,
		_w2569_,
		_w2579_
	);
	LUT2 #(
		.INIT('h9)
	) name1577 (
		_w2576_,
		_w2579_,
		_w2580_
	);
	LUT3 #(
		.INIT('h14)
	) name1578 (
		_w2575_,
		_w2576_,
		_w2579_,
		_w2581_
	);
	LUT3 #(
		.INIT('h17)
	) name1579 (
		\A[247] ,
		\A[248] ,
		\A[249] ,
		_w2582_
	);
	LUT3 #(
		.INIT('h80)
	) name1580 (
		_w2572_,
		_w2573_,
		_w2574_,
		_w2583_
	);
	LUT3 #(
		.INIT('h17)
	) name1581 (
		\A[250] ,
		\A[251] ,
		\A[252] ,
		_w2584_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1582 (
		\A[250] ,
		\A[251] ,
		\A[252] ,
		_w2572_,
		_w2585_
	);
	LUT2 #(
		.INIT('h9)
	) name1583 (
		_w2582_,
		_w2585_,
		_w2586_
	);
	LUT3 #(
		.INIT('h82)
	) name1584 (
		_w2575_,
		_w2576_,
		_w2579_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		_w2576_,
		_w2577_,
		_w2588_
	);
	LUT4 #(
		.INIT('h0080)
	) name1586 (
		_w2572_,
		_w2573_,
		_w2574_,
		_w2582_,
		_w2589_
	);
	LUT2 #(
		.INIT('h1)
	) name1587 (
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT4 #(
		.INIT('h171f)
	) name1588 (
		_w2575_,
		_w2580_,
		_w2586_,
		_w2590_,
		_w2591_
	);
	LUT4 #(
		.INIT('h080f)
	) name1589 (
		_w2569_,
		_w2571_,
		_w2576_,
		_w2577_,
		_w2592_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w2578_,
		_w2592_,
		_w2593_
	);
	LUT4 #(
		.INIT('h080f)
	) name1591 (
		_w2572_,
		_w2574_,
		_w2582_,
		_w2584_,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name1592 (
		_w2583_,
		_w2594_,
		_w2595_
	);
	LUT3 #(
		.INIT('he8)
	) name1593 (
		_w2591_,
		_w2593_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name1594 (
		_w2568_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h8)
	) name1595 (
		_w2568_,
		_w2596_,
		_w2598_
	);
	LUT3 #(
		.INIT('h69)
	) name1596 (
		_w2591_,
		_w2593_,
		_w2595_,
		_w2599_
	);
	LUT4 #(
		.INIT('hf20d)
	) name1597 (
		_w2547_,
		_w2558_,
		_w2561_,
		_w2563_,
		_w2600_
	);
	LUT2 #(
		.INIT('h9)
	) name1598 (
		_w2566_,
		_w2600_,
		_w2601_
	);
	LUT4 #(
		.INIT('h6996)
	) name1599 (
		_w2542_,
		_w2543_,
		_w2548_,
		_w2550_,
		_w2602_
	);
	LUT4 #(
		.INIT('h6996)
	) name1600 (
		_w2569_,
		_w2571_,
		_w2572_,
		_w2574_,
		_w2603_
	);
	LUT2 #(
		.INIT('h8)
	) name1601 (
		_w2602_,
		_w2603_,
		_w2604_
	);
	LUT4 #(
		.INIT('h89a9)
	) name1602 (
		_w2547_,
		_w2558_,
		_w2559_,
		_w2560_,
		_w2605_
	);
	LUT4 #(
		.INIT('hc989)
	) name1603 (
		_w2581_,
		_w2586_,
		_w2587_,
		_w2590_,
		_w2606_
	);
	LUT3 #(
		.INIT('he8)
	) name1604 (
		_w2604_,
		_w2605_,
		_w2606_,
		_w2607_
	);
	LUT3 #(
		.INIT('he8)
	) name1605 (
		_w2599_,
		_w2601_,
		_w2607_,
		_w2608_
	);
	LUT3 #(
		.INIT('h45)
	) name1606 (
		_w2597_,
		_w2598_,
		_w2608_,
		_w2609_
	);
	LUT3 #(
		.INIT('h17)
	) name1607 (
		\A[235] ,
		\A[236] ,
		\A[237] ,
		_w2610_
	);
	LUT2 #(
		.INIT('h8)
	) name1608 (
		\A[238] ,
		\A[239] ,
		_w2611_
	);
	LUT3 #(
		.INIT('h96)
	) name1609 (
		\A[235] ,
		\A[236] ,
		\A[237] ,
		_w2612_
	);
	LUT3 #(
		.INIT('h96)
	) name1610 (
		\A[238] ,
		\A[239] ,
		\A[240] ,
		_w2613_
	);
	LUT3 #(
		.INIT('h80)
	) name1611 (
		_w2611_,
		_w2612_,
		_w2613_,
		_w2614_
	);
	LUT3 #(
		.INIT('h17)
	) name1612 (
		\A[238] ,
		\A[239] ,
		\A[240] ,
		_w2615_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1613 (
		\A[238] ,
		\A[239] ,
		\A[240] ,
		_w2612_,
		_w2616_
	);
	LUT2 #(
		.INIT('h9)
	) name1614 (
		_w2610_,
		_w2616_,
		_w2617_
	);
	LUT3 #(
		.INIT('h96)
	) name1615 (
		\A[241] ,
		\A[242] ,
		\A[243] ,
		_w2618_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		\A[244] ,
		\A[245] ,
		_w2619_
	);
	LUT3 #(
		.INIT('h96)
	) name1617 (
		\A[244] ,
		\A[245] ,
		\A[246] ,
		_w2620_
	);
	LUT3 #(
		.INIT('h17)
	) name1618 (
		\A[244] ,
		\A[245] ,
		\A[246] ,
		_w2621_
	);
	LUT3 #(
		.INIT('h17)
	) name1619 (
		\A[241] ,
		\A[242] ,
		\A[243] ,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w2621_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h6)
	) name1621 (
		_w2621_,
		_w2622_,
		_w2624_
	);
	LUT4 #(
		.INIT('h8008)
	) name1622 (
		_w2618_,
		_w2620_,
		_w2621_,
		_w2622_,
		_w2625_
	);
	LUT4 #(
		.INIT('h0770)
	) name1623 (
		_w2618_,
		_w2620_,
		_w2621_,
		_w2622_,
		_w2626_
	);
	LUT4 #(
		.INIT('h0660)
	) name1624 (
		_w2612_,
		_w2613_,
		_w2618_,
		_w2620_,
		_w2627_
	);
	LUT3 #(
		.INIT('h01)
	) name1625 (
		_w2626_,
		_w2627_,
		_w2625_,
		_w2628_
	);
	LUT2 #(
		.INIT('h8)
	) name1626 (
		_w2624_,
		_w2627_,
		_w2629_
	);
	LUT4 #(
		.INIT('h4000)
	) name1627 (
		_w2610_,
		_w2611_,
		_w2612_,
		_w2613_,
		_w2630_
	);
	LUT3 #(
		.INIT('h08)
	) name1628 (
		_w2624_,
		_w2627_,
		_w2630_,
		_w2631_
	);
	LUT3 #(
		.INIT('h0d)
	) name1629 (
		_w2617_,
		_w2628_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1630 (
		_w2618_,
		_w2619_,
		_w2620_,
		_w2622_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w2623_,
		_w2633_,
		_w2634_
	);
	LUT4 #(
		.INIT('h00f2)
	) name1632 (
		_w2617_,
		_w2628_,
		_w2631_,
		_w2634_,
		_w2635_
	);
	LUT4 #(
		.INIT('h4055)
	) name1633 (
		_w2610_,
		_w2612_,
		_w2613_,
		_w2615_,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name1634 (
		_w2614_,
		_w2636_,
		_w2637_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1635 (
		_w2617_,
		_w2628_,
		_w2631_,
		_w2634_,
		_w2638_
	);
	LUT3 #(
		.INIT('h96)
	) name1636 (
		\A[229] ,
		\A[230] ,
		\A[231] ,
		_w2639_
	);
	LUT3 #(
		.INIT('h96)
	) name1637 (
		\A[232] ,
		\A[233] ,
		\A[234] ,
		_w2640_
	);
	LUT2 #(
		.INIT('h8)
	) name1638 (
		_w2639_,
		_w2640_,
		_w2641_
	);
	LUT3 #(
		.INIT('h96)
	) name1639 (
		\A[223] ,
		\A[224] ,
		\A[225] ,
		_w2642_
	);
	LUT3 #(
		.INIT('h96)
	) name1640 (
		\A[226] ,
		\A[227] ,
		\A[228] ,
		_w2643_
	);
	LUT4 #(
		.INIT('h0660)
	) name1641 (
		_w2639_,
		_w2640_,
		_w2642_,
		_w2643_,
		_w2644_
	);
	LUT3 #(
		.INIT('h17)
	) name1642 (
		\A[232] ,
		\A[233] ,
		\A[234] ,
		_w2645_
	);
	LUT3 #(
		.INIT('h17)
	) name1643 (
		\A[229] ,
		\A[230] ,
		\A[231] ,
		_w2646_
	);
	LUT2 #(
		.INIT('h6)
	) name1644 (
		_w2645_,
		_w2646_,
		_w2647_
	);
	LUT3 #(
		.INIT('h17)
	) name1645 (
		\A[226] ,
		\A[227] ,
		\A[228] ,
		_w2648_
	);
	LUT3 #(
		.INIT('h17)
	) name1646 (
		\A[223] ,
		\A[224] ,
		\A[225] ,
		_w2649_
	);
	LUT4 #(
		.INIT('h7887)
	) name1647 (
		_w2642_,
		_w2643_,
		_w2648_,
		_w2649_,
		_w2650_
	);
	LUT4 #(
		.INIT('hc0de)
	) name1648 (
		_w2641_,
		_w2644_,
		_w2647_,
		_w2650_,
		_w2651_
	);
	LUT4 #(
		.INIT('h088f)
	) name1649 (
		_w2639_,
		_w2640_,
		_w2645_,
		_w2646_,
		_w2652_
	);
	LUT4 #(
		.INIT('h088f)
	) name1650 (
		_w2642_,
		_w2643_,
		_w2648_,
		_w2649_,
		_w2653_
	);
	LUT3 #(
		.INIT('he8)
	) name1651 (
		_w2651_,
		_w2652_,
		_w2653_,
		_w2654_
	);
	LUT4 #(
		.INIT('h1700)
	) name1652 (
		_w2632_,
		_w2634_,
		_w2637_,
		_w2654_,
		_w2655_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1653 (
		_w2632_,
		_w2634_,
		_w2637_,
		_w2654_,
		_w2656_
	);
	LUT4 #(
		.INIT('hf20d)
	) name1654 (
		_w2617_,
		_w2628_,
		_w2631_,
		_w2634_,
		_w2657_
	);
	LUT3 #(
		.INIT('h69)
	) name1655 (
		_w2651_,
		_w2652_,
		_w2653_,
		_w2658_
	);
	LUT3 #(
		.INIT('h09)
	) name1656 (
		_w2637_,
		_w2657_,
		_w2658_,
		_w2659_
	);
	LUT3 #(
		.INIT('h60)
	) name1657 (
		_w2637_,
		_w2657_,
		_w2658_,
		_w2660_
	);
	LUT4 #(
		.INIT('h6996)
	) name1658 (
		_w2612_,
		_w2613_,
		_w2618_,
		_w2620_,
		_w2661_
	);
	LUT4 #(
		.INIT('h6996)
	) name1659 (
		_w2639_,
		_w2640_,
		_w2642_,
		_w2643_,
		_w2662_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT4 #(
		.INIT('h89a9)
	) name1661 (
		_w2617_,
		_w2628_,
		_w2629_,
		_w2630_,
		_w2664_
	);
	LUT4 #(
		.INIT('he11e)
	) name1662 (
		_w2641_,
		_w2644_,
		_w2647_,
		_w2650_,
		_w2665_
	);
	LUT3 #(
		.INIT('h71)
	) name1663 (
		_w2663_,
		_w2664_,
		_w2665_,
		_w2666_
	);
	LUT4 #(
		.INIT('h4445)
	) name1664 (
		_w2656_,
		_w2659_,
		_w2660_,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		_w2655_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h1)
	) name1666 (
		_w2609_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h8)
	) name1667 (
		_w2609_,
		_w2668_,
		_w2670_
	);
	LUT2 #(
		.INIT('h6)
	) name1668 (
		_w2568_,
		_w2596_,
		_w2671_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1669 (
		_w2635_,
		_w2637_,
		_w2638_,
		_w2654_,
		_w2672_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1670 (
		_w2659_,
		_w2660_,
		_w2666_,
		_w2672_,
		_w2673_
	);
	LUT3 #(
		.INIT('h09)
	) name1671 (
		_w2608_,
		_w2671_,
		_w2673_,
		_w2674_
	);
	LUT3 #(
		.INIT('h60)
	) name1672 (
		_w2608_,
		_w2671_,
		_w2673_,
		_w2675_
	);
	LUT3 #(
		.INIT('h96)
	) name1673 (
		_w2599_,
		_w2601_,
		_w2607_,
		_w2676_
	);
	LUT3 #(
		.INIT('h96)
	) name1674 (
		_w2637_,
		_w2657_,
		_w2658_,
		_w2677_
	);
	LUT2 #(
		.INIT('h9)
	) name1675 (
		_w2666_,
		_w2677_,
		_w2678_
	);
	LUT4 #(
		.INIT('h0660)
	) name1676 (
		_w2602_,
		_w2603_,
		_w2661_,
		_w2662_,
		_w2679_
	);
	LUT4 #(
		.INIT('h9600)
	) name1677 (
		_w2604_,
		_w2605_,
		_w2606_,
		_w2679_,
		_w2680_
	);
	LUT4 #(
		.INIT('h0069)
	) name1678 (
		_w2604_,
		_w2605_,
		_w2606_,
		_w2679_,
		_w2681_
	);
	LUT3 #(
		.INIT('h69)
	) name1679 (
		_w2663_,
		_w2664_,
		_w2665_,
		_w2682_
	);
	LUT3 #(
		.INIT('h45)
	) name1680 (
		_w2680_,
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT3 #(
		.INIT('h71)
	) name1681 (
		_w2676_,
		_w2678_,
		_w2683_,
		_w2684_
	);
	LUT3 #(
		.INIT('h45)
	) name1682 (
		_w2674_,
		_w2675_,
		_w2684_,
		_w2685_
	);
	LUT3 #(
		.INIT('h45)
	) name1683 (
		_w2669_,
		_w2670_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w2539_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h8)
	) name1685 (
		_w2539_,
		_w2686_,
		_w2688_
	);
	LUT2 #(
		.INIT('h6)
	) name1686 (
		_w2609_,
		_w2668_,
		_w2689_
	);
	LUT2 #(
		.INIT('h6)
	) name1687 (
		_w2459_,
		_w2521_,
		_w2690_
	);
	LUT4 #(
		.INIT('h4182)
	) name1688 (
		_w2538_,
		_w2685_,
		_w2689_,
		_w2690_,
		_w2691_
	);
	LUT4 #(
		.INIT('h2814)
	) name1689 (
		_w2538_,
		_w2685_,
		_w2689_,
		_w2690_,
		_w2692_
	);
	LUT4 #(
		.INIT('h6996)
	) name1690 (
		_w2458_,
		_w2520_,
		_w2524_,
		_w2525_,
		_w2693_
	);
	LUT3 #(
		.INIT('h96)
	) name1691 (
		_w2608_,
		_w2671_,
		_w2673_,
		_w2694_
	);
	LUT4 #(
		.INIT('h1248)
	) name1692 (
		_w2537_,
		_w2684_,
		_w2693_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h8421)
	) name1693 (
		_w2537_,
		_w2684_,
		_w2693_,
		_w2694_,
		_w2696_
	);
	LUT3 #(
		.INIT('h69)
	) name1694 (
		_w2528_,
		_w2530_,
		_w2536_,
		_w2697_
	);
	LUT3 #(
		.INIT('h69)
	) name1695 (
		_w2676_,
		_w2678_,
		_w2683_,
		_w2698_
	);
	LUT4 #(
		.INIT('h6996)
	) name1696 (
		_w2602_,
		_w2603_,
		_w2661_,
		_w2662_,
		_w2699_
	);
	LUT4 #(
		.INIT('h6996)
	) name1697 (
		_w2452_,
		_w2453_,
		_w2509_,
		_w2510_,
		_w2700_
	);
	LUT2 #(
		.INIT('h8)
	) name1698 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT4 #(
		.INIT('h6996)
	) name1699 (
		_w2604_,
		_w2605_,
		_w2606_,
		_w2679_,
		_w2702_
	);
	LUT3 #(
		.INIT('h48)
	) name1700 (
		_w2682_,
		_w2701_,
		_w2702_,
		_w2703_
	);
	LUT3 #(
		.INIT('h21)
	) name1701 (
		_w2682_,
		_w2701_,
		_w2702_,
		_w2704_
	);
	LUT4 #(
		.INIT('h6996)
	) name1702 (
		_w2454_,
		_w2455_,
		_w2456_,
		_w2531_,
		_w2705_
	);
	LUT2 #(
		.INIT('h9)
	) name1703 (
		_w2535_,
		_w2705_,
		_w2706_
	);
	LUT3 #(
		.INIT('h54)
	) name1704 (
		_w2703_,
		_w2704_,
		_w2706_,
		_w2707_
	);
	LUT3 #(
		.INIT('h8e)
	) name1705 (
		_w2697_,
		_w2698_,
		_w2707_,
		_w2708_
	);
	LUT3 #(
		.INIT('h54)
	) name1706 (
		_w2695_,
		_w2696_,
		_w2708_,
		_w2709_
	);
	LUT3 #(
		.INIT('h54)
	) name1707 (
		_w2691_,
		_w2692_,
		_w2709_,
		_w2710_
	);
	LUT3 #(
		.INIT('h45)
	) name1708 (
		_w2687_,
		_w2688_,
		_w2710_,
		_w2711_
	);
	LUT3 #(
		.INIT('h96)
	) name1709 (
		\A[145] ,
		\A[146] ,
		\A[147] ,
		_w2712_
	);
	LUT3 #(
		.INIT('h96)
	) name1710 (
		\A[148] ,
		\A[149] ,
		\A[150] ,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		_w2712_,
		_w2713_,
		_w2714_
	);
	LUT3 #(
		.INIT('h96)
	) name1712 (
		\A[139] ,
		\A[140] ,
		\A[141] ,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name1713 (
		\A[142] ,
		\A[143] ,
		_w2716_
	);
	LUT3 #(
		.INIT('h96)
	) name1714 (
		\A[142] ,
		\A[143] ,
		\A[144] ,
		_w2717_
	);
	LUT4 #(
		.INIT('h0660)
	) name1715 (
		_w2712_,
		_w2713_,
		_w2715_,
		_w2717_,
		_w2718_
	);
	LUT3 #(
		.INIT('h17)
	) name1716 (
		\A[148] ,
		\A[149] ,
		\A[150] ,
		_w2719_
	);
	LUT3 #(
		.INIT('h17)
	) name1717 (
		\A[145] ,
		\A[146] ,
		\A[147] ,
		_w2720_
	);
	LUT2 #(
		.INIT('h6)
	) name1718 (
		_w2719_,
		_w2720_,
		_w2721_
	);
	LUT3 #(
		.INIT('h17)
	) name1719 (
		\A[139] ,
		\A[140] ,
		\A[141] ,
		_w2722_
	);
	LUT3 #(
		.INIT('h17)
	) name1720 (
		\A[142] ,
		\A[143] ,
		\A[144] ,
		_w2723_
	);
	LUT3 #(
		.INIT('h80)
	) name1721 (
		_w2715_,
		_w2716_,
		_w2717_,
		_w2724_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1722 (
		\A[142] ,
		\A[143] ,
		\A[144] ,
		_w2715_,
		_w2725_
	);
	LUT2 #(
		.INIT('h9)
	) name1723 (
		_w2722_,
		_w2725_,
		_w2726_
	);
	LUT4 #(
		.INIT('h0770)
	) name1724 (
		_w2718_,
		_w2721_,
		_w2722_,
		_w2725_,
		_w2727_
	);
	LUT4 #(
		.INIT('h8008)
	) name1725 (
		_w2712_,
		_w2713_,
		_w2719_,
		_w2720_,
		_w2728_
	);
	LUT4 #(
		.INIT('h0770)
	) name1726 (
		_w2712_,
		_w2713_,
		_w2719_,
		_w2720_,
		_w2729_
	);
	LUT3 #(
		.INIT('h01)
	) name1727 (
		_w2718_,
		_w2729_,
		_w2728_,
		_w2730_
	);
	LUT4 #(
		.INIT('h088f)
	) name1728 (
		_w2712_,
		_w2713_,
		_w2719_,
		_w2720_,
		_w2731_
	);
	LUT4 #(
		.INIT('h080f)
	) name1729 (
		_w2715_,
		_w2717_,
		_w2722_,
		_w2723_,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name1730 (
		_w2724_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h10f1)
	) name1731 (
		_w2727_,
		_w2730_,
		_w2731_,
		_w2733_,
		_w2734_
	);
	LUT4 #(
		.INIT('he11e)
	) name1732 (
		_w2727_,
		_w2730_,
		_w2731_,
		_w2733_,
		_w2735_
	);
	LUT2 #(
		.INIT('h8)
	) name1733 (
		\A[130] ,
		\A[131] ,
		_w2736_
	);
	LUT3 #(
		.INIT('h96)
	) name1734 (
		\A[127] ,
		\A[128] ,
		\A[129] ,
		_w2737_
	);
	LUT3 #(
		.INIT('h96)
	) name1735 (
		\A[130] ,
		\A[131] ,
		\A[132] ,
		_w2738_
	);
	LUT3 #(
		.INIT('h80)
	) name1736 (
		_w2736_,
		_w2737_,
		_w2738_,
		_w2739_
	);
	LUT3 #(
		.INIT('h17)
	) name1737 (
		\A[127] ,
		\A[128] ,
		\A[129] ,
		_w2740_
	);
	LUT3 #(
		.INIT('h17)
	) name1738 (
		\A[130] ,
		\A[131] ,
		\A[132] ,
		_w2741_
	);
	LUT4 #(
		.INIT('h080f)
	) name1739 (
		_w2737_,
		_w2738_,
		_w2740_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w2739_,
		_w2742_,
		_w2743_
	);
	LUT3 #(
		.INIT('h96)
	) name1741 (
		\A[133] ,
		\A[134] ,
		\A[135] ,
		_w2744_
	);
	LUT3 #(
		.INIT('h96)
	) name1742 (
		\A[136] ,
		\A[137] ,
		\A[138] ,
		_w2745_
	);
	LUT2 #(
		.INIT('h8)
	) name1743 (
		_w2744_,
		_w2745_,
		_w2746_
	);
	LUT4 #(
		.INIT('h0660)
	) name1744 (
		_w2737_,
		_w2738_,
		_w2744_,
		_w2745_,
		_w2747_
	);
	LUT3 #(
		.INIT('h17)
	) name1745 (
		\A[136] ,
		\A[137] ,
		\A[138] ,
		_w2748_
	);
	LUT3 #(
		.INIT('h17)
	) name1746 (
		\A[133] ,
		\A[134] ,
		\A[135] ,
		_w2749_
	);
	LUT2 #(
		.INIT('h6)
	) name1747 (
		_w2748_,
		_w2749_,
		_w2750_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1748 (
		\A[130] ,
		\A[131] ,
		\A[132] ,
		_w2737_,
		_w2751_
	);
	LUT2 #(
		.INIT('h9)
	) name1749 (
		_w2740_,
		_w2751_,
		_w2752_
	);
	LUT4 #(
		.INIT('h152a)
	) name1750 (
		_w2740_,
		_w2747_,
		_w2750_,
		_w2751_,
		_w2753_
	);
	LUT4 #(
		.INIT('h8008)
	) name1751 (
		_w2744_,
		_w2745_,
		_w2748_,
		_w2749_,
		_w2754_
	);
	LUT4 #(
		.INIT('h0770)
	) name1752 (
		_w2744_,
		_w2745_,
		_w2748_,
		_w2749_,
		_w2755_
	);
	LUT3 #(
		.INIT('h01)
	) name1753 (
		_w2747_,
		_w2755_,
		_w2754_,
		_w2756_
	);
	LUT4 #(
		.INIT('h088f)
	) name1754 (
		_w2744_,
		_w2745_,
		_w2748_,
		_w2749_,
		_w2757_
	);
	LUT4 #(
		.INIT('ha956)
	) name1755 (
		_w2743_,
		_w2753_,
		_w2756_,
		_w2757_,
		_w2758_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		_w2735_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w2735_,
		_w2758_,
		_w2760_
	);
	LUT4 #(
		.INIT('h6996)
	) name1758 (
		_w2712_,
		_w2713_,
		_w2715_,
		_w2717_,
		_w2761_
	);
	LUT4 #(
		.INIT('h6996)
	) name1759 (
		_w2737_,
		_w2738_,
		_w2744_,
		_w2745_,
		_w2762_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		_w2761_,
		_w2762_,
		_w2763_
	);
	LUT3 #(
		.INIT('h1e)
	) name1761 (
		_w2714_,
		_w2718_,
		_w2721_,
		_w2764_
	);
	LUT3 #(
		.INIT('h48)
	) name1762 (
		_w2726_,
		_w2763_,
		_w2764_,
		_w2765_
	);
	LUT3 #(
		.INIT('h21)
	) name1763 (
		_w2726_,
		_w2763_,
		_w2764_,
		_w2766_
	);
	LUT3 #(
		.INIT('h1e)
	) name1764 (
		_w2746_,
		_w2747_,
		_w2750_,
		_w2767_
	);
	LUT2 #(
		.INIT('h9)
	) name1765 (
		_w2752_,
		_w2767_,
		_w2768_
	);
	LUT3 #(
		.INIT('h54)
	) name1766 (
		_w2765_,
		_w2766_,
		_w2768_,
		_w2769_
	);
	LUT4 #(
		.INIT('h1501)
	) name1767 (
		_w2734_,
		_w2735_,
		_w2758_,
		_w2769_,
		_w2770_
	);
	LUT4 #(
		.INIT('h80a8)
	) name1768 (
		_w2734_,
		_w2735_,
		_w2758_,
		_w2769_,
		_w2771_
	);
	LUT4 #(
		.INIT('h5701)
	) name1769 (
		_w2743_,
		_w2753_,
		_w2756_,
		_w2757_,
		_w2772_
	);
	LUT3 #(
		.INIT('h54)
	) name1770 (
		_w2770_,
		_w2771_,
		_w2772_,
		_w2773_
	);
	LUT3 #(
		.INIT('h96)
	) name1771 (
		\A[169] ,
		\A[170] ,
		\A[171] ,
		_w2774_
	);
	LUT3 #(
		.INIT('h96)
	) name1772 (
		\A[172] ,
		\A[173] ,
		\A[174] ,
		_w2775_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		_w2774_,
		_w2775_,
		_w2776_
	);
	LUT3 #(
		.INIT('h96)
	) name1774 (
		\A[163] ,
		\A[164] ,
		\A[165] ,
		_w2777_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		\A[166] ,
		\A[167] ,
		_w2778_
	);
	LUT3 #(
		.INIT('h96)
	) name1776 (
		\A[166] ,
		\A[167] ,
		\A[168] ,
		_w2779_
	);
	LUT4 #(
		.INIT('h0660)
	) name1777 (
		_w2774_,
		_w2775_,
		_w2777_,
		_w2779_,
		_w2780_
	);
	LUT3 #(
		.INIT('h17)
	) name1778 (
		\A[172] ,
		\A[173] ,
		\A[174] ,
		_w2781_
	);
	LUT3 #(
		.INIT('h17)
	) name1779 (
		\A[169] ,
		\A[170] ,
		\A[171] ,
		_w2782_
	);
	LUT2 #(
		.INIT('h6)
	) name1780 (
		_w2781_,
		_w2782_,
		_w2783_
	);
	LUT3 #(
		.INIT('h17)
	) name1781 (
		\A[163] ,
		\A[164] ,
		\A[165] ,
		_w2784_
	);
	LUT3 #(
		.INIT('h17)
	) name1782 (
		\A[166] ,
		\A[167] ,
		\A[168] ,
		_w2785_
	);
	LUT3 #(
		.INIT('h80)
	) name1783 (
		_w2777_,
		_w2778_,
		_w2779_,
		_w2786_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1784 (
		\A[166] ,
		\A[167] ,
		\A[168] ,
		_w2777_,
		_w2787_
	);
	LUT2 #(
		.INIT('h9)
	) name1785 (
		_w2784_,
		_w2787_,
		_w2788_
	);
	LUT4 #(
		.INIT('h0770)
	) name1786 (
		_w2780_,
		_w2783_,
		_w2784_,
		_w2787_,
		_w2789_
	);
	LUT4 #(
		.INIT('h8008)
	) name1787 (
		_w2774_,
		_w2775_,
		_w2781_,
		_w2782_,
		_w2790_
	);
	LUT4 #(
		.INIT('h0770)
	) name1788 (
		_w2774_,
		_w2775_,
		_w2781_,
		_w2782_,
		_w2791_
	);
	LUT3 #(
		.INIT('h01)
	) name1789 (
		_w2780_,
		_w2791_,
		_w2790_,
		_w2792_
	);
	LUT4 #(
		.INIT('h088f)
	) name1790 (
		_w2774_,
		_w2775_,
		_w2781_,
		_w2782_,
		_w2793_
	);
	LUT4 #(
		.INIT('h080f)
	) name1791 (
		_w2777_,
		_w2779_,
		_w2784_,
		_w2785_,
		_w2794_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w2786_,
		_w2794_,
		_w2795_
	);
	LUT4 #(
		.INIT('h10f1)
	) name1793 (
		_w2789_,
		_w2792_,
		_w2793_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('he11e)
	) name1794 (
		_w2789_,
		_w2792_,
		_w2793_,
		_w2795_,
		_w2797_
	);
	LUT2 #(
		.INIT('h8)
	) name1795 (
		\A[154] ,
		\A[155] ,
		_w2798_
	);
	LUT3 #(
		.INIT('h96)
	) name1796 (
		\A[151] ,
		\A[152] ,
		\A[153] ,
		_w2799_
	);
	LUT3 #(
		.INIT('h96)
	) name1797 (
		\A[154] ,
		\A[155] ,
		\A[156] ,
		_w2800_
	);
	LUT3 #(
		.INIT('h80)
	) name1798 (
		_w2798_,
		_w2799_,
		_w2800_,
		_w2801_
	);
	LUT3 #(
		.INIT('h17)
	) name1799 (
		\A[151] ,
		\A[152] ,
		\A[153] ,
		_w2802_
	);
	LUT3 #(
		.INIT('h17)
	) name1800 (
		\A[154] ,
		\A[155] ,
		\A[156] ,
		_w2803_
	);
	LUT4 #(
		.INIT('h080f)
	) name1801 (
		_w2799_,
		_w2800_,
		_w2802_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		_w2801_,
		_w2804_,
		_w2805_
	);
	LUT3 #(
		.INIT('h96)
	) name1803 (
		\A[157] ,
		\A[158] ,
		\A[159] ,
		_w2806_
	);
	LUT3 #(
		.INIT('h96)
	) name1804 (
		\A[160] ,
		\A[161] ,
		\A[162] ,
		_w2807_
	);
	LUT2 #(
		.INIT('h8)
	) name1805 (
		_w2806_,
		_w2807_,
		_w2808_
	);
	LUT4 #(
		.INIT('h0660)
	) name1806 (
		_w2799_,
		_w2800_,
		_w2806_,
		_w2807_,
		_w2809_
	);
	LUT3 #(
		.INIT('h17)
	) name1807 (
		\A[160] ,
		\A[161] ,
		\A[162] ,
		_w2810_
	);
	LUT3 #(
		.INIT('h17)
	) name1808 (
		\A[157] ,
		\A[158] ,
		\A[159] ,
		_w2811_
	);
	LUT2 #(
		.INIT('h6)
	) name1809 (
		_w2810_,
		_w2811_,
		_w2812_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1810 (
		\A[154] ,
		\A[155] ,
		\A[156] ,
		_w2799_,
		_w2813_
	);
	LUT2 #(
		.INIT('h9)
	) name1811 (
		_w2802_,
		_w2813_,
		_w2814_
	);
	LUT4 #(
		.INIT('h152a)
	) name1812 (
		_w2802_,
		_w2809_,
		_w2812_,
		_w2813_,
		_w2815_
	);
	LUT4 #(
		.INIT('h8008)
	) name1813 (
		_w2806_,
		_w2807_,
		_w2810_,
		_w2811_,
		_w2816_
	);
	LUT4 #(
		.INIT('h0770)
	) name1814 (
		_w2806_,
		_w2807_,
		_w2810_,
		_w2811_,
		_w2817_
	);
	LUT3 #(
		.INIT('h01)
	) name1815 (
		_w2809_,
		_w2817_,
		_w2816_,
		_w2818_
	);
	LUT4 #(
		.INIT('h088f)
	) name1816 (
		_w2806_,
		_w2807_,
		_w2810_,
		_w2811_,
		_w2819_
	);
	LUT4 #(
		.INIT('ha956)
	) name1817 (
		_w2805_,
		_w2815_,
		_w2818_,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		_w2797_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		_w2797_,
		_w2820_,
		_w2822_
	);
	LUT4 #(
		.INIT('h6996)
	) name1820 (
		_w2774_,
		_w2775_,
		_w2777_,
		_w2779_,
		_w2823_
	);
	LUT4 #(
		.INIT('h6996)
	) name1821 (
		_w2799_,
		_w2800_,
		_w2806_,
		_w2807_,
		_w2824_
	);
	LUT2 #(
		.INIT('h8)
	) name1822 (
		_w2823_,
		_w2824_,
		_w2825_
	);
	LUT3 #(
		.INIT('h1e)
	) name1823 (
		_w2776_,
		_w2780_,
		_w2783_,
		_w2826_
	);
	LUT3 #(
		.INIT('h48)
	) name1824 (
		_w2788_,
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT3 #(
		.INIT('h21)
	) name1825 (
		_w2788_,
		_w2825_,
		_w2826_,
		_w2828_
	);
	LUT3 #(
		.INIT('h1e)
	) name1826 (
		_w2808_,
		_w2809_,
		_w2812_,
		_w2829_
	);
	LUT2 #(
		.INIT('h9)
	) name1827 (
		_w2814_,
		_w2829_,
		_w2830_
	);
	LUT3 #(
		.INIT('h54)
	) name1828 (
		_w2827_,
		_w2828_,
		_w2830_,
		_w2831_
	);
	LUT4 #(
		.INIT('h1501)
	) name1829 (
		_w2796_,
		_w2797_,
		_w2820_,
		_w2831_,
		_w2832_
	);
	LUT4 #(
		.INIT('h80a8)
	) name1830 (
		_w2796_,
		_w2797_,
		_w2820_,
		_w2831_,
		_w2833_
	);
	LUT4 #(
		.INIT('h5701)
	) name1831 (
		_w2805_,
		_w2815_,
		_w2818_,
		_w2819_,
		_w2834_
	);
	LUT3 #(
		.INIT('h54)
	) name1832 (
		_w2832_,
		_w2833_,
		_w2834_,
		_w2835_
	);
	LUT2 #(
		.INIT('h1)
	) name1833 (
		_w2773_,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		_w2773_,
		_w2835_,
		_w2837_
	);
	LUT4 #(
		.INIT('h6665)
	) name1835 (
		_w2796_,
		_w2821_,
		_w2822_,
		_w2831_,
		_w2838_
	);
	LUT4 #(
		.INIT('h6665)
	) name1836 (
		_w2734_,
		_w2759_,
		_w2760_,
		_w2769_,
		_w2839_
	);
	LUT4 #(
		.INIT('h8241)
	) name1837 (
		_w2772_,
		_w2834_,
		_w2838_,
		_w2839_,
		_w2840_
	);
	LUT4 #(
		.INIT('h1428)
	) name1838 (
		_w2772_,
		_w2834_,
		_w2838_,
		_w2839_,
		_w2841_
	);
	LUT2 #(
		.INIT('h6)
	) name1839 (
		_w2735_,
		_w2758_,
		_w2842_
	);
	LUT2 #(
		.INIT('h6)
	) name1840 (
		_w2797_,
		_w2820_,
		_w2843_
	);
	LUT4 #(
		.INIT('h1248)
	) name1841 (
		_w2769_,
		_w2831_,
		_w2842_,
		_w2843_,
		_w2844_
	);
	LUT4 #(
		.INIT('h8421)
	) name1842 (
		_w2769_,
		_w2831_,
		_w2842_,
		_w2843_,
		_w2845_
	);
	LUT4 #(
		.INIT('h0660)
	) name1843 (
		_w2761_,
		_w2762_,
		_w2823_,
		_w2824_,
		_w2846_
	);
	LUT3 #(
		.INIT('h96)
	) name1844 (
		_w2788_,
		_w2825_,
		_w2826_,
		_w2847_
	);
	LUT3 #(
		.INIT('h84)
	) name1845 (
		_w2830_,
		_w2846_,
		_w2847_,
		_w2848_
	);
	LUT3 #(
		.INIT('h12)
	) name1846 (
		_w2830_,
		_w2846_,
		_w2847_,
		_w2849_
	);
	LUT3 #(
		.INIT('h96)
	) name1847 (
		_w2726_,
		_w2763_,
		_w2764_,
		_w2850_
	);
	LUT2 #(
		.INIT('h9)
	) name1848 (
		_w2768_,
		_w2850_,
		_w2851_
	);
	LUT3 #(
		.INIT('h45)
	) name1849 (
		_w2848_,
		_w2849_,
		_w2851_,
		_w2852_
	);
	LUT3 #(
		.INIT('h45)
	) name1850 (
		_w2844_,
		_w2845_,
		_w2852_,
		_w2853_
	);
	LUT3 #(
		.INIT('h54)
	) name1851 (
		_w2840_,
		_w2841_,
		_w2853_,
		_w2854_
	);
	LUT3 #(
		.INIT('h54)
	) name1852 (
		_w2836_,
		_w2837_,
		_w2854_,
		_w2855_
	);
	LUT3 #(
		.INIT('h96)
	) name1853 (
		\A[97] ,
		\A[98] ,
		\A[99] ,
		_w2856_
	);
	LUT3 #(
		.INIT('h96)
	) name1854 (
		\A[100] ,
		\A[101] ,
		\A[102] ,
		_w2857_
	);
	LUT2 #(
		.INIT('h8)
	) name1855 (
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT3 #(
		.INIT('h96)
	) name1856 (
		\A[91] ,
		\A[92] ,
		\A[93] ,
		_w2859_
	);
	LUT2 #(
		.INIT('h8)
	) name1857 (
		\A[94] ,
		\A[95] ,
		_w2860_
	);
	LUT3 #(
		.INIT('h96)
	) name1858 (
		\A[94] ,
		\A[95] ,
		\A[96] ,
		_w2861_
	);
	LUT4 #(
		.INIT('h0660)
	) name1859 (
		_w2856_,
		_w2857_,
		_w2859_,
		_w2861_,
		_w2862_
	);
	LUT3 #(
		.INIT('h17)
	) name1860 (
		\A[100] ,
		\A[101] ,
		\A[102] ,
		_w2863_
	);
	LUT3 #(
		.INIT('h17)
	) name1861 (
		\A[97] ,
		\A[98] ,
		\A[99] ,
		_w2864_
	);
	LUT2 #(
		.INIT('h6)
	) name1862 (
		_w2863_,
		_w2864_,
		_w2865_
	);
	LUT3 #(
		.INIT('h17)
	) name1863 (
		\A[91] ,
		\A[92] ,
		\A[93] ,
		_w2866_
	);
	LUT3 #(
		.INIT('h17)
	) name1864 (
		\A[94] ,
		\A[95] ,
		\A[96] ,
		_w2867_
	);
	LUT3 #(
		.INIT('h80)
	) name1865 (
		_w2859_,
		_w2860_,
		_w2861_,
		_w2868_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1866 (
		\A[94] ,
		\A[95] ,
		\A[96] ,
		_w2859_,
		_w2869_
	);
	LUT2 #(
		.INIT('h9)
	) name1867 (
		_w2866_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('h0770)
	) name1868 (
		_w2862_,
		_w2865_,
		_w2866_,
		_w2869_,
		_w2871_
	);
	LUT4 #(
		.INIT('h8008)
	) name1869 (
		_w2856_,
		_w2857_,
		_w2863_,
		_w2864_,
		_w2872_
	);
	LUT4 #(
		.INIT('h0770)
	) name1870 (
		_w2856_,
		_w2857_,
		_w2863_,
		_w2864_,
		_w2873_
	);
	LUT3 #(
		.INIT('h01)
	) name1871 (
		_w2862_,
		_w2873_,
		_w2872_,
		_w2874_
	);
	LUT4 #(
		.INIT('h088f)
	) name1872 (
		_w2856_,
		_w2857_,
		_w2863_,
		_w2864_,
		_w2875_
	);
	LUT4 #(
		.INIT('h080f)
	) name1873 (
		_w2859_,
		_w2861_,
		_w2866_,
		_w2867_,
		_w2876_
	);
	LUT2 #(
		.INIT('h1)
	) name1874 (
		_w2868_,
		_w2876_,
		_w2877_
	);
	LUT4 #(
		.INIT('h10f1)
	) name1875 (
		_w2871_,
		_w2874_,
		_w2875_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('he11e)
	) name1876 (
		_w2871_,
		_w2874_,
		_w2875_,
		_w2877_,
		_w2879_
	);
	LUT2 #(
		.INIT('h8)
	) name1877 (
		\A[82] ,
		\A[83] ,
		_w2880_
	);
	LUT3 #(
		.INIT('h96)
	) name1878 (
		\A[79] ,
		\A[80] ,
		\A[81] ,
		_w2881_
	);
	LUT3 #(
		.INIT('h96)
	) name1879 (
		\A[82] ,
		\A[83] ,
		\A[84] ,
		_w2882_
	);
	LUT3 #(
		.INIT('h80)
	) name1880 (
		_w2880_,
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT3 #(
		.INIT('h17)
	) name1881 (
		\A[79] ,
		\A[80] ,
		\A[81] ,
		_w2884_
	);
	LUT3 #(
		.INIT('h17)
	) name1882 (
		\A[82] ,
		\A[83] ,
		\A[84] ,
		_w2885_
	);
	LUT4 #(
		.INIT('h080f)
	) name1883 (
		_w2881_,
		_w2882_,
		_w2884_,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h1)
	) name1884 (
		_w2883_,
		_w2886_,
		_w2887_
	);
	LUT3 #(
		.INIT('h96)
	) name1885 (
		\A[85] ,
		\A[86] ,
		\A[87] ,
		_w2888_
	);
	LUT3 #(
		.INIT('h96)
	) name1886 (
		\A[88] ,
		\A[89] ,
		\A[90] ,
		_w2889_
	);
	LUT2 #(
		.INIT('h8)
	) name1887 (
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT4 #(
		.INIT('h0660)
	) name1888 (
		_w2881_,
		_w2882_,
		_w2888_,
		_w2889_,
		_w2891_
	);
	LUT3 #(
		.INIT('h17)
	) name1889 (
		\A[88] ,
		\A[89] ,
		\A[90] ,
		_w2892_
	);
	LUT3 #(
		.INIT('h17)
	) name1890 (
		\A[85] ,
		\A[86] ,
		\A[87] ,
		_w2893_
	);
	LUT2 #(
		.INIT('h6)
	) name1891 (
		_w2892_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1892 (
		\A[82] ,
		\A[83] ,
		\A[84] ,
		_w2881_,
		_w2895_
	);
	LUT2 #(
		.INIT('h9)
	) name1893 (
		_w2884_,
		_w2895_,
		_w2896_
	);
	LUT4 #(
		.INIT('h152a)
	) name1894 (
		_w2884_,
		_w2891_,
		_w2894_,
		_w2895_,
		_w2897_
	);
	LUT4 #(
		.INIT('h8008)
	) name1895 (
		_w2888_,
		_w2889_,
		_w2892_,
		_w2893_,
		_w2898_
	);
	LUT4 #(
		.INIT('h0770)
	) name1896 (
		_w2888_,
		_w2889_,
		_w2892_,
		_w2893_,
		_w2899_
	);
	LUT3 #(
		.INIT('h01)
	) name1897 (
		_w2891_,
		_w2899_,
		_w2898_,
		_w2900_
	);
	LUT4 #(
		.INIT('h088f)
	) name1898 (
		_w2888_,
		_w2889_,
		_w2892_,
		_w2893_,
		_w2901_
	);
	LUT4 #(
		.INIT('ha956)
	) name1899 (
		_w2887_,
		_w2897_,
		_w2900_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h8)
	) name1900 (
		_w2879_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w2879_,
		_w2902_,
		_w2904_
	);
	LUT4 #(
		.INIT('h6996)
	) name1902 (
		_w2856_,
		_w2857_,
		_w2859_,
		_w2861_,
		_w2905_
	);
	LUT4 #(
		.INIT('h6996)
	) name1903 (
		_w2881_,
		_w2882_,
		_w2888_,
		_w2889_,
		_w2906_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		_w2905_,
		_w2906_,
		_w2907_
	);
	LUT3 #(
		.INIT('h1e)
	) name1905 (
		_w2858_,
		_w2862_,
		_w2865_,
		_w2908_
	);
	LUT3 #(
		.INIT('h48)
	) name1906 (
		_w2870_,
		_w2907_,
		_w2908_,
		_w2909_
	);
	LUT3 #(
		.INIT('h21)
	) name1907 (
		_w2870_,
		_w2907_,
		_w2908_,
		_w2910_
	);
	LUT3 #(
		.INIT('h1e)
	) name1908 (
		_w2890_,
		_w2891_,
		_w2894_,
		_w2911_
	);
	LUT2 #(
		.INIT('h9)
	) name1909 (
		_w2896_,
		_w2911_,
		_w2912_
	);
	LUT3 #(
		.INIT('h54)
	) name1910 (
		_w2909_,
		_w2910_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('h1501)
	) name1911 (
		_w2878_,
		_w2879_,
		_w2902_,
		_w2913_,
		_w2914_
	);
	LUT4 #(
		.INIT('h80a8)
	) name1912 (
		_w2878_,
		_w2879_,
		_w2902_,
		_w2913_,
		_w2915_
	);
	LUT4 #(
		.INIT('h5701)
	) name1913 (
		_w2887_,
		_w2897_,
		_w2900_,
		_w2901_,
		_w2916_
	);
	LUT3 #(
		.INIT('h54)
	) name1914 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2917_
	);
	LUT3 #(
		.INIT('h96)
	) name1915 (
		\A[121] ,
		\A[122] ,
		\A[123] ,
		_w2918_
	);
	LUT3 #(
		.INIT('h96)
	) name1916 (
		\A[124] ,
		\A[125] ,
		\A[126] ,
		_w2919_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		_w2918_,
		_w2919_,
		_w2920_
	);
	LUT3 #(
		.INIT('h96)
	) name1918 (
		\A[115] ,
		\A[116] ,
		\A[117] ,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name1919 (
		\A[118] ,
		\A[119] ,
		_w2922_
	);
	LUT3 #(
		.INIT('h96)
	) name1920 (
		\A[118] ,
		\A[119] ,
		\A[120] ,
		_w2923_
	);
	LUT4 #(
		.INIT('h0660)
	) name1921 (
		_w2918_,
		_w2919_,
		_w2921_,
		_w2923_,
		_w2924_
	);
	LUT3 #(
		.INIT('h17)
	) name1922 (
		\A[124] ,
		\A[125] ,
		\A[126] ,
		_w2925_
	);
	LUT3 #(
		.INIT('h17)
	) name1923 (
		\A[121] ,
		\A[122] ,
		\A[123] ,
		_w2926_
	);
	LUT2 #(
		.INIT('h6)
	) name1924 (
		_w2925_,
		_w2926_,
		_w2927_
	);
	LUT3 #(
		.INIT('h17)
	) name1925 (
		\A[115] ,
		\A[116] ,
		\A[117] ,
		_w2928_
	);
	LUT3 #(
		.INIT('h17)
	) name1926 (
		\A[118] ,
		\A[119] ,
		\A[120] ,
		_w2929_
	);
	LUT3 #(
		.INIT('h80)
	) name1927 (
		_w2921_,
		_w2922_,
		_w2923_,
		_w2930_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1928 (
		\A[118] ,
		\A[119] ,
		\A[120] ,
		_w2921_,
		_w2931_
	);
	LUT2 #(
		.INIT('h9)
	) name1929 (
		_w2928_,
		_w2931_,
		_w2932_
	);
	LUT4 #(
		.INIT('h0770)
	) name1930 (
		_w2924_,
		_w2927_,
		_w2928_,
		_w2931_,
		_w2933_
	);
	LUT4 #(
		.INIT('h8008)
	) name1931 (
		_w2918_,
		_w2919_,
		_w2925_,
		_w2926_,
		_w2934_
	);
	LUT4 #(
		.INIT('h0770)
	) name1932 (
		_w2918_,
		_w2919_,
		_w2925_,
		_w2926_,
		_w2935_
	);
	LUT3 #(
		.INIT('h01)
	) name1933 (
		_w2924_,
		_w2935_,
		_w2934_,
		_w2936_
	);
	LUT4 #(
		.INIT('h088f)
	) name1934 (
		_w2918_,
		_w2919_,
		_w2925_,
		_w2926_,
		_w2937_
	);
	LUT4 #(
		.INIT('h080f)
	) name1935 (
		_w2921_,
		_w2923_,
		_w2928_,
		_w2929_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name1936 (
		_w2930_,
		_w2938_,
		_w2939_
	);
	LUT4 #(
		.INIT('h10f1)
	) name1937 (
		_w2933_,
		_w2936_,
		_w2937_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('he11e)
	) name1938 (
		_w2933_,
		_w2936_,
		_w2937_,
		_w2939_,
		_w2941_
	);
	LUT2 #(
		.INIT('h8)
	) name1939 (
		\A[106] ,
		\A[107] ,
		_w2942_
	);
	LUT3 #(
		.INIT('h96)
	) name1940 (
		\A[103] ,
		\A[104] ,
		\A[105] ,
		_w2943_
	);
	LUT3 #(
		.INIT('h96)
	) name1941 (
		\A[106] ,
		\A[107] ,
		\A[108] ,
		_w2944_
	);
	LUT3 #(
		.INIT('h80)
	) name1942 (
		_w2942_,
		_w2943_,
		_w2944_,
		_w2945_
	);
	LUT3 #(
		.INIT('h17)
	) name1943 (
		\A[103] ,
		\A[104] ,
		\A[105] ,
		_w2946_
	);
	LUT3 #(
		.INIT('h17)
	) name1944 (
		\A[106] ,
		\A[107] ,
		\A[108] ,
		_w2947_
	);
	LUT4 #(
		.INIT('h080f)
	) name1945 (
		_w2943_,
		_w2944_,
		_w2946_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w2945_,
		_w2948_,
		_w2949_
	);
	LUT3 #(
		.INIT('h96)
	) name1947 (
		\A[109] ,
		\A[110] ,
		\A[111] ,
		_w2950_
	);
	LUT3 #(
		.INIT('h96)
	) name1948 (
		\A[112] ,
		\A[113] ,
		\A[114] ,
		_w2951_
	);
	LUT2 #(
		.INIT('h8)
	) name1949 (
		_w2950_,
		_w2951_,
		_w2952_
	);
	LUT4 #(
		.INIT('h0660)
	) name1950 (
		_w2943_,
		_w2944_,
		_w2950_,
		_w2951_,
		_w2953_
	);
	LUT3 #(
		.INIT('h17)
	) name1951 (
		\A[112] ,
		\A[113] ,
		\A[114] ,
		_w2954_
	);
	LUT3 #(
		.INIT('h17)
	) name1952 (
		\A[109] ,
		\A[110] ,
		\A[111] ,
		_w2955_
	);
	LUT2 #(
		.INIT('h6)
	) name1953 (
		_w2954_,
		_w2955_,
		_w2956_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name1954 (
		\A[106] ,
		\A[107] ,
		\A[108] ,
		_w2943_,
		_w2957_
	);
	LUT2 #(
		.INIT('h9)
	) name1955 (
		_w2946_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h152a)
	) name1956 (
		_w2946_,
		_w2953_,
		_w2956_,
		_w2957_,
		_w2959_
	);
	LUT4 #(
		.INIT('h8008)
	) name1957 (
		_w2950_,
		_w2951_,
		_w2954_,
		_w2955_,
		_w2960_
	);
	LUT4 #(
		.INIT('h0770)
	) name1958 (
		_w2950_,
		_w2951_,
		_w2954_,
		_w2955_,
		_w2961_
	);
	LUT3 #(
		.INIT('h01)
	) name1959 (
		_w2953_,
		_w2961_,
		_w2960_,
		_w2962_
	);
	LUT4 #(
		.INIT('h088f)
	) name1960 (
		_w2950_,
		_w2951_,
		_w2954_,
		_w2955_,
		_w2963_
	);
	LUT4 #(
		.INIT('ha956)
	) name1961 (
		_w2949_,
		_w2959_,
		_w2962_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h8)
	) name1962 (
		_w2941_,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h1)
	) name1963 (
		_w2941_,
		_w2964_,
		_w2966_
	);
	LUT4 #(
		.INIT('h6996)
	) name1964 (
		_w2918_,
		_w2919_,
		_w2921_,
		_w2923_,
		_w2967_
	);
	LUT4 #(
		.INIT('h6996)
	) name1965 (
		_w2943_,
		_w2944_,
		_w2950_,
		_w2951_,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name1966 (
		_w2967_,
		_w2968_,
		_w2969_
	);
	LUT3 #(
		.INIT('h1e)
	) name1967 (
		_w2920_,
		_w2924_,
		_w2927_,
		_w2970_
	);
	LUT3 #(
		.INIT('h48)
	) name1968 (
		_w2932_,
		_w2969_,
		_w2970_,
		_w2971_
	);
	LUT3 #(
		.INIT('h21)
	) name1969 (
		_w2932_,
		_w2969_,
		_w2970_,
		_w2972_
	);
	LUT3 #(
		.INIT('h1e)
	) name1970 (
		_w2952_,
		_w2953_,
		_w2956_,
		_w2973_
	);
	LUT2 #(
		.INIT('h9)
	) name1971 (
		_w2958_,
		_w2973_,
		_w2974_
	);
	LUT3 #(
		.INIT('h54)
	) name1972 (
		_w2971_,
		_w2972_,
		_w2974_,
		_w2975_
	);
	LUT4 #(
		.INIT('h1501)
	) name1973 (
		_w2940_,
		_w2941_,
		_w2964_,
		_w2975_,
		_w2976_
	);
	LUT4 #(
		.INIT('h80a8)
	) name1974 (
		_w2940_,
		_w2941_,
		_w2964_,
		_w2975_,
		_w2977_
	);
	LUT4 #(
		.INIT('h5701)
	) name1975 (
		_w2949_,
		_w2959_,
		_w2962_,
		_w2963_,
		_w2978_
	);
	LUT3 #(
		.INIT('h54)
	) name1976 (
		_w2976_,
		_w2977_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w2917_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		_w2917_,
		_w2979_,
		_w2981_
	);
	LUT4 #(
		.INIT('h6665)
	) name1979 (
		_w2940_,
		_w2965_,
		_w2966_,
		_w2975_,
		_w2982_
	);
	LUT4 #(
		.INIT('h6665)
	) name1980 (
		_w2878_,
		_w2903_,
		_w2904_,
		_w2913_,
		_w2983_
	);
	LUT4 #(
		.INIT('h8241)
	) name1981 (
		_w2916_,
		_w2978_,
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT4 #(
		.INIT('h1428)
	) name1982 (
		_w2916_,
		_w2978_,
		_w2982_,
		_w2983_,
		_w2985_
	);
	LUT2 #(
		.INIT('h6)
	) name1983 (
		_w2879_,
		_w2902_,
		_w2986_
	);
	LUT2 #(
		.INIT('h6)
	) name1984 (
		_w2941_,
		_w2964_,
		_w2987_
	);
	LUT4 #(
		.INIT('h1248)
	) name1985 (
		_w2913_,
		_w2975_,
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('h8421)
	) name1986 (
		_w2913_,
		_w2975_,
		_w2986_,
		_w2987_,
		_w2989_
	);
	LUT4 #(
		.INIT('h0660)
	) name1987 (
		_w2905_,
		_w2906_,
		_w2967_,
		_w2968_,
		_w2990_
	);
	LUT3 #(
		.INIT('h96)
	) name1988 (
		_w2932_,
		_w2969_,
		_w2970_,
		_w2991_
	);
	LUT3 #(
		.INIT('h84)
	) name1989 (
		_w2974_,
		_w2990_,
		_w2991_,
		_w2992_
	);
	LUT3 #(
		.INIT('h12)
	) name1990 (
		_w2974_,
		_w2990_,
		_w2991_,
		_w2993_
	);
	LUT3 #(
		.INIT('h96)
	) name1991 (
		_w2870_,
		_w2907_,
		_w2908_,
		_w2994_
	);
	LUT2 #(
		.INIT('h9)
	) name1992 (
		_w2912_,
		_w2994_,
		_w2995_
	);
	LUT3 #(
		.INIT('h45)
	) name1993 (
		_w2992_,
		_w2993_,
		_w2995_,
		_w2996_
	);
	LUT3 #(
		.INIT('h45)
	) name1994 (
		_w2988_,
		_w2989_,
		_w2996_,
		_w2997_
	);
	LUT3 #(
		.INIT('h54)
	) name1995 (
		_w2984_,
		_w2985_,
		_w2997_,
		_w2998_
	);
	LUT3 #(
		.INIT('h54)
	) name1996 (
		_w2980_,
		_w2981_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h1)
	) name1997 (
		_w2855_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h8)
	) name1998 (
		_w2855_,
		_w2999_,
		_w3001_
	);
	LUT2 #(
		.INIT('h6)
	) name1999 (
		_w2917_,
		_w2979_,
		_w3002_
	);
	LUT2 #(
		.INIT('h6)
	) name2000 (
		_w2773_,
		_w2835_,
		_w3003_
	);
	LUT4 #(
		.INIT('h1428)
	) name2001 (
		_w2854_,
		_w2998_,
		_w3002_,
		_w3003_,
		_w3004_
	);
	LUT4 #(
		.INIT('h8241)
	) name2002 (
		_w2854_,
		_w2998_,
		_w3002_,
		_w3003_,
		_w3005_
	);
	LUT4 #(
		.INIT('h6996)
	) name2003 (
		_w2772_,
		_w2834_,
		_w2838_,
		_w2839_,
		_w3006_
	);
	LUT4 #(
		.INIT('h6996)
	) name2004 (
		_w2916_,
		_w2978_,
		_w2982_,
		_w2983_,
		_w3007_
	);
	LUT4 #(
		.INIT('h1248)
	) name2005 (
		_w2853_,
		_w2997_,
		_w3006_,
		_w3007_,
		_w3008_
	);
	LUT4 #(
		.INIT('h8421)
	) name2006 (
		_w2853_,
		_w2997_,
		_w3006_,
		_w3007_,
		_w3009_
	);
	LUT4 #(
		.INIT('h6996)
	) name2007 (
		_w2913_,
		_w2975_,
		_w2986_,
		_w2987_,
		_w3010_
	);
	LUT4 #(
		.INIT('h6996)
	) name2008 (
		_w2769_,
		_w2831_,
		_w2842_,
		_w2843_,
		_w3011_
	);
	LUT4 #(
		.INIT('h1428)
	) name2009 (
		_w2852_,
		_w2996_,
		_w3010_,
		_w3011_,
		_w3012_
	);
	LUT4 #(
		.INIT('h8241)
	) name2010 (
		_w2852_,
		_w2996_,
		_w3010_,
		_w3011_,
		_w3013_
	);
	LUT4 #(
		.INIT('h6996)
	) name2011 (
		_w2761_,
		_w2762_,
		_w2823_,
		_w2824_,
		_w3014_
	);
	LUT4 #(
		.INIT('h6996)
	) name2012 (
		_w2905_,
		_w2906_,
		_w2967_,
		_w2968_,
		_w3015_
	);
	LUT2 #(
		.INIT('h8)
	) name2013 (
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT3 #(
		.INIT('h69)
	) name2014 (
		_w2830_,
		_w2846_,
		_w2847_,
		_w3017_
	);
	LUT3 #(
		.INIT('h48)
	) name2015 (
		_w2851_,
		_w3016_,
		_w3017_,
		_w3018_
	);
	LUT3 #(
		.INIT('h21)
	) name2016 (
		_w2851_,
		_w3016_,
		_w3017_,
		_w3019_
	);
	LUT3 #(
		.INIT('h69)
	) name2017 (
		_w2974_,
		_w2990_,
		_w2991_,
		_w3020_
	);
	LUT2 #(
		.INIT('h9)
	) name2018 (
		_w2995_,
		_w3020_,
		_w3021_
	);
	LUT3 #(
		.INIT('h54)
	) name2019 (
		_w3018_,
		_w3019_,
		_w3021_,
		_w3022_
	);
	LUT3 #(
		.INIT('h45)
	) name2020 (
		_w3012_,
		_w3013_,
		_w3022_,
		_w3023_
	);
	LUT3 #(
		.INIT('h45)
	) name2021 (
		_w3008_,
		_w3009_,
		_w3023_,
		_w3024_
	);
	LUT3 #(
		.INIT('h54)
	) name2022 (
		_w3004_,
		_w3005_,
		_w3024_,
		_w3025_
	);
	LUT3 #(
		.INIT('h45)
	) name2023 (
		_w3000_,
		_w3001_,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h4)
	) name2024 (
		_w2711_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h2)
	) name2025 (
		_w2711_,
		_w3026_,
		_w3028_
	);
	LUT2 #(
		.INIT('h6)
	) name2026 (
		_w2855_,
		_w2999_,
		_w3029_
	);
	LUT2 #(
		.INIT('h6)
	) name2027 (
		_w2539_,
		_w2686_,
		_w3030_
	);
	LUT4 #(
		.INIT('h4182)
	) name2028 (
		_w2710_,
		_w3025_,
		_w3029_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('h2814)
	) name2029 (
		_w2710_,
		_w3025_,
		_w3029_,
		_w3030_,
		_w3032_
	);
	LUT4 #(
		.INIT('h6996)
	) name2030 (
		_w2854_,
		_w2998_,
		_w3002_,
		_w3003_,
		_w3033_
	);
	LUT4 #(
		.INIT('h9669)
	) name2031 (
		_w2538_,
		_w2685_,
		_w2689_,
		_w2690_,
		_w3034_
	);
	LUT4 #(
		.INIT('h2814)
	) name2032 (
		_w2709_,
		_w3024_,
		_w3033_,
		_w3034_,
		_w3035_
	);
	LUT4 #(
		.INIT('h4182)
	) name2033 (
		_w2709_,
		_w3024_,
		_w3033_,
		_w3034_,
		_w3036_
	);
	LUT4 #(
		.INIT('h6996)
	) name2034 (
		_w2537_,
		_w2684_,
		_w2693_,
		_w2694_,
		_w3037_
	);
	LUT4 #(
		.INIT('h6996)
	) name2035 (
		_w2853_,
		_w2997_,
		_w3006_,
		_w3007_,
		_w3038_
	);
	LUT4 #(
		.INIT('h8421)
	) name2036 (
		_w2708_,
		_w3023_,
		_w3037_,
		_w3038_,
		_w3039_
	);
	LUT4 #(
		.INIT('h1248)
	) name2037 (
		_w2708_,
		_w3023_,
		_w3037_,
		_w3038_,
		_w3040_
	);
	LUT4 #(
		.INIT('h6996)
	) name2038 (
		_w2852_,
		_w2996_,
		_w3010_,
		_w3011_,
		_w3041_
	);
	LUT2 #(
		.INIT('h9)
	) name2039 (
		_w3022_,
		_w3041_,
		_w3042_
	);
	LUT3 #(
		.INIT('h69)
	) name2040 (
		_w2697_,
		_w2698_,
		_w2707_,
		_w3043_
	);
	LUT4 #(
		.INIT('h0660)
	) name2041 (
		_w2699_,
		_w2700_,
		_w3014_,
		_w3015_,
		_w3044_
	);
	LUT3 #(
		.INIT('h96)
	) name2042 (
		_w2682_,
		_w2701_,
		_w2702_,
		_w3045_
	);
	LUT3 #(
		.INIT('h84)
	) name2043 (
		_w2706_,
		_w3044_,
		_w3045_,
		_w3046_
	);
	LUT3 #(
		.INIT('h12)
	) name2044 (
		_w2706_,
		_w3044_,
		_w3045_,
		_w3047_
	);
	LUT3 #(
		.INIT('h96)
	) name2045 (
		_w2851_,
		_w3016_,
		_w3017_,
		_w3048_
	);
	LUT2 #(
		.INIT('h9)
	) name2046 (
		_w3021_,
		_w3048_,
		_w3049_
	);
	LUT3 #(
		.INIT('h45)
	) name2047 (
		_w3046_,
		_w3047_,
		_w3049_,
		_w3050_
	);
	LUT3 #(
		.INIT('h8e)
	) name2048 (
		_w3042_,
		_w3043_,
		_w3050_,
		_w3051_
	);
	LUT3 #(
		.INIT('h54)
	) name2049 (
		_w3039_,
		_w3040_,
		_w3051_,
		_w3052_
	);
	LUT3 #(
		.INIT('h54)
	) name2050 (
		_w3035_,
		_w3036_,
		_w3052_,
		_w3053_
	);
	LUT3 #(
		.INIT('h45)
	) name2051 (
		_w3031_,
		_w3032_,
		_w3053_,
		_w3054_
	);
	LUT3 #(
		.INIT('h54)
	) name2052 (
		_w3027_,
		_w3028_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w2389_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w2389_,
		_w3055_,
		_w3057_
	);
	LUT2 #(
		.INIT('h6)
	) name2055 (
		_w2088_,
		_w2362_,
		_w3058_
	);
	LUT2 #(
		.INIT('h9)
	) name2056 (
		_w2711_,
		_w3026_,
		_w3059_
	);
	LUT4 #(
		.INIT('h2184)
	) name2057 (
		_w2388_,
		_w3054_,
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('h4812)
	) name2058 (
		_w2388_,
		_w3054_,
		_w3058_,
		_w3059_,
		_w3061_
	);
	LUT4 #(
		.INIT('h9669)
	) name2059 (
		_w2710_,
		_w3025_,
		_w3029_,
		_w3030_,
		_w3062_
	);
	LUT3 #(
		.INIT('h96)
	) name2060 (
		_w2087_,
		_w2365_,
		_w2367_,
		_w3063_
	);
	LUT4 #(
		.INIT('h1428)
	) name2061 (
		_w2387_,
		_w3053_,
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT4 #(
		.INIT('h8241)
	) name2062 (
		_w2387_,
		_w3053_,
		_w3062_,
		_w3063_,
		_w3065_
	);
	LUT4 #(
		.INIT('h9669)
	) name2063 (
		_w2709_,
		_w3024_,
		_w3033_,
		_w3034_,
		_w3066_
	);
	LUT4 #(
		.INIT('h9669)
	) name2064 (
		_w2086_,
		_w2360_,
		_w2370_,
		_w2371_,
		_w3067_
	);
	LUT4 #(
		.INIT('h1428)
	) name2065 (
		_w2386_,
		_w3052_,
		_w3066_,
		_w3067_,
		_w3068_
	);
	LUT4 #(
		.INIT('h8241)
	) name2066 (
		_w2386_,
		_w3052_,
		_w3066_,
		_w3067_,
		_w3069_
	);
	LUT4 #(
		.INIT('h6996)
	) name2067 (
		_w2085_,
		_w2359_,
		_w2374_,
		_w2375_,
		_w3070_
	);
	LUT4 #(
		.INIT('h6996)
	) name2068 (
		_w2708_,
		_w3023_,
		_w3037_,
		_w3038_,
		_w3071_
	);
	LUT4 #(
		.INIT('h1248)
	) name2069 (
		_w2385_,
		_w3051_,
		_w3070_,
		_w3071_,
		_w3072_
	);
	LUT4 #(
		.INIT('h8421)
	) name2070 (
		_w2385_,
		_w3051_,
		_w3070_,
		_w3071_,
		_w3073_
	);
	LUT3 #(
		.INIT('h69)
	) name2071 (
		_w3042_,
		_w3043_,
		_w3050_,
		_w3074_
	);
	LUT3 #(
		.INIT('h69)
	) name2072 (
		_w2379_,
		_w2380_,
		_w2384_,
		_w3075_
	);
	LUT4 #(
		.INIT('h6996)
	) name2073 (
		_w2076_,
		_w2077_,
		_w2352_,
		_w2353_,
		_w3076_
	);
	LUT4 #(
		.INIT('h6996)
	) name2074 (
		_w2699_,
		_w2700_,
		_w3014_,
		_w3015_,
		_w3077_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		_w3076_,
		_w3077_,
		_w3078_
	);
	LUT4 #(
		.INIT('h6996)
	) name2076 (
		_w2083_,
		_w2381_,
		_w2382_,
		_w2383_,
		_w3079_
	);
	LUT3 #(
		.INIT('h69)
	) name2077 (
		_w2706_,
		_w3044_,
		_w3045_,
		_w3080_
	);
	LUT4 #(
		.INIT('hb271)
	) name2078 (
		_w3049_,
		_w3078_,
		_w3079_,
		_w3080_,
		_w3081_
	);
	LUT3 #(
		.INIT('h8e)
	) name2079 (
		_w3074_,
		_w3075_,
		_w3081_,
		_w3082_
	);
	LUT3 #(
		.INIT('h45)
	) name2080 (
		_w3072_,
		_w3073_,
		_w3082_,
		_w3083_
	);
	LUT3 #(
		.INIT('h54)
	) name2081 (
		_w3068_,
		_w3069_,
		_w3083_,
		_w3084_
	);
	LUT3 #(
		.INIT('h54)
	) name2082 (
		_w3064_,
		_w3065_,
		_w3084_,
		_w3085_
	);
	LUT3 #(
		.INIT('h45)
	) name2083 (
		_w3060_,
		_w3061_,
		_w3085_,
		_w3086_
	);
	LUT4 #(
		.INIT('h4054)
	) name2084 (
		_w1769_,
		_w2389_,
		_w3055_,
		_w3086_,
		_w3087_
	);
	LUT4 #(
		.INIT('h2a02)
	) name2085 (
		_w1769_,
		_w2389_,
		_w3055_,
		_w3086_,
		_w3088_
	);
	LUT4 #(
		.INIT('h6566)
	) name2086 (
		_w1769_,
		_w3056_,
		_w3057_,
		_w3086_,
		_w3089_
	);
	LUT3 #(
		.INIT('h60)
	) name2087 (
		_w1406_,
		_w1408_,
		_w1743_,
		_w3090_
	);
	LUT4 #(
		.INIT('h0065)
	) name2088 (
		_w1409_,
		_w1744_,
		_w1768_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h6)
	) name2089 (
		_w2389_,
		_w3055_,
		_w3092_
	);
	LUT2 #(
		.INIT('h9)
	) name2090 (
		_w3086_,
		_w3092_,
		_w3093_
	);
	LUT3 #(
		.INIT('h84)
	) name2091 (
		_w3086_,
		_w3091_,
		_w3092_,
		_w3094_
	);
	LUT3 #(
		.INIT('h12)
	) name2092 (
		_w3086_,
		_w3091_,
		_w3092_,
		_w3095_
	);
	LUT3 #(
		.INIT('h96)
	) name2093 (
		_w1406_,
		_w1408_,
		_w1743_,
		_w3096_
	);
	LUT2 #(
		.INIT('h9)
	) name2094 (
		_w1768_,
		_w3096_,
		_w3097_
	);
	LUT4 #(
		.INIT('h9669)
	) name2095 (
		_w2388_,
		_w3054_,
		_w3058_,
		_w3059_,
		_w3098_
	);
	LUT3 #(
		.INIT('h48)
	) name2096 (
		_w3085_,
		_w3097_,
		_w3098_,
		_w3099_
	);
	LUT3 #(
		.INIT('h21)
	) name2097 (
		_w3085_,
		_w3097_,
		_w3098_,
		_w3100_
	);
	LUT3 #(
		.INIT('h69)
	) name2098 (
		_w1745_,
		_w1747_,
		_w1767_,
		_w3101_
	);
	LUT4 #(
		.INIT('h6996)
	) name2099 (
		_w2387_,
		_w3053_,
		_w3062_,
		_w3063_,
		_w3102_
	);
	LUT3 #(
		.INIT('h48)
	) name2100 (
		_w3084_,
		_w3101_,
		_w3102_,
		_w3103_
	);
	LUT3 #(
		.INIT('h21)
	) name2101 (
		_w3084_,
		_w3101_,
		_w3102_,
		_w3104_
	);
	LUT3 #(
		.INIT('h96)
	) name2102 (
		_w1749_,
		_w1750_,
		_w1766_,
		_w3105_
	);
	LUT4 #(
		.INIT('h6996)
	) name2103 (
		_w2386_,
		_w3052_,
		_w3066_,
		_w3067_,
		_w3106_
	);
	LUT3 #(
		.INIT('h48)
	) name2104 (
		_w3083_,
		_w3105_,
		_w3106_,
		_w3107_
	);
	LUT3 #(
		.INIT('h21)
	) name2105 (
		_w3083_,
		_w3105_,
		_w3106_,
		_w3108_
	);
	LUT4 #(
		.INIT('h6996)
	) name2106 (
		_w2385_,
		_w3051_,
		_w3070_,
		_w3071_,
		_w3109_
	);
	LUT3 #(
		.INIT('h96)
	) name2107 (
		_w1751_,
		_w1753_,
		_w1765_,
		_w3110_
	);
	LUT3 #(
		.INIT('h06)
	) name2108 (
		_w3082_,
		_w3109_,
		_w3110_,
		_w3111_
	);
	LUT3 #(
		.INIT('h90)
	) name2109 (
		_w3082_,
		_w3109_,
		_w3110_,
		_w3112_
	);
	LUT3 #(
		.INIT('h69)
	) name2110 (
		_w1755_,
		_w1756_,
		_w1764_,
		_w3113_
	);
	LUT4 #(
		.INIT('h0096)
	) name2111 (
		_w3074_,
		_w3075_,
		_w3081_,
		_w3113_,
		_w3114_
	);
	LUT4 #(
		.INIT('h6900)
	) name2112 (
		_w3074_,
		_w3075_,
		_w3081_,
		_w3113_,
		_w3115_
	);
	LUT4 #(
		.INIT('h0660)
	) name2113 (
		_w1757_,
		_w1758_,
		_w3076_,
		_w3077_,
		_w3116_
	);
	LUT4 #(
		.INIT('h6996)
	) name2114 (
		_w3049_,
		_w3078_,
		_w3079_,
		_w3080_,
		_w3117_
	);
	LUT4 #(
		.INIT('h9669)
	) name2115 (
		_w1398_,
		_w1399_,
		_w1401_,
		_w1759_,
		_w3118_
	);
	LUT2 #(
		.INIT('h9)
	) name2116 (
		_w1763_,
		_w3118_,
		_w3119_
	);
	LUT3 #(
		.INIT('h4d)
	) name2117 (
		_w3116_,
		_w3117_,
		_w3119_,
		_w3120_
	);
	LUT3 #(
		.INIT('h45)
	) name2118 (
		_w3114_,
		_w3115_,
		_w3120_,
		_w3121_
	);
	LUT3 #(
		.INIT('h45)
	) name2119 (
		_w3111_,
		_w3112_,
		_w3121_,
		_w3122_
	);
	LUT3 #(
		.INIT('h45)
	) name2120 (
		_w3107_,
		_w3108_,
		_w3122_,
		_w3123_
	);
	LUT3 #(
		.INIT('h54)
	) name2121 (
		_w3103_,
		_w3104_,
		_w3123_,
		_w3124_
	);
	LUT3 #(
		.INIT('h54)
	) name2122 (
		_w3099_,
		_w3100_,
		_w3124_,
		_w3125_
	);
	LUT4 #(
		.INIT('h6665)
	) name2123 (
		_w3089_,
		_w3094_,
		_w3095_,
		_w3125_,
		_w3126_
	);
	LUT3 #(
		.INIT('h96)
	) name2124 (
		\A[835] ,
		\A[836] ,
		\A[837] ,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name2125 (
		\A[838] ,
		\A[839] ,
		_w3128_
	);
	LUT3 #(
		.INIT('h96)
	) name2126 (
		\A[838] ,
		\A[839] ,
		\A[840] ,
		_w3129_
	);
	LUT3 #(
		.INIT('h96)
	) name2127 (
		\A[841] ,
		\A[842] ,
		\A[843] ,
		_w3130_
	);
	LUT3 #(
		.INIT('h96)
	) name2128 (
		\A[844] ,
		\A[845] ,
		\A[846] ,
		_w3131_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		_w3130_,
		_w3131_,
		_w3132_
	);
	LUT4 #(
		.INIT('h0660)
	) name2130 (
		_w3127_,
		_w3129_,
		_w3130_,
		_w3131_,
		_w3133_
	);
	LUT3 #(
		.INIT('h17)
	) name2131 (
		\A[844] ,
		\A[845] ,
		\A[846] ,
		_w3134_
	);
	LUT3 #(
		.INIT('h17)
	) name2132 (
		\A[841] ,
		\A[842] ,
		\A[843] ,
		_w3135_
	);
	LUT2 #(
		.INIT('h6)
	) name2133 (
		_w3134_,
		_w3135_,
		_w3136_
	);
	LUT3 #(
		.INIT('h17)
	) name2134 (
		\A[835] ,
		\A[836] ,
		\A[837] ,
		_w3137_
	);
	LUT3 #(
		.INIT('h80)
	) name2135 (
		_w3127_,
		_w3128_,
		_w3129_,
		_w3138_
	);
	LUT3 #(
		.INIT('h17)
	) name2136 (
		\A[838] ,
		\A[839] ,
		\A[840] ,
		_w3139_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2137 (
		\A[838] ,
		\A[839] ,
		\A[840] ,
		_w3127_,
		_w3140_
	);
	LUT2 #(
		.INIT('h9)
	) name2138 (
		_w3137_,
		_w3140_,
		_w3141_
	);
	LUT4 #(
		.INIT('h0770)
	) name2139 (
		_w3133_,
		_w3136_,
		_w3137_,
		_w3140_,
		_w3142_
	);
	LUT4 #(
		.INIT('h8008)
	) name2140 (
		_w3130_,
		_w3131_,
		_w3134_,
		_w3135_,
		_w3143_
	);
	LUT4 #(
		.INIT('h0770)
	) name2141 (
		_w3130_,
		_w3131_,
		_w3134_,
		_w3135_,
		_w3144_
	);
	LUT3 #(
		.INIT('h01)
	) name2142 (
		_w3133_,
		_w3144_,
		_w3143_,
		_w3145_
	);
	LUT4 #(
		.INIT('hf770)
	) name2143 (
		_w3130_,
		_w3131_,
		_w3134_,
		_w3135_,
		_w3146_
	);
	LUT4 #(
		.INIT('h080f)
	) name2144 (
		_w3127_,
		_w3129_,
		_w3137_,
		_w3139_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		_w3138_,
		_w3147_,
		_w3148_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2146 (
		_w3142_,
		_w3145_,
		_w3146_,
		_w3148_,
		_w3149_
	);
	LUT3 #(
		.INIT('h96)
	) name2147 (
		\A[823] ,
		\A[824] ,
		\A[825] ,
		_w3150_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		\A[826] ,
		\A[827] ,
		_w3151_
	);
	LUT3 #(
		.INIT('h96)
	) name2149 (
		\A[826] ,
		\A[827] ,
		\A[828] ,
		_w3152_
	);
	LUT3 #(
		.INIT('h96)
	) name2150 (
		\A[829] ,
		\A[830] ,
		\A[831] ,
		_w3153_
	);
	LUT3 #(
		.INIT('h96)
	) name2151 (
		\A[832] ,
		\A[833] ,
		\A[834] ,
		_w3154_
	);
	LUT2 #(
		.INIT('h8)
	) name2152 (
		_w3153_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('h0660)
	) name2153 (
		_w3150_,
		_w3152_,
		_w3153_,
		_w3154_,
		_w3156_
	);
	LUT3 #(
		.INIT('h17)
	) name2154 (
		\A[832] ,
		\A[833] ,
		\A[834] ,
		_w3157_
	);
	LUT3 #(
		.INIT('h17)
	) name2155 (
		\A[829] ,
		\A[830] ,
		\A[831] ,
		_w3158_
	);
	LUT2 #(
		.INIT('h6)
	) name2156 (
		_w3157_,
		_w3158_,
		_w3159_
	);
	LUT3 #(
		.INIT('h17)
	) name2157 (
		\A[823] ,
		\A[824] ,
		\A[825] ,
		_w3160_
	);
	LUT3 #(
		.INIT('h80)
	) name2158 (
		_w3150_,
		_w3151_,
		_w3152_,
		_w3161_
	);
	LUT3 #(
		.INIT('h17)
	) name2159 (
		\A[826] ,
		\A[827] ,
		\A[828] ,
		_w3162_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2160 (
		\A[826] ,
		\A[827] ,
		\A[828] ,
		_w3150_,
		_w3163_
	);
	LUT2 #(
		.INIT('h9)
	) name2161 (
		_w3160_,
		_w3163_,
		_w3164_
	);
	LUT4 #(
		.INIT('h0770)
	) name2162 (
		_w3156_,
		_w3159_,
		_w3160_,
		_w3163_,
		_w3165_
	);
	LUT4 #(
		.INIT('h8008)
	) name2163 (
		_w3153_,
		_w3154_,
		_w3157_,
		_w3158_,
		_w3166_
	);
	LUT4 #(
		.INIT('h0770)
	) name2164 (
		_w3153_,
		_w3154_,
		_w3157_,
		_w3158_,
		_w3167_
	);
	LUT3 #(
		.INIT('h01)
	) name2165 (
		_w3156_,
		_w3167_,
		_w3166_,
		_w3168_
	);
	LUT4 #(
		.INIT('hf770)
	) name2166 (
		_w3153_,
		_w3154_,
		_w3157_,
		_w3158_,
		_w3169_
	);
	LUT4 #(
		.INIT('h080f)
	) name2167 (
		_w3150_,
		_w3152_,
		_w3160_,
		_w3162_,
		_w3170_
	);
	LUT2 #(
		.INIT('h1)
	) name2168 (
		_w3161_,
		_w3170_,
		_w3171_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2169 (
		_w3165_,
		_w3168_,
		_w3169_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w3149_,
		_w3172_,
		_w3173_
	);
	LUT2 #(
		.INIT('h8)
	) name2171 (
		_w3149_,
		_w3172_,
		_w3174_
	);
	LUT2 #(
		.INIT('h6)
	) name2172 (
		_w3149_,
		_w3172_,
		_w3175_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2173 (
		_w3165_,
		_w3168_,
		_w3169_,
		_w3171_,
		_w3176_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2174 (
		_w3142_,
		_w3145_,
		_w3146_,
		_w3148_,
		_w3177_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h8)
	) name2176 (
		_w3176_,
		_w3177_,
		_w3179_
	);
	LUT4 #(
		.INIT('h6996)
	) name2177 (
		_w3127_,
		_w3129_,
		_w3130_,
		_w3131_,
		_w3180_
	);
	LUT4 #(
		.INIT('h6996)
	) name2178 (
		_w3150_,
		_w3152_,
		_w3153_,
		_w3154_,
		_w3181_
	);
	LUT2 #(
		.INIT('h8)
	) name2179 (
		_w3180_,
		_w3181_,
		_w3182_
	);
	LUT3 #(
		.INIT('h1e)
	) name2180 (
		_w3132_,
		_w3133_,
		_w3136_,
		_w3183_
	);
	LUT3 #(
		.INIT('h48)
	) name2181 (
		_w3141_,
		_w3182_,
		_w3183_,
		_w3184_
	);
	LUT3 #(
		.INIT('h21)
	) name2182 (
		_w3141_,
		_w3182_,
		_w3183_,
		_w3185_
	);
	LUT3 #(
		.INIT('h1e)
	) name2183 (
		_w3155_,
		_w3156_,
		_w3159_,
		_w3186_
	);
	LUT2 #(
		.INIT('h9)
	) name2184 (
		_w3164_,
		_w3186_,
		_w3187_
	);
	LUT3 #(
		.INIT('h54)
	) name2185 (
		_w3184_,
		_w3185_,
		_w3187_,
		_w3188_
	);
	LUT4 #(
		.INIT('h6566)
	) name2186 (
		_w3175_,
		_w3178_,
		_w3179_,
		_w3188_,
		_w3189_
	);
	LUT3 #(
		.INIT('h96)
	) name2187 (
		\A[811] ,
		\A[812] ,
		\A[813] ,
		_w3190_
	);
	LUT2 #(
		.INIT('h8)
	) name2188 (
		\A[814] ,
		\A[815] ,
		_w3191_
	);
	LUT3 #(
		.INIT('h96)
	) name2189 (
		\A[814] ,
		\A[815] ,
		\A[816] ,
		_w3192_
	);
	LUT3 #(
		.INIT('h96)
	) name2190 (
		\A[817] ,
		\A[818] ,
		\A[819] ,
		_w3193_
	);
	LUT3 #(
		.INIT('h96)
	) name2191 (
		\A[820] ,
		\A[821] ,
		\A[822] ,
		_w3194_
	);
	LUT2 #(
		.INIT('h8)
	) name2192 (
		_w3193_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h0660)
	) name2193 (
		_w3190_,
		_w3192_,
		_w3193_,
		_w3194_,
		_w3196_
	);
	LUT3 #(
		.INIT('h17)
	) name2194 (
		\A[820] ,
		\A[821] ,
		\A[822] ,
		_w3197_
	);
	LUT3 #(
		.INIT('h17)
	) name2195 (
		\A[817] ,
		\A[818] ,
		\A[819] ,
		_w3198_
	);
	LUT2 #(
		.INIT('h6)
	) name2196 (
		_w3197_,
		_w3198_,
		_w3199_
	);
	LUT3 #(
		.INIT('h17)
	) name2197 (
		\A[811] ,
		\A[812] ,
		\A[813] ,
		_w3200_
	);
	LUT3 #(
		.INIT('h80)
	) name2198 (
		_w3190_,
		_w3191_,
		_w3192_,
		_w3201_
	);
	LUT3 #(
		.INIT('h17)
	) name2199 (
		\A[814] ,
		\A[815] ,
		\A[816] ,
		_w3202_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2200 (
		\A[814] ,
		\A[815] ,
		\A[816] ,
		_w3190_,
		_w3203_
	);
	LUT2 #(
		.INIT('h9)
	) name2201 (
		_w3200_,
		_w3203_,
		_w3204_
	);
	LUT4 #(
		.INIT('h0770)
	) name2202 (
		_w3196_,
		_w3199_,
		_w3200_,
		_w3203_,
		_w3205_
	);
	LUT4 #(
		.INIT('h8008)
	) name2203 (
		_w3193_,
		_w3194_,
		_w3197_,
		_w3198_,
		_w3206_
	);
	LUT4 #(
		.INIT('h0770)
	) name2204 (
		_w3193_,
		_w3194_,
		_w3197_,
		_w3198_,
		_w3207_
	);
	LUT3 #(
		.INIT('h01)
	) name2205 (
		_w3196_,
		_w3207_,
		_w3206_,
		_w3208_
	);
	LUT4 #(
		.INIT('hf770)
	) name2206 (
		_w3193_,
		_w3194_,
		_w3197_,
		_w3198_,
		_w3209_
	);
	LUT4 #(
		.INIT('h080f)
	) name2207 (
		_w3190_,
		_w3192_,
		_w3200_,
		_w3202_,
		_w3210_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		_w3201_,
		_w3210_,
		_w3211_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2209 (
		_w3205_,
		_w3208_,
		_w3209_,
		_w3211_,
		_w3212_
	);
	LUT3 #(
		.INIT('h96)
	) name2210 (
		\A[805] ,
		\A[806] ,
		\A[807] ,
		_w3213_
	);
	LUT3 #(
		.INIT('h96)
	) name2211 (
		\A[808] ,
		\A[809] ,
		\A[810] ,
		_w3214_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		_w3213_,
		_w3214_,
		_w3215_
	);
	LUT3 #(
		.INIT('h96)
	) name2213 (
		\A[799] ,
		\A[800] ,
		\A[801] ,
		_w3216_
	);
	LUT3 #(
		.INIT('h96)
	) name2214 (
		\A[802] ,
		\A[803] ,
		\A[804] ,
		_w3217_
	);
	LUT4 #(
		.INIT('h0660)
	) name2215 (
		_w3213_,
		_w3214_,
		_w3216_,
		_w3217_,
		_w3218_
	);
	LUT3 #(
		.INIT('h17)
	) name2216 (
		\A[808] ,
		\A[809] ,
		\A[810] ,
		_w3219_
	);
	LUT3 #(
		.INIT('h17)
	) name2217 (
		\A[805] ,
		\A[806] ,
		\A[807] ,
		_w3220_
	);
	LUT2 #(
		.INIT('h6)
	) name2218 (
		_w3219_,
		_w3220_,
		_w3221_
	);
	LUT3 #(
		.INIT('h17)
	) name2219 (
		\A[802] ,
		\A[803] ,
		\A[804] ,
		_w3222_
	);
	LUT3 #(
		.INIT('h17)
	) name2220 (
		\A[799] ,
		\A[800] ,
		\A[801] ,
		_w3223_
	);
	LUT4 #(
		.INIT('h7887)
	) name2221 (
		_w3216_,
		_w3217_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT4 #(
		.INIT('hc0de)
	) name2222 (
		_w3215_,
		_w3218_,
		_w3221_,
		_w3224_,
		_w3225_
	);
	LUT4 #(
		.INIT('h088f)
	) name2223 (
		_w3213_,
		_w3214_,
		_w3219_,
		_w3220_,
		_w3226_
	);
	LUT4 #(
		.INIT('h088f)
	) name2224 (
		_w3216_,
		_w3217_,
		_w3222_,
		_w3223_,
		_w3227_
	);
	LUT3 #(
		.INIT('he8)
	) name2225 (
		_w3225_,
		_w3226_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h4)
	) name2226 (
		_w3212_,
		_w3228_,
		_w3229_
	);
	LUT2 #(
		.INIT('h2)
	) name2227 (
		_w3212_,
		_w3228_,
		_w3230_
	);
	LUT2 #(
		.INIT('h9)
	) name2228 (
		_w3212_,
		_w3228_,
		_w3231_
	);
	LUT3 #(
		.INIT('h69)
	) name2229 (
		_w3225_,
		_w3226_,
		_w3227_,
		_w3232_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2230 (
		_w3205_,
		_w3208_,
		_w3209_,
		_w3211_,
		_w3233_
	);
	LUT4 #(
		.INIT('h6996)
	) name2231 (
		_w3190_,
		_w3192_,
		_w3193_,
		_w3194_,
		_w3234_
	);
	LUT4 #(
		.INIT('h6996)
	) name2232 (
		_w3213_,
		_w3214_,
		_w3216_,
		_w3217_,
		_w3235_
	);
	LUT2 #(
		.INIT('h8)
	) name2233 (
		_w3234_,
		_w3235_,
		_w3236_
	);
	LUT3 #(
		.INIT('h1e)
	) name2234 (
		_w3195_,
		_w3196_,
		_w3199_,
		_w3237_
	);
	LUT4 #(
		.INIT('he11e)
	) name2235 (
		_w3215_,
		_w3218_,
		_w3221_,
		_w3224_,
		_w3238_
	);
	LUT4 #(
		.INIT('hb721)
	) name2236 (
		_w3204_,
		_w3236_,
		_w3237_,
		_w3238_,
		_w3239_
	);
	LUT3 #(
		.INIT('hb2)
	) name2237 (
		_w3232_,
		_w3233_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h9)
	) name2238 (
		_w3231_,
		_w3240_,
		_w3241_
	);
	LUT3 #(
		.INIT('h96)
	) name2239 (
		_w3232_,
		_w3233_,
		_w3239_,
		_w3242_
	);
	LUT2 #(
		.INIT('h6)
	) name2240 (
		_w3176_,
		_w3177_,
		_w3243_
	);
	LUT4 #(
		.INIT('h0660)
	) name2241 (
		_w3180_,
		_w3181_,
		_w3234_,
		_w3235_,
		_w3244_
	);
	LUT3 #(
		.INIT('h96)
	) name2242 (
		_w3141_,
		_w3182_,
		_w3183_,
		_w3245_
	);
	LUT4 #(
		.INIT('h9669)
	) name2243 (
		_w3204_,
		_w3236_,
		_w3237_,
		_w3238_,
		_w3246_
	);
	LUT4 #(
		.INIT('h127b)
	) name2244 (
		_w3187_,
		_w3244_,
		_w3245_,
		_w3246_,
		_w3247_
	);
	LUT4 #(
		.INIT('h84ed)
	) name2245 (
		_w3188_,
		_w3242_,
		_w3243_,
		_w3247_,
		_w3248_
	);
	LUT3 #(
		.INIT('hd4)
	) name2246 (
		_w3189_,
		_w3241_,
		_w3248_,
		_w3249_
	);
	LUT4 #(
		.INIT('h4054)
	) name2247 (
		_w3174_,
		_w3176_,
		_w3177_,
		_w3188_,
		_w3250_
	);
	LUT2 #(
		.INIT('h1)
	) name2248 (
		_w3173_,
		_w3250_,
		_w3251_
	);
	LUT3 #(
		.INIT('h54)
	) name2249 (
		_w3229_,
		_w3230_,
		_w3240_,
		_w3252_
	);
	LUT3 #(
		.INIT('hd4)
	) name2250 (
		_w3249_,
		_w3251_,
		_w3252_,
		_w3253_
	);
	LUT3 #(
		.INIT('h96)
	) name2251 (
		\A[787] ,
		\A[788] ,
		\A[789] ,
		_w3254_
	);
	LUT2 #(
		.INIT('h8)
	) name2252 (
		\A[790] ,
		\A[791] ,
		_w3255_
	);
	LUT3 #(
		.INIT('h96)
	) name2253 (
		\A[790] ,
		\A[791] ,
		\A[792] ,
		_w3256_
	);
	LUT3 #(
		.INIT('h96)
	) name2254 (
		\A[793] ,
		\A[794] ,
		\A[795] ,
		_w3257_
	);
	LUT3 #(
		.INIT('h96)
	) name2255 (
		\A[796] ,
		\A[797] ,
		\A[798] ,
		_w3258_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		_w3257_,
		_w3258_,
		_w3259_
	);
	LUT4 #(
		.INIT('h0660)
	) name2257 (
		_w3254_,
		_w3256_,
		_w3257_,
		_w3258_,
		_w3260_
	);
	LUT3 #(
		.INIT('h17)
	) name2258 (
		\A[796] ,
		\A[797] ,
		\A[798] ,
		_w3261_
	);
	LUT3 #(
		.INIT('h17)
	) name2259 (
		\A[793] ,
		\A[794] ,
		\A[795] ,
		_w3262_
	);
	LUT2 #(
		.INIT('h6)
	) name2260 (
		_w3261_,
		_w3262_,
		_w3263_
	);
	LUT3 #(
		.INIT('h17)
	) name2261 (
		\A[787] ,
		\A[788] ,
		\A[789] ,
		_w3264_
	);
	LUT3 #(
		.INIT('h80)
	) name2262 (
		_w3254_,
		_w3255_,
		_w3256_,
		_w3265_
	);
	LUT3 #(
		.INIT('h17)
	) name2263 (
		\A[790] ,
		\A[791] ,
		\A[792] ,
		_w3266_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2264 (
		\A[790] ,
		\A[791] ,
		\A[792] ,
		_w3254_,
		_w3267_
	);
	LUT2 #(
		.INIT('h9)
	) name2265 (
		_w3264_,
		_w3267_,
		_w3268_
	);
	LUT4 #(
		.INIT('h0770)
	) name2266 (
		_w3260_,
		_w3263_,
		_w3264_,
		_w3267_,
		_w3269_
	);
	LUT4 #(
		.INIT('h8008)
	) name2267 (
		_w3257_,
		_w3258_,
		_w3261_,
		_w3262_,
		_w3270_
	);
	LUT4 #(
		.INIT('h0770)
	) name2268 (
		_w3257_,
		_w3258_,
		_w3261_,
		_w3262_,
		_w3271_
	);
	LUT3 #(
		.INIT('h01)
	) name2269 (
		_w3260_,
		_w3271_,
		_w3270_,
		_w3272_
	);
	LUT4 #(
		.INIT('hf770)
	) name2270 (
		_w3257_,
		_w3258_,
		_w3261_,
		_w3262_,
		_w3273_
	);
	LUT4 #(
		.INIT('h080f)
	) name2271 (
		_w3254_,
		_w3256_,
		_w3264_,
		_w3266_,
		_w3274_
	);
	LUT2 #(
		.INIT('h1)
	) name2272 (
		_w3265_,
		_w3274_,
		_w3275_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2273 (
		_w3269_,
		_w3272_,
		_w3273_,
		_w3275_,
		_w3276_
	);
	LUT3 #(
		.INIT('h96)
	) name2274 (
		\A[775] ,
		\A[776] ,
		\A[777] ,
		_w3277_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		\A[778] ,
		\A[779] ,
		_w3278_
	);
	LUT3 #(
		.INIT('h96)
	) name2276 (
		\A[778] ,
		\A[779] ,
		\A[780] ,
		_w3279_
	);
	LUT3 #(
		.INIT('h96)
	) name2277 (
		\A[781] ,
		\A[782] ,
		\A[783] ,
		_w3280_
	);
	LUT3 #(
		.INIT('h96)
	) name2278 (
		\A[784] ,
		\A[785] ,
		\A[786] ,
		_w3281_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w3280_,
		_w3281_,
		_w3282_
	);
	LUT4 #(
		.INIT('h0660)
	) name2280 (
		_w3277_,
		_w3279_,
		_w3280_,
		_w3281_,
		_w3283_
	);
	LUT3 #(
		.INIT('h17)
	) name2281 (
		\A[784] ,
		\A[785] ,
		\A[786] ,
		_w3284_
	);
	LUT3 #(
		.INIT('h17)
	) name2282 (
		\A[781] ,
		\A[782] ,
		\A[783] ,
		_w3285_
	);
	LUT2 #(
		.INIT('h6)
	) name2283 (
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT3 #(
		.INIT('h17)
	) name2284 (
		\A[775] ,
		\A[776] ,
		\A[777] ,
		_w3287_
	);
	LUT3 #(
		.INIT('h80)
	) name2285 (
		_w3277_,
		_w3278_,
		_w3279_,
		_w3288_
	);
	LUT3 #(
		.INIT('h17)
	) name2286 (
		\A[778] ,
		\A[779] ,
		\A[780] ,
		_w3289_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2287 (
		\A[778] ,
		\A[779] ,
		\A[780] ,
		_w3277_,
		_w3290_
	);
	LUT2 #(
		.INIT('h9)
	) name2288 (
		_w3287_,
		_w3290_,
		_w3291_
	);
	LUT4 #(
		.INIT('h0770)
	) name2289 (
		_w3283_,
		_w3286_,
		_w3287_,
		_w3290_,
		_w3292_
	);
	LUT4 #(
		.INIT('h8008)
	) name2290 (
		_w3280_,
		_w3281_,
		_w3284_,
		_w3285_,
		_w3293_
	);
	LUT4 #(
		.INIT('h0770)
	) name2291 (
		_w3280_,
		_w3281_,
		_w3284_,
		_w3285_,
		_w3294_
	);
	LUT3 #(
		.INIT('h01)
	) name2292 (
		_w3283_,
		_w3294_,
		_w3293_,
		_w3295_
	);
	LUT4 #(
		.INIT('hf770)
	) name2293 (
		_w3280_,
		_w3281_,
		_w3284_,
		_w3285_,
		_w3296_
	);
	LUT4 #(
		.INIT('h080f)
	) name2294 (
		_w3277_,
		_w3279_,
		_w3287_,
		_w3289_,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w3288_,
		_w3297_,
		_w3298_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2296 (
		_w3292_,
		_w3295_,
		_w3296_,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w3276_,
		_w3299_,
		_w3300_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		_w3276_,
		_w3299_,
		_w3301_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2299 (
		_w3292_,
		_w3295_,
		_w3296_,
		_w3298_,
		_w3302_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2300 (
		_w3269_,
		_w3272_,
		_w3273_,
		_w3275_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name2301 (
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		_w3302_,
		_w3303_,
		_w3305_
	);
	LUT4 #(
		.INIT('h6996)
	) name2303 (
		_w3254_,
		_w3256_,
		_w3257_,
		_w3258_,
		_w3306_
	);
	LUT4 #(
		.INIT('h6996)
	) name2304 (
		_w3277_,
		_w3279_,
		_w3280_,
		_w3281_,
		_w3307_
	);
	LUT2 #(
		.INIT('h8)
	) name2305 (
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT3 #(
		.INIT('h1e)
	) name2306 (
		_w3259_,
		_w3260_,
		_w3263_,
		_w3309_
	);
	LUT3 #(
		.INIT('h48)
	) name2307 (
		_w3268_,
		_w3308_,
		_w3309_,
		_w3310_
	);
	LUT3 #(
		.INIT('h21)
	) name2308 (
		_w3268_,
		_w3308_,
		_w3309_,
		_w3311_
	);
	LUT3 #(
		.INIT('h1e)
	) name2309 (
		_w3282_,
		_w3283_,
		_w3286_,
		_w3312_
	);
	LUT2 #(
		.INIT('h9)
	) name2310 (
		_w3291_,
		_w3312_,
		_w3313_
	);
	LUT3 #(
		.INIT('h54)
	) name2311 (
		_w3310_,
		_w3311_,
		_w3313_,
		_w3314_
	);
	LUT4 #(
		.INIT('h4054)
	) name2312 (
		_w3301_,
		_w3302_,
		_w3303_,
		_w3314_,
		_w3315_
	);
	LUT3 #(
		.INIT('h96)
	) name2313 (
		\A[757] ,
		\A[758] ,
		\A[759] ,
		_w3316_
	);
	LUT3 #(
		.INIT('h96)
	) name2314 (
		\A[760] ,
		\A[761] ,
		\A[762] ,
		_w3317_
	);
	LUT2 #(
		.INIT('h8)
	) name2315 (
		_w3316_,
		_w3317_,
		_w3318_
	);
	LUT3 #(
		.INIT('h96)
	) name2316 (
		\A[751] ,
		\A[752] ,
		\A[753] ,
		_w3319_
	);
	LUT3 #(
		.INIT('h96)
	) name2317 (
		\A[754] ,
		\A[755] ,
		\A[756] ,
		_w3320_
	);
	LUT4 #(
		.INIT('h0660)
	) name2318 (
		_w3316_,
		_w3317_,
		_w3319_,
		_w3320_,
		_w3321_
	);
	LUT3 #(
		.INIT('h17)
	) name2319 (
		\A[760] ,
		\A[761] ,
		\A[762] ,
		_w3322_
	);
	LUT3 #(
		.INIT('h17)
	) name2320 (
		\A[757] ,
		\A[758] ,
		\A[759] ,
		_w3323_
	);
	LUT2 #(
		.INIT('h6)
	) name2321 (
		_w3322_,
		_w3323_,
		_w3324_
	);
	LUT3 #(
		.INIT('h17)
	) name2322 (
		\A[754] ,
		\A[755] ,
		\A[756] ,
		_w3325_
	);
	LUT3 #(
		.INIT('h17)
	) name2323 (
		\A[751] ,
		\A[752] ,
		\A[753] ,
		_w3326_
	);
	LUT4 #(
		.INIT('h7887)
	) name2324 (
		_w3319_,
		_w3320_,
		_w3325_,
		_w3326_,
		_w3327_
	);
	LUT4 #(
		.INIT('hc0de)
	) name2325 (
		_w3318_,
		_w3321_,
		_w3324_,
		_w3327_,
		_w3328_
	);
	LUT4 #(
		.INIT('h088f)
	) name2326 (
		_w3319_,
		_w3320_,
		_w3325_,
		_w3326_,
		_w3329_
	);
	LUT4 #(
		.INIT('h088f)
	) name2327 (
		_w3316_,
		_w3317_,
		_w3322_,
		_w3323_,
		_w3330_
	);
	LUT3 #(
		.INIT('h69)
	) name2328 (
		_w3328_,
		_w3329_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		\A[766] ,
		\A[767] ,
		_w3332_
	);
	LUT3 #(
		.INIT('h96)
	) name2330 (
		\A[763] ,
		\A[764] ,
		\A[765] ,
		_w3333_
	);
	LUT3 #(
		.INIT('h96)
	) name2331 (
		\A[766] ,
		\A[767] ,
		\A[768] ,
		_w3334_
	);
	LUT3 #(
		.INIT('h80)
	) name2332 (
		_w3332_,
		_w3333_,
		_w3334_,
		_w3335_
	);
	LUT3 #(
		.INIT('h17)
	) name2333 (
		\A[763] ,
		\A[764] ,
		\A[765] ,
		_w3336_
	);
	LUT3 #(
		.INIT('h17)
	) name2334 (
		\A[766] ,
		\A[767] ,
		\A[768] ,
		_w3337_
	);
	LUT4 #(
		.INIT('h080f)
	) name2335 (
		_w3333_,
		_w3334_,
		_w3336_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w3335_,
		_w3338_,
		_w3339_
	);
	LUT3 #(
		.INIT('h17)
	) name2337 (
		\A[772] ,
		\A[773] ,
		\A[774] ,
		_w3340_
	);
	LUT3 #(
		.INIT('h17)
	) name2338 (
		\A[769] ,
		\A[770] ,
		\A[771] ,
		_w3341_
	);
	LUT3 #(
		.INIT('h96)
	) name2339 (
		\A[769] ,
		\A[770] ,
		\A[771] ,
		_w3342_
	);
	LUT3 #(
		.INIT('h96)
	) name2340 (
		\A[772] ,
		\A[773] ,
		\A[774] ,
		_w3343_
	);
	LUT4 #(
		.INIT('h7111)
	) name2341 (
		_w3340_,
		_w3341_,
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT4 #(
		.INIT('h0660)
	) name2342 (
		_w3333_,
		_w3334_,
		_w3342_,
		_w3343_,
		_w3345_
	);
	LUT4 #(
		.INIT('h0080)
	) name2343 (
		_w3332_,
		_w3333_,
		_w3334_,
		_w3336_,
		_w3346_
	);
	LUT2 #(
		.INIT('h2)
	) name2344 (
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT4 #(
		.INIT('h6999)
	) name2345 (
		_w3340_,
		_w3341_,
		_w3342_,
		_w3343_,
		_w3348_
	);
	LUT3 #(
		.INIT('h02)
	) name2346 (
		_w3345_,
		_w3346_,
		_w3348_,
		_w3349_
	);
	LUT3 #(
		.INIT('hd0)
	) name2347 (
		_w3345_,
		_w3346_,
		_w3348_,
		_w3350_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2348 (
		\A[766] ,
		\A[767] ,
		\A[768] ,
		_w3333_,
		_w3351_
	);
	LUT2 #(
		.INIT('h9)
	) name2349 (
		_w3336_,
		_w3351_,
		_w3352_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2350 (
		_w3344_,
		_w3347_,
		_w3348_,
		_w3352_,
		_w3353_
	);
	LUT4 #(
		.INIT('h1051)
	) name2351 (
		_w3344_,
		_w3347_,
		_w3348_,
		_w3352_,
		_w3354_
	);
	LUT4 #(
		.INIT('h6566)
	) name2352 (
		_w3344_,
		_w3349_,
		_w3350_,
		_w3352_,
		_w3355_
	);
	LUT4 #(
		.INIT('h6996)
	) name2353 (
		_w3333_,
		_w3334_,
		_w3342_,
		_w3343_,
		_w3356_
	);
	LUT4 #(
		.INIT('h6996)
	) name2354 (
		_w3316_,
		_w3317_,
		_w3319_,
		_w3320_,
		_w3357_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		_w3356_,
		_w3357_,
		_w3358_
	);
	LUT3 #(
		.INIT('h2d)
	) name2356 (
		_w3345_,
		_w3346_,
		_w3348_,
		_w3359_
	);
	LUT4 #(
		.INIT('he11e)
	) name2357 (
		_w3318_,
		_w3321_,
		_w3324_,
		_w3327_,
		_w3360_
	);
	LUT4 #(
		.INIT('hb721)
	) name2358 (
		_w3352_,
		_w3358_,
		_w3359_,
		_w3360_,
		_w3361_
	);
	LUT4 #(
		.INIT('hbe28)
	) name2359 (
		_w3331_,
		_w3339_,
		_w3355_,
		_w3361_,
		_w3362_
	);
	LUT3 #(
		.INIT('h32)
	) name2360 (
		_w3339_,
		_w3353_,
		_w3354_,
		_w3363_
	);
	LUT3 #(
		.INIT('he8)
	) name2361 (
		_w3328_,
		_w3329_,
		_w3330_,
		_w3364_
	);
	LUT3 #(
		.INIT('h71)
	) name2362 (
		_w3362_,
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT3 #(
		.INIT('he0)
	) name2363 (
		_w3300_,
		_w3315_,
		_w3365_,
		_w3366_
	);
	LUT3 #(
		.INIT('h01)
	) name2364 (
		_w3300_,
		_w3315_,
		_w3365_,
		_w3367_
	);
	LUT2 #(
		.INIT('h6)
	) name2365 (
		_w3276_,
		_w3299_,
		_w3368_
	);
	LUT4 #(
		.INIT('h45ba)
	) name2366 (
		_w3304_,
		_w3305_,
		_w3314_,
		_w3368_,
		_w3369_
	);
	LUT3 #(
		.INIT('h69)
	) name2367 (
		_w3362_,
		_w3363_,
		_w3364_,
		_w3370_
	);
	LUT4 #(
		.INIT('h9669)
	) name2368 (
		_w3331_,
		_w3339_,
		_w3355_,
		_w3361_,
		_w3371_
	);
	LUT2 #(
		.INIT('h6)
	) name2369 (
		_w3302_,
		_w3303_,
		_w3372_
	);
	LUT4 #(
		.INIT('h0660)
	) name2370 (
		_w3306_,
		_w3307_,
		_w3356_,
		_w3357_,
		_w3373_
	);
	LUT3 #(
		.INIT('h96)
	) name2371 (
		_w3268_,
		_w3308_,
		_w3309_,
		_w3374_
	);
	LUT4 #(
		.INIT('h9669)
	) name2372 (
		_w3352_,
		_w3358_,
		_w3359_,
		_w3360_,
		_w3375_
	);
	LUT4 #(
		.INIT('h127b)
	) name2373 (
		_w3313_,
		_w3373_,
		_w3374_,
		_w3375_,
		_w3376_
	);
	LUT4 #(
		.INIT('h84ed)
	) name2374 (
		_w3314_,
		_w3371_,
		_w3372_,
		_w3376_,
		_w3377_
	);
	LUT3 #(
		.INIT('h8e)
	) name2375 (
		_w3369_,
		_w3370_,
		_w3377_,
		_w3378_
	);
	LUT3 #(
		.INIT('h54)
	) name2376 (
		_w3366_,
		_w3367_,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w3253_,
		_w3379_,
		_w3380_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		_w3253_,
		_w3379_,
		_w3381_
	);
	LUT3 #(
		.INIT('h1e)
	) name2379 (
		_w3300_,
		_w3315_,
		_w3365_,
		_w3382_
	);
	LUT2 #(
		.INIT('h9)
	) name2380 (
		_w3378_,
		_w3382_,
		_w3383_
	);
	LUT3 #(
		.INIT('h69)
	) name2381 (
		_w3249_,
		_w3251_,
		_w3252_,
		_w3384_
	);
	LUT3 #(
		.INIT('h96)
	) name2382 (
		_w3189_,
		_w3241_,
		_w3248_,
		_w3385_
	);
	LUT3 #(
		.INIT('h96)
	) name2383 (
		_w3369_,
		_w3370_,
		_w3377_,
		_w3386_
	);
	LUT4 #(
		.INIT('h6996)
	) name2384 (
		_w3314_,
		_w3371_,
		_w3372_,
		_w3376_,
		_w3387_
	);
	LUT4 #(
		.INIT('h6996)
	) name2385 (
		_w3188_,
		_w3242_,
		_w3243_,
		_w3247_,
		_w3388_
	);
	LUT4 #(
		.INIT('h6996)
	) name2386 (
		_w3180_,
		_w3181_,
		_w3234_,
		_w3235_,
		_w3389_
	);
	LUT4 #(
		.INIT('h6996)
	) name2387 (
		_w3306_,
		_w3307_,
		_w3356_,
		_w3357_,
		_w3390_
	);
	LUT2 #(
		.INIT('h8)
	) name2388 (
		_w3389_,
		_w3390_,
		_w3391_
	);
	LUT4 #(
		.INIT('h6996)
	) name2389 (
		_w3187_,
		_w3244_,
		_w3245_,
		_w3246_,
		_w3392_
	);
	LUT4 #(
		.INIT('h6996)
	) name2390 (
		_w3313_,
		_w3373_,
		_w3374_,
		_w3375_,
		_w3393_
	);
	LUT3 #(
		.INIT('hd4)
	) name2391 (
		_w3391_,
		_w3392_,
		_w3393_,
		_w3394_
	);
	LUT3 #(
		.INIT('h8e)
	) name2392 (
		_w3387_,
		_w3388_,
		_w3394_,
		_w3395_
	);
	LUT3 #(
		.INIT('hd4)
	) name2393 (
		_w3385_,
		_w3386_,
		_w3395_,
		_w3396_
	);
	LUT3 #(
		.INIT('h4d)
	) name2394 (
		_w3383_,
		_w3384_,
		_w3396_,
		_w3397_
	);
	LUT3 #(
		.INIT('h54)
	) name2395 (
		_w3380_,
		_w3381_,
		_w3397_,
		_w3398_
	);
	LUT3 #(
		.INIT('h96)
	) name2396 (
		\A[739] ,
		\A[740] ,
		\A[741] ,
		_w3399_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		\A[742] ,
		\A[743] ,
		_w3400_
	);
	LUT3 #(
		.INIT('h96)
	) name2398 (
		\A[742] ,
		\A[743] ,
		\A[744] ,
		_w3401_
	);
	LUT3 #(
		.INIT('h96)
	) name2399 (
		\A[745] ,
		\A[746] ,
		\A[747] ,
		_w3402_
	);
	LUT3 #(
		.INIT('h96)
	) name2400 (
		\A[748] ,
		\A[749] ,
		\A[750] ,
		_w3403_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		_w3402_,
		_w3403_,
		_w3404_
	);
	LUT4 #(
		.INIT('h0660)
	) name2402 (
		_w3399_,
		_w3401_,
		_w3402_,
		_w3403_,
		_w3405_
	);
	LUT3 #(
		.INIT('h17)
	) name2403 (
		\A[748] ,
		\A[749] ,
		\A[750] ,
		_w3406_
	);
	LUT3 #(
		.INIT('h17)
	) name2404 (
		\A[745] ,
		\A[746] ,
		\A[747] ,
		_w3407_
	);
	LUT2 #(
		.INIT('h6)
	) name2405 (
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT3 #(
		.INIT('h17)
	) name2406 (
		\A[739] ,
		\A[740] ,
		\A[741] ,
		_w3409_
	);
	LUT3 #(
		.INIT('h80)
	) name2407 (
		_w3399_,
		_w3400_,
		_w3401_,
		_w3410_
	);
	LUT3 #(
		.INIT('h17)
	) name2408 (
		\A[742] ,
		\A[743] ,
		\A[744] ,
		_w3411_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2409 (
		\A[742] ,
		\A[743] ,
		\A[744] ,
		_w3399_,
		_w3412_
	);
	LUT2 #(
		.INIT('h9)
	) name2410 (
		_w3409_,
		_w3412_,
		_w3413_
	);
	LUT4 #(
		.INIT('h0770)
	) name2411 (
		_w3405_,
		_w3408_,
		_w3409_,
		_w3412_,
		_w3414_
	);
	LUT4 #(
		.INIT('h8008)
	) name2412 (
		_w3402_,
		_w3403_,
		_w3406_,
		_w3407_,
		_w3415_
	);
	LUT4 #(
		.INIT('h0770)
	) name2413 (
		_w3402_,
		_w3403_,
		_w3406_,
		_w3407_,
		_w3416_
	);
	LUT3 #(
		.INIT('h01)
	) name2414 (
		_w3405_,
		_w3416_,
		_w3415_,
		_w3417_
	);
	LUT4 #(
		.INIT('hf770)
	) name2415 (
		_w3402_,
		_w3403_,
		_w3406_,
		_w3407_,
		_w3418_
	);
	LUT4 #(
		.INIT('h080f)
	) name2416 (
		_w3399_,
		_w3401_,
		_w3409_,
		_w3411_,
		_w3419_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		_w3410_,
		_w3419_,
		_w3420_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2418 (
		_w3414_,
		_w3417_,
		_w3418_,
		_w3420_,
		_w3421_
	);
	LUT3 #(
		.INIT('h96)
	) name2419 (
		\A[727] ,
		\A[728] ,
		\A[729] ,
		_w3422_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		\A[730] ,
		\A[731] ,
		_w3423_
	);
	LUT3 #(
		.INIT('h96)
	) name2421 (
		\A[730] ,
		\A[731] ,
		\A[732] ,
		_w3424_
	);
	LUT3 #(
		.INIT('h96)
	) name2422 (
		\A[733] ,
		\A[734] ,
		\A[735] ,
		_w3425_
	);
	LUT3 #(
		.INIT('h96)
	) name2423 (
		\A[736] ,
		\A[737] ,
		\A[738] ,
		_w3426_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		_w3425_,
		_w3426_,
		_w3427_
	);
	LUT4 #(
		.INIT('h0660)
	) name2425 (
		_w3422_,
		_w3424_,
		_w3425_,
		_w3426_,
		_w3428_
	);
	LUT3 #(
		.INIT('h17)
	) name2426 (
		\A[736] ,
		\A[737] ,
		\A[738] ,
		_w3429_
	);
	LUT3 #(
		.INIT('h17)
	) name2427 (
		\A[733] ,
		\A[734] ,
		\A[735] ,
		_w3430_
	);
	LUT2 #(
		.INIT('h6)
	) name2428 (
		_w3429_,
		_w3430_,
		_w3431_
	);
	LUT3 #(
		.INIT('h17)
	) name2429 (
		\A[727] ,
		\A[728] ,
		\A[729] ,
		_w3432_
	);
	LUT3 #(
		.INIT('h80)
	) name2430 (
		_w3422_,
		_w3423_,
		_w3424_,
		_w3433_
	);
	LUT3 #(
		.INIT('h17)
	) name2431 (
		\A[730] ,
		\A[731] ,
		\A[732] ,
		_w3434_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2432 (
		\A[730] ,
		\A[731] ,
		\A[732] ,
		_w3422_,
		_w3435_
	);
	LUT2 #(
		.INIT('h9)
	) name2433 (
		_w3432_,
		_w3435_,
		_w3436_
	);
	LUT4 #(
		.INIT('h0770)
	) name2434 (
		_w3428_,
		_w3431_,
		_w3432_,
		_w3435_,
		_w3437_
	);
	LUT4 #(
		.INIT('h8008)
	) name2435 (
		_w3425_,
		_w3426_,
		_w3429_,
		_w3430_,
		_w3438_
	);
	LUT4 #(
		.INIT('h0770)
	) name2436 (
		_w3425_,
		_w3426_,
		_w3429_,
		_w3430_,
		_w3439_
	);
	LUT3 #(
		.INIT('h01)
	) name2437 (
		_w3428_,
		_w3439_,
		_w3438_,
		_w3440_
	);
	LUT4 #(
		.INIT('hf770)
	) name2438 (
		_w3425_,
		_w3426_,
		_w3429_,
		_w3430_,
		_w3441_
	);
	LUT4 #(
		.INIT('h080f)
	) name2439 (
		_w3422_,
		_w3424_,
		_w3432_,
		_w3434_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		_w3433_,
		_w3442_,
		_w3443_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2441 (
		_w3437_,
		_w3440_,
		_w3441_,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h1)
	) name2442 (
		_w3421_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h8)
	) name2443 (
		_w3421_,
		_w3444_,
		_w3446_
	);
	LUT2 #(
		.INIT('h6)
	) name2444 (
		_w3421_,
		_w3444_,
		_w3447_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2445 (
		_w3437_,
		_w3440_,
		_w3441_,
		_w3443_,
		_w3448_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2446 (
		_w3414_,
		_w3417_,
		_w3418_,
		_w3420_,
		_w3449_
	);
	LUT2 #(
		.INIT('h1)
	) name2447 (
		_w3448_,
		_w3449_,
		_w3450_
	);
	LUT2 #(
		.INIT('h8)
	) name2448 (
		_w3448_,
		_w3449_,
		_w3451_
	);
	LUT4 #(
		.INIT('h6996)
	) name2449 (
		_w3399_,
		_w3401_,
		_w3402_,
		_w3403_,
		_w3452_
	);
	LUT4 #(
		.INIT('h6996)
	) name2450 (
		_w3422_,
		_w3424_,
		_w3425_,
		_w3426_,
		_w3453_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		_w3452_,
		_w3453_,
		_w3454_
	);
	LUT3 #(
		.INIT('h1e)
	) name2452 (
		_w3404_,
		_w3405_,
		_w3408_,
		_w3455_
	);
	LUT3 #(
		.INIT('h48)
	) name2453 (
		_w3413_,
		_w3454_,
		_w3455_,
		_w3456_
	);
	LUT3 #(
		.INIT('h21)
	) name2454 (
		_w3413_,
		_w3454_,
		_w3455_,
		_w3457_
	);
	LUT3 #(
		.INIT('h1e)
	) name2455 (
		_w3427_,
		_w3428_,
		_w3431_,
		_w3458_
	);
	LUT2 #(
		.INIT('h9)
	) name2456 (
		_w3436_,
		_w3458_,
		_w3459_
	);
	LUT3 #(
		.INIT('h54)
	) name2457 (
		_w3456_,
		_w3457_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('h6566)
	) name2458 (
		_w3447_,
		_w3450_,
		_w3451_,
		_w3460_,
		_w3461_
	);
	LUT3 #(
		.INIT('h96)
	) name2459 (
		\A[715] ,
		\A[716] ,
		\A[717] ,
		_w3462_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		\A[718] ,
		\A[719] ,
		_w3463_
	);
	LUT3 #(
		.INIT('h96)
	) name2461 (
		\A[718] ,
		\A[719] ,
		\A[720] ,
		_w3464_
	);
	LUT3 #(
		.INIT('h96)
	) name2462 (
		\A[721] ,
		\A[722] ,
		\A[723] ,
		_w3465_
	);
	LUT3 #(
		.INIT('h96)
	) name2463 (
		\A[724] ,
		\A[725] ,
		\A[726] ,
		_w3466_
	);
	LUT2 #(
		.INIT('h8)
	) name2464 (
		_w3465_,
		_w3466_,
		_w3467_
	);
	LUT4 #(
		.INIT('h0660)
	) name2465 (
		_w3462_,
		_w3464_,
		_w3465_,
		_w3466_,
		_w3468_
	);
	LUT3 #(
		.INIT('h17)
	) name2466 (
		\A[724] ,
		\A[725] ,
		\A[726] ,
		_w3469_
	);
	LUT3 #(
		.INIT('h17)
	) name2467 (
		\A[721] ,
		\A[722] ,
		\A[723] ,
		_w3470_
	);
	LUT2 #(
		.INIT('h6)
	) name2468 (
		_w3469_,
		_w3470_,
		_w3471_
	);
	LUT3 #(
		.INIT('h17)
	) name2469 (
		\A[715] ,
		\A[716] ,
		\A[717] ,
		_w3472_
	);
	LUT3 #(
		.INIT('h80)
	) name2470 (
		_w3462_,
		_w3463_,
		_w3464_,
		_w3473_
	);
	LUT3 #(
		.INIT('h17)
	) name2471 (
		\A[718] ,
		\A[719] ,
		\A[720] ,
		_w3474_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2472 (
		\A[718] ,
		\A[719] ,
		\A[720] ,
		_w3462_,
		_w3475_
	);
	LUT2 #(
		.INIT('h9)
	) name2473 (
		_w3472_,
		_w3475_,
		_w3476_
	);
	LUT4 #(
		.INIT('h0770)
	) name2474 (
		_w3468_,
		_w3471_,
		_w3472_,
		_w3475_,
		_w3477_
	);
	LUT4 #(
		.INIT('h8008)
	) name2475 (
		_w3465_,
		_w3466_,
		_w3469_,
		_w3470_,
		_w3478_
	);
	LUT4 #(
		.INIT('h0770)
	) name2476 (
		_w3465_,
		_w3466_,
		_w3469_,
		_w3470_,
		_w3479_
	);
	LUT3 #(
		.INIT('h01)
	) name2477 (
		_w3468_,
		_w3479_,
		_w3478_,
		_w3480_
	);
	LUT4 #(
		.INIT('hf770)
	) name2478 (
		_w3465_,
		_w3466_,
		_w3469_,
		_w3470_,
		_w3481_
	);
	LUT4 #(
		.INIT('h080f)
	) name2479 (
		_w3462_,
		_w3464_,
		_w3472_,
		_w3474_,
		_w3482_
	);
	LUT2 #(
		.INIT('h1)
	) name2480 (
		_w3473_,
		_w3482_,
		_w3483_
	);
	LUT4 #(
		.INIT('hfee0)
	) name2481 (
		_w3477_,
		_w3480_,
		_w3481_,
		_w3483_,
		_w3484_
	);
	LUT3 #(
		.INIT('h96)
	) name2482 (
		\A[709] ,
		\A[710] ,
		\A[711] ,
		_w3485_
	);
	LUT3 #(
		.INIT('h96)
	) name2483 (
		\A[712] ,
		\A[713] ,
		\A[714] ,
		_w3486_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		_w3485_,
		_w3486_,
		_w3487_
	);
	LUT3 #(
		.INIT('h96)
	) name2485 (
		\A[703] ,
		\A[704] ,
		\A[705] ,
		_w3488_
	);
	LUT3 #(
		.INIT('h96)
	) name2486 (
		\A[706] ,
		\A[707] ,
		\A[708] ,
		_w3489_
	);
	LUT4 #(
		.INIT('h0660)
	) name2487 (
		_w3485_,
		_w3486_,
		_w3488_,
		_w3489_,
		_w3490_
	);
	LUT3 #(
		.INIT('h17)
	) name2488 (
		\A[712] ,
		\A[713] ,
		\A[714] ,
		_w3491_
	);
	LUT3 #(
		.INIT('h17)
	) name2489 (
		\A[709] ,
		\A[710] ,
		\A[711] ,
		_w3492_
	);
	LUT2 #(
		.INIT('h6)
	) name2490 (
		_w3491_,
		_w3492_,
		_w3493_
	);
	LUT3 #(
		.INIT('h17)
	) name2491 (
		\A[706] ,
		\A[707] ,
		\A[708] ,
		_w3494_
	);
	LUT3 #(
		.INIT('h17)
	) name2492 (
		\A[703] ,
		\A[704] ,
		\A[705] ,
		_w3495_
	);
	LUT4 #(
		.INIT('h7887)
	) name2493 (
		_w3488_,
		_w3489_,
		_w3494_,
		_w3495_,
		_w3496_
	);
	LUT4 #(
		.INIT('hc0de)
	) name2494 (
		_w3487_,
		_w3490_,
		_w3493_,
		_w3496_,
		_w3497_
	);
	LUT4 #(
		.INIT('h088f)
	) name2495 (
		_w3485_,
		_w3486_,
		_w3491_,
		_w3492_,
		_w3498_
	);
	LUT4 #(
		.INIT('h088f)
	) name2496 (
		_w3488_,
		_w3489_,
		_w3494_,
		_w3495_,
		_w3499_
	);
	LUT3 #(
		.INIT('he8)
	) name2497 (
		_w3497_,
		_w3498_,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('h4)
	) name2498 (
		_w3484_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h2)
	) name2499 (
		_w3484_,
		_w3500_,
		_w3502_
	);
	LUT2 #(
		.INIT('h9)
	) name2500 (
		_w3484_,
		_w3500_,
		_w3503_
	);
	LUT3 #(
		.INIT('h69)
	) name2501 (
		_w3497_,
		_w3498_,
		_w3499_,
		_w3504_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2502 (
		_w3477_,
		_w3480_,
		_w3481_,
		_w3483_,
		_w3505_
	);
	LUT4 #(
		.INIT('h6996)
	) name2503 (
		_w3462_,
		_w3464_,
		_w3465_,
		_w3466_,
		_w3506_
	);
	LUT4 #(
		.INIT('h6996)
	) name2504 (
		_w3485_,
		_w3486_,
		_w3488_,
		_w3489_,
		_w3507_
	);
	LUT2 #(
		.INIT('h8)
	) name2505 (
		_w3506_,
		_w3507_,
		_w3508_
	);
	LUT3 #(
		.INIT('h1e)
	) name2506 (
		_w3467_,
		_w3468_,
		_w3471_,
		_w3509_
	);
	LUT4 #(
		.INIT('he11e)
	) name2507 (
		_w3487_,
		_w3490_,
		_w3493_,
		_w3496_,
		_w3510_
	);
	LUT4 #(
		.INIT('hb721)
	) name2508 (
		_w3476_,
		_w3508_,
		_w3509_,
		_w3510_,
		_w3511_
	);
	LUT3 #(
		.INIT('hb2)
	) name2509 (
		_w3504_,
		_w3505_,
		_w3511_,
		_w3512_
	);
	LUT2 #(
		.INIT('h9)
	) name2510 (
		_w3503_,
		_w3512_,
		_w3513_
	);
	LUT3 #(
		.INIT('h96)
	) name2511 (
		_w3504_,
		_w3505_,
		_w3511_,
		_w3514_
	);
	LUT2 #(
		.INIT('h6)
	) name2512 (
		_w3448_,
		_w3449_,
		_w3515_
	);
	LUT4 #(
		.INIT('h0660)
	) name2513 (
		_w3452_,
		_w3453_,
		_w3506_,
		_w3507_,
		_w3516_
	);
	LUT3 #(
		.INIT('h96)
	) name2514 (
		_w3413_,
		_w3454_,
		_w3455_,
		_w3517_
	);
	LUT4 #(
		.INIT('h9669)
	) name2515 (
		_w3476_,
		_w3508_,
		_w3509_,
		_w3510_,
		_w3518_
	);
	LUT4 #(
		.INIT('h127b)
	) name2516 (
		_w3459_,
		_w3516_,
		_w3517_,
		_w3518_,
		_w3519_
	);
	LUT4 #(
		.INIT('h84ed)
	) name2517 (
		_w3460_,
		_w3514_,
		_w3515_,
		_w3519_,
		_w3520_
	);
	LUT3 #(
		.INIT('hd4)
	) name2518 (
		_w3461_,
		_w3513_,
		_w3520_,
		_w3521_
	);
	LUT4 #(
		.INIT('h4054)
	) name2519 (
		_w3446_,
		_w3448_,
		_w3449_,
		_w3460_,
		_w3522_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w3445_,
		_w3522_,
		_w3523_
	);
	LUT3 #(
		.INIT('h54)
	) name2521 (
		_w3501_,
		_w3502_,
		_w3512_,
		_w3524_
	);
	LUT3 #(
		.INIT('hd4)
	) name2522 (
		_w3521_,
		_w3523_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h8)
	) name2523 (
		\A[658] ,
		\A[659] ,
		_w3526_
	);
	LUT3 #(
		.INIT('h96)
	) name2524 (
		\A[655] ,
		\A[656] ,
		\A[657] ,
		_w3527_
	);
	LUT3 #(
		.INIT('h96)
	) name2525 (
		\A[658] ,
		\A[659] ,
		\A[660] ,
		_w3528_
	);
	LUT3 #(
		.INIT('h80)
	) name2526 (
		_w3526_,
		_w3527_,
		_w3528_,
		_w3529_
	);
	LUT3 #(
		.INIT('h17)
	) name2527 (
		\A[655] ,
		\A[656] ,
		\A[657] ,
		_w3530_
	);
	LUT3 #(
		.INIT('h17)
	) name2528 (
		\A[658] ,
		\A[659] ,
		\A[660] ,
		_w3531_
	);
	LUT4 #(
		.INIT('h080f)
	) name2529 (
		_w3527_,
		_w3528_,
		_w3530_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name2530 (
		_w3529_,
		_w3532_,
		_w3533_
	);
	LUT3 #(
		.INIT('h17)
	) name2531 (
		\A[664] ,
		\A[665] ,
		\A[666] ,
		_w3534_
	);
	LUT3 #(
		.INIT('h17)
	) name2532 (
		\A[661] ,
		\A[662] ,
		\A[663] ,
		_w3535_
	);
	LUT3 #(
		.INIT('h96)
	) name2533 (
		\A[661] ,
		\A[662] ,
		\A[663] ,
		_w3536_
	);
	LUT3 #(
		.INIT('h96)
	) name2534 (
		\A[664] ,
		\A[665] ,
		\A[666] ,
		_w3537_
	);
	LUT4 #(
		.INIT('h7111)
	) name2535 (
		_w3534_,
		_w3535_,
		_w3536_,
		_w3537_,
		_w3538_
	);
	LUT4 #(
		.INIT('h0660)
	) name2536 (
		_w3527_,
		_w3528_,
		_w3536_,
		_w3537_,
		_w3539_
	);
	LUT4 #(
		.INIT('h0080)
	) name2537 (
		_w3526_,
		_w3527_,
		_w3528_,
		_w3530_,
		_w3540_
	);
	LUT2 #(
		.INIT('h2)
	) name2538 (
		_w3539_,
		_w3540_,
		_w3541_
	);
	LUT4 #(
		.INIT('h6999)
	) name2539 (
		_w3534_,
		_w3535_,
		_w3536_,
		_w3537_,
		_w3542_
	);
	LUT3 #(
		.INIT('h02)
	) name2540 (
		_w3539_,
		_w3540_,
		_w3542_,
		_w3543_
	);
	LUT3 #(
		.INIT('hd0)
	) name2541 (
		_w3539_,
		_w3540_,
		_w3542_,
		_w3544_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2542 (
		\A[658] ,
		\A[659] ,
		\A[660] ,
		_w3527_,
		_w3545_
	);
	LUT2 #(
		.INIT('h9)
	) name2543 (
		_w3530_,
		_w3545_,
		_w3546_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2544 (
		_w3538_,
		_w3541_,
		_w3542_,
		_w3546_,
		_w3547_
	);
	LUT4 #(
		.INIT('h1051)
	) name2545 (
		_w3538_,
		_w3541_,
		_w3542_,
		_w3546_,
		_w3548_
	);
	LUT4 #(
		.INIT('h6566)
	) name2546 (
		_w3538_,
		_w3543_,
		_w3544_,
		_w3546_,
		_w3549_
	);
	LUT2 #(
		.INIT('h6)
	) name2547 (
		_w3533_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		\A[670] ,
		\A[671] ,
		_w3551_
	);
	LUT3 #(
		.INIT('h96)
	) name2549 (
		\A[667] ,
		\A[668] ,
		\A[669] ,
		_w3552_
	);
	LUT3 #(
		.INIT('h96)
	) name2550 (
		\A[670] ,
		\A[671] ,
		\A[672] ,
		_w3553_
	);
	LUT3 #(
		.INIT('h80)
	) name2551 (
		_w3551_,
		_w3552_,
		_w3553_,
		_w3554_
	);
	LUT3 #(
		.INIT('h17)
	) name2552 (
		\A[667] ,
		\A[668] ,
		\A[669] ,
		_w3555_
	);
	LUT3 #(
		.INIT('h17)
	) name2553 (
		\A[670] ,
		\A[671] ,
		\A[672] ,
		_w3556_
	);
	LUT4 #(
		.INIT('h080f)
	) name2554 (
		_w3552_,
		_w3553_,
		_w3555_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w3554_,
		_w3557_,
		_w3558_
	);
	LUT3 #(
		.INIT('h17)
	) name2556 (
		\A[676] ,
		\A[677] ,
		\A[678] ,
		_w3559_
	);
	LUT3 #(
		.INIT('h17)
	) name2557 (
		\A[673] ,
		\A[674] ,
		\A[675] ,
		_w3560_
	);
	LUT3 #(
		.INIT('h96)
	) name2558 (
		\A[673] ,
		\A[674] ,
		\A[675] ,
		_w3561_
	);
	LUT3 #(
		.INIT('h96)
	) name2559 (
		\A[676] ,
		\A[677] ,
		\A[678] ,
		_w3562_
	);
	LUT4 #(
		.INIT('h7111)
	) name2560 (
		_w3559_,
		_w3560_,
		_w3561_,
		_w3562_,
		_w3563_
	);
	LUT4 #(
		.INIT('h0660)
	) name2561 (
		_w3552_,
		_w3553_,
		_w3561_,
		_w3562_,
		_w3564_
	);
	LUT4 #(
		.INIT('h0080)
	) name2562 (
		_w3551_,
		_w3552_,
		_w3553_,
		_w3555_,
		_w3565_
	);
	LUT2 #(
		.INIT('h2)
	) name2563 (
		_w3564_,
		_w3565_,
		_w3566_
	);
	LUT4 #(
		.INIT('h6999)
	) name2564 (
		_w3559_,
		_w3560_,
		_w3561_,
		_w3562_,
		_w3567_
	);
	LUT3 #(
		.INIT('h02)
	) name2565 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w3568_
	);
	LUT3 #(
		.INIT('hd0)
	) name2566 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w3569_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2567 (
		\A[670] ,
		\A[671] ,
		\A[672] ,
		_w3552_,
		_w3570_
	);
	LUT2 #(
		.INIT('h9)
	) name2568 (
		_w3555_,
		_w3570_,
		_w3571_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2569 (
		_w3563_,
		_w3566_,
		_w3567_,
		_w3571_,
		_w3572_
	);
	LUT4 #(
		.INIT('h1051)
	) name2570 (
		_w3563_,
		_w3566_,
		_w3567_,
		_w3571_,
		_w3573_
	);
	LUT4 #(
		.INIT('h6566)
	) name2571 (
		_w3563_,
		_w3568_,
		_w3569_,
		_w3571_,
		_w3574_
	);
	LUT2 #(
		.INIT('h6)
	) name2572 (
		_w3558_,
		_w3574_,
		_w3575_
	);
	LUT4 #(
		.INIT('h9009)
	) name2573 (
		_w3533_,
		_w3549_,
		_w3558_,
		_w3574_,
		_w3576_
	);
	LUT4 #(
		.INIT('h0660)
	) name2574 (
		_w3533_,
		_w3549_,
		_w3558_,
		_w3574_,
		_w3577_
	);
	LUT4 #(
		.INIT('h6996)
	) name2575 (
		_w3552_,
		_w3553_,
		_w3561_,
		_w3562_,
		_w3578_
	);
	LUT4 #(
		.INIT('h6996)
	) name2576 (
		_w3527_,
		_w3528_,
		_w3536_,
		_w3537_,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name2577 (
		_w3578_,
		_w3579_,
		_w3580_
	);
	LUT3 #(
		.INIT('h2d)
	) name2578 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w3581_
	);
	LUT3 #(
		.INIT('h48)
	) name2579 (
		_w3571_,
		_w3580_,
		_w3581_,
		_w3582_
	);
	LUT3 #(
		.INIT('h21)
	) name2580 (
		_w3571_,
		_w3580_,
		_w3581_,
		_w3583_
	);
	LUT3 #(
		.INIT('h2d)
	) name2581 (
		_w3539_,
		_w3540_,
		_w3542_,
		_w3584_
	);
	LUT2 #(
		.INIT('h6)
	) name2582 (
		_w3546_,
		_w3584_,
		_w3585_
	);
	LUT3 #(
		.INIT('h45)
	) name2583 (
		_w3582_,
		_w3583_,
		_w3585_,
		_w3586_
	);
	LUT3 #(
		.INIT('h32)
	) name2584 (
		_w3558_,
		_w3572_,
		_w3573_,
		_w3587_
	);
	LUT4 #(
		.INIT('h0017)
	) name2585 (
		_w3550_,
		_w3575_,
		_w3586_,
		_w3587_,
		_w3588_
	);
	LUT4 #(
		.INIT('he800)
	) name2586 (
		_w3550_,
		_w3575_,
		_w3586_,
		_w3587_,
		_w3589_
	);
	LUT3 #(
		.INIT('h32)
	) name2587 (
		_w3533_,
		_w3547_,
		_w3548_,
		_w3590_
	);
	LUT3 #(
		.INIT('h54)
	) name2588 (
		_w3588_,
		_w3589_,
		_w3590_,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		\A[682] ,
		\A[683] ,
		_w3592_
	);
	LUT3 #(
		.INIT('h96)
	) name2590 (
		\A[679] ,
		\A[680] ,
		\A[681] ,
		_w3593_
	);
	LUT3 #(
		.INIT('h96)
	) name2591 (
		\A[682] ,
		\A[683] ,
		\A[684] ,
		_w3594_
	);
	LUT3 #(
		.INIT('h80)
	) name2592 (
		_w3592_,
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT3 #(
		.INIT('h17)
	) name2593 (
		\A[679] ,
		\A[680] ,
		\A[681] ,
		_w3596_
	);
	LUT3 #(
		.INIT('h17)
	) name2594 (
		\A[682] ,
		\A[683] ,
		\A[684] ,
		_w3597_
	);
	LUT4 #(
		.INIT('h080f)
	) name2595 (
		_w3593_,
		_w3594_,
		_w3596_,
		_w3597_,
		_w3598_
	);
	LUT2 #(
		.INIT('h1)
	) name2596 (
		_w3595_,
		_w3598_,
		_w3599_
	);
	LUT3 #(
		.INIT('h17)
	) name2597 (
		\A[688] ,
		\A[689] ,
		\A[690] ,
		_w3600_
	);
	LUT3 #(
		.INIT('h17)
	) name2598 (
		\A[685] ,
		\A[686] ,
		\A[687] ,
		_w3601_
	);
	LUT3 #(
		.INIT('h96)
	) name2599 (
		\A[685] ,
		\A[686] ,
		\A[687] ,
		_w3602_
	);
	LUT3 #(
		.INIT('h96)
	) name2600 (
		\A[688] ,
		\A[689] ,
		\A[690] ,
		_w3603_
	);
	LUT4 #(
		.INIT('h7111)
	) name2601 (
		_w3600_,
		_w3601_,
		_w3602_,
		_w3603_,
		_w3604_
	);
	LUT4 #(
		.INIT('h0660)
	) name2602 (
		_w3593_,
		_w3594_,
		_w3602_,
		_w3603_,
		_w3605_
	);
	LUT4 #(
		.INIT('h0080)
	) name2603 (
		_w3592_,
		_w3593_,
		_w3594_,
		_w3596_,
		_w3606_
	);
	LUT2 #(
		.INIT('h2)
	) name2604 (
		_w3605_,
		_w3606_,
		_w3607_
	);
	LUT4 #(
		.INIT('h6999)
	) name2605 (
		_w3600_,
		_w3601_,
		_w3602_,
		_w3603_,
		_w3608_
	);
	LUT3 #(
		.INIT('h02)
	) name2606 (
		_w3605_,
		_w3606_,
		_w3608_,
		_w3609_
	);
	LUT3 #(
		.INIT('hd0)
	) name2607 (
		_w3605_,
		_w3606_,
		_w3608_,
		_w3610_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2608 (
		\A[682] ,
		\A[683] ,
		\A[684] ,
		_w3593_,
		_w3611_
	);
	LUT2 #(
		.INIT('h9)
	) name2609 (
		_w3596_,
		_w3611_,
		_w3612_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2610 (
		_w3604_,
		_w3607_,
		_w3608_,
		_w3612_,
		_w3613_
	);
	LUT4 #(
		.INIT('h1051)
	) name2611 (
		_w3604_,
		_w3607_,
		_w3608_,
		_w3612_,
		_w3614_
	);
	LUT4 #(
		.INIT('h6566)
	) name2612 (
		_w3604_,
		_w3609_,
		_w3610_,
		_w3612_,
		_w3615_
	);
	LUT2 #(
		.INIT('h6)
	) name2613 (
		_w3599_,
		_w3615_,
		_w3616_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		\A[694] ,
		\A[695] ,
		_w3617_
	);
	LUT3 #(
		.INIT('h96)
	) name2615 (
		\A[691] ,
		\A[692] ,
		\A[693] ,
		_w3618_
	);
	LUT3 #(
		.INIT('h96)
	) name2616 (
		\A[694] ,
		\A[695] ,
		\A[696] ,
		_w3619_
	);
	LUT3 #(
		.INIT('h80)
	) name2617 (
		_w3617_,
		_w3618_,
		_w3619_,
		_w3620_
	);
	LUT3 #(
		.INIT('h17)
	) name2618 (
		\A[691] ,
		\A[692] ,
		\A[693] ,
		_w3621_
	);
	LUT3 #(
		.INIT('h17)
	) name2619 (
		\A[694] ,
		\A[695] ,
		\A[696] ,
		_w3622_
	);
	LUT4 #(
		.INIT('h080f)
	) name2620 (
		_w3618_,
		_w3619_,
		_w3621_,
		_w3622_,
		_w3623_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		_w3620_,
		_w3623_,
		_w3624_
	);
	LUT3 #(
		.INIT('h17)
	) name2622 (
		\A[700] ,
		\A[701] ,
		\A[702] ,
		_w3625_
	);
	LUT3 #(
		.INIT('h17)
	) name2623 (
		\A[697] ,
		\A[698] ,
		\A[699] ,
		_w3626_
	);
	LUT3 #(
		.INIT('h96)
	) name2624 (
		\A[697] ,
		\A[698] ,
		\A[699] ,
		_w3627_
	);
	LUT3 #(
		.INIT('h96)
	) name2625 (
		\A[700] ,
		\A[701] ,
		\A[702] ,
		_w3628_
	);
	LUT4 #(
		.INIT('h7111)
	) name2626 (
		_w3625_,
		_w3626_,
		_w3627_,
		_w3628_,
		_w3629_
	);
	LUT4 #(
		.INIT('h0660)
	) name2627 (
		_w3618_,
		_w3619_,
		_w3627_,
		_w3628_,
		_w3630_
	);
	LUT4 #(
		.INIT('h0080)
	) name2628 (
		_w3617_,
		_w3618_,
		_w3619_,
		_w3621_,
		_w3631_
	);
	LUT2 #(
		.INIT('h2)
	) name2629 (
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT4 #(
		.INIT('h6999)
	) name2630 (
		_w3625_,
		_w3626_,
		_w3627_,
		_w3628_,
		_w3633_
	);
	LUT3 #(
		.INIT('h02)
	) name2631 (
		_w3630_,
		_w3631_,
		_w3633_,
		_w3634_
	);
	LUT3 #(
		.INIT('hd0)
	) name2632 (
		_w3630_,
		_w3631_,
		_w3633_,
		_w3635_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2633 (
		\A[694] ,
		\A[695] ,
		\A[696] ,
		_w3618_,
		_w3636_
	);
	LUT2 #(
		.INIT('h9)
	) name2634 (
		_w3621_,
		_w3636_,
		_w3637_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2635 (
		_w3629_,
		_w3632_,
		_w3633_,
		_w3637_,
		_w3638_
	);
	LUT4 #(
		.INIT('h1051)
	) name2636 (
		_w3629_,
		_w3632_,
		_w3633_,
		_w3637_,
		_w3639_
	);
	LUT4 #(
		.INIT('h6566)
	) name2637 (
		_w3629_,
		_w3634_,
		_w3635_,
		_w3637_,
		_w3640_
	);
	LUT2 #(
		.INIT('h6)
	) name2638 (
		_w3624_,
		_w3640_,
		_w3641_
	);
	LUT4 #(
		.INIT('h9009)
	) name2639 (
		_w3599_,
		_w3615_,
		_w3624_,
		_w3640_,
		_w3642_
	);
	LUT4 #(
		.INIT('h0660)
	) name2640 (
		_w3599_,
		_w3615_,
		_w3624_,
		_w3640_,
		_w3643_
	);
	LUT4 #(
		.INIT('h6996)
	) name2641 (
		_w3618_,
		_w3619_,
		_w3627_,
		_w3628_,
		_w3644_
	);
	LUT4 #(
		.INIT('h6996)
	) name2642 (
		_w3593_,
		_w3594_,
		_w3602_,
		_w3603_,
		_w3645_
	);
	LUT2 #(
		.INIT('h8)
	) name2643 (
		_w3644_,
		_w3645_,
		_w3646_
	);
	LUT3 #(
		.INIT('h2d)
	) name2644 (
		_w3630_,
		_w3631_,
		_w3633_,
		_w3647_
	);
	LUT3 #(
		.INIT('h48)
	) name2645 (
		_w3637_,
		_w3646_,
		_w3647_,
		_w3648_
	);
	LUT3 #(
		.INIT('h21)
	) name2646 (
		_w3637_,
		_w3646_,
		_w3647_,
		_w3649_
	);
	LUT3 #(
		.INIT('h2d)
	) name2647 (
		_w3605_,
		_w3606_,
		_w3608_,
		_w3650_
	);
	LUT2 #(
		.INIT('h6)
	) name2648 (
		_w3612_,
		_w3650_,
		_w3651_
	);
	LUT3 #(
		.INIT('h45)
	) name2649 (
		_w3648_,
		_w3649_,
		_w3651_,
		_w3652_
	);
	LUT3 #(
		.INIT('h32)
	) name2650 (
		_w3624_,
		_w3638_,
		_w3639_,
		_w3653_
	);
	LUT4 #(
		.INIT('h0017)
	) name2651 (
		_w3616_,
		_w3641_,
		_w3652_,
		_w3653_,
		_w3654_
	);
	LUT4 #(
		.INIT('he800)
	) name2652 (
		_w3616_,
		_w3641_,
		_w3652_,
		_w3653_,
		_w3655_
	);
	LUT4 #(
		.INIT('hab54)
	) name2653 (
		_w3642_,
		_w3643_,
		_w3652_,
		_w3653_,
		_w3656_
	);
	LUT3 #(
		.INIT('h32)
	) name2654 (
		_w3599_,
		_w3613_,
		_w3614_,
		_w3657_
	);
	LUT2 #(
		.INIT('h9)
	) name2655 (
		_w3656_,
		_w3657_,
		_w3658_
	);
	LUT4 #(
		.INIT('hab54)
	) name2656 (
		_w3576_,
		_w3577_,
		_w3586_,
		_w3587_,
		_w3659_
	);
	LUT2 #(
		.INIT('h9)
	) name2657 (
		_w3590_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('h1428)
	) name2658 (
		_w3590_,
		_w3656_,
		_w3657_,
		_w3659_,
		_w3661_
	);
	LUT4 #(
		.INIT('h8241)
	) name2659 (
		_w3590_,
		_w3656_,
		_w3657_,
		_w3659_,
		_w3662_
	);
	LUT4 #(
		.INIT('h6996)
	) name2660 (
		_w3533_,
		_w3549_,
		_w3558_,
		_w3574_,
		_w3663_
	);
	LUT4 #(
		.INIT('h6996)
	) name2661 (
		_w3599_,
		_w3615_,
		_w3624_,
		_w3640_,
		_w3664_
	);
	LUT4 #(
		.INIT('h1248)
	) name2662 (
		_w3586_,
		_w3652_,
		_w3663_,
		_w3664_,
		_w3665_
	);
	LUT4 #(
		.INIT('h8421)
	) name2663 (
		_w3586_,
		_w3652_,
		_w3663_,
		_w3664_,
		_w3666_
	);
	LUT4 #(
		.INIT('h0660)
	) name2664 (
		_w3578_,
		_w3579_,
		_w3644_,
		_w3645_,
		_w3667_
	);
	LUT3 #(
		.INIT('h96)
	) name2665 (
		_w3637_,
		_w3646_,
		_w3647_,
		_w3668_
	);
	LUT3 #(
		.INIT('h48)
	) name2666 (
		_w3651_,
		_w3667_,
		_w3668_,
		_w3669_
	);
	LUT3 #(
		.INIT('h21)
	) name2667 (
		_w3651_,
		_w3667_,
		_w3668_,
		_w3670_
	);
	LUT3 #(
		.INIT('h96)
	) name2668 (
		_w3571_,
		_w3580_,
		_w3581_,
		_w3671_
	);
	LUT2 #(
		.INIT('h9)
	) name2669 (
		_w3585_,
		_w3671_,
		_w3672_
	);
	LUT3 #(
		.INIT('h54)
	) name2670 (
		_w3669_,
		_w3670_,
		_w3672_,
		_w3673_
	);
	LUT3 #(
		.INIT('h45)
	) name2671 (
		_w3665_,
		_w3666_,
		_w3673_,
		_w3674_
	);
	LUT3 #(
		.INIT('h54)
	) name2672 (
		_w3661_,
		_w3662_,
		_w3674_,
		_w3675_
	);
	LUT4 #(
		.INIT('h022a)
	) name2673 (
		_w3591_,
		_w3658_,
		_w3660_,
		_w3674_,
		_w3676_
	);
	LUT4 #(
		.INIT('h5440)
	) name2674 (
		_w3591_,
		_w3658_,
		_w3660_,
		_w3674_,
		_w3677_
	);
	LUT3 #(
		.INIT('h54)
	) name2675 (
		_w3654_,
		_w3655_,
		_w3657_,
		_w3678_
	);
	LUT4 #(
		.INIT('h1051)
	) name2676 (
		_w3525_,
		_w3591_,
		_w3675_,
		_w3678_,
		_w3679_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2677 (
		_w3525_,
		_w3591_,
		_w3675_,
		_w3678_,
		_w3680_
	);
	LUT4 #(
		.INIT('h6665)
	) name2678 (
		_w3591_,
		_w3661_,
		_w3662_,
		_w3674_,
		_w3681_
	);
	LUT3 #(
		.INIT('h96)
	) name2679 (
		_w3521_,
		_w3523_,
		_w3524_,
		_w3682_
	);
	LUT3 #(
		.INIT('h96)
	) name2680 (
		_w3461_,
		_w3513_,
		_w3520_,
		_w3683_
	);
	LUT4 #(
		.INIT('h6996)
	) name2681 (
		_w3590_,
		_w3656_,
		_w3657_,
		_w3659_,
		_w3684_
	);
	LUT4 #(
		.INIT('h6996)
	) name2682 (
		_w3586_,
		_w3652_,
		_w3663_,
		_w3664_,
		_w3685_
	);
	LUT4 #(
		.INIT('h6996)
	) name2683 (
		_w3460_,
		_w3514_,
		_w3515_,
		_w3519_,
		_w3686_
	);
	LUT4 #(
		.INIT('h6996)
	) name2684 (
		_w3452_,
		_w3453_,
		_w3506_,
		_w3507_,
		_w3687_
	);
	LUT4 #(
		.INIT('h6996)
	) name2685 (
		_w3578_,
		_w3579_,
		_w3644_,
		_w3645_,
		_w3688_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		_w3687_,
		_w3688_,
		_w3689_
	);
	LUT4 #(
		.INIT('h6996)
	) name2687 (
		_w3459_,
		_w3516_,
		_w3517_,
		_w3518_,
		_w3690_
	);
	LUT3 #(
		.INIT('h96)
	) name2688 (
		_w3651_,
		_w3667_,
		_w3668_,
		_w3691_
	);
	LUT4 #(
		.INIT('h71b2)
	) name2689 (
		_w3672_,
		_w3689_,
		_w3690_,
		_w3691_,
		_w3692_
	);
	LUT4 #(
		.INIT('h90f9)
	) name2690 (
		_w3673_,
		_w3685_,
		_w3686_,
		_w3692_,
		_w3693_
	);
	LUT4 #(
		.INIT('h84ed)
	) name2691 (
		_w3674_,
		_w3683_,
		_w3684_,
		_w3693_,
		_w3694_
	);
	LUT4 #(
		.INIT('h6f06)
	) name2692 (
		_w3678_,
		_w3681_,
		_w3682_,
		_w3694_,
		_w3695_
	);
	LUT3 #(
		.INIT('h54)
	) name2693 (
		_w3679_,
		_w3680_,
		_w3695_,
		_w3696_
	);
	LUT2 #(
		.INIT('h1)
	) name2694 (
		_w3398_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		_w3398_,
		_w3696_,
		_w3698_
	);
	LUT2 #(
		.INIT('h6)
	) name2696 (
		_w3253_,
		_w3379_,
		_w3699_
	);
	LUT4 #(
		.INIT('h6566)
	) name2697 (
		_w3525_,
		_w3676_,
		_w3677_,
		_w3678_,
		_w3700_
	);
	LUT4 #(
		.INIT('h1248)
	) name2698 (
		_w3397_,
		_w3695_,
		_w3699_,
		_w3700_,
		_w3701_
	);
	LUT4 #(
		.INIT('h8421)
	) name2699 (
		_w3397_,
		_w3695_,
		_w3699_,
		_w3700_,
		_w3702_
	);
	LUT3 #(
		.INIT('h96)
	) name2700 (
		_w3383_,
		_w3384_,
		_w3396_,
		_w3703_
	);
	LUT4 #(
		.INIT('h6996)
	) name2701 (
		_w3678_,
		_w3681_,
		_w3682_,
		_w3694_,
		_w3704_
	);
	LUT3 #(
		.INIT('h96)
	) name2702 (
		_w3385_,
		_w3386_,
		_w3395_,
		_w3705_
	);
	LUT4 #(
		.INIT('h9669)
	) name2703 (
		_w3674_,
		_w3683_,
		_w3684_,
		_w3693_,
		_w3706_
	);
	LUT4 #(
		.INIT('h6996)
	) name2704 (
		_w3673_,
		_w3685_,
		_w3686_,
		_w3692_,
		_w3707_
	);
	LUT3 #(
		.INIT('h69)
	) name2705 (
		_w3387_,
		_w3388_,
		_w3394_,
		_w3708_
	);
	LUT4 #(
		.INIT('h0660)
	) name2706 (
		_w3389_,
		_w3390_,
		_w3687_,
		_w3688_,
		_w3709_
	);
	LUT4 #(
		.INIT('h9600)
	) name2707 (
		_w3391_,
		_w3392_,
		_w3393_,
		_w3709_,
		_w3710_
	);
	LUT4 #(
		.INIT('h0069)
	) name2708 (
		_w3391_,
		_w3392_,
		_w3393_,
		_w3709_,
		_w3711_
	);
	LUT4 #(
		.INIT('h9669)
	) name2709 (
		_w3672_,
		_w3689_,
		_w3690_,
		_w3691_,
		_w3712_
	);
	LUT3 #(
		.INIT('h54)
	) name2710 (
		_w3710_,
		_w3711_,
		_w3712_,
		_w3713_
	);
	LUT3 #(
		.INIT('h8e)
	) name2711 (
		_w3707_,
		_w3708_,
		_w3713_,
		_w3714_
	);
	LUT3 #(
		.INIT('hd4)
	) name2712 (
		_w3705_,
		_w3706_,
		_w3714_,
		_w3715_
	);
	LUT3 #(
		.INIT('hd4)
	) name2713 (
		_w3703_,
		_w3704_,
		_w3715_,
		_w3716_
	);
	LUT3 #(
		.INIT('h54)
	) name2714 (
		_w3701_,
		_w3702_,
		_w3716_,
		_w3717_
	);
	LUT3 #(
		.INIT('h45)
	) name2715 (
		_w3697_,
		_w3698_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h8)
	) name2716 (
		\A[562] ,
		\A[563] ,
		_w3719_
	);
	LUT3 #(
		.INIT('h96)
	) name2717 (
		\A[559] ,
		\A[560] ,
		\A[561] ,
		_w3720_
	);
	LUT3 #(
		.INIT('h96)
	) name2718 (
		\A[562] ,
		\A[563] ,
		\A[564] ,
		_w3721_
	);
	LUT3 #(
		.INIT('h80)
	) name2719 (
		_w3719_,
		_w3720_,
		_w3721_,
		_w3722_
	);
	LUT3 #(
		.INIT('h17)
	) name2720 (
		\A[559] ,
		\A[560] ,
		\A[561] ,
		_w3723_
	);
	LUT3 #(
		.INIT('h17)
	) name2721 (
		\A[562] ,
		\A[563] ,
		\A[564] ,
		_w3724_
	);
	LUT4 #(
		.INIT('h080f)
	) name2722 (
		_w3720_,
		_w3721_,
		_w3723_,
		_w3724_,
		_w3725_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w3722_,
		_w3725_,
		_w3726_
	);
	LUT3 #(
		.INIT('h17)
	) name2724 (
		\A[568] ,
		\A[569] ,
		\A[570] ,
		_w3727_
	);
	LUT3 #(
		.INIT('h17)
	) name2725 (
		\A[565] ,
		\A[566] ,
		\A[567] ,
		_w3728_
	);
	LUT3 #(
		.INIT('h96)
	) name2726 (
		\A[565] ,
		\A[566] ,
		\A[567] ,
		_w3729_
	);
	LUT3 #(
		.INIT('h96)
	) name2727 (
		\A[568] ,
		\A[569] ,
		\A[570] ,
		_w3730_
	);
	LUT4 #(
		.INIT('h7111)
	) name2728 (
		_w3727_,
		_w3728_,
		_w3729_,
		_w3730_,
		_w3731_
	);
	LUT4 #(
		.INIT('h0660)
	) name2729 (
		_w3720_,
		_w3721_,
		_w3729_,
		_w3730_,
		_w3732_
	);
	LUT4 #(
		.INIT('h0080)
	) name2730 (
		_w3719_,
		_w3720_,
		_w3721_,
		_w3723_,
		_w3733_
	);
	LUT2 #(
		.INIT('h2)
	) name2731 (
		_w3732_,
		_w3733_,
		_w3734_
	);
	LUT4 #(
		.INIT('h6999)
	) name2732 (
		_w3727_,
		_w3728_,
		_w3729_,
		_w3730_,
		_w3735_
	);
	LUT3 #(
		.INIT('h02)
	) name2733 (
		_w3732_,
		_w3733_,
		_w3735_,
		_w3736_
	);
	LUT3 #(
		.INIT('hd0)
	) name2734 (
		_w3732_,
		_w3733_,
		_w3735_,
		_w3737_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2735 (
		\A[562] ,
		\A[563] ,
		\A[564] ,
		_w3720_,
		_w3738_
	);
	LUT2 #(
		.INIT('h9)
	) name2736 (
		_w3723_,
		_w3738_,
		_w3739_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2737 (
		_w3731_,
		_w3734_,
		_w3735_,
		_w3739_,
		_w3740_
	);
	LUT4 #(
		.INIT('h1051)
	) name2738 (
		_w3731_,
		_w3734_,
		_w3735_,
		_w3739_,
		_w3741_
	);
	LUT4 #(
		.INIT('h6566)
	) name2739 (
		_w3731_,
		_w3736_,
		_w3737_,
		_w3739_,
		_w3742_
	);
	LUT2 #(
		.INIT('h6)
	) name2740 (
		_w3726_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h8)
	) name2741 (
		\A[574] ,
		\A[575] ,
		_w3744_
	);
	LUT3 #(
		.INIT('h96)
	) name2742 (
		\A[571] ,
		\A[572] ,
		\A[573] ,
		_w3745_
	);
	LUT3 #(
		.INIT('h96)
	) name2743 (
		\A[574] ,
		\A[575] ,
		\A[576] ,
		_w3746_
	);
	LUT3 #(
		.INIT('h80)
	) name2744 (
		_w3744_,
		_w3745_,
		_w3746_,
		_w3747_
	);
	LUT3 #(
		.INIT('h17)
	) name2745 (
		\A[571] ,
		\A[572] ,
		\A[573] ,
		_w3748_
	);
	LUT3 #(
		.INIT('h17)
	) name2746 (
		\A[574] ,
		\A[575] ,
		\A[576] ,
		_w3749_
	);
	LUT4 #(
		.INIT('h080f)
	) name2747 (
		_w3745_,
		_w3746_,
		_w3748_,
		_w3749_,
		_w3750_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w3747_,
		_w3750_,
		_w3751_
	);
	LUT3 #(
		.INIT('h17)
	) name2749 (
		\A[580] ,
		\A[581] ,
		\A[582] ,
		_w3752_
	);
	LUT3 #(
		.INIT('h17)
	) name2750 (
		\A[577] ,
		\A[578] ,
		\A[579] ,
		_w3753_
	);
	LUT3 #(
		.INIT('h96)
	) name2751 (
		\A[577] ,
		\A[578] ,
		\A[579] ,
		_w3754_
	);
	LUT3 #(
		.INIT('h96)
	) name2752 (
		\A[580] ,
		\A[581] ,
		\A[582] ,
		_w3755_
	);
	LUT4 #(
		.INIT('h7111)
	) name2753 (
		_w3752_,
		_w3753_,
		_w3754_,
		_w3755_,
		_w3756_
	);
	LUT4 #(
		.INIT('h0660)
	) name2754 (
		_w3745_,
		_w3746_,
		_w3754_,
		_w3755_,
		_w3757_
	);
	LUT4 #(
		.INIT('h0080)
	) name2755 (
		_w3744_,
		_w3745_,
		_w3746_,
		_w3748_,
		_w3758_
	);
	LUT2 #(
		.INIT('h2)
	) name2756 (
		_w3757_,
		_w3758_,
		_w3759_
	);
	LUT4 #(
		.INIT('h6999)
	) name2757 (
		_w3752_,
		_w3753_,
		_w3754_,
		_w3755_,
		_w3760_
	);
	LUT3 #(
		.INIT('h02)
	) name2758 (
		_w3757_,
		_w3758_,
		_w3760_,
		_w3761_
	);
	LUT3 #(
		.INIT('hd0)
	) name2759 (
		_w3757_,
		_w3758_,
		_w3760_,
		_w3762_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2760 (
		\A[574] ,
		\A[575] ,
		\A[576] ,
		_w3745_,
		_w3763_
	);
	LUT2 #(
		.INIT('h9)
	) name2761 (
		_w3748_,
		_w3763_,
		_w3764_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2762 (
		_w3756_,
		_w3759_,
		_w3760_,
		_w3764_,
		_w3765_
	);
	LUT4 #(
		.INIT('h1051)
	) name2763 (
		_w3756_,
		_w3759_,
		_w3760_,
		_w3764_,
		_w3766_
	);
	LUT4 #(
		.INIT('h6566)
	) name2764 (
		_w3756_,
		_w3761_,
		_w3762_,
		_w3764_,
		_w3767_
	);
	LUT2 #(
		.INIT('h6)
	) name2765 (
		_w3751_,
		_w3767_,
		_w3768_
	);
	LUT4 #(
		.INIT('h9009)
	) name2766 (
		_w3726_,
		_w3742_,
		_w3751_,
		_w3767_,
		_w3769_
	);
	LUT4 #(
		.INIT('h0660)
	) name2767 (
		_w3726_,
		_w3742_,
		_w3751_,
		_w3767_,
		_w3770_
	);
	LUT4 #(
		.INIT('h6996)
	) name2768 (
		_w3745_,
		_w3746_,
		_w3754_,
		_w3755_,
		_w3771_
	);
	LUT4 #(
		.INIT('h6996)
	) name2769 (
		_w3720_,
		_w3721_,
		_w3729_,
		_w3730_,
		_w3772_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		_w3771_,
		_w3772_,
		_w3773_
	);
	LUT3 #(
		.INIT('h2d)
	) name2771 (
		_w3757_,
		_w3758_,
		_w3760_,
		_w3774_
	);
	LUT3 #(
		.INIT('h48)
	) name2772 (
		_w3764_,
		_w3773_,
		_w3774_,
		_w3775_
	);
	LUT3 #(
		.INIT('h21)
	) name2773 (
		_w3764_,
		_w3773_,
		_w3774_,
		_w3776_
	);
	LUT3 #(
		.INIT('h2d)
	) name2774 (
		_w3732_,
		_w3733_,
		_w3735_,
		_w3777_
	);
	LUT2 #(
		.INIT('h6)
	) name2775 (
		_w3739_,
		_w3777_,
		_w3778_
	);
	LUT3 #(
		.INIT('h45)
	) name2776 (
		_w3775_,
		_w3776_,
		_w3778_,
		_w3779_
	);
	LUT3 #(
		.INIT('h32)
	) name2777 (
		_w3751_,
		_w3765_,
		_w3766_,
		_w3780_
	);
	LUT4 #(
		.INIT('h0017)
	) name2778 (
		_w3743_,
		_w3768_,
		_w3779_,
		_w3780_,
		_w3781_
	);
	LUT4 #(
		.INIT('he800)
	) name2779 (
		_w3743_,
		_w3768_,
		_w3779_,
		_w3780_,
		_w3782_
	);
	LUT3 #(
		.INIT('h32)
	) name2780 (
		_w3726_,
		_w3740_,
		_w3741_,
		_w3783_
	);
	LUT3 #(
		.INIT('h54)
	) name2781 (
		_w3781_,
		_w3782_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h8)
	) name2782 (
		\A[586] ,
		\A[587] ,
		_w3785_
	);
	LUT3 #(
		.INIT('h96)
	) name2783 (
		\A[583] ,
		\A[584] ,
		\A[585] ,
		_w3786_
	);
	LUT3 #(
		.INIT('h96)
	) name2784 (
		\A[586] ,
		\A[587] ,
		\A[588] ,
		_w3787_
	);
	LUT3 #(
		.INIT('h80)
	) name2785 (
		_w3785_,
		_w3786_,
		_w3787_,
		_w3788_
	);
	LUT3 #(
		.INIT('h17)
	) name2786 (
		\A[583] ,
		\A[584] ,
		\A[585] ,
		_w3789_
	);
	LUT3 #(
		.INIT('h17)
	) name2787 (
		\A[586] ,
		\A[587] ,
		\A[588] ,
		_w3790_
	);
	LUT4 #(
		.INIT('h080f)
	) name2788 (
		_w3786_,
		_w3787_,
		_w3789_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h1)
	) name2789 (
		_w3788_,
		_w3791_,
		_w3792_
	);
	LUT3 #(
		.INIT('h17)
	) name2790 (
		\A[592] ,
		\A[593] ,
		\A[594] ,
		_w3793_
	);
	LUT3 #(
		.INIT('h17)
	) name2791 (
		\A[589] ,
		\A[590] ,
		\A[591] ,
		_w3794_
	);
	LUT3 #(
		.INIT('h96)
	) name2792 (
		\A[589] ,
		\A[590] ,
		\A[591] ,
		_w3795_
	);
	LUT3 #(
		.INIT('h96)
	) name2793 (
		\A[592] ,
		\A[593] ,
		\A[594] ,
		_w3796_
	);
	LUT4 #(
		.INIT('h7111)
	) name2794 (
		_w3793_,
		_w3794_,
		_w3795_,
		_w3796_,
		_w3797_
	);
	LUT4 #(
		.INIT('h0660)
	) name2795 (
		_w3786_,
		_w3787_,
		_w3795_,
		_w3796_,
		_w3798_
	);
	LUT4 #(
		.INIT('h0080)
	) name2796 (
		_w3785_,
		_w3786_,
		_w3787_,
		_w3789_,
		_w3799_
	);
	LUT2 #(
		.INIT('h2)
	) name2797 (
		_w3798_,
		_w3799_,
		_w3800_
	);
	LUT4 #(
		.INIT('h6999)
	) name2798 (
		_w3793_,
		_w3794_,
		_w3795_,
		_w3796_,
		_w3801_
	);
	LUT3 #(
		.INIT('h02)
	) name2799 (
		_w3798_,
		_w3799_,
		_w3801_,
		_w3802_
	);
	LUT3 #(
		.INIT('hd0)
	) name2800 (
		_w3798_,
		_w3799_,
		_w3801_,
		_w3803_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2801 (
		\A[586] ,
		\A[587] ,
		\A[588] ,
		_w3786_,
		_w3804_
	);
	LUT2 #(
		.INIT('h9)
	) name2802 (
		_w3789_,
		_w3804_,
		_w3805_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2803 (
		_w3797_,
		_w3800_,
		_w3801_,
		_w3805_,
		_w3806_
	);
	LUT4 #(
		.INIT('h1051)
	) name2804 (
		_w3797_,
		_w3800_,
		_w3801_,
		_w3805_,
		_w3807_
	);
	LUT4 #(
		.INIT('h6566)
	) name2805 (
		_w3797_,
		_w3802_,
		_w3803_,
		_w3805_,
		_w3808_
	);
	LUT2 #(
		.INIT('h6)
	) name2806 (
		_w3792_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name2807 (
		\A[598] ,
		\A[599] ,
		_w3810_
	);
	LUT3 #(
		.INIT('h96)
	) name2808 (
		\A[595] ,
		\A[596] ,
		\A[597] ,
		_w3811_
	);
	LUT3 #(
		.INIT('h96)
	) name2809 (
		\A[598] ,
		\A[599] ,
		\A[600] ,
		_w3812_
	);
	LUT3 #(
		.INIT('h80)
	) name2810 (
		_w3810_,
		_w3811_,
		_w3812_,
		_w3813_
	);
	LUT3 #(
		.INIT('h17)
	) name2811 (
		\A[595] ,
		\A[596] ,
		\A[597] ,
		_w3814_
	);
	LUT3 #(
		.INIT('h17)
	) name2812 (
		\A[598] ,
		\A[599] ,
		\A[600] ,
		_w3815_
	);
	LUT4 #(
		.INIT('h080f)
	) name2813 (
		_w3811_,
		_w3812_,
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		_w3813_,
		_w3816_,
		_w3817_
	);
	LUT3 #(
		.INIT('h17)
	) name2815 (
		\A[604] ,
		\A[605] ,
		\A[606] ,
		_w3818_
	);
	LUT3 #(
		.INIT('h17)
	) name2816 (
		\A[601] ,
		\A[602] ,
		\A[603] ,
		_w3819_
	);
	LUT3 #(
		.INIT('h96)
	) name2817 (
		\A[601] ,
		\A[602] ,
		\A[603] ,
		_w3820_
	);
	LUT3 #(
		.INIT('h96)
	) name2818 (
		\A[604] ,
		\A[605] ,
		\A[606] ,
		_w3821_
	);
	LUT4 #(
		.INIT('h7111)
	) name2819 (
		_w3818_,
		_w3819_,
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('h0660)
	) name2820 (
		_w3811_,
		_w3812_,
		_w3820_,
		_w3821_,
		_w3823_
	);
	LUT4 #(
		.INIT('h0080)
	) name2821 (
		_w3810_,
		_w3811_,
		_w3812_,
		_w3814_,
		_w3824_
	);
	LUT2 #(
		.INIT('h2)
	) name2822 (
		_w3823_,
		_w3824_,
		_w3825_
	);
	LUT4 #(
		.INIT('h6999)
	) name2823 (
		_w3818_,
		_w3819_,
		_w3820_,
		_w3821_,
		_w3826_
	);
	LUT3 #(
		.INIT('h02)
	) name2824 (
		_w3823_,
		_w3824_,
		_w3826_,
		_w3827_
	);
	LUT3 #(
		.INIT('hd0)
	) name2825 (
		_w3823_,
		_w3824_,
		_w3826_,
		_w3828_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2826 (
		\A[598] ,
		\A[599] ,
		\A[600] ,
		_w3811_,
		_w3829_
	);
	LUT2 #(
		.INIT('h9)
	) name2827 (
		_w3814_,
		_w3829_,
		_w3830_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2828 (
		_w3822_,
		_w3825_,
		_w3826_,
		_w3830_,
		_w3831_
	);
	LUT4 #(
		.INIT('h1051)
	) name2829 (
		_w3822_,
		_w3825_,
		_w3826_,
		_w3830_,
		_w3832_
	);
	LUT4 #(
		.INIT('h6566)
	) name2830 (
		_w3822_,
		_w3827_,
		_w3828_,
		_w3830_,
		_w3833_
	);
	LUT2 #(
		.INIT('h6)
	) name2831 (
		_w3817_,
		_w3833_,
		_w3834_
	);
	LUT4 #(
		.INIT('h9009)
	) name2832 (
		_w3792_,
		_w3808_,
		_w3817_,
		_w3833_,
		_w3835_
	);
	LUT4 #(
		.INIT('h0660)
	) name2833 (
		_w3792_,
		_w3808_,
		_w3817_,
		_w3833_,
		_w3836_
	);
	LUT4 #(
		.INIT('h6996)
	) name2834 (
		_w3811_,
		_w3812_,
		_w3820_,
		_w3821_,
		_w3837_
	);
	LUT4 #(
		.INIT('h6996)
	) name2835 (
		_w3786_,
		_w3787_,
		_w3795_,
		_w3796_,
		_w3838_
	);
	LUT2 #(
		.INIT('h8)
	) name2836 (
		_w3837_,
		_w3838_,
		_w3839_
	);
	LUT3 #(
		.INIT('h2d)
	) name2837 (
		_w3823_,
		_w3824_,
		_w3826_,
		_w3840_
	);
	LUT3 #(
		.INIT('h48)
	) name2838 (
		_w3830_,
		_w3839_,
		_w3840_,
		_w3841_
	);
	LUT3 #(
		.INIT('h21)
	) name2839 (
		_w3830_,
		_w3839_,
		_w3840_,
		_w3842_
	);
	LUT3 #(
		.INIT('h2d)
	) name2840 (
		_w3798_,
		_w3799_,
		_w3801_,
		_w3843_
	);
	LUT2 #(
		.INIT('h6)
	) name2841 (
		_w3805_,
		_w3843_,
		_w3844_
	);
	LUT3 #(
		.INIT('h45)
	) name2842 (
		_w3841_,
		_w3842_,
		_w3844_,
		_w3845_
	);
	LUT3 #(
		.INIT('h32)
	) name2843 (
		_w3817_,
		_w3831_,
		_w3832_,
		_w3846_
	);
	LUT4 #(
		.INIT('h0017)
	) name2844 (
		_w3809_,
		_w3834_,
		_w3845_,
		_w3846_,
		_w3847_
	);
	LUT4 #(
		.INIT('he800)
	) name2845 (
		_w3809_,
		_w3834_,
		_w3845_,
		_w3846_,
		_w3848_
	);
	LUT4 #(
		.INIT('hab54)
	) name2846 (
		_w3835_,
		_w3836_,
		_w3845_,
		_w3846_,
		_w3849_
	);
	LUT3 #(
		.INIT('h32)
	) name2847 (
		_w3792_,
		_w3806_,
		_w3807_,
		_w3850_
	);
	LUT2 #(
		.INIT('h9)
	) name2848 (
		_w3849_,
		_w3850_,
		_w3851_
	);
	LUT4 #(
		.INIT('hab54)
	) name2849 (
		_w3769_,
		_w3770_,
		_w3779_,
		_w3780_,
		_w3852_
	);
	LUT2 #(
		.INIT('h9)
	) name2850 (
		_w3783_,
		_w3852_,
		_w3853_
	);
	LUT4 #(
		.INIT('h1428)
	) name2851 (
		_w3783_,
		_w3849_,
		_w3850_,
		_w3852_,
		_w3854_
	);
	LUT4 #(
		.INIT('h8241)
	) name2852 (
		_w3783_,
		_w3849_,
		_w3850_,
		_w3852_,
		_w3855_
	);
	LUT4 #(
		.INIT('h6996)
	) name2853 (
		_w3726_,
		_w3742_,
		_w3751_,
		_w3767_,
		_w3856_
	);
	LUT4 #(
		.INIT('h6996)
	) name2854 (
		_w3792_,
		_w3808_,
		_w3817_,
		_w3833_,
		_w3857_
	);
	LUT4 #(
		.INIT('h1248)
	) name2855 (
		_w3779_,
		_w3845_,
		_w3856_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('h8421)
	) name2856 (
		_w3779_,
		_w3845_,
		_w3856_,
		_w3857_,
		_w3859_
	);
	LUT4 #(
		.INIT('h0660)
	) name2857 (
		_w3771_,
		_w3772_,
		_w3837_,
		_w3838_,
		_w3860_
	);
	LUT3 #(
		.INIT('h96)
	) name2858 (
		_w3830_,
		_w3839_,
		_w3840_,
		_w3861_
	);
	LUT3 #(
		.INIT('h48)
	) name2859 (
		_w3844_,
		_w3860_,
		_w3861_,
		_w3862_
	);
	LUT3 #(
		.INIT('h21)
	) name2860 (
		_w3844_,
		_w3860_,
		_w3861_,
		_w3863_
	);
	LUT3 #(
		.INIT('h96)
	) name2861 (
		_w3764_,
		_w3773_,
		_w3774_,
		_w3864_
	);
	LUT2 #(
		.INIT('h9)
	) name2862 (
		_w3778_,
		_w3864_,
		_w3865_
	);
	LUT3 #(
		.INIT('h54)
	) name2863 (
		_w3862_,
		_w3863_,
		_w3865_,
		_w3866_
	);
	LUT3 #(
		.INIT('h45)
	) name2864 (
		_w3858_,
		_w3859_,
		_w3866_,
		_w3867_
	);
	LUT4 #(
		.INIT('h022a)
	) name2865 (
		_w3784_,
		_w3851_,
		_w3853_,
		_w3867_,
		_w3868_
	);
	LUT4 #(
		.INIT('h5440)
	) name2866 (
		_w3784_,
		_w3851_,
		_w3853_,
		_w3867_,
		_w3869_
	);
	LUT4 #(
		.INIT('h6665)
	) name2867 (
		_w3784_,
		_w3854_,
		_w3855_,
		_w3867_,
		_w3870_
	);
	LUT3 #(
		.INIT('h54)
	) name2868 (
		_w3847_,
		_w3848_,
		_w3850_,
		_w3871_
	);
	LUT2 #(
		.INIT('h6)
	) name2869 (
		_w3870_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		\A[634] ,
		\A[635] ,
		_w3873_
	);
	LUT3 #(
		.INIT('h96)
	) name2871 (
		\A[631] ,
		\A[632] ,
		\A[633] ,
		_w3874_
	);
	LUT3 #(
		.INIT('h96)
	) name2872 (
		\A[634] ,
		\A[635] ,
		\A[636] ,
		_w3875_
	);
	LUT3 #(
		.INIT('h80)
	) name2873 (
		_w3873_,
		_w3874_,
		_w3875_,
		_w3876_
	);
	LUT3 #(
		.INIT('h17)
	) name2874 (
		\A[631] ,
		\A[632] ,
		\A[633] ,
		_w3877_
	);
	LUT3 #(
		.INIT('h17)
	) name2875 (
		\A[634] ,
		\A[635] ,
		\A[636] ,
		_w3878_
	);
	LUT4 #(
		.INIT('h080f)
	) name2876 (
		_w3874_,
		_w3875_,
		_w3877_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w3876_,
		_w3879_,
		_w3880_
	);
	LUT3 #(
		.INIT('h17)
	) name2878 (
		\A[640] ,
		\A[641] ,
		\A[642] ,
		_w3881_
	);
	LUT3 #(
		.INIT('h17)
	) name2879 (
		\A[637] ,
		\A[638] ,
		\A[639] ,
		_w3882_
	);
	LUT3 #(
		.INIT('h96)
	) name2880 (
		\A[637] ,
		\A[638] ,
		\A[639] ,
		_w3883_
	);
	LUT3 #(
		.INIT('h96)
	) name2881 (
		\A[640] ,
		\A[641] ,
		\A[642] ,
		_w3884_
	);
	LUT4 #(
		.INIT('h7111)
	) name2882 (
		_w3881_,
		_w3882_,
		_w3883_,
		_w3884_,
		_w3885_
	);
	LUT4 #(
		.INIT('h0660)
	) name2883 (
		_w3874_,
		_w3875_,
		_w3883_,
		_w3884_,
		_w3886_
	);
	LUT4 #(
		.INIT('h0080)
	) name2884 (
		_w3873_,
		_w3874_,
		_w3875_,
		_w3877_,
		_w3887_
	);
	LUT2 #(
		.INIT('h2)
	) name2885 (
		_w3886_,
		_w3887_,
		_w3888_
	);
	LUT4 #(
		.INIT('h6999)
	) name2886 (
		_w3881_,
		_w3882_,
		_w3883_,
		_w3884_,
		_w3889_
	);
	LUT3 #(
		.INIT('h02)
	) name2887 (
		_w3886_,
		_w3887_,
		_w3889_,
		_w3890_
	);
	LUT3 #(
		.INIT('hd0)
	) name2888 (
		_w3886_,
		_w3887_,
		_w3889_,
		_w3891_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2889 (
		\A[634] ,
		\A[635] ,
		\A[636] ,
		_w3874_,
		_w3892_
	);
	LUT2 #(
		.INIT('h9)
	) name2890 (
		_w3877_,
		_w3892_,
		_w3893_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2891 (
		_w3885_,
		_w3888_,
		_w3889_,
		_w3893_,
		_w3894_
	);
	LUT4 #(
		.INIT('h1051)
	) name2892 (
		_w3885_,
		_w3888_,
		_w3889_,
		_w3893_,
		_w3895_
	);
	LUT4 #(
		.INIT('h6566)
	) name2893 (
		_w3885_,
		_w3890_,
		_w3891_,
		_w3893_,
		_w3896_
	);
	LUT2 #(
		.INIT('h6)
	) name2894 (
		_w3880_,
		_w3896_,
		_w3897_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		\A[646] ,
		\A[647] ,
		_w3898_
	);
	LUT3 #(
		.INIT('h96)
	) name2896 (
		\A[643] ,
		\A[644] ,
		\A[645] ,
		_w3899_
	);
	LUT3 #(
		.INIT('h96)
	) name2897 (
		\A[646] ,
		\A[647] ,
		\A[648] ,
		_w3900_
	);
	LUT3 #(
		.INIT('h80)
	) name2898 (
		_w3898_,
		_w3899_,
		_w3900_,
		_w3901_
	);
	LUT3 #(
		.INIT('h17)
	) name2899 (
		\A[643] ,
		\A[644] ,
		\A[645] ,
		_w3902_
	);
	LUT3 #(
		.INIT('h17)
	) name2900 (
		\A[646] ,
		\A[647] ,
		\A[648] ,
		_w3903_
	);
	LUT4 #(
		.INIT('h080f)
	) name2901 (
		_w3899_,
		_w3900_,
		_w3902_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h1)
	) name2902 (
		_w3901_,
		_w3904_,
		_w3905_
	);
	LUT3 #(
		.INIT('h17)
	) name2903 (
		\A[652] ,
		\A[653] ,
		\A[654] ,
		_w3906_
	);
	LUT3 #(
		.INIT('h17)
	) name2904 (
		\A[649] ,
		\A[650] ,
		\A[651] ,
		_w3907_
	);
	LUT3 #(
		.INIT('h96)
	) name2905 (
		\A[649] ,
		\A[650] ,
		\A[651] ,
		_w3908_
	);
	LUT3 #(
		.INIT('h96)
	) name2906 (
		\A[652] ,
		\A[653] ,
		\A[654] ,
		_w3909_
	);
	LUT4 #(
		.INIT('h7111)
	) name2907 (
		_w3906_,
		_w3907_,
		_w3908_,
		_w3909_,
		_w3910_
	);
	LUT4 #(
		.INIT('h0660)
	) name2908 (
		_w3899_,
		_w3900_,
		_w3908_,
		_w3909_,
		_w3911_
	);
	LUT4 #(
		.INIT('h0080)
	) name2909 (
		_w3898_,
		_w3899_,
		_w3900_,
		_w3902_,
		_w3912_
	);
	LUT2 #(
		.INIT('h2)
	) name2910 (
		_w3911_,
		_w3912_,
		_w3913_
	);
	LUT4 #(
		.INIT('h6999)
	) name2911 (
		_w3906_,
		_w3907_,
		_w3908_,
		_w3909_,
		_w3914_
	);
	LUT3 #(
		.INIT('h02)
	) name2912 (
		_w3911_,
		_w3912_,
		_w3914_,
		_w3915_
	);
	LUT3 #(
		.INIT('hd0)
	) name2913 (
		_w3911_,
		_w3912_,
		_w3914_,
		_w3916_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2914 (
		\A[646] ,
		\A[647] ,
		\A[648] ,
		_w3899_,
		_w3917_
	);
	LUT2 #(
		.INIT('h9)
	) name2915 (
		_w3902_,
		_w3917_,
		_w3918_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2916 (
		_w3910_,
		_w3913_,
		_w3914_,
		_w3918_,
		_w3919_
	);
	LUT4 #(
		.INIT('h1051)
	) name2917 (
		_w3910_,
		_w3913_,
		_w3914_,
		_w3918_,
		_w3920_
	);
	LUT4 #(
		.INIT('h6566)
	) name2918 (
		_w3910_,
		_w3915_,
		_w3916_,
		_w3918_,
		_w3921_
	);
	LUT2 #(
		.INIT('h6)
	) name2919 (
		_w3905_,
		_w3921_,
		_w3922_
	);
	LUT4 #(
		.INIT('h9009)
	) name2920 (
		_w3880_,
		_w3896_,
		_w3905_,
		_w3921_,
		_w3923_
	);
	LUT4 #(
		.INIT('h0660)
	) name2921 (
		_w3880_,
		_w3896_,
		_w3905_,
		_w3921_,
		_w3924_
	);
	LUT4 #(
		.INIT('h6996)
	) name2922 (
		_w3899_,
		_w3900_,
		_w3908_,
		_w3909_,
		_w3925_
	);
	LUT4 #(
		.INIT('h6996)
	) name2923 (
		_w3874_,
		_w3875_,
		_w3883_,
		_w3884_,
		_w3926_
	);
	LUT2 #(
		.INIT('h8)
	) name2924 (
		_w3925_,
		_w3926_,
		_w3927_
	);
	LUT3 #(
		.INIT('h2d)
	) name2925 (
		_w3911_,
		_w3912_,
		_w3914_,
		_w3928_
	);
	LUT3 #(
		.INIT('h48)
	) name2926 (
		_w3918_,
		_w3927_,
		_w3928_,
		_w3929_
	);
	LUT3 #(
		.INIT('h21)
	) name2927 (
		_w3918_,
		_w3927_,
		_w3928_,
		_w3930_
	);
	LUT3 #(
		.INIT('h2d)
	) name2928 (
		_w3886_,
		_w3887_,
		_w3889_,
		_w3931_
	);
	LUT2 #(
		.INIT('h6)
	) name2929 (
		_w3893_,
		_w3931_,
		_w3932_
	);
	LUT3 #(
		.INIT('h45)
	) name2930 (
		_w3929_,
		_w3930_,
		_w3932_,
		_w3933_
	);
	LUT3 #(
		.INIT('h32)
	) name2931 (
		_w3905_,
		_w3919_,
		_w3920_,
		_w3934_
	);
	LUT4 #(
		.INIT('h0017)
	) name2932 (
		_w3897_,
		_w3922_,
		_w3933_,
		_w3934_,
		_w3935_
	);
	LUT4 #(
		.INIT('he800)
	) name2933 (
		_w3897_,
		_w3922_,
		_w3933_,
		_w3934_,
		_w3936_
	);
	LUT3 #(
		.INIT('h32)
	) name2934 (
		_w3880_,
		_w3894_,
		_w3895_,
		_w3937_
	);
	LUT3 #(
		.INIT('h54)
	) name2935 (
		_w3935_,
		_w3936_,
		_w3937_,
		_w3938_
	);
	LUT4 #(
		.INIT('hab54)
	) name2936 (
		_w3923_,
		_w3924_,
		_w3933_,
		_w3934_,
		_w3939_
	);
	LUT2 #(
		.INIT('h9)
	) name2937 (
		_w3937_,
		_w3939_,
		_w3940_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		\A[610] ,
		\A[611] ,
		_w3941_
	);
	LUT3 #(
		.INIT('h96)
	) name2939 (
		\A[607] ,
		\A[608] ,
		\A[609] ,
		_w3942_
	);
	LUT3 #(
		.INIT('h96)
	) name2940 (
		\A[610] ,
		\A[611] ,
		\A[612] ,
		_w3943_
	);
	LUT3 #(
		.INIT('h80)
	) name2941 (
		_w3941_,
		_w3942_,
		_w3943_,
		_w3944_
	);
	LUT3 #(
		.INIT('h17)
	) name2942 (
		\A[607] ,
		\A[608] ,
		\A[609] ,
		_w3945_
	);
	LUT3 #(
		.INIT('h17)
	) name2943 (
		\A[610] ,
		\A[611] ,
		\A[612] ,
		_w3946_
	);
	LUT4 #(
		.INIT('h080f)
	) name2944 (
		_w3942_,
		_w3943_,
		_w3945_,
		_w3946_,
		_w3947_
	);
	LUT2 #(
		.INIT('h1)
	) name2945 (
		_w3944_,
		_w3947_,
		_w3948_
	);
	LUT3 #(
		.INIT('h17)
	) name2946 (
		\A[616] ,
		\A[617] ,
		\A[618] ,
		_w3949_
	);
	LUT3 #(
		.INIT('h17)
	) name2947 (
		\A[613] ,
		\A[614] ,
		\A[615] ,
		_w3950_
	);
	LUT3 #(
		.INIT('h96)
	) name2948 (
		\A[613] ,
		\A[614] ,
		\A[615] ,
		_w3951_
	);
	LUT3 #(
		.INIT('h96)
	) name2949 (
		\A[616] ,
		\A[617] ,
		\A[618] ,
		_w3952_
	);
	LUT4 #(
		.INIT('h7111)
	) name2950 (
		_w3949_,
		_w3950_,
		_w3951_,
		_w3952_,
		_w3953_
	);
	LUT4 #(
		.INIT('h0660)
	) name2951 (
		_w3942_,
		_w3943_,
		_w3951_,
		_w3952_,
		_w3954_
	);
	LUT4 #(
		.INIT('h0080)
	) name2952 (
		_w3941_,
		_w3942_,
		_w3943_,
		_w3945_,
		_w3955_
	);
	LUT2 #(
		.INIT('h2)
	) name2953 (
		_w3954_,
		_w3955_,
		_w3956_
	);
	LUT4 #(
		.INIT('h6999)
	) name2954 (
		_w3949_,
		_w3950_,
		_w3951_,
		_w3952_,
		_w3957_
	);
	LUT3 #(
		.INIT('h02)
	) name2955 (
		_w3954_,
		_w3955_,
		_w3957_,
		_w3958_
	);
	LUT3 #(
		.INIT('hd0)
	) name2956 (
		_w3954_,
		_w3955_,
		_w3957_,
		_w3959_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2957 (
		\A[610] ,
		\A[611] ,
		\A[612] ,
		_w3942_,
		_w3960_
	);
	LUT2 #(
		.INIT('h9)
	) name2958 (
		_w3945_,
		_w3960_,
		_w3961_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2959 (
		_w3953_,
		_w3956_,
		_w3957_,
		_w3961_,
		_w3962_
	);
	LUT4 #(
		.INIT('h1051)
	) name2960 (
		_w3953_,
		_w3956_,
		_w3957_,
		_w3961_,
		_w3963_
	);
	LUT4 #(
		.INIT('h6566)
	) name2961 (
		_w3953_,
		_w3958_,
		_w3959_,
		_w3961_,
		_w3964_
	);
	LUT2 #(
		.INIT('h6)
	) name2962 (
		_w3948_,
		_w3964_,
		_w3965_
	);
	LUT2 #(
		.INIT('h8)
	) name2963 (
		\A[622] ,
		\A[623] ,
		_w3966_
	);
	LUT3 #(
		.INIT('h96)
	) name2964 (
		\A[619] ,
		\A[620] ,
		\A[621] ,
		_w3967_
	);
	LUT3 #(
		.INIT('h96)
	) name2965 (
		\A[622] ,
		\A[623] ,
		\A[624] ,
		_w3968_
	);
	LUT3 #(
		.INIT('h80)
	) name2966 (
		_w3966_,
		_w3967_,
		_w3968_,
		_w3969_
	);
	LUT3 #(
		.INIT('h17)
	) name2967 (
		\A[619] ,
		\A[620] ,
		\A[621] ,
		_w3970_
	);
	LUT3 #(
		.INIT('h17)
	) name2968 (
		\A[622] ,
		\A[623] ,
		\A[624] ,
		_w3971_
	);
	LUT4 #(
		.INIT('h080f)
	) name2969 (
		_w3967_,
		_w3968_,
		_w3970_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h1)
	) name2970 (
		_w3969_,
		_w3972_,
		_w3973_
	);
	LUT3 #(
		.INIT('h17)
	) name2971 (
		\A[628] ,
		\A[629] ,
		\A[630] ,
		_w3974_
	);
	LUT3 #(
		.INIT('h17)
	) name2972 (
		\A[625] ,
		\A[626] ,
		\A[627] ,
		_w3975_
	);
	LUT3 #(
		.INIT('h96)
	) name2973 (
		\A[625] ,
		\A[626] ,
		\A[627] ,
		_w3976_
	);
	LUT3 #(
		.INIT('h96)
	) name2974 (
		\A[628] ,
		\A[629] ,
		\A[630] ,
		_w3977_
	);
	LUT4 #(
		.INIT('h7111)
	) name2975 (
		_w3974_,
		_w3975_,
		_w3976_,
		_w3977_,
		_w3978_
	);
	LUT4 #(
		.INIT('h0660)
	) name2976 (
		_w3967_,
		_w3968_,
		_w3976_,
		_w3977_,
		_w3979_
	);
	LUT4 #(
		.INIT('h0080)
	) name2977 (
		_w3966_,
		_w3967_,
		_w3968_,
		_w3970_,
		_w3980_
	);
	LUT2 #(
		.INIT('h2)
	) name2978 (
		_w3979_,
		_w3980_,
		_w3981_
	);
	LUT4 #(
		.INIT('h6999)
	) name2979 (
		_w3974_,
		_w3975_,
		_w3976_,
		_w3977_,
		_w3982_
	);
	LUT3 #(
		.INIT('h02)
	) name2980 (
		_w3979_,
		_w3980_,
		_w3982_,
		_w3983_
	);
	LUT3 #(
		.INIT('hd0)
	) name2981 (
		_w3979_,
		_w3980_,
		_w3982_,
		_w3984_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name2982 (
		\A[622] ,
		\A[623] ,
		\A[624] ,
		_w3967_,
		_w3985_
	);
	LUT2 #(
		.INIT('h9)
	) name2983 (
		_w3970_,
		_w3985_,
		_w3986_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2984 (
		_w3978_,
		_w3981_,
		_w3982_,
		_w3986_,
		_w3987_
	);
	LUT4 #(
		.INIT('h1051)
	) name2985 (
		_w3978_,
		_w3981_,
		_w3982_,
		_w3986_,
		_w3988_
	);
	LUT4 #(
		.INIT('h6566)
	) name2986 (
		_w3978_,
		_w3983_,
		_w3984_,
		_w3986_,
		_w3989_
	);
	LUT2 #(
		.INIT('h6)
	) name2987 (
		_w3973_,
		_w3989_,
		_w3990_
	);
	LUT4 #(
		.INIT('h9009)
	) name2988 (
		_w3948_,
		_w3964_,
		_w3973_,
		_w3989_,
		_w3991_
	);
	LUT4 #(
		.INIT('h0660)
	) name2989 (
		_w3948_,
		_w3964_,
		_w3973_,
		_w3989_,
		_w3992_
	);
	LUT4 #(
		.INIT('h6996)
	) name2990 (
		_w3967_,
		_w3968_,
		_w3976_,
		_w3977_,
		_w3993_
	);
	LUT4 #(
		.INIT('h6996)
	) name2991 (
		_w3942_,
		_w3943_,
		_w3951_,
		_w3952_,
		_w3994_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		_w3993_,
		_w3994_,
		_w3995_
	);
	LUT3 #(
		.INIT('h2d)
	) name2993 (
		_w3979_,
		_w3980_,
		_w3982_,
		_w3996_
	);
	LUT3 #(
		.INIT('h48)
	) name2994 (
		_w3986_,
		_w3995_,
		_w3996_,
		_w3997_
	);
	LUT3 #(
		.INIT('h21)
	) name2995 (
		_w3986_,
		_w3995_,
		_w3996_,
		_w3998_
	);
	LUT3 #(
		.INIT('h2d)
	) name2996 (
		_w3954_,
		_w3955_,
		_w3957_,
		_w3999_
	);
	LUT2 #(
		.INIT('h6)
	) name2997 (
		_w3961_,
		_w3999_,
		_w4000_
	);
	LUT3 #(
		.INIT('h45)
	) name2998 (
		_w3997_,
		_w3998_,
		_w4000_,
		_w4001_
	);
	LUT3 #(
		.INIT('h32)
	) name2999 (
		_w3973_,
		_w3987_,
		_w3988_,
		_w4002_
	);
	LUT4 #(
		.INIT('h0017)
	) name3000 (
		_w3965_,
		_w3990_,
		_w4001_,
		_w4002_,
		_w4003_
	);
	LUT4 #(
		.INIT('he800)
	) name3001 (
		_w3965_,
		_w3990_,
		_w4001_,
		_w4002_,
		_w4004_
	);
	LUT4 #(
		.INIT('hab54)
	) name3002 (
		_w3991_,
		_w3992_,
		_w4001_,
		_w4002_,
		_w4005_
	);
	LUT3 #(
		.INIT('h32)
	) name3003 (
		_w3948_,
		_w3962_,
		_w3963_,
		_w4006_
	);
	LUT2 #(
		.INIT('h9)
	) name3004 (
		_w4005_,
		_w4006_,
		_w4007_
	);
	LUT4 #(
		.INIT('h0660)
	) name3005 (
		_w3937_,
		_w3939_,
		_w4005_,
		_w4006_,
		_w4008_
	);
	LUT4 #(
		.INIT('h9009)
	) name3006 (
		_w3937_,
		_w3939_,
		_w4005_,
		_w4006_,
		_w4009_
	);
	LUT4 #(
		.INIT('h6996)
	) name3007 (
		_w3948_,
		_w3964_,
		_w3973_,
		_w3989_,
		_w4010_
	);
	LUT4 #(
		.INIT('h6996)
	) name3008 (
		_w3880_,
		_w3896_,
		_w3905_,
		_w3921_,
		_w4011_
	);
	LUT4 #(
		.INIT('h1428)
	) name3009 (
		_w3933_,
		_w4001_,
		_w4010_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('h8241)
	) name3010 (
		_w3933_,
		_w4001_,
		_w4010_,
		_w4011_,
		_w4013_
	);
	LUT4 #(
		.INIT('h0660)
	) name3011 (
		_w3925_,
		_w3926_,
		_w3993_,
		_w3994_,
		_w4014_
	);
	LUT3 #(
		.INIT('h96)
	) name3012 (
		_w3918_,
		_w3927_,
		_w3928_,
		_w4015_
	);
	LUT3 #(
		.INIT('h48)
	) name3013 (
		_w3932_,
		_w4014_,
		_w4015_,
		_w4016_
	);
	LUT3 #(
		.INIT('h21)
	) name3014 (
		_w3932_,
		_w4014_,
		_w4015_,
		_w4017_
	);
	LUT3 #(
		.INIT('h96)
	) name3015 (
		_w3986_,
		_w3995_,
		_w3996_,
		_w4018_
	);
	LUT2 #(
		.INIT('h9)
	) name3016 (
		_w4000_,
		_w4018_,
		_w4019_
	);
	LUT3 #(
		.INIT('h54)
	) name3017 (
		_w4016_,
		_w4017_,
		_w4019_,
		_w4020_
	);
	LUT3 #(
		.INIT('h45)
	) name3018 (
		_w4012_,
		_w4013_,
		_w4020_,
		_w4021_
	);
	LUT4 #(
		.INIT('h022a)
	) name3019 (
		_w3938_,
		_w3940_,
		_w4007_,
		_w4021_,
		_w4022_
	);
	LUT4 #(
		.INIT('h5440)
	) name3020 (
		_w3938_,
		_w3940_,
		_w4007_,
		_w4021_,
		_w4023_
	);
	LUT4 #(
		.INIT('h6665)
	) name3021 (
		_w3938_,
		_w4008_,
		_w4009_,
		_w4021_,
		_w4024_
	);
	LUT3 #(
		.INIT('h54)
	) name3022 (
		_w4003_,
		_w4004_,
		_w4006_,
		_w4025_
	);
	LUT2 #(
		.INIT('h6)
	) name3023 (
		_w4024_,
		_w4025_,
		_w4026_
	);
	LUT4 #(
		.INIT('h9009)
	) name3024 (
		_w3870_,
		_w3871_,
		_w4024_,
		_w4025_,
		_w4027_
	);
	LUT4 #(
		.INIT('h0660)
	) name3025 (
		_w3870_,
		_w3871_,
		_w4024_,
		_w4025_,
		_w4028_
	);
	LUT4 #(
		.INIT('h6996)
	) name3026 (
		_w3937_,
		_w3939_,
		_w4005_,
		_w4006_,
		_w4029_
	);
	LUT4 #(
		.INIT('h6996)
	) name3027 (
		_w3783_,
		_w3849_,
		_w3850_,
		_w3852_,
		_w4030_
	);
	LUT4 #(
		.INIT('h1428)
	) name3028 (
		_w3867_,
		_w4021_,
		_w4029_,
		_w4030_,
		_w4031_
	);
	LUT4 #(
		.INIT('h8241)
	) name3029 (
		_w3867_,
		_w4021_,
		_w4029_,
		_w4030_,
		_w4032_
	);
	LUT4 #(
		.INIT('h6996)
	) name3030 (
		_w3779_,
		_w3845_,
		_w3856_,
		_w3857_,
		_w4033_
	);
	LUT4 #(
		.INIT('h6996)
	) name3031 (
		_w3933_,
		_w4001_,
		_w4010_,
		_w4011_,
		_w4034_
	);
	LUT4 #(
		.INIT('h1248)
	) name3032 (
		_w3866_,
		_w4020_,
		_w4033_,
		_w4034_,
		_w4035_
	);
	LUT4 #(
		.INIT('h8421)
	) name3033 (
		_w3866_,
		_w4020_,
		_w4033_,
		_w4034_,
		_w4036_
	);
	LUT4 #(
		.INIT('h6996)
	) name3034 (
		_w3925_,
		_w3926_,
		_w3993_,
		_w3994_,
		_w4037_
	);
	LUT4 #(
		.INIT('h6996)
	) name3035 (
		_w3771_,
		_w3772_,
		_w3837_,
		_w3838_,
		_w4038_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		_w4037_,
		_w4038_,
		_w4039_
	);
	LUT3 #(
		.INIT('h96)
	) name3037 (
		_w3932_,
		_w4014_,
		_w4015_,
		_w4040_
	);
	LUT3 #(
		.INIT('h84)
	) name3038 (
		_w4019_,
		_w4039_,
		_w4040_,
		_w4041_
	);
	LUT3 #(
		.INIT('h12)
	) name3039 (
		_w4019_,
		_w4039_,
		_w4040_,
		_w4042_
	);
	LUT3 #(
		.INIT('h96)
	) name3040 (
		_w3844_,
		_w3860_,
		_w3861_,
		_w4043_
	);
	LUT2 #(
		.INIT('h9)
	) name3041 (
		_w3865_,
		_w4043_,
		_w4044_
	);
	LUT3 #(
		.INIT('h45)
	) name3042 (
		_w4041_,
		_w4042_,
		_w4044_,
		_w4045_
	);
	LUT3 #(
		.INIT('h45)
	) name3043 (
		_w4035_,
		_w4036_,
		_w4045_,
		_w4046_
	);
	LUT3 #(
		.INIT('h45)
	) name3044 (
		_w4031_,
		_w4032_,
		_w4046_,
		_w4047_
	);
	LUT3 #(
		.INIT('h45)
	) name3045 (
		_w3868_,
		_w3869_,
		_w3871_,
		_w4048_
	);
	LUT4 #(
		.INIT('h00e8)
	) name3046 (
		_w3872_,
		_w4026_,
		_w4047_,
		_w4048_,
		_w4049_
	);
	LUT4 #(
		.INIT('h1700)
	) name3047 (
		_w3872_,
		_w4026_,
		_w4047_,
		_w4048_,
		_w4050_
	);
	LUT3 #(
		.INIT('h45)
	) name3048 (
		_w4022_,
		_w4023_,
		_w4025_,
		_w4051_
	);
	LUT3 #(
		.INIT('h54)
	) name3049 (
		_w4049_,
		_w4050_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		\A[466] ,
		\A[467] ,
		_w4053_
	);
	LUT2 #(
		.INIT('h6)
	) name3051 (
		\A[466] ,
		\A[467] ,
		_w4054_
	);
	LUT3 #(
		.INIT('h96)
	) name3052 (
		\A[466] ,
		\A[467] ,
		\A[468] ,
		_w4055_
	);
	LUT3 #(
		.INIT('h96)
	) name3053 (
		\A[463] ,
		\A[464] ,
		\A[465] ,
		_w4056_
	);
	LUT3 #(
		.INIT('h80)
	) name3054 (
		_w4053_,
		_w4055_,
		_w4056_,
		_w4057_
	);
	LUT3 #(
		.INIT('h17)
	) name3055 (
		\A[463] ,
		\A[464] ,
		\A[465] ,
		_w4058_
	);
	LUT3 #(
		.INIT('h17)
	) name3056 (
		\A[466] ,
		\A[467] ,
		\A[468] ,
		_w4059_
	);
	LUT4 #(
		.INIT('h080f)
	) name3057 (
		_w4055_,
		_w4056_,
		_w4058_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h1)
	) name3058 (
		_w4057_,
		_w4060_,
		_w4061_
	);
	LUT3 #(
		.INIT('h17)
	) name3059 (
		\A[472] ,
		\A[473] ,
		\A[474] ,
		_w4062_
	);
	LUT3 #(
		.INIT('h17)
	) name3060 (
		\A[469] ,
		\A[470] ,
		\A[471] ,
		_w4063_
	);
	LUT3 #(
		.INIT('h96)
	) name3061 (
		\A[469] ,
		\A[470] ,
		\A[471] ,
		_w4064_
	);
	LUT3 #(
		.INIT('h96)
	) name3062 (
		\A[472] ,
		\A[473] ,
		\A[474] ,
		_w4065_
	);
	LUT4 #(
		.INIT('h7111)
	) name3063 (
		_w4062_,
		_w4063_,
		_w4064_,
		_w4065_,
		_w4066_
	);
	LUT4 #(
		.INIT('h0660)
	) name3064 (
		_w4055_,
		_w4056_,
		_w4064_,
		_w4065_,
		_w4067_
	);
	LUT4 #(
		.INIT('h0080)
	) name3065 (
		_w4053_,
		_w4055_,
		_w4056_,
		_w4058_,
		_w4068_
	);
	LUT2 #(
		.INIT('h2)
	) name3066 (
		_w4067_,
		_w4068_,
		_w4069_
	);
	LUT4 #(
		.INIT('h6999)
	) name3067 (
		_w4062_,
		_w4063_,
		_w4064_,
		_w4065_,
		_w4070_
	);
	LUT3 #(
		.INIT('h02)
	) name3068 (
		_w4067_,
		_w4068_,
		_w4070_,
		_w4071_
	);
	LUT3 #(
		.INIT('hd0)
	) name3069 (
		_w4067_,
		_w4068_,
		_w4070_,
		_w4072_
	);
	LUT4 #(
		.INIT('hb6ec)
	) name3070 (
		\A[468] ,
		_w4053_,
		_w4054_,
		_w4056_,
		_w4073_
	);
	LUT2 #(
		.INIT('h9)
	) name3071 (
		_w4058_,
		_w4073_,
		_w4074_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3072 (
		_w4066_,
		_w4069_,
		_w4070_,
		_w4074_,
		_w4075_
	);
	LUT4 #(
		.INIT('h1051)
	) name3073 (
		_w4066_,
		_w4069_,
		_w4070_,
		_w4074_,
		_w4076_
	);
	LUT4 #(
		.INIT('h6566)
	) name3074 (
		_w4066_,
		_w4071_,
		_w4072_,
		_w4074_,
		_w4077_
	);
	LUT2 #(
		.INIT('h6)
	) name3075 (
		_w4061_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h8)
	) name3076 (
		\A[478] ,
		\A[479] ,
		_w4079_
	);
	LUT3 #(
		.INIT('h96)
	) name3077 (
		\A[475] ,
		\A[476] ,
		\A[477] ,
		_w4080_
	);
	LUT3 #(
		.INIT('h96)
	) name3078 (
		\A[478] ,
		\A[479] ,
		\A[480] ,
		_w4081_
	);
	LUT3 #(
		.INIT('h80)
	) name3079 (
		_w4079_,
		_w4080_,
		_w4081_,
		_w4082_
	);
	LUT3 #(
		.INIT('h17)
	) name3080 (
		\A[475] ,
		\A[476] ,
		\A[477] ,
		_w4083_
	);
	LUT3 #(
		.INIT('h17)
	) name3081 (
		\A[478] ,
		\A[479] ,
		\A[480] ,
		_w4084_
	);
	LUT4 #(
		.INIT('h080f)
	) name3082 (
		_w4080_,
		_w4081_,
		_w4083_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name3083 (
		_w4082_,
		_w4085_,
		_w4086_
	);
	LUT3 #(
		.INIT('h17)
	) name3084 (
		\A[484] ,
		\A[485] ,
		\A[486] ,
		_w4087_
	);
	LUT3 #(
		.INIT('h17)
	) name3085 (
		\A[481] ,
		\A[482] ,
		\A[483] ,
		_w4088_
	);
	LUT3 #(
		.INIT('h96)
	) name3086 (
		\A[481] ,
		\A[482] ,
		\A[483] ,
		_w4089_
	);
	LUT3 #(
		.INIT('h96)
	) name3087 (
		\A[484] ,
		\A[485] ,
		\A[486] ,
		_w4090_
	);
	LUT4 #(
		.INIT('h7111)
	) name3088 (
		_w4087_,
		_w4088_,
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT4 #(
		.INIT('h0660)
	) name3089 (
		_w4080_,
		_w4081_,
		_w4089_,
		_w4090_,
		_w4092_
	);
	LUT4 #(
		.INIT('h0080)
	) name3090 (
		_w4079_,
		_w4080_,
		_w4081_,
		_w4083_,
		_w4093_
	);
	LUT2 #(
		.INIT('h2)
	) name3091 (
		_w4092_,
		_w4093_,
		_w4094_
	);
	LUT4 #(
		.INIT('h6999)
	) name3092 (
		_w4087_,
		_w4088_,
		_w4089_,
		_w4090_,
		_w4095_
	);
	LUT3 #(
		.INIT('h02)
	) name3093 (
		_w4092_,
		_w4093_,
		_w4095_,
		_w4096_
	);
	LUT3 #(
		.INIT('hd0)
	) name3094 (
		_w4092_,
		_w4093_,
		_w4095_,
		_w4097_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name3095 (
		\A[478] ,
		\A[479] ,
		\A[480] ,
		_w4080_,
		_w4098_
	);
	LUT2 #(
		.INIT('h9)
	) name3096 (
		_w4083_,
		_w4098_,
		_w4099_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3097 (
		_w4091_,
		_w4094_,
		_w4095_,
		_w4099_,
		_w4100_
	);
	LUT4 #(
		.INIT('h1051)
	) name3098 (
		_w4091_,
		_w4094_,
		_w4095_,
		_w4099_,
		_w4101_
	);
	LUT4 #(
		.INIT('h6566)
	) name3099 (
		_w4091_,
		_w4096_,
		_w4097_,
		_w4099_,
		_w4102_
	);
	LUT2 #(
		.INIT('h6)
	) name3100 (
		_w4086_,
		_w4102_,
		_w4103_
	);
	LUT4 #(
		.INIT('h9009)
	) name3101 (
		_w4061_,
		_w4077_,
		_w4086_,
		_w4102_,
		_w4104_
	);
	LUT4 #(
		.INIT('h0660)
	) name3102 (
		_w4061_,
		_w4077_,
		_w4086_,
		_w4102_,
		_w4105_
	);
	LUT4 #(
		.INIT('h6996)
	) name3103 (
		_w4055_,
		_w4056_,
		_w4064_,
		_w4065_,
		_w4106_
	);
	LUT4 #(
		.INIT('h6996)
	) name3104 (
		_w4080_,
		_w4081_,
		_w4089_,
		_w4090_,
		_w4107_
	);
	LUT2 #(
		.INIT('h8)
	) name3105 (
		_w4106_,
		_w4107_,
		_w4108_
	);
	LUT3 #(
		.INIT('h2d)
	) name3106 (
		_w4092_,
		_w4093_,
		_w4095_,
		_w4109_
	);
	LUT3 #(
		.INIT('h48)
	) name3107 (
		_w4099_,
		_w4108_,
		_w4109_,
		_w4110_
	);
	LUT3 #(
		.INIT('h21)
	) name3108 (
		_w4099_,
		_w4108_,
		_w4109_,
		_w4111_
	);
	LUT3 #(
		.INIT('h2d)
	) name3109 (
		_w4067_,
		_w4068_,
		_w4070_,
		_w4112_
	);
	LUT2 #(
		.INIT('h6)
	) name3110 (
		_w4074_,
		_w4112_,
		_w4113_
	);
	LUT3 #(
		.INIT('h45)
	) name3111 (
		_w4110_,
		_w4111_,
		_w4113_,
		_w4114_
	);
	LUT3 #(
		.INIT('h32)
	) name3112 (
		_w4086_,
		_w4100_,
		_w4101_,
		_w4115_
	);
	LUT4 #(
		.INIT('h0017)
	) name3113 (
		_w4078_,
		_w4103_,
		_w4114_,
		_w4115_,
		_w4116_
	);
	LUT4 #(
		.INIT('he800)
	) name3114 (
		_w4078_,
		_w4103_,
		_w4114_,
		_w4115_,
		_w4117_
	);
	LUT3 #(
		.INIT('h32)
	) name3115 (
		_w4061_,
		_w4075_,
		_w4076_,
		_w4118_
	);
	LUT3 #(
		.INIT('h54)
	) name3116 (
		_w4116_,
		_w4117_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		\A[490] ,
		\A[491] ,
		_w4120_
	);
	LUT3 #(
		.INIT('h96)
	) name3118 (
		\A[487] ,
		\A[488] ,
		\A[489] ,
		_w4121_
	);
	LUT3 #(
		.INIT('h96)
	) name3119 (
		\A[490] ,
		\A[491] ,
		\A[492] ,
		_w4122_
	);
	LUT3 #(
		.INIT('h80)
	) name3120 (
		_w4120_,
		_w4121_,
		_w4122_,
		_w4123_
	);
	LUT3 #(
		.INIT('h17)
	) name3121 (
		\A[487] ,
		\A[488] ,
		\A[489] ,
		_w4124_
	);
	LUT3 #(
		.INIT('h17)
	) name3122 (
		\A[490] ,
		\A[491] ,
		\A[492] ,
		_w4125_
	);
	LUT4 #(
		.INIT('h080f)
	) name3123 (
		_w4121_,
		_w4122_,
		_w4124_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h1)
	) name3124 (
		_w4123_,
		_w4126_,
		_w4127_
	);
	LUT3 #(
		.INIT('h17)
	) name3125 (
		\A[496] ,
		\A[497] ,
		\A[498] ,
		_w4128_
	);
	LUT3 #(
		.INIT('h17)
	) name3126 (
		\A[493] ,
		\A[494] ,
		\A[495] ,
		_w4129_
	);
	LUT3 #(
		.INIT('h96)
	) name3127 (
		\A[493] ,
		\A[494] ,
		\A[495] ,
		_w4130_
	);
	LUT3 #(
		.INIT('h96)
	) name3128 (
		\A[496] ,
		\A[497] ,
		\A[498] ,
		_w4131_
	);
	LUT4 #(
		.INIT('h7111)
	) name3129 (
		_w4128_,
		_w4129_,
		_w4130_,
		_w4131_,
		_w4132_
	);
	LUT4 #(
		.INIT('h0660)
	) name3130 (
		_w4121_,
		_w4122_,
		_w4130_,
		_w4131_,
		_w4133_
	);
	LUT4 #(
		.INIT('h0080)
	) name3131 (
		_w4120_,
		_w4121_,
		_w4122_,
		_w4124_,
		_w4134_
	);
	LUT2 #(
		.INIT('h2)
	) name3132 (
		_w4133_,
		_w4134_,
		_w4135_
	);
	LUT4 #(
		.INIT('h6999)
	) name3133 (
		_w4128_,
		_w4129_,
		_w4130_,
		_w4131_,
		_w4136_
	);
	LUT3 #(
		.INIT('h02)
	) name3134 (
		_w4133_,
		_w4134_,
		_w4136_,
		_w4137_
	);
	LUT3 #(
		.INIT('hd0)
	) name3135 (
		_w4133_,
		_w4134_,
		_w4136_,
		_w4138_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name3136 (
		\A[490] ,
		\A[491] ,
		\A[492] ,
		_w4121_,
		_w4139_
	);
	LUT2 #(
		.INIT('h9)
	) name3137 (
		_w4124_,
		_w4139_,
		_w4140_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3138 (
		_w4132_,
		_w4135_,
		_w4136_,
		_w4140_,
		_w4141_
	);
	LUT4 #(
		.INIT('h1051)
	) name3139 (
		_w4132_,
		_w4135_,
		_w4136_,
		_w4140_,
		_w4142_
	);
	LUT4 #(
		.INIT('h6566)
	) name3140 (
		_w4132_,
		_w4137_,
		_w4138_,
		_w4140_,
		_w4143_
	);
	LUT2 #(
		.INIT('h6)
	) name3141 (
		_w4127_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		\A[502] ,
		\A[503] ,
		_w4145_
	);
	LUT3 #(
		.INIT('h96)
	) name3143 (
		\A[499] ,
		\A[500] ,
		\A[501] ,
		_w4146_
	);
	LUT3 #(
		.INIT('h96)
	) name3144 (
		\A[502] ,
		\A[503] ,
		\A[504] ,
		_w4147_
	);
	LUT3 #(
		.INIT('h80)
	) name3145 (
		_w4145_,
		_w4146_,
		_w4147_,
		_w4148_
	);
	LUT3 #(
		.INIT('h17)
	) name3146 (
		\A[499] ,
		\A[500] ,
		\A[501] ,
		_w4149_
	);
	LUT3 #(
		.INIT('h17)
	) name3147 (
		\A[502] ,
		\A[503] ,
		\A[504] ,
		_w4150_
	);
	LUT4 #(
		.INIT('h080f)
	) name3148 (
		_w4146_,
		_w4147_,
		_w4149_,
		_w4150_,
		_w4151_
	);
	LUT2 #(
		.INIT('h1)
	) name3149 (
		_w4148_,
		_w4151_,
		_w4152_
	);
	LUT3 #(
		.INIT('h17)
	) name3150 (
		\A[508] ,
		\A[509] ,
		\A[510] ,
		_w4153_
	);
	LUT3 #(
		.INIT('h17)
	) name3151 (
		\A[505] ,
		\A[506] ,
		\A[507] ,
		_w4154_
	);
	LUT3 #(
		.INIT('h96)
	) name3152 (
		\A[505] ,
		\A[506] ,
		\A[507] ,
		_w4155_
	);
	LUT3 #(
		.INIT('h96)
	) name3153 (
		\A[508] ,
		\A[509] ,
		\A[510] ,
		_w4156_
	);
	LUT4 #(
		.INIT('h7111)
	) name3154 (
		_w4153_,
		_w4154_,
		_w4155_,
		_w4156_,
		_w4157_
	);
	LUT4 #(
		.INIT('h0660)
	) name3155 (
		_w4146_,
		_w4147_,
		_w4155_,
		_w4156_,
		_w4158_
	);
	LUT4 #(
		.INIT('h0080)
	) name3156 (
		_w4145_,
		_w4146_,
		_w4147_,
		_w4149_,
		_w4159_
	);
	LUT2 #(
		.INIT('h2)
	) name3157 (
		_w4158_,
		_w4159_,
		_w4160_
	);
	LUT4 #(
		.INIT('h6999)
	) name3158 (
		_w4153_,
		_w4154_,
		_w4155_,
		_w4156_,
		_w4161_
	);
	LUT3 #(
		.INIT('h02)
	) name3159 (
		_w4158_,
		_w4159_,
		_w4161_,
		_w4162_
	);
	LUT3 #(
		.INIT('hd0)
	) name3160 (
		_w4158_,
		_w4159_,
		_w4161_,
		_w4163_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name3161 (
		\A[502] ,
		\A[503] ,
		\A[504] ,
		_w4146_,
		_w4164_
	);
	LUT2 #(
		.INIT('h9)
	) name3162 (
		_w4149_,
		_w4164_,
		_w4165_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3163 (
		_w4157_,
		_w4160_,
		_w4161_,
		_w4165_,
		_w4166_
	);
	LUT4 #(
		.INIT('h1051)
	) name3164 (
		_w4157_,
		_w4160_,
		_w4161_,
		_w4165_,
		_w4167_
	);
	LUT4 #(
		.INIT('h6566)
	) name3165 (
		_w4157_,
		_w4162_,
		_w4163_,
		_w4165_,
		_w4168_
	);
	LUT2 #(
		.INIT('h6)
	) name3166 (
		_w4152_,
		_w4168_,
		_w4169_
	);
	LUT4 #(
		.INIT('h9009)
	) name3167 (
		_w4127_,
		_w4143_,
		_w4152_,
		_w4168_,
		_w4170_
	);
	LUT4 #(
		.INIT('h0660)
	) name3168 (
		_w4127_,
		_w4143_,
		_w4152_,
		_w4168_,
		_w4171_
	);
	LUT4 #(
		.INIT('h6996)
	) name3169 (
		_w4146_,
		_w4147_,
		_w4155_,
		_w4156_,
		_w4172_
	);
	LUT4 #(
		.INIT('h6996)
	) name3170 (
		_w4121_,
		_w4122_,
		_w4130_,
		_w4131_,
		_w4173_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		_w4172_,
		_w4173_,
		_w4174_
	);
	LUT3 #(
		.INIT('h2d)
	) name3172 (
		_w4158_,
		_w4159_,
		_w4161_,
		_w4175_
	);
	LUT3 #(
		.INIT('h48)
	) name3173 (
		_w4165_,
		_w4174_,
		_w4175_,
		_w4176_
	);
	LUT3 #(
		.INIT('h21)
	) name3174 (
		_w4165_,
		_w4174_,
		_w4175_,
		_w4177_
	);
	LUT3 #(
		.INIT('h2d)
	) name3175 (
		_w4133_,
		_w4134_,
		_w4136_,
		_w4178_
	);
	LUT2 #(
		.INIT('h6)
	) name3176 (
		_w4140_,
		_w4178_,
		_w4179_
	);
	LUT3 #(
		.INIT('h45)
	) name3177 (
		_w4176_,
		_w4177_,
		_w4179_,
		_w4180_
	);
	LUT3 #(
		.INIT('h32)
	) name3178 (
		_w4152_,
		_w4166_,
		_w4167_,
		_w4181_
	);
	LUT4 #(
		.INIT('h0017)
	) name3179 (
		_w4144_,
		_w4169_,
		_w4180_,
		_w4181_,
		_w4182_
	);
	LUT4 #(
		.INIT('he800)
	) name3180 (
		_w4144_,
		_w4169_,
		_w4180_,
		_w4181_,
		_w4183_
	);
	LUT4 #(
		.INIT('hab54)
	) name3181 (
		_w4170_,
		_w4171_,
		_w4180_,
		_w4181_,
		_w4184_
	);
	LUT3 #(
		.INIT('h32)
	) name3182 (
		_w4127_,
		_w4141_,
		_w4142_,
		_w4185_
	);
	LUT2 #(
		.INIT('h9)
	) name3183 (
		_w4184_,
		_w4185_,
		_w4186_
	);
	LUT4 #(
		.INIT('hab54)
	) name3184 (
		_w4104_,
		_w4105_,
		_w4114_,
		_w4115_,
		_w4187_
	);
	LUT2 #(
		.INIT('h9)
	) name3185 (
		_w4118_,
		_w4187_,
		_w4188_
	);
	LUT4 #(
		.INIT('h1428)
	) name3186 (
		_w4118_,
		_w4184_,
		_w4185_,
		_w4187_,
		_w4189_
	);
	LUT4 #(
		.INIT('h8241)
	) name3187 (
		_w4118_,
		_w4184_,
		_w4185_,
		_w4187_,
		_w4190_
	);
	LUT4 #(
		.INIT('h6996)
	) name3188 (
		_w4061_,
		_w4077_,
		_w4086_,
		_w4102_,
		_w4191_
	);
	LUT4 #(
		.INIT('h6996)
	) name3189 (
		_w4127_,
		_w4143_,
		_w4152_,
		_w4168_,
		_w4192_
	);
	LUT4 #(
		.INIT('h1248)
	) name3190 (
		_w4114_,
		_w4180_,
		_w4191_,
		_w4192_,
		_w4193_
	);
	LUT4 #(
		.INIT('h8421)
	) name3191 (
		_w4114_,
		_w4180_,
		_w4191_,
		_w4192_,
		_w4194_
	);
	LUT4 #(
		.INIT('h0660)
	) name3192 (
		_w4106_,
		_w4107_,
		_w4172_,
		_w4173_,
		_w4195_
	);
	LUT3 #(
		.INIT('h96)
	) name3193 (
		_w4165_,
		_w4174_,
		_w4175_,
		_w4196_
	);
	LUT3 #(
		.INIT('h48)
	) name3194 (
		_w4179_,
		_w4195_,
		_w4196_,
		_w4197_
	);
	LUT3 #(
		.INIT('h21)
	) name3195 (
		_w4179_,
		_w4195_,
		_w4196_,
		_w4198_
	);
	LUT3 #(
		.INIT('h96)
	) name3196 (
		_w4099_,
		_w4108_,
		_w4109_,
		_w4199_
	);
	LUT2 #(
		.INIT('h9)
	) name3197 (
		_w4113_,
		_w4199_,
		_w4200_
	);
	LUT3 #(
		.INIT('h54)
	) name3198 (
		_w4197_,
		_w4198_,
		_w4200_,
		_w4201_
	);
	LUT3 #(
		.INIT('h45)
	) name3199 (
		_w4193_,
		_w4194_,
		_w4201_,
		_w4202_
	);
	LUT4 #(
		.INIT('h022a)
	) name3200 (
		_w4119_,
		_w4186_,
		_w4188_,
		_w4202_,
		_w4203_
	);
	LUT4 #(
		.INIT('h5440)
	) name3201 (
		_w4119_,
		_w4186_,
		_w4188_,
		_w4202_,
		_w4204_
	);
	LUT4 #(
		.INIT('h6665)
	) name3202 (
		_w4119_,
		_w4189_,
		_w4190_,
		_w4202_,
		_w4205_
	);
	LUT3 #(
		.INIT('h54)
	) name3203 (
		_w4182_,
		_w4183_,
		_w4185_,
		_w4206_
	);
	LUT2 #(
		.INIT('h6)
	) name3204 (
		_w4205_,
		_w4206_,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name3205 (
		\A[538] ,
		\A[539] ,
		_w4208_
	);
	LUT3 #(
		.INIT('h96)
	) name3206 (
		\A[535] ,
		\A[536] ,
		\A[537] ,
		_w4209_
	);
	LUT3 #(
		.INIT('h96)
	) name3207 (
		\A[538] ,
		\A[539] ,
		\A[540] ,
		_w4210_
	);
	LUT3 #(
		.INIT('h80)
	) name3208 (
		_w4208_,
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT3 #(
		.INIT('h17)
	) name3209 (
		\A[535] ,
		\A[536] ,
		\A[537] ,
		_w4212_
	);
	LUT3 #(
		.INIT('h17)
	) name3210 (
		\A[538] ,
		\A[539] ,
		\A[540] ,
		_w4213_
	);
	LUT4 #(
		.INIT('h080f)
	) name3211 (
		_w4209_,
		_w4210_,
		_w4212_,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h1)
	) name3212 (
		_w4211_,
		_w4214_,
		_w4215_
	);
	LUT3 #(
		.INIT('h17)
	) name3213 (
		\A[544] ,
		\A[545] ,
		\A[546] ,
		_w4216_
	);
	LUT3 #(
		.INIT('h17)
	) name3214 (
		\A[541] ,
		\A[542] ,
		\A[543] ,
		_w4217_
	);
	LUT3 #(
		.INIT('h96)
	) name3215 (
		\A[541] ,
		\A[542] ,
		\A[543] ,
		_w4218_
	);
	LUT3 #(
		.INIT('h96)
	) name3216 (
		\A[544] ,
		\A[545] ,
		\A[546] ,
		_w4219_
	);
	LUT4 #(
		.INIT('h7111)
	) name3217 (
		_w4216_,
		_w4217_,
		_w4218_,
		_w4219_,
		_w4220_
	);
	LUT4 #(
		.INIT('h0660)
	) name3218 (
		_w4209_,
		_w4210_,
		_w4218_,
		_w4219_,
		_w4221_
	);
	LUT4 #(
		.INIT('h0080)
	) name3219 (
		_w4208_,
		_w4209_,
		_w4210_,
		_w4212_,
		_w4222_
	);
	LUT2 #(
		.INIT('h2)
	) name3220 (
		_w4221_,
		_w4222_,
		_w4223_
	);
	LUT4 #(
		.INIT('h6999)
	) name3221 (
		_w4216_,
		_w4217_,
		_w4218_,
		_w4219_,
		_w4224_
	);
	LUT3 #(
		.INIT('h02)
	) name3222 (
		_w4221_,
		_w4222_,
		_w4224_,
		_w4225_
	);
	LUT3 #(
		.INIT('hd0)
	) name3223 (
		_w4221_,
		_w4222_,
		_w4224_,
		_w4226_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name3224 (
		\A[538] ,
		\A[539] ,
		\A[540] ,
		_w4209_,
		_w4227_
	);
	LUT2 #(
		.INIT('h9)
	) name3225 (
		_w4212_,
		_w4227_,
		_w4228_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3226 (
		_w4220_,
		_w4223_,
		_w4224_,
		_w4228_,
		_w4229_
	);
	LUT4 #(
		.INIT('h1051)
	) name3227 (
		_w4220_,
		_w4223_,
		_w4224_,
		_w4228_,
		_w4230_
	);
	LUT4 #(
		.INIT('h6566)
	) name3228 (
		_w4220_,
		_w4225_,
		_w4226_,
		_w4228_,
		_w4231_
	);
	LUT2 #(
		.INIT('h6)
	) name3229 (
		_w4215_,
		_w4231_,
		_w4232_
	);
	LUT2 #(
		.INIT('h8)
	) name3230 (
		\A[550] ,
		\A[551] ,
		_w4233_
	);
	LUT3 #(
		.INIT('h96)
	) name3231 (
		\A[547] ,
		\A[548] ,
		\A[549] ,
		_w4234_
	);
	LUT3 #(
		.INIT('h96)
	) name3232 (
		\A[550] ,
		\A[551] ,
		\A[552] ,
		_w4235_
	);
	LUT3 #(
		.INIT('h80)
	) name3233 (
		_w4233_,
		_w4234_,
		_w4235_,
		_w4236_
	);
	LUT3 #(
		.INIT('h17)
	) name3234 (
		\A[547] ,
		\A[548] ,
		\A[549] ,
		_w4237_
	);
	LUT3 #(
		.INIT('h17)
	) name3235 (
		\A[550] ,
		\A[551] ,
		\A[552] ,
		_w4238_
	);
	LUT4 #(
		.INIT('h080f)
	) name3236 (
		_w4234_,
		_w4235_,
		_w4237_,
		_w4238_,
		_w4239_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w4236_,
		_w4239_,
		_w4240_
	);
	LUT3 #(
		.INIT('h17)
	) name3238 (
		\A[556] ,
		\A[557] ,
		\A[558] ,
		_w4241_
	);
	LUT3 #(
		.INIT('h17)
	) name3239 (
		\A[553] ,
		\A[554] ,
		\A[555] ,
		_w4242_
	);
	LUT3 #(
		.INIT('h96)
	) name3240 (
		\A[553] ,
		\A[554] ,
		\A[555] ,
		_w4243_
	);
	LUT3 #(
		.INIT('h96)
	) name3241 (
		\A[556] ,
		\A[557] ,
		\A[558] ,
		_w4244_
	);
	LUT4 #(
		.INIT('h7111)
	) name3242 (
		_w4241_,
		_w4242_,
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT4 #(
		.INIT('h0660)
	) name3243 (
		_w4234_,
		_w4235_,
		_w4243_,
		_w4244_,
		_w4246_
	);
	LUT4 #(
		.INIT('h0080)
	) name3244 (
		_w4233_,
		_w4234_,
		_w4235_,
		_w4237_,
		_w4247_
	);
	LUT2 #(
		.INIT('h2)
	) name3245 (
		_w4246_,
		_w4247_,
		_w4248_
	);
	LUT4 #(
		.INIT('h6999)
	) name3246 (
		_w4241_,
		_w4242_,
		_w4243_,
		_w4244_,
		_w4249_
	);
	LUT3 #(
		.INIT('h02)
	) name3247 (
		_w4246_,
		_w4247_,
		_w4249_,
		_w4250_
	);
	LUT3 #(
		.INIT('hd0)
	) name3248 (
		_w4246_,
		_w4247_,
		_w4249_,
		_w4251_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name3249 (
		\A[550] ,
		\A[551] ,
		\A[552] ,
		_w4234_,
		_w4252_
	);
	LUT2 #(
		.INIT('h9)
	) name3250 (
		_w4237_,
		_w4252_,
		_w4253_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3251 (
		_w4245_,
		_w4248_,
		_w4249_,
		_w4253_,
		_w4254_
	);
	LUT4 #(
		.INIT('h1051)
	) name3252 (
		_w4245_,
		_w4248_,
		_w4249_,
		_w4253_,
		_w4255_
	);
	LUT4 #(
		.INIT('h6566)
	) name3253 (
		_w4245_,
		_w4250_,
		_w4251_,
		_w4253_,
		_w4256_
	);
	LUT2 #(
		.INIT('h6)
	) name3254 (
		_w4240_,
		_w4256_,
		_w4257_
	);
	LUT4 #(
		.INIT('h9009)
	) name3255 (
		_w4215_,
		_w4231_,
		_w4240_,
		_w4256_,
		_w4258_
	);
	LUT4 #(
		.INIT('h0660)
	) name3256 (
		_w4215_,
		_w4231_,
		_w4240_,
		_w4256_,
		_w4259_
	);
	LUT4 #(
		.INIT('h6996)
	) name3257 (
		_w4234_,
		_w4235_,
		_w4243_,
		_w4244_,
		_w4260_
	);
	LUT4 #(
		.INIT('h6996)
	) name3258 (
		_w4209_,
		_w4210_,
		_w4218_,
		_w4219_,
		_w4261_
	);
	LUT2 #(
		.INIT('h8)
	) name3259 (
		_w4260_,
		_w4261_,
		_w4262_
	);
	LUT3 #(
		.INIT('h2d)
	) name3260 (
		_w4246_,
		_w4247_,
		_w4249_,
		_w4263_
	);
	LUT3 #(
		.INIT('h48)
	) name3261 (
		_w4253_,
		_w4262_,
		_w4263_,
		_w4264_
	);
	LUT3 #(
		.INIT('h21)
	) name3262 (
		_w4253_,
		_w4262_,
		_w4263_,
		_w4265_
	);
	LUT3 #(
		.INIT('h2d)
	) name3263 (
		_w4221_,
		_w4222_,
		_w4224_,
		_w4266_
	);
	LUT2 #(
		.INIT('h6)
	) name3264 (
		_w4228_,
		_w4266_,
		_w4267_
	);
	LUT3 #(
		.INIT('h45)
	) name3265 (
		_w4264_,
		_w4265_,
		_w4267_,
		_w4268_
	);
	LUT3 #(
		.INIT('h32)
	) name3266 (
		_w4240_,
		_w4254_,
		_w4255_,
		_w4269_
	);
	LUT4 #(
		.INIT('h0017)
	) name3267 (
		_w4232_,
		_w4257_,
		_w4268_,
		_w4269_,
		_w4270_
	);
	LUT4 #(
		.INIT('he800)
	) name3268 (
		_w4232_,
		_w4257_,
		_w4268_,
		_w4269_,
		_w4271_
	);
	LUT3 #(
		.INIT('h32)
	) name3269 (
		_w4215_,
		_w4229_,
		_w4230_,
		_w4272_
	);
	LUT3 #(
		.INIT('h54)
	) name3270 (
		_w4270_,
		_w4271_,
		_w4272_,
		_w4273_
	);
	LUT4 #(
		.INIT('hab54)
	) name3271 (
		_w4258_,
		_w4259_,
		_w4268_,
		_w4269_,
		_w4274_
	);
	LUT2 #(
		.INIT('h9)
	) name3272 (
		_w4272_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name3273 (
		\A[514] ,
		\A[515] ,
		_w4276_
	);
	LUT3 #(
		.INIT('h96)
	) name3274 (
		\A[511] ,
		\A[512] ,
		\A[513] ,
		_w4277_
	);
	LUT3 #(
		.INIT('h96)
	) name3275 (
		\A[514] ,
		\A[515] ,
		\A[516] ,
		_w4278_
	);
	LUT3 #(
		.INIT('h80)
	) name3276 (
		_w4276_,
		_w4277_,
		_w4278_,
		_w4279_
	);
	LUT3 #(
		.INIT('h17)
	) name3277 (
		\A[511] ,
		\A[512] ,
		\A[513] ,
		_w4280_
	);
	LUT3 #(
		.INIT('h17)
	) name3278 (
		\A[514] ,
		\A[515] ,
		\A[516] ,
		_w4281_
	);
	LUT4 #(
		.INIT('h080f)
	) name3279 (
		_w4277_,
		_w4278_,
		_w4280_,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h1)
	) name3280 (
		_w4279_,
		_w4282_,
		_w4283_
	);
	LUT3 #(
		.INIT('h17)
	) name3281 (
		\A[520] ,
		\A[521] ,
		\A[522] ,
		_w4284_
	);
	LUT3 #(
		.INIT('h17)
	) name3282 (
		\A[517] ,
		\A[518] ,
		\A[519] ,
		_w4285_
	);
	LUT3 #(
		.INIT('h96)
	) name3283 (
		\A[517] ,
		\A[518] ,
		\A[519] ,
		_w4286_
	);
	LUT3 #(
		.INIT('h96)
	) name3284 (
		\A[520] ,
		\A[521] ,
		\A[522] ,
		_w4287_
	);
	LUT4 #(
		.INIT('h7111)
	) name3285 (
		_w4284_,
		_w4285_,
		_w4286_,
		_w4287_,
		_w4288_
	);
	LUT4 #(
		.INIT('h0660)
	) name3286 (
		_w4277_,
		_w4278_,
		_w4286_,
		_w4287_,
		_w4289_
	);
	LUT4 #(
		.INIT('h0080)
	) name3287 (
		_w4276_,
		_w4277_,
		_w4278_,
		_w4280_,
		_w4290_
	);
	LUT2 #(
		.INIT('h2)
	) name3288 (
		_w4289_,
		_w4290_,
		_w4291_
	);
	LUT4 #(
		.INIT('h6999)
	) name3289 (
		_w4284_,
		_w4285_,
		_w4286_,
		_w4287_,
		_w4292_
	);
	LUT3 #(
		.INIT('h02)
	) name3290 (
		_w4289_,
		_w4290_,
		_w4292_,
		_w4293_
	);
	LUT3 #(
		.INIT('hd0)
	) name3291 (
		_w4289_,
		_w4290_,
		_w4292_,
		_w4294_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name3292 (
		\A[514] ,
		\A[515] ,
		\A[516] ,
		_w4277_,
		_w4295_
	);
	LUT2 #(
		.INIT('h9)
	) name3293 (
		_w4280_,
		_w4295_,
		_w4296_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3294 (
		_w4288_,
		_w4291_,
		_w4292_,
		_w4296_,
		_w4297_
	);
	LUT4 #(
		.INIT('h1051)
	) name3295 (
		_w4288_,
		_w4291_,
		_w4292_,
		_w4296_,
		_w4298_
	);
	LUT4 #(
		.INIT('h6566)
	) name3296 (
		_w4288_,
		_w4293_,
		_w4294_,
		_w4296_,
		_w4299_
	);
	LUT2 #(
		.INIT('h6)
	) name3297 (
		_w4283_,
		_w4299_,
		_w4300_
	);
	LUT2 #(
		.INIT('h8)
	) name3298 (
		\A[526] ,
		\A[527] ,
		_w4301_
	);
	LUT3 #(
		.INIT('h96)
	) name3299 (
		\A[523] ,
		\A[524] ,
		\A[525] ,
		_w4302_
	);
	LUT3 #(
		.INIT('h96)
	) name3300 (
		\A[526] ,
		\A[527] ,
		\A[528] ,
		_w4303_
	);
	LUT3 #(
		.INIT('h80)
	) name3301 (
		_w4301_,
		_w4302_,
		_w4303_,
		_w4304_
	);
	LUT3 #(
		.INIT('h17)
	) name3302 (
		\A[523] ,
		\A[524] ,
		\A[525] ,
		_w4305_
	);
	LUT3 #(
		.INIT('h17)
	) name3303 (
		\A[526] ,
		\A[527] ,
		\A[528] ,
		_w4306_
	);
	LUT4 #(
		.INIT('h080f)
	) name3304 (
		_w4302_,
		_w4303_,
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT2 #(
		.INIT('h1)
	) name3305 (
		_w4304_,
		_w4307_,
		_w4308_
	);
	LUT3 #(
		.INIT('h17)
	) name3306 (
		\A[532] ,
		\A[533] ,
		\A[534] ,
		_w4309_
	);
	LUT3 #(
		.INIT('h17)
	) name3307 (
		\A[529] ,
		\A[530] ,
		\A[531] ,
		_w4310_
	);
	LUT3 #(
		.INIT('h96)
	) name3308 (
		\A[529] ,
		\A[530] ,
		\A[531] ,
		_w4311_
	);
	LUT3 #(
		.INIT('h96)
	) name3309 (
		\A[532] ,
		\A[533] ,
		\A[534] ,
		_w4312_
	);
	LUT4 #(
		.INIT('h7111)
	) name3310 (
		_w4309_,
		_w4310_,
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT4 #(
		.INIT('h0660)
	) name3311 (
		_w4302_,
		_w4303_,
		_w4311_,
		_w4312_,
		_w4314_
	);
	LUT4 #(
		.INIT('h0080)
	) name3312 (
		_w4301_,
		_w4302_,
		_w4303_,
		_w4305_,
		_w4315_
	);
	LUT2 #(
		.INIT('h2)
	) name3313 (
		_w4314_,
		_w4315_,
		_w4316_
	);
	LUT4 #(
		.INIT('h6999)
	) name3314 (
		_w4309_,
		_w4310_,
		_w4311_,
		_w4312_,
		_w4317_
	);
	LUT3 #(
		.INIT('h02)
	) name3315 (
		_w4314_,
		_w4315_,
		_w4317_,
		_w4318_
	);
	LUT3 #(
		.INIT('hd0)
	) name3316 (
		_w4314_,
		_w4315_,
		_w4317_,
		_w4319_
	);
	LUT4 #(
		.INIT('h7ee8)
	) name3317 (
		\A[526] ,
		\A[527] ,
		\A[528] ,
		_w4302_,
		_w4320_
	);
	LUT2 #(
		.INIT('h9)
	) name3318 (
		_w4305_,
		_w4320_,
		_w4321_
	);
	LUT4 #(
		.INIT('h8a08)
	) name3319 (
		_w4313_,
		_w4316_,
		_w4317_,
		_w4321_,
		_w4322_
	);
	LUT4 #(
		.INIT('h1051)
	) name3320 (
		_w4313_,
		_w4316_,
		_w4317_,
		_w4321_,
		_w4323_
	);
	LUT4 #(
		.INIT('h6566)
	) name3321 (
		_w4313_,
		_w4318_,
		_w4319_,
		_w4321_,
		_w4324_
	);
	LUT2 #(
		.INIT('h6)
	) name3322 (
		_w4308_,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('h9009)
	) name3323 (
		_w4283_,
		_w4299_,
		_w4308_,
		_w4324_,
		_w4326_
	);
	LUT4 #(
		.INIT('h0660)
	) name3324 (
		_w4283_,
		_w4299_,
		_w4308_,
		_w4324_,
		_w4327_
	);
	LUT4 #(
		.INIT('h6996)
	) name3325 (
		_w4302_,
		_w4303_,
		_w4311_,
		_w4312_,
		_w4328_
	);
	LUT4 #(
		.INIT('h6996)
	) name3326 (
		_w4277_,
		_w4278_,
		_w4286_,
		_w4287_,
		_w4329_
	);
	LUT2 #(
		.INIT('h8)
	) name3327 (
		_w4328_,
		_w4329_,
		_w4330_
	);
	LUT3 #(
		.INIT('h2d)
	) name3328 (
		_w4314_,
		_w4315_,
		_w4317_,
		_w4331_
	);
	LUT3 #(
		.INIT('h48)
	) name3329 (
		_w4321_,
		_w4330_,
		_w4331_,
		_w4332_
	);
	LUT3 #(
		.INIT('h21)
	) name3330 (
		_w4321_,
		_w4330_,
		_w4331_,
		_w4333_
	);
	LUT3 #(
		.INIT('h2d)
	) name3331 (
		_w4289_,
		_w4290_,
		_w4292_,
		_w4334_
	);
	LUT2 #(
		.INIT('h6)
	) name3332 (
		_w4296_,
		_w4334_,
		_w4335_
	);
	LUT3 #(
		.INIT('h45)
	) name3333 (
		_w4332_,
		_w4333_,
		_w4335_,
		_w4336_
	);
	LUT3 #(
		.INIT('h32)
	) name3334 (
		_w4308_,
		_w4322_,
		_w4323_,
		_w4337_
	);
	LUT4 #(
		.INIT('h0017)
	) name3335 (
		_w4300_,
		_w4325_,
		_w4336_,
		_w4337_,
		_w4338_
	);
	LUT4 #(
		.INIT('he800)
	) name3336 (
		_w4300_,
		_w4325_,
		_w4336_,
		_w4337_,
		_w4339_
	);
	LUT4 #(
		.INIT('hab54)
	) name3337 (
		_w4326_,
		_w4327_,
		_w4336_,
		_w4337_,
		_w4340_
	);
	LUT3 #(
		.INIT('h32)
	) name3338 (
		_w4283_,
		_w4297_,
		_w4298_,
		_w4341_
	);
	LUT2 #(
		.INIT('h9)
	) name3339 (
		_w4340_,
		_w4341_,
		_w4342_
	);
	LUT4 #(
		.INIT('h0660)
	) name3340 (
		_w4272_,
		_w4274_,
		_w4340_,
		_w4341_,
		_w4343_
	);
	LUT4 #(
		.INIT('h9009)
	) name3341 (
		_w4272_,
		_w4274_,
		_w4340_,
		_w4341_,
		_w4344_
	);
	LUT4 #(
		.INIT('h6996)
	) name3342 (
		_w4283_,
		_w4299_,
		_w4308_,
		_w4324_,
		_w4345_
	);
	LUT4 #(
		.INIT('h6996)
	) name3343 (
		_w4215_,
		_w4231_,
		_w4240_,
		_w4256_,
		_w4346_
	);
	LUT4 #(
		.INIT('h1428)
	) name3344 (
		_w4268_,
		_w4336_,
		_w4345_,
		_w4346_,
		_w4347_
	);
	LUT4 #(
		.INIT('h8241)
	) name3345 (
		_w4268_,
		_w4336_,
		_w4345_,
		_w4346_,
		_w4348_
	);
	LUT4 #(
		.INIT('h0660)
	) name3346 (
		_w4260_,
		_w4261_,
		_w4328_,
		_w4329_,
		_w4349_
	);
	LUT3 #(
		.INIT('h96)
	) name3347 (
		_w4253_,
		_w4262_,
		_w4263_,
		_w4350_
	);
	LUT3 #(
		.INIT('h48)
	) name3348 (
		_w4267_,
		_w4349_,
		_w4350_,
		_w4351_
	);
	LUT3 #(
		.INIT('h21)
	) name3349 (
		_w4267_,
		_w4349_,
		_w4350_,
		_w4352_
	);
	LUT3 #(
		.INIT('h96)
	) name3350 (
		_w4321_,
		_w4330_,
		_w4331_,
		_w4353_
	);
	LUT2 #(
		.INIT('h9)
	) name3351 (
		_w4335_,
		_w4353_,
		_w4354_
	);
	LUT3 #(
		.INIT('h54)
	) name3352 (
		_w4351_,
		_w4352_,
		_w4354_,
		_w4355_
	);
	LUT3 #(
		.INIT('h45)
	) name3353 (
		_w4347_,
		_w4348_,
		_w4355_,
		_w4356_
	);
	LUT4 #(
		.INIT('h022a)
	) name3354 (
		_w4273_,
		_w4275_,
		_w4342_,
		_w4356_,
		_w4357_
	);
	LUT4 #(
		.INIT('h5440)
	) name3355 (
		_w4273_,
		_w4275_,
		_w4342_,
		_w4356_,
		_w4358_
	);
	LUT4 #(
		.INIT('h6665)
	) name3356 (
		_w4273_,
		_w4343_,
		_w4344_,
		_w4356_,
		_w4359_
	);
	LUT3 #(
		.INIT('h54)
	) name3357 (
		_w4338_,
		_w4339_,
		_w4341_,
		_w4360_
	);
	LUT2 #(
		.INIT('h6)
	) name3358 (
		_w4359_,
		_w4360_,
		_w4361_
	);
	LUT4 #(
		.INIT('h9009)
	) name3359 (
		_w4205_,
		_w4206_,
		_w4359_,
		_w4360_,
		_w4362_
	);
	LUT4 #(
		.INIT('h0660)
	) name3360 (
		_w4205_,
		_w4206_,
		_w4359_,
		_w4360_,
		_w4363_
	);
	LUT4 #(
		.INIT('h6996)
	) name3361 (
		_w4272_,
		_w4274_,
		_w4340_,
		_w4341_,
		_w4364_
	);
	LUT4 #(
		.INIT('h6996)
	) name3362 (
		_w4118_,
		_w4184_,
		_w4185_,
		_w4187_,
		_w4365_
	);
	LUT4 #(
		.INIT('h1428)
	) name3363 (
		_w4202_,
		_w4356_,
		_w4364_,
		_w4365_,
		_w4366_
	);
	LUT4 #(
		.INIT('h8241)
	) name3364 (
		_w4202_,
		_w4356_,
		_w4364_,
		_w4365_,
		_w4367_
	);
	LUT4 #(
		.INIT('h6996)
	) name3365 (
		_w4114_,
		_w4180_,
		_w4191_,
		_w4192_,
		_w4368_
	);
	LUT4 #(
		.INIT('h6996)
	) name3366 (
		_w4268_,
		_w4336_,
		_w4345_,
		_w4346_,
		_w4369_
	);
	LUT4 #(
		.INIT('h1248)
	) name3367 (
		_w4201_,
		_w4355_,
		_w4368_,
		_w4369_,
		_w4370_
	);
	LUT4 #(
		.INIT('h8421)
	) name3368 (
		_w4201_,
		_w4355_,
		_w4368_,
		_w4369_,
		_w4371_
	);
	LUT4 #(
		.INIT('h6996)
	) name3369 (
		_w4106_,
		_w4107_,
		_w4172_,
		_w4173_,
		_w4372_
	);
	LUT4 #(
		.INIT('h6996)
	) name3370 (
		_w4260_,
		_w4261_,
		_w4328_,
		_w4329_,
		_w4373_
	);
	LUT2 #(
		.INIT('h8)
	) name3371 (
		_w4372_,
		_w4373_,
		_w4374_
	);
	LUT3 #(
		.INIT('h96)
	) name3372 (
		_w4267_,
		_w4349_,
		_w4350_,
		_w4375_
	);
	LUT3 #(
		.INIT('h84)
	) name3373 (
		_w4354_,
		_w4374_,
		_w4375_,
		_w4376_
	);
	LUT3 #(
		.INIT('h12)
	) name3374 (
		_w4354_,
		_w4374_,
		_w4375_,
		_w4377_
	);
	LUT3 #(
		.INIT('h96)
	) name3375 (
		_w4179_,
		_w4195_,
		_w4196_,
		_w4378_
	);
	LUT2 #(
		.INIT('h9)
	) name3376 (
		_w4200_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('h45)
	) name3377 (
		_w4376_,
		_w4377_,
		_w4379_,
		_w4380_
	);
	LUT3 #(
		.INIT('h45)
	) name3378 (
		_w4370_,
		_w4371_,
		_w4380_,
		_w4381_
	);
	LUT3 #(
		.INIT('h45)
	) name3379 (
		_w4366_,
		_w4367_,
		_w4381_,
		_w4382_
	);
	LUT3 #(
		.INIT('h45)
	) name3380 (
		_w4203_,
		_w4204_,
		_w4206_,
		_w4383_
	);
	LUT4 #(
		.INIT('h00e8)
	) name3381 (
		_w4207_,
		_w4361_,
		_w4382_,
		_w4383_,
		_w4384_
	);
	LUT4 #(
		.INIT('h1700)
	) name3382 (
		_w4207_,
		_w4361_,
		_w4382_,
		_w4383_,
		_w4385_
	);
	LUT3 #(
		.INIT('h45)
	) name3383 (
		_w4357_,
		_w4358_,
		_w4360_,
		_w4386_
	);
	LUT3 #(
		.INIT('h54)
	) name3384 (
		_w4384_,
		_w4385_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h8)
	) name3385 (
		_w4052_,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w4052_,
		_w4387_,
		_w4389_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3387 (
		_w4027_,
		_w4028_,
		_w4047_,
		_w4048_,
		_w4390_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3388 (
		_w4362_,
		_w4363_,
		_w4382_,
		_w4383_,
		_w4391_
	);
	LUT4 #(
		.INIT('h1248)
	) name3389 (
		_w4051_,
		_w4386_,
		_w4390_,
		_w4391_,
		_w4392_
	);
	LUT4 #(
		.INIT('h8421)
	) name3390 (
		_w4051_,
		_w4386_,
		_w4390_,
		_w4391_,
		_w4393_
	);
	LUT4 #(
		.INIT('h6996)
	) name3391 (
		_w4205_,
		_w4206_,
		_w4359_,
		_w4360_,
		_w4394_
	);
	LUT4 #(
		.INIT('h6996)
	) name3392 (
		_w3870_,
		_w3871_,
		_w4024_,
		_w4025_,
		_w4395_
	);
	LUT4 #(
		.INIT('h1428)
	) name3393 (
		_w4047_,
		_w4382_,
		_w4394_,
		_w4395_,
		_w4396_
	);
	LUT4 #(
		.INIT('h8241)
	) name3394 (
		_w4047_,
		_w4382_,
		_w4394_,
		_w4395_,
		_w4397_
	);
	LUT4 #(
		.INIT('h6996)
	) name3395 (
		_w3867_,
		_w4021_,
		_w4029_,
		_w4030_,
		_w4398_
	);
	LUT4 #(
		.INIT('h6996)
	) name3396 (
		_w4202_,
		_w4356_,
		_w4364_,
		_w4365_,
		_w4399_
	);
	LUT4 #(
		.INIT('h8421)
	) name3397 (
		_w4046_,
		_w4381_,
		_w4398_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('h1248)
	) name3398 (
		_w4046_,
		_w4381_,
		_w4398_,
		_w4399_,
		_w4401_
	);
	LUT4 #(
		.INIT('h6996)
	) name3399 (
		_w4201_,
		_w4355_,
		_w4368_,
		_w4369_,
		_w4402_
	);
	LUT4 #(
		.INIT('h6996)
	) name3400 (
		_w3866_,
		_w4020_,
		_w4033_,
		_w4034_,
		_w4403_
	);
	LUT4 #(
		.INIT('h1428)
	) name3401 (
		_w4045_,
		_w4380_,
		_w4402_,
		_w4403_,
		_w4404_
	);
	LUT4 #(
		.INIT('h8241)
	) name3402 (
		_w4045_,
		_w4380_,
		_w4402_,
		_w4403_,
		_w4405_
	);
	LUT4 #(
		.INIT('h0660)
	) name3403 (
		_w4037_,
		_w4038_,
		_w4372_,
		_w4373_,
		_w4406_
	);
	LUT3 #(
		.INIT('h69)
	) name3404 (
		_w4019_,
		_w4039_,
		_w4040_,
		_w4407_
	);
	LUT3 #(
		.INIT('h48)
	) name3405 (
		_w4044_,
		_w4406_,
		_w4407_,
		_w4408_
	);
	LUT3 #(
		.INIT('h21)
	) name3406 (
		_w4044_,
		_w4406_,
		_w4407_,
		_w4409_
	);
	LUT3 #(
		.INIT('h69)
	) name3407 (
		_w4354_,
		_w4374_,
		_w4375_,
		_w4410_
	);
	LUT2 #(
		.INIT('h9)
	) name3408 (
		_w4379_,
		_w4410_,
		_w4411_
	);
	LUT3 #(
		.INIT('h54)
	) name3409 (
		_w4408_,
		_w4409_,
		_w4411_,
		_w4412_
	);
	LUT3 #(
		.INIT('h45)
	) name3410 (
		_w4404_,
		_w4405_,
		_w4412_,
		_w4413_
	);
	LUT3 #(
		.INIT('h54)
	) name3411 (
		_w4400_,
		_w4401_,
		_w4413_,
		_w4414_
	);
	LUT3 #(
		.INIT('h54)
	) name3412 (
		_w4396_,
		_w4397_,
		_w4414_,
		_w4415_
	);
	LUT3 #(
		.INIT('h45)
	) name3413 (
		_w4392_,
		_w4393_,
		_w4415_,
		_w4416_
	);
	LUT4 #(
		.INIT('h4054)
	) name3414 (
		_w3718_,
		_w4052_,
		_w4387_,
		_w4416_,
		_w4417_
	);
	LUT4 #(
		.INIT('h2a02)
	) name3415 (
		_w3718_,
		_w4052_,
		_w4387_,
		_w4416_,
		_w4418_
	);
	LUT2 #(
		.INIT('h6)
	) name3416 (
		_w4052_,
		_w4387_,
		_w4419_
	);
	LUT2 #(
		.INIT('h6)
	) name3417 (
		_w3398_,
		_w3696_,
		_w4420_
	);
	LUT2 #(
		.INIT('h9)
	) name3418 (
		_w3717_,
		_w4420_,
		_w4421_
	);
	LUT4 #(
		.INIT('h6996)
	) name3419 (
		_w3397_,
		_w3695_,
		_w3699_,
		_w3700_,
		_w4422_
	);
	LUT2 #(
		.INIT('h9)
	) name3420 (
		_w3716_,
		_w4422_,
		_w4423_
	);
	LUT4 #(
		.INIT('h6996)
	) name3421 (
		_w4051_,
		_w4386_,
		_w4390_,
		_w4391_,
		_w4424_
	);
	LUT4 #(
		.INIT('h6996)
	) name3422 (
		_w4047_,
		_w4382_,
		_w4394_,
		_w4395_,
		_w4425_
	);
	LUT3 #(
		.INIT('h96)
	) name3423 (
		_w3703_,
		_w3704_,
		_w3715_,
		_w4426_
	);
	LUT3 #(
		.INIT('h96)
	) name3424 (
		_w3705_,
		_w3706_,
		_w3714_,
		_w4427_
	);
	LUT4 #(
		.INIT('h6996)
	) name3425 (
		_w4046_,
		_w4381_,
		_w4398_,
		_w4399_,
		_w4428_
	);
	LUT4 #(
		.INIT('h6996)
	) name3426 (
		_w4045_,
		_w4380_,
		_w4402_,
		_w4403_,
		_w4429_
	);
	LUT3 #(
		.INIT('h69)
	) name3427 (
		_w3707_,
		_w3708_,
		_w3713_,
		_w4430_
	);
	LUT4 #(
		.INIT('h6996)
	) name3428 (
		_w4037_,
		_w4038_,
		_w4372_,
		_w4373_,
		_w4431_
	);
	LUT4 #(
		.INIT('h6996)
	) name3429 (
		_w3389_,
		_w3390_,
		_w3687_,
		_w3688_,
		_w4432_
	);
	LUT2 #(
		.INIT('h8)
	) name3430 (
		_w4431_,
		_w4432_,
		_w4433_
	);
	LUT4 #(
		.INIT('h6996)
	) name3431 (
		_w3391_,
		_w3392_,
		_w3393_,
		_w3709_,
		_w4434_
	);
	LUT3 #(
		.INIT('h84)
	) name3432 (
		_w3712_,
		_w4433_,
		_w4434_,
		_w4435_
	);
	LUT3 #(
		.INIT('h12)
	) name3433 (
		_w3712_,
		_w4433_,
		_w4434_,
		_w4436_
	);
	LUT3 #(
		.INIT('h96)
	) name3434 (
		_w4044_,
		_w4406_,
		_w4407_,
		_w4437_
	);
	LUT4 #(
		.INIT('h3132)
	) name3435 (
		_w4411_,
		_w4435_,
		_w4436_,
		_w4437_,
		_w4438_
	);
	LUT4 #(
		.INIT('h90f9)
	) name3436 (
		_w4412_,
		_w4429_,
		_w4430_,
		_w4438_,
		_w4439_
	);
	LUT4 #(
		.INIT('h84ed)
	) name3437 (
		_w4413_,
		_w4427_,
		_w4428_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('hf990)
	) name3438 (
		_w4414_,
		_w4425_,
		_w4426_,
		_w4440_,
		_w4441_
	);
	LUT4 #(
		.INIT('hed84)
	) name3439 (
		_w4415_,
		_w4423_,
		_w4424_,
		_w4441_,
		_w4442_
	);
	LUT4 #(
		.INIT('hf660)
	) name3440 (
		_w4416_,
		_w4419_,
		_w4421_,
		_w4442_,
		_w4443_
	);
	LUT3 #(
		.INIT('h54)
	) name3441 (
		_w4417_,
		_w4418_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h8)
	) name3442 (
		_w3126_,
		_w4444_,
		_w4445_
	);
	LUT3 #(
		.INIT('h69)
	) name3443 (
		_w3086_,
		_w3091_,
		_w3092_,
		_w4446_
	);
	LUT4 #(
		.INIT('h999a)
	) name3444 (
		_w3718_,
		_w4388_,
		_w4389_,
		_w4416_,
		_w4447_
	);
	LUT2 #(
		.INIT('h9)
	) name3445 (
		_w4443_,
		_w4447_,
		_w4448_
	);
	LUT3 #(
		.INIT('h96)
	) name3446 (
		_w3085_,
		_w3097_,
		_w3098_,
		_w4449_
	);
	LUT4 #(
		.INIT('h9669)
	) name3447 (
		_w4416_,
		_w4419_,
		_w4421_,
		_w4442_,
		_w4450_
	);
	LUT3 #(
		.INIT('h96)
	) name3448 (
		_w3084_,
		_w3101_,
		_w3102_,
		_w4451_
	);
	LUT4 #(
		.INIT('h6996)
	) name3449 (
		_w4415_,
		_w4423_,
		_w4424_,
		_w4441_,
		_w4452_
	);
	LUT3 #(
		.INIT('h96)
	) name3450 (
		_w3083_,
		_w3105_,
		_w3106_,
		_w4453_
	);
	LUT4 #(
		.INIT('h6996)
	) name3451 (
		_w4414_,
		_w4425_,
		_w4426_,
		_w4440_,
		_w4454_
	);
	LUT3 #(
		.INIT('h69)
	) name3452 (
		_w3082_,
		_w3109_,
		_w3110_,
		_w4455_
	);
	LUT4 #(
		.INIT('h9669)
	) name3453 (
		_w4413_,
		_w4427_,
		_w4428_,
		_w4439_,
		_w4456_
	);
	LUT4 #(
		.INIT('h9669)
	) name3454 (
		_w3074_,
		_w3075_,
		_w3081_,
		_w3113_,
		_w4457_
	);
	LUT4 #(
		.INIT('h6996)
	) name3455 (
		_w4412_,
		_w4429_,
		_w4430_,
		_w4438_,
		_w4458_
	);
	LUT2 #(
		.INIT('h6)
	) name3456 (
		_w4431_,
		_w4432_,
		_w4459_
	);
	LUT4 #(
		.INIT('h6996)
	) name3457 (
		_w1757_,
		_w1758_,
		_w3076_,
		_w3077_,
		_w4460_
	);
	LUT2 #(
		.INIT('h8)
	) name3458 (
		_w4459_,
		_w4460_,
		_w4461_
	);
	LUT4 #(
		.INIT('h0096)
	) name3459 (
		_w3116_,
		_w3117_,
		_w3119_,
		_w4461_,
		_w4462_
	);
	LUT4 #(
		.INIT('h6900)
	) name3460 (
		_w3116_,
		_w3117_,
		_w3119_,
		_w4461_,
		_w4463_
	);
	LUT3 #(
		.INIT('h69)
	) name3461 (
		_w3712_,
		_w4433_,
		_w4434_,
		_w4464_
	);
	LUT3 #(
		.INIT('h96)
	) name3462 (
		_w4411_,
		_w4437_,
		_w4464_,
		_w4465_
	);
	LUT3 #(
		.INIT('h45)
	) name3463 (
		_w4462_,
		_w4463_,
		_w4465_,
		_w4466_
	);
	LUT4 #(
		.INIT('h066f)
	) name3464 (
		_w3120_,
		_w4457_,
		_w4458_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('h60f6)
	) name3465 (
		_w3121_,
		_w4455_,
		_w4456_,
		_w4467_,
		_w4468_
	);
	LUT4 #(
		.INIT('hf990)
	) name3466 (
		_w3122_,
		_w4453_,
		_w4454_,
		_w4468_,
		_w4469_
	);
	LUT4 #(
		.INIT('h099f)
	) name3467 (
		_w3123_,
		_w4451_,
		_w4452_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('h60f6)
	) name3468 (
		_w3124_,
		_w4449_,
		_w4450_,
		_w4470_,
		_w4471_
	);
	LUT4 #(
		.INIT('hf660)
	) name3469 (
		_w3125_,
		_w4446_,
		_w4448_,
		_w4471_,
		_w4472_
	);
	LUT4 #(
		.INIT('h9669)
	) name3470 (
		_w3125_,
		_w4446_,
		_w4448_,
		_w4471_,
		_w4473_
	);
	LUT4 #(
		.INIT('h0096)
	) name3471 (
		_w3124_,
		_w4449_,
		_w4450_,
		_w4470_,
		_w4474_
	);
	LUT4 #(
		.INIT('h6900)
	) name3472 (
		_w3124_,
		_w4449_,
		_w4450_,
		_w4470_,
		_w4475_
	);
	LUT4 #(
		.INIT('h0069)
	) name3473 (
		_w3123_,
		_w4451_,
		_w4452_,
		_w4469_,
		_w4476_
	);
	LUT4 #(
		.INIT('h9600)
	) name3474 (
		_w3123_,
		_w4451_,
		_w4452_,
		_w4469_,
		_w4477_
	);
	LUT4 #(
		.INIT('h6996)
	) name3475 (
		_w3122_,
		_w4453_,
		_w4454_,
		_w4468_,
		_w4478_
	);
	LUT4 #(
		.INIT('h9600)
	) name3476 (
		_w3121_,
		_w4455_,
		_w4456_,
		_w4467_,
		_w4479_
	);
	LUT4 #(
		.INIT('h6900)
	) name3477 (
		_w3120_,
		_w4457_,
		_w4458_,
		_w4466_,
		_w4480_
	);
	LUT4 #(
		.INIT('h0096)
	) name3478 (
		_w3120_,
		_w4457_,
		_w4458_,
		_w4466_,
		_w4481_
	);
	LUT3 #(
		.INIT('h41)
	) name3479 (
		\A[1000] ,
		_w4459_,
		_w4460_,
		_w4482_
	);
	LUT4 #(
		.INIT('he100)
	) name3480 (
		_w4462_,
		_w4463_,
		_w4465_,
		_w4482_,
		_w4483_
	);
	LUT3 #(
		.INIT('h01)
	) name3481 (
		_w4481_,
		_w4483_,
		_w4480_,
		_w4484_
	);
	LUT4 #(
		.INIT('h0069)
	) name3482 (
		_w3121_,
		_w4455_,
		_w4456_,
		_w4467_,
		_w4485_
	);
	LUT3 #(
		.INIT('h01)
	) name3483 (
		_w4484_,
		_w4485_,
		_w4479_,
		_w4486_
	);
	LUT2 #(
		.INIT('h1)
	) name3484 (
		_w4478_,
		_w4486_,
		_w4487_
	);
	LUT3 #(
		.INIT('h10)
	) name3485 (
		_w4477_,
		_w4476_,
		_w4487_,
		_w4488_
	);
	LUT3 #(
		.INIT('h10)
	) name3486 (
		_w4475_,
		_w4474_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h4)
	) name3487 (
		_w4473_,
		_w4489_,
		_w4490_
	);
	LUT4 #(
		.INIT('h1501)
	) name3488 (
		_w3087_,
		_w3091_,
		_w3093_,
		_w3125_,
		_w4491_
	);
	LUT4 #(
		.INIT('h0054)
	) name3489 (
		_w3088_,
		_w3126_,
		_w4444_,
		_w4491_,
		_w4492_
	);
	LUT4 #(
		.INIT('hd4ff)
	) name3490 (
		_w4445_,
		_w4472_,
		_w4490_,
		_w4492_,
		_w4493_
	);
	assign maj = _w4493_ ;
endmodule;