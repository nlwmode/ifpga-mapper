module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  output q_pad ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n17 = ~b_pad & ~c_pad ;
  assign n18 = b_pad & c_pad ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = a_pad & ~d_pad ;
  assign n21 = ~a_pad & d_pad ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = ~n19 & ~n22 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = e_pad & ~f_pad ;
  assign n27 = ~e_pad & f_pad ;
  assign n28 = ~n26 & ~n27 ;
  assign n29 = g_pad & ~h_pad ;
  assign n30 = ~g_pad & h_pad ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = ~n28 & n31 ;
  assign n34 = ~n32 & ~n33 ;
  assign n35 = n25 & n34 ;
  assign n36 = ~n25 & ~n34 ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = ~j_pad & ~k_pad ;
  assign n39 = j_pad & k_pad ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = i_pad & ~l_pad ;
  assign n42 = ~i_pad & l_pad ;
  assign n43 = ~n41 & ~n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = ~n40 & ~n43 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = m_pad & ~n_pad ;
  assign n48 = ~m_pad & n_pad ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = o_pad & ~p_pad ;
  assign n51 = ~o_pad & p_pad ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = n49 & ~n52 ;
  assign n54 = ~n49 & n52 ;
  assign n55 = ~n53 & ~n54 ;
  assign n56 = n46 & ~n55 ;
  assign n57 = ~n46 & n55 ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = n37 & n58 ;
  assign n60 = ~n37 & ~n58 ;
  assign n61 = ~n59 & ~n60 ;
  assign q_pad = ~n61 ;
endmodule
