module top( \C3_Q0_reg/NET0131  , \C3_Q1_reg/NET0131  , \C3_Q2_reg/NET0131  , \C3_Q3_reg/NET0131  , CLR_pad , \FML_reg/NET0131  , FM_pad , \OLATCHVUC_5_reg/NET0131  , \OLATCHVUC_6_reg/NET0131  , \OLATCH_FEL_reg/NET0131  , \TESTL_reg/NET0131  , TEST_pad , \UC_10_reg/NET0131  , \UC_11_reg/NET0131  , \UC_16_reg/NET0131  , \UC_17_reg/NET0131  , \UC_18_reg/NET0131  , \UC_19_reg/NET0131  , \UC_8_reg/NET0131  , \UC_9_reg/NET0131  , \RED2_pad  , \YLW1_pad  , \_al_n0  , \_al_n1  , \g19/_0_  , \g28/_2_  , \g706/_0_  , \g726/_0_  , \g727/_0_  , \g738/_0_  , \g740/_0_  , \g747/_0_  , \g755/_0_  , \g759/_0_  , \g762/_0_  , \g765/_0_  , \g768/_0_  , \g776/_0_  , \g778/_0_  , \g780/_0_  , \g781/_0_  , \g787/_0_  , \g909/_0_  , \g928/_2_  , \g978/_1_  );
  input \C3_Q0_reg/NET0131  ;
  input \C3_Q1_reg/NET0131  ;
  input \C3_Q2_reg/NET0131  ;
  input \C3_Q3_reg/NET0131  ;
  input CLR_pad ;
  input \FML_reg/NET0131  ;
  input FM_pad ;
  input \OLATCHVUC_5_reg/NET0131  ;
  input \OLATCHVUC_6_reg/NET0131  ;
  input \OLATCH_FEL_reg/NET0131  ;
  input \TESTL_reg/NET0131  ;
  input TEST_pad ;
  input \UC_10_reg/NET0131  ;
  input \UC_11_reg/NET0131  ;
  input \UC_16_reg/NET0131  ;
  input \UC_17_reg/NET0131  ;
  input \UC_18_reg/NET0131  ;
  input \UC_19_reg/NET0131  ;
  input \UC_8_reg/NET0131  ;
  input \UC_9_reg/NET0131  ;
  output \RED2_pad  ;
  output \YLW1_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g19/_0_  ;
  output \g28/_2_  ;
  output \g706/_0_  ;
  output \g726/_0_  ;
  output \g727/_0_  ;
  output \g738/_0_  ;
  output \g740/_0_  ;
  output \g747/_0_  ;
  output \g755/_0_  ;
  output \g759/_0_  ;
  output \g762/_0_  ;
  output \g765/_0_  ;
  output \g768/_0_  ;
  output \g776/_0_  ;
  output \g778/_0_  ;
  output \g780/_0_  ;
  output \g781/_0_  ;
  output \g787/_0_  ;
  output \g909/_0_  ;
  output \g928/_2_  ;
  output \g978/_1_  ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 ;
  assign n21 = ~\UC_10_reg/NET0131  & ~\UC_11_reg/NET0131  ;
  assign n22 = ~\UC_9_reg/NET0131  & n21 ;
  assign n23 = \UC_8_reg/NET0131  & ~n22 ;
  assign n24 = ~\TESTL_reg/NET0131  & ~n23 ;
  assign n30 = \UC_18_reg/NET0131  & \UC_19_reg/NET0131  ;
  assign n31 = ~n24 & n30 ;
  assign n32 = \UC_17_reg/NET0131  & n31 ;
  assign n34 = \UC_16_reg/NET0131  & n32 ;
  assign n25 = ~\UC_17_reg/NET0131  & ~\UC_18_reg/NET0131  ;
  assign n26 = ~\UC_19_reg/NET0131  & n25 ;
  assign n27 = \UC_16_reg/NET0131  & ~n26 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = ~CLR_pad & ~n28 ;
  assign n33 = ~\UC_16_reg/NET0131  & ~n32 ;
  assign n35 = n29 & ~n33 ;
  assign n36 = ~n34 & n35 ;
  assign n42 = \C3_Q0_reg/NET0131  & \C3_Q1_reg/NET0131  ;
  assign n43 = n28 & n42 ;
  assign n45 = \C3_Q2_reg/NET0131  & n43 ;
  assign n37 = ~\C3_Q0_reg/NET0131  & ~\C3_Q1_reg/NET0131  ;
  assign n38 = ~\C3_Q2_reg/NET0131  & n37 ;
  assign n39 = \C3_Q3_reg/NET0131  & ~n38 ;
  assign n40 = n28 & n39 ;
  assign n41 = ~CLR_pad & ~n40 ;
  assign n44 = ~\C3_Q2_reg/NET0131  & ~n43 ;
  assign n46 = n41 & ~n44 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~\UC_17_reg/NET0131  & ~n31 ;
  assign n49 = n29 & ~n32 ;
  assign n50 = ~n48 & n49 ;
  assign n51 = \UC_19_reg/NET0131  & ~n24 ;
  assign n52 = ~\UC_18_reg/NET0131  & ~n51 ;
  assign n53 = n29 & ~n31 ;
  assign n54 = ~n52 & n53 ;
  assign n55 = ~\UC_19_reg/NET0131  & n24 ;
  assign n56 = ~n51 & ~n55 ;
  assign n57 = n29 & n56 ;
  assign n58 = \C3_Q2_reg/NET0131  & ~CLR_pad ;
  assign n59 = \FML_reg/NET0131  & n37 ;
  assign n60 = n58 & n59 ;
  assign n61 = \C3_Q0_reg/NET0131  & ~\C3_Q1_reg/NET0131  ;
  assign n62 = ~\C3_Q3_reg/NET0131  & ~\FML_reg/NET0131  ;
  assign n63 = n61 & n62 ;
  assign n64 = \C3_Q2_reg/NET0131  & n63 ;
  assign n65 = ~CLR_pad & \OLATCH_FEL_reg/NET0131  ;
  assign n66 = ~n64 & n65 ;
  assign n67 = ~n60 & ~n66 ;
  assign n68 = \UC_17_reg/NET0131  & ~n67 ;
  assign n69 = ~\C3_Q2_reg/NET0131  & ~\OLATCH_FEL_reg/NET0131  ;
  assign n70 = \C3_Q3_reg/NET0131  & n37 ;
  assign n71 = n69 & ~n70 ;
  assign n72 = ~CLR_pad & ~n71 ;
  assign n73 = ~n68 & n72 ;
  assign n75 = ~\C3_Q3_reg/NET0131  & \FML_reg/NET0131  ;
  assign n76 = \C3_Q2_reg/NET0131  & ~n75 ;
  assign n74 = ~\C3_Q2_reg/NET0131  & ~\C3_Q3_reg/NET0131  ;
  assign n77 = ~CLR_pad & n37 ;
  assign n78 = ~n74 & n77 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = ~n66 & ~n79 ;
  assign n81 = ~n68 & ~n80 ;
  assign n83 = \OLATCH_FEL_reg/NET0131  & ~n63 ;
  assign n82 = \C3_Q3_reg/NET0131  & \FML_reg/NET0131  ;
  assign n84 = n58 & ~n82 ;
  assign n85 = ~n59 & n84 ;
  assign n86 = ~n83 & n85 ;
  assign n87 = ~CLR_pad & ~n23 ;
  assign n88 = \UC_10_reg/NET0131  & \UC_11_reg/NET0131  ;
  assign n89 = \UC_9_reg/NET0131  & n88 ;
  assign n90 = ~\UC_8_reg/NET0131  & ~n89 ;
  assign n91 = \UC_8_reg/NET0131  & n89 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = n87 & n92 ;
  assign n94 = ~\UC_9_reg/NET0131  & ~n88 ;
  assign n95 = ~n89 & ~n94 ;
  assign n96 = n87 & n95 ;
  assign n97 = ~n21 & ~n88 ;
  assign n98 = n87 & n97 ;
  assign n99 = ~\C3_Q0_reg/NET0131  & \C3_Q3_reg/NET0131  ;
  assign n100 = ~n42 & n69 ;
  assign n101 = ~n99 & n100 ;
  assign n102 = ~CLR_pad & ~n101 ;
  assign n103 = ~\UC_11_reg/NET0131  & n87 ;
  assign n104 = \C3_Q3_reg/NET0131  & ~n61 ;
  assign n105 = n69 & ~n104 ;
  assign n106 = ~CLR_pad & ~n105 ;
  assign n107 = \FML_reg/NET0131  & ~FM_pad ;
  assign n108 = ~\FML_reg/NET0131  & FM_pad ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = ~CLR_pad & ~n109 ;
  assign n111 = \TESTL_reg/NET0131  & ~TEST_pad ;
  assign n112 = ~\TESTL_reg/NET0131  & TEST_pad ;
  assign n113 = ~n111 & ~n112 ;
  assign n114 = ~CLR_pad & ~n113 ;
  assign n115 = ~CLR_pad & n42 ;
  assign n116 = n69 & n115 ;
  assign n117 = \C3_Q0_reg/NET0131  & n28 ;
  assign n118 = ~\C3_Q1_reg/NET0131  & ~n117 ;
  assign n119 = n41 & ~n43 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = ~\C3_Q0_reg/NET0131  & ~n28 ;
  assign n122 = ~n117 & ~n121 ;
  assign n123 = n41 & n122 ;
  assign n124 = ~\C3_Q3_reg/NET0131  & ~n45 ;
  assign n125 = n41 & ~n124 ;
  assign \RED2_pad  = ~\OLATCHVUC_5_reg/NET0131  ;
  assign \YLW1_pad  = ~\OLATCHVUC_6_reg/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g19/_0_  = n36 ;
  assign \g28/_2_  = n47 ;
  assign \g706/_0_  = n50 ;
  assign \g726/_0_  = n54 ;
  assign \g727/_0_  = n57 ;
  assign \g738/_0_  = ~n73 ;
  assign \g740/_0_  = ~n81 ;
  assign \g747/_0_  = n86 ;
  assign \g755/_0_  = ~n67 ;
  assign \g759/_0_  = n93 ;
  assign \g762/_0_  = n96 ;
  assign \g765/_0_  = n98 ;
  assign \g768/_0_  = ~n102 ;
  assign \g776/_0_  = n103 ;
  assign \g778/_0_  = ~n106 ;
  assign \g780/_0_  = n110 ;
  assign \g781/_0_  = n114 ;
  assign \g787/_0_  = n116 ;
  assign \g909/_0_  = n120 ;
  assign \g928/_2_  = n123 ;
  assign \g978/_1_  = n125 ;
endmodule
