module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  output e_pad ;
  output f_pad ;
  output g_pad ;
  output h_pad ;
  output i_pad ;
  output j_pad ;
  output k_pad ;
  output l_pad ;
  output m_pad ;
  output n_pad ;
  wire n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n5 = ~c_pad & ~d_pad ;
  assign n6 = ~a_pad & ~b_pad ;
  assign n7 = n5 & n6 ;
  assign n8 = a_pad & ~b_pad ;
  assign n9 = n5 & n8 ;
  assign n10 = ~a_pad & b_pad ;
  assign n11 = n5 & n10 ;
  assign n12 = a_pad & b_pad ;
  assign n13 = n5 & n12 ;
  assign n14 = c_pad & ~d_pad ;
  assign n15 = n6 & n14 ;
  assign n16 = n8 & n14 ;
  assign n17 = n10 & n14 ;
  assign n18 = n12 & n14 ;
  assign n19 = ~b_pad & ~c_pad ;
  assign n20 = ~a_pad & d_pad ;
  assign n21 = n19 & n20 ;
  assign n22 = a_pad & d_pad ;
  assign n23 = n19 & n22 ;
  assign e_pad = ~n7 ;
  assign f_pad = ~n9 ;
  assign g_pad = ~n11 ;
  assign h_pad = ~n13 ;
  assign i_pad = ~n15 ;
  assign j_pad = ~n16 ;
  assign k_pad = ~n17 ;
  assign l_pad = ~n18 ;
  assign m_pad = ~n21 ;
  assign n_pad = ~n23 ;
endmodule
