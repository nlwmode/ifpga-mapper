module top( \G0_pad  , \G11_reg/NET0131  , \G12_reg/NET0131  , \G13_reg/NET0131  , \G14_reg/NET0131  , \G15_reg/NET0131  , \G16_reg/NET0131  , \G17_reg/NET0131  , \G18_reg/NET0131  , \G19_reg/NET0131  , \G1_pad  , \G20_reg/NET0131  , \G21_reg/NET0131  , \G22_reg/NET0131  , \G23_reg/NET0131  , \G24_reg/NET0131  , \G28_reg/NET0131  , \G29_reg/NET0131  , \G2_pad  , \G31_reg/NET0131  , \G119_pad  , \G167_pad  , \_al_n0  , \_al_n1  , \g43/_3_  , \g754/_0_  , \g757/_0_  , \g760/_0_  , \g768/_2_  , \g770/_2_  , \g773/_0_  , \g786/_2_  , \g792/_0_  , \g793/_0_  , \g796/_0_  , \g804/_0_  , \g808/_0_  , \g817/_0_  , \g825/_0_  , \g834/_0_  , \g837/_0_  , \g838/_0_  , \g839/_0_  , \g840/_0_  , \g843/_0_  );
  input \G0_pad  ;
  input \G11_reg/NET0131  ;
  input \G12_reg/NET0131  ;
  input \G13_reg/NET0131  ;
  input \G14_reg/NET0131  ;
  input \G15_reg/NET0131  ;
  input \G16_reg/NET0131  ;
  input \G17_reg/NET0131  ;
  input \G18_reg/NET0131  ;
  input \G19_reg/NET0131  ;
  input \G1_pad  ;
  input \G20_reg/NET0131  ;
  input \G21_reg/NET0131  ;
  input \G22_reg/NET0131  ;
  input \G23_reg/NET0131  ;
  input \G24_reg/NET0131  ;
  input \G28_reg/NET0131  ;
  input \G29_reg/NET0131  ;
  input \G2_pad  ;
  input \G31_reg/NET0131  ;
  output \G119_pad  ;
  output \G167_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g43/_3_  ;
  output \g754/_0_  ;
  output \g757/_0_  ;
  output \g760/_0_  ;
  output \g768/_2_  ;
  output \g770/_2_  ;
  output \g773/_0_  ;
  output \g786/_2_  ;
  output \g792/_0_  ;
  output \g793/_0_  ;
  output \g796/_0_  ;
  output \g804/_0_  ;
  output \g808/_0_  ;
  output \g817/_0_  ;
  output \g825/_0_  ;
  output \g834/_0_  ;
  output \g837/_0_  ;
  output \g838/_0_  ;
  output \g839/_0_  ;
  output \g840/_0_  ;
  output \g843/_0_  ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 ;
  assign n21 = ~\G11_reg/NET0131  & ~\G12_reg/NET0131  ;
  assign n22 = ~\G13_reg/NET0131  & n21 ;
  assign n23 = \G14_reg/NET0131  & ~n22 ;
  assign n24 = ~\G31_reg/NET0131  & ~n23 ;
  assign n25 = ~\G15_reg/NET0131  & ~\G16_reg/NET0131  ;
  assign n26 = ~\G17_reg/NET0131  & n25 ;
  assign n27 = \G18_reg/NET0131  & ~n26 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = ~\G19_reg/NET0131  & ~\G20_reg/NET0131  ;
  assign n30 = ~\G21_reg/NET0131  & n29 ;
  assign n31 = n28 & ~n30 ;
  assign n32 = \G22_reg/NET0131  & n31 ;
  assign n33 = ~\G0_pad  & ~n32 ;
  assign n34 = \G19_reg/NET0131  & \G20_reg/NET0131  ;
  assign n35 = n28 & n34 ;
  assign n36 = \G19_reg/NET0131  & n28 ;
  assign n37 = ~\G20_reg/NET0131  & ~n36 ;
  assign n38 = ~n35 & ~n37 ;
  assign n39 = n33 & n38 ;
  assign n40 = \G15_reg/NET0131  & ~n24 ;
  assign n41 = \G16_reg/NET0131  & n40 ;
  assign n42 = \G17_reg/NET0131  & n41 ;
  assign n43 = ~\G0_pad  & ~n28 ;
  assign n44 = \G18_reg/NET0131  & n43 ;
  assign n45 = ~n42 & n44 ;
  assign n46 = ~\G0_pad  & ~\G18_reg/NET0131  ;
  assign n47 = n42 & n46 ;
  assign n48 = ~n45 & ~n47 ;
  assign n49 = \G22_reg/NET0131  & ~n31 ;
  assign n50 = \G21_reg/NET0131  & ~\G22_reg/NET0131  ;
  assign n51 = n35 & n50 ;
  assign n52 = ~n49 & ~n51 ;
  assign n53 = ~\G0_pad  & ~n52 ;
  assign n54 = ~\G17_reg/NET0131  & ~n41 ;
  assign n55 = ~n42 & n43 ;
  assign n56 = ~n54 & n55 ;
  assign n57 = ~\G21_reg/NET0131  & ~n35 ;
  assign n58 = \G21_reg/NET0131  & n35 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = n33 & n59 ;
  assign n61 = ~\G19_reg/NET0131  & ~n28 ;
  assign n62 = ~n36 & ~n61 ;
  assign n63 = n33 & n62 ;
  assign n64 = ~\G16_reg/NET0131  & ~n40 ;
  assign n65 = ~n41 & n43 ;
  assign n66 = ~n64 & n65 ;
  assign n67 = \G11_reg/NET0131  & \G12_reg/NET0131  ;
  assign n68 = \G13_reg/NET0131  & n67 ;
  assign n69 = ~\G14_reg/NET0131  & ~n68 ;
  assign n70 = ~\G0_pad  & ~n23 ;
  assign n71 = ~n69 & n70 ;
  assign n75 = \G19_reg/NET0131  & ~\G20_reg/NET0131  ;
  assign n76 = ~\G23_reg/NET0131  & n50 ;
  assign n77 = n75 & n76 ;
  assign n78 = \G24_reg/NET0131  & ~n77 ;
  assign n79 = ~\G0_pad  & n78 ;
  assign n80 = ~\G0_pad  & \G21_reg/NET0131  ;
  assign n81 = \G23_reg/NET0131  & n29 ;
  assign n82 = n80 & n81 ;
  assign n83 = ~n79 & ~n82 ;
  assign n84 = \G17_reg/NET0131  & ~n83 ;
  assign n72 = ~\G21_reg/NET0131  & ~\G24_reg/NET0131  ;
  assign n73 = \G22_reg/NET0131  & n29 ;
  assign n74 = n72 & ~n73 ;
  assign n85 = ~\G0_pad  & ~n74 ;
  assign n86 = ~n84 & n85 ;
  assign n87 = ~\G15_reg/NET0131  & n24 ;
  assign n88 = ~n40 & ~n87 ;
  assign n89 = n43 & n88 ;
  assign n90 = ~\G21_reg/NET0131  & \G22_reg/NET0131  ;
  assign n91 = \G23_reg/NET0131  & n50 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = ~\G0_pad  & n29 ;
  assign n94 = ~n92 & n93 ;
  assign n95 = ~n79 & ~n94 ;
  assign n96 = ~n84 & ~n95 ;
  assign n97 = ~\G13_reg/NET0131  & ~n67 ;
  assign n98 = ~n68 & ~n97 ;
  assign n99 = n70 & n98 ;
  assign n100 = ~\G22_reg/NET0131  & ~n29 ;
  assign n101 = \G23_reg/NET0131  & ~n100 ;
  assign n102 = n80 & ~n101 ;
  assign n103 = ~n78 & n102 ;
  assign n104 = ~n21 & ~n67 ;
  assign n105 = n70 & n104 ;
  assign n106 = ~\G19_reg/NET0131  & \G22_reg/NET0131  ;
  assign n107 = ~n34 & n72 ;
  assign n108 = ~n106 & n107 ;
  assign n109 = ~\G0_pad  & ~n108 ;
  assign n110 = \G22_reg/NET0131  & ~n75 ;
  assign n111 = n72 & ~n110 ;
  assign n112 = ~\G0_pad  & ~n111 ;
  assign n113 = ~\G11_reg/NET0131  & n70 ;
  assign n114 = \G1_pad  & ~\G31_reg/NET0131  ;
  assign n115 = ~\G1_pad  & \G31_reg/NET0131  ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = ~\G0_pad  & ~n116 ;
  assign n118 = \G23_reg/NET0131  & ~\G2_pad  ;
  assign n119 = ~\G23_reg/NET0131  & \G2_pad  ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = ~\G0_pad  & ~n120 ;
  assign n122 = ~\G0_pad  & n34 ;
  assign n123 = n72 & n122 ;
  assign \G119_pad  = ~\G28_reg/NET0131  ;
  assign \G167_pad  = ~\G29_reg/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g43/_3_  = n39 ;
  assign \g754/_0_  = ~n48 ;
  assign \g757/_0_  = n53 ;
  assign \g760/_0_  = n56 ;
  assign \g768/_2_  = n60 ;
  assign \g770/_2_  = n63 ;
  assign \g773/_0_  = n66 ;
  assign \g786/_2_  = n71 ;
  assign \g792/_0_  = ~n86 ;
  assign \g793/_0_  = n89 ;
  assign \g796/_0_  = ~n96 ;
  assign \g804/_0_  = n99 ;
  assign \g808/_0_  = n103 ;
  assign \g817/_0_  = ~n83 ;
  assign \g825/_0_  = n105 ;
  assign \g834/_0_  = ~n109 ;
  assign \g837/_0_  = ~n112 ;
  assign \g838/_0_  = n113 ;
  assign \g839/_0_  = n117 ;
  assign \g840/_0_  = n121 ;
  assign \g843/_0_  = n123 ;
endmodule
