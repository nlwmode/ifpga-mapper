module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	output q_pad ;
	output r_pad ;
	output s_pad ;
	output t_pad ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		h_pad,
		i_pad,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		k_pad,
		l_pad,
		_w18_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		f_pad,
		g_pad,
		_w19_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		a_pad,
		b_pad,
		_w20_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		c_pad,
		d_pad,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		e_pad,
		j_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w21_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w17_,
		_w20_,
		_w24_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w18_,
		_w19_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w24_,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w23_,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		i_pad,
		j_pad,
		_w28_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w17_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		l_pad,
		m_pad,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w18_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		n_pad,
		o_pad,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		m_pad,
		n_pad,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		j_pad,
		k_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		g_pad,
		h_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w19_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		e_pad,
		f_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		e_pad,
		p_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w29_,
		_w35_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w31_,
		_w34_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w37_,
		_w40_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w41_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		p_pad,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		o_pad,
		_w45_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		k_pad,
		p_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w28_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w30_,
		_w32_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w36_,
		_w38_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w49_,
		_w52_,
		_w53_
	);
	assign q_pad = _w27_ ;
	assign r_pad = _w46_ ;
	assign s_pad = _w47_ ;
	assign t_pad = _w53_ ;
endmodule;