module top( \pi0000  , \pi0001  , \pi0002  , \pi0003  , \pi0004  , \pi0005  , \pi0006  , \pi0007  , \pi0008  , \pi0009  , \pi0010  , \pi0011  , \pi0012  , \pi0013  , \pi0014  , \pi0015  , \pi0016  , \pi0017  , \pi0018  , \pi0019  , \pi0020  , \pi0021  , \pi0022  , \pi0023  , \pi0024  , \pi0025  , \pi0026  , \pi0027  , \pi0028  , \pi0029  , \pi0030  , \pi0031  , \pi0032  , \pi0033  , \pi0034  , \pi0035  , \pi0036  , \pi0037  , \pi0038  , \pi0039  , \pi0040  , \pi0041  , \pi0042  , \pi0043  , \pi0044  , \pi0045  , \pi0046  , \pi0047  , \pi0048  , \pi0049  , \pi0050  , \pi0051  , \pi0052  , \pi0053  , \pi0054  , \pi0055  , \pi0056  , \pi0057  , \pi0058  , \pi0059  , \pi0060  , \pi0061  , \pi0062  , \pi0063  , \pi0064  , \pi0065  , \pi0066  , \pi0067  , \pi0068  , \pi0069  , \pi0070  , \pi0071  , \pi0072  , \pi0073  , \pi0074  , \pi0075  , \pi0076  , \pi0077  , \pi0078  , \pi0079  , \pi0080  , \pi0081  , \pi0082  , \pi0083  , \pi0084  , \pi0085  , \pi0086  , \pi0087  , \pi0088  , \pi0089  , \pi0090  , \pi0091  , \pi0092  , \pi0093  , \pi0094  , \pi0095  , \pi0096  , \pi0097  , \pi0098  , \pi0099  , \pi0100  , \pi0101  , \pi0102  , \pi0103  , \pi0104  , \pi0105  , \pi0106  , \pi0107  , \pi0108  , \pi0109  , \pi0110  , \pi0111  , \pi0112  , \pi0113  , \pi0114  , \pi0115  , \pi0116  , \pi0117  , \pi0118  , \pi0119  , \pi0120  , \pi0121  , \pi0122  , \pi0123  , \pi0124  , \pi0125  , \pi0126  , \pi0127  , \pi0128  , \pi0129  , \pi0130  , \pi0131  , \pi0132  , \pi0133  , \pi0134  , \pi0135  , \pi0136  , \pi0137  , \pi0138  , \pi0139  , \pi0140  , \pi0141  , \pi0142  , \pi0143  , \pi0144  , \pi0145  , \pi0146  , \pi0147  , \pi0148  , \pi0149  , \pi0150  , \pi0151  , \pi0152  , \pi0153  , \pi0154  , \pi0155  , \pi0156  , \pi0157  , \pi0158  , \pi0159  , \pi0160  , \pi0161  , \pi0162  , \pi0163  , \pi0164  , \pi0165  , \pi0166  , \pi0167  , \pi0168  , \pi0169  , \pi0170  , \pi0171  , \pi0172  , \pi0173  , \pi0174  , \pi0175  , \pi0176  , \pi0177  , \pi0178  , \pi0179  , \pi0180  , \pi0181  , \pi0182  , \pi0183  , \pi0184  , \pi0185  , \pi0186  , \pi0187  , \pi0188  , \pi0189  , \pi0190  , \pi0191  , \pi0192  , \pi0193  , \pi0194  , \pi0195  , \pi0196  , \pi0197  , \pi0198  , \pi0199  , \pi0200  , \pi0201  , \pi0202  , \pi0203  , \pi0204  , \pi0205  , \pi0206  , \pi0207  , \pi0208  , \pi0209  , \pi0210  , \pi0211  , \pi0212  , \pi0213  , \pi0214  , \pi0215  , \pi0216  , \pi0217  , \pi0218  , \pi0219  , \pi0220  , \pi0221  , \pi0222  , \pi0223  , \pi0224  , \pi0225  , \pi0226  , \pi0227  , \pi0228  , \pi0229  , \pi0230  , \pi0231  , \pi0232  , \pi0233  , \pi0234  , \pi0235  , \pi0236  , \pi0237  , \pi0238  , \pi0239  , \pi0240  , \pi0241  , \pi0242  , \pi0243  , \pi0244  , \pi0245  , \pi0246  , \pi0247  , \pi0248  , \pi0249  , \pi0250  , \pi0251  , \pi0252  , \pi0253  , \pi0254  , \pi0255  , \pi0256  , \pi0257  , \pi0258  , \pi0259  , \pi0260  , \pi0261  , \pi0262  , \pi0263  , \pi0264  , \pi0265  , \pi0266  , \pi0267  , \pi0268  , \pi0269  , \pi0270  , \pi0271  , \pi0272  , \pi0273  , \pi0274  , \pi0275  , \pi0276  , \pi0277  , \pi0278  , \pi0279  , \pi0280  , \pi0281  , \pi0282  , \pi0283  , \pi0284  , \pi0285  , \pi0286  , \pi0287  , \pi0288  , \pi0289  , \pi0290  , \pi0291  , \pi0292  , \pi0293  , \pi0294  , \pi0295  , \pi0296  , \pi0297  , \pi0298  , \pi0299  , \pi0300  , \pi0301  , \pi0302  , \pi0303  , \pi0304  , \pi0305  , \pi0306  , \pi0307  , \pi0308  , \pi0309  , \pi0310  , \pi0311  , \pi0312  , \pi0313  , \pi0314  , \pi0315  , \pi0316  , \pi0317  , \pi0318  , \pi0319  , \pi0320  , \pi0321  , \pi0322  , \pi0323  , \pi0324  , \pi0325  , \pi0326  , \pi0327  , \pi0328  , \pi0329  , \pi0330  , \pi0331  , \pi0332  , \pi0333  , \pi0334  , \pi0335  , \pi0336  , \pi0337  , \pi0338  , \pi0339  , \pi0340  , \pi0341  , \pi0342  , \pi0343  , \pi0344  , \pi0345  , \pi0346  , \pi0347  , \pi0348  , \pi0349  , \pi0350  , \pi0351  , \pi0352  , \pi0353  , \pi0354  , \pi0355  , \pi0356  , \pi0357  , \pi0358  , \pi0359  , \pi0360  , \pi0361  , \pi0362  , \pi0363  , \pi0364  , \pi0365  , \pi0366  , \pi0367  , \pi0368  , \pi0369  , \pi0370  , \pi0371  , \pi0372  , \pi0373  , \pi0374  , \pi0375  , \pi0376  , \pi0377  , \pi0378  , \pi0379  , \pi0380  , \pi0381  , \pi0382  , \pi0383  , \pi0384  , \pi0385  , \pi0386  , \pi0387  , \pi0388  , \pi0389  , \pi0390  , \pi0391  , \pi0392  , \pi0393  , \pi0394  , \pi0395  , \pi0396  , \pi0397  , \pi0398  , \pi0399  , \pi0400  , \pi0401  , \pi0402  , \pi0403  , \pi0404  , \pi0405  , \pi0406  , \pi0407  , \pi0408  , \pi0409  , \pi0410  , \pi0411  , \pi0412  , \pi0413  , \pi0414  , \pi0415  , \pi0416  , \pi0417  , \pi0418  , \pi0419  , \pi0420  , \pi0421  , \pi0422  , \pi0423  , \pi0424  , \pi0425  , \pi0426  , \pi0427  , \pi0428  , \pi0429  , \pi0430  , \pi0431  , \pi0432  , \pi0433  , \pi0434  , \pi0435  , \pi0436  , \pi0437  , \pi0438  , \pi0439  , \pi0440  , \pi0441  , \pi0442  , \pi0443  , \pi0444  , \pi0445  , \pi0446  , \pi0447  , \pi0448  , \pi0449  , \pi0450  , \pi0451  , \pi0452  , \pi0453  , \pi0454  , \pi0455  , \pi0456  , \pi0457  , \pi0458  , \pi0459  , \pi0460  , \pi0461  , \pi0462  , \pi0463  , \pi0464  , \pi0465  , \pi0466  , \pi0467  , \pi0468  , \pi0469  , \pi0470  , \pi0471  , \pi0472  , \pi0473  , \pi0474  , \pi0475  , \pi0476  , \pi0477  , \pi0478  , \pi0479  , \pi0480  , \pi0481  , \pi0482  , \pi0483  , \pi0484  , \pi0485  , \pi0486  , \pi0487  , \pi0488  , \pi0489  , \pi0490  , \pi0491  , \pi0492  , \pi0493  , \pi0494  , \pi0495  , \pi0496  , \pi0497  , \pi0498  , \pi0499  , \pi0500  , \pi0501  , \pi0502  , \pi0503  , \pi0504  , \pi0505  , \pi0506  , \pi0507  , \pi0508  , \pi0509  , \pi0510  , \pi0511  , \pi0512  , \pi0513  , \pi0514  , \pi0515  , \pi0516  , \pi0517  , \pi0518  , \pi0519  , \pi0520  , \pi0521  , \pi0522  , \pi0523  , \pi0524  , \pi0525  , \pi0526  , \pi0527  , \pi0528  , \pi0529  , \pi0530  , \pi0531  , \pi0532  , \pi0533  , \pi0534  , \pi0535  , \pi0536  , \pi0537  , \pi0538  , \pi0539  , \pi0540  , \pi0541  , \pi0542  , \pi0543  , \pi0544  , \pi0545  , \pi0546  , \pi0547  , \pi0548  , \pi0549  , \pi0550  , \pi0551  , \pi0552  , \pi0553  , \pi0554  , \pi0555  , \pi0556  , \pi0557  , \pi0558  , \pi0559  , \pi0560  , \pi0561  , \pi0562  , \pi0563  , \pi0564  , \pi0565  , \pi0566  , \pi0567  , \pi0568  , \pi0569  , \pi0570  , \pi0571  , \pi0572  , \pi0573  , \pi0574  , \pi0575  , \pi0576  , \pi0577  , \pi0578  , \pi0579  , \pi0580  , \pi0581  , \pi0582  , \pi0583  , \pi0584  , \pi0585  , \pi0586  , \pi0587  , \pi0588  , \pi0589  , \pi0590  , \pi0591  , \pi0592  , \pi0593  , \pi0594  , \pi0595  , \pi0596  , \pi0597  , \pi0598  , \pi0599  , \pi0600  , \pi0601  , \pi0602  , \pi0603  , \pi0604  , \pi0605  , \pi0606  , \pi0607  , \pi0608  , \pi0609  , \pi0610  , \pi0611  , \pi0612  , \pi0613  , \pi0614  , \pi0615  , \pi0616  , \pi0617  , \pi0618  , \pi0619  , \pi0620  , \pi0621  , \pi0622  , \pi0623  , \pi0624  , \pi0625  , \pi0626  , \pi0627  , \pi0628  , \pi0629  , \pi0630  , \pi0631  , \pi0632  , \pi0633  , \pi0634  , \pi0635  , \pi0636  , \pi0637  , \pi0638  , \pi0639  , \pi0640  , \pi0641  , \pi0642  , \pi0643  , \pi0644  , \pi0645  , \pi0646  , \pi0647  , \pi0648  , \pi0649  , \pi0650  , \pi0651  , \pi0652  , \pi0653  , \pi0654  , \pi0655  , \pi0656  , \pi0657  , \pi0658  , \pi0659  , \pi0660  , \pi0661  , \pi0662  , \pi0663  , \pi0664  , \pi0665  , \pi0666  , \pi0667  , \pi0668  , \pi0669  , \pi0670  , \pi0671  , \pi0672  , \pi0673  , \pi0674  , \pi0675  , \pi0676  , \pi0677  , \pi0678  , \pi0679  , \pi0680  , \pi0681  , \pi0682  , \pi0683  , \pi0684  , \pi0685  , \pi0686  , \pi0687  , \pi0688  , \pi0689  , \pi0690  , \pi0691  , \pi0692  , \pi0693  , \pi0694  , \pi0695  , \pi0696  , \pi0697  , \pi0698  , \pi0699  , \pi0700  , \pi0701  , \pi0702  , \pi0703  , \pi0704  , \pi0705  , \pi0706  , \pi0707  , \pi0708  , \pi0709  , \pi0710  , \pi0711  , \pi0712  , \pi0713  , \pi0714  , \pi0715  , \pi0716  , \pi0717  , \pi0718  , \pi0719  , \pi0720  , \pi0721  , \pi0722  , \pi0723  , \pi0724  , \pi0725  , \pi0726  , \pi0727  , \pi0728  , \pi0729  , \pi0730  , \pi0731  , \pi0732  , \pi0733  , \pi0734  , \pi0735  , \pi0736  , \pi0737  , \pi0738  , \pi0739  , \pi0740  , \pi0741  , \pi0742  , \pi0743  , \pi0744  , \pi0745  , \pi0746  , \pi0747  , \pi0748  , \pi0749  , \pi0750  , \pi0751  , \pi0752  , \pi0753  , \pi0754  , \pi0755  , \pi0756  , \pi0757  , \pi0758  , \pi0759  , \pi0760  , \pi0761  , \pi0762  , \pi0763  , \pi0764  , \pi0765  , \pi0766  , \pi0767  , \pi0768  , \pi0769  , \pi0770  , \pi0771  , \pi0772  , \pi0773  , \pi0774  , \pi0775  , \pi0776  , \pi0777  , \pi0778  , \pi0779  , \pi0780  , \pi0781  , \pi0782  , \pi0783  , \pi0784  , \pi0785  , \pi0786  , \pi0787  , \pi0788  , \pi0789  , \pi0790  , \pi0791  , \pi0792  , \pi0793  , \pi0794  , \pi0795  , \pi0796  , \pi0797  , \pi0798  , \pi0799  , \pi0800  , \pi0801  , \pi0802  , \pi0803  , \pi0804  , \pi0805  , \pi0806  , \pi0807  , \pi0808  , \pi0809  , \pi0810  , \pi0811  , \pi0812  , \pi0813  , \pi0814  , \pi0815  , \pi0816  , \pi0817  , \pi0818  , \pi0819  , \pi0820  , \pi0821  , \pi0822  , \pi0823  , \pi0824  , \pi0825  , \pi0826  , \pi0827  , \pi0828  , \pi0829  , \pi0830  , \pi0831  , \pi0832  , \pi0833  , \pi0834  , \pi0835  , \pi0836  , \pi0837  , \pi0838  , \pi0839  , \pi0840  , \pi0841  , \pi0842  , \pi0843  , \pi0844  , \pi0845  , \pi0846  , \pi0847  , \pi0848  , \pi0849  , \pi0850  , \pi0851  , \pi0852  , \pi0853  , \pi0854  , \pi0855  , \pi0856  , \pi0857  , \pi0858  , \pi0859  , \pi0860  , \pi0861  , \pi0862  , \pi0863  , \pi0864  , \pi0865  , \pi0866  , \pi0867  , \pi0868  , \pi0869  , \pi0870  , \pi0871  , \pi0872  , \pi0873  , \pi0874  , \pi0875  , \pi0876  , \pi0877  , \pi0878  , \pi0879  , \pi0880  , \pi0881  , \pi0882  , \pi0883  , \pi0884  , \pi0885  , \pi0886  , \pi0887  , \pi0888  , \pi0889  , \pi0890  , \pi0891  , \pi0892  , \pi0893  , \pi0894  , \pi0895  , \pi0896  , \pi0897  , \pi0898  , \pi0899  , \pi0900  , \pi0901  , \pi0902  , \pi0903  , \pi0904  , \pi0905  , \pi0906  , \pi0907  , \pi0908  , \pi0909  , \pi0910  , \pi0911  , \pi0912  , \pi0913  , \pi0914  , \pi0915  , \pi0916  , \pi0917  , \pi0918  , \pi0919  , \pi0920  , \pi0921  , \pi0922  , \pi0923  , \pi0924  , \pi0925  , \pi0926  , \pi0927  , \pi0928  , \pi0929  , \pi0930  , \pi0931  , \pi0932  , \pi0933  , \pi0934  , \pi0935  , \pi0936  , \pi0937  , \pi0938  , \pi0939  , \pi0940  , \pi0941  , \pi0942  , \pi0943  , \pi0944  , \pi0945  , \pi0946  , \pi0947  , \pi0948  , \pi0949  , \pi0950  , \pi0951  , \pi0952  , \pi0953  , \pi0954  , \pi0955  , \pi0956  , \pi0957  , \pi0958  , \pi0959  , \pi0960  , \pi0961  , \pi0962  , \pi0963  , \pi0964  , \pi0965  , \pi0966  , \pi0967  , \pi0968  , \pi0969  , \pi0970  , \pi0971  , \pi0972  , \pi0973  , \pi0974  , \pi0975  , \pi0976  , \pi0977  , \pi0978  , \pi0979  , \pi0980  , \pi0981  , \pi0982  , \pi0983  , \pi0984  , \pi0985  , \pi0986  , \pi0987  , \pi0988  , \pi0989  , \pi0990  , \pi0991  , \pi0992  , \pi0993  , \pi0994  , \pi0995  , \pi0996  , \pi0997  , \pi0998  , \pi0999  , \pi1000  , \pi1001  , \pi1002  , \pi1003  , \pi1004  , \pi1005  , \pi1006  , \pi1007  , \pi1008  , \pi1009  , \pi1010  , \pi1011  , \pi1012  , \pi1013  , \pi1014  , \pi1015  , \pi1016  , \pi1017  , \pi1018  , \pi1019  , \pi1020  , \pi1021  , \pi1022  , \pi1023  , \pi1024  , \pi1025  , \pi1026  , \pi1027  , \pi1028  , \pi1029  , \pi1030  , \pi1031  , \pi1032  , \pi1033  , \pi1034  , \pi1035  , \pi1036  , \pi1037  , \pi1038  , \pi1039  , \pi1040  , \pi1041  , \pi1042  , \pi1043  , \pi1044  , \pi1045  , \pi1046  , \pi1047  , \pi1048  , \pi1049  , \pi1050  , \pi1051  , \pi1052  , \pi1053  , \pi1054  , \pi1055  , \pi1056  , \pi1057  , \pi1058  , \pi1059  , \pi1060  , \pi1061  , \pi1062  , \pi1063  , \pi1064  , \pi1065  , \pi1066  , \pi1067  , \pi1068  , \pi1069  , \pi1070  , \pi1071  , \pi1072  , \pi1073  , \pi1074  , \pi1075  , \pi1076  , \pi1077  , \pi1078  , \pi1079  , \pi1080  , \pi1081  , \pi1082  , \pi1083  , \pi1084  , \pi1085  , \pi1086  , \pi1087  , \pi1088  , \pi1089  , \pi1090  , \pi1091  , \pi1092  , \pi1093  , \pi1094  , \pi1095  , \pi1096  , \pi1097  , \pi1098  , \pi1099  , \pi1100  , \pi1101  , \pi1102  , \pi1103  , \pi1104  , \pi1105  , \pi1106  , \pi1107  , \pi1108  , \pi1109  , \pi1110  , \pi1111  , \pi1112  , \pi1113  , \pi1114  , \pi1115  , \pi1116  , \pi1117  , \pi1118  , \pi1119  , \pi1120  , \pi1121  , \pi1122  , \pi1123  , \pi1124  , \pi1125  , \pi1126  , \pi1127  , \pi1128  , \pi1129  , \pi1130  , \pi1131  , \pi1132  , \pi1133  , \pi1134  , \pi1135  , \pi1136  , \pi1137  , \pi1138  , \pi1139  , \pi1140  , \pi1141  , \pi1142  , \pi1143  , \pi1144  , \pi1145  , \pi1146  , \pi1147  , \pi1148  , \pi1149  , \pi1150  , \pi1151  , \pi1152  , \pi1153  , \pi1154  , \pi1155  , \pi1156  , \pi1157  , \pi1158  , \pi1159  , \pi1160  , \pi1161  , \pi1162  , \pi1163  , \pi1164  , \pi1165  , \pi1166  , \pi1167  , \pi1168  , \pi1169  , \pi1170  , \pi1171  , \pi1172  , \pi1173  , \pi1174  , \pi1175  , \pi1176  , \pi1177  , \pi1178  , \pi1179  , \pi1180  , \pi1181  , \pi1182  , \pi1183  , \pi1184  , \pi1185  , \pi1186  , \pi1187  , \pi1188  , \pi1189  , \pi1190  , \pi1191  , \pi1192  , \pi1193  , \pi1194  , \pi1195  , \pi1196  , \pi1197  , \pi1198  , \pi1199  , \pi1200  , \pi1201  , \pi1202  , \pi1203  , \po0000  , \po0001  , \po0002  , \po0003  , \po0004  , \po0005  , \po0006  , \po0007  , \po0008  , \po0009  , \po0010  , \po0011  , \po0012  , \po0013  , \po0014  , \po0015  , \po0016  , \po0017  , \po0018  , \po0019  , \po0020  , \po0021  , \po0022  , \po0023  , \po0024  , \po0025  , \po0026  , \po0027  , \po0028  , \po0029  , \po0030  , \po0031  , \po0032  , \po0033  , \po0034  , \po0035  , \po0036  , \po0037  , \po0038  , \po0039  , \po0040  , \po0041  , \po0042  , \po0043  , \po0044  , \po0045  , \po0046  , \po0047  , \po0048  , \po0049  , \po0050  , \po0051  , \po0052  , \po0053  , \po0054  , \po0055  , \po0056  , \po0057  , \po0058  , \po0059  , \po0060  , \po0061  , \po0062  , \po0063  , \po0064  , \po0065  , \po0066  , \po0067  , \po0068  , \po0069  , \po0070  , \po0071  , \po0072  , \po0073  , \po0074  , \po0075  , \po0076  , \po0077  , \po0078  , \po0079  , \po0080  , \po0081  , \po0082  , \po0083  , \po0084  , \po0085  , \po0086  , \po0087  , \po0088  , \po0089  , \po0090  , \po0091  , \po0092  , \po0093  , \po0094  , \po0095  , \po0096  , \po0097  , \po0098  , \po0099  , \po0100  , \po0101  , \po0102  , \po0103  , \po0104  , \po0105  , \po0106  , \po0107  , \po0108  , \po0109  , \po0110  , \po0111  , \po0112  , \po0113  , \po0114  , \po0115  , \po0116  , \po0117  , \po0118  , \po0119  , \po0120  , \po0121  , \po0122  , \po0123  , \po0124  , \po0125  , \po0126  , \po0127  , \po0128  , \po0129  , \po0130  , \po0131  , \po0132  , \po0133  , \po0134  , \po0135  , \po0136  , \po0137  , \po0138  , \po0139  , \po0140  , \po0141  , \po0142  , \po0143  , \po0144  , \po0145  , \po0146  , \po0147  , \po0148  , \po0149  , \po0150  , \po0151  , \po0152  , \po0153  , \po0154  , \po0155  , \po0156  , \po0157  , \po0158  , \po0159  , \po0160  , \po0161  , \po0162  , \po0163  , \po0164  , \po0165  , \po0166  , \po0167  , \po0168  , \po0169  , \po0170  , \po0171  , \po0172  , \po0173  , \po0174  , \po0175  , \po0176  , \po0177  , \po0178  , \po0179  , \po0180  , \po0181  , \po0182  , \po0183  , \po0184  , \po0185  , \po0186  , \po0187  , \po0188  , \po0189  , \po0190  , \po0191  , \po0192  , \po0193  , \po0194  , \po0195  , \po0196  , \po0197  , \po0198  , \po0199  , \po0200  , \po0201  , \po0202  , \po0203  , \po0204  , \po0205  , \po0206  , \po0207  , \po0208  , \po0209  , \po0210  , \po0211  , \po0212  , \po0213  , \po0214  , \po0215  , \po0216  , \po0217  , \po0218  , \po0219  , \po0220  , \po0221  , \po0222  , \po0223  , \po0224  , \po0225  , \po0226  , \po0227  , \po0228  , \po0229  , \po0230  , \po0231  , \po0232  , \po0233  , \po0234  , \po0235  , \po0236  , \po0237  , \po0238  , \po0239  , \po0240  , \po0241  , \po0242  , \po0243  , \po0244  , \po0245  , \po0246  , \po0247  , \po0248  , \po0249  , \po0250  , \po0251  , \po0252  , \po0253  , \po0254  , \po0255  , \po0256  , \po0257  , \po0258  , \po0259  , \po0260  , \po0261  , \po0262  , \po0263  , \po0264  , \po0265  , \po0266  , \po0267  , \po0268  , \po0269  , \po0270  , \po0271  , \po0272  , \po0273  , \po0274  , \po0275  , \po0276  , \po0277  , \po0278  , \po0279  , \po0280  , \po0281  , \po0282  , \po0283  , \po0284  , \po0285  , \po0286  , \po0287  , \po0288  , \po0289  , \po0290  , \po0291  , \po0292  , \po0293  , \po0294  , \po0295  , \po0296  , \po0297  , \po0298  , \po0299  , \po0300  , \po0301  , \po0302  , \po0303  , \po0304  , \po0305  , \po0306  , \po0307  , \po0308  , \po0309  , \po0310  , \po0311  , \po0312  , \po0313  , \po0314  , \po0315  , \po0316  , \po0317  , \po0318  , \po0319  , \po0320  , \po0321  , \po0322  , \po0323  , \po0324  , \po0325  , \po0326  , \po0327  , \po0328  , \po0329  , \po0330  , \po0331  , \po0332  , \po0333  , \po0334  , \po0335  , \po0336  , \po0337  , \po0338  , \po0339  , \po0340  , \po0341  , \po0342  , \po0343  , \po0344  , \po0345  , \po0346  , \po0347  , \po0348  , \po0349  , \po0350  , \po0351  , \po0352  , \po0353  , \po0354  , \po0355  , \po0356  , \po0357  , \po0358  , \po0359  , \po0360  , \po0361  , \po0362  , \po0363  , \po0364  , \po0365  , \po0366  , \po0367  , \po0368  , \po0369  , \po0370  , \po0371  , \po0372  , \po0373  , \po0374  , \po0375  , \po0376  , \po0377  , \po0378  , \po0379  , \po0380  , \po0381  , \po0382  , \po0383  , \po0384  , \po0385  , \po0386  , \po0387  , \po0388  , \po0389  , \po0390  , \po0391  , \po0392  , \po0393  , \po0394  , \po0395  , \po0396  , \po0397  , \po0398  , \po0399  , \po0400  , \po0401  , \po0402  , \po0403  , \po0404  , \po0405  , \po0406  , \po0407  , \po0408  , \po0409  , \po0410  , \po0411  , \po0412  , \po0413  , \po0414  , \po0415  , \po0416  , \po0417  , \po0418  , \po0419  , \po0420  , \po0421  , \po0422  , \po0423  , \po0424  , \po0425  , \po0426  , \po0427  , \po0428  , \po0429  , \po0430  , \po0431  , \po0432  , \po0433  , \po0434  , \po0435  , \po0436  , \po0437  , \po0438  , \po0439  , \po0440  , \po0441  , \po0442  , \po0443  , \po0444  , \po0445  , \po0446  , \po0447  , \po0448  , \po0449  , \po0450  , \po0451  , \po0452  , \po0453  , \po0454  , \po0455  , \po0456  , \po0457  , \po0458  , \po0459  , \po0460  , \po0461  , \po0462  , \po0463  , \po0464  , \po0465  , \po0466  , \po0467  , \po0468  , \po0469  , \po0470  , \po0471  , \po0472  , \po0473  , \po0474  , \po0475  , \po0476  , \po0477  , \po0478  , \po0479  , \po0480  , \po0481  , \po0482  , \po0483  , \po0484  , \po0485  , \po0486  , \po0487  , \po0488  , \po0489  , \po0490  , \po0491  , \po0492  , \po0493  , \po0494  , \po0495  , \po0496  , \po0497  , \po0498  , \po0499  , \po0500  , \po0501  , \po0502  , \po0503  , \po0504  , \po0505  , \po0506  , \po0507  , \po0508  , \po0509  , \po0510  , \po0511  , \po0512  , \po0513  , \po0514  , \po0515  , \po0516  , \po0517  , \po0518  , \po0519  , \po0520  , \po0521  , \po0522  , \po0523  , \po0524  , \po0525  , \po0526  , \po0527  , \po0528  , \po0529  , \po0530  , \po0531  , \po0532  , \po0533  , \po0534  , \po0535  , \po0536  , \po0537  , \po0538  , \po0539  , \po0540  , \po0541  , \po0542  , \po0543  , \po0544  , \po0545  , \po0546  , \po0547  , \po0548  , \po0549  , \po0550  , \po0551  , \po0552  , \po0553  , \po0554  , \po0555  , \po0556  , \po0557  , \po0558  , \po0559  , \po0560  , \po0561  , \po0562  , \po0563  , \po0564  , \po0565  , \po0566  , \po0567  , \po0568  , \po0569  , \po0570  , \po0571  , \po0572  , \po0573  , \po0574  , \po0575  , \po0576  , \po0577  , \po0578  , \po0579  , \po0580  , \po0581  , \po0582  , \po0583  , \po0584  , \po0585  , \po0586  , \po0587  , \po0588  , \po0589  , \po0590  , \po0591  , \po0592  , \po0593  , \po0594  , \po0595  , \po0596  , \po0597  , \po0598  , \po0599  , \po0600  , \po0601  , \po0602  , \po0603  , \po0604  , \po0605  , \po0606  , \po0607  , \po0608  , \po0609  , \po0610  , \po0611  , \po0612  , \po0613  , \po0614  , \po0615  , \po0616  , \po0617  , \po0618  , \po0619  , \po0620  , \po0621  , \po0622  , \po0623  , \po0624  , \po0625  , \po0626  , \po0627  , \po0628  , \po0629  , \po0630  , \po0631  , \po0632  , \po0633  , \po0634  , \po0635  , \po0636  , \po0637  , \po0638  , \po0639  , \po0640  , \po0641  , \po0642  , \po0643  , \po0644  , \po0645  , \po0646  , \po0647  , \po0648  , \po0649  , \po0650  , \po0651  , \po0652  , \po0653  , \po0654  , \po0655  , \po0656  , \po0657  , \po0658  , \po0659  , \po0660  , \po0661  , \po0662  , \po0663  , \po0664  , \po0665  , \po0666  , \po0667  , \po0668  , \po0669  , \po0670  , \po0671  , \po0672  , \po0673  , \po0674  , \po0675  , \po0676  , \po0677  , \po0678  , \po0679  , \po0680  , \po0681  , \po0682  , \po0683  , \po0684  , \po0685  , \po0686  , \po0687  , \po0688  , \po0689  , \po0690  , \po0691  , \po0692  , \po0693  , \po0694  , \po0695  , \po0696  , \po0697  , \po0698  , \po0699  , \po0700  , \po0701  , \po0702  , \po0703  , \po0704  , \po0705  , \po0706  , \po0707  , \po0708  , \po0709  , \po0710  , \po0711  , \po0712  , \po0713  , \po0714  , \po0715  , \po0716  , \po0717  , \po0718  , \po0719  , \po0720  , \po0721  , \po0722  , \po0723  , \po0724  , \po0725  , \po0726  , \po0727  , \po0728  , \po0729  , \po0730  , \po0731  , \po0732  , \po0733  , \po0734  , \po0735  , \po0736  , \po0737  , \po0738  , \po0739  , \po0740  , \po0741  , \po0742  , \po0743  , \po0744  , \po0745  , \po0746  , \po0747  , \po0748  , \po0749  , \po0750  , \po0751  , \po0752  , \po0753  , \po0754  , \po0755  , \po0756  , \po0757  , \po0758  , \po0759  , \po0760  , \po0761  , \po0762  , \po0763  , \po0764  , \po0765  , \po0766  , \po0767  , \po0768  , \po0769  , \po0770  , \po0771  , \po0772  , \po0773  , \po0774  , \po0775  , \po0776  , \po0777  , \po0778  , \po0779  , \po0780  , \po0781  , \po0782  , \po0783  , \po0784  , \po0785  , \po0786  , \po0787  , \po0788  , \po0789  , \po0790  , \po0791  , \po0792  , \po0793  , \po0794  , \po0795  , \po0796  , \po0797  , \po0798  , \po0799  , \po0800  , \po0801  , \po0802  , \po0803  , \po0804  , \po0805  , \po0806  , \po0807  , \po0808  , \po0809  , \po0810  , \po0811  , \po0812  , \po0813  , \po0814  , \po0815  , \po0816  , \po0817  , \po0818  , \po0819  , \po0820  , \po0821  , \po0822  , \po0823  , \po0824  , \po0825  , \po0826  , \po0827  , \po0828  , \po0829  , \po0830  , \po0831  , \po0832  , \po0833  , \po0834  , \po0835  , \po0836  , \po0837  , \po0838  , \po0839  , \po0840  , \po0841  , \po0842  , \po0843  , \po0844  , \po0845  , \po0846  , \po0847  , \po0848  , \po0849  , \po0850  , \po0851  , \po0852  , \po0853  , \po0854  , \po0855  , \po0856  , \po0857  , \po0858  , \po0859  , \po0860  , \po0861  , \po0862  , \po0863  , \po0864  , \po0865  , \po0866  , \po0867  , \po0868  , \po0869  , \po0870  , \po0871  , \po0872  , \po0873  , \po0874  , \po0875  , \po0876  , \po0877  , \po0878  , \po0879  , \po0880  , \po0881  , \po0882  , \po0883  , \po0884  , \po0885  , \po0886  , \po0887  , \po0888  , \po0889  , \po0890  , \po0891  , \po0892  , \po0893  , \po0894  , \po0895  , \po0896  , \po0897  , \po0898  , \po0899  , \po0900  , \po0901  , \po0902  , \po0903  , \po0904  , \po0905  , \po0906  , \po0907  , \po0908  , \po0909  , \po0910  , \po0911  , \po0912  , \po0913  , \po0914  , \po0915  , \po0916  , \po0917  , \po0918  , \po0919  , \po0920  , \po0921  , \po0922  , \po0923  , \po0924  , \po0925  , \po0926  , \po0927  , \po0928  , \po0929  , \po0930  , \po0931  , \po0932  , \po0933  , \po0934  , \po0935  , \po0936  , \po0937  , \po0938  , \po0939  , \po0940  , \po0941  , \po0942  , \po0943  , \po0944  , \po0945  , \po0946  , \po0947  , \po0948  , \po0949  , \po0950  , \po0951  , \po0952  , \po0953  , \po0954  , \po0955  , \po0956  , \po0957  , \po0958  , \po0959  , \po0960  , \po0961  , \po0962  , \po0963  , \po0964  , \po0965  , \po0966  , \po0967  , \po0968  , \po0969  , \po0970  , \po0971  , \po0972  , \po0973  , \po0974  , \po0975  , \po0976  , \po0977  , \po0978  , \po0979  , \po0980  , \po0981  , \po0982  , \po0983  , \po0984  , \po0985  , \po0986  , \po0987  , \po0988  , \po0989  , \po0990  , \po0991  , \po0992  , \po0993  , \po0994  , \po0995  , \po0996  , \po0997  , \po0998  , \po0999  , \po1000  , \po1001  , \po1002  , \po1003  , \po1004  , \po1005  , \po1006  , \po1007  , \po1008  , \po1009  , \po1010  , \po1011  , \po1012  , \po1013  , \po1014  , \po1015  , \po1016  , \po1017  , \po1018  , \po1019  , \po1020  , \po1021  , \po1022  , \po1023  , \po1024  , \po1025  , \po1026  , \po1027  , \po1028  , \po1029  , \po1030  , \po1031  , \po1032  , \po1033  , \po1034  , \po1035  , \po1036  , \po1037  , \po1038  , \po1039  , \po1040  , \po1041  , \po1042  , \po1043  , \po1044  , \po1045  , \po1046  , \po1047  , \po1048  , \po1049  , \po1050  , \po1051  , \po1052  , \po1053  , \po1054  , \po1055  , \po1056  , \po1057  , \po1058  , \po1059  , \po1060  , \po1061  , \po1062  , \po1063  , \po1064  , \po1065  , \po1066  , \po1067  , \po1068  , \po1069  , \po1070  , \po1071  , \po1072  , \po1073  , \po1074  , \po1075  , \po1076  , \po1077  , \po1078  , \po1079  , \po1080  , \po1081  , \po1082  , \po1083  , \po1084  , \po1085  , \po1086  , \po1087  , \po1088  , \po1089  , \po1090  , \po1091  , \po1092  , \po1093  , \po1094  , \po1095  , \po1096  , \po1097  , \po1098  , \po1099  , \po1100  , \po1101  , \po1102  , \po1103  , \po1104  , \po1105  , \po1106  , \po1107  , \po1108  , \po1109  , \po1110  , \po1111  , \po1112  , \po1113  , \po1114  , \po1115  , \po1116  , \po1117  , \po1118  , \po1119  , \po1120  , \po1121  , \po1122  , \po1123  , \po1124  , \po1125  , \po1126  , \po1127  , \po1128  , \po1129  , \po1130  , \po1131  , \po1132  , \po1133  , \po1134  , \po1135  , \po1136  , \po1137  , \po1138  , \po1139  , \po1140  , \po1141  , \po1142  , \po1143  , \po1144  , \po1145  , \po1146  , \po1147  , \po1148  , \po1149  , \po1150  , \po1151  , \po1152  , \po1153  , \po1154  , \po1155  , \po1156  , \po1157  , \po1158  , \po1159  , \po1160  , \po1161  , \po1162  , \po1163  , \po1164  , \po1165  , \po1166  , \po1167  , \po1168  , \po1169  , \po1170  , \po1171  , \po1172  , \po1173  , \po1174  , \po1175  , \po1176  , \po1177  , \po1178  , \po1179  , \po1180  , \po1181  , \po1182  , \po1183  , \po1184  , \po1185  , \po1186  , \po1187  , \po1188  , \po1189  , \po1190  , \po1191  , \po1192  , \po1193  , \po1194  , \po1195  , \po1196  , \po1197  , \po1198  , \po1199  , \po1200  , \po1201  , \po1202  , \po1203  , \po1204  , \po1205  , \po1206  , \po1207  , \po1208  , \po1209  , \po1210  , \po1211  , \po1212  , \po1213  , \po1214  , \po1215  , \po1216  , \po1217  , \po1218  , \po1219  , \po1220  , \po1221  , \po1222  , \po1223  , \po1224  , \po1225  , \po1226  , \po1227  , \po1228  , \po1229  , \po1230  );
  input \pi0000  ;
  input \pi0001  ;
  input \pi0002  ;
  input \pi0003  ;
  input \pi0004  ;
  input \pi0005  ;
  input \pi0006  ;
  input \pi0007  ;
  input \pi0008  ;
  input \pi0009  ;
  input \pi0010  ;
  input \pi0011  ;
  input \pi0012  ;
  input \pi0013  ;
  input \pi0014  ;
  input \pi0015  ;
  input \pi0016  ;
  input \pi0017  ;
  input \pi0018  ;
  input \pi0019  ;
  input \pi0020  ;
  input \pi0021  ;
  input \pi0022  ;
  input \pi0023  ;
  input \pi0024  ;
  input \pi0025  ;
  input \pi0026  ;
  input \pi0027  ;
  input \pi0028  ;
  input \pi0029  ;
  input \pi0030  ;
  input \pi0031  ;
  input \pi0032  ;
  input \pi0033  ;
  input \pi0034  ;
  input \pi0035  ;
  input \pi0036  ;
  input \pi0037  ;
  input \pi0038  ;
  input \pi0039  ;
  input \pi0040  ;
  input \pi0041  ;
  input \pi0042  ;
  input \pi0043  ;
  input \pi0044  ;
  input \pi0045  ;
  input \pi0046  ;
  input \pi0047  ;
  input \pi0048  ;
  input \pi0049  ;
  input \pi0050  ;
  input \pi0051  ;
  input \pi0052  ;
  input \pi0053  ;
  input \pi0054  ;
  input \pi0055  ;
  input \pi0056  ;
  input \pi0057  ;
  input \pi0058  ;
  input \pi0059  ;
  input \pi0060  ;
  input \pi0061  ;
  input \pi0062  ;
  input \pi0063  ;
  input \pi0064  ;
  input \pi0065  ;
  input \pi0066  ;
  input \pi0067  ;
  input \pi0068  ;
  input \pi0069  ;
  input \pi0070  ;
  input \pi0071  ;
  input \pi0072  ;
  input \pi0073  ;
  input \pi0074  ;
  input \pi0075  ;
  input \pi0076  ;
  input \pi0077  ;
  input \pi0078  ;
  input \pi0079  ;
  input \pi0080  ;
  input \pi0081  ;
  input \pi0082  ;
  input \pi0083  ;
  input \pi0084  ;
  input \pi0085  ;
  input \pi0086  ;
  input \pi0087  ;
  input \pi0088  ;
  input \pi0089  ;
  input \pi0090  ;
  input \pi0091  ;
  input \pi0092  ;
  input \pi0093  ;
  input \pi0094  ;
  input \pi0095  ;
  input \pi0096  ;
  input \pi0097  ;
  input \pi0098  ;
  input \pi0099  ;
  input \pi0100  ;
  input \pi0101  ;
  input \pi0102  ;
  input \pi0103  ;
  input \pi0104  ;
  input \pi0105  ;
  input \pi0106  ;
  input \pi0107  ;
  input \pi0108  ;
  input \pi0109  ;
  input \pi0110  ;
  input \pi0111  ;
  input \pi0112  ;
  input \pi0113  ;
  input \pi0114  ;
  input \pi0115  ;
  input \pi0116  ;
  input \pi0117  ;
  input \pi0118  ;
  input \pi0119  ;
  input \pi0120  ;
  input \pi0121  ;
  input \pi0122  ;
  input \pi0123  ;
  input \pi0124  ;
  input \pi0125  ;
  input \pi0126  ;
  input \pi0127  ;
  input \pi0128  ;
  input \pi0129  ;
  input \pi0130  ;
  input \pi0131  ;
  input \pi0132  ;
  input \pi0133  ;
  input \pi0134  ;
  input \pi0135  ;
  input \pi0136  ;
  input \pi0137  ;
  input \pi0138  ;
  input \pi0139  ;
  input \pi0140  ;
  input \pi0141  ;
  input \pi0142  ;
  input \pi0143  ;
  input \pi0144  ;
  input \pi0145  ;
  input \pi0146  ;
  input \pi0147  ;
  input \pi0148  ;
  input \pi0149  ;
  input \pi0150  ;
  input \pi0151  ;
  input \pi0152  ;
  input \pi0153  ;
  input \pi0154  ;
  input \pi0155  ;
  input \pi0156  ;
  input \pi0157  ;
  input \pi0158  ;
  input \pi0159  ;
  input \pi0160  ;
  input \pi0161  ;
  input \pi0162  ;
  input \pi0163  ;
  input \pi0164  ;
  input \pi0165  ;
  input \pi0166  ;
  input \pi0167  ;
  input \pi0168  ;
  input \pi0169  ;
  input \pi0170  ;
  input \pi0171  ;
  input \pi0172  ;
  input \pi0173  ;
  input \pi0174  ;
  input \pi0175  ;
  input \pi0176  ;
  input \pi0177  ;
  input \pi0178  ;
  input \pi0179  ;
  input \pi0180  ;
  input \pi0181  ;
  input \pi0182  ;
  input \pi0183  ;
  input \pi0184  ;
  input \pi0185  ;
  input \pi0186  ;
  input \pi0187  ;
  input \pi0188  ;
  input \pi0189  ;
  input \pi0190  ;
  input \pi0191  ;
  input \pi0192  ;
  input \pi0193  ;
  input \pi0194  ;
  input \pi0195  ;
  input \pi0196  ;
  input \pi0197  ;
  input \pi0198  ;
  input \pi0199  ;
  input \pi0200  ;
  input \pi0201  ;
  input \pi0202  ;
  input \pi0203  ;
  input \pi0204  ;
  input \pi0205  ;
  input \pi0206  ;
  input \pi0207  ;
  input \pi0208  ;
  input \pi0209  ;
  input \pi0210  ;
  input \pi0211  ;
  input \pi0212  ;
  input \pi0213  ;
  input \pi0214  ;
  input \pi0215  ;
  input \pi0216  ;
  input \pi0217  ;
  input \pi0218  ;
  input \pi0219  ;
  input \pi0220  ;
  input \pi0221  ;
  input \pi0222  ;
  input \pi0223  ;
  input \pi0224  ;
  input \pi0225  ;
  input \pi0226  ;
  input \pi0227  ;
  input \pi0228  ;
  input \pi0229  ;
  input \pi0230  ;
  input \pi0231  ;
  input \pi0232  ;
  input \pi0233  ;
  input \pi0234  ;
  input \pi0235  ;
  input \pi0236  ;
  input \pi0237  ;
  input \pi0238  ;
  input \pi0239  ;
  input \pi0240  ;
  input \pi0241  ;
  input \pi0242  ;
  input \pi0243  ;
  input \pi0244  ;
  input \pi0245  ;
  input \pi0246  ;
  input \pi0247  ;
  input \pi0248  ;
  input \pi0249  ;
  input \pi0250  ;
  input \pi0251  ;
  input \pi0252  ;
  input \pi0253  ;
  input \pi0254  ;
  input \pi0255  ;
  input \pi0256  ;
  input \pi0257  ;
  input \pi0258  ;
  input \pi0259  ;
  input \pi0260  ;
  input \pi0261  ;
  input \pi0262  ;
  input \pi0263  ;
  input \pi0264  ;
  input \pi0265  ;
  input \pi0266  ;
  input \pi0267  ;
  input \pi0268  ;
  input \pi0269  ;
  input \pi0270  ;
  input \pi0271  ;
  input \pi0272  ;
  input \pi0273  ;
  input \pi0274  ;
  input \pi0275  ;
  input \pi0276  ;
  input \pi0277  ;
  input \pi0278  ;
  input \pi0279  ;
  input \pi0280  ;
  input \pi0281  ;
  input \pi0282  ;
  input \pi0283  ;
  input \pi0284  ;
  input \pi0285  ;
  input \pi0286  ;
  input \pi0287  ;
  input \pi0288  ;
  input \pi0289  ;
  input \pi0290  ;
  input \pi0291  ;
  input \pi0292  ;
  input \pi0293  ;
  input \pi0294  ;
  input \pi0295  ;
  input \pi0296  ;
  input \pi0297  ;
  input \pi0298  ;
  input \pi0299  ;
  input \pi0300  ;
  input \pi0301  ;
  input \pi0302  ;
  input \pi0303  ;
  input \pi0304  ;
  input \pi0305  ;
  input \pi0306  ;
  input \pi0307  ;
  input \pi0308  ;
  input \pi0309  ;
  input \pi0310  ;
  input \pi0311  ;
  input \pi0312  ;
  input \pi0313  ;
  input \pi0314  ;
  input \pi0315  ;
  input \pi0316  ;
  input \pi0317  ;
  input \pi0318  ;
  input \pi0319  ;
  input \pi0320  ;
  input \pi0321  ;
  input \pi0322  ;
  input \pi0323  ;
  input \pi0324  ;
  input \pi0325  ;
  input \pi0326  ;
  input \pi0327  ;
  input \pi0328  ;
  input \pi0329  ;
  input \pi0330  ;
  input \pi0331  ;
  input \pi0332  ;
  input \pi0333  ;
  input \pi0334  ;
  input \pi0335  ;
  input \pi0336  ;
  input \pi0337  ;
  input \pi0338  ;
  input \pi0339  ;
  input \pi0340  ;
  input \pi0341  ;
  input \pi0342  ;
  input \pi0343  ;
  input \pi0344  ;
  input \pi0345  ;
  input \pi0346  ;
  input \pi0347  ;
  input \pi0348  ;
  input \pi0349  ;
  input \pi0350  ;
  input \pi0351  ;
  input \pi0352  ;
  input \pi0353  ;
  input \pi0354  ;
  input \pi0355  ;
  input \pi0356  ;
  input \pi0357  ;
  input \pi0358  ;
  input \pi0359  ;
  input \pi0360  ;
  input \pi0361  ;
  input \pi0362  ;
  input \pi0363  ;
  input \pi0364  ;
  input \pi0365  ;
  input \pi0366  ;
  input \pi0367  ;
  input \pi0368  ;
  input \pi0369  ;
  input \pi0370  ;
  input \pi0371  ;
  input \pi0372  ;
  input \pi0373  ;
  input \pi0374  ;
  input \pi0375  ;
  input \pi0376  ;
  input \pi0377  ;
  input \pi0378  ;
  input \pi0379  ;
  input \pi0380  ;
  input \pi0381  ;
  input \pi0382  ;
  input \pi0383  ;
  input \pi0384  ;
  input \pi0385  ;
  input \pi0386  ;
  input \pi0387  ;
  input \pi0388  ;
  input \pi0389  ;
  input \pi0390  ;
  input \pi0391  ;
  input \pi0392  ;
  input \pi0393  ;
  input \pi0394  ;
  input \pi0395  ;
  input \pi0396  ;
  input \pi0397  ;
  input \pi0398  ;
  input \pi0399  ;
  input \pi0400  ;
  input \pi0401  ;
  input \pi0402  ;
  input \pi0403  ;
  input \pi0404  ;
  input \pi0405  ;
  input \pi0406  ;
  input \pi0407  ;
  input \pi0408  ;
  input \pi0409  ;
  input \pi0410  ;
  input \pi0411  ;
  input \pi0412  ;
  input \pi0413  ;
  input \pi0414  ;
  input \pi0415  ;
  input \pi0416  ;
  input \pi0417  ;
  input \pi0418  ;
  input \pi0419  ;
  input \pi0420  ;
  input \pi0421  ;
  input \pi0422  ;
  input \pi0423  ;
  input \pi0424  ;
  input \pi0425  ;
  input \pi0426  ;
  input \pi0427  ;
  input \pi0428  ;
  input \pi0429  ;
  input \pi0430  ;
  input \pi0431  ;
  input \pi0432  ;
  input \pi0433  ;
  input \pi0434  ;
  input \pi0435  ;
  input \pi0436  ;
  input \pi0437  ;
  input \pi0438  ;
  input \pi0439  ;
  input \pi0440  ;
  input \pi0441  ;
  input \pi0442  ;
  input \pi0443  ;
  input \pi0444  ;
  input \pi0445  ;
  input \pi0446  ;
  input \pi0447  ;
  input \pi0448  ;
  input \pi0449  ;
  input \pi0450  ;
  input \pi0451  ;
  input \pi0452  ;
  input \pi0453  ;
  input \pi0454  ;
  input \pi0455  ;
  input \pi0456  ;
  input \pi0457  ;
  input \pi0458  ;
  input \pi0459  ;
  input \pi0460  ;
  input \pi0461  ;
  input \pi0462  ;
  input \pi0463  ;
  input \pi0464  ;
  input \pi0465  ;
  input \pi0466  ;
  input \pi0467  ;
  input \pi0468  ;
  input \pi0469  ;
  input \pi0470  ;
  input \pi0471  ;
  input \pi0472  ;
  input \pi0473  ;
  input \pi0474  ;
  input \pi0475  ;
  input \pi0476  ;
  input \pi0477  ;
  input \pi0478  ;
  input \pi0479  ;
  input \pi0480  ;
  input \pi0481  ;
  input \pi0482  ;
  input \pi0483  ;
  input \pi0484  ;
  input \pi0485  ;
  input \pi0486  ;
  input \pi0487  ;
  input \pi0488  ;
  input \pi0489  ;
  input \pi0490  ;
  input \pi0491  ;
  input \pi0492  ;
  input \pi0493  ;
  input \pi0494  ;
  input \pi0495  ;
  input \pi0496  ;
  input \pi0497  ;
  input \pi0498  ;
  input \pi0499  ;
  input \pi0500  ;
  input \pi0501  ;
  input \pi0502  ;
  input \pi0503  ;
  input \pi0504  ;
  input \pi0505  ;
  input \pi0506  ;
  input \pi0507  ;
  input \pi0508  ;
  input \pi0509  ;
  input \pi0510  ;
  input \pi0511  ;
  input \pi0512  ;
  input \pi0513  ;
  input \pi0514  ;
  input \pi0515  ;
  input \pi0516  ;
  input \pi0517  ;
  input \pi0518  ;
  input \pi0519  ;
  input \pi0520  ;
  input \pi0521  ;
  input \pi0522  ;
  input \pi0523  ;
  input \pi0524  ;
  input \pi0525  ;
  input \pi0526  ;
  input \pi0527  ;
  input \pi0528  ;
  input \pi0529  ;
  input \pi0530  ;
  input \pi0531  ;
  input \pi0532  ;
  input \pi0533  ;
  input \pi0534  ;
  input \pi0535  ;
  input \pi0536  ;
  input \pi0537  ;
  input \pi0538  ;
  input \pi0539  ;
  input \pi0540  ;
  input \pi0541  ;
  input \pi0542  ;
  input \pi0543  ;
  input \pi0544  ;
  input \pi0545  ;
  input \pi0546  ;
  input \pi0547  ;
  input \pi0548  ;
  input \pi0549  ;
  input \pi0550  ;
  input \pi0551  ;
  input \pi0552  ;
  input \pi0553  ;
  input \pi0554  ;
  input \pi0555  ;
  input \pi0556  ;
  input \pi0557  ;
  input \pi0558  ;
  input \pi0559  ;
  input \pi0560  ;
  input \pi0561  ;
  input \pi0562  ;
  input \pi0563  ;
  input \pi0564  ;
  input \pi0565  ;
  input \pi0566  ;
  input \pi0567  ;
  input \pi0568  ;
  input \pi0569  ;
  input \pi0570  ;
  input \pi0571  ;
  input \pi0572  ;
  input \pi0573  ;
  input \pi0574  ;
  input \pi0575  ;
  input \pi0576  ;
  input \pi0577  ;
  input \pi0578  ;
  input \pi0579  ;
  input \pi0580  ;
  input \pi0581  ;
  input \pi0582  ;
  input \pi0583  ;
  input \pi0584  ;
  input \pi0585  ;
  input \pi0586  ;
  input \pi0587  ;
  input \pi0588  ;
  input \pi0589  ;
  input \pi0590  ;
  input \pi0591  ;
  input \pi0592  ;
  input \pi0593  ;
  input \pi0594  ;
  input \pi0595  ;
  input \pi0596  ;
  input \pi0597  ;
  input \pi0598  ;
  input \pi0599  ;
  input \pi0600  ;
  input \pi0601  ;
  input \pi0602  ;
  input \pi0603  ;
  input \pi0604  ;
  input \pi0605  ;
  input \pi0606  ;
  input \pi0607  ;
  input \pi0608  ;
  input \pi0609  ;
  input \pi0610  ;
  input \pi0611  ;
  input \pi0612  ;
  input \pi0613  ;
  input \pi0614  ;
  input \pi0615  ;
  input \pi0616  ;
  input \pi0617  ;
  input \pi0618  ;
  input \pi0619  ;
  input \pi0620  ;
  input \pi0621  ;
  input \pi0622  ;
  input \pi0623  ;
  input \pi0624  ;
  input \pi0625  ;
  input \pi0626  ;
  input \pi0627  ;
  input \pi0628  ;
  input \pi0629  ;
  input \pi0630  ;
  input \pi0631  ;
  input \pi0632  ;
  input \pi0633  ;
  input \pi0634  ;
  input \pi0635  ;
  input \pi0636  ;
  input \pi0637  ;
  input \pi0638  ;
  input \pi0639  ;
  input \pi0640  ;
  input \pi0641  ;
  input \pi0642  ;
  input \pi0643  ;
  input \pi0644  ;
  input \pi0645  ;
  input \pi0646  ;
  input \pi0647  ;
  input \pi0648  ;
  input \pi0649  ;
  input \pi0650  ;
  input \pi0651  ;
  input \pi0652  ;
  input \pi0653  ;
  input \pi0654  ;
  input \pi0655  ;
  input \pi0656  ;
  input \pi0657  ;
  input \pi0658  ;
  input \pi0659  ;
  input \pi0660  ;
  input \pi0661  ;
  input \pi0662  ;
  input \pi0663  ;
  input \pi0664  ;
  input \pi0665  ;
  input \pi0666  ;
  input \pi0667  ;
  input \pi0668  ;
  input \pi0669  ;
  input \pi0670  ;
  input \pi0671  ;
  input \pi0672  ;
  input \pi0673  ;
  input \pi0674  ;
  input \pi0675  ;
  input \pi0676  ;
  input \pi0677  ;
  input \pi0678  ;
  input \pi0679  ;
  input \pi0680  ;
  input \pi0681  ;
  input \pi0682  ;
  input \pi0683  ;
  input \pi0684  ;
  input \pi0685  ;
  input \pi0686  ;
  input \pi0687  ;
  input \pi0688  ;
  input \pi0689  ;
  input \pi0690  ;
  input \pi0691  ;
  input \pi0692  ;
  input \pi0693  ;
  input \pi0694  ;
  input \pi0695  ;
  input \pi0696  ;
  input \pi0697  ;
  input \pi0698  ;
  input \pi0699  ;
  input \pi0700  ;
  input \pi0701  ;
  input \pi0702  ;
  input \pi0703  ;
  input \pi0704  ;
  input \pi0705  ;
  input \pi0706  ;
  input \pi0707  ;
  input \pi0708  ;
  input \pi0709  ;
  input \pi0710  ;
  input \pi0711  ;
  input \pi0712  ;
  input \pi0713  ;
  input \pi0714  ;
  input \pi0715  ;
  input \pi0716  ;
  input \pi0717  ;
  input \pi0718  ;
  input \pi0719  ;
  input \pi0720  ;
  input \pi0721  ;
  input \pi0722  ;
  input \pi0723  ;
  input \pi0724  ;
  input \pi0725  ;
  input \pi0726  ;
  input \pi0727  ;
  input \pi0728  ;
  input \pi0729  ;
  input \pi0730  ;
  input \pi0731  ;
  input \pi0732  ;
  input \pi0733  ;
  input \pi0734  ;
  input \pi0735  ;
  input \pi0736  ;
  input \pi0737  ;
  input \pi0738  ;
  input \pi0739  ;
  input \pi0740  ;
  input \pi0741  ;
  input \pi0742  ;
  input \pi0743  ;
  input \pi0744  ;
  input \pi0745  ;
  input \pi0746  ;
  input \pi0747  ;
  input \pi0748  ;
  input \pi0749  ;
  input \pi0750  ;
  input \pi0751  ;
  input \pi0752  ;
  input \pi0753  ;
  input \pi0754  ;
  input \pi0755  ;
  input \pi0756  ;
  input \pi0757  ;
  input \pi0758  ;
  input \pi0759  ;
  input \pi0760  ;
  input \pi0761  ;
  input \pi0762  ;
  input \pi0763  ;
  input \pi0764  ;
  input \pi0765  ;
  input \pi0766  ;
  input \pi0767  ;
  input \pi0768  ;
  input \pi0769  ;
  input \pi0770  ;
  input \pi0771  ;
  input \pi0772  ;
  input \pi0773  ;
  input \pi0774  ;
  input \pi0775  ;
  input \pi0776  ;
  input \pi0777  ;
  input \pi0778  ;
  input \pi0779  ;
  input \pi0780  ;
  input \pi0781  ;
  input \pi0782  ;
  input \pi0783  ;
  input \pi0784  ;
  input \pi0785  ;
  input \pi0786  ;
  input \pi0787  ;
  input \pi0788  ;
  input \pi0789  ;
  input \pi0790  ;
  input \pi0791  ;
  input \pi0792  ;
  input \pi0793  ;
  input \pi0794  ;
  input \pi0795  ;
  input \pi0796  ;
  input \pi0797  ;
  input \pi0798  ;
  input \pi0799  ;
  input \pi0800  ;
  input \pi0801  ;
  input \pi0802  ;
  input \pi0803  ;
  input \pi0804  ;
  input \pi0805  ;
  input \pi0806  ;
  input \pi0807  ;
  input \pi0808  ;
  input \pi0809  ;
  input \pi0810  ;
  input \pi0811  ;
  input \pi0812  ;
  input \pi0813  ;
  input \pi0814  ;
  input \pi0815  ;
  input \pi0816  ;
  input \pi0817  ;
  input \pi0818  ;
  input \pi0819  ;
  input \pi0820  ;
  input \pi0821  ;
  input \pi0822  ;
  input \pi0823  ;
  input \pi0824  ;
  input \pi0825  ;
  input \pi0826  ;
  input \pi0827  ;
  input \pi0828  ;
  input \pi0829  ;
  input \pi0830  ;
  input \pi0831  ;
  input \pi0832  ;
  input \pi0833  ;
  input \pi0834  ;
  input \pi0835  ;
  input \pi0836  ;
  input \pi0837  ;
  input \pi0838  ;
  input \pi0839  ;
  input \pi0840  ;
  input \pi0841  ;
  input \pi0842  ;
  input \pi0843  ;
  input \pi0844  ;
  input \pi0845  ;
  input \pi0846  ;
  input \pi0847  ;
  input \pi0848  ;
  input \pi0849  ;
  input \pi0850  ;
  input \pi0851  ;
  input \pi0852  ;
  input \pi0853  ;
  input \pi0854  ;
  input \pi0855  ;
  input \pi0856  ;
  input \pi0857  ;
  input \pi0858  ;
  input \pi0859  ;
  input \pi0860  ;
  input \pi0861  ;
  input \pi0862  ;
  input \pi0863  ;
  input \pi0864  ;
  input \pi0865  ;
  input \pi0866  ;
  input \pi0867  ;
  input \pi0868  ;
  input \pi0869  ;
  input \pi0870  ;
  input \pi0871  ;
  input \pi0872  ;
  input \pi0873  ;
  input \pi0874  ;
  input \pi0875  ;
  input \pi0876  ;
  input \pi0877  ;
  input \pi0878  ;
  input \pi0879  ;
  input \pi0880  ;
  input \pi0881  ;
  input \pi0882  ;
  input \pi0883  ;
  input \pi0884  ;
  input \pi0885  ;
  input \pi0886  ;
  input \pi0887  ;
  input \pi0888  ;
  input \pi0889  ;
  input \pi0890  ;
  input \pi0891  ;
  input \pi0892  ;
  input \pi0893  ;
  input \pi0894  ;
  input \pi0895  ;
  input \pi0896  ;
  input \pi0897  ;
  input \pi0898  ;
  input \pi0899  ;
  input \pi0900  ;
  input \pi0901  ;
  input \pi0902  ;
  input \pi0903  ;
  input \pi0904  ;
  input \pi0905  ;
  input \pi0906  ;
  input \pi0907  ;
  input \pi0908  ;
  input \pi0909  ;
  input \pi0910  ;
  input \pi0911  ;
  input \pi0912  ;
  input \pi0913  ;
  input \pi0914  ;
  input \pi0915  ;
  input \pi0916  ;
  input \pi0917  ;
  input \pi0918  ;
  input \pi0919  ;
  input \pi0920  ;
  input \pi0921  ;
  input \pi0922  ;
  input \pi0923  ;
  input \pi0924  ;
  input \pi0925  ;
  input \pi0926  ;
  input \pi0927  ;
  input \pi0928  ;
  input \pi0929  ;
  input \pi0930  ;
  input \pi0931  ;
  input \pi0932  ;
  input \pi0933  ;
  input \pi0934  ;
  input \pi0935  ;
  input \pi0936  ;
  input \pi0937  ;
  input \pi0938  ;
  input \pi0939  ;
  input \pi0940  ;
  input \pi0941  ;
  input \pi0942  ;
  input \pi0943  ;
  input \pi0944  ;
  input \pi0945  ;
  input \pi0946  ;
  input \pi0947  ;
  input \pi0948  ;
  input \pi0949  ;
  input \pi0950  ;
  input \pi0951  ;
  input \pi0952  ;
  input \pi0953  ;
  input \pi0954  ;
  input \pi0955  ;
  input \pi0956  ;
  input \pi0957  ;
  input \pi0958  ;
  input \pi0959  ;
  input \pi0960  ;
  input \pi0961  ;
  input \pi0962  ;
  input \pi0963  ;
  input \pi0964  ;
  input \pi0965  ;
  input \pi0966  ;
  input \pi0967  ;
  input \pi0968  ;
  input \pi0969  ;
  input \pi0970  ;
  input \pi0971  ;
  input \pi0972  ;
  input \pi0973  ;
  input \pi0974  ;
  input \pi0975  ;
  input \pi0976  ;
  input \pi0977  ;
  input \pi0978  ;
  input \pi0979  ;
  input \pi0980  ;
  input \pi0981  ;
  input \pi0982  ;
  input \pi0983  ;
  input \pi0984  ;
  input \pi0985  ;
  input \pi0986  ;
  input \pi0987  ;
  input \pi0988  ;
  input \pi0989  ;
  input \pi0990  ;
  input \pi0991  ;
  input \pi0992  ;
  input \pi0993  ;
  input \pi0994  ;
  input \pi0995  ;
  input \pi0996  ;
  input \pi0997  ;
  input \pi0998  ;
  input \pi0999  ;
  input \pi1000  ;
  input \pi1001  ;
  input \pi1002  ;
  input \pi1003  ;
  input \pi1004  ;
  input \pi1005  ;
  input \pi1006  ;
  input \pi1007  ;
  input \pi1008  ;
  input \pi1009  ;
  input \pi1010  ;
  input \pi1011  ;
  input \pi1012  ;
  input \pi1013  ;
  input \pi1014  ;
  input \pi1015  ;
  input \pi1016  ;
  input \pi1017  ;
  input \pi1018  ;
  input \pi1019  ;
  input \pi1020  ;
  input \pi1021  ;
  input \pi1022  ;
  input \pi1023  ;
  input \pi1024  ;
  input \pi1025  ;
  input \pi1026  ;
  input \pi1027  ;
  input \pi1028  ;
  input \pi1029  ;
  input \pi1030  ;
  input \pi1031  ;
  input \pi1032  ;
  input \pi1033  ;
  input \pi1034  ;
  input \pi1035  ;
  input \pi1036  ;
  input \pi1037  ;
  input \pi1038  ;
  input \pi1039  ;
  input \pi1040  ;
  input \pi1041  ;
  input \pi1042  ;
  input \pi1043  ;
  input \pi1044  ;
  input \pi1045  ;
  input \pi1046  ;
  input \pi1047  ;
  input \pi1048  ;
  input \pi1049  ;
  input \pi1050  ;
  input \pi1051  ;
  input \pi1052  ;
  input \pi1053  ;
  input \pi1054  ;
  input \pi1055  ;
  input \pi1056  ;
  input \pi1057  ;
  input \pi1058  ;
  input \pi1059  ;
  input \pi1060  ;
  input \pi1061  ;
  input \pi1062  ;
  input \pi1063  ;
  input \pi1064  ;
  input \pi1065  ;
  input \pi1066  ;
  input \pi1067  ;
  input \pi1068  ;
  input \pi1069  ;
  input \pi1070  ;
  input \pi1071  ;
  input \pi1072  ;
  input \pi1073  ;
  input \pi1074  ;
  input \pi1075  ;
  input \pi1076  ;
  input \pi1077  ;
  input \pi1078  ;
  input \pi1079  ;
  input \pi1080  ;
  input \pi1081  ;
  input \pi1082  ;
  input \pi1083  ;
  input \pi1084  ;
  input \pi1085  ;
  input \pi1086  ;
  input \pi1087  ;
  input \pi1088  ;
  input \pi1089  ;
  input \pi1090  ;
  input \pi1091  ;
  input \pi1092  ;
  input \pi1093  ;
  input \pi1094  ;
  input \pi1095  ;
  input \pi1096  ;
  input \pi1097  ;
  input \pi1098  ;
  input \pi1099  ;
  input \pi1100  ;
  input \pi1101  ;
  input \pi1102  ;
  input \pi1103  ;
  input \pi1104  ;
  input \pi1105  ;
  input \pi1106  ;
  input \pi1107  ;
  input \pi1108  ;
  input \pi1109  ;
  input \pi1110  ;
  input \pi1111  ;
  input \pi1112  ;
  input \pi1113  ;
  input \pi1114  ;
  input \pi1115  ;
  input \pi1116  ;
  input \pi1117  ;
  input \pi1118  ;
  input \pi1119  ;
  input \pi1120  ;
  input \pi1121  ;
  input \pi1122  ;
  input \pi1123  ;
  input \pi1124  ;
  input \pi1125  ;
  input \pi1126  ;
  input \pi1127  ;
  input \pi1128  ;
  input \pi1129  ;
  input \pi1130  ;
  input \pi1131  ;
  input \pi1132  ;
  input \pi1133  ;
  input \pi1134  ;
  input \pi1135  ;
  input \pi1136  ;
  input \pi1137  ;
  input \pi1138  ;
  input \pi1139  ;
  input \pi1140  ;
  input \pi1141  ;
  input \pi1142  ;
  input \pi1143  ;
  input \pi1144  ;
  input \pi1145  ;
  input \pi1146  ;
  input \pi1147  ;
  input \pi1148  ;
  input \pi1149  ;
  input \pi1150  ;
  input \pi1151  ;
  input \pi1152  ;
  input \pi1153  ;
  input \pi1154  ;
  input \pi1155  ;
  input \pi1156  ;
  input \pi1157  ;
  input \pi1158  ;
  input \pi1159  ;
  input \pi1160  ;
  input \pi1161  ;
  input \pi1162  ;
  input \pi1163  ;
  input \pi1164  ;
  input \pi1165  ;
  input \pi1166  ;
  input \pi1167  ;
  input \pi1168  ;
  input \pi1169  ;
  input \pi1170  ;
  input \pi1171  ;
  input \pi1172  ;
  input \pi1173  ;
  input \pi1174  ;
  input \pi1175  ;
  input \pi1176  ;
  input \pi1177  ;
  input \pi1178  ;
  input \pi1179  ;
  input \pi1180  ;
  input \pi1181  ;
  input \pi1182  ;
  input \pi1183  ;
  input \pi1184  ;
  input \pi1185  ;
  input \pi1186  ;
  input \pi1187  ;
  input \pi1188  ;
  input \pi1189  ;
  input \pi1190  ;
  input \pi1191  ;
  input \pi1192  ;
  input \pi1193  ;
  input \pi1194  ;
  input \pi1195  ;
  input \pi1196  ;
  input \pi1197  ;
  input \pi1198  ;
  input \pi1199  ;
  input \pi1200  ;
  input \pi1201  ;
  input \pi1202  ;
  input \pi1203  ;
  output \po0000  ;
  output \po0001  ;
  output \po0002  ;
  output \po0003  ;
  output \po0004  ;
  output \po0005  ;
  output \po0006  ;
  output \po0007  ;
  output \po0008  ;
  output \po0009  ;
  output \po0010  ;
  output \po0011  ;
  output \po0012  ;
  output \po0013  ;
  output \po0014  ;
  output \po0015  ;
  output \po0016  ;
  output \po0017  ;
  output \po0018  ;
  output \po0019  ;
  output \po0020  ;
  output \po0021  ;
  output \po0022  ;
  output \po0023  ;
  output \po0024  ;
  output \po0025  ;
  output \po0026  ;
  output \po0027  ;
  output \po0028  ;
  output \po0029  ;
  output \po0030  ;
  output \po0031  ;
  output \po0032  ;
  output \po0033  ;
  output \po0034  ;
  output \po0035  ;
  output \po0036  ;
  output \po0037  ;
  output \po0038  ;
  output \po0039  ;
  output \po0040  ;
  output \po0041  ;
  output \po0042  ;
  output \po0043  ;
  output \po0044  ;
  output \po0045  ;
  output \po0046  ;
  output \po0047  ;
  output \po0048  ;
  output \po0049  ;
  output \po0050  ;
  output \po0051  ;
  output \po0052  ;
  output \po0053  ;
  output \po0054  ;
  output \po0055  ;
  output \po0056  ;
  output \po0057  ;
  output \po0058  ;
  output \po0059  ;
  output \po0060  ;
  output \po0061  ;
  output \po0062  ;
  output \po0063  ;
  output \po0064  ;
  output \po0065  ;
  output \po0066  ;
  output \po0067  ;
  output \po0068  ;
  output \po0069  ;
  output \po0070  ;
  output \po0071  ;
  output \po0072  ;
  output \po0073  ;
  output \po0074  ;
  output \po0075  ;
  output \po0076  ;
  output \po0077  ;
  output \po0078  ;
  output \po0079  ;
  output \po0080  ;
  output \po0081  ;
  output \po0082  ;
  output \po0083  ;
  output \po0084  ;
  output \po0085  ;
  output \po0086  ;
  output \po0087  ;
  output \po0088  ;
  output \po0089  ;
  output \po0090  ;
  output \po0091  ;
  output \po0092  ;
  output \po0093  ;
  output \po0094  ;
  output \po0095  ;
  output \po0096  ;
  output \po0097  ;
  output \po0098  ;
  output \po0099  ;
  output \po0100  ;
  output \po0101  ;
  output \po0102  ;
  output \po0103  ;
  output \po0104  ;
  output \po0105  ;
  output \po0106  ;
  output \po0107  ;
  output \po0108  ;
  output \po0109  ;
  output \po0110  ;
  output \po0111  ;
  output \po0112  ;
  output \po0113  ;
  output \po0114  ;
  output \po0115  ;
  output \po0116  ;
  output \po0117  ;
  output \po0118  ;
  output \po0119  ;
  output \po0120  ;
  output \po0121  ;
  output \po0122  ;
  output \po0123  ;
  output \po0124  ;
  output \po0125  ;
  output \po0126  ;
  output \po0127  ;
  output \po0128  ;
  output \po0129  ;
  output \po0130  ;
  output \po0131  ;
  output \po0132  ;
  output \po0133  ;
  output \po0134  ;
  output \po0135  ;
  output \po0136  ;
  output \po0137  ;
  output \po0138  ;
  output \po0139  ;
  output \po0140  ;
  output \po0141  ;
  output \po0142  ;
  output \po0143  ;
  output \po0144  ;
  output \po0145  ;
  output \po0146  ;
  output \po0147  ;
  output \po0148  ;
  output \po0149  ;
  output \po0150  ;
  output \po0151  ;
  output \po0152  ;
  output \po0153  ;
  output \po0154  ;
  output \po0155  ;
  output \po0156  ;
  output \po0157  ;
  output \po0158  ;
  output \po0159  ;
  output \po0160  ;
  output \po0161  ;
  output \po0162  ;
  output \po0163  ;
  output \po0164  ;
  output \po0165  ;
  output \po0166  ;
  output \po0167  ;
  output \po0168  ;
  output \po0169  ;
  output \po0170  ;
  output \po0171  ;
  output \po0172  ;
  output \po0173  ;
  output \po0174  ;
  output \po0175  ;
  output \po0176  ;
  output \po0177  ;
  output \po0178  ;
  output \po0179  ;
  output \po0180  ;
  output \po0181  ;
  output \po0182  ;
  output \po0183  ;
  output \po0184  ;
  output \po0185  ;
  output \po0186  ;
  output \po0187  ;
  output \po0188  ;
  output \po0189  ;
  output \po0190  ;
  output \po0191  ;
  output \po0192  ;
  output \po0193  ;
  output \po0194  ;
  output \po0195  ;
  output \po0196  ;
  output \po0197  ;
  output \po0198  ;
  output \po0199  ;
  output \po0200  ;
  output \po0201  ;
  output \po0202  ;
  output \po0203  ;
  output \po0204  ;
  output \po0205  ;
  output \po0206  ;
  output \po0207  ;
  output \po0208  ;
  output \po0209  ;
  output \po0210  ;
  output \po0211  ;
  output \po0212  ;
  output \po0213  ;
  output \po0214  ;
  output \po0215  ;
  output \po0216  ;
  output \po0217  ;
  output \po0218  ;
  output \po0219  ;
  output \po0220  ;
  output \po0221  ;
  output \po0222  ;
  output \po0223  ;
  output \po0224  ;
  output \po0225  ;
  output \po0226  ;
  output \po0227  ;
  output \po0228  ;
  output \po0229  ;
  output \po0230  ;
  output \po0231  ;
  output \po0232  ;
  output \po0233  ;
  output \po0234  ;
  output \po0235  ;
  output \po0236  ;
  output \po0237  ;
  output \po0238  ;
  output \po0239  ;
  output \po0240  ;
  output \po0241  ;
  output \po0242  ;
  output \po0243  ;
  output \po0244  ;
  output \po0245  ;
  output \po0246  ;
  output \po0247  ;
  output \po0248  ;
  output \po0249  ;
  output \po0250  ;
  output \po0251  ;
  output \po0252  ;
  output \po0253  ;
  output \po0254  ;
  output \po0255  ;
  output \po0256  ;
  output \po0257  ;
  output \po0258  ;
  output \po0259  ;
  output \po0260  ;
  output \po0261  ;
  output \po0262  ;
  output \po0263  ;
  output \po0264  ;
  output \po0265  ;
  output \po0266  ;
  output \po0267  ;
  output \po0268  ;
  output \po0269  ;
  output \po0270  ;
  output \po0271  ;
  output \po0272  ;
  output \po0273  ;
  output \po0274  ;
  output \po0275  ;
  output \po0276  ;
  output \po0277  ;
  output \po0278  ;
  output \po0279  ;
  output \po0280  ;
  output \po0281  ;
  output \po0282  ;
  output \po0283  ;
  output \po0284  ;
  output \po0285  ;
  output \po0286  ;
  output \po0287  ;
  output \po0288  ;
  output \po0289  ;
  output \po0290  ;
  output \po0291  ;
  output \po0292  ;
  output \po0293  ;
  output \po0294  ;
  output \po0295  ;
  output \po0296  ;
  output \po0297  ;
  output \po0298  ;
  output \po0299  ;
  output \po0300  ;
  output \po0301  ;
  output \po0302  ;
  output \po0303  ;
  output \po0304  ;
  output \po0305  ;
  output \po0306  ;
  output \po0307  ;
  output \po0308  ;
  output \po0309  ;
  output \po0310  ;
  output \po0311  ;
  output \po0312  ;
  output \po0313  ;
  output \po0314  ;
  output \po0315  ;
  output \po0316  ;
  output \po0317  ;
  output \po0318  ;
  output \po0319  ;
  output \po0320  ;
  output \po0321  ;
  output \po0322  ;
  output \po0323  ;
  output \po0324  ;
  output \po0325  ;
  output \po0326  ;
  output \po0327  ;
  output \po0328  ;
  output \po0329  ;
  output \po0330  ;
  output \po0331  ;
  output \po0332  ;
  output \po0333  ;
  output \po0334  ;
  output \po0335  ;
  output \po0336  ;
  output \po0337  ;
  output \po0338  ;
  output \po0339  ;
  output \po0340  ;
  output \po0341  ;
  output \po0342  ;
  output \po0343  ;
  output \po0344  ;
  output \po0345  ;
  output \po0346  ;
  output \po0347  ;
  output \po0348  ;
  output \po0349  ;
  output \po0350  ;
  output \po0351  ;
  output \po0352  ;
  output \po0353  ;
  output \po0354  ;
  output \po0355  ;
  output \po0356  ;
  output \po0357  ;
  output \po0358  ;
  output \po0359  ;
  output \po0360  ;
  output \po0361  ;
  output \po0362  ;
  output \po0363  ;
  output \po0364  ;
  output \po0365  ;
  output \po0366  ;
  output \po0367  ;
  output \po0368  ;
  output \po0369  ;
  output \po0370  ;
  output \po0371  ;
  output \po0372  ;
  output \po0373  ;
  output \po0374  ;
  output \po0375  ;
  output \po0376  ;
  output \po0377  ;
  output \po0378  ;
  output \po0379  ;
  output \po0380  ;
  output \po0381  ;
  output \po0382  ;
  output \po0383  ;
  output \po0384  ;
  output \po0385  ;
  output \po0386  ;
  output \po0387  ;
  output \po0388  ;
  output \po0389  ;
  output \po0390  ;
  output \po0391  ;
  output \po0392  ;
  output \po0393  ;
  output \po0394  ;
  output \po0395  ;
  output \po0396  ;
  output \po0397  ;
  output \po0398  ;
  output \po0399  ;
  output \po0400  ;
  output \po0401  ;
  output \po0402  ;
  output \po0403  ;
  output \po0404  ;
  output \po0405  ;
  output \po0406  ;
  output \po0407  ;
  output \po0408  ;
  output \po0409  ;
  output \po0410  ;
  output \po0411  ;
  output \po0412  ;
  output \po0413  ;
  output \po0414  ;
  output \po0415  ;
  output \po0416  ;
  output \po0417  ;
  output \po0418  ;
  output \po0419  ;
  output \po0420  ;
  output \po0421  ;
  output \po0422  ;
  output \po0423  ;
  output \po0424  ;
  output \po0425  ;
  output \po0426  ;
  output \po0427  ;
  output \po0428  ;
  output \po0429  ;
  output \po0430  ;
  output \po0431  ;
  output \po0432  ;
  output \po0433  ;
  output \po0434  ;
  output \po0435  ;
  output \po0436  ;
  output \po0437  ;
  output \po0438  ;
  output \po0439  ;
  output \po0440  ;
  output \po0441  ;
  output \po0442  ;
  output \po0443  ;
  output \po0444  ;
  output \po0445  ;
  output \po0446  ;
  output \po0447  ;
  output \po0448  ;
  output \po0449  ;
  output \po0450  ;
  output \po0451  ;
  output \po0452  ;
  output \po0453  ;
  output \po0454  ;
  output \po0455  ;
  output \po0456  ;
  output \po0457  ;
  output \po0458  ;
  output \po0459  ;
  output \po0460  ;
  output \po0461  ;
  output \po0462  ;
  output \po0463  ;
  output \po0464  ;
  output \po0465  ;
  output \po0466  ;
  output \po0467  ;
  output \po0468  ;
  output \po0469  ;
  output \po0470  ;
  output \po0471  ;
  output \po0472  ;
  output \po0473  ;
  output \po0474  ;
  output \po0475  ;
  output \po0476  ;
  output \po0477  ;
  output \po0478  ;
  output \po0479  ;
  output \po0480  ;
  output \po0481  ;
  output \po0482  ;
  output \po0483  ;
  output \po0484  ;
  output \po0485  ;
  output \po0486  ;
  output \po0487  ;
  output \po0488  ;
  output \po0489  ;
  output \po0490  ;
  output \po0491  ;
  output \po0492  ;
  output \po0493  ;
  output \po0494  ;
  output \po0495  ;
  output \po0496  ;
  output \po0497  ;
  output \po0498  ;
  output \po0499  ;
  output \po0500  ;
  output \po0501  ;
  output \po0502  ;
  output \po0503  ;
  output \po0504  ;
  output \po0505  ;
  output \po0506  ;
  output \po0507  ;
  output \po0508  ;
  output \po0509  ;
  output \po0510  ;
  output \po0511  ;
  output \po0512  ;
  output \po0513  ;
  output \po0514  ;
  output \po0515  ;
  output \po0516  ;
  output \po0517  ;
  output \po0518  ;
  output \po0519  ;
  output \po0520  ;
  output \po0521  ;
  output \po0522  ;
  output \po0523  ;
  output \po0524  ;
  output \po0525  ;
  output \po0526  ;
  output \po0527  ;
  output \po0528  ;
  output \po0529  ;
  output \po0530  ;
  output \po0531  ;
  output \po0532  ;
  output \po0533  ;
  output \po0534  ;
  output \po0535  ;
  output \po0536  ;
  output \po0537  ;
  output \po0538  ;
  output \po0539  ;
  output \po0540  ;
  output \po0541  ;
  output \po0542  ;
  output \po0543  ;
  output \po0544  ;
  output \po0545  ;
  output \po0546  ;
  output \po0547  ;
  output \po0548  ;
  output \po0549  ;
  output \po0550  ;
  output \po0551  ;
  output \po0552  ;
  output \po0553  ;
  output \po0554  ;
  output \po0555  ;
  output \po0556  ;
  output \po0557  ;
  output \po0558  ;
  output \po0559  ;
  output \po0560  ;
  output \po0561  ;
  output \po0562  ;
  output \po0563  ;
  output \po0564  ;
  output \po0565  ;
  output \po0566  ;
  output \po0567  ;
  output \po0568  ;
  output \po0569  ;
  output \po0570  ;
  output \po0571  ;
  output \po0572  ;
  output \po0573  ;
  output \po0574  ;
  output \po0575  ;
  output \po0576  ;
  output \po0577  ;
  output \po0578  ;
  output \po0579  ;
  output \po0580  ;
  output \po0581  ;
  output \po0582  ;
  output \po0583  ;
  output \po0584  ;
  output \po0585  ;
  output \po0586  ;
  output \po0587  ;
  output \po0588  ;
  output \po0589  ;
  output \po0590  ;
  output \po0591  ;
  output \po0592  ;
  output \po0593  ;
  output \po0594  ;
  output \po0595  ;
  output \po0596  ;
  output \po0597  ;
  output \po0598  ;
  output \po0599  ;
  output \po0600  ;
  output \po0601  ;
  output \po0602  ;
  output \po0603  ;
  output \po0604  ;
  output \po0605  ;
  output \po0606  ;
  output \po0607  ;
  output \po0608  ;
  output \po0609  ;
  output \po0610  ;
  output \po0611  ;
  output \po0612  ;
  output \po0613  ;
  output \po0614  ;
  output \po0615  ;
  output \po0616  ;
  output \po0617  ;
  output \po0618  ;
  output \po0619  ;
  output \po0620  ;
  output \po0621  ;
  output \po0622  ;
  output \po0623  ;
  output \po0624  ;
  output \po0625  ;
  output \po0626  ;
  output \po0627  ;
  output \po0628  ;
  output \po0629  ;
  output \po0630  ;
  output \po0631  ;
  output \po0632  ;
  output \po0633  ;
  output \po0634  ;
  output \po0635  ;
  output \po0636  ;
  output \po0637  ;
  output \po0638  ;
  output \po0639  ;
  output \po0640  ;
  output \po0641  ;
  output \po0642  ;
  output \po0643  ;
  output \po0644  ;
  output \po0645  ;
  output \po0646  ;
  output \po0647  ;
  output \po0648  ;
  output \po0649  ;
  output \po0650  ;
  output \po0651  ;
  output \po0652  ;
  output \po0653  ;
  output \po0654  ;
  output \po0655  ;
  output \po0656  ;
  output \po0657  ;
  output \po0658  ;
  output \po0659  ;
  output \po0660  ;
  output \po0661  ;
  output \po0662  ;
  output \po0663  ;
  output \po0664  ;
  output \po0665  ;
  output \po0666  ;
  output \po0667  ;
  output \po0668  ;
  output \po0669  ;
  output \po0670  ;
  output \po0671  ;
  output \po0672  ;
  output \po0673  ;
  output \po0674  ;
  output \po0675  ;
  output \po0676  ;
  output \po0677  ;
  output \po0678  ;
  output \po0679  ;
  output \po0680  ;
  output \po0681  ;
  output \po0682  ;
  output \po0683  ;
  output \po0684  ;
  output \po0685  ;
  output \po0686  ;
  output \po0687  ;
  output \po0688  ;
  output \po0689  ;
  output \po0690  ;
  output \po0691  ;
  output \po0692  ;
  output \po0693  ;
  output \po0694  ;
  output \po0695  ;
  output \po0696  ;
  output \po0697  ;
  output \po0698  ;
  output \po0699  ;
  output \po0700  ;
  output \po0701  ;
  output \po0702  ;
  output \po0703  ;
  output \po0704  ;
  output \po0705  ;
  output \po0706  ;
  output \po0707  ;
  output \po0708  ;
  output \po0709  ;
  output \po0710  ;
  output \po0711  ;
  output \po0712  ;
  output \po0713  ;
  output \po0714  ;
  output \po0715  ;
  output \po0716  ;
  output \po0717  ;
  output \po0718  ;
  output \po0719  ;
  output \po0720  ;
  output \po0721  ;
  output \po0722  ;
  output \po0723  ;
  output \po0724  ;
  output \po0725  ;
  output \po0726  ;
  output \po0727  ;
  output \po0728  ;
  output \po0729  ;
  output \po0730  ;
  output \po0731  ;
  output \po0732  ;
  output \po0733  ;
  output \po0734  ;
  output \po0735  ;
  output \po0736  ;
  output \po0737  ;
  output \po0738  ;
  output \po0739  ;
  output \po0740  ;
  output \po0741  ;
  output \po0742  ;
  output \po0743  ;
  output \po0744  ;
  output \po0745  ;
  output \po0746  ;
  output \po0747  ;
  output \po0748  ;
  output \po0749  ;
  output \po0750  ;
  output \po0751  ;
  output \po0752  ;
  output \po0753  ;
  output \po0754  ;
  output \po0755  ;
  output \po0756  ;
  output \po0757  ;
  output \po0758  ;
  output \po0759  ;
  output \po0760  ;
  output \po0761  ;
  output \po0762  ;
  output \po0763  ;
  output \po0764  ;
  output \po0765  ;
  output \po0766  ;
  output \po0767  ;
  output \po0768  ;
  output \po0769  ;
  output \po0770  ;
  output \po0771  ;
  output \po0772  ;
  output \po0773  ;
  output \po0774  ;
  output \po0775  ;
  output \po0776  ;
  output \po0777  ;
  output \po0778  ;
  output \po0779  ;
  output \po0780  ;
  output \po0781  ;
  output \po0782  ;
  output \po0783  ;
  output \po0784  ;
  output \po0785  ;
  output \po0786  ;
  output \po0787  ;
  output \po0788  ;
  output \po0789  ;
  output \po0790  ;
  output \po0791  ;
  output \po0792  ;
  output \po0793  ;
  output \po0794  ;
  output \po0795  ;
  output \po0796  ;
  output \po0797  ;
  output \po0798  ;
  output \po0799  ;
  output \po0800  ;
  output \po0801  ;
  output \po0802  ;
  output \po0803  ;
  output \po0804  ;
  output \po0805  ;
  output \po0806  ;
  output \po0807  ;
  output \po0808  ;
  output \po0809  ;
  output \po0810  ;
  output \po0811  ;
  output \po0812  ;
  output \po0813  ;
  output \po0814  ;
  output \po0815  ;
  output \po0816  ;
  output \po0817  ;
  output \po0818  ;
  output \po0819  ;
  output \po0820  ;
  output \po0821  ;
  output \po0822  ;
  output \po0823  ;
  output \po0824  ;
  output \po0825  ;
  output \po0826  ;
  output \po0827  ;
  output \po0828  ;
  output \po0829  ;
  output \po0830  ;
  output \po0831  ;
  output \po0832  ;
  output \po0833  ;
  output \po0834  ;
  output \po0835  ;
  output \po0836  ;
  output \po0837  ;
  output \po0838  ;
  output \po0839  ;
  output \po0840  ;
  output \po0841  ;
  output \po0842  ;
  output \po0843  ;
  output \po0844  ;
  output \po0845  ;
  output \po0846  ;
  output \po0847  ;
  output \po0848  ;
  output \po0849  ;
  output \po0850  ;
  output \po0851  ;
  output \po0852  ;
  output \po0853  ;
  output \po0854  ;
  output \po0855  ;
  output \po0856  ;
  output \po0857  ;
  output \po0858  ;
  output \po0859  ;
  output \po0860  ;
  output \po0861  ;
  output \po0862  ;
  output \po0863  ;
  output \po0864  ;
  output \po0865  ;
  output \po0866  ;
  output \po0867  ;
  output \po0868  ;
  output \po0869  ;
  output \po0870  ;
  output \po0871  ;
  output \po0872  ;
  output \po0873  ;
  output \po0874  ;
  output \po0875  ;
  output \po0876  ;
  output \po0877  ;
  output \po0878  ;
  output \po0879  ;
  output \po0880  ;
  output \po0881  ;
  output \po0882  ;
  output \po0883  ;
  output \po0884  ;
  output \po0885  ;
  output \po0886  ;
  output \po0887  ;
  output \po0888  ;
  output \po0889  ;
  output \po0890  ;
  output \po0891  ;
  output \po0892  ;
  output \po0893  ;
  output \po0894  ;
  output \po0895  ;
  output \po0896  ;
  output \po0897  ;
  output \po0898  ;
  output \po0899  ;
  output \po0900  ;
  output \po0901  ;
  output \po0902  ;
  output \po0903  ;
  output \po0904  ;
  output \po0905  ;
  output \po0906  ;
  output \po0907  ;
  output \po0908  ;
  output \po0909  ;
  output \po0910  ;
  output \po0911  ;
  output \po0912  ;
  output \po0913  ;
  output \po0914  ;
  output \po0915  ;
  output \po0916  ;
  output \po0917  ;
  output \po0918  ;
  output \po0919  ;
  output \po0920  ;
  output \po0921  ;
  output \po0922  ;
  output \po0923  ;
  output \po0924  ;
  output \po0925  ;
  output \po0926  ;
  output \po0927  ;
  output \po0928  ;
  output \po0929  ;
  output \po0930  ;
  output \po0931  ;
  output \po0932  ;
  output \po0933  ;
  output \po0934  ;
  output \po0935  ;
  output \po0936  ;
  output \po0937  ;
  output \po0938  ;
  output \po0939  ;
  output \po0940  ;
  output \po0941  ;
  output \po0942  ;
  output \po0943  ;
  output \po0944  ;
  output \po0945  ;
  output \po0946  ;
  output \po0947  ;
  output \po0948  ;
  output \po0949  ;
  output \po0950  ;
  output \po0951  ;
  output \po0952  ;
  output \po0953  ;
  output \po0954  ;
  output \po0955  ;
  output \po0956  ;
  output \po0957  ;
  output \po0958  ;
  output \po0959  ;
  output \po0960  ;
  output \po0961  ;
  output \po0962  ;
  output \po0963  ;
  output \po0964  ;
  output \po0965  ;
  output \po0966  ;
  output \po0967  ;
  output \po0968  ;
  output \po0969  ;
  output \po0970  ;
  output \po0971  ;
  output \po0972  ;
  output \po0973  ;
  output \po0974  ;
  output \po0975  ;
  output \po0976  ;
  output \po0977  ;
  output \po0978  ;
  output \po0979  ;
  output \po0980  ;
  output \po0981  ;
  output \po0982  ;
  output \po0983  ;
  output \po0984  ;
  output \po0985  ;
  output \po0986  ;
  output \po0987  ;
  output \po0988  ;
  output \po0989  ;
  output \po0990  ;
  output \po0991  ;
  output \po0992  ;
  output \po0993  ;
  output \po0994  ;
  output \po0995  ;
  output \po0996  ;
  output \po0997  ;
  output \po0998  ;
  output \po0999  ;
  output \po1000  ;
  output \po1001  ;
  output \po1002  ;
  output \po1003  ;
  output \po1004  ;
  output \po1005  ;
  output \po1006  ;
  output \po1007  ;
  output \po1008  ;
  output \po1009  ;
  output \po1010  ;
  output \po1011  ;
  output \po1012  ;
  output \po1013  ;
  output \po1014  ;
  output \po1015  ;
  output \po1016  ;
  output \po1017  ;
  output \po1018  ;
  output \po1019  ;
  output \po1020  ;
  output \po1021  ;
  output \po1022  ;
  output \po1023  ;
  output \po1024  ;
  output \po1025  ;
  output \po1026  ;
  output \po1027  ;
  output \po1028  ;
  output \po1029  ;
  output \po1030  ;
  output \po1031  ;
  output \po1032  ;
  output \po1033  ;
  output \po1034  ;
  output \po1035  ;
  output \po1036  ;
  output \po1037  ;
  output \po1038  ;
  output \po1039  ;
  output \po1040  ;
  output \po1041  ;
  output \po1042  ;
  output \po1043  ;
  output \po1044  ;
  output \po1045  ;
  output \po1046  ;
  output \po1047  ;
  output \po1048  ;
  output \po1049  ;
  output \po1050  ;
  output \po1051  ;
  output \po1052  ;
  output \po1053  ;
  output \po1054  ;
  output \po1055  ;
  output \po1056  ;
  output \po1057  ;
  output \po1058  ;
  output \po1059  ;
  output \po1060  ;
  output \po1061  ;
  output \po1062  ;
  output \po1063  ;
  output \po1064  ;
  output \po1065  ;
  output \po1066  ;
  output \po1067  ;
  output \po1068  ;
  output \po1069  ;
  output \po1070  ;
  output \po1071  ;
  output \po1072  ;
  output \po1073  ;
  output \po1074  ;
  output \po1075  ;
  output \po1076  ;
  output \po1077  ;
  output \po1078  ;
  output \po1079  ;
  output \po1080  ;
  output \po1081  ;
  output \po1082  ;
  output \po1083  ;
  output \po1084  ;
  output \po1085  ;
  output \po1086  ;
  output \po1087  ;
  output \po1088  ;
  output \po1089  ;
  output \po1090  ;
  output \po1091  ;
  output \po1092  ;
  output \po1093  ;
  output \po1094  ;
  output \po1095  ;
  output \po1096  ;
  output \po1097  ;
  output \po1098  ;
  output \po1099  ;
  output \po1100  ;
  output \po1101  ;
  output \po1102  ;
  output \po1103  ;
  output \po1104  ;
  output \po1105  ;
  output \po1106  ;
  output \po1107  ;
  output \po1108  ;
  output \po1109  ;
  output \po1110  ;
  output \po1111  ;
  output \po1112  ;
  output \po1113  ;
  output \po1114  ;
  output \po1115  ;
  output \po1116  ;
  output \po1117  ;
  output \po1118  ;
  output \po1119  ;
  output \po1120  ;
  output \po1121  ;
  output \po1122  ;
  output \po1123  ;
  output \po1124  ;
  output \po1125  ;
  output \po1126  ;
  output \po1127  ;
  output \po1128  ;
  output \po1129  ;
  output \po1130  ;
  output \po1131  ;
  output \po1132  ;
  output \po1133  ;
  output \po1134  ;
  output \po1135  ;
  output \po1136  ;
  output \po1137  ;
  output \po1138  ;
  output \po1139  ;
  output \po1140  ;
  output \po1141  ;
  output \po1142  ;
  output \po1143  ;
  output \po1144  ;
  output \po1145  ;
  output \po1146  ;
  output \po1147  ;
  output \po1148  ;
  output \po1149  ;
  output \po1150  ;
  output \po1151  ;
  output \po1152  ;
  output \po1153  ;
  output \po1154  ;
  output \po1155  ;
  output \po1156  ;
  output \po1157  ;
  output \po1158  ;
  output \po1159  ;
  output \po1160  ;
  output \po1161  ;
  output \po1162  ;
  output \po1163  ;
  output \po1164  ;
  output \po1165  ;
  output \po1166  ;
  output \po1167  ;
  output \po1168  ;
  output \po1169  ;
  output \po1170  ;
  output \po1171  ;
  output \po1172  ;
  output \po1173  ;
  output \po1174  ;
  output \po1175  ;
  output \po1176  ;
  output \po1177  ;
  output \po1178  ;
  output \po1179  ;
  output \po1180  ;
  output \po1181  ;
  output \po1182  ;
  output \po1183  ;
  output \po1184  ;
  output \po1185  ;
  output \po1186  ;
  output \po1187  ;
  output \po1188  ;
  output \po1189  ;
  output \po1190  ;
  output \po1191  ;
  output \po1192  ;
  output \po1193  ;
  output \po1194  ;
  output \po1195  ;
  output \po1196  ;
  output \po1197  ;
  output \po1198  ;
  output \po1199  ;
  output \po1200  ;
  output \po1201  ;
  output \po1202  ;
  output \po1203  ;
  output \po1204  ;
  output \po1205  ;
  output \po1206  ;
  output \po1207  ;
  output \po1208  ;
  output \po1209  ;
  output \po1210  ;
  output \po1211  ;
  output \po1212  ;
  output \po1213  ;
  output \po1214  ;
  output \po1215  ;
  output \po1216  ;
  output \po1217  ;
  output \po1218  ;
  output \po1219  ;
  output \po1220  ;
  output \po1221  ;
  output \po1222  ;
  output \po1223  ;
  output \po1224  ;
  output \po1225  ;
  output \po1226  ;
  output \po1227  ;
  output \po1228  ;
  output \po1229  ;
  output \po1230  ;
  wire n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , n64765 , n64766 ;
  assign n1205 = ~\pi0332  & ~\pi1144  ;
  assign n1206 = \pi0215  & ~n1205 ;
  assign n1207 = \pi0095  & \pi0234  ;
  assign n1208 = ~\pi0479  & n1207 ;
  assign n1209 = \pi0105  & \pi0228  ;
  assign n1210 = ~\pi0332  & n1209 ;
  assign n1211 = ~n1208 & n1210 ;
  assign n1212 = \pi0153  & ~\pi0332  ;
  assign n1213 = ~n1209 & n1212 ;
  assign n1214 = ~\pi0216  & ~n1213 ;
  assign n1215 = ~n1211 & n1214 ;
  assign n1216 = \pi0265  & ~\pi0332  ;
  assign n1217 = \pi0216  & ~n1216 ;
  assign n1218 = ~\pi0221  & ~n1217 ;
  assign n1219 = ~n1215 & n1218 ;
  assign n1220 = ~\pi0216  & \pi0833  ;
  assign n1221 = n1205 & ~n1220 ;
  assign n1222 = ~\pi0332  & ~\pi0929  ;
  assign n1223 = n1220 & n1222 ;
  assign n1224 = ~n1221 & ~n1223 ;
  assign n1225 = \pi0221  & ~n1224 ;
  assign n1226 = ~\pi0215  & ~n1225 ;
  assign n1227 = ~n1219 & n1226 ;
  assign n1228 = ~n1206 & ~n1227 ;
  assign n1229 = \pi0057  & ~n1228 ;
  assign n1230 = ~\pi0332  & ~n1208 ;
  assign n1231 = ~\pi0082  & ~\pi0111  ;
  assign n1232 = ~\pi0036  & n1231 ;
  assign n1233 = ~\pi0068  & ~\pi0084  ;
  assign n1234 = ~\pi0066  & ~\pi0073  ;
  assign n1235 = n1233 & n1234 ;
  assign n1236 = n1232 & n1235 ;
  assign n1237 = ~\pi0061  & ~\pi0076  ;
  assign n1238 = ~\pi0085  & ~\pi0106  ;
  assign n1239 = n1237 & n1238 ;
  assign n1240 = ~\pi0048  & ~\pi0089  ;
  assign n1241 = ~\pi0049  & n1240 ;
  assign n1242 = n1239 & n1241 ;
  assign n1243 = ~\pi0045  & ~\pi0104  ;
  assign n1244 = ~\pi0083  & ~\pi0103  ;
  assign n1245 = ~\pi0067  & ~\pi0069  ;
  assign n1246 = n1244 & n1245 ;
  assign n1247 = n1243 & n1246 ;
  assign n1248 = n1242 & n1247 ;
  assign n1249 = n1236 & n1248 ;
  assign n1250 = ~\pi0064  & ~\pi0102  ;
  assign n1251 = ~\pi0081  & n1250 ;
  assign n1252 = ~\pi0050  & ~\pi0077  ;
  assign n1253 = ~\pi0088  & ~\pi0098  ;
  assign n1254 = n1252 & n1253 ;
  assign n1255 = n1251 & n1254 ;
  assign n1256 = ~\pi0063  & ~\pi0107  ;
  assign n1257 = ~\pi0065  & ~\pi0071  ;
  assign n1258 = n1256 & n1257 ;
  assign n1259 = n1255 & n1258 ;
  assign n1260 = n1249 & n1259 ;
  assign n1261 = ~\pi0035  & ~\pi0051  ;
  assign n1262 = ~\pi0072  & ~\pi0096  ;
  assign n1263 = ~\pi0040  & n1262 ;
  assign n1264 = ~\pi0032  & ~\pi0095  ;
  assign n1265 = ~\pi0070  & n1264 ;
  assign n1266 = n1263 & n1265 ;
  assign n1267 = n1261 & n1266 ;
  assign n1268 = ~\pi0046  & ~\pi0097  ;
  assign n1269 = ~\pi0108  & n1268 ;
  assign n1270 = ~\pi0109  & ~\pi0110  ;
  assign n1271 = ~\pi0047  & ~\pi0091  ;
  assign n1272 = n1270 & n1271 ;
  assign n1273 = n1269 & n1272 ;
  assign n1274 = ~\pi0086  & ~\pi0094  ;
  assign n1275 = ~\pi0053  & ~\pi0060  ;
  assign n1276 = n1274 & n1275 ;
  assign n1277 = ~\pi0058  & ~\pi0090  ;
  assign n1278 = ~\pi0093  & n1277 ;
  assign n1279 = n1276 & n1278 ;
  assign n1280 = n1273 & n1279 ;
  assign n1281 = n1267 & n1280 ;
  assign n1282 = \pi0137  & n1281 ;
  assign n1283 = n1260 & n1282 ;
  assign n1284 = n1230 & ~n1283 ;
  assign n1285 = ~\pi0054  & ~\pi0092  ;
  assign n1286 = ~\pi0075  & ~\pi0087  ;
  assign n1287 = n1285 & n1286 ;
  assign n1288 = ~\pi0038  & ~\pi0039  ;
  assign n1289 = ~\pi0074  & ~\pi0100  ;
  assign n1290 = n1288 & n1289 ;
  assign n1291 = n1287 & n1290 ;
  assign n1292 = ~\pi0056  & ~\pi0062  ;
  assign n1293 = ~\pi0055  & n1292 ;
  assign n1294 = n1291 & n1293 ;
  assign n1295 = ~\pi0215  & ~\pi0221  ;
  assign n1296 = ~\pi0059  & ~\pi0216  ;
  assign n1297 = n1295 & n1296 ;
  assign n1298 = ~n1213 & n1297 ;
  assign n1299 = n1294 & n1298 ;
  assign n1300 = \pi0057  & n1299 ;
  assign n1301 = ~n1284 & n1300 ;
  assign n1302 = ~n1229 & ~n1301 ;
  assign n1303 = ~\pi0216  & n1295 ;
  assign n1304 = ~n1213 & n1303 ;
  assign n1305 = n1294 & n1304 ;
  assign n1306 = ~n1284 & n1305 ;
  assign n1307 = \pi0059  & ~n1206 ;
  assign n1308 = ~n1227 & n1307 ;
  assign n1309 = ~n1306 & n1308 ;
  assign n1310 = ~\pi0057  & ~n1309 ;
  assign n1311 = n1302 & ~n1310 ;
  assign n1312 = ~\pi0234  & ~\pi0332  ;
  assign n1313 = \pi0095  & ~\pi0137  ;
  assign n1314 = n1255 & n1257 ;
  assign n1315 = n1269 & n1276 ;
  assign n1316 = n1314 & n1315 ;
  assign n1317 = n1236 & n1256 ;
  assign n1318 = n1248 & n1317 ;
  assign n1319 = n1316 & n1318 ;
  assign n1320 = ~\pi0090  & ~\pi0093  ;
  assign n1321 = ~\pi0035  & ~\pi0070  ;
  assign n1322 = n1320 & n1321 ;
  assign n1323 = ~\pi0051  & ~\pi0096  ;
  assign n1324 = n1322 & n1323 ;
  assign n1325 = ~\pi0047  & ~\pi0110  ;
  assign n1326 = ~\pi0058  & ~\pi0091  ;
  assign n1327 = n1325 & n1326 ;
  assign n1328 = ~\pi0109  & n1327 ;
  assign n1329 = ~\pi0040  & ~\pi0072  ;
  assign n1330 = \pi0225  & n1329 ;
  assign n1331 = n1328 & n1330 ;
  assign n1332 = n1324 & n1331 ;
  assign n1333 = n1319 & n1332 ;
  assign n1334 = \pi0032  & ~\pi0137  ;
  assign n1335 = ~n1333 & n1334 ;
  assign n1336 = ~n1313 & ~n1335 ;
  assign n1337 = \pi0210  & ~n1336 ;
  assign n1338 = ~\pi0060  & n1257 ;
  assign n1339 = n1256 & n1338 ;
  assign n1340 = n1255 & n1339 ;
  assign n1341 = \pi0053  & n1274 ;
  assign n1342 = n1340 & n1341 ;
  assign n1343 = n1249 & n1342 ;
  assign n1344 = ~\pi0053  & n1274 ;
  assign n1345 = \pi0060  & n1257 ;
  assign n1346 = n1256 & n1345 ;
  assign n1347 = n1255 & n1346 ;
  assign n1348 = n1344 & n1347 ;
  assign n1349 = n1249 & n1348 ;
  assign n1350 = ~n1343 & ~n1349 ;
  assign n1351 = n1273 & n1278 ;
  assign n1352 = ~n1350 & n1351 ;
  assign n1353 = ~\pi0035  & ~n1352 ;
  assign n1354 = n1256 & n1278 ;
  assign n1355 = n1255 & n1338 ;
  assign n1356 = n1273 & n1344 ;
  assign n1357 = n1355 & n1356 ;
  assign n1358 = n1249 & n1357 ;
  assign n1359 = n1354 & n1358 ;
  assign n1360 = \pi0035  & ~n1359 ;
  assign n1361 = \pi0035  & ~\pi0225  ;
  assign n1362 = n1354 & n1361 ;
  assign n1363 = n1358 & n1362 ;
  assign n1364 = ~\pi0051  & ~\pi0070  ;
  assign n1365 = n1263 & n1364 ;
  assign n1366 = ~n1363 & n1365 ;
  assign n1367 = ~n1360 & n1366 ;
  assign n1368 = ~n1353 & n1367 ;
  assign n1369 = ~\pi0032  & ~\pi0137  ;
  assign n1370 = \pi0210  & n1369 ;
  assign n1371 = ~n1368 & n1370 ;
  assign n1372 = ~n1337 & ~n1371 ;
  assign n1373 = \pi0225  & n1354 ;
  assign n1374 = n1358 & n1373 ;
  assign n1375 = \pi0035  & ~n1374 ;
  assign n1376 = ~\pi0070  & ~\pi0096  ;
  assign n1377 = ~\pi0035  & n1354 ;
  assign n1378 = n1358 & n1377 ;
  assign n1379 = \pi0051  & ~n1378 ;
  assign n1380 = n1376 & ~n1379 ;
  assign n1381 = \pi0093  & n1277 ;
  assign n1382 = n1256 & n1381 ;
  assign n1383 = n1358 & n1382 ;
  assign n1384 = ~\pi0035  & ~n1383 ;
  assign n1385 = n1380 & ~n1384 ;
  assign n1386 = \pi0047  & n1257 ;
  assign n1387 = n1256 & n1386 ;
  assign n1388 = n1255 & n1387 ;
  assign n1389 = n1270 & n1315 ;
  assign n1390 = n1388 & n1389 ;
  assign n1391 = n1249 & n1390 ;
  assign n1392 = \pi0047  & ~n1391 ;
  assign n1393 = ~\pi0091  & ~\pi0110  ;
  assign n1394 = ~\pi0091  & ~\pi0109  ;
  assign n1395 = n1319 & n1394 ;
  assign n1396 = ~n1393 & ~n1395 ;
  assign n1397 = ~n1392 & ~n1396 ;
  assign n1398 = \pi0091  & ~\pi0109  ;
  assign n1399 = n1325 & n1398 ;
  assign n1400 = n1319 & n1399 ;
  assign n1401 = n1277 & ~n1400 ;
  assign n1402 = ~n1397 & n1401 ;
  assign n1403 = ~\pi0065  & n1236 ;
  assign n1404 = n1248 & n1403 ;
  assign n1405 = ~n1257 & ~n1404 ;
  assign n1406 = \pi0065  & ~\pi0071  ;
  assign n1407 = n1236 & n1406 ;
  assign n1408 = n1248 & n1407 ;
  assign n1409 = ~\pi0107  & ~n1408 ;
  assign n1410 = n1405 & n1409 ;
  assign n1411 = n1235 & n1243 ;
  assign n1412 = n1242 & n1411 ;
  assign n1413 = \pi0111  & ~n1412 ;
  assign n1414 = ~\pi0082  & ~n1413 ;
  assign n1415 = ~\pi0084  & n1234 ;
  assign n1416 = n1243 & n1415 ;
  assign n1417 = n1242 & n1416 ;
  assign n1418 = \pi0068  & ~n1417 ;
  assign n1419 = n1414 & ~n1418 ;
  assign n1420 = ~\pi0068  & ~\pi0111  ;
  assign n1421 = \pi0082  & n1420 ;
  assign n1422 = n1417 & n1421 ;
  assign n1423 = ~\pi0069  & ~\pi0083  ;
  assign n1424 = ~\pi0036  & ~\pi0067  ;
  assign n1425 = n1423 & n1424 ;
  assign n1426 = ~n1422 & n1425 ;
  assign n1427 = ~n1419 & n1426 ;
  assign n1428 = \pi0085  & \pi0106  ;
  assign n1429 = n1237 & ~n1428 ;
  assign n1430 = \pi0061  & \pi0076  ;
  assign n1431 = n1238 & ~n1430 ;
  assign n1432 = ~n1429 & ~n1431 ;
  assign n1433 = ~\pi0048  & ~n1432 ;
  assign n1434 = ~n1239 & ~n1433 ;
  assign n1435 = n1239 & n1240 ;
  assign n1436 = ~\pi0049  & ~\pi0089  ;
  assign n1437 = ~\pi0048  & ~\pi0049  ;
  assign n1438 = n1239 & n1437 ;
  assign n1439 = ~n1436 & ~n1438 ;
  assign n1440 = ~n1435 & n1439 ;
  assign n1441 = \pi0104  & ~n1242 ;
  assign n1442 = ~\pi0049  & ~\pi0104  ;
  assign n1443 = n1240 & n1442 ;
  assign n1444 = n1239 & n1443 ;
  assign n1445 = ~\pi0045  & ~n1444 ;
  assign n1446 = ~n1441 & n1445 ;
  assign n1447 = ~n1440 & n1446 ;
  assign n1448 = ~n1434 & n1447 ;
  assign n1449 = ~n1243 & n1444 ;
  assign n1450 = n1415 & ~n1449 ;
  assign n1451 = ~n1448 & n1450 ;
  assign n1452 = \pi0066  & \pi0073  ;
  assign n1453 = n1234 & ~n1452 ;
  assign n1454 = n1243 & ~n1452 ;
  assign n1455 = n1242 & n1454 ;
  assign n1456 = ~n1453 & ~n1455 ;
  assign n1457 = ~\pi0084  & n1456 ;
  assign n1458 = n1234 & n1243 ;
  assign n1459 = n1242 & n1458 ;
  assign n1460 = \pi0084  & ~n1459 ;
  assign n1461 = ~n1457 & ~n1460 ;
  assign n1462 = ~n1451 & n1461 ;
  assign n1463 = n1420 & n1426 ;
  assign n1464 = ~n1462 & n1463 ;
  assign n1465 = ~n1427 & ~n1464 ;
  assign n1466 = n1231 & n1233 ;
  assign n1467 = n1458 & n1466 ;
  assign n1468 = n1242 & n1467 ;
  assign n1469 = \pi0036  & ~n1468 ;
  assign n1470 = n1423 & n1469 ;
  assign n1471 = n1242 & n1243 ;
  assign n1472 = n1236 & n1471 ;
  assign n1473 = \pi0067  & n1423 ;
  assign n1474 = ~n1472 & n1473 ;
  assign n1475 = ~n1470 & ~n1474 ;
  assign n1476 = n1231 & n1424 ;
  assign n1477 = n1235 & n1476 ;
  assign n1478 = n1471 & n1477 ;
  assign n1479 = \pi0069  & ~n1478 ;
  assign n1480 = n1236 & n1245 ;
  assign n1481 = n1471 & n1480 ;
  assign n1482 = \pi0083  & ~n1481 ;
  assign n1483 = ~\pi0103  & ~n1482 ;
  assign n1484 = ~n1479 & n1483 ;
  assign n1485 = n1475 & n1484 ;
  assign n1486 = n1465 & n1485 ;
  assign n1487 = ~\pi0083  & \pi0103  ;
  assign n1488 = n1243 & n1487 ;
  assign n1489 = n1242 & n1488 ;
  assign n1490 = n1480 & n1489 ;
  assign n1491 = ~\pi0071  & ~n1490 ;
  assign n1492 = n1409 & n1491 ;
  assign n1493 = ~n1486 & n1492 ;
  assign n1494 = ~n1410 & ~n1493 ;
  assign n1495 = n1236 & n1258 ;
  assign n1496 = n1248 & n1495 ;
  assign n1497 = \pi0064  & ~n1496 ;
  assign n1498 = ~\pi0063  & n1257 ;
  assign n1499 = n1236 & n1498 ;
  assign n1500 = n1248 & n1499 ;
  assign n1501 = ~n1256 & ~n1500 ;
  assign n1502 = ~n1497 & ~n1501 ;
  assign n1503 = n1494 & n1502 ;
  assign n1504 = ~\pi0081  & ~\pi0102  ;
  assign n1505 = \pi0064  & n1258 ;
  assign n1506 = n1236 & n1505 ;
  assign n1507 = n1248 & n1506 ;
  assign n1508 = n1504 & ~n1507 ;
  assign n1509 = ~n1503 & n1508 ;
  assign n1510 = \pi0063  & ~\pi0107  ;
  assign n1511 = n1257 & n1510 ;
  assign n1512 = n1236 & n1511 ;
  assign n1513 = n1248 & n1512 ;
  assign n1514 = ~\pi0064  & ~n1513 ;
  assign n1515 = n1405 & n1514 ;
  assign n1516 = n1491 & n1514 ;
  assign n1517 = ~n1486 & n1516 ;
  assign n1518 = ~n1515 & ~n1517 ;
  assign n1519 = ~\pi0107  & ~n1518 ;
  assign n1520 = n1501 & n1514 ;
  assign n1521 = ~n1497 & ~n1520 ;
  assign n1522 = ~n1519 & n1521 ;
  assign n1523 = n1253 & ~n1522 ;
  assign n1524 = n1509 & n1523 ;
  assign n1525 = ~\pi0064  & n1256 ;
  assign n1526 = n1257 & n1525 ;
  assign n1527 = n1236 & n1526 ;
  assign n1528 = n1248 & n1527 ;
  assign n1529 = \pi0081  & ~n1528 ;
  assign n1530 = ~\pi0064  & ~\pi0081  ;
  assign n1531 = n1256 & n1530 ;
  assign n1532 = n1257 & n1531 ;
  assign n1533 = n1236 & n1532 ;
  assign n1534 = n1248 & n1533 ;
  assign n1535 = \pi0102  & ~n1534 ;
  assign n1536 = ~n1529 & ~n1535 ;
  assign n1537 = n1253 & ~n1536 ;
  assign n1538 = ~\pi0050  & ~\pi0060  ;
  assign n1539 = ~\pi0102  & n1257 ;
  assign n1540 = n1531 & n1539 ;
  assign n1541 = n1236 & n1540 ;
  assign n1542 = n1248 & n1541 ;
  assign n1543 = ~\pi0077  & n1253 ;
  assign n1544 = ~\pi0060  & n1543 ;
  assign n1545 = n1542 & n1544 ;
  assign n1546 = ~n1538 & ~n1545 ;
  assign n1547 = ~\pi0098  & n1542 ;
  assign n1548 = \pi0088  & ~n1547 ;
  assign n1549 = \pi0098  & ~n1542 ;
  assign n1550 = ~\pi0077  & ~n1549 ;
  assign n1551 = ~n1548 & n1550 ;
  assign n1552 = ~n1546 & n1551 ;
  assign n1553 = ~n1537 & n1552 ;
  assign n1554 = ~n1524 & n1553 ;
  assign n1555 = \pi0077  & n1253 ;
  assign n1556 = n1542 & n1555 ;
  assign n1557 = ~\pi0050  & ~n1556 ;
  assign n1558 = ~n1546 & ~n1557 ;
  assign n1559 = n1249 & n1347 ;
  assign n1560 = ~\pi0053  & ~\pi0086  ;
  assign n1561 = ~n1559 & n1560 ;
  assign n1562 = ~n1558 & n1561 ;
  assign n1563 = ~n1554 & n1562 ;
  assign n1564 = n1249 & n1340 ;
  assign n1565 = \pi0053  & ~\pi0086  ;
  assign n1566 = ~n1564 & n1565 ;
  assign n1567 = ~\pi0050  & n1275 ;
  assign n1568 = n1543 & n1567 ;
  assign n1569 = n1274 & n1568 ;
  assign n1570 = n1542 & n1569 ;
  assign n1571 = \pi0097  & ~n1570 ;
  assign n1572 = ~\pi0094  & n1568 ;
  assign n1573 = n1542 & n1572 ;
  assign n1574 = ~n1274 & ~n1573 ;
  assign n1575 = ~n1571 & ~n1574 ;
  assign n1576 = ~n1566 & n1575 ;
  assign n1577 = ~n1563 & n1576 ;
  assign n1578 = ~\pi0086  & \pi0094  ;
  assign n1579 = n1568 & n1578 ;
  assign n1580 = n1542 & n1579 ;
  assign n1581 = ~\pi0097  & ~n1580 ;
  assign n1582 = ~n1571 & ~n1581 ;
  assign n1583 = ~\pi0108  & n1274 ;
  assign n1584 = \pi0046  & n1583 ;
  assign n1585 = n1568 & n1584 ;
  assign n1586 = n1542 & n1585 ;
  assign n1587 = ~\pi0097  & n1586 ;
  assign n1588 = ~\pi0108  & ~\pi0109  ;
  assign n1589 = ~n1587 & n1588 ;
  assign n1590 = ~n1582 & n1589 ;
  assign n1591 = ~n1577 & n1590 ;
  assign n1592 = ~\pi0097  & n1274 ;
  assign n1593 = n1568 & n1592 ;
  assign n1594 = n1542 & n1593 ;
  assign n1595 = \pi0108  & ~n1594 ;
  assign n1596 = ~\pi0046  & ~n1595 ;
  assign n1597 = ~\pi0109  & ~n1587 ;
  assign n1598 = ~n1596 & n1597 ;
  assign n1599 = \pi0109  & ~n1319 ;
  assign n1600 = ~n1598 & ~n1599 ;
  assign n1601 = ~n1591 & n1600 ;
  assign n1602 = n1325 & n1401 ;
  assign n1603 = ~n1601 & n1602 ;
  assign n1604 = ~n1402 & ~n1603 ;
  assign n1605 = n1256 & n1358 ;
  assign n1606 = \pi0058  & ~n1605 ;
  assign n1607 = ~\pi0093  & n1328 ;
  assign n1608 = n1319 & n1607 ;
  assign n1609 = ~n1320 & ~n1608 ;
  assign n1610 = ~n1606 & ~n1609 ;
  assign n1611 = n1380 & n1610 ;
  assign n1612 = n1604 & n1611 ;
  assign n1613 = ~n1385 & ~n1612 ;
  assign n1614 = ~n1375 & ~n1613 ;
  assign n1615 = \pi0051  & n1376 ;
  assign n1616 = n1378 & n1615 ;
  assign n1617 = ~\pi0035  & \pi0040  ;
  assign n1618 = n1262 & n1364 ;
  assign n1619 = n1617 & n1618 ;
  assign n1620 = n1354 & n1619 ;
  assign n1621 = n1358 & n1620 ;
  assign n1622 = ~\pi0032  & ~\pi0072  ;
  assign n1623 = ~n1621 & n1622 ;
  assign n1624 = ~n1616 & n1623 ;
  assign n1625 = ~n1614 & n1624 ;
  assign n1626 = ~\pi0032  & ~n1621 ;
  assign n1627 = n1324 & n1328 ;
  assign n1628 = n1319 & n1627 ;
  assign n1629 = \pi0072  & ~n1628 ;
  assign n1630 = ~\pi0040  & ~n1629 ;
  assign n1631 = n1626 & ~n1630 ;
  assign n1632 = \pi0032  & ~n1333 ;
  assign n1633 = \pi0095  & ~\pi0479  ;
  assign n1634 = ~\pi0032  & ~\pi0040  ;
  assign n1635 = ~\pi0035  & n1634 ;
  assign n1636 = n1618 & n1635 ;
  assign n1637 = n1354 & n1636 ;
  assign n1638 = n1358 & n1637 ;
  assign n1639 = \pi0095  & ~n1638 ;
  assign n1640 = ~n1633 & ~n1639 ;
  assign n1641 = ~n1632 & n1640 ;
  assign n1642 = ~n1631 & n1641 ;
  assign n1643 = ~n1625 & n1642 ;
  assign n1644 = \pi0095  & \pi0479  ;
  assign n1645 = n1638 & n1644 ;
  assign n1646 = \pi0137  & \pi0210  ;
  assign n1647 = ~n1645 & n1646 ;
  assign n1648 = ~n1643 & n1647 ;
  assign n1649 = n1372 & ~n1648 ;
  assign n1650 = \pi0841  & n1329 ;
  assign n1651 = n1261 & n1376 ;
  assign n1652 = n1650 & n1651 ;
  assign n1653 = n1373 & n1652 ;
  assign n1654 = n1358 & n1653 ;
  assign n1655 = \pi0032  & ~n1654 ;
  assign n1656 = n1640 & ~n1655 ;
  assign n1657 = ~n1631 & n1656 ;
  assign n1658 = ~n1625 & n1657 ;
  assign n1659 = \pi0137  & ~\pi0210  ;
  assign n1660 = ~n1645 & n1659 ;
  assign n1661 = ~n1658 & n1660 ;
  assign n1662 = ~\pi0095  & \pi0225  ;
  assign n1663 = n1652 & n1662 ;
  assign n1664 = n1354 & n1663 ;
  assign n1665 = n1358 & n1664 ;
  assign n1666 = ~\pi0137  & ~n1264 ;
  assign n1667 = ~n1665 & n1666 ;
  assign n1668 = ~\pi0210  & n1667 ;
  assign n1669 = ~\pi0210  & n1369 ;
  assign n1670 = ~n1368 & n1669 ;
  assign n1671 = ~n1668 & ~n1670 ;
  assign n1672 = ~\pi0146  & n1671 ;
  assign n1673 = ~n1661 & n1672 ;
  assign n1674 = n1649 & n1673 ;
  assign n1675 = n1568 & n1583 ;
  assign n1676 = n1542 & n1675 ;
  assign n1677 = ~\pi0097  & ~\pi0108  ;
  assign n1678 = ~n1676 & ~n1677 ;
  assign n1679 = ~\pi0110  & ~n1678 ;
  assign n1680 = ~\pi0097  & n1350 ;
  assign n1681 = ~\pi0046  & ~\pi0109  ;
  assign n1682 = n1271 & n1681 ;
  assign n1683 = n1278 & n1682 ;
  assign n1684 = ~n1680 & n1683 ;
  assign n1685 = n1679 & n1684 ;
  assign n1686 = ~\pi0833  & \pi0957  ;
  assign n1687 = \pi0829  & \pi0950  ;
  assign n1688 = ~n1686 & n1687 ;
  assign n1689 = \pi1092  & \pi1093  ;
  assign n1690 = ~\pi0035  & \pi1091  ;
  assign n1691 = n1689 & n1690 ;
  assign n1692 = n1688 & n1691 ;
  assign n1693 = ~n1685 & n1692 ;
  assign n1694 = ~n1264 & ~n1665 ;
  assign n1695 = \pi1091  & n1689 ;
  assign n1696 = n1688 & n1695 ;
  assign n1697 = ~\pi0035  & ~n1696 ;
  assign n1698 = ~n1352 & n1697 ;
  assign n1699 = n1367 & ~n1698 ;
  assign n1700 = ~n1694 & n1699 ;
  assign n1701 = ~n1693 & n1700 ;
  assign n1702 = \pi0032  & n1665 ;
  assign n1703 = ~\pi0137  & ~\pi0210  ;
  assign n1704 = ~n1702 & n1703 ;
  assign n1705 = ~n1701 & n1704 ;
  assign n1706 = \pi0146  & ~n1705 ;
  assign n1707 = ~n1661 & n1706 ;
  assign n1708 = n1649 & n1707 ;
  assign n1709 = ~n1674 & ~n1708 ;
  assign n1710 = n1312 & n1709 ;
  assign n1711 = ~n1363 & n1364 ;
  assign n1712 = ~n1360 & n1711 ;
  assign n1713 = ~n1353 & n1712 ;
  assign n1714 = ~\pi0032  & ~\pi0096  ;
  assign n1715 = ~n1713 & n1714 ;
  assign n1716 = ~\pi0096  & n1329 ;
  assign n1717 = ~\pi0109  & n1325 ;
  assign n1718 = ~\pi0035  & n1320 ;
  assign n1719 = n1326 & n1364 ;
  assign n1720 = n1718 & n1719 ;
  assign n1721 = n1717 & n1720 ;
  assign n1722 = n1329 & n1721 ;
  assign n1723 = n1319 & n1722 ;
  assign n1724 = ~n1716 & ~n1723 ;
  assign n1725 = ~\pi0032  & n1724 ;
  assign n1726 = ~n1644 & ~n1655 ;
  assign n1727 = ~n1725 & n1726 ;
  assign n1728 = ~n1715 & n1727 ;
  assign n1729 = ~\pi0137  & ~n1633 ;
  assign n1730 = ~n1728 & n1729 ;
  assign n1731 = ~\pi0137  & ~n1730 ;
  assign n1732 = \pi0096  & n1329 ;
  assign n1733 = n1721 & n1732 ;
  assign n1734 = n1319 & n1733 ;
  assign n1735 = n1261 & n1354 ;
  assign n1736 = n1358 & n1735 ;
  assign n1737 = n1734 & n1736 ;
  assign n1738 = ~\pi0095  & ~n1737 ;
  assign n1739 = \pi0032  & ~\pi0095  ;
  assign n1740 = ~n1654 & n1739 ;
  assign n1741 = ~n1738 & ~n1740 ;
  assign n1742 = ~n1631 & ~n1740 ;
  assign n1743 = ~n1625 & n1742 ;
  assign n1744 = ~n1741 & ~n1743 ;
  assign n1745 = ~n1638 & n1644 ;
  assign n1746 = ~n1730 & ~n1745 ;
  assign n1747 = ~n1744 & n1746 ;
  assign n1748 = ~n1731 & ~n1747 ;
  assign n1749 = ~\pi0146  & ~\pi0210  ;
  assign n1750 = ~n1748 & n1749 ;
  assign n1751 = ~\pi0095  & ~n1632 ;
  assign n1752 = ~n1725 & n1751 ;
  assign n1753 = ~n1715 & n1752 ;
  assign n1754 = n1729 & ~n1753 ;
  assign n1755 = ~\pi0137  & ~n1754 ;
  assign n1756 = ~\pi0146  & \pi0210  ;
  assign n1757 = n1755 & n1756 ;
  assign n1758 = ~n1333 & n1739 ;
  assign n1759 = ~n1738 & ~n1758 ;
  assign n1760 = ~n1631 & ~n1758 ;
  assign n1761 = ~n1625 & n1760 ;
  assign n1762 = ~n1759 & ~n1761 ;
  assign n1763 = ~n1745 & ~n1754 ;
  assign n1764 = n1756 & n1763 ;
  assign n1765 = ~n1762 & n1764 ;
  assign n1766 = ~n1757 & ~n1765 ;
  assign n1767 = ~n1750 & n1766 ;
  assign n1768 = \pi0234  & ~\pi0332  ;
  assign n1769 = \pi0146  & ~\pi0210  ;
  assign n1770 = ~\pi0035  & ~\pi0096  ;
  assign n1771 = ~n1685 & n1770 ;
  assign n1772 = ~\pi0096  & ~n1712 ;
  assign n1773 = ~n1655 & ~n1724 ;
  assign n1774 = ~n1772 & n1773 ;
  assign n1775 = ~n1771 & n1774 ;
  assign n1776 = \pi0032  & n1654 ;
  assign n1777 = ~\pi0095  & ~n1776 ;
  assign n1778 = ~n1775 & n1777 ;
  assign n1779 = ~n1644 & n1696 ;
  assign n1780 = ~n1778 & n1779 ;
  assign n1781 = ~\pi0137  & n1696 ;
  assign n1782 = ~n1730 & ~n1781 ;
  assign n1783 = ~n1780 & ~n1782 ;
  assign n1784 = ~\pi0137  & ~n1783 ;
  assign n1785 = n1769 & n1784 ;
  assign n1786 = ~n1745 & ~n1783 ;
  assign n1787 = n1769 & n1786 ;
  assign n1788 = ~n1744 & n1787 ;
  assign n1789 = ~n1785 & ~n1788 ;
  assign n1790 = \pi0146  & \pi0210  ;
  assign n1791 = n1755 & n1790 ;
  assign n1792 = n1763 & n1790 ;
  assign n1793 = ~n1762 & n1792 ;
  assign n1794 = ~n1791 & ~n1793 ;
  assign n1795 = n1789 & n1794 ;
  assign n1796 = n1768 & n1795 ;
  assign n1797 = n1767 & n1796 ;
  assign n1798 = ~n1710 & ~n1797 ;
  assign n1799 = ~\pi0105  & ~n1212 ;
  assign n1800 = ~\pi0152  & ~\pi0161  ;
  assign n1801 = ~\pi0166  & n1800 ;
  assign n1802 = ~n1799 & ~n1801 ;
  assign n1803 = ~n1798 & n1802 ;
  assign n1804 = ~\pi0210  & \pi0234  ;
  assign n1805 = n1784 & n1804 ;
  assign n1806 = n1786 & n1804 ;
  assign n1807 = ~n1744 & n1806 ;
  assign n1808 = ~n1805 & ~n1807 ;
  assign n1809 = \pi0210  & \pi0234  ;
  assign n1810 = n1755 & n1809 ;
  assign n1811 = n1763 & n1809 ;
  assign n1812 = ~n1762 & n1811 ;
  assign n1813 = ~n1810 & ~n1812 ;
  assign n1814 = n1808 & n1813 ;
  assign n1815 = ~\pi0234  & ~n1705 ;
  assign n1816 = ~n1661 & n1815 ;
  assign n1817 = n1649 & n1816 ;
  assign n1818 = ~\pi0166  & ~\pi0332  ;
  assign n1819 = n1800 & n1818 ;
  assign n1820 = ~n1817 & n1819 ;
  assign n1821 = n1814 & n1820 ;
  assign n1822 = \pi0105  & ~n1821 ;
  assign n1823 = ~n1799 & ~n1822 ;
  assign n1824 = ~\pi0216  & \pi0228  ;
  assign n1825 = ~n1823 & n1824 ;
  assign n1826 = ~n1803 & n1825 ;
  assign n1827 = \pi0221  & n1224 ;
  assign n1828 = ~n1217 & ~n1827 ;
  assign n1829 = n1256 & n1277 ;
  assign n1830 = n1358 & n1829 ;
  assign n1831 = \pi0093  & ~n1830 ;
  assign n1832 = ~\pi0035  & ~n1831 ;
  assign n1833 = ~\pi0072  & n1364 ;
  assign n1834 = ~n1363 & n1833 ;
  assign n1835 = ~n1832 & n1834 ;
  assign n1836 = \pi0086  & ~\pi0094  ;
  assign n1837 = n1568 & n1836 ;
  assign n1838 = n1542 & n1837 ;
  assign n1839 = ~\pi0053  & ~n1574 ;
  assign n1840 = ~n1838 & ~n1839 ;
  assign n1841 = ~n1558 & ~n1838 ;
  assign n1842 = ~n1554 & n1841 ;
  assign n1843 = ~n1840 & ~n1842 ;
  assign n1844 = ~n1580 & n1677 ;
  assign n1845 = ~n1843 & n1844 ;
  assign n1846 = \pi0097  & ~\pi0108  ;
  assign n1847 = ~n1570 & n1846 ;
  assign n1848 = n1596 & ~n1599 ;
  assign n1849 = ~n1847 & n1848 ;
  assign n1850 = ~n1845 & n1849 ;
  assign n1851 = \pi0109  & n1319 ;
  assign n1852 = n1277 & n1325 ;
  assign n1853 = ~n1400 & n1852 ;
  assign n1854 = ~n1851 & n1853 ;
  assign n1855 = ~n1850 & n1854 ;
  assign n1856 = n1319 & n1328 ;
  assign n1857 = \pi0090  & ~n1856 ;
  assign n1858 = ~n1606 & ~n1857 ;
  assign n1859 = ~n1402 & n1858 ;
  assign n1860 = ~n1855 & n1859 ;
  assign n1861 = ~\pi0093  & n1834 ;
  assign n1862 = ~n1860 & n1861 ;
  assign n1863 = ~n1835 & ~n1862 ;
  assign n1864 = \pi0070  & ~n1378 ;
  assign n1865 = ~\pi0096  & n1321 ;
  assign n1866 = n1354 & n1865 ;
  assign n1867 = n1358 & n1866 ;
  assign n1868 = ~n1323 & ~n1867 ;
  assign n1869 = ~n1864 & ~n1868 ;
  assign n1870 = ~\pi0072  & ~n1869 ;
  assign n1871 = n1630 & ~n1870 ;
  assign n1872 = n1863 & n1871 ;
  assign n1873 = ~\pi0032  & ~n1696 ;
  assign n1874 = ~n1621 & n1873 ;
  assign n1875 = ~n1872 & n1874 ;
  assign n1876 = \pi0225  & \pi0841  ;
  assign n1877 = n1328 & ~n1876 ;
  assign n1878 = n1324 & n1877 ;
  assign n1879 = n1319 & n1878 ;
  assign n1880 = n1329 & n1879 ;
  assign n1881 = \pi0032  & ~n1880 ;
  assign n1882 = ~\pi0032  & \pi1091  ;
  assign n1883 = n1689 & n1882 ;
  assign n1884 = n1688 & n1883 ;
  assign n1885 = ~n1621 & n1884 ;
  assign n1886 = ~n1881 & ~n1885 ;
  assign n1887 = n1832 & n1858 ;
  assign n1888 = ~n1402 & ~n1854 ;
  assign n1889 = ~\pi0108  & ~n1580 ;
  assign n1890 = ~n1843 & n1889 ;
  assign n1891 = ~n1846 & ~n1890 ;
  assign n1892 = ~n1402 & n1848 ;
  assign n1893 = n1891 & n1892 ;
  assign n1894 = ~n1888 & ~n1893 ;
  assign n1895 = n1887 & ~n1894 ;
  assign n1896 = ~\pi0035  & \pi0093  ;
  assign n1897 = n1830 & n1896 ;
  assign n1898 = n1834 & ~n1897 ;
  assign n1899 = ~n1895 & n1898 ;
  assign n1900 = n1630 & ~n1881 ;
  assign n1901 = ~n1870 & n1900 ;
  assign n1902 = ~n1899 & n1901 ;
  assign n1903 = ~n1886 & ~n1902 ;
  assign n1904 = ~n1875 & ~n1903 ;
  assign n1905 = ~\pi0095  & ~\pi0137  ;
  assign n1906 = ~n1904 & n1905 ;
  assign n1907 = ~\pi0095  & n1329 ;
  assign n1908 = n1879 & n1907 ;
  assign n1909 = ~n1264 & ~n1908 ;
  assign n1910 = \pi0137  & n1909 ;
  assign n1911 = n1323 & ~n1864 ;
  assign n1912 = ~\pi0070  & ~n1363 ;
  assign n1913 = n1329 & ~n1912 ;
  assign n1914 = n1911 & n1913 ;
  assign n1915 = ~\pi0032  & \pi0137  ;
  assign n1916 = ~n1914 & n1915 ;
  assign n1917 = ~n1910 & ~n1916 ;
  assign n1918 = ~\pi0137  & n1633 ;
  assign n1919 = n1313 & ~n1638 ;
  assign n1920 = ~n1918 & ~n1919 ;
  assign n1921 = n1917 & n1920 ;
  assign n1922 = ~n1906 & n1921 ;
  assign n1923 = n1769 & ~n1922 ;
  assign n1924 = ~\pi0225  & n1329 ;
  assign n1925 = n1328 & n1924 ;
  assign n1926 = n1324 & n1925 ;
  assign n1927 = n1319 & n1926 ;
  assign n1928 = \pi0032  & ~n1927 ;
  assign n1929 = n1630 & ~n1928 ;
  assign n1930 = ~n1870 & n1929 ;
  assign n1931 = n1863 & n1930 ;
  assign n1932 = ~n1626 & ~n1928 ;
  assign n1933 = ~\pi0095  & \pi0137  ;
  assign n1934 = \pi0210  & ~n1933 ;
  assign n1935 = \pi0032  & \pi0210  ;
  assign n1936 = ~n1927 & n1935 ;
  assign n1937 = ~n1934 & ~n1936 ;
  assign n1938 = ~\pi0032  & \pi0210  ;
  assign n1939 = ~n1914 & n1938 ;
  assign n1940 = n1937 & ~n1939 ;
  assign n1941 = ~\pi0095  & ~n1940 ;
  assign n1942 = ~n1932 & n1941 ;
  assign n1943 = ~n1931 & n1942 ;
  assign n1944 = ~n1639 & n1729 ;
  assign n1945 = n1768 & n1944 ;
  assign n1946 = n1768 & n1937 ;
  assign n1947 = ~n1939 & n1946 ;
  assign n1948 = ~n1945 & ~n1947 ;
  assign n1949 = ~n1943 & ~n1948 ;
  assign n1950 = n1863 & n1901 ;
  assign n1951 = ~\pi0032  & n1621 ;
  assign n1952 = \pi0032  & n1329 ;
  assign n1953 = n1879 & n1952 ;
  assign n1954 = ~n1951 & ~n1953 ;
  assign n1955 = n1905 & n1954 ;
  assign n1956 = ~n1950 & n1955 ;
  assign n1957 = n1921 & ~n1956 ;
  assign n1958 = n1749 & ~n1957 ;
  assign n1959 = n1949 & ~n1958 ;
  assign n1960 = ~n1923 & n1959 ;
  assign n1961 = \pi0096  & n1721 ;
  assign n1962 = n1319 & n1961 ;
  assign n1963 = ~\pi0072  & ~n1962 ;
  assign n1964 = n1711 & n1963 ;
  assign n1965 = ~n1832 & n1964 ;
  assign n1966 = ~\pi0093  & n1964 ;
  assign n1967 = ~n1860 & n1966 ;
  assign n1968 = ~n1965 & ~n1967 ;
  assign n1969 = ~n1869 & n1963 ;
  assign n1970 = n1929 & ~n1969 ;
  assign n1971 = n1968 & n1970 ;
  assign n1972 = ~n1928 & n1933 ;
  assign n1973 = \pi0210  & ~n1972 ;
  assign n1974 = ~\pi0032  & ~n1734 ;
  assign n1975 = \pi0210  & n1974 ;
  assign n1976 = ~n1914 & n1975 ;
  assign n1977 = ~n1973 & ~n1976 ;
  assign n1978 = ~\pi0032  & n1633 ;
  assign n1979 = n1618 & n1978 ;
  assign n1980 = ~\pi0035  & ~\pi0040  ;
  assign n1981 = n1979 & n1980 ;
  assign n1982 = n1354 & n1981 ;
  assign n1983 = n1358 & n1982 ;
  assign n1984 = \pi0137  & n1983 ;
  assign n1985 = ~\pi0095  & ~n1984 ;
  assign n1986 = ~n1932 & n1985 ;
  assign n1987 = ~n1977 & n1986 ;
  assign n1988 = ~n1971 & n1987 ;
  assign n1989 = ~\pi0137  & ~n1639 ;
  assign n1990 = ~n1984 & ~n1989 ;
  assign n1991 = ~n1977 & n1990 ;
  assign n1992 = n1312 & ~n1991 ;
  assign n1993 = ~n1988 & n1992 ;
  assign n1994 = \pi0137  & ~n1983 ;
  assign n1995 = n1909 & n1994 ;
  assign n1996 = n1974 & n1994 ;
  assign n1997 = ~n1914 & n1996 ;
  assign n1998 = ~n1995 & ~n1997 ;
  assign n1999 = ~n1919 & n1998 ;
  assign n2000 = n1900 & ~n1969 ;
  assign n2001 = n1968 & n2000 ;
  assign n2002 = n1955 & ~n2001 ;
  assign n2003 = n1999 & ~n2002 ;
  assign n2004 = n1749 & ~n2003 ;
  assign n2005 = n1993 & ~n2004 ;
  assign n2006 = ~n1801 & ~n2005 ;
  assign n2007 = n1630 & ~n1969 ;
  assign n2008 = n1968 & n2007 ;
  assign n2009 = n1874 & ~n2008 ;
  assign n2010 = ~n1897 & n1964 ;
  assign n2011 = ~n1895 & n2010 ;
  assign n2012 = n2000 & ~n2011 ;
  assign n2013 = ~n1886 & ~n2012 ;
  assign n2014 = ~n2009 & ~n2013 ;
  assign n2015 = n1905 & ~n2014 ;
  assign n2016 = n1999 & ~n2015 ;
  assign n2017 = n1769 & ~n1801 ;
  assign n2018 = ~n2016 & n2017 ;
  assign n2019 = ~n2006 & ~n2018 ;
  assign n2020 = ~n1960 & ~n2019 ;
  assign n2021 = ~\pi0210  & ~n2016 ;
  assign n2022 = n1993 & ~n2021 ;
  assign n2023 = n1801 & ~n1949 ;
  assign n2024 = ~\pi0166  & ~\pi0210  ;
  assign n2025 = n1800 & n2024 ;
  assign n2026 = ~n1922 & n2025 ;
  assign n2027 = ~n2023 & ~n2026 ;
  assign n2028 = ~n2022 & ~n2027 ;
  assign n2029 = ~\pi0153  & ~n2028 ;
  assign n2030 = ~n2020 & n2029 ;
  assign n2031 = ~n1582 & n1588 ;
  assign n2032 = ~n1577 & n2031 ;
  assign n2033 = ~n1392 & ~n1599 ;
  assign n2034 = ~n1396 & n2033 ;
  assign n2035 = \pi0046  & ~\pi0109  ;
  assign n2036 = \pi0108  & ~\pi0109  ;
  assign n2037 = ~n1594 & n2036 ;
  assign n2038 = ~n2035 & ~n2037 ;
  assign n2039 = n2034 & n2038 ;
  assign n2040 = ~n2032 & n2039 ;
  assign n2041 = n1384 & n1401 ;
  assign n2042 = ~n1325 & ~n1392 ;
  assign n2043 = ~n1396 & n2042 ;
  assign n2044 = n2041 & ~n2043 ;
  assign n2045 = ~n2040 & n2044 ;
  assign n2046 = ~n1360 & ~n1363 ;
  assign n2047 = n1380 & n2046 ;
  assign n2048 = n1384 & ~n1610 ;
  assign n2049 = n2047 & ~n2048 ;
  assign n2050 = ~n2045 & n2049 ;
  assign n2051 = n1624 & ~n2050 ;
  assign n2052 = n1760 & ~n2051 ;
  assign n2053 = ~n1759 & ~n2052 ;
  assign n2054 = \pi0137  & ~n1639 ;
  assign n2055 = ~n2053 & n2054 ;
  assign n2056 = n1752 & n1989 ;
  assign n2057 = ~n1715 & n2056 ;
  assign n2058 = n1638 & n1918 ;
  assign n2059 = n1809 & ~n2058 ;
  assign n2060 = ~n2057 & n2059 ;
  assign n2061 = ~n2055 & n2060 ;
  assign n2062 = n1212 & n2061 ;
  assign n2063 = \pi0032  & n1933 ;
  assign n2064 = ~n1654 & n2063 ;
  assign n2065 = ~n1737 & n1933 ;
  assign n2066 = ~n2064 & ~n2065 ;
  assign n2067 = ~n1631 & ~n2064 ;
  assign n2068 = ~n2051 & n2067 ;
  assign n2069 = ~n2066 & ~n2068 ;
  assign n2070 = ~\pi0146  & ~n1801 ;
  assign n2071 = n1696 & ~n2070 ;
  assign n2072 = ~n1644 & n2071 ;
  assign n2073 = ~n1778 & n2072 ;
  assign n2074 = ~\pi0137  & n2071 ;
  assign n2075 = ~n1730 & ~n2074 ;
  assign n2076 = ~n2073 & ~n2075 ;
  assign n2077 = \pi0234  & ~n1639 ;
  assign n2078 = ~n2076 & n2077 ;
  assign n2079 = ~n2069 & n2078 ;
  assign n2080 = ~n1809 & ~n2079 ;
  assign n2081 = ~\pi0210  & ~\pi0234  ;
  assign n2082 = n1667 & n2070 ;
  assign n2083 = n1369 & n2070 ;
  assign n2084 = ~n1368 & n2083 ;
  assign n2085 = ~n2082 & ~n2084 ;
  assign n2086 = n2081 & n2085 ;
  assign n2087 = n1632 & ~n2086 ;
  assign n2088 = ~n1368 & n1369 ;
  assign n2089 = \pi0210  & n1333 ;
  assign n2090 = n1336 & n2089 ;
  assign n2091 = ~n2088 & n2090 ;
  assign n2092 = n1655 & ~n2091 ;
  assign n2093 = n1640 & ~n2092 ;
  assign n2094 = ~n2087 & n2093 ;
  assign n2095 = ~n1631 & n2094 ;
  assign n2096 = ~n2051 & n2095 ;
  assign n2097 = \pi0137  & ~n1645 ;
  assign n2098 = ~n2096 & n2097 ;
  assign n2099 = \pi0210  & n1336 ;
  assign n2100 = ~n2088 & n2099 ;
  assign n2101 = ~\pi0137  & \pi0146  ;
  assign n2102 = ~\pi0137  & ~\pi0166  ;
  assign n2103 = n1800 & n2102 ;
  assign n2104 = ~n2101 & ~n2103 ;
  assign n2105 = ~n1702 & ~n2104 ;
  assign n2106 = ~n1701 & n2105 ;
  assign n2107 = n2086 & ~n2106 ;
  assign n2108 = ~n2100 & ~n2107 ;
  assign n2109 = ~n2098 & ~n2108 ;
  assign n2110 = n1212 & ~n2109 ;
  assign n2111 = n2080 & n2110 ;
  assign n2112 = ~n2062 & ~n2111 ;
  assign n2113 = ~\pi0228  & n2112 ;
  assign n2114 = ~\pi0216  & n2113 ;
  assign n2115 = ~n2030 & n2114 ;
  assign n2116 = n1828 & ~n2115 ;
  assign n2117 = ~n1826 & n2116 ;
  assign n2118 = ~\pi0142  & ~\pi0198  ;
  assign n2119 = ~n1748 & n2118 ;
  assign n2120 = ~\pi0142  & \pi0198  ;
  assign n2121 = n1755 & n2120 ;
  assign n2122 = n1763 & n2120 ;
  assign n2123 = ~n1762 & n2122 ;
  assign n2124 = ~n2121 & ~n2123 ;
  assign n2125 = ~n2119 & n2124 ;
  assign n2126 = \pi0142  & ~\pi0198  ;
  assign n2127 = n1784 & n2126 ;
  assign n2128 = n1786 & n2126 ;
  assign n2129 = ~n1744 & n2128 ;
  assign n2130 = ~n2127 & ~n2129 ;
  assign n2131 = \pi0142  & \pi0198  ;
  assign n2132 = n1755 & n2131 ;
  assign n2133 = n1763 & n2131 ;
  assign n2134 = ~n1762 & n2133 ;
  assign n2135 = ~n2132 & ~n2134 ;
  assign n2136 = n2130 & n2135 ;
  assign n2137 = n1768 & n2136 ;
  assign n2138 = n2125 & n2137 ;
  assign n2139 = \pi0198  & ~n1336 ;
  assign n2140 = \pi0198  & n1369 ;
  assign n2141 = ~n1368 & n2140 ;
  assign n2142 = ~n2139 & ~n2141 ;
  assign n2143 = \pi0137  & \pi0198  ;
  assign n2144 = ~n1645 & n2143 ;
  assign n2145 = ~n1643 & n2144 ;
  assign n2146 = n2142 & ~n2145 ;
  assign n2147 = \pi0137  & ~\pi0198  ;
  assign n2148 = ~n1645 & n2147 ;
  assign n2149 = ~n1658 & n2148 ;
  assign n2150 = ~\pi0198  & n1667 ;
  assign n2151 = ~\pi0198  & n1369 ;
  assign n2152 = ~n1368 & n2151 ;
  assign n2153 = ~n2150 & ~n2152 ;
  assign n2154 = ~\pi0142  & n2153 ;
  assign n2155 = ~n2149 & n2154 ;
  assign n2156 = n2146 & n2155 ;
  assign n2157 = ~\pi0137  & ~\pi0198  ;
  assign n2158 = ~n1702 & n2157 ;
  assign n2159 = ~n1701 & n2158 ;
  assign n2160 = \pi0142  & ~n2159 ;
  assign n2161 = ~n2149 & n2160 ;
  assign n2162 = n2146 & n2161 ;
  assign n2163 = ~n2156 & ~n2162 ;
  assign n2164 = n1312 & n2163 ;
  assign n2165 = ~\pi0222  & ~\pi0224  ;
  assign n2166 = ~\pi0144  & ~\pi0174  ;
  assign n2167 = ~\pi0189  & n2166 ;
  assign n2168 = ~\pi0223  & ~n2167 ;
  assign n2169 = n2165 & n2168 ;
  assign n2170 = ~n2164 & n2169 ;
  assign n2171 = ~n2138 & n2170 ;
  assign n2172 = ~\pi0198  & \pi0234  ;
  assign n2173 = n1784 & n2172 ;
  assign n2174 = n1786 & n2172 ;
  assign n2175 = ~n1744 & n2174 ;
  assign n2176 = ~n2173 & ~n2175 ;
  assign n2177 = \pi0198  & \pi0234  ;
  assign n2178 = n1755 & n2177 ;
  assign n2179 = n1763 & n2177 ;
  assign n2180 = ~n1762 & n2179 ;
  assign n2181 = ~n2178 & ~n2180 ;
  assign n2182 = n2176 & n2181 ;
  assign n2183 = ~\pi0234  & ~n2159 ;
  assign n2184 = ~n2149 & n2183 ;
  assign n2185 = n2146 & n2184 ;
  assign n2186 = ~\pi0332  & ~n2185 ;
  assign n2187 = n2182 & n2186 ;
  assign n2188 = ~\pi0189  & ~\pi0223  ;
  assign n2189 = n2165 & n2188 ;
  assign n2190 = n2166 & n2189 ;
  assign n2191 = ~n2187 & n2190 ;
  assign n2192 = ~\pi0224  & \pi0833  ;
  assign n2193 = \pi0222  & ~n2192 ;
  assign n2194 = ~\pi0223  & ~n2193 ;
  assign n2195 = n1205 & ~n2194 ;
  assign n2196 = ~\pi0223  & n2192 ;
  assign n2197 = n1222 & n2196 ;
  assign n2198 = \pi0224  & ~n1216 ;
  assign n2199 = ~\pi0222  & ~\pi0223  ;
  assign n2200 = ~n2198 & n2199 ;
  assign n2201 = ~n2197 & ~n2200 ;
  assign n2202 = ~n2195 & n2201 ;
  assign n2203 = ~\pi0299  & ~n2202 ;
  assign n2204 = ~n2191 & n2203 ;
  assign n2205 = ~n2171 & n2204 ;
  assign n2206 = ~\pi0039  & ~\pi0215  ;
  assign n2207 = ~n1225 & n2206 ;
  assign n2208 = ~n2205 & n2207 ;
  assign n2209 = ~n2117 & n2208 ;
  assign n2210 = \pi0299  & ~n1206 ;
  assign n2211 = ~\pi0039  & ~n2210 ;
  assign n2212 = ~n2205 & n2211 ;
  assign n2213 = ~n1227 & n2210 ;
  assign n2214 = ~\pi0223  & n2165 ;
  assign n2215 = ~\pi0299  & ~n2214 ;
  assign n2216 = ~\pi0299  & ~\pi0332  ;
  assign n2217 = ~n1208 & n2216 ;
  assign n2218 = ~n2215 & ~n2217 ;
  assign n2219 = ~n2202 & ~n2218 ;
  assign n2220 = \pi0100  & ~n2219 ;
  assign n2221 = ~n2213 & n2220 ;
  assign n2222 = \pi0100  & n1288 ;
  assign n2223 = ~\pi0087  & ~n2222 ;
  assign n2224 = ~n2221 & n2223 ;
  assign n2225 = ~\pi0105  & \pi0228  ;
  assign n2226 = n1212 & n2225 ;
  assign n2227 = ~n1769 & ~n2025 ;
  assign n2228 = ~\pi0137  & ~n1207 ;
  assign n2229 = n2227 & n2228 ;
  assign n2230 = n1208 & ~n2229 ;
  assign n2231 = n1281 & ~n2229 ;
  assign n2232 = n1260 & n2231 ;
  assign n2233 = ~n2230 & ~n2232 ;
  assign n2234 = \pi0228  & ~\pi0332  ;
  assign n2235 = ~n1799 & n2234 ;
  assign n2236 = n2233 & n2235 ;
  assign n2237 = ~n2226 & ~n2236 ;
  assign n2238 = \pi0146  & \pi0252  ;
  assign n2239 = ~\pi0166  & \pi0252  ;
  assign n2240 = n1800 & n2239 ;
  assign n2241 = ~n2238 & ~n2240 ;
  assign n2242 = n1281 & n2241 ;
  assign n2243 = n1260 & n2242 ;
  assign n2244 = ~\pi0153  & ~n2243 ;
  assign n2245 = ~\pi0228  & ~\pi0332  ;
  assign n2246 = ~\pi0137  & ~n1769 ;
  assign n2247 = ~n2025 & n2246 ;
  assign n2248 = n2241 & ~n2247 ;
  assign n2249 = n1281 & n2248 ;
  assign n2250 = n1260 & n2249 ;
  assign n2251 = n2245 & ~n2250 ;
  assign n2252 = ~n2244 & n2251 ;
  assign n2253 = ~\pi0216  & ~n2252 ;
  assign n2254 = n2237 & n2253 ;
  assign n2255 = n1828 & ~n2254 ;
  assign n2256 = ~\pi0215  & \pi0299  ;
  assign n2257 = ~n1225 & n2256 ;
  assign n2258 = ~n2255 & n2257 ;
  assign n2259 = \pi0215  & \pi0299  ;
  assign n2260 = ~n1205 & n2259 ;
  assign n2261 = ~n2202 & ~n2214 ;
  assign n2262 = ~\pi0299  & ~n2261 ;
  assign n2263 = ~\pi0087  & ~n2262 ;
  assign n2264 = n1207 & n2167 ;
  assign n2265 = ~\pi0189  & ~\pi0198  ;
  assign n2266 = n2166 & n2265 ;
  assign n2267 = ~\pi0137  & ~n2126 ;
  assign n2268 = ~n2266 & n2267 ;
  assign n2269 = ~n2264 & n2268 ;
  assign n2270 = n1281 & ~n2269 ;
  assign n2271 = n1260 & n2270 ;
  assign n2272 = n1230 & ~n2202 ;
  assign n2273 = ~\pi0087  & n2272 ;
  assign n2274 = ~n2271 & n2273 ;
  assign n2275 = ~n2263 & ~n2274 ;
  assign n2276 = n1288 & ~n2275 ;
  assign n2277 = ~n2260 & n2276 ;
  assign n2278 = ~n2258 & n2277 ;
  assign n2279 = ~n2224 & ~n2278 ;
  assign n2280 = n1260 & n1281 ;
  assign n2281 = ~\pi0153  & ~n2280 ;
  assign n2282 = ~n1283 & n2245 ;
  assign n2283 = ~n2281 & n2282 ;
  assign n2284 = \pi0228  & ~n1799 ;
  assign n2285 = n1230 & n2284 ;
  assign n2286 = ~n1283 & n2285 ;
  assign n2287 = ~\pi0221  & ~n2226 ;
  assign n2288 = ~\pi0216  & n2287 ;
  assign n2289 = ~n2286 & n2288 ;
  assign n2290 = ~n2283 & n2289 ;
  assign n2291 = \pi0216  & ~\pi0221  ;
  assign n2292 = ~n1216 & n2291 ;
  assign n2293 = ~n1206 & ~n1827 ;
  assign n2294 = ~n2292 & n2293 ;
  assign n2295 = ~n2290 & n2294 ;
  assign n2296 = \pi0215  & n1205 ;
  assign n2297 = \pi0039  & \pi0299  ;
  assign n2298 = ~n2296 & n2297 ;
  assign n2299 = ~n2295 & n2298 ;
  assign n2300 = ~n1283 & n2272 ;
  assign n2301 = \pi0039  & n2262 ;
  assign n2302 = ~n2300 & n2301 ;
  assign n2303 = ~\pi0038  & ~n2302 ;
  assign n2304 = ~n2299 & n2303 ;
  assign n2305 = ~n2279 & n2304 ;
  assign n2306 = ~n2212 & n2305 ;
  assign n2307 = ~n2209 & n2306 ;
  assign n2308 = \pi0039  & ~n2219 ;
  assign n2309 = ~n2213 & n2308 ;
  assign n2310 = \pi0038  & ~n2309 ;
  assign n2311 = ~\pi0100  & ~n2310 ;
  assign n2312 = n2262 & ~n2300 ;
  assign n2313 = \pi0299  & ~n1228 ;
  assign n2314 = ~\pi0216  & \pi0299  ;
  assign n2315 = n1295 & n2314 ;
  assign n2316 = ~n1213 & n2315 ;
  assign n2317 = ~n1284 & n2316 ;
  assign n2318 = ~n2313 & ~n2317 ;
  assign n2319 = ~n2312 & n2318 ;
  assign n2320 = ~\pi0039  & ~\pi0100  ;
  assign n2321 = ~n2319 & n2320 ;
  assign n2322 = ~n2311 & ~n2321 ;
  assign n2323 = ~n2279 & n2322 ;
  assign n2324 = ~\pi0092  & n1286 ;
  assign n2325 = \pi0299  & ~n2296 ;
  assign n2326 = ~n2295 & n2325 ;
  assign n2327 = ~\pi0038  & ~\pi0100  ;
  assign n2328 = ~\pi0039  & n2327 ;
  assign n2329 = ~n2312 & n2328 ;
  assign n2330 = ~n2326 & n2329 ;
  assign n2331 = n2219 & ~n2328 ;
  assign n2332 = n2210 & ~n2328 ;
  assign n2333 = ~n1227 & n2332 ;
  assign n2334 = ~n2331 & ~n2333 ;
  assign n2335 = ~\pi0075  & n2334 ;
  assign n2336 = ~\pi0092  & n2335 ;
  assign n2337 = ~n2330 & n2336 ;
  assign n2338 = ~n2324 & ~n2337 ;
  assign n2339 = ~n2323 & ~n2338 ;
  assign n2340 = ~n2307 & n2339 ;
  assign n2341 = ~\pi0039  & ~\pi0087  ;
  assign n2342 = n2327 & n2341 ;
  assign n2343 = ~n2262 & n2342 ;
  assign n2344 = n2272 & n2342 ;
  assign n2345 = ~n2271 & n2344 ;
  assign n2346 = ~n2343 & ~n2345 ;
  assign n2347 = \pi0075  & n2342 ;
  assign n2348 = \pi0075  & ~n2219 ;
  assign n2349 = ~n2213 & n2348 ;
  assign n2350 = ~n2347 & ~n2349 ;
  assign n2351 = n2346 & ~n2350 ;
  assign n2352 = ~\pi0216  & ~\pi0221  ;
  assign n2353 = ~n1213 & n2352 ;
  assign n2354 = ~n2226 & n2353 ;
  assign n2355 = ~n2236 & n2354 ;
  assign n2356 = n2294 & ~n2355 ;
  assign n2357 = \pi0299  & ~n2350 ;
  assign n2358 = ~n2296 & n2357 ;
  assign n2359 = ~n2356 & n2358 ;
  assign n2360 = ~n2351 & ~n2359 ;
  assign n2361 = ~\pi0092  & ~n2360 ;
  assign n2362 = ~\pi0087  & ~\pi0100  ;
  assign n2363 = ~\pi0038  & n2362 ;
  assign n2364 = ~\pi0075  & ~\pi0092  ;
  assign n2365 = ~\pi0039  & n2364 ;
  assign n2366 = n2363 & n2365 ;
  assign n2367 = n2342 & n2364 ;
  assign n2368 = ~n2219 & ~n2367 ;
  assign n2369 = ~n2213 & n2368 ;
  assign n2370 = ~n2366 & ~n2369 ;
  assign n2371 = ~n2312 & ~n2369 ;
  assign n2372 = n2318 & n2371 ;
  assign n2373 = ~n2370 & ~n2372 ;
  assign n2374 = ~\pi0054  & ~n2373 ;
  assign n2375 = ~\pi0054  & \pi0074  ;
  assign n2376 = \pi0074  & ~n2219 ;
  assign n2377 = ~n2213 & n2376 ;
  assign n2378 = ~n2375 & ~n2377 ;
  assign n2379 = ~n2374 & ~n2378 ;
  assign n2380 = ~n1286 & n2219 ;
  assign n2381 = ~n1286 & n2210 ;
  assign n2382 = ~n1227 & n2381 ;
  assign n2383 = ~n2380 & ~n2382 ;
  assign n2384 = \pi0092  & n2383 ;
  assign n2385 = n2334 & n2384 ;
  assign n2386 = ~n2330 & n2385 ;
  assign n2387 = \pi0092  & ~n1286 ;
  assign n2388 = ~n2219 & n2387 ;
  assign n2389 = ~n2213 & n2388 ;
  assign n2390 = ~\pi0054  & ~n2389 ;
  assign n2391 = ~n2386 & n2390 ;
  assign n2392 = ~n2379 & n2391 ;
  assign n2393 = ~n2361 & n2392 ;
  assign n2394 = ~n2340 & n2393 ;
  assign n2395 = \pi0054  & ~n2369 ;
  assign n2396 = ~n2366 & n2395 ;
  assign n2397 = ~n2312 & n2395 ;
  assign n2398 = n2318 & n2397 ;
  assign n2399 = ~n2396 & ~n2398 ;
  assign n2400 = ~\pi0074  & n2399 ;
  assign n2401 = ~n2379 & ~n2400 ;
  assign n2402 = ~\pi0100  & n1288 ;
  assign n2403 = n1287 & n2402 ;
  assign n2404 = ~\pi0055  & ~\pi0074  ;
  assign n2405 = \pi0056  & n2404 ;
  assign n2406 = n2403 & n2405 ;
  assign n2407 = n2403 & n2404 ;
  assign n2408 = \pi0056  & ~n1206 ;
  assign n2409 = ~n2407 & n2408 ;
  assign n2410 = ~n1227 & n2409 ;
  assign n2411 = ~\pi0062  & ~n2410 ;
  assign n2412 = ~n2406 & n2411 ;
  assign n2413 = ~n2296 & n2411 ;
  assign n2414 = ~n2295 & n2413 ;
  assign n2415 = ~n2412 & ~n2414 ;
  assign n2416 = ~\pi0055  & ~n2415 ;
  assign n2417 = ~n2401 & n2416 ;
  assign n2418 = ~n2394 & n2417 ;
  assign n2419 = ~n2406 & ~n2410 ;
  assign n2420 = ~n2296 & ~n2410 ;
  assign n2421 = ~n2295 & n2420 ;
  assign n2422 = ~n2419 & ~n2421 ;
  assign n2423 = ~\pi0055  & ~\pi0056  ;
  assign n2424 = ~n1206 & ~n1291 ;
  assign n2425 = ~\pi0056  & n2424 ;
  assign n2426 = ~n1227 & n2425 ;
  assign n2427 = ~n2423 & ~n2426 ;
  assign n2428 = \pi0105  & ~n1230 ;
  assign n2429 = \pi0105  & n1281 ;
  assign n2430 = n1260 & n2429 ;
  assign n2431 = ~n2428 & ~n2430 ;
  assign n2432 = ~n1217 & n2284 ;
  assign n2433 = n2431 & n2432 ;
  assign n2434 = ~\pi0216  & n1281 ;
  assign n2435 = n1260 & n2434 ;
  assign n2436 = ~\pi0228  & n1212 ;
  assign n2437 = ~\pi0216  & ~n2436 ;
  assign n2438 = ~n1217 & ~n2437 ;
  assign n2439 = ~n2435 & n2438 ;
  assign n2440 = n1295 & ~n2439 ;
  assign n2441 = ~n2433 & n2440 ;
  assign n2442 = ~\pi0215  & \pi0221  ;
  assign n2443 = n1224 & n2442 ;
  assign n2444 = ~\pi0056  & ~n1206 ;
  assign n2445 = n1291 & n2444 ;
  assign n2446 = ~n2443 & n2445 ;
  assign n2447 = ~n2441 & n2446 ;
  assign n2448 = n2427 & ~n2447 ;
  assign n2449 = ~\pi0062  & n2448 ;
  assign n2450 = ~n2422 & n2449 ;
  assign n2451 = ~n2407 & n2444 ;
  assign n2452 = ~n1227 & n2451 ;
  assign n2453 = ~\pi0056  & n2404 ;
  assign n2454 = n2403 & n2453 ;
  assign n2455 = ~n2452 & ~n2454 ;
  assign n2456 = ~n2296 & ~n2452 ;
  assign n2457 = ~n2295 & n2456 ;
  assign n2458 = ~n2455 & ~n2457 ;
  assign n2459 = ~n1227 & n2408 ;
  assign n2460 = \pi0062  & ~n2459 ;
  assign n2461 = ~n2458 & n2460 ;
  assign n2462 = ~\pi0059  & n1302 ;
  assign n2463 = ~n2461 & n2462 ;
  assign n2464 = ~n2450 & n2463 ;
  assign n2465 = ~n2418 & n2464 ;
  assign n2466 = ~n1311 & ~n2465 ;
  assign n2467 = ~\pi0057  & ~\pi0059  ;
  assign n2468 = ~\pi0055  & \pi0056  ;
  assign n2469 = \pi0215  & \pi1146  ;
  assign n2470 = ~\pi0154  & n2469 ;
  assign n2471 = \pi0221  & \pi1146  ;
  assign n2472 = ~n1220 & n2471 ;
  assign n2473 = \pi0221  & \pi0939  ;
  assign n2474 = n1220 & n2473 ;
  assign n2475 = ~n2472 & ~n2474 ;
  assign n2476 = \pi0276  & n2291 ;
  assign n2477 = ~n1209 & n2352 ;
  assign n2478 = ~n2476 & ~n2477 ;
  assign n2479 = n2475 & n2478 ;
  assign n2480 = ~\pi0154  & ~\pi0215  ;
  assign n2481 = ~n2479 & n2480 ;
  assign n2482 = ~n2470 & ~n2481 ;
  assign n2483 = ~n2469 & ~n2476 ;
  assign n2484 = n2475 & n2483 ;
  assign n2485 = \pi0215  & ~\pi1146  ;
  assign n2486 = \pi0154  & ~n2485 ;
  assign n2487 = ~n2484 & n2486 ;
  assign n2488 = \pi0056  & ~n2487 ;
  assign n2489 = n2482 & n2488 ;
  assign n2490 = ~n2468 & ~n2489 ;
  assign n2491 = ~\pi0062  & n2490 ;
  assign n2492 = ~\pi0216  & ~\pi0228  ;
  assign n2493 = ~n2469 & n2492 ;
  assign n2494 = n2475 & n2493 ;
  assign n2495 = n1259 & n2494 ;
  assign n2496 = n1249 & n2495 ;
  assign n2497 = n1281 & n2496 ;
  assign n2498 = n1291 & ~n2487 ;
  assign n2499 = n2497 & n2498 ;
  assign n2500 = n2482 & ~n2487 ;
  assign n2501 = ~\pi0062  & ~n2500 ;
  assign n2502 = ~n2499 & n2501 ;
  assign n2503 = ~n2491 & ~n2502 ;
  assign n2504 = n1291 & n2423 ;
  assign n2505 = n1281 & ~n2487 ;
  assign n2506 = n2496 & n2505 ;
  assign n2507 = n2504 & n2506 ;
  assign n2508 = \pi0062  & ~n2500 ;
  assign n2509 = ~n2507 & n2508 ;
  assign n2510 = n2503 & ~n2509 ;
  assign n2511 = ~\pi0054  & ~\pi0074  ;
  assign n2512 = \pi0299  & n2469 ;
  assign n2513 = n2256 & ~n2479 ;
  assign n2514 = ~n2512 & ~n2513 ;
  assign n2515 = ~\pi0154  & ~n2514 ;
  assign n2516 = ~n2497 & n2515 ;
  assign n2517 = \pi0222  & \pi1146  ;
  assign n2518 = ~n2192 & n2517 ;
  assign n2519 = \pi0222  & \pi0939  ;
  assign n2520 = n2192 & n2519 ;
  assign n2521 = ~n2518 & ~n2520 ;
  assign n2522 = ~\pi0222  & \pi0224  ;
  assign n2523 = \pi0276  & n2522 ;
  assign n2524 = ~\pi0223  & ~n2523 ;
  assign n2525 = n2521 & n2524 ;
  assign n2526 = \pi0223  & ~\pi1146  ;
  assign n2527 = ~\pi0299  & ~n2526 ;
  assign n2528 = ~\pi0154  & n2527 ;
  assign n2529 = ~n2525 & n2528 ;
  assign n2530 = \pi0154  & n2527 ;
  assign n2531 = ~n2525 & n2530 ;
  assign n2532 = \pi0154  & \pi0299  ;
  assign n2533 = ~n2485 & n2532 ;
  assign n2534 = ~n2484 & n2533 ;
  assign n2535 = ~n2531 & ~n2534 ;
  assign n2536 = n1286 & n2402 ;
  assign n2537 = n2535 & n2536 ;
  assign n2538 = ~n2529 & n2537 ;
  assign n2539 = ~n2516 & n2538 ;
  assign n2540 = ~n2525 & n2527 ;
  assign n2541 = ~\pi0299  & ~n2540 ;
  assign n2542 = ~n2487 & ~n2540 ;
  assign n2543 = n2482 & n2542 ;
  assign n2544 = ~n2541 & ~n2543 ;
  assign n2545 = ~n2536 & ~n2544 ;
  assign n2546 = \pi0092  & ~n2545 ;
  assign n2547 = ~n2539 & n2546 ;
  assign n2548 = n2511 & ~n2547 ;
  assign n2549 = ~n2511 & ~n2544 ;
  assign n2550 = ~\pi0055  & ~n2549 ;
  assign n2551 = ~n2548 & n2550 ;
  assign n2552 = \pi0087  & ~n2328 ;
  assign n2553 = ~n2544 & n2552 ;
  assign n2554 = \pi0087  & n2402 ;
  assign n2555 = n2535 & n2554 ;
  assign n2556 = ~n2529 & n2555 ;
  assign n2557 = ~n2516 & n2556 ;
  assign n2558 = ~n2553 & ~n2557 ;
  assign n2559 = ~\pi0075  & ~n2558 ;
  assign n2560 = ~\pi0038  & n2535 ;
  assign n2561 = \pi0038  & ~n2540 ;
  assign n2562 = ~\pi0100  & ~n2561 ;
  assign n2563 = ~\pi0100  & \pi0299  ;
  assign n2564 = ~n2500 & n2563 ;
  assign n2565 = ~n2562 & ~n2564 ;
  assign n2566 = ~n2560 & ~n2565 ;
  assign n2567 = ~n1360 & ~n1864 ;
  assign n2568 = ~\pi0051  & ~n2567 ;
  assign n2569 = ~n1629 & ~n1868 ;
  assign n2570 = ~n2568 & n2569 ;
  assign n2571 = ~n1364 & n2570 ;
  assign n2572 = ~n2048 & n2570 ;
  assign n2573 = ~n2045 & n2572 ;
  assign n2574 = ~n2571 & ~n2573 ;
  assign n2575 = ~\pi0095  & n1634 ;
  assign n2576 = ~\pi0072  & n2575 ;
  assign n2577 = ~n1962 & n2576 ;
  assign n2578 = \pi0072  & n2575 ;
  assign n2579 = ~n1628 & n2578 ;
  assign n2580 = ~n2577 & ~n2579 ;
  assign n2581 = n2574 & ~n2580 ;
  assign n2582 = ~\pi0035  & n1618 ;
  assign n2583 = n1354 & n2582 ;
  assign n2584 = n1358 & n2583 ;
  assign n2585 = \pi0040  & ~n2584 ;
  assign n2586 = n1324 & n1329 ;
  assign n2587 = n1328 & n2586 ;
  assign n2588 = n1319 & n2587 ;
  assign n2589 = \pi0032  & ~n2588 ;
  assign n2590 = ~n2585 & ~n2589 ;
  assign n2591 = ~\pi0095  & ~n2590 ;
  assign n2592 = ~\pi0039  & ~n1639 ;
  assign n2593 = ~n2591 & n2592 ;
  assign n2594 = ~n2581 & n2593 ;
  assign n2595 = \pi0039  & n1281 ;
  assign n2596 = n1260 & n2595 ;
  assign n2597 = ~n2514 & ~n2596 ;
  assign n2598 = ~n2594 & n2597 ;
  assign n2599 = ~n2494 & ~n2514 ;
  assign n2600 = ~n2540 & ~n2599 ;
  assign n2601 = ~n2598 & n2600 ;
  assign n2602 = ~\pi0154  & ~n2565 ;
  assign n2603 = ~n2601 & n2602 ;
  assign n2604 = ~n2566 & ~n2603 ;
  assign n2605 = ~\pi0161  & ~\pi0166  ;
  assign n2606 = ~n2238 & ~n2605 ;
  assign n2607 = n1259 & n2606 ;
  assign n2608 = n1249 & n2607 ;
  assign n2609 = n1281 & n2608 ;
  assign n2610 = ~\pi0252  & n2605 ;
  assign n2611 = n1259 & n2610 ;
  assign n2612 = n1281 & n2611 ;
  assign n2613 = n1249 & n2612 ;
  assign n2614 = ~\pi0152  & ~n2613 ;
  assign n2615 = ~n2609 & n2614 ;
  assign n2616 = n1281 & ~n2238 ;
  assign n2617 = n1260 & n2616 ;
  assign n2618 = \pi0152  & ~n2617 ;
  assign n2619 = ~\pi0154  & \pi0299  ;
  assign n2620 = n1288 & n2619 ;
  assign n2621 = n2493 & n2620 ;
  assign n2622 = n2475 & n2621 ;
  assign n2623 = ~n2618 & n2622 ;
  assign n2624 = ~n2615 & n2623 ;
  assign n2625 = \pi0100  & n2544 ;
  assign n2626 = ~n2624 & n2625 ;
  assign n2627 = ~\pi0087  & ~n2626 ;
  assign n2628 = ~\pi0075  & n2627 ;
  assign n2629 = n2604 & n2628 ;
  assign n2630 = ~n2559 & ~n2629 ;
  assign n2631 = \pi0075  & ~n2540 ;
  assign n2632 = ~\pi0092  & ~n2631 ;
  assign n2633 = ~\pi0092  & \pi0299  ;
  assign n2634 = ~n2500 & n2633 ;
  assign n2635 = ~n2632 & ~n2634 ;
  assign n2636 = n2550 & ~n2635 ;
  assign n2637 = n2630 & n2636 ;
  assign n2638 = ~n2551 & ~n2637 ;
  assign n2639 = \pi0055  & ~n2500 ;
  assign n2640 = ~n2499 & n2639 ;
  assign n2641 = ~\pi0056  & ~n2640 ;
  assign n2642 = ~n2509 & n2641 ;
  assign n2643 = n2638 & n2642 ;
  assign n2644 = ~n2510 & ~n2643 ;
  assign n2645 = n2467 & ~n2644 ;
  assign n2646 = ~n2467 & ~n2487 ;
  assign n2647 = n2482 & n2646 ;
  assign n2648 = ~\pi0239  & ~n2647 ;
  assign n2649 = ~n2645 & n2648 ;
  assign n2650 = ~\pi0215  & n2352 ;
  assign n2651 = n1209 & n1633 ;
  assign n2652 = n2650 & n2651 ;
  assign n2653 = \pi0154  & n2652 ;
  assign n2654 = ~n2487 & ~n2653 ;
  assign n2655 = n2406 & n2654 ;
  assign n2656 = n2497 & n2655 ;
  assign n2657 = n2475 & ~n2476 ;
  assign n2658 = ~\pi0215  & ~n2657 ;
  assign n2659 = ~n2652 & ~n2658 ;
  assign n2660 = n2654 & n2659 ;
  assign n2661 = \pi0056  & n2482 ;
  assign n2662 = n2660 & n2661 ;
  assign n2663 = ~\pi0062  & ~n2662 ;
  assign n2664 = ~n2656 & n2663 ;
  assign n2665 = ~\pi0299  & n1633 ;
  assign n2666 = n2214 & n2665 ;
  assign n2667 = ~n2540 & ~n2666 ;
  assign n2668 = ~\pi0299  & n2667 ;
  assign n2669 = n2482 & n2667 ;
  assign n2670 = n2660 & n2669 ;
  assign n2671 = ~n2668 & ~n2670 ;
  assign n2672 = \pi0092  & n2671 ;
  assign n2673 = n2497 & n2654 ;
  assign n2674 = n2482 & n2660 ;
  assign n2675 = ~n2673 & ~n2674 ;
  assign n2676 = \pi0299  & n1286 ;
  assign n2677 = n2328 & n2676 ;
  assign n2678 = ~n2675 & n2677 ;
  assign n2679 = n2672 & ~n2678 ;
  assign n2680 = ~\pi0224  & ~n1633 ;
  assign n2681 = \pi0224  & ~\pi0276  ;
  assign n2682 = ~\pi0222  & ~n2681 ;
  assign n2683 = ~n2680 & n2682 ;
  assign n2684 = ~\pi0032  & n1732 ;
  assign n2685 = n1721 & n2684 ;
  assign n2686 = n1319 & n2685 ;
  assign n2687 = ~\pi0095  & n2682 ;
  assign n2688 = n2686 & n2687 ;
  assign n2689 = ~n2683 & ~n2688 ;
  assign n2690 = n2527 & ~n2689 ;
  assign n2691 = ~\pi0039  & ~n2527 ;
  assign n2692 = ~\pi0039  & ~\pi0223  ;
  assign n2693 = n2521 & n2692 ;
  assign n2694 = ~n2691 & ~n2693 ;
  assign n2695 = ~n2690 & ~n2694 ;
  assign n2696 = \pi0039  & ~n2671 ;
  assign n2697 = n2297 & ~n2675 ;
  assign n2698 = ~n2696 & ~n2697 ;
  assign n2699 = ~n2695 & n2698 ;
  assign n2700 = \pi0072  & n1324 ;
  assign n2701 = n1328 & n2700 ;
  assign n2702 = n1319 & n2701 ;
  assign n2703 = n2575 & ~n2702 ;
  assign n2704 = n2574 & n2703 ;
  assign n2705 = ~\pi0228  & ~n1633 ;
  assign n2706 = ~n1639 & n2705 ;
  assign n2707 = ~n2591 & n2706 ;
  assign n2708 = ~n2704 & n2707 ;
  assign n2709 = \pi0228  & ~n1633 ;
  assign n2710 = ~n2225 & ~n2709 ;
  assign n2711 = ~\pi0095  & ~n2225 ;
  assign n2712 = n2686 & n2711 ;
  assign n2713 = ~n2710 & ~n2712 ;
  assign n2714 = \pi0154  & n2713 ;
  assign n2715 = n2650 & ~n2714 ;
  assign n2716 = ~\pi0095  & n2686 ;
  assign n2717 = n1633 & n1638 ;
  assign n2718 = ~n2716 & ~n2717 ;
  assign n2719 = \pi0154  & ~\pi0228  ;
  assign n2720 = n2718 & n2719 ;
  assign n2721 = n1209 & ~n1633 ;
  assign n2722 = ~n2716 & n2721 ;
  assign n2723 = ~n2720 & ~n2722 ;
  assign n2724 = n2715 & n2723 ;
  assign n2725 = ~n2708 & n2724 ;
  assign n2726 = ~n2484 & ~n2485 ;
  assign n2727 = \pi0154  & n2650 ;
  assign n2728 = ~n2713 & n2727 ;
  assign n2729 = ~n2720 & n2728 ;
  assign n2730 = ~n2726 & ~n2729 ;
  assign n2731 = ~n2725 & n2730 ;
  assign n2732 = \pi0299  & n2698 ;
  assign n2733 = ~n2731 & n2732 ;
  assign n2734 = ~n2699 & ~n2733 ;
  assign n2735 = ~\pi0087  & n2327 ;
  assign n2736 = ~n2734 & n2735 ;
  assign n2737 = \pi0087  & n2671 ;
  assign n2738 = ~\pi0039  & \pi0299  ;
  assign n2739 = n2327 & n2738 ;
  assign n2740 = ~n2675 & n2739 ;
  assign n2741 = n2737 & ~n2740 ;
  assign n2742 = ~\pi0075  & ~n2741 ;
  assign n2743 = \pi0100  & n2622 ;
  assign n2744 = ~n2618 & n2743 ;
  assign n2745 = ~n2615 & n2744 ;
  assign n2746 = ~\pi0087  & ~n2327 ;
  assign n2747 = n2671 & n2746 ;
  assign n2748 = ~n2745 & n2747 ;
  assign n2749 = n2511 & ~n2748 ;
  assign n2750 = n2742 & n2749 ;
  assign n2751 = ~n2736 & n2750 ;
  assign n2752 = ~n2679 & n2751 ;
  assign n2753 = \pi0075  & ~n2666 ;
  assign n2754 = ~n2540 & n2753 ;
  assign n2755 = ~\pi0299  & n2754 ;
  assign n2756 = n2482 & n2754 ;
  assign n2757 = n2660 & n2756 ;
  assign n2758 = ~n2755 & ~n2757 ;
  assign n2759 = ~\pi0092  & n2758 ;
  assign n2760 = n2511 & ~n2759 ;
  assign n2761 = ~n2679 & n2760 ;
  assign n2762 = ~n2511 & ~n2671 ;
  assign n2763 = ~\pi0055  & ~n2762 ;
  assign n2764 = ~n2761 & n2763 ;
  assign n2765 = ~n2752 & n2764 ;
  assign n2766 = n2664 & n2765 ;
  assign n2767 = n1291 & n2654 ;
  assign n2768 = n2497 & n2767 ;
  assign n2769 = \pi0055  & ~n2674 ;
  assign n2770 = ~n2768 & n2769 ;
  assign n2771 = ~\pi0056  & ~n2770 ;
  assign n2772 = n2664 & ~n2771 ;
  assign n2773 = n2504 & n2654 ;
  assign n2774 = n2497 & n2773 ;
  assign n2775 = \pi0062  & ~n2674 ;
  assign n2776 = ~n2774 & n2775 ;
  assign n2777 = n2467 & ~n2776 ;
  assign n2778 = ~n2772 & n2777 ;
  assign n2779 = ~n2766 & n2778 ;
  assign n2780 = ~n2467 & n2482 ;
  assign n2781 = n2660 & n2780 ;
  assign n2782 = \pi0239  & ~n2781 ;
  assign n2783 = ~n2779 & n2782 ;
  assign n2784 = ~n2649 & ~n2783 ;
  assign n2785 = \pi0221  & \pi1145  ;
  assign n2786 = ~n1220 & n2785 ;
  assign n2787 = \pi0221  & \pi0927  ;
  assign n2788 = n1220 & n2787 ;
  assign n2789 = ~n2786 & ~n2788 ;
  assign n2790 = ~\pi0215  & ~n2789 ;
  assign n2791 = \pi0216  & \pi0274  ;
  assign n2792 = ~\pi0221  & ~n2791 ;
  assign n2793 = ~\pi0215  & \pi0216  ;
  assign n2794 = ~\pi0151  & ~\pi0215  ;
  assign n2795 = ~n1209 & n2794 ;
  assign n2796 = ~n2793 & ~n2795 ;
  assign n2797 = n2792 & ~n2796 ;
  assign n2798 = ~n2790 & ~n2797 ;
  assign n2799 = n1295 & ~n2791 ;
  assign n2800 = n2651 & n2799 ;
  assign n2801 = \pi0235  & n2800 ;
  assign n2802 = \pi0215  & \pi1145  ;
  assign n2803 = ~n2467 & ~n2802 ;
  assign n2804 = ~n2801 & n2803 ;
  assign n2805 = n2798 & n2804 ;
  assign n2806 = ~\pi0235  & n2467 ;
  assign n2807 = ~\pi0062  & n2806 ;
  assign n2808 = ~n2802 & n2806 ;
  assign n2809 = n2798 & n2808 ;
  assign n2810 = ~n2807 & ~n2809 ;
  assign n2811 = n2492 & ~n2802 ;
  assign n2812 = n2789 & n2811 ;
  assign n2813 = n1291 & n2812 ;
  assign n2814 = n1281 & n2813 ;
  assign n2815 = n1260 & n2814 ;
  assign n2816 = n2423 & n2806 ;
  assign n2817 = n2815 & n2816 ;
  assign n2818 = n2810 & ~n2817 ;
  assign n2819 = ~n2805 & n2818 ;
  assign n2820 = n2798 & ~n2802 ;
  assign n2821 = \pi0055  & ~n2820 ;
  assign n2822 = ~n2815 & n2821 ;
  assign n2823 = ~\pi0056  & ~n2822 ;
  assign n2824 = \pi0223  & ~\pi1145  ;
  assign n2825 = \pi0222  & \pi1145  ;
  assign n2826 = ~n2192 & n2825 ;
  assign n2827 = \pi0222  & \pi0927  ;
  assign n2828 = n2192 & n2827 ;
  assign n2829 = ~n2826 & ~n2828 ;
  assign n2830 = \pi0223  & \pi1145  ;
  assign n2831 = \pi0224  & \pi0274  ;
  assign n2832 = n2522 & ~n2831 ;
  assign n2833 = ~n2830 & ~n2832 ;
  assign n2834 = n2829 & n2833 ;
  assign n2835 = ~n2824 & ~n2834 ;
  assign n2836 = ~\pi0299  & ~n2835 ;
  assign n2837 = \pi0299  & ~n2802 ;
  assign n2838 = n2798 & n2837 ;
  assign n2839 = ~n2836 & ~n2838 ;
  assign n2840 = ~n2511 & ~n2839 ;
  assign n2841 = ~\pi0055  & ~n2840 ;
  assign n2842 = n2823 & ~n2841 ;
  assign n2843 = \pi0075  & ~n2839 ;
  assign n2844 = ~\pi0092  & ~n2843 ;
  assign n2845 = \pi0075  & n2844 ;
  assign n2846 = \pi0299  & ~n2820 ;
  assign n2847 = ~\pi0299  & ~n2824 ;
  assign n2848 = ~n2834 & n2847 ;
  assign n2849 = ~\pi0087  & ~n2848 ;
  assign n2850 = ~n2846 & n2849 ;
  assign n2851 = ~\pi0039  & \pi0100  ;
  assign n2852 = ~n2618 & n2851 ;
  assign n2853 = ~n2615 & n2852 ;
  assign n2854 = \pi0100  & ~n2853 ;
  assign n2855 = ~\pi0038  & ~\pi0087  ;
  assign n2856 = n2812 & n2855 ;
  assign n2857 = ~n2848 & n2856 ;
  assign n2858 = ~n2854 & n2857 ;
  assign n2859 = ~n2850 & ~n2858 ;
  assign n2860 = ~n2596 & ~n2853 ;
  assign n2861 = ~n2850 & n2860 ;
  assign n2862 = ~n2594 & n2861 ;
  assign n2863 = ~n2859 & ~n2862 ;
  assign n2864 = n2552 & ~n2839 ;
  assign n2865 = n1281 & n2812 ;
  assign n2866 = n1260 & n2865 ;
  assign n2867 = n2846 & ~n2866 ;
  assign n2868 = n2554 & ~n2848 ;
  assign n2869 = ~n2867 & n2868 ;
  assign n2870 = ~n2864 & ~n2869 ;
  assign n2871 = n2844 & n2870 ;
  assign n2872 = ~n2863 & n2871 ;
  assign n2873 = ~n2845 & ~n2872 ;
  assign n2874 = n2402 & ~n2848 ;
  assign n2875 = n1286 & n2874 ;
  assign n2876 = ~n2867 & n2875 ;
  assign n2877 = ~n2536 & ~n2839 ;
  assign n2878 = \pi0092  & ~n2877 ;
  assign n2879 = ~n2876 & n2878 ;
  assign n2880 = n2511 & ~n2879 ;
  assign n2881 = n2823 & n2880 ;
  assign n2882 = n2873 & n2881 ;
  assign n2883 = ~n2842 & ~n2882 ;
  assign n2884 = n2407 & n2812 ;
  assign n2885 = n1281 & n2884 ;
  assign n2886 = n1260 & n2885 ;
  assign n2887 = ~\pi0062  & ~n2820 ;
  assign n2888 = ~n2886 & n2887 ;
  assign n2889 = ~n1292 & ~n2888 ;
  assign n2890 = ~n2805 & ~n2889 ;
  assign n2891 = n2883 & n2890 ;
  assign n2892 = ~n2819 & ~n2891 ;
  assign n2893 = ~n2800 & ~n2802 ;
  assign n2894 = ~n2504 & n2893 ;
  assign n2895 = n2798 & n2894 ;
  assign n2896 = ~n2504 & ~n2895 ;
  assign n2897 = ~\pi0151  & ~\pi0228  ;
  assign n2898 = n1281 & n2897 ;
  assign n2899 = n1260 & n2898 ;
  assign n2900 = ~\pi0151  & ~n1209 ;
  assign n2901 = ~n2651 & ~n2900 ;
  assign n2902 = n2792 & ~n2901 ;
  assign n2903 = ~n2899 & n2902 ;
  assign n2904 = ~\pi0274  & n2291 ;
  assign n2905 = n2789 & ~n2802 ;
  assign n2906 = ~n2904 & n2905 ;
  assign n2907 = ~n2903 & n2906 ;
  assign n2908 = \pi0215  & ~\pi1145  ;
  assign n2909 = ~n2895 & ~n2908 ;
  assign n2910 = ~n2907 & n2909 ;
  assign n2911 = ~n2896 & ~n2910 ;
  assign n2912 = \pi0062  & ~n2911 ;
  assign n2913 = \pi0235  & n2467 ;
  assign n2914 = ~n2912 & n2913 ;
  assign n2915 = ~\pi0228  & n2718 ;
  assign n2916 = \pi0151  & ~n2713 ;
  assign n2917 = ~n2915 & n2916 ;
  assign n2918 = ~\pi0216  & n2789 ;
  assign n2919 = ~n2917 & n2918 ;
  assign n2920 = n2199 & ~n2831 ;
  assign n2921 = ~n2680 & n2920 ;
  assign n2922 = ~\pi0095  & n2920 ;
  assign n2923 = n2686 & n2922 ;
  assign n2924 = ~n2921 & ~n2923 ;
  assign n2925 = ~\pi0223  & ~n2829 ;
  assign n2926 = ~\pi0299  & ~n2830 ;
  assign n2927 = ~n2925 & n2926 ;
  assign n2928 = n2924 & n2927 ;
  assign n2929 = n2789 & ~n2792 ;
  assign n2930 = n2206 & ~n2929 ;
  assign n2931 = ~n2928 & n2930 ;
  assign n2932 = ~n2919 & n2931 ;
  assign n2933 = ~\pi0151  & ~n2721 ;
  assign n2934 = ~\pi0095  & ~\pi0151  ;
  assign n2935 = n2686 & n2934 ;
  assign n2936 = ~n2933 & ~n2935 ;
  assign n2937 = n2931 & ~n2936 ;
  assign n2938 = ~n2708 & n2937 ;
  assign n2939 = ~n2932 & ~n2938 ;
  assign n2940 = ~\pi0039  & ~n2837 ;
  assign n2941 = ~n2928 & n2940 ;
  assign n2942 = ~\pi0228  & ~n2618 ;
  assign n2943 = ~n2615 & n2942 ;
  assign n2944 = n2933 & ~n2943 ;
  assign n2945 = ~n2899 & ~n2901 ;
  assign n2946 = ~\pi0216  & ~n2945 ;
  assign n2947 = n2789 & n2946 ;
  assign n2948 = ~n2944 & n2947 ;
  assign n2949 = n2256 & ~n2929 ;
  assign n2950 = ~n2948 & n2949 ;
  assign n2951 = \pi0299  & n2802 ;
  assign n2952 = n1288 & ~n2666 ;
  assign n2953 = ~n2848 & n2952 ;
  assign n2954 = ~n2951 & n2953 ;
  assign n2955 = ~n2950 & n2954 ;
  assign n2956 = ~n1288 & ~n2666 ;
  assign n2957 = ~n2848 & n2956 ;
  assign n2958 = \pi0100  & ~n2957 ;
  assign n2959 = n2798 & n2893 ;
  assign n2960 = \pi0100  & \pi0299  ;
  assign n2961 = ~n2959 & n2960 ;
  assign n2962 = ~n2958 & ~n2961 ;
  assign n2963 = ~n2955 & ~n2962 ;
  assign n2964 = n2297 & ~n2908 ;
  assign n2965 = ~n2907 & n2964 ;
  assign n2966 = ~\pi0038  & ~n2666 ;
  assign n2967 = ~n2848 & n2966 ;
  assign n2968 = ~n1288 & ~n2967 ;
  assign n2969 = ~n2965 & ~n2968 ;
  assign n2970 = ~n2963 & n2969 ;
  assign n2971 = ~n2941 & n2970 ;
  assign n2972 = n2939 & n2971 ;
  assign n2973 = \pi0038  & ~n2666 ;
  assign n2974 = ~n2848 & n2973 ;
  assign n2975 = ~\pi0100  & ~n2974 ;
  assign n2976 = n2563 & ~n2959 ;
  assign n2977 = ~n2975 & ~n2976 ;
  assign n2978 = ~n2963 & n2977 ;
  assign n2979 = n2753 & ~n2848 ;
  assign n2980 = ~\pi0092  & ~n2979 ;
  assign n2981 = n2633 & ~n2959 ;
  assign n2982 = ~n2980 & ~n2981 ;
  assign n2983 = ~\pi0087  & ~n2982 ;
  assign n2984 = ~n2978 & n2983 ;
  assign n2985 = ~n2972 & n2984 ;
  assign n2986 = \pi0299  & ~n2908 ;
  assign n2987 = ~n2907 & n2986 ;
  assign n2988 = ~n2666 & ~n2848 ;
  assign n2989 = n2328 & n2988 ;
  assign n2990 = ~n2987 & n2989 ;
  assign n2991 = ~\pi0299  & ~n2328 ;
  assign n2992 = ~n2328 & n2893 ;
  assign n2993 = n2798 & n2992 ;
  assign n2994 = ~n2991 & ~n2993 ;
  assign n2995 = n2988 & ~n2994 ;
  assign n2996 = \pi0087  & ~n2995 ;
  assign n2997 = ~n2990 & n2996 ;
  assign n2998 = ~\pi0075  & ~n2997 ;
  assign n2999 = ~n2982 & ~n2998 ;
  assign n3000 = ~n1286 & ~n2666 ;
  assign n3001 = ~n2848 & n3000 ;
  assign n3002 = \pi0092  & ~n3001 ;
  assign n3003 = \pi0092  & \pi0299  ;
  assign n3004 = ~n2959 & n3003 ;
  assign n3005 = ~n3002 & ~n3004 ;
  assign n3006 = ~n2995 & ~n3005 ;
  assign n3007 = ~n2990 & n3006 ;
  assign n3008 = ~\pi0056  & n1291 ;
  assign n3009 = ~n1291 & n2893 ;
  assign n3010 = n2798 & n3009 ;
  assign n3011 = \pi0055  & ~n3010 ;
  assign n3012 = ~\pi0056  & ~n3011 ;
  assign n3013 = ~n3008 & ~n3012 ;
  assign n3014 = ~n2908 & ~n3012 ;
  assign n3015 = ~n2907 & n3014 ;
  assign n3016 = ~n3013 & ~n3015 ;
  assign n3017 = ~n1286 & ~n3005 ;
  assign n3018 = n2511 & ~n3017 ;
  assign n3019 = n3016 & n3018 ;
  assign n3020 = ~n3007 & n3019 ;
  assign n3021 = ~n2999 & n3020 ;
  assign n3022 = ~n2985 & n3021 ;
  assign n3023 = ~n2511 & ~n2666 ;
  assign n3024 = ~n2848 & n3023 ;
  assign n3025 = ~\pi0055  & ~n3024 ;
  assign n3026 = ~\pi0055  & \pi0299  ;
  assign n3027 = ~n2959 & n3026 ;
  assign n3028 = ~n3025 & ~n3027 ;
  assign n3029 = n3016 & n3028 ;
  assign n3030 = ~\pi0055  & n1291 ;
  assign n3031 = ~n2407 & n2893 ;
  assign n3032 = n2798 & n3031 ;
  assign n3033 = ~\pi0062  & ~n3032 ;
  assign n3034 = ~n3030 & n3033 ;
  assign n3035 = ~n2908 & n3033 ;
  assign n3036 = ~n2907 & n3035 ;
  assign n3037 = ~n3034 & ~n3036 ;
  assign n3038 = ~n1292 & n3037 ;
  assign n3039 = ~n3029 & ~n3038 ;
  assign n3040 = ~n3022 & n3039 ;
  assign n3041 = n2914 & ~n3040 ;
  assign n3042 = ~n2892 & ~n3041 ;
  assign n3043 = \pi0223  & \pi1143  ;
  assign n3044 = ~\pi0299  & n3043 ;
  assign n3045 = n1633 & n2214 ;
  assign n3046 = n3044 & ~n3045 ;
  assign n3047 = \pi0224  & \pi0264  ;
  assign n3048 = ~\pi0222  & ~n3047 ;
  assign n3049 = ~\pi0224  & \pi0284  ;
  assign n3050 = ~n1633 & n3049 ;
  assign n3051 = n3048 & ~n3050 ;
  assign n3052 = \pi0222  & \pi0944  ;
  assign n3053 = n2192 & n3052 ;
  assign n3054 = \pi0222  & \pi1143  ;
  assign n3055 = ~n2192 & n3054 ;
  assign n3056 = ~n3053 & ~n3055 ;
  assign n3057 = ~n3051 & n3056 ;
  assign n3058 = ~\pi0223  & ~\pi0299  ;
  assign n3059 = ~n3045 & n3058 ;
  assign n3060 = ~n3057 & n3059 ;
  assign n3061 = ~n3046 & ~n3060 ;
  assign n3062 = ~\pi0299  & n3061 ;
  assign n3063 = \pi0221  & \pi1143  ;
  assign n3064 = ~n1220 & n3063 ;
  assign n3065 = \pi0221  & \pi0944  ;
  assign n3066 = n1220 & n3065 ;
  assign n3067 = ~n3064 & ~n3066 ;
  assign n3068 = ~\pi0215  & ~n3067 ;
  assign n3069 = ~\pi0146  & ~\pi0228  ;
  assign n3070 = ~n2651 & ~n3069 ;
  assign n3071 = ~\pi0216  & ~n3070 ;
  assign n3072 = ~\pi0105  & ~\pi0146  ;
  assign n3073 = \pi0105  & \pi0284  ;
  assign n3074 = ~n1633 & n3073 ;
  assign n3075 = ~n3072 & ~n3074 ;
  assign n3076 = n1824 & ~n3075 ;
  assign n3077 = ~n3071 & ~n3076 ;
  assign n3078 = \pi0216  & \pi0264  ;
  assign n3079 = ~\pi0221  & ~n3078 ;
  assign n3080 = ~\pi0215  & n3079 ;
  assign n3081 = n3077 & n3080 ;
  assign n3082 = ~n3068 & ~n3081 ;
  assign n3083 = \pi0215  & \pi1143  ;
  assign n3084 = n3061 & ~n3083 ;
  assign n3085 = n3082 & n3084 ;
  assign n3086 = ~n3062 & ~n3085 ;
  assign n3087 = \pi0092  & n3086 ;
  assign n3088 = \pi0092  & n1286 ;
  assign n3089 = n2328 & n3088 ;
  assign n3090 = ~n3087 & ~n3089 ;
  assign n3091 = n2387 & n3086 ;
  assign n3092 = n2511 & ~n3091 ;
  assign n3093 = n3090 & n3092 ;
  assign n3094 = \pi0215  & ~\pi1143  ;
  assign n3095 = \pi0299  & ~n3094 ;
  assign n3096 = n3067 & ~n3083 ;
  assign n3097 = ~\pi0264  & n2291 ;
  assign n3098 = n3096 & ~n3097 ;
  assign n3099 = \pi0146  & ~n2280 ;
  assign n3100 = ~\pi0284  & n1281 ;
  assign n3101 = n1260 & n3100 ;
  assign n3102 = ~\pi0228  & ~n3101 ;
  assign n3103 = ~n3099 & n3102 ;
  assign n3104 = \pi0228  & ~n3075 ;
  assign n3105 = ~n2651 & n3079 ;
  assign n3106 = ~n3104 & n3105 ;
  assign n3107 = ~n3103 & n3106 ;
  assign n3108 = n3098 & ~n3107 ;
  assign n3109 = n3095 & ~n3108 ;
  assign n3110 = n2328 & n3061 ;
  assign n3111 = n3092 & n3110 ;
  assign n3112 = ~n3109 & n3111 ;
  assign n3113 = ~n3093 & ~n3112 ;
  assign n3114 = ~n2511 & ~n3086 ;
  assign n3115 = n3113 & ~n3114 ;
  assign n3116 = ~\pi0146  & ~n1633 ;
  assign n3117 = ~n1639 & n3116 ;
  assign n3118 = ~n2591 & n3117 ;
  assign n3119 = ~n2704 & n3118 ;
  assign n3120 = \pi0146  & n2718 ;
  assign n3121 = ~\pi0284  & ~n3120 ;
  assign n3122 = ~n3119 & n3121 ;
  assign n3123 = n2492 & n3122 ;
  assign n3124 = ~n1639 & ~n2591 ;
  assign n3125 = ~n2581 & n3124 ;
  assign n3126 = \pi0146  & ~n3125 ;
  assign n3127 = \pi0284  & n2492 ;
  assign n3128 = ~n3126 & n3127 ;
  assign n3129 = ~n3123 & ~n3128 ;
  assign n3130 = n1295 & ~n3078 ;
  assign n3131 = ~n1633 & ~n3104 ;
  assign n3132 = ~\pi0105  & \pi0146  ;
  assign n3133 = \pi0228  & ~n3132 ;
  assign n3134 = ~\pi0216  & n3133 ;
  assign n3135 = ~n3131 & n3134 ;
  assign n3136 = ~\pi0095  & n3134 ;
  assign n3137 = n2686 & n3136 ;
  assign n3138 = ~n3135 & ~n3137 ;
  assign n3139 = n3130 & n3138 ;
  assign n3140 = n3129 & n3139 ;
  assign n3141 = \pi0299  & ~n3083 ;
  assign n3142 = ~n3068 & n3141 ;
  assign n3143 = n2297 & ~n3094 ;
  assign n3144 = ~n3108 & n3143 ;
  assign n3145 = \pi0039  & ~n3061 ;
  assign n3146 = ~\pi0038  & ~n3145 ;
  assign n3147 = ~n3144 & n3146 ;
  assign n3148 = n3142 & n3147 ;
  assign n3149 = ~n3140 & n3148 ;
  assign n3150 = ~\pi0299  & ~n3043 ;
  assign n3151 = ~\pi0284  & ~n1633 ;
  assign n3152 = ~\pi0224  & ~n3151 ;
  assign n3153 = ~\pi0095  & ~\pi0224  ;
  assign n3154 = n2686 & n3153 ;
  assign n3155 = ~n3152 & ~n3154 ;
  assign n3156 = n3048 & n3155 ;
  assign n3157 = n1633 & n3048 ;
  assign n3158 = ~\pi0095  & n3048 ;
  assign n3159 = n2686 & n3158 ;
  assign n3160 = ~n3157 & ~n3159 ;
  assign n3161 = n3056 & n3160 ;
  assign n3162 = ~n3156 & n3161 ;
  assign n3163 = ~\pi0223  & ~n3162 ;
  assign n3164 = n3150 & ~n3163 ;
  assign n3165 = n3056 & n3150 ;
  assign n3166 = ~n3156 & n3165 ;
  assign n3167 = ~\pi0039  & ~n3166 ;
  assign n3168 = ~n3164 & n3167 ;
  assign n3169 = n3147 & ~n3168 ;
  assign n3170 = \pi0038  & n3061 ;
  assign n3171 = ~\pi0100  & ~n3170 ;
  assign n3172 = n3082 & ~n3083 ;
  assign n3173 = n2563 & ~n3172 ;
  assign n3174 = ~n3171 & ~n3173 ;
  assign n3175 = ~\pi0087  & ~n3174 ;
  assign n3176 = ~n3169 & n3175 ;
  assign n3177 = ~n3149 & n3176 ;
  assign n3178 = ~n1288 & ~n3086 ;
  assign n3179 = n1288 & n3061 ;
  assign n3180 = \pi0100  & ~n3179 ;
  assign n3181 = ~n3178 & n3180 ;
  assign n3182 = ~\pi0252  & n1281 ;
  assign n3183 = n1260 & n3182 ;
  assign n3184 = \pi0146  & ~n3183 ;
  assign n3185 = ~\pi0284  & ~n2240 ;
  assign n3186 = n1281 & n3185 ;
  assign n3187 = n1260 & n3186 ;
  assign n3188 = ~\pi0228  & ~n3187 ;
  assign n3189 = ~n3184 & n3188 ;
  assign n3190 = n3106 & ~n3189 ;
  assign n3191 = n3098 & ~n3190 ;
  assign n3192 = n2960 & ~n3094 ;
  assign n3193 = ~n3178 & n3192 ;
  assign n3194 = ~n3191 & n3193 ;
  assign n3195 = ~n3181 & ~n3194 ;
  assign n3196 = ~\pi0087  & ~n3195 ;
  assign n3197 = ~n2328 & ~n3086 ;
  assign n3198 = \pi0087  & ~n3197 ;
  assign n3199 = ~\pi0075  & ~n3198 ;
  assign n3200 = ~\pi0075  & n3110 ;
  assign n3201 = ~n3109 & n3200 ;
  assign n3202 = ~n3199 & ~n3201 ;
  assign n3203 = ~n3196 & ~n3202 ;
  assign n3204 = ~n3177 & n3203 ;
  assign n3205 = \pi0075  & n3061 ;
  assign n3206 = ~\pi0092  & ~n3205 ;
  assign n3207 = n2633 & ~n3172 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = ~n3114 & ~n3208 ;
  assign n3210 = ~n3204 & n3209 ;
  assign n3211 = ~n3115 & ~n3210 ;
  assign n3212 = ~n2407 & ~n3083 ;
  assign n3213 = \pi0056  & n3212 ;
  assign n3214 = n3082 & n3213 ;
  assign n3215 = ~\pi0062  & ~n2406 ;
  assign n3216 = ~\pi0062  & ~n3094 ;
  assign n3217 = ~n3108 & n3216 ;
  assign n3218 = ~n3215 & ~n3217 ;
  assign n3219 = ~n3214 & ~n3218 ;
  assign n3220 = ~\pi0055  & n3219 ;
  assign n3221 = ~n3211 & n3220 ;
  assign n3222 = ~n1291 & ~n3083 ;
  assign n3223 = ~\pi0056  & n3222 ;
  assign n3224 = n3082 & n3223 ;
  assign n3225 = ~n2423 & ~n3224 ;
  assign n3226 = ~n3008 & n3225 ;
  assign n3227 = ~n3094 & n3225 ;
  assign n3228 = ~n3108 & n3227 ;
  assign n3229 = ~n3226 & ~n3228 ;
  assign n3230 = n3219 & ~n3229 ;
  assign n3231 = ~\pi0238  & n2467 ;
  assign n3232 = ~n2504 & ~n3083 ;
  assign n3233 = n3082 & n3232 ;
  assign n3234 = \pi0062  & ~n3233 ;
  assign n3235 = ~n2454 & n3234 ;
  assign n3236 = ~n3094 & n3234 ;
  assign n3237 = ~n3108 & n3236 ;
  assign n3238 = ~n3235 & ~n3237 ;
  assign n3239 = n3231 & n3238 ;
  assign n3240 = ~n3230 & n3239 ;
  assign n3241 = ~n3221 & n3240 ;
  assign n3242 = ~\pi0146  & \pi0284  ;
  assign n3243 = n2718 & n3242 ;
  assign n3244 = ~\pi0146  & ~n2718 ;
  assign n3245 = \pi0284  & ~n3244 ;
  assign n3246 = n1640 & ~n2591 ;
  assign n3247 = n3245 & n3246 ;
  assign n3248 = ~n2704 & n3247 ;
  assign n3249 = ~n3243 & ~n3248 ;
  assign n3250 = ~\pi0146  & ~\pi0284  ;
  assign n3251 = ~n3125 & n3250 ;
  assign n3252 = n3249 & ~n3251 ;
  assign n3253 = n2492 & ~n3252 ;
  assign n3254 = n2225 & ~n3132 ;
  assign n3255 = n2709 & ~n3075 ;
  assign n3256 = ~n3254 & ~n3255 ;
  assign n3257 = ~\pi0095  & ~n3254 ;
  assign n3258 = n2686 & n3257 ;
  assign n3259 = ~n3256 & ~n3258 ;
  assign n3260 = ~\pi0216  & n3259 ;
  assign n3261 = n3130 & ~n3260 ;
  assign n3262 = ~n3253 & n3261 ;
  assign n3263 = n3079 & ~n3104 ;
  assign n3264 = ~n3103 & n3263 ;
  assign n3265 = n3098 & ~n3264 ;
  assign n3266 = n3143 & ~n3265 ;
  assign n3267 = \pi0039  & n3044 ;
  assign n3268 = \pi0039  & n3058 ;
  assign n3269 = ~n3057 & n3268 ;
  assign n3270 = ~n3267 & ~n3269 ;
  assign n3271 = ~\pi0038  & n3270 ;
  assign n3272 = ~n3266 & n3271 ;
  assign n3273 = n3142 & n3272 ;
  assign n3274 = ~n3262 & n3273 ;
  assign n3275 = ~\pi0039  & ~n3150 ;
  assign n3276 = n2692 & ~n3162 ;
  assign n3277 = ~n3275 & ~n3276 ;
  assign n3278 = n3272 & n3277 ;
  assign n3279 = ~n3057 & n3058 ;
  assign n3280 = \pi0038  & ~n3044 ;
  assign n3281 = ~n3279 & n3280 ;
  assign n3282 = ~\pi0299  & n3281 ;
  assign n3283 = n2651 & n3130 ;
  assign n3284 = ~n3083 & ~n3283 ;
  assign n3285 = n3281 & n3284 ;
  assign n3286 = n3082 & n3285 ;
  assign n3287 = ~n3282 & ~n3286 ;
  assign n3288 = n2362 & n3287 ;
  assign n3289 = ~n3278 & n3288 ;
  assign n3290 = ~n3274 & n3289 ;
  assign n3291 = n3095 & ~n3265 ;
  assign n3292 = ~n3044 & ~n3279 ;
  assign n3293 = n2328 & n3292 ;
  assign n3294 = ~n3291 & n3293 ;
  assign n3295 = ~n2328 & ~n3044 ;
  assign n3296 = ~n3279 & n3295 ;
  assign n3297 = ~\pi0299  & n3296 ;
  assign n3298 = n3284 & n3296 ;
  assign n3299 = n3082 & n3298 ;
  assign n3300 = ~n3297 & ~n3299 ;
  assign n3301 = \pi0087  & n3300 ;
  assign n3302 = ~n3294 & n3301 ;
  assign n3303 = ~\pi0075  & ~n3302 ;
  assign n3304 = ~n1286 & ~n3044 ;
  assign n3305 = ~n3279 & n3304 ;
  assign n3306 = ~\pi0299  & n3305 ;
  assign n3307 = n3284 & n3305 ;
  assign n3308 = n3082 & n3307 ;
  assign n3309 = ~n3306 & ~n3308 ;
  assign n3310 = \pi0092  & n3309 ;
  assign n3311 = n3300 & n3310 ;
  assign n3312 = ~n3294 & n3311 ;
  assign n3313 = n2387 & n3309 ;
  assign n3314 = n2511 & ~n3313 ;
  assign n3315 = ~n3312 & n3314 ;
  assign n3316 = ~n1288 & ~n3044 ;
  assign n3317 = ~n3279 & n3316 ;
  assign n3318 = ~\pi0299  & n3317 ;
  assign n3319 = n3284 & n3317 ;
  assign n3320 = n3082 & n3319 ;
  assign n3321 = ~n3318 & ~n3320 ;
  assign n3322 = n1288 & ~n3044 ;
  assign n3323 = ~n3279 & n3322 ;
  assign n3324 = \pi0100  & ~n3323 ;
  assign n3325 = n3321 & n3324 ;
  assign n3326 = ~n3189 & n3263 ;
  assign n3327 = n3098 & ~n3326 ;
  assign n3328 = n3192 & n3321 ;
  assign n3329 = ~n3327 & n3328 ;
  assign n3330 = ~n3325 & ~n3329 ;
  assign n3331 = ~\pi0087  & ~n3330 ;
  assign n3332 = n3315 & ~n3331 ;
  assign n3333 = n3303 & n3332 ;
  assign n3334 = ~n3290 & n3333 ;
  assign n3335 = \pi0075  & ~n3044 ;
  assign n3336 = ~n3279 & n3335 ;
  assign n3337 = ~\pi0299  & n3336 ;
  assign n3338 = n3284 & n3336 ;
  assign n3339 = n3082 & n3338 ;
  assign n3340 = ~n3337 & ~n3339 ;
  assign n3341 = ~\pi0092  & n3340 ;
  assign n3342 = n3314 & ~n3341 ;
  assign n3343 = ~n3312 & n3342 ;
  assign n3344 = ~n2407 & n3284 ;
  assign n3345 = n3082 & n3344 ;
  assign n3346 = ~\pi0062  & ~n3345 ;
  assign n3347 = ~n3030 & n3346 ;
  assign n3348 = ~n3094 & n3346 ;
  assign n3349 = ~n3265 & n3348 ;
  assign n3350 = ~n3347 & ~n3349 ;
  assign n3351 = ~n1292 & n3350 ;
  assign n3352 = ~n2511 & ~n3044 ;
  assign n3353 = ~n3279 & n3352 ;
  assign n3354 = ~\pi0299  & n3353 ;
  assign n3355 = n3284 & n3353 ;
  assign n3356 = n3082 & n3355 ;
  assign n3357 = ~n3354 & ~n3356 ;
  assign n3358 = ~\pi0055  & n3357 ;
  assign n3359 = ~n3351 & n3358 ;
  assign n3360 = ~n3343 & n3359 ;
  assign n3361 = ~n3334 & n3360 ;
  assign n3362 = n3222 & ~n3283 ;
  assign n3363 = ~\pi0056  & n3362 ;
  assign n3364 = n3082 & n3363 ;
  assign n3365 = ~n2423 & ~n3364 ;
  assign n3366 = ~n3008 & n3365 ;
  assign n3367 = ~n3094 & n3365 ;
  assign n3368 = ~n3265 & n3367 ;
  assign n3369 = ~n3366 & ~n3368 ;
  assign n3370 = ~n3351 & ~n3369 ;
  assign n3371 = \pi0238  & n2467 ;
  assign n3372 = ~n2504 & n3284 ;
  assign n3373 = n3082 & n3372 ;
  assign n3374 = \pi0062  & ~n3373 ;
  assign n3375 = ~n2504 & n3374 ;
  assign n3376 = ~n3094 & n3374 ;
  assign n3377 = ~n3265 & n3376 ;
  assign n3378 = ~n3375 & ~n3377 ;
  assign n3379 = n3371 & n3378 ;
  assign n3380 = ~n3370 & n3379 ;
  assign n3381 = ~n3361 & n3380 ;
  assign n3382 = \pi0238  & n3283 ;
  assign n3383 = ~n2467 & ~n3083 ;
  assign n3384 = ~n3382 & n3383 ;
  assign n3385 = n3082 & n3384 ;
  assign n3386 = ~n3381 & ~n3385 ;
  assign n3387 = ~n3241 & n3386 ;
  assign n3388 = \pi0105  & \pi0262  ;
  assign n3389 = ~n1633 & n3388 ;
  assign n3390 = ~\pi0105  & \pi0172  ;
  assign n3391 = \pi0172  & ~\pi0228  ;
  assign n3392 = ~n3390 & ~n3391 ;
  assign n3393 = ~n3389 & n3392 ;
  assign n3394 = \pi0221  & \pi0932  ;
  assign n3395 = n1220 & ~n3394 ;
  assign n3396 = \pi0221  & \pi1142  ;
  assign n3397 = ~\pi0216  & ~\pi0833  ;
  assign n3398 = ~n3396 & n3397 ;
  assign n3399 = ~n3395 & ~n3398 ;
  assign n3400 = ~\pi0172  & ~\pi0228  ;
  assign n3401 = ~n3399 & ~n3400 ;
  assign n3402 = ~n3393 & n3401 ;
  assign n3403 = \pi0216  & \pi0277  ;
  assign n3404 = ~\pi0221  & ~n3403 ;
  assign n3405 = ~n1220 & n3396 ;
  assign n3406 = n1220 & n3394 ;
  assign n3407 = ~n3405 & ~n3406 ;
  assign n3408 = ~n3404 & n3407 ;
  assign n3409 = ~\pi0215  & ~n2652 ;
  assign n3410 = ~n3408 & n3409 ;
  assign n3411 = ~n3402 & n3410 ;
  assign n3412 = \pi0215  & \pi1142  ;
  assign n3413 = ~n2467 & ~n3412 ;
  assign n3414 = ~n3411 & n3413 ;
  assign n3415 = ~\pi0249  & ~n3414 ;
  assign n3416 = ~n2504 & ~n3412 ;
  assign n3417 = ~n3411 & n3416 ;
  assign n3418 = \pi0062  & ~n3417 ;
  assign n3419 = n2467 & ~n3418 ;
  assign n3420 = ~\pi0228  & n1281 ;
  assign n3421 = n1260 & n3420 ;
  assign n3422 = ~n3389 & ~n3390 ;
  assign n3423 = \pi0228  & ~n3422 ;
  assign n3424 = ~n2651 & ~n3391 ;
  assign n3425 = ~n3423 & n3424 ;
  assign n3426 = ~n3421 & n3425 ;
  assign n3427 = ~n2651 & ~n3423 ;
  assign n3428 = ~\pi0262  & n1281 ;
  assign n3429 = n1260 & n3428 ;
  assign n3430 = n3427 & n3429 ;
  assign n3431 = ~n3399 & ~n3430 ;
  assign n3432 = ~n3426 & n3431 ;
  assign n3433 = ~\pi0215  & ~n3408 ;
  assign n3434 = ~n3432 & n3433 ;
  assign n3435 = ~\pi0056  & ~n3412 ;
  assign n3436 = n2404 & n3435 ;
  assign n3437 = n2403 & n3436 ;
  assign n3438 = n2467 & n3437 ;
  assign n3439 = ~n3434 & n3438 ;
  assign n3440 = ~n3419 & ~n3439 ;
  assign n3441 = ~n1291 & ~n3412 ;
  assign n3442 = ~n3411 & n3441 ;
  assign n3443 = \pi0055  & ~n3442 ;
  assign n3444 = ~\pi0056  & ~n3443 ;
  assign n3445 = n1291 & ~n3412 ;
  assign n3446 = ~\pi0056  & n3445 ;
  assign n3447 = ~n3434 & n3446 ;
  assign n3448 = ~n3444 & ~n3447 ;
  assign n3449 = ~n2407 & ~n3412 ;
  assign n3450 = ~n3411 & n3449 ;
  assign n3451 = ~\pi0062  & ~n3450 ;
  assign n3452 = ~n1292 & ~n3451 ;
  assign n3453 = n2404 & ~n3412 ;
  assign n3454 = n2403 & n3453 ;
  assign n3455 = ~n1292 & n3454 ;
  assign n3456 = ~n3434 & n3455 ;
  assign n3457 = ~n3452 & ~n3456 ;
  assign n3458 = n3448 & n3457 ;
  assign n3459 = \pi0223  & \pi1142  ;
  assign n3460 = ~\pi0299  & n3459 ;
  assign n3461 = ~n3045 & n3460 ;
  assign n3462 = \pi0224  & \pi0277  ;
  assign n3463 = ~\pi0222  & ~n3462 ;
  assign n3464 = ~\pi0224  & \pi0262  ;
  assign n3465 = ~n1633 & n3464 ;
  assign n3466 = n3463 & ~n3465 ;
  assign n3467 = \pi0222  & \pi0932  ;
  assign n3468 = n2192 & n3467 ;
  assign n3469 = \pi0222  & \pi1142  ;
  assign n3470 = ~n2192 & n3469 ;
  assign n3471 = ~n3468 & ~n3470 ;
  assign n3472 = ~n3466 & n3471 ;
  assign n3473 = n3059 & ~n3472 ;
  assign n3474 = ~n3461 & ~n3473 ;
  assign n3475 = \pi0075  & n3474 ;
  assign n3476 = ~\pi0092  & ~n3475 ;
  assign n3477 = ~n3411 & ~n3412 ;
  assign n3478 = n2633 & ~n3477 ;
  assign n3479 = ~n3476 & ~n3478 ;
  assign n3480 = n2328 & n3474 ;
  assign n3481 = ~\pi0299  & n3480 ;
  assign n3482 = ~n3412 & n3480 ;
  assign n3483 = ~n3434 & n3482 ;
  assign n3484 = ~n3481 & ~n3483 ;
  assign n3485 = \pi0299  & ~n3477 ;
  assign n3486 = ~n2328 & n3474 ;
  assign n3487 = ~n3485 & n3486 ;
  assign n3488 = ~n1286 & n3474 ;
  assign n3489 = \pi0092  & ~n3488 ;
  assign n3490 = n3003 & ~n3477 ;
  assign n3491 = ~n3489 & ~n3490 ;
  assign n3492 = ~n3487 & ~n3491 ;
  assign n3493 = n3484 & n3492 ;
  assign n3494 = ~n1286 & ~n3491 ;
  assign n3495 = n2511 & ~n3494 ;
  assign n3496 = ~n3493 & n3495 ;
  assign n3497 = n3479 & n3496 ;
  assign n3498 = \pi0223  & ~\pi0299  ;
  assign n3499 = ~\pi1142  & n3498 ;
  assign n3500 = ~n3463 & n3471 ;
  assign n3501 = ~\pi0262  & ~n1633 ;
  assign n3502 = n2192 & ~n3467 ;
  assign n3503 = ~\pi0224  & ~\pi0833  ;
  assign n3504 = ~n3469 & n3503 ;
  assign n3505 = ~n3502 & ~n3504 ;
  assign n3506 = ~n3501 & ~n3505 ;
  assign n3507 = ~\pi0095  & ~n3505 ;
  assign n3508 = n2686 & n3507 ;
  assign n3509 = ~n3506 & ~n3508 ;
  assign n3510 = ~n3500 & n3509 ;
  assign n3511 = ~\pi0299  & ~n3459 ;
  assign n3512 = n1633 & n3463 ;
  assign n3513 = ~\pi0095  & n3463 ;
  assign n3514 = n2686 & n3513 ;
  assign n3515 = ~n3512 & ~n3514 ;
  assign n3516 = n3511 & n3515 ;
  assign n3517 = ~n3510 & n3516 ;
  assign n3518 = ~n3499 & ~n3517 ;
  assign n3519 = ~\pi0039  & ~n3511 ;
  assign n3520 = ~\pi0039  & ~n3500 ;
  assign n3521 = n3509 & n3520 ;
  assign n3522 = ~n3519 & ~n3521 ;
  assign n3523 = n3518 & ~n3522 ;
  assign n3524 = ~n2943 & n3425 ;
  assign n3525 = ~\pi0262  & n3427 ;
  assign n3526 = ~n2618 & n3525 ;
  assign n3527 = ~n2615 & n3526 ;
  assign n3528 = ~n3399 & ~n3527 ;
  assign n3529 = ~n3524 & n3528 ;
  assign n3530 = n2256 & ~n3408 ;
  assign n3531 = ~n3529 & n3530 ;
  assign n3532 = \pi0299  & n3412 ;
  assign n3533 = n1288 & n3474 ;
  assign n3534 = ~n3532 & n3533 ;
  assign n3535 = ~n3531 & n3534 ;
  assign n3536 = ~n1288 & n3474 ;
  assign n3537 = \pi0100  & ~n3536 ;
  assign n3538 = n2960 & ~n3477 ;
  assign n3539 = ~n3537 & ~n3538 ;
  assign n3540 = ~n3535 & ~n3539 ;
  assign n3541 = ~\pi0038  & n3474 ;
  assign n3542 = ~\pi0299  & n3541 ;
  assign n3543 = ~n3412 & n3541 ;
  assign n3544 = ~n3434 & n3543 ;
  assign n3545 = ~n3542 & ~n3544 ;
  assign n3546 = ~n1288 & n3545 ;
  assign n3547 = ~n3540 & ~n3546 ;
  assign n3548 = ~n3523 & n3547 ;
  assign n3549 = ~\pi0262  & n1640 ;
  assign n3550 = ~n2591 & n3549 ;
  assign n3551 = ~n2704 & n3550 ;
  assign n3552 = \pi0172  & ~n3551 ;
  assign n3553 = \pi0105  & n1633 ;
  assign n3554 = ~\pi0095  & \pi0105  ;
  assign n3555 = n2686 & n3554 ;
  assign n3556 = ~n3553 & ~n3555 ;
  assign n3557 = \pi0228  & ~n3390 ;
  assign n3558 = ~n3389 & n3557 ;
  assign n3559 = ~\pi0095  & n3557 ;
  assign n3560 = n2686 & n3559 ;
  assign n3561 = ~n3558 & ~n3560 ;
  assign n3562 = n3556 & ~n3561 ;
  assign n3563 = ~\pi0216  & n3407 ;
  assign n3564 = ~n3562 & n3563 ;
  assign n3565 = n3552 & n3564 ;
  assign n3566 = \pi0262  & n2591 ;
  assign n3567 = \pi0262  & ~n2580 ;
  assign n3568 = n2574 & n3567 ;
  assign n3569 = ~n3566 & ~n3568 ;
  assign n3570 = ~\pi0228  & ~n3569 ;
  assign n3571 = ~n2716 & n3501 ;
  assign n3572 = ~\pi0172  & ~n1639 ;
  assign n3573 = ~n3571 & n3572 ;
  assign n3574 = ~\pi0228  & ~n3573 ;
  assign n3575 = n3564 & ~n3574 ;
  assign n3576 = ~n3570 & n3575 ;
  assign n3577 = ~n3565 & ~n3576 ;
  assign n3578 = n3433 & n3577 ;
  assign n3579 = \pi0299  & ~n3412 ;
  assign n3580 = n3547 & n3579 ;
  assign n3581 = ~n3578 & n3580 ;
  assign n3582 = ~n3548 & ~n3581 ;
  assign n3583 = \pi0038  & n3474 ;
  assign n3584 = ~\pi0100  & ~n3583 ;
  assign n3585 = n2563 & ~n3477 ;
  assign n3586 = ~n3584 & ~n3585 ;
  assign n3587 = ~n3540 & n3586 ;
  assign n3588 = ~\pi0087  & ~n3587 ;
  assign n3589 = n3582 & n3588 ;
  assign n3590 = \pi0087  & ~n3486 ;
  assign n3591 = \pi0087  & \pi0299  ;
  assign n3592 = ~n3477 & n3591 ;
  assign n3593 = ~n3590 & ~n3592 ;
  assign n3594 = n3484 & ~n3593 ;
  assign n3595 = ~\pi0075  & ~n3594 ;
  assign n3596 = n3496 & n3595 ;
  assign n3597 = ~n3589 & n3596 ;
  assign n3598 = ~n3497 & ~n3597 ;
  assign n3599 = ~n2511 & n3474 ;
  assign n3600 = ~\pi0055  & ~n3599 ;
  assign n3601 = n3026 & ~n3477 ;
  assign n3602 = ~n3600 & ~n3601 ;
  assign n3603 = n3457 & ~n3602 ;
  assign n3604 = n3598 & n3603 ;
  assign n3605 = ~n3458 & ~n3604 ;
  assign n3606 = ~n3440 & n3605 ;
  assign n3607 = n3415 & ~n3606 ;
  assign n3608 = ~n3402 & n3433 ;
  assign n3609 = n3416 & ~n3608 ;
  assign n3610 = \pi0062  & ~n3609 ;
  assign n3611 = n2467 & ~n3610 ;
  assign n3612 = ~\pi0228  & ~n3391 ;
  assign n3613 = ~n3393 & ~n3612 ;
  assign n3614 = ~n3421 & ~n3613 ;
  assign n3615 = n1259 & ~n3423 ;
  assign n3616 = n1249 & n3615 ;
  assign n3617 = n3428 & n3616 ;
  assign n3618 = ~n3399 & ~n3617 ;
  assign n3619 = ~n3614 & n3618 ;
  assign n3620 = n3433 & ~n3619 ;
  assign n3621 = n3438 & ~n3620 ;
  assign n3622 = ~n3611 & ~n3621 ;
  assign n3623 = n3413 & ~n3608 ;
  assign n3624 = \pi0249  & ~n3623 ;
  assign n3625 = n3622 & n3624 ;
  assign n3626 = ~n3402 & n3530 ;
  assign n3627 = ~n3532 & ~n3626 ;
  assign n3628 = n3058 & ~n3472 ;
  assign n3629 = ~n2511 & ~n3460 ;
  assign n3630 = ~n3628 & n3629 ;
  assign n3631 = n3627 & n3630 ;
  assign n3632 = ~\pi0055  & ~n3631 ;
  assign n3633 = n3441 & ~n3608 ;
  assign n3634 = \pi0055  & ~n3633 ;
  assign n3635 = ~\pi0056  & ~n3634 ;
  assign n3636 = n3446 & ~n3620 ;
  assign n3637 = ~n3635 & ~n3636 ;
  assign n3638 = ~n3632 & ~n3637 ;
  assign n3639 = n3530 & ~n3619 ;
  assign n3640 = n2328 & ~n3460 ;
  assign n3641 = ~n3628 & n3640 ;
  assign n3642 = ~n3532 & n3641 ;
  assign n3643 = ~n3639 & n3642 ;
  assign n3644 = ~n3460 & ~n3628 ;
  assign n3645 = ~n2328 & ~n3532 ;
  assign n3646 = ~n3626 & n3645 ;
  assign n3647 = n3644 & n3646 ;
  assign n3648 = \pi0087  & ~n3647 ;
  assign n3649 = ~n3643 & n3648 ;
  assign n3650 = ~\pi0075  & ~n3649 ;
  assign n3651 = \pi0075  & ~n3532 ;
  assign n3652 = ~n3626 & n3651 ;
  assign n3653 = n3644 & n3652 ;
  assign n3654 = ~\pi0092  & ~n3653 ;
  assign n3655 = ~n3650 & n3654 ;
  assign n3656 = \pi0262  & n1640 ;
  assign n3657 = ~n2591 & n3656 ;
  assign n3658 = ~n2704 & n3657 ;
  assign n3659 = ~\pi0172  & ~n3658 ;
  assign n3660 = \pi0262  & n2718 ;
  assign n3661 = \pi0172  & ~n3660 ;
  assign n3662 = n3124 & n3661 ;
  assign n3663 = ~n2581 & n3662 ;
  assign n3664 = \pi0172  & \pi0262  ;
  assign n3665 = ~n2718 & n3664 ;
  assign n3666 = ~n3663 & ~n3665 ;
  assign n3667 = ~n3659 & n3666 ;
  assign n3668 = ~\pi0221  & ~\pi0228  ;
  assign n3669 = ~n3403 & n3668 ;
  assign n3670 = ~n3667 & n3669 ;
  assign n3671 = ~\pi0216  & n3561 ;
  assign n3672 = n3404 & ~n3671 ;
  assign n3673 = n3407 & n3579 ;
  assign n3674 = ~n3672 & n3673 ;
  assign n3675 = ~n3670 & n3674 ;
  assign n3676 = ~\pi1142  & n2259 ;
  assign n3677 = \pi0038  & ~n3532 ;
  assign n3678 = ~n3626 & n3677 ;
  assign n3679 = n3644 & n3678 ;
  assign n3680 = n2320 & ~n3499 ;
  assign n3681 = ~n3679 & n3680 ;
  assign n3682 = ~n3517 & n3681 ;
  assign n3683 = ~n3676 & n3682 ;
  assign n3684 = ~n3675 & n3683 ;
  assign n3685 = ~\pi0038  & ~n3532 ;
  assign n3686 = n3644 & n3685 ;
  assign n3687 = ~n3639 & n3686 ;
  assign n3688 = ~\pi0100  & ~n1288 ;
  assign n3689 = ~n3679 & n3688 ;
  assign n3690 = ~n3687 & n3689 ;
  assign n3691 = ~n2943 & ~n3613 ;
  assign n3692 = ~\pi0262  & ~n3423 ;
  assign n3693 = ~n2618 & n3692 ;
  assign n3694 = ~n2615 & n3693 ;
  assign n3695 = ~n3399 & ~n3694 ;
  assign n3696 = ~n3691 & n3695 ;
  assign n3697 = n3530 & ~n3696 ;
  assign n3698 = n1288 & ~n3532 ;
  assign n3699 = n3644 & n3698 ;
  assign n3700 = ~n3697 & n3699 ;
  assign n3701 = ~n1288 & ~n3460 ;
  assign n3702 = ~n3628 & n3701 ;
  assign n3703 = n3627 & n3702 ;
  assign n3704 = \pi0100  & ~n3703 ;
  assign n3705 = ~n3700 & n3704 ;
  assign n3706 = ~n3690 & ~n3705 ;
  assign n3707 = ~n3684 & n3706 ;
  assign n3708 = ~\pi0087  & n3654 ;
  assign n3709 = ~n3707 & n3708 ;
  assign n3710 = ~n3655 & ~n3709 ;
  assign n3711 = ~n1286 & ~n3460 ;
  assign n3712 = ~n3628 & n3711 ;
  assign n3713 = n3627 & n3712 ;
  assign n3714 = \pi0092  & ~n3713 ;
  assign n3715 = ~n3647 & n3714 ;
  assign n3716 = ~n3643 & n3715 ;
  assign n3717 = n2387 & ~n3713 ;
  assign n3718 = n2511 & ~n3717 ;
  assign n3719 = ~n3716 & n3718 ;
  assign n3720 = ~n3637 & n3719 ;
  assign n3721 = n3710 & n3720 ;
  assign n3722 = ~n3638 & ~n3721 ;
  assign n3723 = n3449 & ~n3608 ;
  assign n3724 = \pi0056  & n3723 ;
  assign n3725 = \pi0056  & n3454 ;
  assign n3726 = ~n3620 & n3725 ;
  assign n3727 = ~n3724 & ~n3726 ;
  assign n3728 = ~\pi0062  & n3727 ;
  assign n3729 = n3624 & n3728 ;
  assign n3730 = n3722 & n3729 ;
  assign n3731 = ~n3625 & ~n3730 ;
  assign n3732 = ~n3607 & n3731 ;
  assign n3733 = \pi0216  & \pi0270  ;
  assign n3734 = ~\pi0221  & ~n3733 ;
  assign n3735 = \pi0221  & \pi1141  ;
  assign n3736 = ~n1220 & n3735 ;
  assign n3737 = \pi0221  & \pi0935  ;
  assign n3738 = n1220 & n3737 ;
  assign n3739 = ~n3736 & ~n3738 ;
  assign n3740 = ~n3734 & n3739 ;
  assign n3741 = ~\pi0215  & ~n3740 ;
  assign n3742 = ~\pi0105  & \pi0171  ;
  assign n3743 = \pi0228  & ~n3742 ;
  assign n3744 = ~\pi0216  & ~n3743 ;
  assign n3745 = \pi0861  & ~n1633 ;
  assign n3746 = \pi0105  & ~\pi0216  ;
  assign n3747 = ~n3745 & n3746 ;
  assign n3748 = ~n3744 & ~n3747 ;
  assign n3749 = ~\pi0171  & ~\pi0228  ;
  assign n3750 = n3739 & ~n3749 ;
  assign n3751 = ~n3748 & n3750 ;
  assign n3752 = n3741 & ~n3751 ;
  assign n3753 = \pi0215  & \pi1141  ;
  assign n3754 = n1295 & ~n3733 ;
  assign n3755 = n2651 & n3754 ;
  assign n3756 = ~n3753 & ~n3755 ;
  assign n3757 = ~n3752 & n3756 ;
  assign n3758 = \pi0299  & ~n3757 ;
  assign n3759 = \pi0222  & \pi1141  ;
  assign n3760 = ~n2192 & n3759 ;
  assign n3761 = \pi0222  & \pi0935  ;
  assign n3762 = n2192 & n3761 ;
  assign n3763 = ~n3760 & ~n3762 ;
  assign n3764 = ~\pi0223  & ~n3763 ;
  assign n3765 = ~\pi0224  & ~n3745 ;
  assign n3766 = \pi0224  & \pi0270  ;
  assign n3767 = ~\pi0222  & ~n3766 ;
  assign n3768 = ~\pi0223  & n3767 ;
  assign n3769 = ~n3765 & n3768 ;
  assign n3770 = ~n3764 & ~n3769 ;
  assign n3771 = \pi0223  & \pi1141  ;
  assign n3772 = ~n3045 & ~n3771 ;
  assign n3773 = n3770 & n3772 ;
  assign n3774 = ~\pi0299  & ~n3773 ;
  assign n3775 = ~n2511 & ~n3774 ;
  assign n3776 = ~n3758 & n3775 ;
  assign n3777 = ~\pi0055  & ~n3776 ;
  assign n3778 = \pi0171  & ~n2280 ;
  assign n3779 = ~\pi0861  & n1281 ;
  assign n3780 = n1260 & n3779 ;
  assign n3781 = ~\pi0228  & ~n3780 ;
  assign n3782 = ~n3778 & n3781 ;
  assign n3783 = ~n2651 & n3739 ;
  assign n3784 = ~n3748 & n3783 ;
  assign n3785 = ~n3782 & n3784 ;
  assign n3786 = n3741 & ~n3785 ;
  assign n3787 = n1291 & ~n3753 ;
  assign n3788 = ~n3786 & n3787 ;
  assign n3789 = ~n1291 & ~n3753 ;
  assign n3790 = ~n3755 & n3789 ;
  assign n3791 = ~n3752 & n3790 ;
  assign n3792 = \pi0055  & ~n3791 ;
  assign n3793 = ~n3788 & n3792 ;
  assign n3794 = ~n3777 & ~n3793 ;
  assign n3795 = n2328 & ~n3774 ;
  assign n3796 = ~\pi0299  & n3795 ;
  assign n3797 = ~n3753 & n3795 ;
  assign n3798 = ~n3786 & n3797 ;
  assign n3799 = ~n3796 & ~n3798 ;
  assign n3800 = ~n2328 & ~n3774 ;
  assign n3801 = ~n3758 & n3800 ;
  assign n3802 = \pi0087  & ~n3801 ;
  assign n3803 = n3799 & n3802 ;
  assign n3804 = ~\pi0075  & ~n3803 ;
  assign n3805 = \pi0075  & ~n3774 ;
  assign n3806 = ~n3758 & n3805 ;
  assign n3807 = ~\pi0092  & ~n3806 ;
  assign n3808 = ~n3804 & n3807 ;
  assign n3809 = \pi0038  & ~n3774 ;
  assign n3810 = ~n3758 & n3809 ;
  assign n3811 = ~\pi0100  & ~n3810 ;
  assign n3812 = ~n1288 & ~n3774 ;
  assign n3813 = ~n3758 & n3812 ;
  assign n3814 = n1288 & ~n3774 ;
  assign n3815 = \pi0100  & ~n3814 ;
  assign n3816 = ~n3813 & n3815 ;
  assign n3817 = ~n2651 & ~n3748 ;
  assign n3818 = n3734 & ~n3817 ;
  assign n3819 = ~\pi0861  & ~n2618 ;
  assign n3820 = ~n2615 & n3819 ;
  assign n3821 = ~\pi0228  & ~n3820 ;
  assign n3822 = \pi0171  & n2618 ;
  assign n3823 = \pi0171  & ~n2609 ;
  assign n3824 = n2614 & n3823 ;
  assign n3825 = ~n3822 & ~n3824 ;
  assign n3826 = n3734 & n3825 ;
  assign n3827 = n3821 & n3826 ;
  assign n3828 = ~n3818 & ~n3827 ;
  assign n3829 = n3739 & ~n3753 ;
  assign n3830 = n3828 & n3829 ;
  assign n3831 = \pi0215  & ~\pi1141  ;
  assign n3832 = n2960 & ~n3831 ;
  assign n3833 = ~n3813 & n3832 ;
  assign n3834 = ~n3830 & n3833 ;
  assign n3835 = ~n3816 & ~n3834 ;
  assign n3836 = ~n3811 & n3835 ;
  assign n3837 = ~\pi0861  & n1640 ;
  assign n3838 = ~n2591 & n3837 ;
  assign n3839 = ~n2704 & n3838 ;
  assign n3840 = ~\pi0171  & ~n3839 ;
  assign n3841 = ~\pi0861  & n2718 ;
  assign n3842 = \pi0171  & ~n3841 ;
  assign n3843 = n3124 & n3842 ;
  assign n3844 = ~n2581 & n3843 ;
  assign n3845 = \pi0171  & ~\pi0861  ;
  assign n3846 = ~n2718 & n3845 ;
  assign n3847 = ~n3844 & ~n3846 ;
  assign n3848 = ~n3840 & n3847 ;
  assign n3849 = n3668 & ~n3733 ;
  assign n3850 = ~n3848 & n3849 ;
  assign n3851 = ~\pi0095  & n1209 ;
  assign n3852 = n2686 & n3851 ;
  assign n3853 = ~n2651 & ~n3852 ;
  assign n3854 = ~n3748 & n3853 ;
  assign n3855 = n3734 & ~n3854 ;
  assign n3856 = \pi0299  & ~n3753 ;
  assign n3857 = n3739 & n3856 ;
  assign n3858 = ~n3855 & n3857 ;
  assign n3859 = ~n3850 & n3858 ;
  assign n3860 = ~\pi1141  & n2259 ;
  assign n3861 = n3763 & ~n3767 ;
  assign n3862 = n2192 & ~n3761 ;
  assign n3863 = n3503 & ~n3759 ;
  assign n3864 = ~n3862 & ~n3863 ;
  assign n3865 = ~n3745 & ~n3864 ;
  assign n3866 = ~\pi0095  & ~n3864 ;
  assign n3867 = n2686 & n3866 ;
  assign n3868 = ~n3865 & ~n3867 ;
  assign n3869 = ~n3861 & n3868 ;
  assign n3870 = ~\pi0299  & ~n3771 ;
  assign n3871 = n1633 & n3767 ;
  assign n3872 = ~\pi0095  & n3767 ;
  assign n3873 = n2686 & n3872 ;
  assign n3874 = ~n3871 & ~n3873 ;
  assign n3875 = n3870 & n3874 ;
  assign n3876 = ~n3869 & n3875 ;
  assign n3877 = ~\pi1141  & n3498 ;
  assign n3878 = ~\pi0039  & ~n3877 ;
  assign n3879 = ~n3876 & n3878 ;
  assign n3880 = ~n3860 & n3879 ;
  assign n3881 = ~n3859 & n3880 ;
  assign n3882 = ~\pi0038  & ~n3774 ;
  assign n3883 = ~\pi0299  & n3882 ;
  assign n3884 = ~n3753 & n3882 ;
  assign n3885 = ~n3786 & n3884 ;
  assign n3886 = ~n3883 & ~n3885 ;
  assign n3887 = ~n1288 & n3886 ;
  assign n3888 = n3835 & ~n3887 ;
  assign n3889 = ~n3881 & n3888 ;
  assign n3890 = ~n3836 & ~n3889 ;
  assign n3891 = ~\pi0087  & n3807 ;
  assign n3892 = n3890 & n3891 ;
  assign n3893 = ~n3808 & ~n3892 ;
  assign n3894 = ~n1286 & ~n3774 ;
  assign n3895 = ~n3758 & n3894 ;
  assign n3896 = \pi0092  & ~n3895 ;
  assign n3897 = ~n3801 & n3896 ;
  assign n3898 = n3799 & n3897 ;
  assign n3899 = n2387 & ~n3895 ;
  assign n3900 = n2511 & ~n3899 ;
  assign n3901 = ~n3898 & n3900 ;
  assign n3902 = ~n3793 & n3901 ;
  assign n3903 = n3893 & n3902 ;
  assign n3904 = ~n3794 & ~n3903 ;
  assign n3905 = n2504 & ~n3753 ;
  assign n3906 = ~n3786 & n3905 ;
  assign n3907 = ~n2504 & n3756 ;
  assign n3908 = ~n3752 & n3907 ;
  assign n3909 = \pi0062  & ~n3908 ;
  assign n3910 = ~n3906 & n3909 ;
  assign n3911 = \pi0241  & n2467 ;
  assign n3912 = ~n3910 & n3911 ;
  assign n3913 = ~\pi0056  & n3912 ;
  assign n3914 = ~n3904 & n3913 ;
  assign n3915 = \pi0299  & n2328 ;
  assign n3916 = n2328 & ~n3771 ;
  assign n3917 = n3770 & n3916 ;
  assign n3918 = ~n3915 & ~n3917 ;
  assign n3919 = ~\pi0299  & ~n3918 ;
  assign n3920 = n3739 & ~n3748 ;
  assign n3921 = ~n3782 & n3920 ;
  assign n3922 = n3741 & ~n3921 ;
  assign n3923 = ~n3753 & ~n3918 ;
  assign n3924 = ~n3922 & n3923 ;
  assign n3925 = ~n3919 & ~n3924 ;
  assign n3926 = n3770 & ~n3771 ;
  assign n3927 = ~\pi0299  & n3926 ;
  assign n3928 = ~n3752 & n3856 ;
  assign n3929 = ~n3927 & ~n3928 ;
  assign n3930 = \pi0092  & n3929 ;
  assign n3931 = ~n3089 & ~n3930 ;
  assign n3932 = n3925 & ~n3931 ;
  assign n3933 = n2387 & n3929 ;
  assign n3934 = n2511 & ~n3933 ;
  assign n3935 = ~n3932 & n3934 ;
  assign n3936 = ~n2511 & ~n3929 ;
  assign n3937 = ~\pi0055  & ~n3936 ;
  assign n3938 = n1292 & n3937 ;
  assign n3939 = n2407 & ~n3753 ;
  assign n3940 = ~n3922 & n3939 ;
  assign n3941 = ~n2407 & ~n3753 ;
  assign n3942 = ~n3752 & n3941 ;
  assign n3943 = ~\pi0062  & ~n3942 ;
  assign n3944 = n3937 & n3943 ;
  assign n3945 = ~n3940 & n3944 ;
  assign n3946 = ~n3938 & ~n3945 ;
  assign n3947 = ~n3935 & ~n3946 ;
  assign n3948 = \pi0105  & ~n3745 ;
  assign n3949 = n3743 & ~n3948 ;
  assign n3950 = ~n1633 & n3949 ;
  assign n3951 = ~n2716 & n3950 ;
  assign n3952 = n2225 & ~n3742 ;
  assign n3953 = ~\pi0216  & ~n3952 ;
  assign n3954 = ~n3951 & n3953 ;
  assign n3955 = \pi0171  & n1640 ;
  assign n3956 = ~n2591 & n3955 ;
  assign n3957 = ~n2704 & n3956 ;
  assign n3958 = \pi0861  & n3957 ;
  assign n3959 = ~\pi0228  & n3958 ;
  assign n3960 = ~n2716 & n3745 ;
  assign n3961 = ~n1639 & ~n3960 ;
  assign n3962 = ~\pi0861  & n2591 ;
  assign n3963 = ~\pi0861  & ~n2580 ;
  assign n3964 = n2574 & n3963 ;
  assign n3965 = ~n3962 & ~n3964 ;
  assign n3966 = n3961 & n3965 ;
  assign n3967 = n3749 & ~n3966 ;
  assign n3968 = ~n3959 & ~n3967 ;
  assign n3969 = n3954 & n3968 ;
  assign n3970 = ~\pi0215  & n3734 ;
  assign n3971 = ~n3969 & n3970 ;
  assign n3972 = ~\pi0038  & \pi0299  ;
  assign n3973 = ~\pi0038  & ~n3771 ;
  assign n3974 = n3770 & n3973 ;
  assign n3975 = ~n3972 & ~n3974 ;
  assign n3976 = ~\pi0299  & ~n3975 ;
  assign n3977 = ~n3753 & ~n3975 ;
  assign n3978 = ~n3922 & n3977 ;
  assign n3979 = ~n3976 & ~n3978 ;
  assign n3980 = ~n1288 & n3979 ;
  assign n3981 = ~\pi0215  & ~n3739 ;
  assign n3982 = n3856 & ~n3981 ;
  assign n3983 = ~n3980 & n3982 ;
  assign n3984 = ~n3971 & n3983 ;
  assign n3985 = ~n3869 & n3870 ;
  assign n3986 = n3879 & ~n3985 ;
  assign n3987 = \pi0038  & \pi0299  ;
  assign n3988 = \pi0038  & ~n3771 ;
  assign n3989 = n3770 & n3988 ;
  assign n3990 = ~n3987 & ~n3989 ;
  assign n3991 = ~\pi0100  & n3990 ;
  assign n3992 = ~n3752 & ~n3753 ;
  assign n3993 = n2563 & ~n3992 ;
  assign n3994 = ~n3991 & ~n3993 ;
  assign n3995 = ~\pi0087  & ~n3994 ;
  assign n3996 = n3986 & n3995 ;
  assign n3997 = ~n1288 & n3995 ;
  assign n3998 = n3979 & n3997 ;
  assign n3999 = ~n3996 & ~n3998 ;
  assign n4000 = ~n3984 & ~n3999 ;
  assign n4001 = ~n1288 & ~n3929 ;
  assign n4002 = \pi0299  & n1288 ;
  assign n4003 = n1288 & ~n3771 ;
  assign n4004 = n3770 & n4003 ;
  assign n4005 = ~n4002 & ~n4004 ;
  assign n4006 = \pi0100  & n4005 ;
  assign n4007 = ~n4001 & n4006 ;
  assign n4008 = n3734 & n3748 ;
  assign n4009 = ~n3827 & ~n4008 ;
  assign n4010 = n3829 & n4009 ;
  assign n4011 = n3832 & ~n4001 ;
  assign n4012 = ~n4010 & n4011 ;
  assign n4013 = ~n4007 & ~n4012 ;
  assign n4014 = ~\pi0087  & ~n4013 ;
  assign n4015 = ~n2328 & ~n3929 ;
  assign n4016 = \pi0087  & ~n4015 ;
  assign n4017 = n3925 & n4016 ;
  assign n4018 = ~\pi0075  & ~n4017 ;
  assign n4019 = ~n4014 & n4018 ;
  assign n4020 = ~n4000 & n4019 ;
  assign n4021 = \pi0075  & \pi0299  ;
  assign n4022 = \pi0075  & ~n3771 ;
  assign n4023 = n3770 & n4022 ;
  assign n4024 = ~n4021 & ~n4023 ;
  assign n4025 = ~\pi0092  & n4024 ;
  assign n4026 = n2633 & ~n3992 ;
  assign n4027 = ~n4025 & ~n4026 ;
  assign n4028 = ~n3946 & ~n4027 ;
  assign n4029 = ~n4020 & n4028 ;
  assign n4030 = ~n3947 & ~n4029 ;
  assign n4031 = ~n3752 & n3789 ;
  assign n4032 = \pi0055  & ~n4031 ;
  assign n4033 = ~\pi0056  & ~n4032 ;
  assign n4034 = ~\pi0056  & n3787 ;
  assign n4035 = ~n3922 & n4034 ;
  assign n4036 = ~n4033 & ~n4035 ;
  assign n4037 = ~n3940 & n3943 ;
  assign n4038 = ~n1292 & ~n4037 ;
  assign n4039 = n4036 & ~n4038 ;
  assign n4040 = ~\pi0241  & n2467 ;
  assign n4041 = ~n2504 & ~n3753 ;
  assign n4042 = ~n3752 & n4041 ;
  assign n4043 = \pi0062  & ~n4042 ;
  assign n4044 = ~\pi0056  & ~n3753 ;
  assign n4045 = n2404 & n4044 ;
  assign n4046 = n2403 & n4045 ;
  assign n4047 = ~n3922 & n4046 ;
  assign n4048 = n4043 & ~n4047 ;
  assign n4049 = n4040 & ~n4048 ;
  assign n4050 = ~n4039 & n4049 ;
  assign n4051 = n4030 & n4050 ;
  assign n4052 = ~\pi0055  & ~n3753 ;
  assign n4053 = n1291 & n4052 ;
  assign n4054 = ~n3786 & n4053 ;
  assign n4055 = ~n2407 & n3756 ;
  assign n4056 = ~n3752 & n4055 ;
  assign n4057 = ~\pi0062  & ~n4056 ;
  assign n4058 = ~n4054 & n4057 ;
  assign n4059 = ~n1292 & ~n4058 ;
  assign n4060 = n3912 & n4059 ;
  assign n4061 = \pi0241  & n3755 ;
  assign n4062 = ~n2467 & ~n4061 ;
  assign n4063 = ~n3753 & n4062 ;
  assign n4064 = ~n3752 & n4063 ;
  assign n4065 = ~n4060 & ~n4064 ;
  assign n4066 = ~n4051 & n4065 ;
  assign n4067 = ~n3914 & n4066 ;
  assign n4068 = \pi0216  & \pi0282  ;
  assign n4069 = ~\pi0221  & ~n4068 ;
  assign n4070 = \pi0221  & \pi1140  ;
  assign n4071 = ~n1220 & n4070 ;
  assign n4072 = \pi0221  & \pi0921  ;
  assign n4073 = n1220 & n4072 ;
  assign n4074 = ~n4071 & ~n4073 ;
  assign n4075 = ~n4069 & n4074 ;
  assign n4076 = ~\pi0215  & ~n4075 ;
  assign n4077 = ~\pi0105  & \pi0170  ;
  assign n4078 = \pi0228  & ~n4077 ;
  assign n4079 = ~\pi0216  & ~n4078 ;
  assign n4080 = \pi0869  & ~n1633 ;
  assign n4081 = n3746 & ~n4080 ;
  assign n4082 = ~n4079 & ~n4081 ;
  assign n4083 = ~\pi0170  & ~\pi0228  ;
  assign n4084 = n4074 & ~n4083 ;
  assign n4085 = ~n4082 & n4084 ;
  assign n4086 = n4076 & ~n4085 ;
  assign n4087 = \pi0215  & \pi1140  ;
  assign n4088 = n1295 & ~n4068 ;
  assign n4089 = n2651 & n4088 ;
  assign n4090 = ~n4087 & ~n4089 ;
  assign n4091 = ~n4086 & n4090 ;
  assign n4092 = \pi0299  & ~n4091 ;
  assign n4093 = \pi0222  & \pi1140  ;
  assign n4094 = ~n2192 & n4093 ;
  assign n4095 = \pi0222  & \pi0921  ;
  assign n4096 = n2192 & n4095 ;
  assign n4097 = ~n4094 & ~n4096 ;
  assign n4098 = ~\pi0223  & ~n4097 ;
  assign n4099 = ~\pi0224  & ~n4080 ;
  assign n4100 = \pi0224  & \pi0282  ;
  assign n4101 = ~\pi0222  & ~n4100 ;
  assign n4102 = ~\pi0223  & n4101 ;
  assign n4103 = ~n4099 & n4102 ;
  assign n4104 = ~n4098 & ~n4103 ;
  assign n4105 = \pi0223  & \pi1140  ;
  assign n4106 = ~n3045 & ~n4105 ;
  assign n4107 = n4104 & n4106 ;
  assign n4108 = ~\pi0299  & ~n4107 ;
  assign n4109 = ~n2511 & ~n4108 ;
  assign n4110 = ~n4092 & n4109 ;
  assign n4111 = ~\pi0055  & ~n4110 ;
  assign n4112 = \pi0170  & ~n2280 ;
  assign n4113 = ~\pi0869  & n1281 ;
  assign n4114 = n1260 & n4113 ;
  assign n4115 = ~\pi0228  & ~n4114 ;
  assign n4116 = ~n4112 & n4115 ;
  assign n4117 = ~n2651 & n4074 ;
  assign n4118 = ~n4082 & n4117 ;
  assign n4119 = ~n4116 & n4118 ;
  assign n4120 = n4076 & ~n4119 ;
  assign n4121 = n1291 & ~n4087 ;
  assign n4122 = ~n4120 & n4121 ;
  assign n4123 = ~n1291 & ~n4087 ;
  assign n4124 = ~n4089 & n4123 ;
  assign n4125 = ~n4086 & n4124 ;
  assign n4126 = \pi0055  & ~n4125 ;
  assign n4127 = ~n4122 & n4126 ;
  assign n4128 = ~n4111 & ~n4127 ;
  assign n4129 = n2328 & ~n4108 ;
  assign n4130 = ~\pi0299  & n4129 ;
  assign n4131 = ~n4087 & n4129 ;
  assign n4132 = ~n4120 & n4131 ;
  assign n4133 = ~n4130 & ~n4132 ;
  assign n4134 = ~n2328 & ~n4108 ;
  assign n4135 = ~n4092 & n4134 ;
  assign n4136 = \pi0087  & ~n4135 ;
  assign n4137 = n4133 & n4136 ;
  assign n4138 = ~\pi0075  & ~n4137 ;
  assign n4139 = \pi0075  & ~n4108 ;
  assign n4140 = ~n4092 & n4139 ;
  assign n4141 = ~\pi0092  & ~n4140 ;
  assign n4142 = ~n4138 & n4141 ;
  assign n4143 = \pi0038  & ~n4108 ;
  assign n4144 = ~n4092 & n4143 ;
  assign n4145 = ~\pi0100  & ~n4144 ;
  assign n4146 = ~n1288 & ~n4108 ;
  assign n4147 = ~n4092 & n4146 ;
  assign n4148 = n1288 & ~n4108 ;
  assign n4149 = \pi0100  & ~n4148 ;
  assign n4150 = ~n4147 & n4149 ;
  assign n4151 = ~n2651 & ~n4082 ;
  assign n4152 = n4069 & ~n4151 ;
  assign n4153 = ~\pi0869  & ~n2618 ;
  assign n4154 = ~n2615 & n4153 ;
  assign n4155 = ~\pi0228  & ~n4154 ;
  assign n4156 = \pi0170  & n2618 ;
  assign n4157 = \pi0170  & ~n2609 ;
  assign n4158 = n2614 & n4157 ;
  assign n4159 = ~n4156 & ~n4158 ;
  assign n4160 = n4069 & n4159 ;
  assign n4161 = n4155 & n4160 ;
  assign n4162 = ~n4152 & ~n4161 ;
  assign n4163 = n4074 & ~n4087 ;
  assign n4164 = n4162 & n4163 ;
  assign n4165 = \pi0215  & ~\pi1140  ;
  assign n4166 = n2960 & ~n4165 ;
  assign n4167 = ~n4147 & n4166 ;
  assign n4168 = ~n4164 & n4167 ;
  assign n4169 = ~n4150 & ~n4168 ;
  assign n4170 = ~n4145 & n4169 ;
  assign n4171 = ~\pi0869  & n1640 ;
  assign n4172 = ~n2591 & n4171 ;
  assign n4173 = ~n2704 & n4172 ;
  assign n4174 = ~\pi0170  & ~n4173 ;
  assign n4175 = ~\pi0869  & n2718 ;
  assign n4176 = \pi0170  & ~n4175 ;
  assign n4177 = n3124 & n4176 ;
  assign n4178 = ~n2581 & n4177 ;
  assign n4179 = \pi0170  & ~\pi0869  ;
  assign n4180 = ~n2718 & n4179 ;
  assign n4181 = ~n4178 & ~n4180 ;
  assign n4182 = ~n4174 & n4181 ;
  assign n4183 = n3668 & ~n4068 ;
  assign n4184 = ~n4182 & n4183 ;
  assign n4185 = n3853 & ~n4082 ;
  assign n4186 = n4069 & ~n4185 ;
  assign n4187 = \pi0299  & ~n4087 ;
  assign n4188 = n4074 & n4187 ;
  assign n4189 = ~n4186 & n4188 ;
  assign n4190 = ~n4184 & n4189 ;
  assign n4191 = ~\pi1140  & n2259 ;
  assign n4192 = n4097 & ~n4101 ;
  assign n4193 = n2192 & ~n4095 ;
  assign n4194 = n3503 & ~n4093 ;
  assign n4195 = ~n4193 & ~n4194 ;
  assign n4196 = ~n4080 & ~n4195 ;
  assign n4197 = ~\pi0095  & ~n4195 ;
  assign n4198 = n2686 & n4197 ;
  assign n4199 = ~n4196 & ~n4198 ;
  assign n4200 = ~n4192 & n4199 ;
  assign n4201 = ~\pi0299  & ~n4105 ;
  assign n4202 = n1633 & n4101 ;
  assign n4203 = ~\pi0095  & n4101 ;
  assign n4204 = n2686 & n4203 ;
  assign n4205 = ~n4202 & ~n4204 ;
  assign n4206 = n4201 & n4205 ;
  assign n4207 = ~n4200 & n4206 ;
  assign n4208 = ~\pi1140  & n3498 ;
  assign n4209 = ~\pi0039  & ~n4208 ;
  assign n4210 = ~n4207 & n4209 ;
  assign n4211 = ~n4191 & n4210 ;
  assign n4212 = ~n4190 & n4211 ;
  assign n4213 = ~\pi0038  & ~n4108 ;
  assign n4214 = ~\pi0299  & n4213 ;
  assign n4215 = ~n4087 & n4213 ;
  assign n4216 = ~n4120 & n4215 ;
  assign n4217 = ~n4214 & ~n4216 ;
  assign n4218 = ~n1288 & n4217 ;
  assign n4219 = n4169 & ~n4218 ;
  assign n4220 = ~n4212 & n4219 ;
  assign n4221 = ~n4170 & ~n4220 ;
  assign n4222 = ~\pi0087  & n4141 ;
  assign n4223 = n4221 & n4222 ;
  assign n4224 = ~n4142 & ~n4223 ;
  assign n4225 = ~n1286 & ~n4108 ;
  assign n4226 = ~n4092 & n4225 ;
  assign n4227 = \pi0092  & ~n4226 ;
  assign n4228 = ~n4135 & n4227 ;
  assign n4229 = n4133 & n4228 ;
  assign n4230 = n2387 & ~n4226 ;
  assign n4231 = n2511 & ~n4230 ;
  assign n4232 = ~n4229 & n4231 ;
  assign n4233 = ~n4127 & n4232 ;
  assign n4234 = n4224 & n4233 ;
  assign n4235 = ~n4128 & ~n4234 ;
  assign n4236 = n2504 & ~n4087 ;
  assign n4237 = ~n4120 & n4236 ;
  assign n4238 = ~n2504 & n4090 ;
  assign n4239 = ~n4086 & n4238 ;
  assign n4240 = \pi0062  & ~n4239 ;
  assign n4241 = ~n4237 & n4240 ;
  assign n4242 = \pi0248  & n2467 ;
  assign n4243 = ~n4241 & n4242 ;
  assign n4244 = ~\pi0056  & n4243 ;
  assign n4245 = ~n4235 & n4244 ;
  assign n4246 = n4104 & ~n4105 ;
  assign n4247 = ~\pi0299  & n4246 ;
  assign n4248 = ~n4086 & n4187 ;
  assign n4249 = ~n4247 & ~n4248 ;
  assign n4250 = \pi0092  & n4249 ;
  assign n4251 = ~n3089 & ~n4250 ;
  assign n4252 = n2387 & n4249 ;
  assign n4253 = n2511 & ~n4252 ;
  assign n4254 = n4251 & n4253 ;
  assign n4255 = \pi0299  & n4087 ;
  assign n4256 = n4074 & ~n4082 ;
  assign n4257 = ~n4116 & n4256 ;
  assign n4258 = ~n4075 & ~n4257 ;
  assign n4259 = n2256 & n4258 ;
  assign n4260 = ~n4255 & ~n4259 ;
  assign n4261 = n2328 & ~n4105 ;
  assign n4262 = n4104 & n4261 ;
  assign n4263 = ~n3915 & ~n4262 ;
  assign n4264 = n4253 & ~n4263 ;
  assign n4265 = n4260 & n4264 ;
  assign n4266 = ~n4254 & ~n4265 ;
  assign n4267 = ~n2511 & ~n4249 ;
  assign n4268 = ~\pi0055  & ~n4267 ;
  assign n4269 = n1292 & n4268 ;
  assign n4270 = ~\pi0215  & n4258 ;
  assign n4271 = n2407 & ~n4087 ;
  assign n4272 = ~n4270 & n4271 ;
  assign n4273 = ~n2407 & ~n4087 ;
  assign n4274 = ~n4086 & n4273 ;
  assign n4275 = ~\pi0062  & ~n4274 ;
  assign n4276 = n4268 & n4275 ;
  assign n4277 = ~n4272 & n4276 ;
  assign n4278 = ~n4269 & ~n4277 ;
  assign n4279 = n4266 & ~n4278 ;
  assign n4280 = \pi0105  & ~n4080 ;
  assign n4281 = n4078 & ~n4280 ;
  assign n4282 = ~n1633 & n4281 ;
  assign n4283 = ~n2716 & n4282 ;
  assign n4284 = n2225 & ~n4077 ;
  assign n4285 = ~\pi0216  & ~n4284 ;
  assign n4286 = ~n4283 & n4285 ;
  assign n4287 = \pi0170  & n1640 ;
  assign n4288 = ~n2591 & n4287 ;
  assign n4289 = ~n2704 & n4288 ;
  assign n4290 = \pi0869  & n4289 ;
  assign n4291 = ~\pi0228  & n4290 ;
  assign n4292 = ~n2716 & n4080 ;
  assign n4293 = ~n1639 & ~n4292 ;
  assign n4294 = ~\pi0869  & n2591 ;
  assign n4295 = ~\pi0869  & ~n2580 ;
  assign n4296 = n2574 & n4295 ;
  assign n4297 = ~n4294 & ~n4296 ;
  assign n4298 = n4293 & n4297 ;
  assign n4299 = n4083 & ~n4298 ;
  assign n4300 = ~n4291 & ~n4299 ;
  assign n4301 = n4286 & n4300 ;
  assign n4302 = ~\pi0215  & n4069 ;
  assign n4303 = ~n4301 & n4302 ;
  assign n4304 = ~\pi0038  & ~n4105 ;
  assign n4305 = n4104 & n4304 ;
  assign n4306 = ~n3972 & ~n4305 ;
  assign n4307 = n4260 & ~n4306 ;
  assign n4308 = ~n1288 & ~n4307 ;
  assign n4309 = ~\pi0215  & ~n4074 ;
  assign n4310 = n4187 & ~n4309 ;
  assign n4311 = ~n4308 & n4310 ;
  assign n4312 = ~n4303 & n4311 ;
  assign n4313 = ~n4200 & n4201 ;
  assign n4314 = n4210 & ~n4313 ;
  assign n4315 = \pi0038  & ~n4105 ;
  assign n4316 = n4104 & n4315 ;
  assign n4317 = ~n3987 & ~n4316 ;
  assign n4318 = ~\pi0100  & n4317 ;
  assign n4319 = ~n4086 & ~n4087 ;
  assign n4320 = n2563 & ~n4319 ;
  assign n4321 = ~n4318 & ~n4320 ;
  assign n4322 = ~\pi0087  & ~n4321 ;
  assign n4323 = n4314 & n4322 ;
  assign n4324 = ~n1288 & n4322 ;
  assign n4325 = ~n4307 & n4324 ;
  assign n4326 = ~n4323 & ~n4325 ;
  assign n4327 = ~n4312 & ~n4326 ;
  assign n4328 = ~n1288 & ~n4249 ;
  assign n4329 = n1288 & ~n4105 ;
  assign n4330 = n4104 & n4329 ;
  assign n4331 = ~n4002 & ~n4330 ;
  assign n4332 = \pi0100  & n4331 ;
  assign n4333 = ~n4328 & n4332 ;
  assign n4334 = n4069 & n4082 ;
  assign n4335 = ~n4161 & ~n4334 ;
  assign n4336 = n4163 & n4335 ;
  assign n4337 = n4166 & ~n4328 ;
  assign n4338 = ~n4336 & n4337 ;
  assign n4339 = ~n4333 & ~n4338 ;
  assign n4340 = ~\pi0087  & ~n4339 ;
  assign n4341 = ~n2328 & ~n4249 ;
  assign n4342 = \pi0087  & ~n4341 ;
  assign n4343 = ~\pi0075  & ~n4342 ;
  assign n4344 = ~\pi0075  & ~n4263 ;
  assign n4345 = n4260 & n4344 ;
  assign n4346 = ~n4343 & ~n4345 ;
  assign n4347 = ~n4340 & ~n4346 ;
  assign n4348 = ~n4327 & n4347 ;
  assign n4349 = \pi0075  & ~n4105 ;
  assign n4350 = n4104 & n4349 ;
  assign n4351 = ~n4021 & ~n4350 ;
  assign n4352 = ~\pi0092  & n4351 ;
  assign n4353 = n2633 & ~n4319 ;
  assign n4354 = ~n4352 & ~n4353 ;
  assign n4355 = ~n4278 & ~n4354 ;
  assign n4356 = ~n4348 & n4355 ;
  assign n4357 = ~n4279 & ~n4356 ;
  assign n4358 = ~n4086 & n4123 ;
  assign n4359 = \pi0055  & ~n4358 ;
  assign n4360 = ~n4121 & n4359 ;
  assign n4361 = ~\pi0215  & n4359 ;
  assign n4362 = n4258 & n4361 ;
  assign n4363 = ~n4360 & ~n4362 ;
  assign n4364 = ~\pi0056  & n4363 ;
  assign n4365 = ~n4272 & n4275 ;
  assign n4366 = ~n1292 & ~n4365 ;
  assign n4367 = ~n4364 & ~n4366 ;
  assign n4368 = ~\pi0248  & n2467 ;
  assign n4369 = ~n2504 & ~n4087 ;
  assign n4370 = ~n4086 & n4369 ;
  assign n4371 = \pi0062  & ~n4370 ;
  assign n4372 = ~\pi0056  & ~n4087 ;
  assign n4373 = n2404 & n4372 ;
  assign n4374 = n2403 & n4373 ;
  assign n4375 = n4371 & ~n4374 ;
  assign n4376 = ~\pi0215  & n4371 ;
  assign n4377 = n4258 & n4376 ;
  assign n4378 = ~n4375 & ~n4377 ;
  assign n4379 = n4368 & n4378 ;
  assign n4380 = ~n4367 & n4379 ;
  assign n4381 = n4357 & n4380 ;
  assign n4382 = ~\pi0055  & ~n4087 ;
  assign n4383 = n1291 & n4382 ;
  assign n4384 = ~n4120 & n4383 ;
  assign n4385 = ~n2407 & n4090 ;
  assign n4386 = ~n4086 & n4385 ;
  assign n4387 = ~\pi0062  & ~n4386 ;
  assign n4388 = ~n4384 & n4387 ;
  assign n4389 = ~n1292 & ~n4388 ;
  assign n4390 = n4243 & n4389 ;
  assign n4391 = \pi0248  & n4089 ;
  assign n4392 = ~n2467 & ~n4391 ;
  assign n4393 = ~n4087 & n4392 ;
  assign n4394 = ~n4086 & n4393 ;
  assign n4395 = ~n4390 & ~n4394 ;
  assign n4396 = ~n4381 & n4395 ;
  assign n4397 = ~n4245 & n4396 ;
  assign n4398 = \pi0148  & ~n1209 ;
  assign n4399 = ~\pi0215  & ~n4398 ;
  assign n4400 = \pi0833  & \pi0920  ;
  assign n4401 = ~\pi0833  & \pi1139  ;
  assign n4402 = ~\pi0216  & ~n4401 ;
  assign n4403 = ~n4400 & n4402 ;
  assign n4404 = ~\pi0215  & ~n2352 ;
  assign n4405 = ~n4403 & n4404 ;
  assign n4406 = ~n4399 & ~n4405 ;
  assign n4407 = \pi0216  & ~\pi1139  ;
  assign n4408 = \pi0221  & ~n4407 ;
  assign n4409 = ~n4403 & n4408 ;
  assign n4410 = \pi0216  & \pi0281  ;
  assign n4411 = ~\pi0221  & ~n4410 ;
  assign n4412 = ~\pi0216  & ~\pi0862  ;
  assign n4413 = n2721 & n4412 ;
  assign n4414 = n4411 & ~n4413 ;
  assign n4415 = ~n4409 & ~n4414 ;
  assign n4416 = ~n4406 & ~n4415 ;
  assign n4417 = \pi0215  & \pi1139  ;
  assign n4418 = ~n2467 & ~n4417 ;
  assign n4419 = ~n4416 & n4418 ;
  assign n4420 = \pi0247  & ~n4419 ;
  assign n4421 = ~n2721 & n4411 ;
  assign n4422 = ~n3421 & n4421 ;
  assign n4423 = n4411 & ~n4412 ;
  assign n4424 = ~n4409 & ~n4423 ;
  assign n4425 = ~n4422 & n4424 ;
  assign n4426 = \pi0148  & ~\pi0215  ;
  assign n4427 = ~n2352 & ~n4403 ;
  assign n4428 = ~n2721 & ~n4427 ;
  assign n4429 = ~n3421 & n4428 ;
  assign n4430 = n4426 & ~n4429 ;
  assign n4431 = ~n4425 & n4430 ;
  assign n4432 = ~n4406 & ~n4424 ;
  assign n4433 = ~n4406 & n4421 ;
  assign n4434 = ~n3421 & n4433 ;
  assign n4435 = ~n4432 & ~n4434 ;
  assign n4436 = n2454 & ~n4417 ;
  assign n4437 = n4435 & n4436 ;
  assign n4438 = ~n4431 & n4437 ;
  assign n4439 = ~n2504 & ~n4417 ;
  assign n4440 = ~n4416 & n4439 ;
  assign n4441 = \pi0062  & ~n4440 ;
  assign n4442 = ~n4438 & n4441 ;
  assign n4443 = n2467 & ~n4442 ;
  assign n4444 = ~n4416 & ~n4417 ;
  assign n4445 = \pi0299  & ~n4444 ;
  assign n4446 = \pi0223  & ~\pi1139  ;
  assign n4447 = \pi0222  & \pi1139  ;
  assign n4448 = ~n2192 & n4447 ;
  assign n4449 = \pi0222  & \pi0920  ;
  assign n4450 = n2192 & n4449 ;
  assign n4451 = ~n4448 & ~n4450 ;
  assign n4452 = \pi0223  & \pi1139  ;
  assign n4453 = \pi0224  & \pi0281  ;
  assign n4454 = ~\pi0222  & ~n4453 ;
  assign n4455 = ~n4452 & ~n4454 ;
  assign n4456 = n4451 & n4455 ;
  assign n4457 = ~n4446 & ~n4456 ;
  assign n4458 = ~\pi0224  & ~n4452 ;
  assign n4459 = ~\pi0862  & n4458 ;
  assign n4460 = n4451 & n4459 ;
  assign n4461 = ~\pi0299  & ~n4460 ;
  assign n4462 = n4457 & n4461 ;
  assign n4463 = ~n2666 & ~n4462 ;
  assign n4464 = \pi0075  & n4463 ;
  assign n4465 = ~n4445 & n4464 ;
  assign n4466 = ~n1288 & n4463 ;
  assign n4467 = ~n4445 & n4466 ;
  assign n4468 = n2952 & ~n4462 ;
  assign n4469 = \pi0100  & ~n4468 ;
  assign n4470 = ~n4467 & n4469 ;
  assign n4471 = ~\pi0148  & ~\pi0215  ;
  assign n4472 = ~n4425 & n4471 ;
  assign n4473 = n4421 & n4471 ;
  assign n4474 = ~n2943 & n4473 ;
  assign n4475 = ~n4472 & ~n4474 ;
  assign n4476 = ~n1209 & ~n4400 ;
  assign n4477 = n4402 & n4476 ;
  assign n4478 = ~n2477 & ~n4477 ;
  assign n4479 = ~n2943 & ~n4478 ;
  assign n4480 = ~n4425 & n4426 ;
  assign n4481 = ~n4479 & n4480 ;
  assign n4482 = ~n4417 & ~n4481 ;
  assign n4483 = n4475 & n4482 ;
  assign n4484 = n2960 & ~n4467 ;
  assign n4485 = ~n4483 & n4484 ;
  assign n4486 = ~n4470 & ~n4485 ;
  assign n4487 = ~n4465 & ~n4486 ;
  assign n4488 = n4408 & n4426 ;
  assign n4489 = ~n4403 & n4488 ;
  assign n4490 = ~\pi0228  & ~n1639 ;
  assign n4491 = ~n2591 & n4490 ;
  assign n4492 = ~n2581 & n4491 ;
  assign n4493 = ~\pi0862  & ~n2713 ;
  assign n4494 = ~n2915 & n4493 ;
  assign n4495 = ~\pi0216  & ~n4494 ;
  assign n4496 = ~n1209 & n4495 ;
  assign n4497 = ~n4492 & n4496 ;
  assign n4498 = ~n2713 & ~n2915 ;
  assign n4499 = n4412 & ~n4498 ;
  assign n4500 = n4411 & n4426 ;
  assign n4501 = ~n4499 & n4500 ;
  assign n4502 = ~n4497 & n4501 ;
  assign n4503 = ~n4489 & ~n4502 ;
  assign n4504 = ~n4417 & ~n4471 ;
  assign n4505 = ~\pi0095  & n4411 ;
  assign n4506 = n2686 & n4505 ;
  assign n4507 = ~n4421 & ~n4506 ;
  assign n4508 = ~n2708 & ~n4507 ;
  assign n4509 = ~n4417 & n4424 ;
  assign n4510 = ~n4508 & n4509 ;
  assign n4511 = ~n4504 & ~n4510 ;
  assign n4512 = n4503 & ~n4511 ;
  assign n4513 = n2738 & ~n4512 ;
  assign n4514 = ~\pi0299  & ~n4446 ;
  assign n4515 = ~n4456 & n4514 ;
  assign n4516 = ~\pi0862  & ~n1633 ;
  assign n4517 = n4458 & n4516 ;
  assign n4518 = n4451 & n4517 ;
  assign n4519 = ~\pi0039  & ~n4518 ;
  assign n4520 = ~\pi0039  & ~\pi0095  ;
  assign n4521 = n2686 & n4520 ;
  assign n4522 = ~n4519 & ~n4521 ;
  assign n4523 = n4515 & ~n4522 ;
  assign n4524 = \pi0039  & ~n4463 ;
  assign n4525 = ~n4417 & n4435 ;
  assign n4526 = ~n4431 & n4525 ;
  assign n4527 = n2297 & ~n4526 ;
  assign n4528 = ~n4524 & ~n4527 ;
  assign n4529 = ~\pi0038  & n4528 ;
  assign n4530 = ~n4523 & n4529 ;
  assign n4531 = ~n4513 & n4530 ;
  assign n4532 = n2973 & ~n4462 ;
  assign n4533 = ~\pi0100  & ~n4532 ;
  assign n4534 = n2563 & ~n4444 ;
  assign n4535 = ~n4533 & ~n4534 ;
  assign n4536 = ~n4465 & ~n4535 ;
  assign n4537 = ~n4531 & n4536 ;
  assign n4538 = ~n4487 & ~n4537 ;
  assign n4539 = ~\pi0087  & ~\pi0092  ;
  assign n4540 = ~n4538 & n4539 ;
  assign n4541 = \pi0299  & ~n4526 ;
  assign n4542 = n2328 & n4463 ;
  assign n4543 = ~n4541 & n4542 ;
  assign n4544 = ~n2328 & n4463 ;
  assign n4545 = ~n4445 & n4544 ;
  assign n4546 = \pi0087  & ~n4545 ;
  assign n4547 = ~n4543 & n4546 ;
  assign n4548 = ~\pi0075  & ~n4547 ;
  assign n4549 = n2753 & ~n4462 ;
  assign n4550 = ~\pi0092  & ~n4549 ;
  assign n4551 = n2633 & ~n4444 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = ~n4548 & ~n4552 ;
  assign n4554 = ~n1286 & n4463 ;
  assign n4555 = ~n4445 & n4554 ;
  assign n4556 = \pi0092  & ~n4555 ;
  assign n4557 = ~n1286 & n4556 ;
  assign n4558 = ~n4545 & n4556 ;
  assign n4559 = ~n4543 & n4558 ;
  assign n4560 = ~n4557 & ~n4559 ;
  assign n4561 = n1291 & ~n4417 ;
  assign n4562 = n4435 & n4561 ;
  assign n4563 = ~n4431 & n4562 ;
  assign n4564 = ~n1291 & ~n4417 ;
  assign n4565 = ~n4416 & n4564 ;
  assign n4566 = \pi0055  & ~n4565 ;
  assign n4567 = ~n4563 & n4566 ;
  assign n4568 = ~\pi0056  & ~n4567 ;
  assign n4569 = n2511 & n4568 ;
  assign n4570 = n4560 & n4569 ;
  assign n4571 = ~n4553 & n4570 ;
  assign n4572 = ~n4540 & n4571 ;
  assign n4573 = ~n2511 & n4463 ;
  assign n4574 = ~n4445 & n4573 ;
  assign n4575 = ~\pi0055  & ~n4574 ;
  assign n4576 = ~\pi0056  & ~n4575 ;
  assign n4577 = ~n4567 & n4576 ;
  assign n4578 = n2407 & ~n4417 ;
  assign n4579 = n4435 & n4578 ;
  assign n4580 = ~n4431 & n4579 ;
  assign n4581 = ~n2407 & ~n4417 ;
  assign n4582 = ~n4416 & n4581 ;
  assign n4583 = ~\pi0062  & ~n4582 ;
  assign n4584 = ~n4580 & n4583 ;
  assign n4585 = ~n1292 & ~n4584 ;
  assign n4586 = ~n4577 & ~n4585 ;
  assign n4587 = ~n4572 & n4586 ;
  assign n4588 = n4443 & ~n4587 ;
  assign n4589 = n4420 & ~n4588 ;
  assign n4590 = \pi0862  & ~n2651 ;
  assign n4591 = ~\pi0216  & ~n4590 ;
  assign n4592 = n4411 & ~n4591 ;
  assign n4593 = ~n4409 & ~n4592 ;
  assign n4594 = n4471 & ~n4593 ;
  assign n4595 = ~n1209 & n4411 ;
  assign n4596 = n4471 & n4595 ;
  assign n4597 = ~n3421 & n4596 ;
  assign n4598 = ~n4594 & ~n4597 ;
  assign n4599 = n4436 & n4598 ;
  assign n4600 = ~n4431 & n4599 ;
  assign n4601 = n4398 & ~n4427 ;
  assign n4602 = ~n4415 & ~n4601 ;
  assign n4603 = n3409 & n4602 ;
  assign n4604 = n4439 & ~n4603 ;
  assign n4605 = \pi0062  & ~n4604 ;
  assign n4606 = ~n4600 & n4605 ;
  assign n4607 = n2467 & ~n4606 ;
  assign n4608 = n4578 & n4598 ;
  assign n4609 = ~n4431 & n4608 ;
  assign n4610 = n4581 & ~n4603 ;
  assign n4611 = ~\pi0062  & ~n4610 ;
  assign n4612 = ~n4609 & n4611 ;
  assign n4613 = ~n1292 & ~n4612 ;
  assign n4614 = n4607 & n4613 ;
  assign n4615 = \pi0299  & n4417 ;
  assign n4616 = \pi0299  & n3409 ;
  assign n4617 = n4602 & n4616 ;
  assign n4618 = ~n4615 & ~n4617 ;
  assign n4619 = n1633 & n4458 ;
  assign n4620 = n4451 & n4619 ;
  assign n4621 = n4461 & ~n4620 ;
  assign n4622 = n4457 & n4621 ;
  assign n4623 = ~n2511 & ~n4622 ;
  assign n4624 = n4618 & n4623 ;
  assign n4625 = ~\pi0055  & ~n4624 ;
  assign n4626 = ~n4417 & n4598 ;
  assign n4627 = ~n4431 & n4626 ;
  assign n4628 = \pi0299  & ~n4627 ;
  assign n4629 = n1286 & n2328 ;
  assign n4630 = ~n4622 & n4629 ;
  assign n4631 = ~n4628 & n4630 ;
  assign n4632 = n1286 & ~n2328 ;
  assign n4633 = ~n4622 & n4632 ;
  assign n4634 = n4618 & n4633 ;
  assign n4635 = ~n1286 & ~n4622 ;
  assign n4636 = n4618 & n4635 ;
  assign n4637 = \pi0092  & ~n4636 ;
  assign n4638 = ~n4634 & n4637 ;
  assign n4639 = ~n4631 & n4638 ;
  assign n4640 = n2511 & ~n4639 ;
  assign n4641 = n4625 & ~n4640 ;
  assign n4642 = n2328 & ~n4622 ;
  assign n4643 = ~n4628 & n4642 ;
  assign n4644 = ~n2328 & ~n4622 ;
  assign n4645 = n4618 & n4644 ;
  assign n4646 = \pi0087  & ~n4645 ;
  assign n4647 = ~n4643 & n4646 ;
  assign n4648 = ~\pi0075  & ~n4647 ;
  assign n4649 = \pi0087  & n4648 ;
  assign n4650 = \pi0038  & ~n4622 ;
  assign n4651 = n4618 & n4650 ;
  assign n4652 = ~\pi0100  & ~n4651 ;
  assign n4653 = \pi0039  & n4622 ;
  assign n4654 = n2297 & ~n4627 ;
  assign n4655 = ~n4653 & ~n4654 ;
  assign n4656 = ~\pi0038  & n4655 ;
  assign n4657 = n4652 & ~n4656 ;
  assign n4658 = ~n4409 & ~n4411 ;
  assign n4659 = \pi0862  & n2713 ;
  assign n4660 = ~\pi0216  & ~n4659 ;
  assign n4661 = ~\pi0228  & \pi0862  ;
  assign n4662 = n2718 & n4661 ;
  assign n4663 = ~n4409 & ~n4662 ;
  assign n4664 = n4660 & n4663 ;
  assign n4665 = ~n4658 & ~n4664 ;
  assign n4666 = ~\pi0862  & ~n1209 ;
  assign n4667 = ~n4658 & n4666 ;
  assign n4668 = ~n4492 & n4667 ;
  assign n4669 = ~n4665 & ~n4668 ;
  assign n4670 = n4471 & ~n4669 ;
  assign n4671 = \pi0299  & ~n4417 ;
  assign n4672 = ~n4426 & n4671 ;
  assign n4673 = ~\pi0095  & ~n4427 ;
  assign n4674 = n2686 & n4673 ;
  assign n4675 = ~n4428 & ~n4674 ;
  assign n4676 = n4671 & ~n4675 ;
  assign n4677 = ~n2708 & n4676 ;
  assign n4678 = ~n4672 & ~n4677 ;
  assign n4679 = n4424 & n4671 ;
  assign n4680 = ~n4508 & n4679 ;
  assign n4681 = n4678 & ~n4680 ;
  assign n4682 = ~n4670 & ~n4681 ;
  assign n4683 = n4457 & ~n4460 ;
  assign n4684 = ~n1633 & n4683 ;
  assign n4685 = ~n2716 & n4684 ;
  assign n4686 = n4451 & n4458 ;
  assign n4687 = n4457 & ~n4686 ;
  assign n4688 = ~\pi0299  & ~n4687 ;
  assign n4689 = ~n4685 & n4688 ;
  assign n4690 = ~\pi0039  & ~n4689 ;
  assign n4691 = n4652 & n4690 ;
  assign n4692 = ~n4682 & n4691 ;
  assign n4693 = ~n4657 & ~n4692 ;
  assign n4694 = ~n1288 & ~n4622 ;
  assign n4695 = n4618 & n4694 ;
  assign n4696 = n1288 & ~n4622 ;
  assign n4697 = \pi0100  & ~n4696 ;
  assign n4698 = ~n4695 & n4697 ;
  assign n4699 = ~n2943 & n4421 ;
  assign n4700 = n4425 & ~n4699 ;
  assign n4701 = ~n2943 & n4428 ;
  assign n4702 = n4426 & ~n4701 ;
  assign n4703 = ~n4700 & n4702 ;
  assign n4704 = ~n2943 & n4595 ;
  assign n4705 = ~n3421 & n4595 ;
  assign n4706 = n4593 & ~n4705 ;
  assign n4707 = ~n4417 & n4706 ;
  assign n4708 = ~n4704 & n4707 ;
  assign n4709 = ~n4504 & ~n4708 ;
  assign n4710 = ~n4703 & ~n4709 ;
  assign n4711 = n2960 & ~n4695 ;
  assign n4712 = ~n4710 & n4711 ;
  assign n4713 = ~n4698 & ~n4712 ;
  assign n4714 = n4648 & n4713 ;
  assign n4715 = n4693 & n4714 ;
  assign n4716 = ~n4649 & ~n4715 ;
  assign n4717 = \pi0075  & ~n4622 ;
  assign n4718 = n4618 & n4717 ;
  assign n4719 = ~\pi0092  & ~n4718 ;
  assign n4720 = n4625 & n4719 ;
  assign n4721 = n4716 & n4720 ;
  assign n4722 = ~n4641 & ~n4721 ;
  assign n4723 = n4561 & n4598 ;
  assign n4724 = ~n4431 & n4723 ;
  assign n4725 = n4564 & ~n4603 ;
  assign n4726 = \pi0055  & ~n4725 ;
  assign n4727 = ~n4724 & n4726 ;
  assign n4728 = ~\pi0056  & ~n4727 ;
  assign n4729 = n4607 & n4728 ;
  assign n4730 = n4722 & n4729 ;
  assign n4731 = ~n4614 & ~n4730 ;
  assign n4732 = n4418 & ~n4603 ;
  assign n4733 = ~\pi0247  & ~n4732 ;
  assign n4734 = n4731 & n4733 ;
  assign n4735 = ~n4589 & ~n4734 ;
  assign n4736 = \pi0216  & \pi0269  ;
  assign n4737 = ~\pi0221  & ~n4736 ;
  assign n4738 = \pi0221  & \pi1138  ;
  assign n4739 = ~n1220 & n4738 ;
  assign n4740 = \pi0221  & \pi0940  ;
  assign n4741 = n1220 & n4740 ;
  assign n4742 = ~n4739 & ~n4741 ;
  assign n4743 = ~n4737 & n4742 ;
  assign n4744 = ~\pi0215  & ~n4743 ;
  assign n4745 = ~\pi0105  & \pi0169  ;
  assign n4746 = \pi0228  & ~n4745 ;
  assign n4747 = ~\pi0216  & ~n4746 ;
  assign n4748 = \pi0877  & ~n1633 ;
  assign n4749 = n3746 & ~n4748 ;
  assign n4750 = ~n4747 & ~n4749 ;
  assign n4751 = ~\pi0169  & ~\pi0228  ;
  assign n4752 = n4742 & ~n4751 ;
  assign n4753 = ~n4750 & n4752 ;
  assign n4754 = n4744 & ~n4753 ;
  assign n4755 = \pi0215  & \pi1138  ;
  assign n4756 = n1295 & ~n4736 ;
  assign n4757 = n2651 & n4756 ;
  assign n4758 = ~n4755 & ~n4757 ;
  assign n4759 = ~n4754 & n4758 ;
  assign n4760 = \pi0299  & ~n4759 ;
  assign n4761 = \pi0222  & \pi1138  ;
  assign n4762 = ~n2192 & n4761 ;
  assign n4763 = \pi0222  & \pi0940  ;
  assign n4764 = n2192 & n4763 ;
  assign n4765 = ~n4762 & ~n4764 ;
  assign n4766 = ~\pi0223  & ~n4765 ;
  assign n4767 = ~\pi0224  & ~n4748 ;
  assign n4768 = \pi0224  & \pi0269  ;
  assign n4769 = ~\pi0222  & ~n4768 ;
  assign n4770 = ~\pi0223  & n4769 ;
  assign n4771 = ~n4767 & n4770 ;
  assign n4772 = ~n4766 & ~n4771 ;
  assign n4773 = \pi0223  & \pi1138  ;
  assign n4774 = ~n3045 & ~n4773 ;
  assign n4775 = n4772 & n4774 ;
  assign n4776 = ~\pi0299  & ~n4775 ;
  assign n4777 = ~n2511 & ~n4776 ;
  assign n4778 = ~n4760 & n4777 ;
  assign n4779 = ~\pi0055  & ~n4778 ;
  assign n4780 = \pi0169  & ~n2280 ;
  assign n4781 = ~\pi0877  & n1281 ;
  assign n4782 = n1260 & n4781 ;
  assign n4783 = ~\pi0228  & ~n4782 ;
  assign n4784 = ~n4780 & n4783 ;
  assign n4785 = ~n2651 & n4742 ;
  assign n4786 = ~n4750 & n4785 ;
  assign n4787 = ~n4784 & n4786 ;
  assign n4788 = n4744 & ~n4787 ;
  assign n4789 = n1291 & ~n4755 ;
  assign n4790 = ~n4788 & n4789 ;
  assign n4791 = ~n1291 & ~n4755 ;
  assign n4792 = ~n4757 & n4791 ;
  assign n4793 = ~n4754 & n4792 ;
  assign n4794 = \pi0055  & ~n4793 ;
  assign n4795 = ~n4790 & n4794 ;
  assign n4796 = ~n4779 & ~n4795 ;
  assign n4797 = n2328 & ~n4776 ;
  assign n4798 = ~\pi0299  & n4797 ;
  assign n4799 = ~n4755 & n4797 ;
  assign n4800 = ~n4788 & n4799 ;
  assign n4801 = ~n4798 & ~n4800 ;
  assign n4802 = ~n2328 & ~n4776 ;
  assign n4803 = ~n4760 & n4802 ;
  assign n4804 = \pi0087  & ~n4803 ;
  assign n4805 = n4801 & n4804 ;
  assign n4806 = ~\pi0075  & ~n4805 ;
  assign n4807 = \pi0075  & ~n4776 ;
  assign n4808 = ~n4760 & n4807 ;
  assign n4809 = ~\pi0092  & ~n4808 ;
  assign n4810 = ~n4806 & n4809 ;
  assign n4811 = \pi0038  & ~n4776 ;
  assign n4812 = ~n4760 & n4811 ;
  assign n4813 = ~\pi0100  & ~n4812 ;
  assign n4814 = ~n1288 & ~n4776 ;
  assign n4815 = ~n4760 & n4814 ;
  assign n4816 = n1288 & ~n4776 ;
  assign n4817 = \pi0100  & ~n4816 ;
  assign n4818 = ~n4815 & n4817 ;
  assign n4819 = ~n2651 & ~n4750 ;
  assign n4820 = n4737 & ~n4819 ;
  assign n4821 = ~\pi0877  & ~n2618 ;
  assign n4822 = ~n2615 & n4821 ;
  assign n4823 = ~\pi0228  & ~n4822 ;
  assign n4824 = \pi0169  & n2618 ;
  assign n4825 = \pi0169  & ~n2609 ;
  assign n4826 = n2614 & n4825 ;
  assign n4827 = ~n4824 & ~n4826 ;
  assign n4828 = n4737 & n4827 ;
  assign n4829 = n4823 & n4828 ;
  assign n4830 = ~n4820 & ~n4829 ;
  assign n4831 = n4742 & ~n4755 ;
  assign n4832 = n4830 & n4831 ;
  assign n4833 = \pi0215  & ~\pi1138  ;
  assign n4834 = n2960 & ~n4833 ;
  assign n4835 = ~n4815 & n4834 ;
  assign n4836 = ~n4832 & n4835 ;
  assign n4837 = ~n4818 & ~n4836 ;
  assign n4838 = ~n4813 & n4837 ;
  assign n4839 = ~\pi0877  & ~n1633 ;
  assign n4840 = ~n1639 & n4839 ;
  assign n4841 = ~n2591 & n4840 ;
  assign n4842 = ~n2704 & n4841 ;
  assign n4843 = ~\pi0169  & ~n4842 ;
  assign n4844 = n3668 & ~n4736 ;
  assign n4845 = n4843 & n4844 ;
  assign n4846 = \pi0877  & ~n3125 ;
  assign n4847 = ~\pi0877  & n2718 ;
  assign n4848 = \pi0169  & ~n4847 ;
  assign n4849 = n4844 & n4848 ;
  assign n4850 = ~n4846 & n4849 ;
  assign n4851 = ~n4845 & ~n4850 ;
  assign n4852 = n3853 & ~n4750 ;
  assign n4853 = n4737 & ~n4852 ;
  assign n4854 = \pi0299  & ~n4755 ;
  assign n4855 = n4742 & n4854 ;
  assign n4856 = ~n4853 & n4855 ;
  assign n4857 = n4851 & n4856 ;
  assign n4858 = ~\pi1138  & n2259 ;
  assign n4859 = n4765 & ~n4769 ;
  assign n4860 = n2192 & ~n4763 ;
  assign n4861 = n3503 & ~n4761 ;
  assign n4862 = ~n4860 & ~n4861 ;
  assign n4863 = ~n4748 & ~n4862 ;
  assign n4864 = ~\pi0095  & ~n4862 ;
  assign n4865 = n2686 & n4864 ;
  assign n4866 = ~n4863 & ~n4865 ;
  assign n4867 = ~n4859 & n4866 ;
  assign n4868 = ~\pi0299  & ~n4773 ;
  assign n4869 = n1633 & n4769 ;
  assign n4870 = ~\pi0095  & n4769 ;
  assign n4871 = n2686 & n4870 ;
  assign n4872 = ~n4869 & ~n4871 ;
  assign n4873 = n4868 & n4872 ;
  assign n4874 = ~n4867 & n4873 ;
  assign n4875 = ~\pi1138  & n3498 ;
  assign n4876 = ~\pi0039  & ~n4875 ;
  assign n4877 = ~n4874 & n4876 ;
  assign n4878 = ~n4858 & n4877 ;
  assign n4879 = ~n4857 & n4878 ;
  assign n4880 = ~\pi0038  & ~n4776 ;
  assign n4881 = ~\pi0299  & n4880 ;
  assign n4882 = ~n4755 & n4880 ;
  assign n4883 = ~n4788 & n4882 ;
  assign n4884 = ~n4881 & ~n4883 ;
  assign n4885 = ~n1288 & n4884 ;
  assign n4886 = n4837 & ~n4885 ;
  assign n4887 = ~n4879 & n4886 ;
  assign n4888 = ~n4838 & ~n4887 ;
  assign n4889 = ~\pi0087  & n4809 ;
  assign n4890 = n4888 & n4889 ;
  assign n4891 = ~n4810 & ~n4890 ;
  assign n4892 = ~n1286 & ~n4776 ;
  assign n4893 = ~n4760 & n4892 ;
  assign n4894 = \pi0092  & ~n4893 ;
  assign n4895 = ~n4803 & n4894 ;
  assign n4896 = n4801 & n4895 ;
  assign n4897 = n2387 & ~n4893 ;
  assign n4898 = n2511 & ~n4897 ;
  assign n4899 = ~n4896 & n4898 ;
  assign n4900 = ~n4795 & n4899 ;
  assign n4901 = n4891 & n4900 ;
  assign n4902 = ~n4796 & ~n4901 ;
  assign n4903 = n2504 & ~n4755 ;
  assign n4904 = ~n4788 & n4903 ;
  assign n4905 = ~n2504 & n4758 ;
  assign n4906 = ~n4754 & n4905 ;
  assign n4907 = \pi0062  & ~n4906 ;
  assign n4908 = ~n4904 & n4907 ;
  assign n4909 = \pi0246  & n2467 ;
  assign n4910 = ~n4908 & n4909 ;
  assign n4911 = ~\pi0056  & n4910 ;
  assign n4912 = ~n4902 & n4911 ;
  assign n4913 = n2328 & ~n4773 ;
  assign n4914 = n4772 & n4913 ;
  assign n4915 = ~n3915 & ~n4914 ;
  assign n4916 = ~\pi0299  & ~n4915 ;
  assign n4917 = n4742 & ~n4750 ;
  assign n4918 = ~n4784 & n4917 ;
  assign n4919 = n4744 & ~n4918 ;
  assign n4920 = ~n4755 & ~n4915 ;
  assign n4921 = ~n4919 & n4920 ;
  assign n4922 = ~n4916 & ~n4921 ;
  assign n4923 = n4772 & ~n4773 ;
  assign n4924 = ~\pi0299  & n4923 ;
  assign n4925 = ~n4754 & n4854 ;
  assign n4926 = ~n4924 & ~n4925 ;
  assign n4927 = \pi0092  & n4926 ;
  assign n4928 = ~n3089 & ~n4927 ;
  assign n4929 = n4922 & ~n4928 ;
  assign n4930 = n2387 & n4926 ;
  assign n4931 = n2511 & ~n4930 ;
  assign n4932 = ~n4929 & n4931 ;
  assign n4933 = ~n2511 & ~n4926 ;
  assign n4934 = ~\pi0055  & ~n4933 ;
  assign n4935 = n1292 & n4934 ;
  assign n4936 = n2407 & ~n4755 ;
  assign n4937 = ~n4919 & n4936 ;
  assign n4938 = ~n2407 & ~n4755 ;
  assign n4939 = ~n4754 & n4938 ;
  assign n4940 = ~\pi0062  & ~n4939 ;
  assign n4941 = n4934 & n4940 ;
  assign n4942 = ~n4937 & n4941 ;
  assign n4943 = ~n4935 & ~n4942 ;
  assign n4944 = ~n4932 & ~n4943 ;
  assign n4945 = \pi0105  & ~n4748 ;
  assign n4946 = n4746 & ~n4945 ;
  assign n4947 = ~n1633 & n4946 ;
  assign n4948 = ~n2716 & n4947 ;
  assign n4949 = n2225 & ~n4745 ;
  assign n4950 = ~\pi0216  & ~n4949 ;
  assign n4951 = ~n4948 & n4950 ;
  assign n4952 = \pi0169  & n1640 ;
  assign n4953 = ~n2591 & n4952 ;
  assign n4954 = ~n2704 & n4953 ;
  assign n4955 = \pi0877  & n4954 ;
  assign n4956 = ~\pi0228  & n4955 ;
  assign n4957 = ~n2716 & n4748 ;
  assign n4958 = ~n1639 & ~n4957 ;
  assign n4959 = ~\pi0877  & n2591 ;
  assign n4960 = ~\pi0877  & ~n2580 ;
  assign n4961 = n2574 & n4960 ;
  assign n4962 = ~n4959 & ~n4961 ;
  assign n4963 = n4958 & n4962 ;
  assign n4964 = n4751 & ~n4963 ;
  assign n4965 = ~n4956 & ~n4964 ;
  assign n4966 = n4951 & n4965 ;
  assign n4967 = ~\pi0215  & n4737 ;
  assign n4968 = ~n4966 & n4967 ;
  assign n4969 = ~\pi0038  & ~n4773 ;
  assign n4970 = n4772 & n4969 ;
  assign n4971 = ~n3972 & ~n4970 ;
  assign n4972 = ~\pi0299  & ~n4971 ;
  assign n4973 = ~n4755 & ~n4971 ;
  assign n4974 = ~n4919 & n4973 ;
  assign n4975 = ~n4972 & ~n4974 ;
  assign n4976 = ~n1288 & n4975 ;
  assign n4977 = ~\pi0215  & ~n4742 ;
  assign n4978 = n4854 & ~n4977 ;
  assign n4979 = ~n4976 & n4978 ;
  assign n4980 = ~n4968 & n4979 ;
  assign n4981 = ~n4874 & ~n4875 ;
  assign n4982 = ~\pi0039  & ~n4868 ;
  assign n4983 = ~\pi0039  & ~n4859 ;
  assign n4984 = n4866 & n4983 ;
  assign n4985 = ~n4982 & ~n4984 ;
  assign n4986 = n4981 & ~n4985 ;
  assign n4987 = \pi0038  & ~n4773 ;
  assign n4988 = n4772 & n4987 ;
  assign n4989 = ~n3987 & ~n4988 ;
  assign n4990 = ~\pi0100  & n4989 ;
  assign n4991 = ~n4754 & ~n4755 ;
  assign n4992 = n2563 & ~n4991 ;
  assign n4993 = ~n4990 & ~n4992 ;
  assign n4994 = ~\pi0087  & ~n4993 ;
  assign n4995 = n4986 & n4994 ;
  assign n4996 = ~n1288 & n4994 ;
  assign n4997 = n4975 & n4996 ;
  assign n4998 = ~n4995 & ~n4997 ;
  assign n4999 = ~n4980 & ~n4998 ;
  assign n5000 = ~n1288 & ~n4926 ;
  assign n5001 = n1288 & ~n4773 ;
  assign n5002 = n4772 & n5001 ;
  assign n5003 = ~n4002 & ~n5002 ;
  assign n5004 = \pi0100  & n5003 ;
  assign n5005 = ~n5000 & n5004 ;
  assign n5006 = n4737 & n4750 ;
  assign n5007 = n4831 & ~n5006 ;
  assign n5008 = ~n4829 & n5007 ;
  assign n5009 = n4834 & ~n5000 ;
  assign n5010 = ~n5008 & n5009 ;
  assign n5011 = ~n5005 & ~n5010 ;
  assign n5012 = ~\pi0087  & ~n5011 ;
  assign n5013 = ~n2328 & ~n4926 ;
  assign n5014 = \pi0087  & ~n5013 ;
  assign n5015 = n4922 & n5014 ;
  assign n5016 = ~\pi0075  & ~n5015 ;
  assign n5017 = ~n5012 & n5016 ;
  assign n5018 = ~n4999 & n5017 ;
  assign n5019 = \pi0075  & ~n4773 ;
  assign n5020 = n4772 & n5019 ;
  assign n5021 = ~n4021 & ~n5020 ;
  assign n5022 = ~\pi0092  & n5021 ;
  assign n5023 = n2633 & ~n4991 ;
  assign n5024 = ~n5022 & ~n5023 ;
  assign n5025 = ~n4943 & ~n5024 ;
  assign n5026 = ~n5018 & n5025 ;
  assign n5027 = ~n4944 & ~n5026 ;
  assign n5028 = ~n4754 & n4791 ;
  assign n5029 = \pi0055  & ~n5028 ;
  assign n5030 = ~\pi0056  & ~n5029 ;
  assign n5031 = ~\pi0056  & n4789 ;
  assign n5032 = ~n4919 & n5031 ;
  assign n5033 = ~n5030 & ~n5032 ;
  assign n5034 = ~n4937 & n4940 ;
  assign n5035 = ~n1292 & ~n5034 ;
  assign n5036 = n5033 & ~n5035 ;
  assign n5037 = ~\pi0246  & n2467 ;
  assign n5038 = ~n2504 & ~n4755 ;
  assign n5039 = ~n4754 & n5038 ;
  assign n5040 = \pi0062  & ~n5039 ;
  assign n5041 = ~\pi0056  & ~n4755 ;
  assign n5042 = n2404 & n5041 ;
  assign n5043 = n2403 & n5042 ;
  assign n5044 = ~n4919 & n5043 ;
  assign n5045 = n5040 & ~n5044 ;
  assign n5046 = n5037 & ~n5045 ;
  assign n5047 = ~n5036 & n5046 ;
  assign n5048 = n5027 & n5047 ;
  assign n5049 = ~\pi0055  & ~n4755 ;
  assign n5050 = n1291 & n5049 ;
  assign n5051 = ~n4788 & n5050 ;
  assign n5052 = ~n2407 & n4758 ;
  assign n5053 = ~n4754 & n5052 ;
  assign n5054 = ~\pi0062  & ~n5053 ;
  assign n5055 = ~n5051 & n5054 ;
  assign n5056 = ~n1292 & ~n5055 ;
  assign n5057 = n4910 & n5056 ;
  assign n5058 = \pi0246  & n4757 ;
  assign n5059 = ~n2467 & ~n5058 ;
  assign n5060 = ~n4755 & n5059 ;
  assign n5061 = ~n4754 & n5060 ;
  assign n5062 = ~n5057 & ~n5061 ;
  assign n5063 = ~n5048 & n5062 ;
  assign n5064 = ~n4912 & n5063 ;
  assign n5065 = \pi0216  & \pi0280  ;
  assign n5066 = ~\pi0221  & ~n5065 ;
  assign n5067 = \pi0221  & \pi1137  ;
  assign n5068 = ~n1220 & n5067 ;
  assign n5069 = \pi0221  & \pi0933  ;
  assign n5070 = n1220 & n5069 ;
  assign n5071 = ~n5068 & ~n5070 ;
  assign n5072 = ~n5066 & n5071 ;
  assign n5073 = ~\pi0215  & ~n5072 ;
  assign n5074 = ~\pi0105  & \pi0168  ;
  assign n5075 = \pi0228  & ~n5074 ;
  assign n5076 = ~\pi0216  & ~n5075 ;
  assign n5077 = \pi0878  & ~n1633 ;
  assign n5078 = n3746 & ~n5077 ;
  assign n5079 = ~n5076 & ~n5078 ;
  assign n5080 = ~\pi0168  & ~\pi0228  ;
  assign n5081 = n5071 & ~n5080 ;
  assign n5082 = ~n5079 & n5081 ;
  assign n5083 = n5073 & ~n5082 ;
  assign n5084 = \pi0215  & \pi1137  ;
  assign n5085 = n1295 & ~n5065 ;
  assign n5086 = n2651 & n5085 ;
  assign n5087 = ~n5084 & ~n5086 ;
  assign n5088 = ~n5083 & n5087 ;
  assign n5089 = \pi0299  & ~n5088 ;
  assign n5090 = \pi0222  & \pi1137  ;
  assign n5091 = ~n2192 & n5090 ;
  assign n5092 = \pi0222  & \pi0933  ;
  assign n5093 = n2192 & n5092 ;
  assign n5094 = ~n5091 & ~n5093 ;
  assign n5095 = ~\pi0223  & ~n5094 ;
  assign n5096 = ~\pi0224  & ~n5077 ;
  assign n5097 = \pi0224  & \pi0280  ;
  assign n5098 = ~\pi0222  & ~n5097 ;
  assign n5099 = ~\pi0223  & n5098 ;
  assign n5100 = ~n5096 & n5099 ;
  assign n5101 = ~n5095 & ~n5100 ;
  assign n5102 = \pi0223  & \pi1137  ;
  assign n5103 = ~n3045 & ~n5102 ;
  assign n5104 = n5101 & n5103 ;
  assign n5105 = ~\pi0299  & ~n5104 ;
  assign n5106 = ~n2511 & ~n5105 ;
  assign n5107 = ~n5089 & n5106 ;
  assign n5108 = ~\pi0055  & ~n5107 ;
  assign n5109 = \pi0168  & ~n2280 ;
  assign n5110 = ~\pi0878  & n1281 ;
  assign n5111 = n1260 & n5110 ;
  assign n5112 = ~\pi0228  & ~n5111 ;
  assign n5113 = ~n5109 & n5112 ;
  assign n5114 = ~n2651 & n5071 ;
  assign n5115 = ~n5079 & n5114 ;
  assign n5116 = ~n5113 & n5115 ;
  assign n5117 = n5073 & ~n5116 ;
  assign n5118 = n1291 & ~n5084 ;
  assign n5119 = ~n5117 & n5118 ;
  assign n5120 = ~n1291 & ~n5084 ;
  assign n5121 = ~n5086 & n5120 ;
  assign n5122 = ~n5083 & n5121 ;
  assign n5123 = \pi0055  & ~n5122 ;
  assign n5124 = ~n5119 & n5123 ;
  assign n5125 = ~n5108 & ~n5124 ;
  assign n5126 = n2328 & ~n5105 ;
  assign n5127 = ~\pi0299  & n5126 ;
  assign n5128 = ~n5084 & n5126 ;
  assign n5129 = ~n5117 & n5128 ;
  assign n5130 = ~n5127 & ~n5129 ;
  assign n5131 = ~n2328 & ~n5105 ;
  assign n5132 = ~n5089 & n5131 ;
  assign n5133 = \pi0087  & ~n5132 ;
  assign n5134 = n5130 & n5133 ;
  assign n5135 = ~\pi0075  & ~n5134 ;
  assign n5136 = \pi0075  & ~n5105 ;
  assign n5137 = ~n5089 & n5136 ;
  assign n5138 = ~\pi0092  & ~n5137 ;
  assign n5139 = ~n5135 & n5138 ;
  assign n5140 = \pi0038  & ~n5105 ;
  assign n5141 = ~n5089 & n5140 ;
  assign n5142 = ~\pi0100  & ~n5141 ;
  assign n5143 = ~n1288 & ~n5105 ;
  assign n5144 = ~n5089 & n5143 ;
  assign n5145 = n1288 & ~n5105 ;
  assign n5146 = \pi0100  & ~n5145 ;
  assign n5147 = ~n5144 & n5146 ;
  assign n5148 = ~n2651 & ~n5079 ;
  assign n5149 = n5066 & ~n5148 ;
  assign n5150 = ~\pi0878  & ~n2618 ;
  assign n5151 = ~n2615 & n5150 ;
  assign n5152 = ~\pi0228  & ~n5151 ;
  assign n5153 = \pi0168  & n2618 ;
  assign n5154 = \pi0168  & ~n2609 ;
  assign n5155 = n2614 & n5154 ;
  assign n5156 = ~n5153 & ~n5155 ;
  assign n5157 = n5066 & n5156 ;
  assign n5158 = n5152 & n5157 ;
  assign n5159 = ~n5149 & ~n5158 ;
  assign n5160 = n5071 & ~n5084 ;
  assign n5161 = n5159 & n5160 ;
  assign n5162 = \pi0215  & ~\pi1137  ;
  assign n5163 = n2960 & ~n5162 ;
  assign n5164 = ~n5144 & n5163 ;
  assign n5165 = ~n5161 & n5164 ;
  assign n5166 = ~n5147 & ~n5165 ;
  assign n5167 = ~n5142 & n5166 ;
  assign n5168 = ~\pi0878  & n1640 ;
  assign n5169 = ~n2591 & n5168 ;
  assign n5170 = ~n2704 & n5169 ;
  assign n5171 = ~\pi0168  & ~n5170 ;
  assign n5172 = ~\pi0878  & n2718 ;
  assign n5173 = \pi0168  & ~n5172 ;
  assign n5174 = n3124 & n5173 ;
  assign n5175 = ~n2581 & n5174 ;
  assign n5176 = \pi0168  & ~\pi0878  ;
  assign n5177 = ~n2718 & n5176 ;
  assign n5178 = ~n5175 & ~n5177 ;
  assign n5179 = ~n5171 & n5178 ;
  assign n5180 = n3668 & ~n5065 ;
  assign n5181 = ~n5179 & n5180 ;
  assign n5182 = n3853 & ~n5079 ;
  assign n5183 = n5066 & ~n5182 ;
  assign n5184 = \pi0299  & ~n5084 ;
  assign n5185 = n5071 & n5184 ;
  assign n5186 = ~n5183 & n5185 ;
  assign n5187 = ~n5181 & n5186 ;
  assign n5188 = ~\pi1137  & n2259 ;
  assign n5189 = n5094 & ~n5098 ;
  assign n5190 = n2192 & ~n5092 ;
  assign n5191 = n3503 & ~n5090 ;
  assign n5192 = ~n5190 & ~n5191 ;
  assign n5193 = ~n5077 & ~n5192 ;
  assign n5194 = ~\pi0095  & ~n5192 ;
  assign n5195 = n2686 & n5194 ;
  assign n5196 = ~n5193 & ~n5195 ;
  assign n5197 = ~n5189 & n5196 ;
  assign n5198 = ~\pi0299  & ~n5102 ;
  assign n5199 = n1633 & n5098 ;
  assign n5200 = ~\pi0095  & n5098 ;
  assign n5201 = n2686 & n5200 ;
  assign n5202 = ~n5199 & ~n5201 ;
  assign n5203 = n5198 & n5202 ;
  assign n5204 = ~n5197 & n5203 ;
  assign n5205 = ~\pi1137  & n3498 ;
  assign n5206 = ~\pi0039  & ~n5205 ;
  assign n5207 = ~n5204 & n5206 ;
  assign n5208 = ~n5188 & n5207 ;
  assign n5209 = ~n5187 & n5208 ;
  assign n5210 = ~\pi0038  & ~n5105 ;
  assign n5211 = ~\pi0299  & n5210 ;
  assign n5212 = ~n5084 & n5210 ;
  assign n5213 = ~n5117 & n5212 ;
  assign n5214 = ~n5211 & ~n5213 ;
  assign n5215 = ~n1288 & n5214 ;
  assign n5216 = n5166 & ~n5215 ;
  assign n5217 = ~n5209 & n5216 ;
  assign n5218 = ~n5167 & ~n5217 ;
  assign n5219 = ~\pi0087  & n5138 ;
  assign n5220 = n5218 & n5219 ;
  assign n5221 = ~n5139 & ~n5220 ;
  assign n5222 = ~n1286 & ~n5105 ;
  assign n5223 = ~n5089 & n5222 ;
  assign n5224 = \pi0092  & ~n5223 ;
  assign n5225 = ~n5132 & n5224 ;
  assign n5226 = n5130 & n5225 ;
  assign n5227 = n2387 & ~n5223 ;
  assign n5228 = n2511 & ~n5227 ;
  assign n5229 = ~n5226 & n5228 ;
  assign n5230 = ~n5124 & n5229 ;
  assign n5231 = n5221 & n5230 ;
  assign n5232 = ~n5125 & ~n5231 ;
  assign n5233 = n2504 & ~n5084 ;
  assign n5234 = ~n5117 & n5233 ;
  assign n5235 = ~n2504 & n5087 ;
  assign n5236 = ~n5083 & n5235 ;
  assign n5237 = \pi0062  & ~n5236 ;
  assign n5238 = ~n5234 & n5237 ;
  assign n5239 = \pi0240  & n2467 ;
  assign n5240 = ~n5238 & n5239 ;
  assign n5241 = ~\pi0056  & n5240 ;
  assign n5242 = ~n5232 & n5241 ;
  assign n5243 = n2328 & ~n5102 ;
  assign n5244 = n5101 & n5243 ;
  assign n5245 = ~n3915 & ~n5244 ;
  assign n5246 = ~\pi0299  & ~n5245 ;
  assign n5247 = n5071 & ~n5079 ;
  assign n5248 = ~n5113 & n5247 ;
  assign n5249 = n5073 & ~n5248 ;
  assign n5250 = ~n5084 & ~n5245 ;
  assign n5251 = ~n5249 & n5250 ;
  assign n5252 = ~n5246 & ~n5251 ;
  assign n5253 = n5101 & ~n5102 ;
  assign n5254 = ~\pi0299  & ~n5253 ;
  assign n5255 = n2256 & ~n5072 ;
  assign n5256 = ~n5082 & n5255 ;
  assign n5257 = \pi0299  & n5084 ;
  assign n5258 = ~n1286 & ~n5257 ;
  assign n5259 = ~n5256 & n5258 ;
  assign n5260 = ~n5254 & n5259 ;
  assign n5261 = \pi0092  & ~n5260 ;
  assign n5262 = ~n2328 & ~n5257 ;
  assign n5263 = ~n5256 & n5262 ;
  assign n5264 = ~n5254 & n5263 ;
  assign n5265 = n5261 & ~n5264 ;
  assign n5266 = n5252 & n5265 ;
  assign n5267 = ~n5256 & ~n5257 ;
  assign n5268 = ~n5254 & n5267 ;
  assign n5269 = n2387 & ~n5268 ;
  assign n5270 = n2511 & ~n5269 ;
  assign n5271 = ~n5266 & n5270 ;
  assign n5272 = ~n2511 & ~n5257 ;
  assign n5273 = ~n5256 & n5272 ;
  assign n5274 = ~n5254 & n5273 ;
  assign n5275 = ~\pi0055  & ~n5274 ;
  assign n5276 = n1292 & n5275 ;
  assign n5277 = n2407 & ~n5084 ;
  assign n5278 = ~n5249 & n5277 ;
  assign n5279 = ~n2407 & ~n5084 ;
  assign n5280 = ~n5083 & n5279 ;
  assign n5281 = ~\pi0062  & ~n5280 ;
  assign n5282 = n5275 & n5281 ;
  assign n5283 = ~n5278 & n5282 ;
  assign n5284 = ~n5276 & ~n5283 ;
  assign n5285 = ~n5271 & ~n5284 ;
  assign n5286 = \pi0105  & ~n5077 ;
  assign n5287 = n5075 & ~n5286 ;
  assign n5288 = ~n1633 & n5287 ;
  assign n5289 = ~n2716 & n5288 ;
  assign n5290 = n2225 & ~n5074 ;
  assign n5291 = ~\pi0216  & ~n5290 ;
  assign n5292 = ~n5289 & n5291 ;
  assign n5293 = \pi0168  & n1640 ;
  assign n5294 = ~n2591 & n5293 ;
  assign n5295 = ~n2704 & n5294 ;
  assign n5296 = \pi0878  & n5295 ;
  assign n5297 = ~\pi0228  & n5296 ;
  assign n5298 = ~n2716 & n5077 ;
  assign n5299 = ~n1639 & ~n5298 ;
  assign n5300 = ~\pi0878  & n2591 ;
  assign n5301 = ~\pi0878  & ~n2580 ;
  assign n5302 = n2574 & n5301 ;
  assign n5303 = ~n5300 & ~n5302 ;
  assign n5304 = n5299 & n5303 ;
  assign n5305 = n5080 & ~n5304 ;
  assign n5306 = ~n5297 & ~n5305 ;
  assign n5307 = n5292 & n5306 ;
  assign n5308 = ~\pi0215  & n5066 ;
  assign n5309 = ~n5307 & n5308 ;
  assign n5310 = ~\pi0038  & ~n5102 ;
  assign n5311 = n5101 & n5310 ;
  assign n5312 = ~n3972 & ~n5311 ;
  assign n5313 = ~\pi0299  & ~n5312 ;
  assign n5314 = ~n5084 & ~n5312 ;
  assign n5315 = ~n5249 & n5314 ;
  assign n5316 = ~n5313 & ~n5315 ;
  assign n5317 = ~n1288 & n5316 ;
  assign n5318 = ~\pi0215  & ~n5071 ;
  assign n5319 = n5184 & ~n5318 ;
  assign n5320 = ~n5317 & n5319 ;
  assign n5321 = ~n5309 & n5320 ;
  assign n5322 = ~n5197 & n5198 ;
  assign n5323 = n5207 & ~n5322 ;
  assign n5324 = \pi0038  & ~n5102 ;
  assign n5325 = n5101 & n5324 ;
  assign n5326 = ~n3987 & ~n5325 ;
  assign n5327 = n5267 & ~n5326 ;
  assign n5328 = n2362 & ~n5327 ;
  assign n5329 = n5323 & n5328 ;
  assign n5330 = ~n1288 & n5328 ;
  assign n5331 = n5316 & n5330 ;
  assign n5332 = ~n5329 & ~n5331 ;
  assign n5333 = ~n5321 & ~n5332 ;
  assign n5334 = ~n1288 & ~n5257 ;
  assign n5335 = ~n5256 & n5334 ;
  assign n5336 = ~n5254 & n5335 ;
  assign n5337 = n1288 & ~n5102 ;
  assign n5338 = n5101 & n5337 ;
  assign n5339 = ~n4002 & ~n5338 ;
  assign n5340 = \pi0100  & n5339 ;
  assign n5341 = ~n5336 & n5340 ;
  assign n5342 = n5066 & n5079 ;
  assign n5343 = ~n5158 & ~n5342 ;
  assign n5344 = n5160 & n5343 ;
  assign n5345 = n5163 & ~n5336 ;
  assign n5346 = ~n5344 & n5345 ;
  assign n5347 = ~n5341 & ~n5346 ;
  assign n5348 = ~\pi0087  & ~n5347 ;
  assign n5349 = \pi0087  & ~n5264 ;
  assign n5350 = n5252 & n5349 ;
  assign n5351 = ~\pi0075  & ~n5350 ;
  assign n5352 = ~n5348 & n5351 ;
  assign n5353 = ~n5333 & n5352 ;
  assign n5354 = \pi0075  & ~n5102 ;
  assign n5355 = n5101 & n5354 ;
  assign n5356 = ~n4021 & ~n5355 ;
  assign n5357 = n5267 & ~n5356 ;
  assign n5358 = ~\pi0092  & ~n5357 ;
  assign n5359 = ~n5284 & n5358 ;
  assign n5360 = ~n5353 & n5359 ;
  assign n5361 = ~n5285 & ~n5360 ;
  assign n5362 = ~n5083 & n5120 ;
  assign n5363 = \pi0055  & ~n5362 ;
  assign n5364 = ~\pi0056  & ~n5363 ;
  assign n5365 = ~\pi0056  & n5118 ;
  assign n5366 = ~n5249 & n5365 ;
  assign n5367 = ~n5364 & ~n5366 ;
  assign n5368 = ~n5278 & n5281 ;
  assign n5369 = ~n1292 & ~n5368 ;
  assign n5370 = n5367 & ~n5369 ;
  assign n5371 = ~\pi0240  & n2467 ;
  assign n5372 = ~n2504 & ~n5084 ;
  assign n5373 = ~n5083 & n5372 ;
  assign n5374 = \pi0062  & ~n5373 ;
  assign n5375 = ~\pi0056  & ~n5084 ;
  assign n5376 = n2404 & n5375 ;
  assign n5377 = n2403 & n5376 ;
  assign n5378 = ~n5249 & n5377 ;
  assign n5379 = n5374 & ~n5378 ;
  assign n5380 = n5371 & ~n5379 ;
  assign n5381 = ~n5370 & n5380 ;
  assign n5382 = n5361 & n5381 ;
  assign n5383 = ~\pi0055  & ~n5084 ;
  assign n5384 = n1291 & n5383 ;
  assign n5385 = ~n5117 & n5384 ;
  assign n5386 = ~n2407 & n5087 ;
  assign n5387 = ~n5083 & n5386 ;
  assign n5388 = ~\pi0062  & ~n5387 ;
  assign n5389 = ~n5385 & n5388 ;
  assign n5390 = ~n1292 & ~n5389 ;
  assign n5391 = n5240 & n5390 ;
  assign n5392 = \pi0240  & n5086 ;
  assign n5393 = ~n2467 & ~n5392 ;
  assign n5394 = ~n5084 & n5393 ;
  assign n5395 = ~n5083 & n5394 ;
  assign n5396 = ~n5391 & ~n5395 ;
  assign n5397 = ~n5382 & n5396 ;
  assign n5398 = ~n5242 & n5397 ;
  assign n5399 = ~\pi0245  & n2467 ;
  assign n5400 = \pi0875  & ~n1633 ;
  assign n5401 = n1209 & ~n5400 ;
  assign n5402 = ~\pi0105  & ~\pi0166  ;
  assign n5403 = ~\pi0166  & ~\pi0228  ;
  assign n5404 = ~n5402 & ~n5403 ;
  assign n5405 = n2352 & n5404 ;
  assign n5406 = ~n5401 & n5405 ;
  assign n5407 = \pi0221  & \pi1136  ;
  assign n5408 = ~n1220 & n5407 ;
  assign n5409 = \pi0221  & \pi0928  ;
  assign n5410 = n1220 & n5409 ;
  assign n5411 = ~n5408 & ~n5410 ;
  assign n5412 = \pi0215  & \pi1136  ;
  assign n5413 = \pi0216  & \pi0266  ;
  assign n5414 = ~\pi0221  & n5413 ;
  assign n5415 = ~n5412 & ~n5414 ;
  assign n5416 = n5411 & n5415 ;
  assign n5417 = ~n5406 & n5416 ;
  assign n5418 = \pi0215  & ~\pi1136  ;
  assign n5419 = ~\pi0245  & ~n5418 ;
  assign n5420 = ~n5417 & n5419 ;
  assign n5421 = ~n5399 & ~n5420 ;
  assign n5422 = ~\pi0224  & ~\pi0875  ;
  assign n5423 = ~n1633 & n5422 ;
  assign n5424 = \pi0224  & ~\pi0266  ;
  assign n5425 = ~\pi0222  & ~n5424 ;
  assign n5426 = ~n5423 & n5425 ;
  assign n5427 = \pi0222  & \pi1136  ;
  assign n5428 = ~n2192 & n5427 ;
  assign n5429 = \pi0222  & \pi0928  ;
  assign n5430 = n2192 & n5429 ;
  assign n5431 = ~n5428 & ~n5430 ;
  assign n5432 = ~n5426 & n5431 ;
  assign n5433 = n3058 & ~n5432 ;
  assign n5434 = \pi0223  & \pi1136  ;
  assign n5435 = ~\pi0299  & n5434 ;
  assign n5436 = n2328 & ~n5435 ;
  assign n5437 = ~n5433 & n5436 ;
  assign n5438 = ~\pi0299  & n5437 ;
  assign n5439 = \pi0221  & n5411 ;
  assign n5440 = ~\pi0215  & ~n5439 ;
  assign n5441 = \pi0166  & ~\pi0228  ;
  assign n5442 = ~n3421 & ~n5441 ;
  assign n5443 = ~\pi0875  & n1259 ;
  assign n5444 = n1281 & n5443 ;
  assign n5445 = n1249 & n5444 ;
  assign n5446 = ~\pi0216  & ~n5445 ;
  assign n5447 = ~n5442 & n5446 ;
  assign n5448 = n5411 & ~n5413 ;
  assign n5449 = ~\pi0105  & \pi0166  ;
  assign n5450 = \pi0105  & \pi0875  ;
  assign n5451 = ~n1633 & n5450 ;
  assign n5452 = ~n5449 & ~n5451 ;
  assign n5453 = n1824 & ~n5452 ;
  assign n5454 = ~\pi0216  & n2651 ;
  assign n5455 = ~n5453 & ~n5454 ;
  assign n5456 = n5448 & n5455 ;
  assign n5457 = ~n5447 & n5456 ;
  assign n5458 = n5440 & ~n5457 ;
  assign n5459 = ~n5412 & n5437 ;
  assign n5460 = ~n5458 & n5459 ;
  assign n5461 = ~n5438 & ~n5460 ;
  assign n5462 = ~n5417 & ~n5418 ;
  assign n5463 = ~n2652 & ~n5435 ;
  assign n5464 = ~n5433 & n5463 ;
  assign n5465 = ~n5462 & n5464 ;
  assign n5466 = ~\pi0299  & ~n5434 ;
  assign n5467 = ~n5433 & n5466 ;
  assign n5468 = \pi0092  & ~n5467 ;
  assign n5469 = ~n5465 & n5468 ;
  assign n5470 = ~n3088 & ~n5469 ;
  assign n5471 = ~n5465 & ~n5467 ;
  assign n5472 = ~n2328 & ~n5471 ;
  assign n5473 = ~n5470 & ~n5472 ;
  assign n5474 = n5461 & n5473 ;
  assign n5475 = n2387 & ~n5467 ;
  assign n5476 = ~n5465 & n5475 ;
  assign n5477 = n2511 & ~n5476 ;
  assign n5478 = ~n5474 & n5477 ;
  assign n5479 = ~\pi0055  & n2511 ;
  assign n5480 = ~\pi0055  & ~n5467 ;
  assign n5481 = ~n5465 & n5480 ;
  assign n5482 = ~n5479 & ~n5481 ;
  assign n5483 = n1292 & ~n5482 ;
  assign n5484 = n1291 & ~n5412 ;
  assign n5485 = ~\pi0055  & n5484 ;
  assign n5486 = ~n5458 & n5485 ;
  assign n5487 = ~\pi0062  & ~n5418 ;
  assign n5488 = ~n5417 & n5487 ;
  assign n5489 = ~n2407 & ~n2652 ;
  assign n5490 = ~\pi0062  & ~n5489 ;
  assign n5491 = ~n5488 & ~n5490 ;
  assign n5492 = ~n5482 & ~n5491 ;
  assign n5493 = ~n5486 & n5492 ;
  assign n5494 = ~n5483 & ~n5493 ;
  assign n5495 = ~n5478 & ~n5494 ;
  assign n5496 = ~\pi0215  & ~n5411 ;
  assign n5497 = \pi0216  & ~n5413 ;
  assign n5498 = ~n5413 & n5452 ;
  assign n5499 = n2713 & n5498 ;
  assign n5500 = ~n5497 & ~n5499 ;
  assign n5501 = n1295 & n5500 ;
  assign n5502 = ~n5496 & ~n5501 ;
  assign n5503 = \pi0166  & ~n1633 ;
  assign n5504 = ~n1639 & n5503 ;
  assign n5505 = ~n2591 & n5504 ;
  assign n5506 = ~n2704 & n5505 ;
  assign n5507 = ~\pi0166  & n2718 ;
  assign n5508 = ~\pi0875  & ~n5507 ;
  assign n5509 = ~n5506 & n5508 ;
  assign n5510 = ~\pi0228  & ~n5509 ;
  assign n5511 = \pi0875  & ~n1639 ;
  assign n5512 = ~n2591 & n5511 ;
  assign n5513 = ~n2581 & n5512 ;
  assign n5514 = \pi0166  & \pi0875  ;
  assign n5515 = ~n5413 & ~n5514 ;
  assign n5516 = ~n5513 & n5515 ;
  assign n5517 = ~n5496 & n5516 ;
  assign n5518 = n5510 & n5517 ;
  assign n5519 = ~n5502 & ~n5518 ;
  assign n5520 = \pi0299  & ~n5412 ;
  assign n5521 = ~n5433 & ~n5435 ;
  assign n5522 = ~\pi0038  & ~\pi0299  ;
  assign n5523 = ~\pi0038  & ~n5412 ;
  assign n5524 = ~n5458 & n5523 ;
  assign n5525 = ~n5522 & ~n5524 ;
  assign n5526 = n5521 & ~n5525 ;
  assign n5527 = ~n1288 & ~n5526 ;
  assign n5528 = n5520 & ~n5527 ;
  assign n5529 = ~n5519 & n5528 ;
  assign n5530 = ~\pi0039  & ~n5466 ;
  assign n5531 = ~n1633 & n5432 ;
  assign n5532 = ~n2716 & n5531 ;
  assign n5533 = ~n2165 & n5432 ;
  assign n5534 = n2692 & ~n5533 ;
  assign n5535 = ~n5532 & n5534 ;
  assign n5536 = ~n5530 & ~n5535 ;
  assign n5537 = n1288 & n5536 ;
  assign n5538 = n5521 & n5536 ;
  assign n5539 = ~n5525 & n5538 ;
  assign n5540 = ~n5537 & ~n5539 ;
  assign n5541 = ~\pi0100  & ~n5467 ;
  assign n5542 = ~n5465 & n5541 ;
  assign n5543 = ~n2327 & ~n5542 ;
  assign n5544 = ~\pi0087  & ~n5543 ;
  assign n5545 = n5540 & n5544 ;
  assign n5546 = ~n5529 & n5545 ;
  assign n5547 = n1288 & ~n5435 ;
  assign n5548 = ~n5433 & n5547 ;
  assign n5549 = \pi0100  & ~n5467 ;
  assign n5550 = ~n5465 & n5549 ;
  assign n5551 = ~n2222 & ~n5550 ;
  assign n5552 = ~n5548 & ~n5551 ;
  assign n5553 = n5411 & ~n5412 ;
  assign n5554 = ~n5414 & n5553 ;
  assign n5555 = \pi0875  & n1259 ;
  assign n5556 = n1249 & n5555 ;
  assign n5557 = n3182 & n5556 ;
  assign n5558 = n1800 & n5557 ;
  assign n5559 = n1259 & ~n1800 ;
  assign n5560 = n1249 & n5559 ;
  assign n5561 = n2616 & n5560 ;
  assign n5562 = \pi0875  & n5561 ;
  assign n5563 = ~n5558 & ~n5562 ;
  assign n5564 = ~\pi0875  & ~n2238 ;
  assign n5565 = n1281 & n5564 ;
  assign n5566 = n1260 & n5565 ;
  assign n5567 = \pi0166  & ~n5566 ;
  assign n5568 = \pi0228  & ~n5452 ;
  assign n5569 = ~n2651 & ~n5568 ;
  assign n5570 = ~n5567 & n5569 ;
  assign n5571 = n5563 & n5570 ;
  assign n5572 = \pi0228  & ~n2651 ;
  assign n5573 = n5452 & n5572 ;
  assign n5574 = n2352 & ~n5573 ;
  assign n5575 = ~n5571 & n5574 ;
  assign n5576 = n5554 & ~n5575 ;
  assign n5577 = n2960 & ~n5418 ;
  assign n5578 = ~n1288 & ~n5471 ;
  assign n5579 = n5577 & ~n5578 ;
  assign n5580 = ~n5576 & n5579 ;
  assign n5581 = ~n5552 & ~n5580 ;
  assign n5582 = ~\pi0087  & ~n5581 ;
  assign n5583 = \pi0087  & n2328 ;
  assign n5584 = \pi0087  & ~n5467 ;
  assign n5585 = ~n5465 & n5584 ;
  assign n5586 = ~n5583 & ~n5585 ;
  assign n5587 = n5461 & ~n5586 ;
  assign n5588 = ~\pi0075  & ~n5587 ;
  assign n5589 = ~n5582 & n5588 ;
  assign n5590 = ~n5546 & n5589 ;
  assign n5591 = ~\pi0092  & ~n5467 ;
  assign n5592 = ~n5465 & n5591 ;
  assign n5593 = ~n2364 & ~n5592 ;
  assign n5594 = ~n5494 & ~n5593 ;
  assign n5595 = ~n5590 & n5594 ;
  assign n5596 = ~n5495 & ~n5595 ;
  assign n5597 = \pi0055  & ~n5418 ;
  assign n5598 = ~n5417 & n5597 ;
  assign n5599 = ~n1291 & ~n2652 ;
  assign n5600 = \pi0055  & ~n5599 ;
  assign n5601 = ~n5598 & ~n5600 ;
  assign n5602 = ~\pi0056  & n5601 ;
  assign n5603 = ~\pi0056  & n5484 ;
  assign n5604 = ~n5458 & n5603 ;
  assign n5605 = ~n5602 & ~n5604 ;
  assign n5606 = ~n5486 & ~n5491 ;
  assign n5607 = ~n1292 & ~n5606 ;
  assign n5608 = n5605 & ~n5607 ;
  assign n5609 = n2504 & ~n5412 ;
  assign n5610 = ~n5458 & n5609 ;
  assign n5611 = \pi0062  & ~n5418 ;
  assign n5612 = ~n5417 & n5611 ;
  assign n5613 = ~n2504 & ~n2652 ;
  assign n5614 = \pi0062  & ~n5613 ;
  assign n5615 = ~n5612 & ~n5614 ;
  assign n5616 = ~n5610 & ~n5615 ;
  assign n5617 = n2467 & ~n5616 ;
  assign n5618 = ~n5608 & n5617 ;
  assign n5619 = n5596 & n5618 ;
  assign n5620 = ~n2467 & ~n2652 ;
  assign n5621 = \pi0245  & ~n5620 ;
  assign n5622 = \pi0245  & ~n5418 ;
  assign n5623 = ~n5417 & n5622 ;
  assign n5624 = ~n5621 & ~n5623 ;
  assign n5625 = ~n5619 & ~n5624 ;
  assign n5626 = n5421 & ~n5625 ;
  assign n5627 = \pi0055  & n1291 ;
  assign n5628 = ~n5598 & ~n5627 ;
  assign n5629 = ~\pi0056  & n5628 ;
  assign n5630 = ~n5413 & ~n5453 ;
  assign n5631 = ~n5447 & n5630 ;
  assign n5632 = n1295 & ~n5631 ;
  assign n5633 = ~n5496 & ~n5632 ;
  assign n5634 = n5603 & n5633 ;
  assign n5635 = ~n5629 & ~n5634 ;
  assign n5636 = n2407 & ~n5412 ;
  assign n5637 = n5633 & n5636 ;
  assign n5638 = ~\pi0062  & n2407 ;
  assign n5639 = ~n5488 & ~n5638 ;
  assign n5640 = ~n5637 & ~n5639 ;
  assign n5641 = ~n1292 & ~n5640 ;
  assign n5642 = n5635 & ~n5641 ;
  assign n5643 = \pi0299  & ~n5418 ;
  assign n5644 = ~n5417 & n5643 ;
  assign n5645 = n2214 & ~n5400 ;
  assign n5646 = n5435 & ~n5645 ;
  assign n5647 = n3058 & ~n5645 ;
  assign n5648 = ~n5432 & n5647 ;
  assign n5649 = ~n5646 & ~n5648 ;
  assign n5650 = ~n5644 & n5649 ;
  assign n5651 = \pi0075  & n5650 ;
  assign n5652 = \pi0100  & ~n5649 ;
  assign n5653 = \pi0100  & ~n1288 ;
  assign n5654 = n5644 & n5653 ;
  assign n5655 = ~n5652 & ~n5654 ;
  assign n5656 = ~n5567 & ~n5568 ;
  assign n5657 = n5563 & n5656 ;
  assign n5658 = \pi0228  & ~n5449 ;
  assign n5659 = ~n5451 & n5658 ;
  assign n5660 = n2352 & ~n5659 ;
  assign n5661 = ~n5657 & n5660 ;
  assign n5662 = n5554 & ~n5661 ;
  assign n5663 = ~n1288 & n5650 ;
  assign n5664 = n5577 & ~n5663 ;
  assign n5665 = ~n5662 & n5664 ;
  assign n5666 = n5655 & ~n5665 ;
  assign n5667 = ~n5651 & ~n5666 ;
  assign n5668 = n1633 & n2165 ;
  assign n5669 = ~\pi0095  & n2165 ;
  assign n5670 = n2686 & n5669 ;
  assign n5671 = ~n5668 & ~n5670 ;
  assign n5672 = n5426 & n5671 ;
  assign n5673 = n5431 & n5466 ;
  assign n5674 = ~n5672 & n5673 ;
  assign n5675 = ~n5536 & ~n5674 ;
  assign n5676 = ~\pi0038  & n5649 ;
  assign n5677 = ~\pi0299  & n5676 ;
  assign n5678 = ~n5412 & n5676 ;
  assign n5679 = n5633 & n5678 ;
  assign n5680 = ~n5677 & ~n5679 ;
  assign n5681 = ~n1288 & n5680 ;
  assign n5682 = ~n5675 & ~n5681 ;
  assign n5683 = \pi0166  & ~\pi0875  ;
  assign n5684 = ~n3125 & n5683 ;
  assign n5685 = n2713 & n5452 ;
  assign n5686 = n2492 & ~n5685 ;
  assign n5687 = n5684 & n5686 ;
  assign n5688 = ~n2704 & n3246 ;
  assign n5689 = ~\pi0166  & ~n5688 ;
  assign n5690 = \pi0166  & ~n2718 ;
  assign n5691 = \pi0875  & ~n5690 ;
  assign n5692 = n5686 & n5691 ;
  assign n5693 = ~n5689 & n5692 ;
  assign n5694 = ~n5687 & ~n5693 ;
  assign n5695 = ~\pi0216  & ~n5452 ;
  assign n5696 = n2713 & n5695 ;
  assign n5697 = n5448 & ~n5696 ;
  assign n5698 = n5694 & n5697 ;
  assign n5699 = n5440 & ~n5698 ;
  assign n5700 = n5520 & ~n5681 ;
  assign n5701 = ~n5699 & n5700 ;
  assign n5702 = ~n5682 & ~n5701 ;
  assign n5703 = \pi0038  & n5649 ;
  assign n5704 = ~n5644 & n5703 ;
  assign n5705 = ~\pi0100  & ~n5704 ;
  assign n5706 = ~n5651 & n5705 ;
  assign n5707 = n5702 & n5706 ;
  assign n5708 = ~n5667 & ~n5707 ;
  assign n5709 = n4539 & ~n5708 ;
  assign n5710 = \pi0075  & n5649 ;
  assign n5711 = ~n5644 & n5710 ;
  assign n5712 = ~\pi0092  & ~n5711 ;
  assign n5713 = \pi0075  & n5712 ;
  assign n5714 = n2328 & n5649 ;
  assign n5715 = ~\pi0299  & n5714 ;
  assign n5716 = ~n5412 & n5714 ;
  assign n5717 = n5633 & n5716 ;
  assign n5718 = ~n5715 & ~n5717 ;
  assign n5719 = ~n2328 & n5650 ;
  assign n5720 = \pi0087  & ~n5719 ;
  assign n5721 = n5712 & n5720 ;
  assign n5722 = n5718 & n5721 ;
  assign n5723 = ~n5713 & ~n5722 ;
  assign n5724 = \pi0092  & ~n5650 ;
  assign n5725 = ~n3089 & ~n5724 ;
  assign n5726 = n5718 & ~n5725 ;
  assign n5727 = n2387 & ~n5650 ;
  assign n5728 = n2511 & ~n5727 ;
  assign n5729 = ~n5726 & n5728 ;
  assign n5730 = n5723 & n5729 ;
  assign n5731 = ~n5709 & n5730 ;
  assign n5732 = ~n2511 & n5649 ;
  assign n5733 = ~n5644 & n5732 ;
  assign n5734 = ~\pi0055  & ~n5733 ;
  assign n5735 = ~n5641 & n5734 ;
  assign n5736 = ~n5731 & n5735 ;
  assign n5737 = ~n5642 & ~n5736 ;
  assign n5738 = ~\pi0056  & ~n5412 ;
  assign n5739 = n2407 & n5738 ;
  assign n5740 = n5633 & n5739 ;
  assign n5741 = \pi0062  & n2504 ;
  assign n5742 = ~n5612 & ~n5741 ;
  assign n5743 = ~n5740 & ~n5742 ;
  assign n5744 = n2467 & ~n5743 ;
  assign n5745 = ~n5625 & n5744 ;
  assign n5746 = n5737 & n5745 ;
  assign n5747 = ~n5626 & ~n5746 ;
  assign n5748 = ~\pi0244  & n2467 ;
  assign n5749 = \pi0221  & \pi1135  ;
  assign n5750 = ~n1220 & n5749 ;
  assign n5751 = \pi0221  & \pi0938  ;
  assign n5752 = n1220 & n5751 ;
  assign n5753 = ~n5750 & ~n5752 ;
  assign n5754 = \pi0215  & \pi1135  ;
  assign n5755 = \pi0216  & \pi0279  ;
  assign n5756 = ~\pi0221  & n5755 ;
  assign n5757 = ~n5754 & ~n5756 ;
  assign n5758 = n5753 & n5757 ;
  assign n5759 = \pi0879  & ~n1633 ;
  assign n5760 = n1209 & ~n5759 ;
  assign n5761 = ~\pi0105  & ~\pi0161  ;
  assign n5762 = ~\pi0161  & ~\pi0228  ;
  assign n5763 = ~n5761 & ~n5762 ;
  assign n5764 = n2352 & n5763 ;
  assign n5765 = ~n5760 & n5764 ;
  assign n5766 = n5758 & ~n5765 ;
  assign n5767 = \pi0215  & ~\pi1135  ;
  assign n5768 = ~\pi0244  & ~n5767 ;
  assign n5769 = ~n5766 & n5768 ;
  assign n5770 = ~n5748 & ~n5769 ;
  assign n5771 = ~\pi0215  & ~n5753 ;
  assign n5772 = \pi0216  & ~n5755 ;
  assign n5773 = ~\pi0105  & \pi0161  ;
  assign n5774 = \pi0105  & \pi0879  ;
  assign n5775 = ~n1633 & n5774 ;
  assign n5776 = ~n5773 & ~n5775 ;
  assign n5777 = ~n5755 & n5776 ;
  assign n5778 = n2713 & n5777 ;
  assign n5779 = ~n5772 & ~n5778 ;
  assign n5780 = n1295 & n5779 ;
  assign n5781 = ~n5771 & ~n5780 ;
  assign n5782 = \pi0161  & ~n1633 ;
  assign n5783 = ~n1639 & n5782 ;
  assign n5784 = ~n2591 & n5783 ;
  assign n5785 = ~n2704 & n5784 ;
  assign n5786 = ~\pi0161  & n2718 ;
  assign n5787 = ~\pi0879  & ~n5786 ;
  assign n5788 = ~n5785 & n5787 ;
  assign n5789 = ~\pi0228  & ~n5788 ;
  assign n5790 = \pi0879  & ~n1639 ;
  assign n5791 = ~n2591 & n5790 ;
  assign n5792 = ~n2581 & n5791 ;
  assign n5793 = \pi0161  & \pi0879  ;
  assign n5794 = ~n5755 & ~n5793 ;
  assign n5795 = ~n5792 & n5794 ;
  assign n5796 = ~n5771 & n5795 ;
  assign n5797 = n5789 & n5796 ;
  assign n5798 = ~n5781 & ~n5797 ;
  assign n5799 = \pi0299  & ~n5754 ;
  assign n5800 = ~n5758 & ~n5767 ;
  assign n5801 = ~\pi0879  & n1281 ;
  assign n5802 = n1260 & n5801 ;
  assign n5803 = \pi0228  & ~n5776 ;
  assign n5804 = ~n2651 & ~n5803 ;
  assign n5805 = n5802 & n5804 ;
  assign n5806 = n2352 & ~n5805 ;
  assign n5807 = \pi0161  & ~\pi0228  ;
  assign n5808 = ~n2651 & ~n5807 ;
  assign n5809 = ~n5803 & n5808 ;
  assign n5810 = ~n3421 & n5809 ;
  assign n5811 = ~n5767 & ~n5810 ;
  assign n5812 = n5806 & n5811 ;
  assign n5813 = ~n5800 & ~n5812 ;
  assign n5814 = n2297 & ~n5813 ;
  assign n5815 = \pi0223  & \pi1135  ;
  assign n5816 = ~\pi0299  & n5815 ;
  assign n5817 = \pi0039  & n5816 ;
  assign n5818 = \pi0222  & \pi1135  ;
  assign n5819 = ~n2192 & n5818 ;
  assign n5820 = \pi0222  & \pi0938  ;
  assign n5821 = n2192 & n5820 ;
  assign n5822 = ~n5819 & ~n5821 ;
  assign n5823 = ~\pi0224  & ~\pi0879  ;
  assign n5824 = ~n1633 & n5823 ;
  assign n5825 = \pi0224  & ~\pi0279  ;
  assign n5826 = ~\pi0222  & ~n5825 ;
  assign n5827 = ~n5824 & n5826 ;
  assign n5828 = n5822 & ~n5827 ;
  assign n5829 = n3268 & ~n5828 ;
  assign n5830 = ~n5817 & ~n5829 ;
  assign n5831 = ~\pi0038  & n5830 ;
  assign n5832 = ~n5814 & n5831 ;
  assign n5833 = n5799 & n5832 ;
  assign n5834 = ~n5798 & n5833 ;
  assign n5835 = ~n1633 & n5828 ;
  assign n5836 = ~n2716 & n5835 ;
  assign n5837 = ~n2165 & n5828 ;
  assign n5838 = n2692 & ~n5837 ;
  assign n5839 = ~n5836 & n5838 ;
  assign n5840 = ~\pi0299  & ~n5815 ;
  assign n5841 = ~\pi0039  & ~n5840 ;
  assign n5842 = n5831 & ~n5841 ;
  assign n5843 = ~n5839 & n5842 ;
  assign n5844 = ~n5814 & n5843 ;
  assign n5845 = ~n5766 & ~n5767 ;
  assign n5846 = n3058 & ~n5828 ;
  assign n5847 = ~n2652 & ~n5816 ;
  assign n5848 = ~n5846 & n5847 ;
  assign n5849 = ~n5845 & n5848 ;
  assign n5850 = n5840 & ~n5846 ;
  assign n5851 = ~\pi0100  & ~n5850 ;
  assign n5852 = ~n5849 & n5851 ;
  assign n5853 = ~n2327 & ~n5852 ;
  assign n5854 = ~\pi0087  & ~n5853 ;
  assign n5855 = ~n5844 & n5854 ;
  assign n5856 = ~n5834 & n5855 ;
  assign n5857 = \pi0299  & ~n5813 ;
  assign n5858 = ~n5816 & ~n5846 ;
  assign n5859 = n2328 & n5858 ;
  assign n5860 = ~n5857 & n5859 ;
  assign n5861 = \pi0087  & ~n5850 ;
  assign n5862 = ~n5849 & n5861 ;
  assign n5863 = ~n5583 & ~n5862 ;
  assign n5864 = ~n5860 & ~n5863 ;
  assign n5865 = ~\pi0075  & ~n5864 ;
  assign n5866 = \pi0092  & ~n5850 ;
  assign n5867 = ~n5849 & n5866 ;
  assign n5868 = ~n3088 & ~n5867 ;
  assign n5869 = ~n5849 & ~n5850 ;
  assign n5870 = ~n2328 & ~n5869 ;
  assign n5871 = ~n5868 & ~n5870 ;
  assign n5872 = ~n5860 & n5871 ;
  assign n5873 = n2387 & ~n5850 ;
  assign n5874 = ~n5849 & n5873 ;
  assign n5875 = n2511 & ~n5874 ;
  assign n5876 = ~n5872 & n5875 ;
  assign n5877 = n1288 & ~n5816 ;
  assign n5878 = ~n5846 & n5877 ;
  assign n5879 = \pi0100  & ~n5850 ;
  assign n5880 = ~n5849 & n5879 ;
  assign n5881 = ~n2222 & ~n5880 ;
  assign n5882 = ~n5878 & ~n5881 ;
  assign n5883 = ~\pi0152  & ~\pi0166  ;
  assign n5884 = n1259 & ~n5883 ;
  assign n5885 = n1249 & n5884 ;
  assign n5886 = n2616 & n5885 ;
  assign n5887 = \pi0879  & n5886 ;
  assign n5888 = \pi0879  & n1259 ;
  assign n5889 = n1249 & n5888 ;
  assign n5890 = n3182 & n5889 ;
  assign n5891 = n5883 & n5890 ;
  assign n5892 = ~n5887 & ~n5891 ;
  assign n5893 = ~\pi0879  & ~n2238 ;
  assign n5894 = n1281 & n5893 ;
  assign n5895 = n1260 & n5894 ;
  assign n5896 = \pi0161  & ~n5895 ;
  assign n5897 = n5804 & ~n5896 ;
  assign n5898 = n5892 & n5897 ;
  assign n5899 = n5572 & n5776 ;
  assign n5900 = n2352 & ~n5899 ;
  assign n5901 = ~n5767 & n5900 ;
  assign n5902 = ~n5898 & n5901 ;
  assign n5903 = ~n5800 & ~n5902 ;
  assign n5904 = ~n1288 & ~n5869 ;
  assign n5905 = n2960 & ~n5904 ;
  assign n5906 = ~n5903 & n5905 ;
  assign n5907 = ~n5882 & ~n5906 ;
  assign n5908 = ~\pi0087  & ~n5907 ;
  assign n5909 = n5876 & ~n5908 ;
  assign n5910 = n5865 & n5909 ;
  assign n5911 = ~n5856 & n5910 ;
  assign n5912 = ~\pi0092  & ~n5850 ;
  assign n5913 = ~n5849 & n5912 ;
  assign n5914 = ~n2364 & ~n5913 ;
  assign n5915 = n5875 & n5914 ;
  assign n5916 = ~n5872 & n5915 ;
  assign n5917 = ~\pi0062  & ~n5767 ;
  assign n5918 = ~n5766 & n5917 ;
  assign n5919 = ~n5490 & ~n5918 ;
  assign n5920 = ~n1292 & n5919 ;
  assign n5921 = ~n1292 & n3030 ;
  assign n5922 = n5813 & n5921 ;
  assign n5923 = ~n5920 & ~n5922 ;
  assign n5924 = ~\pi0055  & ~n5850 ;
  assign n5925 = ~n5849 & n5924 ;
  assign n5926 = ~n5479 & ~n5925 ;
  assign n5927 = n5923 & ~n5926 ;
  assign n5928 = ~n5916 & n5927 ;
  assign n5929 = ~n5911 & n5928 ;
  assign n5930 = \pi0055  & ~n5767 ;
  assign n5931 = ~n5766 & n5930 ;
  assign n5932 = ~n5600 & ~n5931 ;
  assign n5933 = ~\pi0056  & n5932 ;
  assign n5934 = n3008 & n5813 ;
  assign n5935 = ~n5933 & ~n5934 ;
  assign n5936 = n5923 & n5935 ;
  assign n5937 = \pi0062  & ~n5767 ;
  assign n5938 = ~n5766 & n5937 ;
  assign n5939 = ~n5614 & ~n5938 ;
  assign n5940 = n2467 & n5939 ;
  assign n5941 = n2423 & n2467 ;
  assign n5942 = n1291 & n5941 ;
  assign n5943 = n5813 & n5942 ;
  assign n5944 = ~n5940 & ~n5943 ;
  assign n5945 = ~n5936 & ~n5944 ;
  assign n5946 = ~n5929 & n5945 ;
  assign n5947 = \pi0244  & ~n5620 ;
  assign n5948 = \pi0244  & ~n5767 ;
  assign n5949 = ~n5766 & n5948 ;
  assign n5950 = ~n5947 & ~n5949 ;
  assign n5951 = ~n5946 & ~n5950 ;
  assign n5952 = n5770 & ~n5951 ;
  assign n5953 = \pi0299  & ~n5767 ;
  assign n5954 = ~n5766 & n5953 ;
  assign n5955 = n2214 & ~n5759 ;
  assign n5956 = n5816 & ~n5955 ;
  assign n5957 = n3058 & ~n5955 ;
  assign n5958 = ~n5828 & n5957 ;
  assign n5959 = ~n5956 & ~n5958 ;
  assign n5960 = \pi0075  & n5959 ;
  assign n5961 = ~n5954 & n5960 ;
  assign n5962 = ~\pi0092  & ~n5961 ;
  assign n5963 = ~n5627 & ~n5931 ;
  assign n5964 = ~\pi0056  & n5963 ;
  assign n5965 = n3008 & n5767 ;
  assign n5966 = ~n5803 & ~n5807 ;
  assign n5967 = ~n3421 & n5966 ;
  assign n5968 = n1259 & ~n5803 ;
  assign n5969 = n1249 & n5968 ;
  assign n5970 = n5801 & n5969 ;
  assign n5971 = n2352 & ~n5970 ;
  assign n5972 = ~n5967 & n5971 ;
  assign n5973 = n3008 & n5758 ;
  assign n5974 = ~n5972 & n5973 ;
  assign n5975 = ~n5965 & ~n5974 ;
  assign n5976 = ~n5964 & n5975 ;
  assign n5977 = ~n5954 & n5959 ;
  assign n5978 = \pi0092  & ~n5977 ;
  assign n5979 = ~n3089 & ~n5978 ;
  assign n5980 = n2387 & ~n5977 ;
  assign n5981 = n2511 & ~n5980 ;
  assign n5982 = n5979 & n5981 ;
  assign n5983 = n5758 & ~n5972 ;
  assign n5984 = n5953 & ~n5983 ;
  assign n5985 = n2328 & n5959 ;
  assign n5986 = n5981 & n5985 ;
  assign n5987 = ~n5984 & n5986 ;
  assign n5988 = ~n5982 & ~n5987 ;
  assign n5989 = ~n5976 & ~n5988 ;
  assign n5990 = ~n5962 & n5989 ;
  assign n5991 = n2165 & n5822 ;
  assign n5992 = n1633 & n5991 ;
  assign n5993 = ~\pi0095  & n5991 ;
  assign n5994 = n2686 & n5993 ;
  assign n5995 = ~n5992 & ~n5994 ;
  assign n5996 = ~\pi0223  & ~n5828 ;
  assign n5997 = ~\pi0039  & n5996 ;
  assign n5998 = n5995 & n5997 ;
  assign n5999 = ~n5841 & ~n5998 ;
  assign n6000 = ~\pi0215  & ~n5999 ;
  assign n6001 = ~n5753 & n6000 ;
  assign n6002 = n2713 & n5776 ;
  assign n6003 = ~\pi0216  & ~n6002 ;
  assign n6004 = \pi0161  & ~\pi0879  ;
  assign n6005 = ~n3125 & n6004 ;
  assign n6006 = n6003 & n6005 ;
  assign n6007 = ~\pi0161  & ~n5688 ;
  assign n6008 = \pi0161  & ~n2718 ;
  assign n6009 = \pi0879  & ~n6008 ;
  assign n6010 = n6003 & n6009 ;
  assign n6011 = ~n6007 & n6010 ;
  assign n6012 = ~n6006 & ~n6011 ;
  assign n6013 = ~\pi0228  & ~n6012 ;
  assign n6014 = ~\pi0216  & ~n5776 ;
  assign n6015 = n2713 & n6014 ;
  assign n6016 = ~n5755 & ~n6015 ;
  assign n6017 = ~n6013 & n6016 ;
  assign n6018 = ~\pi0221  & n6000 ;
  assign n6019 = ~n6017 & n6018 ;
  assign n6020 = ~n6001 & ~n6019 ;
  assign n6021 = ~n5803 & ~n5896 ;
  assign n6022 = n5892 & n6021 ;
  assign n6023 = \pi0228  & ~n5773 ;
  assign n6024 = ~n5775 & n6023 ;
  assign n6025 = n2352 & ~n6024 ;
  assign n6026 = ~n5767 & n6025 ;
  assign n6027 = ~n6022 & n6026 ;
  assign n6028 = ~n5800 & ~n6027 ;
  assign n6029 = ~n1288 & n5977 ;
  assign n6030 = n2960 & ~n6029 ;
  assign n6031 = ~n6028 & n6030 ;
  assign n6032 = ~n5799 & ~n5999 ;
  assign n6033 = n2297 & ~n5767 ;
  assign n6034 = ~n5983 & n6033 ;
  assign n6035 = \pi0100  & ~n5959 ;
  assign n6036 = n5653 & n5954 ;
  assign n6037 = ~n6035 & ~n6036 ;
  assign n6038 = \pi0039  & ~n5959 ;
  assign n6039 = ~\pi0038  & ~n6038 ;
  assign n6040 = n6037 & n6039 ;
  assign n6041 = ~n6034 & n6040 ;
  assign n6042 = ~n6032 & n6041 ;
  assign n6043 = ~n6031 & n6042 ;
  assign n6044 = n6020 & n6043 ;
  assign n6045 = \pi0038  & n5959 ;
  assign n6046 = ~n5954 & n6045 ;
  assign n6047 = ~\pi0100  & ~n6046 ;
  assign n6048 = n6037 & ~n6047 ;
  assign n6049 = ~n6031 & n6048 ;
  assign n6050 = ~\pi0087  & ~n6049 ;
  assign n6051 = ~n6044 & n6050 ;
  assign n6052 = ~n2328 & n5977 ;
  assign n6053 = \pi0087  & ~n6052 ;
  assign n6054 = ~\pi0075  & ~n6053 ;
  assign n6055 = ~\pi0075  & n5985 ;
  assign n6056 = ~n5984 & n6055 ;
  assign n6057 = ~n6054 & ~n6056 ;
  assign n6058 = n5989 & ~n6057 ;
  assign n6059 = ~n6051 & n6058 ;
  assign n6060 = ~n5990 & ~n6059 ;
  assign n6061 = ~n2511 & n5959 ;
  assign n6062 = ~n5954 & n6061 ;
  assign n6063 = ~\pi0055  & ~n6062 ;
  assign n6064 = ~n5976 & ~n6063 ;
  assign n6065 = n2406 & n5767 ;
  assign n6066 = n2406 & n5758 ;
  assign n6067 = ~n5972 & n6066 ;
  assign n6068 = ~n6065 & ~n6067 ;
  assign n6069 = \pi0056  & ~n2407 ;
  assign n6070 = ~n5845 & n6069 ;
  assign n6071 = ~\pi0062  & ~n6070 ;
  assign n6072 = n6068 & n6071 ;
  assign n6073 = ~n6064 & n6072 ;
  assign n6074 = n6060 & n6073 ;
  assign n6075 = n2454 & n5767 ;
  assign n6076 = n2454 & n5758 ;
  assign n6077 = ~n5972 & n6076 ;
  assign n6078 = ~n6075 & ~n6077 ;
  assign n6079 = ~n5741 & ~n5938 ;
  assign n6080 = n6078 & ~n6079 ;
  assign n6081 = n2467 & ~n6080 ;
  assign n6082 = ~n5951 & n6081 ;
  assign n6083 = ~n6074 & n6082 ;
  assign n6084 = ~n5952 & ~n6083 ;
  assign n6085 = \pi0152  & ~\pi0228  ;
  assign n6086 = ~n3421 & ~n6085 ;
  assign n6087 = ~\pi0846  & n1259 ;
  assign n6088 = n1281 & n6087 ;
  assign n6089 = n1249 & n6088 ;
  assign n6090 = ~\pi0216  & ~n6089 ;
  assign n6091 = ~n6086 & n6090 ;
  assign n6092 = \pi0216  & \pi0278  ;
  assign n6093 = ~\pi0221  & ~n6092 ;
  assign n6094 = ~\pi0105  & \pi0152  ;
  assign n6095 = \pi0105  & \pi0846  ;
  assign n6096 = ~n1633 & n6095 ;
  assign n6097 = ~n6094 & ~n6096 ;
  assign n6098 = n1824 & ~n6097 ;
  assign n6099 = ~n5454 & ~n6098 ;
  assign n6100 = n6093 & n6099 ;
  assign n6101 = ~n6091 & n6100 ;
  assign n6102 = \pi0833  & ~\pi0930  ;
  assign n6103 = ~\pi0216  & \pi0221  ;
  assign n6104 = n6102 & n6103 ;
  assign n6105 = ~n6101 & ~n6104 ;
  assign n6106 = ~\pi0215  & n5942 ;
  assign n6107 = ~n6105 & n6106 ;
  assign n6108 = ~n2504 & n3409 ;
  assign n6109 = \pi0062  & ~n6108 ;
  assign n6110 = ~n6085 & ~n6094 ;
  assign n6111 = ~n6096 & n6110 ;
  assign n6112 = ~\pi0152  & ~\pi0228  ;
  assign n6113 = ~\pi0216  & ~n6112 ;
  assign n6114 = ~n6111 & n6113 ;
  assign n6115 = n6093 & ~n6114 ;
  assign n6116 = \pi0062  & ~n6104 ;
  assign n6117 = ~n6115 & n6116 ;
  assign n6118 = ~n6109 & ~n6117 ;
  assign n6119 = n2467 & n6118 ;
  assign n6120 = ~\pi0215  & ~n2467 ;
  assign n6121 = n6104 & n6120 ;
  assign n6122 = n6093 & n6120 ;
  assign n6123 = ~n6114 & n6122 ;
  assign n6124 = ~n6121 & ~n6123 ;
  assign n6125 = ~n2652 & ~n6124 ;
  assign n6126 = \pi0242  & ~n6125 ;
  assign n6127 = ~n6119 & n6126 ;
  assign n6128 = ~n6107 & n6127 ;
  assign n6129 = ~\pi0152  & \pi0846  ;
  assign n6130 = ~n3125 & n6129 ;
  assign n6131 = n6093 & n6130 ;
  assign n6132 = \pi0152  & ~n5688 ;
  assign n6133 = ~\pi0152  & ~n2718 ;
  assign n6134 = ~\pi0846  & ~n6133 ;
  assign n6135 = n6093 & n6134 ;
  assign n6136 = ~n6132 & n6135 ;
  assign n6137 = ~n6131 & ~n6136 ;
  assign n6138 = ~\pi0228  & ~n6137 ;
  assign n6139 = ~\pi0846  & ~n1633 ;
  assign n6140 = n3746 & ~n6139 ;
  assign n6141 = ~\pi0095  & n3746 ;
  assign n6142 = n2686 & n6141 ;
  assign n6143 = ~n6140 & ~n6142 ;
  assign n6144 = \pi0228  & ~n6094 ;
  assign n6145 = ~\pi0216  & ~n6144 ;
  assign n6146 = n6093 & ~n6145 ;
  assign n6147 = n6143 & n6146 ;
  assign n6148 = \pi0222  & ~\pi0224  ;
  assign n6149 = n6102 & n6148 ;
  assign n6150 = ~\pi0224  & ~n6149 ;
  assign n6151 = ~n6139 & n6150 ;
  assign n6152 = ~\pi0095  & n6150 ;
  assign n6153 = n2686 & n6152 ;
  assign n6154 = ~n6151 & ~n6153 ;
  assign n6155 = \pi0224  & \pi0278  ;
  assign n6156 = ~\pi0222  & ~n6155 ;
  assign n6157 = ~n6149 & ~n6156 ;
  assign n6158 = n3058 & ~n6157 ;
  assign n6159 = n6154 & n6158 ;
  assign n6160 = ~\pi0039  & ~n6104 ;
  assign n6161 = ~n6159 & n6160 ;
  assign n6162 = ~n6147 & n6161 ;
  assign n6163 = ~n6138 & n6162 ;
  assign n6164 = ~\pi0039  & ~n2256 ;
  assign n6165 = ~n6159 & n6164 ;
  assign n6166 = ~\pi0228  & n2618 ;
  assign n6167 = ~\pi0228  & \pi0846  ;
  assign n6168 = ~n2615 & n6167 ;
  assign n6169 = ~n6166 & ~n6168 ;
  assign n6170 = \pi0228  & ~n6097 ;
  assign n6171 = ~n2651 & n6093 ;
  assign n6172 = ~n6170 & n6171 ;
  assign n6173 = n6169 & n6172 ;
  assign n6174 = ~\pi0278  & n2291 ;
  assign n6175 = \pi0299  & ~n6104 ;
  assign n6176 = ~n6174 & n6175 ;
  assign n6177 = ~n6173 & n6176 ;
  assign n6178 = ~\pi0224  & \pi0846  ;
  assign n6179 = ~n1633 & n6178 ;
  assign n6180 = n6156 & ~n6179 ;
  assign n6181 = n2194 & ~n6149 ;
  assign n6182 = ~n6180 & n6181 ;
  assign n6183 = ~\pi0299  & ~n3045 ;
  assign n6184 = n2194 & n6183 ;
  assign n6185 = ~n6182 & n6184 ;
  assign n6186 = ~\pi0299  & ~n6185 ;
  assign n6187 = n1288 & ~n6186 ;
  assign n6188 = ~n2259 & n6187 ;
  assign n6189 = ~n6177 & n6188 ;
  assign n6190 = ~\pi0299  & n6185 ;
  assign n6191 = ~\pi0215  & n6104 ;
  assign n6192 = ~\pi0215  & n6093 ;
  assign n6193 = ~n6114 & n6192 ;
  assign n6194 = ~n6191 & ~n6193 ;
  assign n6195 = \pi0299  & ~n2652 ;
  assign n6196 = ~n6194 & n6195 ;
  assign n6197 = ~n6190 & ~n6196 ;
  assign n6198 = ~n1288 & ~n6197 ;
  assign n6199 = \pi0100  & ~n6198 ;
  assign n6200 = ~n6189 & n6199 ;
  assign n6201 = \pi0215  & n2297 ;
  assign n6202 = n2297 & ~n6104 ;
  assign n6203 = ~n6101 & n6202 ;
  assign n6204 = ~n6201 & ~n6203 ;
  assign n6205 = \pi0039  & ~\pi0299  ;
  assign n6206 = ~n6185 & n6205 ;
  assign n6207 = ~\pi0038  & ~n6206 ;
  assign n6208 = n6204 & n6207 ;
  assign n6209 = ~n6200 & n6208 ;
  assign n6210 = ~n6165 & n6209 ;
  assign n6211 = ~n6163 & n6210 ;
  assign n6212 = ~n2652 & ~n6194 ;
  assign n6213 = \pi0299  & ~n6212 ;
  assign n6214 = \pi0038  & ~n6186 ;
  assign n6215 = ~n6213 & n6214 ;
  assign n6216 = ~\pi0100  & ~n6215 ;
  assign n6217 = \pi0075  & ~n6186 ;
  assign n6218 = ~n6213 & n6217 ;
  assign n6219 = n4539 & ~n6218 ;
  assign n6220 = n6216 & n6219 ;
  assign n6221 = n6199 & n6219 ;
  assign n6222 = ~n6189 & n6221 ;
  assign n6223 = ~n6220 & ~n6222 ;
  assign n6224 = ~n6211 & ~n6223 ;
  assign n6225 = ~n2328 & ~n6197 ;
  assign n6226 = \pi0087  & ~n6225 ;
  assign n6227 = ~\pi0075  & ~n6226 ;
  assign n6228 = ~n6101 & n6175 ;
  assign n6229 = ~n2259 & ~n6228 ;
  assign n6230 = n2328 & ~n6186 ;
  assign n6231 = ~\pi0075  & n6230 ;
  assign n6232 = n6229 & n6231 ;
  assign n6233 = ~n6227 & ~n6232 ;
  assign n6234 = ~\pi0092  & ~n6218 ;
  assign n6235 = n6233 & n6234 ;
  assign n6236 = ~n1291 & n3409 ;
  assign n6237 = \pi0055  & ~n6236 ;
  assign n6238 = \pi0055  & ~n6104 ;
  assign n6239 = ~n6115 & n6238 ;
  assign n6240 = ~n6237 & ~n6239 ;
  assign n6241 = ~\pi0056  & n6240 ;
  assign n6242 = ~\pi0215  & n3008 ;
  assign n6243 = ~n6105 & n6242 ;
  assign n6244 = ~n6241 & ~n6243 ;
  assign n6245 = \pi0092  & n6197 ;
  assign n6246 = ~n3089 & ~n6245 ;
  assign n6247 = n2387 & n6197 ;
  assign n6248 = n2511 & ~n6247 ;
  assign n6249 = n6246 & n6248 ;
  assign n6250 = n6230 & n6248 ;
  assign n6251 = n6229 & n6250 ;
  assign n6252 = ~n6249 & ~n6251 ;
  assign n6253 = ~n6244 & ~n6252 ;
  assign n6254 = ~n6235 & n6253 ;
  assign n6255 = ~n6224 & n6254 ;
  assign n6256 = ~n2511 & ~n6197 ;
  assign n6257 = ~\pi0055  & ~n6256 ;
  assign n6258 = ~n6244 & ~n6257 ;
  assign n6259 = n1292 & n6126 ;
  assign n6260 = ~\pi0215  & n3030 ;
  assign n6261 = ~n6105 & n6260 ;
  assign n6262 = ~n6104 & ~n6115 ;
  assign n6263 = ~n2407 & n3409 ;
  assign n6264 = ~n6262 & n6263 ;
  assign n6265 = ~\pi0062  & ~n6264 ;
  assign n6266 = n6126 & n6265 ;
  assign n6267 = ~n6261 & n6266 ;
  assign n6268 = ~n6259 & ~n6267 ;
  assign n6269 = ~n6258 & ~n6268 ;
  assign n6270 = ~n6255 & n6269 ;
  assign n6271 = ~n6128 & ~n6270 ;
  assign n6272 = ~\pi0242  & n6124 ;
  assign n6273 = \pi1134  & ~n6272 ;
  assign n6274 = \pi0152  & ~\pi0846  ;
  assign n6275 = ~\pi0228  & ~n6274 ;
  assign n6276 = ~n4492 & ~n6275 ;
  assign n6277 = n6143 & ~n6145 ;
  assign n6278 = n1633 & n6144 ;
  assign n6279 = ~\pi0095  & n6144 ;
  assign n6280 = n2686 & n6279 ;
  assign n6281 = ~n6278 & ~n6280 ;
  assign n6282 = ~n6104 & n6281 ;
  assign n6283 = ~n6277 & n6282 ;
  assign n6284 = n6276 & n6283 ;
  assign n6285 = ~\pi0152  & ~n5688 ;
  assign n6286 = \pi0152  & ~n2718 ;
  assign n6287 = \pi0846  & ~n6286 ;
  assign n6288 = n6283 & n6287 ;
  assign n6289 = ~n6285 & n6288 ;
  assign n6290 = ~n6284 & ~n6289 ;
  assign n6291 = n6093 & ~n6098 ;
  assign n6292 = ~n6091 & n6291 ;
  assign n6293 = n6202 & ~n6292 ;
  assign n6294 = ~n6201 & ~n6293 ;
  assign n6295 = n2199 & ~n6155 ;
  assign n6296 = ~n6179 & n6295 ;
  assign n6297 = ~\pi0299  & ~n6296 ;
  assign n6298 = \pi0039  & n6297 ;
  assign n6299 = ~n6185 & n6298 ;
  assign n6300 = ~\pi0038  & ~n6299 ;
  assign n6301 = n6294 & n6300 ;
  assign n6302 = ~n6093 & ~n6104 ;
  assign n6303 = n2256 & ~n6302 ;
  assign n6304 = n6301 & n6303 ;
  assign n6305 = n6290 & n6304 ;
  assign n6306 = n3058 & n6156 ;
  assign n6307 = ~n6179 & n6306 ;
  assign n6308 = ~\pi0095  & n6306 ;
  assign n6309 = n2686 & n6308 ;
  assign n6310 = ~n6307 & ~n6309 ;
  assign n6311 = ~\pi0039  & n6310 ;
  assign n6312 = ~n6159 & n6311 ;
  assign n6313 = n6300 & ~n6312 ;
  assign n6314 = n6294 & n6313 ;
  assign n6315 = \pi0299  & n6194 ;
  assign n6316 = ~n6185 & n6297 ;
  assign n6317 = \pi0038  & ~n6316 ;
  assign n6318 = ~n6315 & n6317 ;
  assign n6319 = ~\pi0100  & ~n6318 ;
  assign n6320 = ~\pi0087  & n6319 ;
  assign n6321 = ~n6314 & n6320 ;
  assign n6322 = ~n6305 & n6321 ;
  assign n6323 = n6175 & ~n6292 ;
  assign n6324 = ~n2259 & ~n6323 ;
  assign n6325 = n2328 & ~n6316 ;
  assign n6326 = n6324 & n6325 ;
  assign n6327 = ~n2328 & ~n6316 ;
  assign n6328 = ~n6315 & n6327 ;
  assign n6329 = \pi0087  & ~n6328 ;
  assign n6330 = ~n6326 & n6329 ;
  assign n6331 = ~\pi0075  & ~n6330 ;
  assign n6332 = ~n1286 & ~n6316 ;
  assign n6333 = ~n6315 & n6332 ;
  assign n6334 = \pi0092  & ~n6333 ;
  assign n6335 = ~n6328 & n6334 ;
  assign n6336 = ~n6326 & n6335 ;
  assign n6337 = n2387 & n6316 ;
  assign n6338 = n2387 & n6315 ;
  assign n6339 = ~n6337 & ~n6338 ;
  assign n6340 = n2511 & n6339 ;
  assign n6341 = ~n6336 & n6340 ;
  assign n6342 = n6093 & ~n6170 ;
  assign n6343 = n6169 & n6342 ;
  assign n6344 = n6176 & ~n6343 ;
  assign n6345 = n1288 & ~n2259 ;
  assign n6346 = ~n6316 & n6345 ;
  assign n6347 = ~n6344 & n6346 ;
  assign n6348 = ~n1288 & ~n6316 ;
  assign n6349 = ~n6315 & n6348 ;
  assign n6350 = \pi0100  & ~n6349 ;
  assign n6351 = ~\pi0087  & n6350 ;
  assign n6352 = ~n6347 & n6351 ;
  assign n6353 = n6341 & ~n6352 ;
  assign n6354 = n6331 & n6353 ;
  assign n6355 = ~n6322 & n6354 ;
  assign n6356 = \pi0075  & ~n6316 ;
  assign n6357 = ~n6315 & n6356 ;
  assign n6358 = ~\pi0092  & ~n6357 ;
  assign n6359 = n6340 & ~n6358 ;
  assign n6360 = ~n6336 & n6359 ;
  assign n6361 = ~n6104 & ~n6292 ;
  assign n6362 = ~\pi0215  & n2406 ;
  assign n6363 = ~n6361 & n6362 ;
  assign n6364 = ~\pi0215  & ~n2407 ;
  assign n6365 = \pi0056  & n6104 ;
  assign n6366 = \pi0056  & n6093 ;
  assign n6367 = ~n6114 & n6366 ;
  assign n6368 = ~n6365 & ~n6367 ;
  assign n6369 = n6364 & ~n6368 ;
  assign n6370 = ~\pi0062  & ~n6369 ;
  assign n6371 = ~n2511 & ~n6316 ;
  assign n6372 = ~n6315 & n6371 ;
  assign n6373 = n6370 & ~n6372 ;
  assign n6374 = ~n6363 & n6373 ;
  assign n6375 = ~\pi0055  & n6374 ;
  assign n6376 = ~n6360 & n6375 ;
  assign n6377 = ~n6355 & n6376 ;
  assign n6378 = ~\pi0215  & ~n1291 ;
  assign n6379 = \pi0055  & ~n6378 ;
  assign n6380 = ~n6239 & ~n6379 ;
  assign n6381 = ~\pi0056  & n6380 ;
  assign n6382 = n6242 & ~n6361 ;
  assign n6383 = ~n6381 & ~n6382 ;
  assign n6384 = ~n6363 & n6370 ;
  assign n6385 = n6383 & n6384 ;
  assign n6386 = ~\pi0215  & n2454 ;
  assign n6387 = ~n6361 & n6386 ;
  assign n6388 = ~\pi0215  & ~n2504 ;
  assign n6389 = \pi0062  & ~n6388 ;
  assign n6390 = ~n6117 & ~n6389 ;
  assign n6391 = ~n6387 & ~n6390 ;
  assign n6392 = \pi1134  & ~n6391 ;
  assign n6393 = ~n6385 & n6392 ;
  assign n6394 = ~n6377 & n6393 ;
  assign n6395 = n2467 & n6394 ;
  assign n6396 = ~n6273 & ~n6395 ;
  assign n6397 = n6271 & ~n6396 ;
  assign n6398 = \pi1134  & ~n6397 ;
  assign n6399 = \pi0221  & ~n1220 ;
  assign n6400 = ~\pi0215  & ~n6399 ;
  assign n6401 = ~n6104 & n6400 ;
  assign n6402 = ~n2652 & ~n6401 ;
  assign n6403 = ~n2652 & n6093 ;
  assign n6404 = ~n6114 & n6403 ;
  assign n6405 = ~n6402 & ~n6404 ;
  assign n6406 = ~n2504 & n6405 ;
  assign n6407 = \pi0062  & ~n6406 ;
  assign n6408 = n2467 & ~n6407 ;
  assign n6409 = ~\pi0056  & ~n6104 ;
  assign n6410 = n6400 & n6409 ;
  assign n6411 = n2407 & n6410 ;
  assign n6412 = n2467 & n6411 ;
  assign n6413 = ~n6101 & n6412 ;
  assign n6414 = ~n6408 & ~n6413 ;
  assign n6415 = ~n2467 & n6405 ;
  assign n6416 = \pi0242  & ~n6415 ;
  assign n6417 = n6414 & n6416 ;
  assign n6418 = \pi0299  & ~n6405 ;
  assign n6419 = ~n6182 & n6183 ;
  assign n6420 = ~n2511 & ~n6419 ;
  assign n6421 = ~n6418 & n6420 ;
  assign n6422 = ~\pi0055  & ~n6421 ;
  assign n6423 = ~n1291 & n6405 ;
  assign n6424 = \pi0055  & ~n6423 ;
  assign n6425 = ~\pi0056  & ~n6424 ;
  assign n6426 = n1291 & n6401 ;
  assign n6427 = ~\pi0056  & n6426 ;
  assign n6428 = ~n6101 & n6427 ;
  assign n6429 = ~n6425 & ~n6428 ;
  assign n6430 = ~n6422 & ~n6429 ;
  assign n6431 = n2328 & ~n6183 ;
  assign n6432 = n2328 & ~n6180 ;
  assign n6433 = n6181 & n6432 ;
  assign n6434 = ~n6431 & ~n6433 ;
  assign n6435 = ~\pi0299  & ~n6434 ;
  assign n6436 = n6401 & ~n6434 ;
  assign n6437 = ~n6101 & n6436 ;
  assign n6438 = ~n6435 & ~n6437 ;
  assign n6439 = ~n2328 & ~n6419 ;
  assign n6440 = ~n6418 & n6439 ;
  assign n6441 = \pi0087  & ~n6440 ;
  assign n6442 = n6438 & n6441 ;
  assign n6443 = ~\pi0075  & ~n6442 ;
  assign n6444 = \pi0075  & ~n6183 ;
  assign n6445 = \pi0075  & ~n6180 ;
  assign n6446 = n6181 & n6445 ;
  assign n6447 = ~n6444 & ~n6446 ;
  assign n6448 = ~\pi0092  & n6447 ;
  assign n6449 = n2633 & ~n6405 ;
  assign n6450 = ~n6448 & ~n6449 ;
  assign n6451 = ~n6443 & ~n6450 ;
  assign n6452 = n2256 & ~n6399 ;
  assign n6453 = ~n6104 & n6452 ;
  assign n6454 = ~n6147 & n6453 ;
  assign n6455 = ~n6138 & n6454 ;
  assign n6456 = ~n2193 & n3058 ;
  assign n6457 = n6150 & n6456 ;
  assign n6458 = ~n6139 & n6457 ;
  assign n6459 = ~\pi0095  & n6457 ;
  assign n6460 = n2686 & n6459 ;
  assign n6461 = ~n6458 & ~n6460 ;
  assign n6462 = \pi0038  & ~n6183 ;
  assign n6463 = \pi0038  & ~n6180 ;
  assign n6464 = n6181 & n6463 ;
  assign n6465 = ~n6462 & ~n6464 ;
  assign n6466 = ~\pi0100  & n6465 ;
  assign n6467 = n2563 & ~n6405 ;
  assign n6468 = ~n6466 & ~n6467 ;
  assign n6469 = n6157 & n6456 ;
  assign n6470 = ~\pi0039  & ~n6469 ;
  assign n6471 = ~n6468 & n6470 ;
  assign n6472 = n6461 & n6471 ;
  assign n6473 = ~n6455 & n6472 ;
  assign n6474 = ~\pi0038  & ~n6183 ;
  assign n6475 = ~\pi0038  & ~n6180 ;
  assign n6476 = n6181 & n6475 ;
  assign n6477 = ~n6474 & ~n6476 ;
  assign n6478 = ~\pi0299  & ~n6477 ;
  assign n6479 = n6401 & ~n6477 ;
  assign n6480 = ~n6101 & n6479 ;
  assign n6481 = ~n6478 & ~n6480 ;
  assign n6482 = ~n1288 & ~n6468 ;
  assign n6483 = n6481 & n6482 ;
  assign n6484 = n1288 & ~n6183 ;
  assign n6485 = n1288 & ~n6180 ;
  assign n6486 = n6181 & n6485 ;
  assign n6487 = ~n6484 & ~n6486 ;
  assign n6488 = n6401 & ~n6487 ;
  assign n6489 = ~n6174 & n6488 ;
  assign n6490 = ~n6173 & n6489 ;
  assign n6491 = ~n1288 & ~n6419 ;
  assign n6492 = ~n6418 & n6491 ;
  assign n6493 = ~\pi0299  & ~n6487 ;
  assign n6494 = \pi0100  & ~n6493 ;
  assign n6495 = ~n6492 & n6494 ;
  assign n6496 = ~n6490 & n6495 ;
  assign n6497 = ~n6483 & ~n6496 ;
  assign n6498 = ~n6473 & n6497 ;
  assign n6499 = ~\pi0087  & ~n6450 ;
  assign n6500 = ~n6498 & n6499 ;
  assign n6501 = ~n6451 & ~n6500 ;
  assign n6502 = ~n1286 & ~n6183 ;
  assign n6503 = ~n1286 & ~n6180 ;
  assign n6504 = n6181 & n6503 ;
  assign n6505 = ~n6502 & ~n6504 ;
  assign n6506 = \pi0092  & n6505 ;
  assign n6507 = n3003 & ~n6405 ;
  assign n6508 = ~n6506 & ~n6507 ;
  assign n6509 = ~n6440 & ~n6508 ;
  assign n6510 = n6438 & n6509 ;
  assign n6511 = ~n1286 & ~n6508 ;
  assign n6512 = n2511 & ~n6511 ;
  assign n6513 = ~n6510 & n6512 ;
  assign n6514 = ~n6429 & n6513 ;
  assign n6515 = n6501 & n6514 ;
  assign n6516 = ~n6430 & ~n6515 ;
  assign n6517 = ~n2407 & n6405 ;
  assign n6518 = ~\pi0062  & ~n6517 ;
  assign n6519 = ~n1292 & ~n6518 ;
  assign n6520 = n2407 & n6401 ;
  assign n6521 = ~n1292 & n6520 ;
  assign n6522 = ~n6101 & n6521 ;
  assign n6523 = ~n6519 & ~n6522 ;
  assign n6524 = n6416 & n6523 ;
  assign n6525 = n6516 & n6524 ;
  assign n6526 = ~n6417 & ~n6525 ;
  assign n6527 = ~n3915 & ~n6433 ;
  assign n6528 = ~\pi0299  & ~n6527 ;
  assign n6529 = n6401 & ~n6527 ;
  assign n6530 = ~n6292 & n6529 ;
  assign n6531 = ~n6528 & ~n6530 ;
  assign n6532 = ~\pi0299  & ~n6182 ;
  assign n6533 = \pi0299  & ~n6401 ;
  assign n6534 = \pi0299  & n6093 ;
  assign n6535 = ~n6114 & n6534 ;
  assign n6536 = ~n6533 & ~n6535 ;
  assign n6537 = ~n6532 & n6536 ;
  assign n6538 = \pi0092  & ~n6537 ;
  assign n6539 = ~n3089 & ~n6538 ;
  assign n6540 = n6531 & ~n6539 ;
  assign n6541 = n2387 & ~n6537 ;
  assign n6542 = n2511 & ~n6541 ;
  assign n6543 = ~n6540 & n6542 ;
  assign n6544 = ~n2407 & n6401 ;
  assign n6545 = ~n6115 & n6544 ;
  assign n6546 = ~\pi0062  & ~n6545 ;
  assign n6547 = ~n1292 & ~n6546 ;
  assign n6548 = ~n6292 & n6521 ;
  assign n6549 = ~n6547 & ~n6548 ;
  assign n6550 = ~n2511 & n6537 ;
  assign n6551 = ~\pi0055  & ~n6550 ;
  assign n6552 = n6549 & n6551 ;
  assign n6553 = ~n6543 & n6552 ;
  assign n6554 = ~n6149 & n6178 ;
  assign n6555 = n6456 & n6554 ;
  assign n6556 = ~n1633 & n6555 ;
  assign n6557 = ~n2716 & n6556 ;
  assign n6558 = n6470 & ~n6557 ;
  assign n6559 = ~n3972 & ~n6476 ;
  assign n6560 = ~\pi0299  & ~n6559 ;
  assign n6561 = n6401 & ~n6559 ;
  assign n6562 = ~n6292 & n6561 ;
  assign n6563 = ~n6560 & ~n6562 ;
  assign n6564 = ~n1288 & n6563 ;
  assign n6565 = ~n6558 & ~n6564 ;
  assign n6566 = n6452 & ~n6564 ;
  assign n6567 = ~n3987 & ~n6464 ;
  assign n6568 = n6536 & ~n6567 ;
  assign n6569 = n2362 & ~n6568 ;
  assign n6570 = ~n6566 & n6569 ;
  assign n6571 = ~n6302 & n6569 ;
  assign n6572 = n6290 & n6571 ;
  assign n6573 = ~n6570 & ~n6572 ;
  assign n6574 = ~n6565 & ~n6573 ;
  assign n6575 = ~n4002 & ~n6486 ;
  assign n6576 = n6401 & ~n6575 ;
  assign n6577 = ~n6174 & n6576 ;
  assign n6578 = ~n6343 & n6577 ;
  assign n6579 = ~n1288 & n6537 ;
  assign n6580 = \pi0100  & ~n6579 ;
  assign n6581 = ~\pi0299  & n1288 ;
  assign n6582 = ~n6180 & n6581 ;
  assign n6583 = n6181 & n6582 ;
  assign n6584 = ~\pi0087  & ~n6583 ;
  assign n6585 = n6580 & n6584 ;
  assign n6586 = ~n6578 & n6585 ;
  assign n6587 = ~n2328 & n6537 ;
  assign n6588 = \pi0087  & ~n6587 ;
  assign n6589 = n6531 & n6588 ;
  assign n6590 = ~\pi0075  & ~n6589 ;
  assign n6591 = ~n6586 & n6590 ;
  assign n6592 = ~n6574 & n6591 ;
  assign n6593 = ~n4021 & ~n6446 ;
  assign n6594 = n6536 & ~n6593 ;
  assign n6595 = ~\pi0092  & ~n6594 ;
  assign n6596 = n6552 & n6595 ;
  assign n6597 = ~n6592 & n6596 ;
  assign n6598 = ~n6553 & ~n6597 ;
  assign n6599 = ~n1291 & n6401 ;
  assign n6600 = ~n6115 & n6599 ;
  assign n6601 = \pi0055  & ~n6600 ;
  assign n6602 = ~\pi0056  & ~n6601 ;
  assign n6603 = ~n6292 & n6427 ;
  assign n6604 = ~n6602 & ~n6603 ;
  assign n6605 = n6549 & n6604 ;
  assign n6606 = ~n6292 & n6411 ;
  assign n6607 = ~n2504 & n6401 ;
  assign n6608 = ~n6115 & n6607 ;
  assign n6609 = \pi0062  & ~n6608 ;
  assign n6610 = ~n6606 & n6609 ;
  assign n6611 = n2467 & ~n6610 ;
  assign n6612 = ~n6605 & n6611 ;
  assign n6613 = n6598 & n6612 ;
  assign n6614 = ~n2467 & n6401 ;
  assign n6615 = ~n6115 & n6614 ;
  assign n6616 = ~\pi0242  & ~n6615 ;
  assign n6617 = ~n6613 & n6616 ;
  assign n6618 = ~n6397 & ~n6617 ;
  assign n6619 = n6526 & n6618 ;
  assign n6620 = ~n6398 & ~n6619 ;
  assign n6621 = \pi0057  & \pi0059  ;
  assign n6622 = n1292 & ~n6621 ;
  assign n6623 = ~\pi0055  & \pi0057  ;
  assign n6624 = n6622 & n6623 ;
  assign n6625 = n1291 & n6624 ;
  assign n6626 = n1281 & n6625 ;
  assign n6627 = n1260 & n6626 ;
  assign n6628 = ~n2467 & ~n6627 ;
  assign n6629 = n2327 & n4520 ;
  assign n6630 = n1287 & n6629 ;
  assign n6631 = ~\pi0074  & n2423 ;
  assign n6632 = n6630 & n6631 ;
  assign n6633 = n1638 & n6632 ;
  assign n6634 = \pi0062  & ~n6627 ;
  assign n6635 = ~n6633 & n6634 ;
  assign n6636 = ~n6628 & ~n6635 ;
  assign n6637 = \pi0058  & n1256 ;
  assign n6638 = n1358 & n6637 ;
  assign n6639 = ~\pi0090  & ~n6638 ;
  assign n6640 = ~\pi0841  & n1277 ;
  assign n6641 = n1256 & n6640 ;
  assign n6642 = n1358 & n6641 ;
  assign n6643 = \pi0093  & ~n6642 ;
  assign n6644 = ~n1857 & ~n6643 ;
  assign n6645 = ~n6639 & n6644 ;
  assign n6646 = ~\pi0109  & n1319 ;
  assign n6647 = \pi0110  & ~n6646 ;
  assign n6648 = ~n1599 & ~n6647 ;
  assign n6649 = ~\pi0047  & ~n6648 ;
  assign n6650 = ~\pi0050  & n1276 ;
  assign n6651 = n1551 & n6650 ;
  assign n6652 = ~n1537 & n6651 ;
  assign n6653 = ~n1524 & n6652 ;
  assign n6654 = n1844 & ~n6653 ;
  assign n6655 = n1596 & ~n1847 ;
  assign n6656 = ~n6654 & n6655 ;
  assign n6657 = n1270 & ~n1587 ;
  assign n6658 = ~\pi0047  & n6657 ;
  assign n6659 = ~n6656 & n6658 ;
  assign n6660 = ~n6649 & ~n6659 ;
  assign n6661 = n1326 & ~n1392 ;
  assign n6662 = n6644 & n6661 ;
  assign n6663 = n6660 & n6662 ;
  assign n6664 = ~n6645 & ~n6663 ;
  assign n6665 = \pi0093  & n6642 ;
  assign n6666 = n1261 & ~n6665 ;
  assign n6667 = n6664 & n6666 ;
  assign n6668 = ~\pi0070  & n1354 ;
  assign n6669 = n1358 & n6668 ;
  assign n6670 = ~n1321 & ~n6669 ;
  assign n6671 = ~\pi0051  & n6670 ;
  assign n6672 = n1630 & ~n1868 ;
  assign n6673 = ~n6671 & n6672 ;
  assign n6674 = ~n6667 & n6673 ;
  assign n6675 = n1329 & n1962 ;
  assign n6676 = ~\pi0040  & \pi0072  ;
  assign n6677 = n1628 & n6676 ;
  assign n6678 = ~n6675 & ~n6677 ;
  assign n6679 = n1626 & n6678 ;
  assign n6680 = ~n6674 & n6679 ;
  assign n6681 = ~\pi0095  & n6680 ;
  assign n6682 = ~\pi0198  & ~\pi0299  ;
  assign n6683 = ~\pi0210  & \pi0299  ;
  assign n6684 = ~n6682 & ~n6683 ;
  assign n6685 = n2588 & n6684 ;
  assign n6686 = n1652 & ~n6684 ;
  assign n6687 = n1354 & n6686 ;
  assign n6688 = n1358 & n6687 ;
  assign n6689 = n1739 & ~n6688 ;
  assign n6690 = ~n6685 & n6689 ;
  assign n6691 = ~\pi0100  & n4520 ;
  assign n6692 = n1638 & n6691 ;
  assign n6693 = ~n2327 & ~n6692 ;
  assign n6694 = n2592 & ~n6693 ;
  assign n6695 = ~n6690 & n6694 ;
  assign n6696 = ~n6681 & n6695 ;
  assign n6697 = \pi0038  & ~n6693 ;
  assign n6698 = \pi0829  & \pi1091  ;
  assign n6699 = ~n1686 & n6698 ;
  assign n6700 = \pi0829  & ~\pi1093  ;
  assign n6701 = ~\pi0824  & ~n6700 ;
  assign n6702 = ~n6699 & n6701 ;
  assign n6703 = \pi1091  & \pi1093  ;
  assign n6704 = n1686 & n6703 ;
  assign n6705 = ~n6702 & ~n6704 ;
  assign n6706 = ~\pi0332  & ~\pi0468  ;
  assign n6707 = ~\pi0662  & \pi0680  ;
  assign n6708 = ~\pi0661  & ~\pi0681  ;
  assign n6709 = n6707 & n6708 ;
  assign n6710 = \pi0603  & ~\pi0642  ;
  assign n6711 = ~\pi0614  & ~\pi0616  ;
  assign n6712 = n6710 & n6711 ;
  assign n6713 = ~n6709 & ~n6712 ;
  assign n6714 = ~n6706 & ~n6713 ;
  assign n6715 = ~\pi0252  & ~\pi1001  ;
  assign n6716 = ~\pi0979  & ~n6715 ;
  assign n6717 = \pi0835  & \pi0984  ;
  assign n6718 = ~\pi0287  & ~n6717 ;
  assign n6719 = n6716 & n6718 ;
  assign n6720 = \pi0835  & \pi0950  ;
  assign n6721 = \pi1092  & n6720 ;
  assign n6722 = n6719 & n6721 ;
  assign n6723 = n6714 & n6722 ;
  assign n6724 = n6705 & n6723 ;
  assign n6725 = n2280 & ~n6724 ;
  assign n6726 = ~\pi0975  & ~\pi0978  ;
  assign n6727 = ~\pi0970  & ~\pi0972  ;
  assign n6728 = n6726 & n6727 ;
  assign n6729 = ~\pi0960  & ~\pi0963  ;
  assign n6730 = ~\pi0907  & ~\pi0947  ;
  assign n6731 = n6729 & n6730 ;
  assign n6732 = n6728 & n6731 ;
  assign n6733 = ~n6725 & n6732 ;
  assign n6734 = \pi0215  & n6732 ;
  assign n6735 = ~n6706 & ~n6712 ;
  assign n6736 = ~n6709 & n6735 ;
  assign n6737 = n6705 & ~n6736 ;
  assign n6738 = n6722 & n6737 ;
  assign n6739 = \pi0215  & ~n6738 ;
  assign n6740 = n2280 & n6739 ;
  assign n6741 = ~n6734 & ~n6740 ;
  assign n6742 = ~n6733 & ~n6741 ;
  assign n6743 = n6706 & ~n6732 ;
  assign n6744 = ~n6714 & ~n6743 ;
  assign n6745 = n6719 & n6720 ;
  assign n6746 = \pi0216  & \pi0221  ;
  assign n6747 = n1696 & n6746 ;
  assign n6748 = n6745 & n6747 ;
  assign n6749 = ~n6744 & n6748 ;
  assign n6750 = ~\pi0215  & n1281 ;
  assign n6751 = ~n6749 & n6750 ;
  assign n6752 = n1260 & n6751 ;
  assign n6753 = \pi0299  & ~n6752 ;
  assign n6754 = ~n6742 & n6753 ;
  assign n6755 = ~\pi0974  & ~\pi0977  ;
  assign n6756 = ~\pi0969  & ~\pi0971  ;
  assign n6757 = n6755 & n6756 ;
  assign n6758 = ~\pi0961  & ~\pi0967  ;
  assign n6759 = ~\pi0587  & ~\pi0602  ;
  assign n6760 = n6758 & n6759 ;
  assign n6761 = n6757 & n6760 ;
  assign n6762 = n2280 & ~n6738 ;
  assign n6763 = ~n6761 & ~n6762 ;
  assign n6764 = \pi0223  & ~n6761 ;
  assign n6765 = \pi0223  & ~n6724 ;
  assign n6766 = n2280 & n6765 ;
  assign n6767 = ~n6764 & ~n6766 ;
  assign n6768 = ~n6763 & ~n6767 ;
  assign n6769 = n6706 & ~n6761 ;
  assign n6770 = ~n6714 & ~n6769 ;
  assign n6771 = \pi0222  & \pi0224  ;
  assign n6772 = n1696 & n6771 ;
  assign n6773 = n6745 & n6772 ;
  assign n6774 = ~n6770 & n6773 ;
  assign n6775 = ~\pi0223  & n1281 ;
  assign n6776 = ~n6774 & n6775 ;
  assign n6777 = n1260 & n6776 ;
  assign n6778 = ~\pi0299  & ~n6777 ;
  assign n6779 = ~n6768 & n6778 ;
  assign n6780 = ~n6754 & ~n6779 ;
  assign n6781 = \pi0039  & ~n6693 ;
  assign n6782 = n6780 & n6781 ;
  assign n6783 = ~n6697 & ~n6782 ;
  assign n6784 = ~\pi0039  & n1261 ;
  assign n6785 = ~\pi0038  & \pi0100  ;
  assign n6786 = n6784 & n6785 ;
  assign n6787 = n1266 & n6786 ;
  assign n6788 = n1354 & n6787 ;
  assign n6789 = n1358 & n6788 ;
  assign n6790 = ~\pi0087  & ~n6789 ;
  assign n6791 = ~\pi0142  & ~\pi0299  ;
  assign n6792 = ~n2167 & n6791 ;
  assign n6793 = ~\pi0146  & \pi0299  ;
  assign n6794 = ~n1801 & n6793 ;
  assign n6795 = ~n6792 & ~n6794 ;
  assign n6796 = ~\pi0252  & n6795 ;
  assign n6797 = n1281 & n6796 ;
  assign n6798 = n1260 & n6797 ;
  assign n6799 = ~\pi0113  & ~\pi0116  ;
  assign n6800 = ~\pi0052  & n6799 ;
  assign n6801 = ~\pi0042  & ~\pi0114  ;
  assign n6802 = ~\pi0043  & ~\pi0115  ;
  assign n6803 = n6801 & n6802 ;
  assign n6804 = n6800 & n6803 ;
  assign n6805 = ~\pi0041  & ~\pi0099  ;
  assign n6806 = ~\pi0044  & ~\pi0101  ;
  assign n6807 = n6805 & n6806 ;
  assign n6808 = n6804 & n6807 ;
  assign n6809 = \pi0950  & \pi1092  ;
  assign n6810 = ~\pi0824  & ~\pi0829  ;
  assign n6811 = n6809 & ~n6810 ;
  assign n6812 = \pi0129  & \pi0250  ;
  assign n6813 = ~\pi1093  & ~n6812 ;
  assign n6814 = n6811 & n6813 ;
  assign n6815 = ~\pi0129  & \pi0250  ;
  assign n6816 = \pi0683  & ~n6815 ;
  assign n6817 = ~n6814 & n6816 ;
  assign n6818 = ~n6808 & n6817 ;
  assign n6819 = ~n6795 & ~n6818 ;
  assign n6820 = ~\pi0087  & ~n6819 ;
  assign n6821 = ~n6798 & n6820 ;
  assign n6822 = ~n6790 & ~n6821 ;
  assign n6823 = ~\pi0074  & ~n6822 ;
  assign n6824 = n6783 & n6823 ;
  assign n6825 = ~n6696 & n6824 ;
  assign n6826 = ~\pi0075  & n1285 ;
  assign n6827 = ~\pi0087  & n6826 ;
  assign n6828 = n6629 & n6826 ;
  assign n6829 = n1638 & n6828 ;
  assign n6830 = ~n6827 & ~n6829 ;
  assign n6831 = ~\pi0074  & n6830 ;
  assign n6832 = n2404 & n6630 ;
  assign n6833 = n1638 & n6832 ;
  assign n6834 = \pi0056  & ~n6833 ;
  assign n6835 = ~\pi0055  & n6630 ;
  assign n6836 = n1638 & n6835 ;
  assign n6837 = ~n2404 & ~n6836 ;
  assign n6838 = ~n6834 & ~n6837 ;
  assign n6839 = ~n6831 & n6838 ;
  assign n6840 = ~n6825 & n6839 ;
  assign n6841 = n2405 & n6630 ;
  assign n6842 = n1638 & n6841 ;
  assign n6843 = ~\pi0062  & ~n6627 ;
  assign n6844 = ~n6842 & n6843 ;
  assign n6845 = ~n6840 & n6844 ;
  assign n6846 = n6636 & ~n6845 ;
  assign n6847 = ~\pi0055  & ~\pi0059  ;
  assign n6848 = n1292 & n6847 ;
  assign n6849 = ~\pi0228  & ~n6848 ;
  assign n6850 = \pi0057  & ~n6849 ;
  assign n6851 = ~n6706 & ~n6709 ;
  assign n6852 = ~\pi0907  & n6706 ;
  assign n6853 = \pi0030  & \pi0228  ;
  assign n6854 = ~n6852 & n6853 ;
  assign n6855 = ~n6851 & n6854 ;
  assign n6856 = n6850 & n6855 ;
  assign n6857 = ~\pi0228  & n1288 ;
  assign n6858 = n1281 & n6857 ;
  assign n6859 = n1260 & n6858 ;
  assign n6860 = ~n6851 & ~n6852 ;
  assign n6861 = n1287 & n1289 ;
  assign n6862 = n6860 & n6861 ;
  assign n6863 = n6850 & n6862 ;
  assign n6864 = n6859 & n6863 ;
  assign n6865 = ~n6856 & ~n6864 ;
  assign n6866 = ~\pi0057  & \pi0228  ;
  assign n6867 = ~\pi0055  & ~\pi0057  ;
  assign n6868 = n1292 & n6867 ;
  assign n6869 = ~n6866 & ~n6868 ;
  assign n6870 = n6855 & ~n6869 ;
  assign n6871 = n6862 & ~n6869 ;
  assign n6872 = n6859 & n6871 ;
  assign n6873 = ~n6870 & ~n6872 ;
  assign n6874 = ~n2467 & n6873 ;
  assign n6875 = n6865 & n6874 ;
  assign n6876 = n6859 & n6862 ;
  assign n6877 = \pi0055  & ~n6855 ;
  assign n6878 = ~n6876 & n6877 ;
  assign n6879 = n1292 & ~n6878 ;
  assign n6880 = ~n1292 & n6853 ;
  assign n6881 = ~n6852 & n6880 ;
  assign n6882 = ~n6851 & n6881 ;
  assign n6883 = ~\pi0059  & ~n6882 ;
  assign n6884 = n6865 & n6883 ;
  assign n6885 = ~n6879 & n6884 ;
  assign n6886 = \pi0299  & ~n6852 ;
  assign n6887 = ~n6851 & n6886 ;
  assign n6888 = ~\pi0602  & n6706 ;
  assign n6889 = ~\pi0299  & ~n6888 ;
  assign n6890 = ~n6851 & n6889 ;
  assign n6891 = ~n6887 & ~n6890 ;
  assign n6892 = ~n2342 & n6853 ;
  assign n6893 = ~n6891 & n6892 ;
  assign n6894 = ~\pi0075  & ~n6893 ;
  assign n6895 = ~\pi0075  & \pi0092  ;
  assign n6896 = \pi0092  & n6853 ;
  assign n6897 = ~n6891 & n6896 ;
  assign n6898 = ~n6895 & ~n6897 ;
  assign n6899 = ~n6894 & ~n6898 ;
  assign n6900 = ~n3421 & ~n6853 ;
  assign n6901 = n1288 & n2362 ;
  assign n6902 = ~n6891 & n6901 ;
  assign n6903 = ~n6898 & n6902 ;
  assign n6904 = ~n6900 & n6903 ;
  assign n6905 = ~n6899 & ~n6904 ;
  assign n6906 = ~\pi0054  & n6905 ;
  assign n6907 = ~n6900 & n6902 ;
  assign n6908 = ~\pi0092  & n6894 ;
  assign n6909 = ~n6907 & n6908 ;
  assign n6910 = ~\pi0074  & n2364 ;
  assign n6911 = ~\pi0074  & n6853 ;
  assign n6912 = ~n6891 & n6911 ;
  assign n6913 = ~n6910 & ~n6912 ;
  assign n6914 = ~n6909 & ~n6913 ;
  assign n6915 = ~n2511 & ~n6914 ;
  assign n6916 = ~n6906 & ~n6915 ;
  assign n6917 = \pi0835  & ~\pi0984  ;
  assign n6918 = ~\pi0287  & n6917 ;
  assign n6919 = n6716 & n6918 ;
  assign n6920 = n1281 & n6919 ;
  assign n6921 = n1260 & n6920 ;
  assign n6922 = \pi0824  & \pi1093  ;
  assign n6923 = n6809 & n6922 ;
  assign n6924 = \pi1091  & n1686 ;
  assign n6925 = n6923 & ~n6924 ;
  assign n6926 = \pi1091  & n1689 ;
  assign n6927 = n1688 & n6926 ;
  assign n6928 = ~n6925 & ~n6927 ;
  assign n6929 = \pi0216  & n6928 ;
  assign n6930 = ~\pi0829  & ~n1686 ;
  assign n6931 = \pi1091  & ~n6930 ;
  assign n6932 = n6923 & ~n6931 ;
  assign n6933 = ~\pi0216  & ~n6932 ;
  assign n6934 = ~n6929 & ~n6933 ;
  assign n6935 = n6921 & n6934 ;
  assign n6936 = ~\pi0215  & \pi0221  ;
  assign n6937 = ~n6852 & n6936 ;
  assign n6938 = ~n6851 & n6937 ;
  assign n6939 = ~\pi0228  & n6938 ;
  assign n6940 = n6935 & n6939 ;
  assign n6941 = ~n6855 & ~n6940 ;
  assign n6942 = n2297 & ~n6941 ;
  assign n6943 = n6853 & ~n6888 ;
  assign n6944 = ~n6851 & n6943 ;
  assign n6945 = n6205 & n6944 ;
  assign n6946 = n1259 & n6932 ;
  assign n6947 = n1249 & n6946 ;
  assign n6948 = n6920 & n6947 ;
  assign n6949 = \pi0222  & ~\pi0223  ;
  assign n6950 = ~\pi0224  & n6949 ;
  assign n6951 = n6948 & n6950 ;
  assign n6952 = n1259 & ~n6928 ;
  assign n6953 = n1249 & n6952 ;
  assign n6954 = n6920 & n6953 ;
  assign n6955 = \pi0224  & n6949 ;
  assign n6956 = n6954 & n6955 ;
  assign n6957 = ~n6951 & ~n6956 ;
  assign n6958 = ~\pi0228  & ~n6888 ;
  assign n6959 = ~n6851 & n6958 ;
  assign n6960 = n6205 & n6959 ;
  assign n6961 = ~n6957 & n6960 ;
  assign n6962 = ~n6945 & ~n6961 ;
  assign n6963 = ~\pi0038  & n6962 ;
  assign n6964 = ~n6942 & n6963 ;
  assign n6965 = \pi0039  & n6964 ;
  assign n6966 = ~\pi0030  & \pi0228  ;
  assign n6967 = ~\pi0051  & n1321 ;
  assign n6968 = n1354 & n6967 ;
  assign n6969 = ~\pi0040  & ~\pi0841  ;
  assign n6970 = n1262 & n6969 ;
  assign n6971 = \pi0032  & ~\pi0198  ;
  assign n6972 = ~\pi0095  & n6971 ;
  assign n6973 = n6970 & n6972 ;
  assign n6974 = n6968 & n6973 ;
  assign n6975 = n1358 & n6974 ;
  assign n6976 = ~n6853 & ~n6975 ;
  assign n6977 = ~n6966 & ~n6976 ;
  assign n6978 = n1354 & n1981 ;
  assign n6979 = n1358 & n6978 ;
  assign n6980 = ~\pi0072  & ~n6979 ;
  assign n6981 = ~n1911 & n6980 ;
  assign n6982 = ~\pi0036  & \pi0067  ;
  assign n6983 = n1231 & n6982 ;
  assign n6984 = n1235 & n6983 ;
  assign n6985 = n1471 & n6984 ;
  assign n6986 = n1423 & ~n1424 ;
  assign n6987 = ~n6985 & n6986 ;
  assign n6988 = ~\pi0064  & ~\pi0065  ;
  assign n6989 = n1256 & n6988 ;
  assign n6990 = ~\pi0071  & n6989 ;
  assign n6991 = n1236 & n6989 ;
  assign n6992 = n1248 & n6991 ;
  assign n6993 = ~n6990 & ~n6992 ;
  assign n6994 = ~n1479 & ~n6993 ;
  assign n6995 = n1483 & n6994 ;
  assign n6996 = ~n6987 & n6995 ;
  assign n6997 = \pi0071  & ~n1249 ;
  assign n6998 = n1490 & n6989 ;
  assign n6999 = ~n6997 & n6998 ;
  assign n7000 = \pi0071  & n6989 ;
  assign n7001 = n1236 & n7000 ;
  assign n7002 = n1248 & n7001 ;
  assign n7003 = ~\pi0081  & ~n7002 ;
  assign n7004 = ~n6999 & n7003 ;
  assign n7005 = ~n6996 & n7004 ;
  assign n7006 = ~n1234 & n1243 ;
  assign n7007 = ~n1452 & n7006 ;
  assign n7008 = n1242 & n7007 ;
  assign n7009 = \pi0085  & ~n1456 ;
  assign n7010 = ~n7008 & ~n7009 ;
  assign n7011 = ~n1449 & ~n7008 ;
  assign n7012 = ~n1448 & n7011 ;
  assign n7013 = ~n7010 & ~n7012 ;
  assign n7014 = n1233 & ~n7013 ;
  assign n7015 = ~n1418 & ~n1460 ;
  assign n7016 = n1231 & n7015 ;
  assign n7017 = ~n7014 & n7016 ;
  assign n7018 = n1423 & ~n6985 ;
  assign n7019 = ~n1422 & n7018 ;
  assign n7020 = n7004 & n7019 ;
  assign n7021 = ~n7017 & n7020 ;
  assign n7022 = ~n7005 & ~n7021 ;
  assign n7023 = ~\pi0077  & ~\pi0102  ;
  assign n7024 = n1253 & n7023 ;
  assign n7025 = ~n1529 & n7024 ;
  assign n7026 = n1542 & n1543 ;
  assign n7027 = \pi0050  & ~n7026 ;
  assign n7028 = ~\pi0060  & ~n7027 ;
  assign n7029 = n7025 & n7028 ;
  assign n7030 = n7022 & n7029 ;
  assign n7031 = n1562 & ~n7030 ;
  assign n7032 = n1325 & ~n1599 ;
  assign n7033 = ~\pi0094  & ~\pi0108  ;
  assign n7034 = n1268 & n7033 ;
  assign n7035 = ~\pi0086  & n7034 ;
  assign n7036 = n1568 & n7034 ;
  assign n7037 = n1542 & n7036 ;
  assign n7038 = ~n7035 & ~n7037 ;
  assign n7039 = n7032 & ~n7038 ;
  assign n7040 = ~n1566 & n7039 ;
  assign n7041 = ~n7031 & n7040 ;
  assign n7042 = ~\pi0091  & ~\pi0314  ;
  assign n7043 = ~n1597 & n7032 ;
  assign n7044 = n7042 & ~n7043 ;
  assign n7045 = ~n7041 & n7044 ;
  assign n7046 = n1320 & n7045 ;
  assign n7047 = ~n6996 & ~n7002 ;
  assign n7048 = ~n7002 & n7019 ;
  assign n7049 = ~n7017 & n7048 ;
  assign n7050 = ~n7047 & ~n7049 ;
  assign n7051 = ~\pi0050  & ~\pi0081  ;
  assign n7052 = ~n1556 & n7051 ;
  assign n7053 = ~n7050 & n7052 ;
  assign n7054 = n1557 & ~n7025 ;
  assign n7055 = \pi0053  & ~n1564 ;
  assign n7056 = ~n1546 & ~n7055 ;
  assign n7057 = ~n7054 & n7056 ;
  assign n7058 = ~n7053 & n7057 ;
  assign n7059 = ~\pi0053  & n1347 ;
  assign n7060 = n1249 & n7059 ;
  assign n7061 = \pi0053  & n1340 ;
  assign n7062 = n1249 & n7061 ;
  assign n7063 = ~n7060 & ~n7062 ;
  assign n7064 = ~\pi0086  & ~\pi0109  ;
  assign n7065 = ~n1587 & n7064 ;
  assign n7066 = n7063 & n7065 ;
  assign n7067 = ~n7058 & n7066 ;
  assign n7068 = n1319 & n1717 ;
  assign n7069 = \pi0091  & ~n7068 ;
  assign n7070 = ~\pi0058  & ~n7069 ;
  assign n7071 = n1597 & n7038 ;
  assign n7072 = n7032 & ~n7071 ;
  assign n7073 = n7070 & n7072 ;
  assign n7074 = ~n7067 & n7073 ;
  assign n7075 = ~\pi0091  & \pi0314  ;
  assign n7076 = ~\pi0058  & ~n7075 ;
  assign n7077 = ~n7069 & n7076 ;
  assign n7078 = n1320 & ~n7077 ;
  assign n7079 = ~n7074 & n7078 ;
  assign n7080 = ~n7046 & ~n7079 ;
  assign n7081 = \pi0090  & ~\pi0093  ;
  assign n7082 = ~n1856 & n7081 ;
  assign n7083 = ~\pi0035  & ~\pi0093  ;
  assign n7084 = ~\pi0035  & \pi0841  ;
  assign n7085 = n1829 & n7084 ;
  assign n7086 = n1358 & n7085 ;
  assign n7087 = ~n7083 & ~n7086 ;
  assign n7088 = ~n7082 & ~n7087 ;
  assign n7089 = n7080 & n7088 ;
  assign n7090 = ~\pi0070  & n6980 ;
  assign n7091 = ~n7089 & n7090 ;
  assign n7092 = ~n6981 & ~n7091 ;
  assign n7093 = ~n1629 & n2575 ;
  assign n7094 = ~n6979 & ~n7093 ;
  assign n7095 = ~n6966 & ~n7094 ;
  assign n7096 = n7092 & n7095 ;
  assign n7097 = ~n6977 & ~n7096 ;
  assign n7098 = \pi0181  & \pi0182  ;
  assign n7099 = \pi0145  & \pi0180  ;
  assign n7100 = n7098 & n7099 ;
  assign n7101 = ~n6888 & ~n7100 ;
  assign n7102 = ~n6851 & n7101 ;
  assign n7103 = ~n7097 & n7102 ;
  assign n7104 = ~\pi0299  & ~n7103 ;
  assign n7105 = ~\pi0228  & ~n6706 ;
  assign n7106 = n6709 & n7105 ;
  assign n7107 = n6975 & n7106 ;
  assign n7108 = ~n7094 & n7106 ;
  assign n7109 = n7092 & n7108 ;
  assign n7110 = ~n7107 & ~n7109 ;
  assign n7111 = ~\pi0228  & \pi0602  ;
  assign n7112 = n6706 & n7111 ;
  assign n7113 = n6975 & n7112 ;
  assign n7114 = ~\pi0047  & n1270 ;
  assign n7115 = ~n7038 & n7114 ;
  assign n7116 = ~n1566 & n7115 ;
  assign n7117 = ~n7031 & n7116 ;
  assign n7118 = ~\pi0097  & n7114 ;
  assign n7119 = n1586 & n7118 ;
  assign n7120 = n7042 & ~n7119 ;
  assign n7121 = ~n7117 & n7120 ;
  assign n7122 = n1320 & n7121 ;
  assign n7123 = ~\pi0086  & ~n1587 ;
  assign n7124 = n7063 & n7123 ;
  assign n7125 = ~n7058 & n7124 ;
  assign n7126 = ~n1587 & n7038 ;
  assign n7127 = n7114 & ~n7126 ;
  assign n7128 = n7070 & n7127 ;
  assign n7129 = ~n7125 & n7128 ;
  assign n7130 = n7078 & ~n7129 ;
  assign n7131 = ~n7122 & ~n7130 ;
  assign n7132 = n1911 & ~n7087 ;
  assign n7133 = ~n7082 & n7132 ;
  assign n7134 = n7131 & n7133 ;
  assign n7135 = \pi0070  & n1323 ;
  assign n7136 = n1378 & n7135 ;
  assign n7137 = n6980 & ~n7136 ;
  assign n7138 = ~n7134 & n7137 ;
  assign n7139 = ~n7094 & n7112 ;
  assign n7140 = ~n7138 & n7139 ;
  assign n7141 = ~n7113 & ~n7140 ;
  assign n7142 = ~n6944 & n7141 ;
  assign n7143 = n7110 & n7142 ;
  assign n7144 = n7100 & ~n7143 ;
  assign n7145 = n7104 & ~n7144 ;
  assign n7146 = n7092 & ~n7094 ;
  assign n7147 = \pi0032  & ~\pi0210  ;
  assign n7148 = ~\pi0095  & n7147 ;
  assign n7149 = n6970 & n7148 ;
  assign n7150 = n6968 & n7149 ;
  assign n7151 = n1358 & n7150 ;
  assign n7152 = ~n7146 & ~n7151 ;
  assign n7153 = ~n6706 & n6709 ;
  assign n7154 = ~n7152 & n7153 ;
  assign n7155 = ~n7094 & ~n7138 ;
  assign n7156 = ~n7151 & ~n7155 ;
  assign n7157 = \pi0907  & n6706 ;
  assign n7158 = ~n7156 & n7157 ;
  assign n7159 = \pi0299  & ~n6855 ;
  assign n7160 = \pi0158  & \pi0159  ;
  assign n7161 = \pi0160  & \pi0197  ;
  assign n7162 = n7160 & n7161 ;
  assign n7163 = n7159 & n7162 ;
  assign n7164 = ~n7158 & n7163 ;
  assign n7165 = ~n7154 & n7164 ;
  assign n7166 = \pi0232  & ~n7159 ;
  assign n7167 = ~n7151 & ~n7162 ;
  assign n7168 = ~n7146 & n7167 ;
  assign n7169 = ~\pi0228  & n7162 ;
  assign n7170 = ~\pi0228  & ~n6852 ;
  assign n7171 = ~n6851 & n7170 ;
  assign n7172 = ~n7169 & ~n7171 ;
  assign n7173 = \pi0232  & ~n7172 ;
  assign n7174 = ~n7168 & n7173 ;
  assign n7175 = ~n7166 & ~n7174 ;
  assign n7176 = ~n7165 & ~n7175 ;
  assign n7177 = ~n7145 & n7176 ;
  assign n7178 = ~n6851 & ~n6888 ;
  assign n7179 = ~n7097 & n7178 ;
  assign n7180 = ~\pi0299  & ~n7179 ;
  assign n7181 = n7151 & n7171 ;
  assign n7182 = ~n7094 & n7171 ;
  assign n7183 = n7092 & n7182 ;
  assign n7184 = ~n7181 & ~n7183 ;
  assign n7185 = n7159 & n7184 ;
  assign n7186 = ~\pi0232  & ~n7185 ;
  assign n7187 = ~n7180 & n7186 ;
  assign n7188 = n6964 & ~n7187 ;
  assign n7189 = ~n7177 & n7188 ;
  assign n7190 = ~n6965 & ~n7189 ;
  assign n7191 = ~n1288 & n6853 ;
  assign n7192 = ~\pi0087  & n7191 ;
  assign n7193 = ~n6891 & n7192 ;
  assign n7194 = ~n2362 & ~n7193 ;
  assign n7195 = ~\pi0039  & ~n6891 ;
  assign n7196 = ~n6900 & n7195 ;
  assign n7197 = n6853 & ~n6891 ;
  assign n7198 = \pi0038  & ~n7197 ;
  assign n7199 = ~n7196 & n7198 ;
  assign n7200 = ~n7194 & ~n7199 ;
  assign n7201 = n1288 & ~n7159 ;
  assign n7202 = ~\pi0095  & \pi0252  ;
  assign n7203 = n1634 & n7202 ;
  assign n7204 = n1618 & n7203 ;
  assign n7205 = ~\pi0035  & n1354 ;
  assign n7206 = n7204 & n7205 ;
  assign n7207 = n1358 & n7206 ;
  assign n7208 = n6709 & n7207 ;
  assign n7209 = \pi0252  & n6706 ;
  assign n7210 = n1281 & n7209 ;
  assign n7211 = n1259 & ~n6709 ;
  assign n7212 = n1249 & n7211 ;
  assign n7213 = n7210 & n7212 ;
  assign n7214 = ~n2070 & ~n7213 ;
  assign n7215 = ~n7208 & n7214 ;
  assign n7216 = n1281 & n6817 ;
  assign n7217 = n1260 & n7216 ;
  assign n7218 = ~n6808 & ~n6851 ;
  assign n7219 = n7217 & n7218 ;
  assign n7220 = n2070 & ~n7219 ;
  assign n7221 = ~n7215 & ~n7220 ;
  assign n7222 = n1288 & n7170 ;
  assign n7223 = n7221 & n7222 ;
  assign n7224 = ~n7201 & ~n7223 ;
  assign n7225 = \pi0142  & \pi0252  ;
  assign n7226 = ~\pi0189  & \pi0252  ;
  assign n7227 = n2166 & n7226 ;
  assign n7228 = ~n7225 & ~n7227 ;
  assign n7229 = n7213 & ~n7228 ;
  assign n7230 = n6709 & ~n7228 ;
  assign n7231 = n7207 & n7230 ;
  assign n7232 = ~n7229 & ~n7231 ;
  assign n7233 = ~\pi0299  & ~n6944 ;
  assign n7234 = ~\pi0142  & ~n2167 ;
  assign n7235 = ~n6851 & n7234 ;
  assign n7236 = ~n6808 & n7235 ;
  assign n7237 = n7217 & n7236 ;
  assign n7238 = n7233 & ~n7237 ;
  assign n7239 = n7232 & n7238 ;
  assign n7240 = ~\pi0299  & ~n6958 ;
  assign n7241 = ~n6944 & n7240 ;
  assign n7242 = ~\pi0087  & ~n7241 ;
  assign n7243 = ~n7239 & n7242 ;
  assign n7244 = ~n7199 & n7243 ;
  assign n7245 = ~n7224 & n7244 ;
  assign n7246 = ~n7200 & ~n7245 ;
  assign n7247 = n7190 & ~n7246 ;
  assign n7248 = \pi0100  & ~n7194 ;
  assign n7249 = \pi0100  & n7243 ;
  assign n7250 = ~n7224 & n7249 ;
  assign n7251 = ~n7248 & ~n7250 ;
  assign n7252 = \pi0087  & n6853 ;
  assign n7253 = ~n6891 & n7252 ;
  assign n7254 = ~\pi0075  & ~n7253 ;
  assign n7255 = n7251 & n7254 ;
  assign n7256 = ~n7247 & n7255 ;
  assign n7257 = \pi0075  & ~n6893 ;
  assign n7258 = ~\pi0092  & ~n7257 ;
  assign n7259 = ~\pi0092  & n6902 ;
  assign n7260 = ~n6900 & n7259 ;
  assign n7261 = ~n7258 & ~n7260 ;
  assign n7262 = ~n6915 & ~n7261 ;
  assign n7263 = ~n7256 & n7262 ;
  assign n7264 = ~n6916 & ~n7263 ;
  assign n7265 = ~\pi0054  & n2364 ;
  assign n7266 = ~n6893 & n7265 ;
  assign n7267 = n2364 & n2375 ;
  assign n7268 = \pi0074  & n6853 ;
  assign n7269 = ~n6891 & n7268 ;
  assign n7270 = ~n7267 & ~n7269 ;
  assign n7271 = ~n7266 & ~n7270 ;
  assign n7272 = n6902 & ~n7270 ;
  assign n7273 = ~n6900 & n7272 ;
  assign n7274 = ~n7271 & ~n7273 ;
  assign n7275 = ~\pi0055  & n7274 ;
  assign n7276 = n6884 & n7275 ;
  assign n7277 = n7264 & n7276 ;
  assign n7278 = ~n6885 & ~n7277 ;
  assign n7279 = ~n6875 & n7278 ;
  assign n7280 = ~\pi0947  & n6706 ;
  assign n7281 = n6853 & ~n7280 ;
  assign n7282 = ~n6735 & n7281 ;
  assign n7283 = n6850 & n7282 ;
  assign n7284 = ~n6735 & ~n7280 ;
  assign n7285 = n1259 & n7284 ;
  assign n7286 = n1249 & n7285 ;
  assign n7287 = n6858 & n7286 ;
  assign n7288 = n6850 & n6861 ;
  assign n7289 = n7287 & n7288 ;
  assign n7290 = ~n7283 & ~n7289 ;
  assign n7291 = ~n6869 & n7282 ;
  assign n7292 = n6861 & ~n6869 ;
  assign n7293 = n7287 & n7292 ;
  assign n7294 = ~n7291 & ~n7293 ;
  assign n7295 = ~n2467 & n7294 ;
  assign n7296 = n7290 & n7295 ;
  assign n7297 = n6880 & ~n7280 ;
  assign n7298 = ~n6735 & n7297 ;
  assign n7299 = ~\pi0059  & ~n7298 ;
  assign n7300 = n7290 & n7299 ;
  assign n7301 = ~n7296 & ~n7300 ;
  assign n7302 = ~n6706 & n6853 ;
  assign n7303 = n6712 & n7302 ;
  assign n7304 = \pi0299  & \pi0947  ;
  assign n7305 = ~\pi0299  & \pi0587  ;
  assign n7306 = ~n7304 & ~n7305 ;
  assign n7307 = n6706 & n6853 ;
  assign n7308 = ~n7306 & n7307 ;
  assign n7309 = ~n7303 & ~n7308 ;
  assign n7310 = ~n7265 & n7309 ;
  assign n7311 = \pi0074  & ~n7310 ;
  assign n7312 = ~\pi0055  & ~n7311 ;
  assign n7313 = ~n6706 & n6712 ;
  assign n7314 = n6706 & ~n7306 ;
  assign n7315 = ~n7313 & ~n7314 ;
  assign n7316 = n6901 & ~n7315 ;
  assign n7317 = ~n6900 & n7316 ;
  assign n7318 = ~n2342 & ~n7309 ;
  assign n7319 = n7265 & ~n7318 ;
  assign n7320 = ~\pi0055  & n7319 ;
  assign n7321 = ~n7317 & n7320 ;
  assign n7322 = ~n7312 & ~n7321 ;
  assign n7323 = ~\pi0075  & ~n7318 ;
  assign n7324 = ~\pi0092  & n7323 ;
  assign n7325 = ~n7317 & n7324 ;
  assign n7326 = ~n2364 & n7309 ;
  assign n7327 = ~\pi0074  & ~n7326 ;
  assign n7328 = ~n7325 & n7327 ;
  assign n7329 = ~n2511 & ~n7328 ;
  assign n7330 = ~n7322 & n7329 ;
  assign n7331 = \pi0075  & ~n7318 ;
  assign n7332 = ~n7317 & n7331 ;
  assign n7333 = ~\pi0092  & ~n7332 ;
  assign n7334 = \pi0087  & ~n7309 ;
  assign n7335 = ~\pi0075  & ~n7334 ;
  assign n7336 = n7333 & ~n7335 ;
  assign n7337 = ~\pi0039  & ~n7315 ;
  assign n7338 = ~n6900 & n7337 ;
  assign n7339 = \pi0038  & n7309 ;
  assign n7340 = ~n7338 & n7339 ;
  assign n7341 = ~\pi0100  & n7340 ;
  assign n7342 = ~\pi0587  & n6706 ;
  assign n7343 = ~n6735 & ~n7342 ;
  assign n7344 = ~n7097 & n7343 ;
  assign n7345 = ~\pi0299  & ~n7344 ;
  assign n7346 = \pi0299  & ~n7282 ;
  assign n7347 = ~\pi0228  & n7151 ;
  assign n7348 = ~\pi0228  & ~n7094 ;
  assign n7349 = n7092 & n7348 ;
  assign n7350 = ~n7347 & ~n7349 ;
  assign n7351 = n7284 & ~n7350 ;
  assign n7352 = n7346 & ~n7351 ;
  assign n7353 = ~\pi0232  & ~n7352 ;
  assign n7354 = ~n7345 & n7353 ;
  assign n7355 = ~\pi0039  & n7354 ;
  assign n7356 = n6853 & ~n7342 ;
  assign n7357 = ~n6735 & n7356 ;
  assign n7358 = ~\pi0228  & ~n7342 ;
  assign n7359 = ~n6735 & n7358 ;
  assign n7360 = n6975 & n7359 ;
  assign n7361 = ~n7094 & n7359 ;
  assign n7362 = ~n7138 & n7361 ;
  assign n7363 = ~n7360 & ~n7362 ;
  assign n7364 = n6706 & ~n7363 ;
  assign n7365 = n6712 & n7105 ;
  assign n7366 = n6975 & n7365 ;
  assign n7367 = ~n7094 & n7365 ;
  assign n7368 = n7092 & n7367 ;
  assign n7369 = ~n7366 & ~n7368 ;
  assign n7370 = ~n7364 & n7369 ;
  assign n7371 = ~n7357 & n7370 ;
  assign n7372 = n7100 & ~n7371 ;
  assign n7373 = ~n7100 & ~n7342 ;
  assign n7374 = ~n6735 & n7373 ;
  assign n7375 = ~n7097 & n7374 ;
  assign n7376 = ~\pi0299  & ~n7375 ;
  assign n7377 = ~n7372 & n7376 ;
  assign n7378 = n7151 & n7284 ;
  assign n7379 = ~n7094 & n7284 ;
  assign n7380 = ~n7138 & n7379 ;
  assign n7381 = ~n7378 & ~n7380 ;
  assign n7382 = n6706 & ~n7381 ;
  assign n7383 = n7151 & n7313 ;
  assign n7384 = ~n7094 & n7313 ;
  assign n7385 = n7092 & n7384 ;
  assign n7386 = ~n7383 & ~n7385 ;
  assign n7387 = ~n7382 & n7386 ;
  assign n7388 = n7162 & n7346 ;
  assign n7389 = n7387 & n7388 ;
  assign n7390 = \pi0232  & ~n7346 ;
  assign n7391 = ~\pi0228  & ~n7280 ;
  assign n7392 = ~n6735 & n7391 ;
  assign n7393 = ~n7169 & ~n7392 ;
  assign n7394 = \pi0232  & ~n7393 ;
  assign n7395 = ~n7168 & n7394 ;
  assign n7396 = ~n7390 & ~n7395 ;
  assign n7397 = ~n7389 & ~n7396 ;
  assign n7398 = ~\pi0039  & n7397 ;
  assign n7399 = ~n7377 & n7398 ;
  assign n7400 = ~n7355 & ~n7399 ;
  assign n7401 = ~\pi0299  & ~n7357 ;
  assign n7402 = \pi0039  & ~n7401 ;
  assign n7403 = \pi0039  & n7359 ;
  assign n7404 = ~n6957 & n7403 ;
  assign n7405 = ~n7402 & ~n7404 ;
  assign n7406 = ~\pi0038  & n7405 ;
  assign n7407 = n6853 & n7284 ;
  assign n7408 = ~\pi0228  & n7284 ;
  assign n7409 = n6935 & n7408 ;
  assign n7410 = ~n7407 & ~n7409 ;
  assign n7411 = n6936 & ~n7410 ;
  assign n7412 = \pi0299  & n6936 ;
  assign n7413 = ~n7346 & ~n7412 ;
  assign n7414 = ~\pi0038  & ~n7413 ;
  assign n7415 = ~n7411 & n7414 ;
  assign n7416 = ~n7406 & ~n7415 ;
  assign n7417 = ~\pi0100  & ~n7416 ;
  assign n7418 = n7400 & n7417 ;
  assign n7419 = ~n7341 & ~n7418 ;
  assign n7420 = ~\pi0228  & \pi0587  ;
  assign n7421 = ~n7365 & ~n7420 ;
  assign n7422 = n1260 & n7210 ;
  assign n7423 = \pi0142  & ~n6712 ;
  assign n7424 = ~n7422 & n7423 ;
  assign n7425 = \pi0142  & n6712 ;
  assign n7426 = ~n7207 & n7425 ;
  assign n7427 = ~n7424 & ~n7426 ;
  assign n7428 = ~n6735 & ~n6808 ;
  assign n7429 = n7217 & n7428 ;
  assign n7430 = ~\pi0142  & ~n7429 ;
  assign n7431 = n7427 & ~n7430 ;
  assign n7432 = ~n7421 & n7431 ;
  assign n7433 = ~\pi0189  & ~\pi0228  ;
  assign n7434 = n2166 & n7433 ;
  assign n7435 = ~\pi0299  & ~n7434 ;
  assign n7436 = ~n7357 & n7435 ;
  assign n7437 = ~n7432 & n7436 ;
  assign n7438 = ~n6712 & ~n7342 ;
  assign n7439 = n7422 & n7438 ;
  assign n7440 = n6712 & ~n7342 ;
  assign n7441 = n7207 & n7440 ;
  assign n7442 = ~n7439 & ~n7441 ;
  assign n7443 = ~\pi0299  & n7434 ;
  assign n7444 = n7442 & n7443 ;
  assign n7445 = ~\pi0947  & ~n7313 ;
  assign n7446 = ~n2070 & ~n7445 ;
  assign n7447 = ~n6712 & n7446 ;
  assign n7448 = n7422 & n7447 ;
  assign n7449 = n6712 & n7446 ;
  assign n7450 = n7207 & n7449 ;
  assign n7451 = ~n7448 & ~n7450 ;
  assign n7452 = ~n6808 & n7284 ;
  assign n7453 = n2070 & n7452 ;
  assign n7454 = n7217 & n7453 ;
  assign n7455 = n7346 & ~n7454 ;
  assign n7456 = n7451 & n7455 ;
  assign n7457 = \pi0228  & \pi0299  ;
  assign n7458 = ~n7282 & n7457 ;
  assign n7459 = n1288 & ~n7458 ;
  assign n7460 = ~n7456 & n7459 ;
  assign n7461 = ~n7444 & n7460 ;
  assign n7462 = ~n7437 & n7461 ;
  assign n7463 = ~n1288 & ~n7309 ;
  assign n7464 = \pi0100  & ~n7463 ;
  assign n7465 = ~n7462 & n7464 ;
  assign n7466 = ~\pi0087  & ~n7465 ;
  assign n7467 = n7333 & n7466 ;
  assign n7468 = n7419 & n7467 ;
  assign n7469 = ~n7336 & ~n7468 ;
  assign n7470 = \pi0075  & n7309 ;
  assign n7471 = \pi0092  & ~n7470 ;
  assign n7472 = ~\pi0054  & ~n7471 ;
  assign n7473 = ~\pi0054  & n7323 ;
  assign n7474 = ~n7317 & n7473 ;
  assign n7475 = ~n7472 & ~n7474 ;
  assign n7476 = ~n7322 & ~n7475 ;
  assign n7477 = n7469 & n7476 ;
  assign n7478 = ~n7330 & ~n7477 ;
  assign n7479 = n6861 & n7287 ;
  assign n7480 = \pi0055  & ~n7282 ;
  assign n7481 = ~n7479 & n7480 ;
  assign n7482 = n1292 & ~n7481 ;
  assign n7483 = ~n7296 & n7482 ;
  assign n7484 = n7478 & n7483 ;
  assign n7485 = ~n7301 & ~n7484 ;
  assign n7486 = \pi0970  & n7307 ;
  assign n7487 = \pi0059  & ~n7486 ;
  assign n7488 = ~\pi0228  & \pi0970  ;
  assign n7489 = n6706 & n7488 ;
  assign n7490 = n1259 & n7489 ;
  assign n7491 = n1249 & n7490 ;
  assign n7492 = n1281 & n1294 ;
  assign n7493 = n7491 & n7492 ;
  assign n7494 = n7487 & ~n7493 ;
  assign n7495 = ~\pi0057  & ~n7494 ;
  assign n7496 = \pi0970  & ~n1292 ;
  assign n7497 = n7307 & n7496 ;
  assign n7498 = ~\pi0059  & ~n7497 ;
  assign n7499 = n7495 & ~n7498 ;
  assign n7500 = \pi0299  & \pi0970  ;
  assign n7501 = ~\pi0299  & \pi0967  ;
  assign n7502 = ~n7500 & ~n7501 ;
  assign n7503 = n7307 & ~n7502 ;
  assign n7504 = ~n2364 & ~n7503 ;
  assign n7505 = ~\pi0074  & ~n7504 ;
  assign n7506 = ~n2511 & ~n7505 ;
  assign n7507 = \pi0967  & n6706 ;
  assign n7508 = ~\pi0299  & ~n7507 ;
  assign n7509 = ~\pi0299  & ~n6853 ;
  assign n7510 = ~n3421 & n7509 ;
  assign n7511 = ~n7508 & ~n7510 ;
  assign n7512 = \pi0299  & ~n7486 ;
  assign n7513 = ~\pi0039  & ~n7512 ;
  assign n7514 = ~\pi0039  & n1281 ;
  assign n7515 = n7491 & n7514 ;
  assign n7516 = ~n7513 & ~n7515 ;
  assign n7517 = n2363 & ~n7516 ;
  assign n7518 = n7511 & n7517 ;
  assign n7519 = ~n2342 & n7503 ;
  assign n7520 = n2364 & ~n7519 ;
  assign n7521 = ~n2511 & n7520 ;
  assign n7522 = ~n7518 & n7521 ;
  assign n7523 = ~n7506 & ~n7522 ;
  assign n7524 = n7265 & ~n7519 ;
  assign n7525 = ~n7518 & n7524 ;
  assign n7526 = ~n7265 & ~n7503 ;
  assign n7527 = \pi0074  & ~n7526 ;
  assign n7528 = ~n7525 & n7527 ;
  assign n7529 = ~\pi0055  & ~n7528 ;
  assign n7530 = ~n7523 & n7529 ;
  assign n7531 = \pi0075  & ~n7519 ;
  assign n7532 = ~n7518 & n7531 ;
  assign n7533 = \pi0087  & n7503 ;
  assign n7534 = ~\pi0075  & ~n7533 ;
  assign n7535 = ~\pi0092  & ~n7534 ;
  assign n7536 = ~n7532 & n7535 ;
  assign n7537 = ~\pi0075  & ~n7519 ;
  assign n7538 = ~n7518 & n7537 ;
  assign n7539 = \pi0075  & ~n7503 ;
  assign n7540 = \pi0092  & ~n7539 ;
  assign n7541 = ~n7538 & n7540 ;
  assign n7542 = ~\pi0054  & ~n7541 ;
  assign n7543 = n7529 & n7542 ;
  assign n7544 = ~n7536 & n7543 ;
  assign n7545 = ~n7530 & ~n7544 ;
  assign n7546 = n6706 & ~n7097 ;
  assign n7547 = ~n7100 & ~n7546 ;
  assign n7548 = n6975 & ~n7100 ;
  assign n7549 = ~n7094 & ~n7100 ;
  assign n7550 = n7092 & n7549 ;
  assign n7551 = ~n7548 & ~n7550 ;
  assign n7552 = ~\pi0228  & n6706 ;
  assign n7553 = n6975 & n7552 ;
  assign n7554 = ~n7094 & n7552 ;
  assign n7555 = ~n7138 & n7554 ;
  assign n7556 = ~n7553 & ~n7555 ;
  assign n7557 = ~n7307 & n7556 ;
  assign n7558 = n7551 & n7557 ;
  assign n7559 = \pi0967  & ~n7558 ;
  assign n7560 = ~n7547 & n7559 ;
  assign n7561 = ~\pi0299  & ~n7560 ;
  assign n7562 = \pi0232  & ~n7561 ;
  assign n7563 = n7151 & n7489 ;
  assign n7564 = ~n7094 & n7489 ;
  assign n7565 = n7092 & n7564 ;
  assign n7566 = ~n7563 & ~n7565 ;
  assign n7567 = n7512 & n7566 ;
  assign n7568 = \pi0299  & n7160 ;
  assign n7569 = ~n7567 & ~n7568 ;
  assign n7570 = n6706 & n7151 ;
  assign n7571 = n6706 & ~n7094 ;
  assign n7572 = ~n7138 & n7571 ;
  assign n7573 = ~n7570 & ~n7572 ;
  assign n7574 = n7161 & n7573 ;
  assign n7575 = ~n7151 & ~n7161 ;
  assign n7576 = n7489 & ~n7575 ;
  assign n7577 = ~n7565 & ~n7576 ;
  assign n7578 = ~n7574 & ~n7577 ;
  assign n7579 = ~n7486 & ~n7578 ;
  assign n7580 = n7160 & ~n7579 ;
  assign n7581 = ~n7569 & ~n7580 ;
  assign n7582 = ~\pi0039  & ~n7581 ;
  assign n7583 = n7562 & n7582 ;
  assign n7584 = ~\pi0232  & ~n7567 ;
  assign n7585 = ~\pi0039  & \pi0299  ;
  assign n7586 = ~\pi0039  & n7507 ;
  assign n7587 = ~n7097 & n7586 ;
  assign n7588 = ~n7585 & ~n7587 ;
  assign n7589 = n7584 & ~n7588 ;
  assign n7590 = \pi0228  & n7500 ;
  assign n7591 = ~\pi0216  & n6923 ;
  assign n7592 = ~n6931 & n7591 ;
  assign n7593 = n1259 & n7592 ;
  assign n7594 = n1249 & n7593 ;
  assign n7595 = n6920 & n7594 ;
  assign n7596 = n6936 & n7595 ;
  assign n7597 = \pi0216  & n6936 ;
  assign n7598 = n6954 & n7597 ;
  assign n7599 = ~n7596 & ~n7598 ;
  assign n7600 = n6706 & n7500 ;
  assign n7601 = ~n7599 & n7600 ;
  assign n7602 = ~n7590 & ~n7601 ;
  assign n7603 = \pi0228  & n7501 ;
  assign n7604 = n6706 & n7501 ;
  assign n7605 = ~n6957 & n7604 ;
  assign n7606 = ~n7603 & ~n7605 ;
  assign n7607 = n7602 & n7606 ;
  assign n7608 = \pi0039  & ~\pi0228  ;
  assign n7609 = \pi0030  & \pi0039  ;
  assign n7610 = n6706 & n7609 ;
  assign n7611 = ~n7608 & ~n7610 ;
  assign n7612 = ~n7607 & ~n7611 ;
  assign n7613 = ~\pi0038  & ~n7612 ;
  assign n7614 = ~n7589 & n7613 ;
  assign n7615 = ~n7583 & n7614 ;
  assign n7616 = ~\pi0100  & n7615 ;
  assign n7617 = n1259 & n7234 ;
  assign n7618 = n1249 & n7617 ;
  assign n7619 = n7216 & n7618 ;
  assign n7620 = n6706 & ~n6808 ;
  assign n7621 = n7619 & n7620 ;
  assign n7622 = n1259 & ~n7234 ;
  assign n7623 = n1249 & n7622 ;
  assign n7624 = n7210 & n7623 ;
  assign n7625 = ~\pi0228  & ~n7624 ;
  assign n7626 = ~n7621 & n7625 ;
  assign n7627 = ~\pi0228  & \pi0967  ;
  assign n7628 = \pi0030  & \pi0967  ;
  assign n7629 = n6706 & n7628 ;
  assign n7630 = ~n7627 & ~n7629 ;
  assign n7631 = ~n7626 & ~n7630 ;
  assign n7632 = ~\pi0299  & ~n7631 ;
  assign n7633 = n1259 & ~n6808 ;
  assign n7634 = n1249 & n7633 ;
  assign n7635 = n7216 & n7634 ;
  assign n7636 = n6706 & n7635 ;
  assign n7637 = n2070 & ~n7636 ;
  assign n7638 = ~n2070 & ~n7422 ;
  assign n7639 = n7488 & ~n7638 ;
  assign n7640 = ~n7637 & n7639 ;
  assign n7641 = n7512 & ~n7640 ;
  assign n7642 = n1288 & ~n7641 ;
  assign n7643 = ~n7632 & n7642 ;
  assign n7644 = ~n1288 & n7503 ;
  assign n7645 = \pi0100  & ~n7644 ;
  assign n7646 = ~n7643 & n7645 ;
  assign n7647 = \pi0039  & n7503 ;
  assign n7648 = \pi0038  & ~n7647 ;
  assign n7649 = n7516 & n7648 ;
  assign n7650 = ~\pi0100  & n7649 ;
  assign n7651 = ~\pi0100  & n7648 ;
  assign n7652 = ~n7511 & n7651 ;
  assign n7653 = ~n7650 & ~n7652 ;
  assign n7654 = ~\pi0087  & n7653 ;
  assign n7655 = ~n7646 & n7654 ;
  assign n7656 = ~n7616 & n7655 ;
  assign n7657 = ~\pi0092  & ~n7532 ;
  assign n7658 = ~n7530 & n7657 ;
  assign n7659 = n7656 & n7658 ;
  assign n7660 = ~n7545 & ~n7659 ;
  assign n7661 = \pi0970  & n1292 ;
  assign n7662 = n7307 & n7661 ;
  assign n7663 = ~n1293 & ~n7662 ;
  assign n7664 = n1291 & n1292 ;
  assign n7665 = n1281 & n7664 ;
  assign n7666 = n7491 & n7665 ;
  assign n7667 = n7663 & ~n7666 ;
  assign n7668 = n7495 & ~n7667 ;
  assign n7669 = ~n7660 & n7668 ;
  assign n7670 = ~n7499 & ~n7669 ;
  assign n7671 = ~n7486 & ~n7493 ;
  assign n7672 = \pi0057  & ~\pi0059  ;
  assign n7673 = \pi0057  & \pi0970  ;
  assign n7674 = n7307 & n7673 ;
  assign n7675 = ~n7672 & ~n7674 ;
  assign n7676 = ~n7671 & ~n7675 ;
  assign n7677 = n7670 & ~n7676 ;
  assign n7678 = \pi0972  & n7307 ;
  assign n7679 = \pi0059  & ~n7678 ;
  assign n7680 = ~\pi0228  & \pi0972  ;
  assign n7681 = n6706 & n7680 ;
  assign n7682 = n1259 & n7681 ;
  assign n7683 = n1249 & n7682 ;
  assign n7684 = n7492 & n7683 ;
  assign n7685 = n7679 & ~n7684 ;
  assign n7686 = ~\pi0057  & ~n7685 ;
  assign n7687 = \pi0972  & ~n1292 ;
  assign n7688 = n7307 & n7687 ;
  assign n7689 = ~\pi0059  & ~n7688 ;
  assign n7690 = n7686 & ~n7689 ;
  assign n7691 = ~\pi0299  & \pi0961  ;
  assign n7692 = \pi0299  & \pi0972  ;
  assign n7693 = ~n7691 & ~n7692 ;
  assign n7694 = n7307 & ~n7693 ;
  assign n7695 = ~n2364 & ~n7694 ;
  assign n7696 = ~\pi0074  & ~n7695 ;
  assign n7697 = ~n2511 & ~n7696 ;
  assign n7698 = \pi0961  & n6706 ;
  assign n7699 = ~\pi0299  & ~n7698 ;
  assign n7700 = ~n7510 & ~n7699 ;
  assign n7701 = \pi0299  & ~n7678 ;
  assign n7702 = ~\pi0039  & ~n7701 ;
  assign n7703 = n7514 & n7683 ;
  assign n7704 = ~n7702 & ~n7703 ;
  assign n7705 = n2363 & ~n7704 ;
  assign n7706 = n7700 & n7705 ;
  assign n7707 = ~n2342 & n7694 ;
  assign n7708 = n2364 & ~n7707 ;
  assign n7709 = ~n2511 & n7708 ;
  assign n7710 = ~n7706 & n7709 ;
  assign n7711 = ~n7697 & ~n7710 ;
  assign n7712 = n7265 & ~n7707 ;
  assign n7713 = ~n7706 & n7712 ;
  assign n7714 = ~n7265 & ~n7694 ;
  assign n7715 = \pi0074  & ~n7714 ;
  assign n7716 = ~n7713 & n7715 ;
  assign n7717 = ~\pi0055  & ~n7716 ;
  assign n7718 = ~n7711 & n7717 ;
  assign n7719 = \pi0075  & ~n7707 ;
  assign n7720 = ~n7706 & n7719 ;
  assign n7721 = \pi0087  & n7694 ;
  assign n7722 = ~\pi0075  & ~n7721 ;
  assign n7723 = ~\pi0092  & ~n7722 ;
  assign n7724 = ~n7720 & n7723 ;
  assign n7725 = ~\pi0075  & ~n7707 ;
  assign n7726 = ~n7706 & n7725 ;
  assign n7727 = \pi0075  & ~n7694 ;
  assign n7728 = \pi0092  & ~n7727 ;
  assign n7729 = ~n7726 & n7728 ;
  assign n7730 = ~\pi0054  & ~n7729 ;
  assign n7731 = n7717 & n7730 ;
  assign n7732 = ~n7724 & n7731 ;
  assign n7733 = ~n7718 & ~n7732 ;
  assign n7734 = \pi0961  & ~n7558 ;
  assign n7735 = ~n7547 & n7734 ;
  assign n7736 = ~\pi0299  & ~n7735 ;
  assign n7737 = \pi0232  & ~n7736 ;
  assign n7738 = n7151 & n7681 ;
  assign n7739 = ~n7094 & n7681 ;
  assign n7740 = n7092 & n7739 ;
  assign n7741 = ~n7738 & ~n7740 ;
  assign n7742 = n7701 & n7741 ;
  assign n7743 = ~n7568 & ~n7742 ;
  assign n7744 = n7160 & n7678 ;
  assign n7745 = ~n7146 & n7575 ;
  assign n7746 = ~n7574 & ~n7745 ;
  assign n7747 = n7160 & n7681 ;
  assign n7748 = n7746 & n7747 ;
  assign n7749 = ~n7744 & ~n7748 ;
  assign n7750 = ~n7743 & n7749 ;
  assign n7751 = ~\pi0039  & ~n7750 ;
  assign n7752 = n7737 & n7751 ;
  assign n7753 = ~\pi0232  & ~n7742 ;
  assign n7754 = ~\pi0039  & n7698 ;
  assign n7755 = ~n7097 & n7754 ;
  assign n7756 = ~n7585 & ~n7755 ;
  assign n7757 = n7753 & ~n7756 ;
  assign n7758 = \pi0228  & n7691 ;
  assign n7759 = n6706 & n7691 ;
  assign n7760 = ~n6957 & n7759 ;
  assign n7761 = ~n7758 & ~n7760 ;
  assign n7762 = \pi0228  & n7692 ;
  assign n7763 = n6706 & n7692 ;
  assign n7764 = ~n7599 & n7763 ;
  assign n7765 = ~n7762 & ~n7764 ;
  assign n7766 = n7761 & n7765 ;
  assign n7767 = ~n7611 & ~n7766 ;
  assign n7768 = ~\pi0038  & ~n7767 ;
  assign n7769 = ~n7757 & n7768 ;
  assign n7770 = ~n7752 & n7769 ;
  assign n7771 = ~\pi0100  & n7770 ;
  assign n7772 = \pi0030  & n6706 ;
  assign n7773 = \pi0228  & ~n7772 ;
  assign n7774 = \pi0961  & ~n7773 ;
  assign n7775 = ~n7626 & n7774 ;
  assign n7776 = ~\pi0299  & ~n7775 ;
  assign n7777 = ~n7638 & n7680 ;
  assign n7778 = ~n7637 & n7777 ;
  assign n7779 = n7701 & ~n7778 ;
  assign n7780 = n1288 & ~n7779 ;
  assign n7781 = ~n7776 & n7780 ;
  assign n7782 = ~n1288 & n7694 ;
  assign n7783 = \pi0100  & ~n7782 ;
  assign n7784 = ~n7781 & n7783 ;
  assign n7785 = \pi0039  & n7694 ;
  assign n7786 = \pi0038  & ~n7785 ;
  assign n7787 = n7704 & n7786 ;
  assign n7788 = ~\pi0100  & n7787 ;
  assign n7789 = ~\pi0100  & n7786 ;
  assign n7790 = ~n7700 & n7789 ;
  assign n7791 = ~n7788 & ~n7790 ;
  assign n7792 = ~\pi0087  & n7791 ;
  assign n7793 = ~n7784 & n7792 ;
  assign n7794 = ~n7771 & n7793 ;
  assign n7795 = ~\pi0092  & ~n7720 ;
  assign n7796 = ~n7718 & n7795 ;
  assign n7797 = n7794 & n7796 ;
  assign n7798 = ~n7733 & ~n7797 ;
  assign n7799 = \pi0972  & n1292 ;
  assign n7800 = n7307 & n7799 ;
  assign n7801 = ~n1293 & ~n7800 ;
  assign n7802 = n7665 & n7683 ;
  assign n7803 = n7801 & ~n7802 ;
  assign n7804 = n7686 & ~n7803 ;
  assign n7805 = ~n7798 & n7804 ;
  assign n7806 = ~n7690 & ~n7805 ;
  assign n7807 = ~n7678 & ~n7684 ;
  assign n7808 = \pi0057  & \pi0972  ;
  assign n7809 = n7307 & n7808 ;
  assign n7810 = ~n7672 & ~n7809 ;
  assign n7811 = ~n7807 & ~n7810 ;
  assign n7812 = n7806 & ~n7811 ;
  assign n7813 = \pi0960  & n7307 ;
  assign n7814 = \pi0059  & ~n7813 ;
  assign n7815 = ~\pi0228  & \pi0960  ;
  assign n7816 = n6706 & n7815 ;
  assign n7817 = n1259 & n7816 ;
  assign n7818 = n1249 & n7817 ;
  assign n7819 = n7492 & n7818 ;
  assign n7820 = n7814 & ~n7819 ;
  assign n7821 = ~\pi0057  & ~n7820 ;
  assign n7822 = \pi0960  & ~n1292 ;
  assign n7823 = n7307 & n7822 ;
  assign n7824 = ~\pi0059  & ~n7823 ;
  assign n7825 = n7821 & ~n7824 ;
  assign n7826 = ~\pi0299  & \pi0977  ;
  assign n7827 = \pi0299  & \pi0960  ;
  assign n7828 = ~n7826 & ~n7827 ;
  assign n7829 = n7307 & ~n7828 ;
  assign n7830 = ~n2364 & ~n7829 ;
  assign n7831 = ~\pi0074  & ~n7830 ;
  assign n7832 = ~n2511 & ~n7831 ;
  assign n7833 = \pi0977  & n6706 ;
  assign n7834 = ~\pi0299  & ~n7833 ;
  assign n7835 = ~n7510 & ~n7834 ;
  assign n7836 = \pi0299  & ~n7813 ;
  assign n7837 = ~\pi0039  & ~n7836 ;
  assign n7838 = n7514 & n7818 ;
  assign n7839 = ~n7837 & ~n7838 ;
  assign n7840 = n2363 & ~n7839 ;
  assign n7841 = n7835 & n7840 ;
  assign n7842 = ~n2342 & n7829 ;
  assign n7843 = n2364 & ~n7842 ;
  assign n7844 = ~n2511 & n7843 ;
  assign n7845 = ~n7841 & n7844 ;
  assign n7846 = ~n7832 & ~n7845 ;
  assign n7847 = n7265 & ~n7842 ;
  assign n7848 = ~n7841 & n7847 ;
  assign n7849 = ~n7265 & ~n7829 ;
  assign n7850 = \pi0074  & ~n7849 ;
  assign n7851 = ~n7848 & n7850 ;
  assign n7852 = ~\pi0055  & ~n7851 ;
  assign n7853 = ~n7846 & n7852 ;
  assign n7854 = \pi0075  & ~n7842 ;
  assign n7855 = ~n7841 & n7854 ;
  assign n7856 = \pi0087  & n7829 ;
  assign n7857 = ~\pi0075  & ~n7856 ;
  assign n7858 = ~\pi0092  & ~n7857 ;
  assign n7859 = ~n7855 & n7858 ;
  assign n7860 = ~\pi0075  & ~n7842 ;
  assign n7861 = ~n7841 & n7860 ;
  assign n7862 = \pi0075  & ~n7829 ;
  assign n7863 = \pi0092  & ~n7862 ;
  assign n7864 = ~n7861 & n7863 ;
  assign n7865 = ~\pi0054  & ~n7864 ;
  assign n7866 = n7852 & n7865 ;
  assign n7867 = ~n7859 & n7866 ;
  assign n7868 = ~n7853 & ~n7867 ;
  assign n7869 = \pi0977  & ~n7558 ;
  assign n7870 = ~n7547 & n7869 ;
  assign n7871 = ~\pi0299  & ~n7870 ;
  assign n7872 = \pi0232  & ~n7871 ;
  assign n7873 = n7151 & n7816 ;
  assign n7874 = ~n7094 & n7816 ;
  assign n7875 = n7092 & n7874 ;
  assign n7876 = ~n7873 & ~n7875 ;
  assign n7877 = n7836 & n7876 ;
  assign n7878 = ~n7568 & ~n7877 ;
  assign n7879 = n7160 & n7813 ;
  assign n7880 = n7160 & n7816 ;
  assign n7881 = n7746 & n7880 ;
  assign n7882 = ~n7879 & ~n7881 ;
  assign n7883 = ~n7878 & n7882 ;
  assign n7884 = ~\pi0039  & ~n7883 ;
  assign n7885 = n7872 & n7884 ;
  assign n7886 = ~\pi0232  & ~n7877 ;
  assign n7887 = ~\pi0039  & n7833 ;
  assign n7888 = ~n7097 & n7887 ;
  assign n7889 = ~n7585 & ~n7888 ;
  assign n7890 = n7886 & ~n7889 ;
  assign n7891 = \pi0228  & n7826 ;
  assign n7892 = n6706 & n7826 ;
  assign n7893 = ~n6957 & n7892 ;
  assign n7894 = ~n7891 & ~n7893 ;
  assign n7895 = \pi0228  & n7827 ;
  assign n7896 = n6706 & n7827 ;
  assign n7897 = ~n7599 & n7896 ;
  assign n7898 = ~n7895 & ~n7897 ;
  assign n7899 = n7894 & n7898 ;
  assign n7900 = ~n7611 & ~n7899 ;
  assign n7901 = ~\pi0038  & ~n7900 ;
  assign n7902 = ~n7890 & n7901 ;
  assign n7903 = ~n7885 & n7902 ;
  assign n7904 = ~\pi0100  & n7903 ;
  assign n7905 = \pi0977  & ~n7773 ;
  assign n7906 = ~n7626 & n7905 ;
  assign n7907 = ~\pi0299  & ~n7906 ;
  assign n7908 = ~n7638 & n7815 ;
  assign n7909 = ~n7637 & n7908 ;
  assign n7910 = n7836 & ~n7909 ;
  assign n7911 = n1288 & ~n7910 ;
  assign n7912 = ~n7907 & n7911 ;
  assign n7913 = ~n1288 & n7829 ;
  assign n7914 = \pi0100  & ~n7913 ;
  assign n7915 = ~n7912 & n7914 ;
  assign n7916 = \pi0039  & n7829 ;
  assign n7917 = \pi0038  & ~n7916 ;
  assign n7918 = n7839 & n7917 ;
  assign n7919 = ~\pi0100  & n7918 ;
  assign n7920 = ~\pi0100  & n7917 ;
  assign n7921 = ~n7835 & n7920 ;
  assign n7922 = ~n7919 & ~n7921 ;
  assign n7923 = ~\pi0087  & n7922 ;
  assign n7924 = ~n7915 & n7923 ;
  assign n7925 = ~n7904 & n7924 ;
  assign n7926 = ~\pi0092  & ~n7855 ;
  assign n7927 = ~n7853 & n7926 ;
  assign n7928 = n7925 & n7927 ;
  assign n7929 = ~n7868 & ~n7928 ;
  assign n7930 = \pi0960  & n1292 ;
  assign n7931 = n7307 & n7930 ;
  assign n7932 = ~n1293 & ~n7931 ;
  assign n7933 = n7665 & n7818 ;
  assign n7934 = n7932 & ~n7933 ;
  assign n7935 = n7821 & ~n7934 ;
  assign n7936 = ~n7929 & n7935 ;
  assign n7937 = ~n7825 & ~n7936 ;
  assign n7938 = ~n7813 & ~n7819 ;
  assign n7939 = \pi0057  & \pi0960  ;
  assign n7940 = n7307 & n7939 ;
  assign n7941 = ~n7672 & ~n7940 ;
  assign n7942 = ~n7938 & ~n7941 ;
  assign n7943 = n7937 & ~n7942 ;
  assign n7944 = \pi0963  & n7307 ;
  assign n7945 = \pi0059  & ~n7944 ;
  assign n7946 = ~\pi0228  & \pi0963  ;
  assign n7947 = n6706 & n7946 ;
  assign n7948 = n1259 & n7947 ;
  assign n7949 = n1249 & n7948 ;
  assign n7950 = n7492 & n7949 ;
  assign n7951 = n7945 & ~n7950 ;
  assign n7952 = ~\pi0057  & ~n7951 ;
  assign n7953 = \pi0963  & ~n1292 ;
  assign n7954 = n7307 & n7953 ;
  assign n7955 = ~\pi0059  & ~n7954 ;
  assign n7956 = n7952 & ~n7955 ;
  assign n7957 = ~\pi0299  & \pi0969  ;
  assign n7958 = \pi0299  & \pi0963  ;
  assign n7959 = ~n7957 & ~n7958 ;
  assign n7960 = n7307 & ~n7959 ;
  assign n7961 = ~n2364 & ~n7960 ;
  assign n7962 = ~\pi0074  & ~n7961 ;
  assign n7963 = ~n2511 & ~n7962 ;
  assign n7964 = \pi0969  & n6706 ;
  assign n7965 = ~\pi0299  & ~n7964 ;
  assign n7966 = ~n7510 & ~n7965 ;
  assign n7967 = \pi0299  & ~n7944 ;
  assign n7968 = ~\pi0039  & ~n7967 ;
  assign n7969 = n7514 & n7949 ;
  assign n7970 = ~n7968 & ~n7969 ;
  assign n7971 = n2363 & ~n7970 ;
  assign n7972 = n7966 & n7971 ;
  assign n7973 = ~n2342 & n7960 ;
  assign n7974 = n2364 & ~n7973 ;
  assign n7975 = ~n2511 & n7974 ;
  assign n7976 = ~n7972 & n7975 ;
  assign n7977 = ~n7963 & ~n7976 ;
  assign n7978 = n7265 & ~n7973 ;
  assign n7979 = ~n7972 & n7978 ;
  assign n7980 = ~n7265 & ~n7960 ;
  assign n7981 = \pi0074  & ~n7980 ;
  assign n7982 = ~n7979 & n7981 ;
  assign n7983 = ~\pi0055  & ~n7982 ;
  assign n7984 = ~n7977 & n7983 ;
  assign n7985 = \pi0075  & ~n7973 ;
  assign n7986 = ~n7972 & n7985 ;
  assign n7987 = \pi0087  & n7960 ;
  assign n7988 = ~\pi0075  & ~n7987 ;
  assign n7989 = ~\pi0092  & ~n7988 ;
  assign n7990 = ~n7986 & n7989 ;
  assign n7991 = ~\pi0075  & ~n7973 ;
  assign n7992 = ~n7972 & n7991 ;
  assign n7993 = \pi0075  & ~n7960 ;
  assign n7994 = \pi0092  & ~n7993 ;
  assign n7995 = ~n7992 & n7994 ;
  assign n7996 = ~\pi0054  & ~n7995 ;
  assign n7997 = n7983 & n7996 ;
  assign n7998 = ~n7990 & n7997 ;
  assign n7999 = ~n7984 & ~n7998 ;
  assign n8000 = \pi0969  & ~n7558 ;
  assign n8001 = ~n7547 & n8000 ;
  assign n8002 = ~\pi0299  & ~n8001 ;
  assign n8003 = \pi0232  & ~n8002 ;
  assign n8004 = n7151 & n7947 ;
  assign n8005 = ~n7094 & n7947 ;
  assign n8006 = n7092 & n8005 ;
  assign n8007 = ~n8004 & ~n8006 ;
  assign n8008 = n7967 & n8007 ;
  assign n8009 = ~n7568 & ~n8008 ;
  assign n8010 = n7160 & n7944 ;
  assign n8011 = n7160 & n7947 ;
  assign n8012 = n7746 & n8011 ;
  assign n8013 = ~n8010 & ~n8012 ;
  assign n8014 = ~n8009 & n8013 ;
  assign n8015 = ~\pi0039  & ~n8014 ;
  assign n8016 = n8003 & n8015 ;
  assign n8017 = ~\pi0232  & ~n8008 ;
  assign n8018 = ~\pi0039  & n7964 ;
  assign n8019 = ~n7097 & n8018 ;
  assign n8020 = ~n7585 & ~n8019 ;
  assign n8021 = n8017 & ~n8020 ;
  assign n8022 = \pi0228  & n7957 ;
  assign n8023 = n6706 & n7957 ;
  assign n8024 = ~n6957 & n8023 ;
  assign n8025 = ~n8022 & ~n8024 ;
  assign n8026 = \pi0228  & n7958 ;
  assign n8027 = n6706 & n7958 ;
  assign n8028 = ~n7599 & n8027 ;
  assign n8029 = ~n8026 & ~n8028 ;
  assign n8030 = n8025 & n8029 ;
  assign n8031 = ~n7611 & ~n8030 ;
  assign n8032 = ~\pi0038  & ~n8031 ;
  assign n8033 = ~n8021 & n8032 ;
  assign n8034 = ~n8016 & n8033 ;
  assign n8035 = ~\pi0100  & n8034 ;
  assign n8036 = \pi0969  & ~n7773 ;
  assign n8037 = ~n7626 & n8036 ;
  assign n8038 = ~\pi0299  & ~n8037 ;
  assign n8039 = ~n7638 & n7946 ;
  assign n8040 = ~n7637 & n8039 ;
  assign n8041 = n7967 & ~n8040 ;
  assign n8042 = n1288 & ~n8041 ;
  assign n8043 = ~n8038 & n8042 ;
  assign n8044 = ~n1288 & n7960 ;
  assign n8045 = \pi0100  & ~n8044 ;
  assign n8046 = ~n8043 & n8045 ;
  assign n8047 = \pi0039  & n7960 ;
  assign n8048 = \pi0038  & ~n8047 ;
  assign n8049 = n7970 & n8048 ;
  assign n8050 = ~\pi0100  & n8049 ;
  assign n8051 = ~\pi0100  & n8048 ;
  assign n8052 = ~n7966 & n8051 ;
  assign n8053 = ~n8050 & ~n8052 ;
  assign n8054 = ~\pi0087  & n8053 ;
  assign n8055 = ~n8046 & n8054 ;
  assign n8056 = ~n8035 & n8055 ;
  assign n8057 = ~\pi0092  & ~n7986 ;
  assign n8058 = ~n7984 & n8057 ;
  assign n8059 = n8056 & n8058 ;
  assign n8060 = ~n7999 & ~n8059 ;
  assign n8061 = \pi0963  & n1292 ;
  assign n8062 = n7307 & n8061 ;
  assign n8063 = ~n1293 & ~n8062 ;
  assign n8064 = n7665 & n7949 ;
  assign n8065 = n8063 & ~n8064 ;
  assign n8066 = n7952 & ~n8065 ;
  assign n8067 = ~n8060 & n8066 ;
  assign n8068 = ~n7956 & ~n8067 ;
  assign n8069 = ~n7944 & ~n7950 ;
  assign n8070 = \pi0057  & \pi0963  ;
  assign n8071 = n7307 & n8070 ;
  assign n8072 = ~n7672 & ~n8071 ;
  assign n8073 = ~n8069 & ~n8072 ;
  assign n8074 = n8068 & ~n8073 ;
  assign n8075 = \pi0975  & n7307 ;
  assign n8076 = \pi0059  & ~n8075 ;
  assign n8077 = ~\pi0228  & \pi0975  ;
  assign n8078 = n6706 & n8077 ;
  assign n8079 = n1259 & n8078 ;
  assign n8080 = n1249 & n8079 ;
  assign n8081 = n7492 & n8080 ;
  assign n8082 = n8076 & ~n8081 ;
  assign n8083 = ~\pi0057  & ~n8082 ;
  assign n8084 = \pi0975  & ~n1292 ;
  assign n8085 = n7307 & n8084 ;
  assign n8086 = ~\pi0059  & ~n8085 ;
  assign n8087 = n8083 & ~n8086 ;
  assign n8088 = ~\pi0299  & \pi0971  ;
  assign n8089 = \pi0299  & \pi0975  ;
  assign n8090 = ~n8088 & ~n8089 ;
  assign n8091 = n7307 & ~n8090 ;
  assign n8092 = ~n2364 & ~n8091 ;
  assign n8093 = ~\pi0074  & ~n8092 ;
  assign n8094 = ~n2511 & ~n8093 ;
  assign n8095 = \pi0971  & n6706 ;
  assign n8096 = ~\pi0299  & ~n8095 ;
  assign n8097 = ~n7510 & ~n8096 ;
  assign n8098 = \pi0299  & ~n8075 ;
  assign n8099 = ~\pi0039  & ~n8098 ;
  assign n8100 = n7514 & n8080 ;
  assign n8101 = ~n8099 & ~n8100 ;
  assign n8102 = n2363 & ~n8101 ;
  assign n8103 = n8097 & n8102 ;
  assign n8104 = ~n2342 & n8091 ;
  assign n8105 = n2364 & ~n8104 ;
  assign n8106 = ~n2511 & n8105 ;
  assign n8107 = ~n8103 & n8106 ;
  assign n8108 = ~n8094 & ~n8107 ;
  assign n8109 = n7265 & ~n8104 ;
  assign n8110 = ~n8103 & n8109 ;
  assign n8111 = ~n7265 & ~n8091 ;
  assign n8112 = \pi0074  & ~n8111 ;
  assign n8113 = ~n8110 & n8112 ;
  assign n8114 = ~\pi0055  & ~n8113 ;
  assign n8115 = ~n8108 & n8114 ;
  assign n8116 = \pi0075  & ~n8104 ;
  assign n8117 = ~n8103 & n8116 ;
  assign n8118 = \pi0087  & n8091 ;
  assign n8119 = ~\pi0075  & ~n8118 ;
  assign n8120 = ~\pi0092  & ~n8119 ;
  assign n8121 = ~n8117 & n8120 ;
  assign n8122 = ~\pi0075  & ~n8104 ;
  assign n8123 = ~n8103 & n8122 ;
  assign n8124 = \pi0075  & ~n8091 ;
  assign n8125 = \pi0092  & ~n8124 ;
  assign n8126 = ~n8123 & n8125 ;
  assign n8127 = ~\pi0054  & ~n8126 ;
  assign n8128 = n8114 & n8127 ;
  assign n8129 = ~n8121 & n8128 ;
  assign n8130 = ~n8115 & ~n8129 ;
  assign n8131 = \pi0971  & ~n7558 ;
  assign n8132 = ~n7547 & n8131 ;
  assign n8133 = ~\pi0299  & ~n8132 ;
  assign n8134 = \pi0232  & ~n8133 ;
  assign n8135 = n7151 & n8078 ;
  assign n8136 = ~n7094 & n8078 ;
  assign n8137 = n7092 & n8136 ;
  assign n8138 = ~n8135 & ~n8137 ;
  assign n8139 = n8098 & n8138 ;
  assign n8140 = ~n7568 & ~n8139 ;
  assign n8141 = n7160 & n8075 ;
  assign n8142 = n7160 & n8078 ;
  assign n8143 = n7746 & n8142 ;
  assign n8144 = ~n8141 & ~n8143 ;
  assign n8145 = ~n8140 & n8144 ;
  assign n8146 = ~\pi0039  & ~n8145 ;
  assign n8147 = n8134 & n8146 ;
  assign n8148 = ~\pi0232  & ~n8139 ;
  assign n8149 = ~\pi0039  & n8095 ;
  assign n8150 = ~n7097 & n8149 ;
  assign n8151 = ~n7585 & ~n8150 ;
  assign n8152 = n8148 & ~n8151 ;
  assign n8153 = \pi0228  & n8088 ;
  assign n8154 = n6706 & n8088 ;
  assign n8155 = ~n6957 & n8154 ;
  assign n8156 = ~n8153 & ~n8155 ;
  assign n8157 = \pi0228  & n8089 ;
  assign n8158 = n6706 & n8089 ;
  assign n8159 = ~n7599 & n8158 ;
  assign n8160 = ~n8157 & ~n8159 ;
  assign n8161 = n8156 & n8160 ;
  assign n8162 = ~n7611 & ~n8161 ;
  assign n8163 = ~\pi0038  & ~n8162 ;
  assign n8164 = ~n8152 & n8163 ;
  assign n8165 = ~n8147 & n8164 ;
  assign n8166 = ~\pi0100  & n8165 ;
  assign n8167 = \pi0971  & ~n7773 ;
  assign n8168 = ~n7626 & n8167 ;
  assign n8169 = ~\pi0299  & ~n8168 ;
  assign n8170 = ~n7638 & n8077 ;
  assign n8171 = ~n7637 & n8170 ;
  assign n8172 = n8098 & ~n8171 ;
  assign n8173 = n1288 & ~n8172 ;
  assign n8174 = ~n8169 & n8173 ;
  assign n8175 = ~n1288 & n8091 ;
  assign n8176 = \pi0100  & ~n8175 ;
  assign n8177 = ~n8174 & n8176 ;
  assign n8178 = \pi0039  & n8091 ;
  assign n8179 = \pi0038  & ~n8178 ;
  assign n8180 = n8101 & n8179 ;
  assign n8181 = ~\pi0100  & n8180 ;
  assign n8182 = ~\pi0100  & n8179 ;
  assign n8183 = ~n8097 & n8182 ;
  assign n8184 = ~n8181 & ~n8183 ;
  assign n8185 = ~\pi0087  & n8184 ;
  assign n8186 = ~n8177 & n8185 ;
  assign n8187 = ~n8166 & n8186 ;
  assign n8188 = ~\pi0092  & ~n8117 ;
  assign n8189 = ~n8115 & n8188 ;
  assign n8190 = n8187 & n8189 ;
  assign n8191 = ~n8130 & ~n8190 ;
  assign n8192 = \pi0975  & n1292 ;
  assign n8193 = n7307 & n8192 ;
  assign n8194 = ~n1293 & ~n8193 ;
  assign n8195 = n7665 & n8080 ;
  assign n8196 = n8194 & ~n8195 ;
  assign n8197 = n8083 & ~n8196 ;
  assign n8198 = ~n8191 & n8197 ;
  assign n8199 = ~n8087 & ~n8198 ;
  assign n8200 = ~n8075 & ~n8081 ;
  assign n8201 = \pi0057  & \pi0975  ;
  assign n8202 = n7307 & n8201 ;
  assign n8203 = ~n7672 & ~n8202 ;
  assign n8204 = ~n8200 & ~n8203 ;
  assign n8205 = n8199 & ~n8204 ;
  assign n8206 = ~\pi0299  & \pi0974  ;
  assign n8207 = \pi0299  & \pi0978  ;
  assign n8208 = ~n8206 & ~n8207 ;
  assign n8209 = n6706 & ~n8208 ;
  assign n8210 = ~\pi0228  & ~n2342 ;
  assign n8211 = n8209 & ~n8210 ;
  assign n8212 = n7265 & ~n8211 ;
  assign n8213 = ~n6853 & n7265 ;
  assign n8214 = ~n3421 & n8213 ;
  assign n8215 = ~n8212 & ~n8214 ;
  assign n8216 = n7307 & ~n8208 ;
  assign n8217 = ~n7265 & ~n8216 ;
  assign n8218 = \pi0074  & ~n8217 ;
  assign n8219 = n8215 & n8218 ;
  assign n8220 = ~\pi0055  & ~n8219 ;
  assign n8221 = ~\pi0057  & \pi0978  ;
  assign n8222 = n7307 & n8221 ;
  assign n8223 = ~n2467 & ~n8222 ;
  assign n8224 = ~\pi0228  & \pi0978  ;
  assign n8225 = n6706 & n8224 ;
  assign n8226 = n1259 & n8225 ;
  assign n8227 = n1249 & n8226 ;
  assign n8228 = ~\pi0057  & n1293 ;
  assign n8229 = n1291 & n8228 ;
  assign n8230 = n1281 & n8229 ;
  assign n8231 = n8227 & n8230 ;
  assign n8232 = n8223 & ~n8231 ;
  assign n8233 = \pi0978  & n1292 ;
  assign n8234 = n7307 & n8233 ;
  assign n8235 = ~n1293 & ~n8234 ;
  assign n8236 = n7665 & n8227 ;
  assign n8237 = n8235 & ~n8236 ;
  assign n8238 = ~n8232 & ~n8237 ;
  assign n8239 = ~n8220 & n8238 ;
  assign n8240 = \pi0075  & ~n8211 ;
  assign n8241 = \pi0075  & ~n6853 ;
  assign n8242 = ~n3421 & n8241 ;
  assign n8243 = ~n8240 & ~n8242 ;
  assign n8244 = ~\pi0092  & n8243 ;
  assign n8245 = ~\pi0054  & \pi0075  ;
  assign n8246 = ~n8216 & n8245 ;
  assign n8247 = ~n1285 & ~n8246 ;
  assign n8248 = ~\pi0054  & ~\pi0075  ;
  assign n8249 = ~n8211 & n8248 ;
  assign n8250 = ~n6853 & n8248 ;
  assign n8251 = ~n3421 & n8250 ;
  assign n8252 = ~n8249 & ~n8251 ;
  assign n8253 = n8247 & n8252 ;
  assign n8254 = ~n8244 & ~n8253 ;
  assign n8255 = \pi0974  & n6706 ;
  assign n8256 = ~n7097 & n8255 ;
  assign n8257 = ~\pi0299  & ~n8256 ;
  assign n8258 = \pi0978  & n7307 ;
  assign n8259 = \pi0299  & ~n8258 ;
  assign n8260 = n7151 & n8225 ;
  assign n8261 = ~n7094 & n8225 ;
  assign n8262 = n7092 & n8261 ;
  assign n8263 = ~n8260 & ~n8262 ;
  assign n8264 = n8259 & n8263 ;
  assign n8265 = ~\pi0232  & ~n8264 ;
  assign n8266 = ~n8257 & n8265 ;
  assign n8267 = ~\pi0039  & n8266 ;
  assign n8268 = \pi0974  & ~n7558 ;
  assign n8269 = ~n7547 & n8268 ;
  assign n8270 = ~\pi0299  & ~n8269 ;
  assign n8271 = \pi0232  & ~n8270 ;
  assign n8272 = ~n7568 & ~n8264 ;
  assign n8273 = n7160 & n8258 ;
  assign n8274 = n7160 & n8225 ;
  assign n8275 = n7746 & n8274 ;
  assign n8276 = ~n8273 & ~n8275 ;
  assign n8277 = ~n8272 & n8276 ;
  assign n8278 = ~\pi0039  & ~n8277 ;
  assign n8279 = n8271 & n8278 ;
  assign n8280 = ~n8267 & ~n8279 ;
  assign n8281 = \pi0228  & n8206 ;
  assign n8282 = n6706 & n8206 ;
  assign n8283 = ~n6957 & n8282 ;
  assign n8284 = ~n8281 & ~n8283 ;
  assign n8285 = \pi0228  & n8207 ;
  assign n8286 = n6706 & n8207 ;
  assign n8287 = ~n7599 & n8286 ;
  assign n8288 = ~n8285 & ~n8287 ;
  assign n8289 = n8284 & n8288 ;
  assign n8290 = ~n7611 & ~n8289 ;
  assign n8291 = n2327 & ~n8290 ;
  assign n8292 = n8280 & n8291 ;
  assign n8293 = \pi0039  & n8216 ;
  assign n8294 = \pi0038  & ~n8293 ;
  assign n8295 = ~\pi0039  & n6706 ;
  assign n8296 = ~n8208 & n8295 ;
  assign n8297 = ~\pi0100  & ~n8296 ;
  assign n8298 = ~\pi0100  & ~n6853 ;
  assign n8299 = ~n3421 & n8298 ;
  assign n8300 = ~n8297 & ~n8299 ;
  assign n8301 = n8294 & ~n8300 ;
  assign n8302 = ~n1288 & n8216 ;
  assign n8303 = \pi0100  & ~n8302 ;
  assign n8304 = ~\pi0087  & ~n8303 ;
  assign n8305 = ~n7638 & n8224 ;
  assign n8306 = ~n7637 & n8305 ;
  assign n8307 = n8259 & ~n8306 ;
  assign n8308 = n1288 & ~n8307 ;
  assign n8309 = \pi0974  & ~n7773 ;
  assign n8310 = ~n7626 & n8309 ;
  assign n8311 = ~\pi0299  & ~n8310 ;
  assign n8312 = ~\pi0087  & ~n8311 ;
  assign n8313 = n8308 & n8312 ;
  assign n8314 = ~n8304 & ~n8313 ;
  assign n8315 = ~n8301 & ~n8314 ;
  assign n8316 = ~n8292 & n8315 ;
  assign n8317 = \pi0087  & n8216 ;
  assign n8318 = ~\pi0075  & ~n8317 ;
  assign n8319 = ~n8253 & n8318 ;
  assign n8320 = ~n8316 & n8319 ;
  assign n8321 = ~n8254 & ~n8320 ;
  assign n8322 = \pi0054  & n2364 ;
  assign n8323 = ~n8211 & n8322 ;
  assign n8324 = ~n6853 & n8322 ;
  assign n8325 = ~n3421 & n8324 ;
  assign n8326 = ~n8323 & ~n8325 ;
  assign n8327 = \pi0054  & ~n2364 ;
  assign n8328 = ~n8216 & n8327 ;
  assign n8329 = ~\pi0074  & ~n8328 ;
  assign n8330 = n8326 & n8329 ;
  assign n8331 = n8238 & n8330 ;
  assign n8332 = n8321 & n8331 ;
  assign n8333 = ~n8239 & ~n8332 ;
  assign n8334 = \pi0978  & ~n1292 ;
  assign n8335 = n7307 & n8334 ;
  assign n8336 = ~\pi0059  & ~n8335 ;
  assign n8337 = ~n8232 & ~n8336 ;
  assign n8338 = \pi0057  & \pi0978  ;
  assign n8339 = n7307 & n8338 ;
  assign n8340 = ~n7672 & ~n8339 ;
  assign n8341 = n1294 & ~n8340 ;
  assign n8342 = n1281 & n8341 ;
  assign n8343 = n8227 & n8342 ;
  assign n8344 = ~n8339 & ~n8343 ;
  assign n8345 = ~n8337 & n8344 ;
  assign n8346 = n8333 & n8345 ;
  assign n8347 = ~n6706 & n7151 ;
  assign n8348 = ~n6706 & ~n7094 ;
  assign n8349 = n7092 & n8348 ;
  assign n8350 = ~n8347 & ~n8349 ;
  assign n8351 = n7568 & n8350 ;
  assign n8352 = ~n7746 & n8351 ;
  assign n8353 = ~n6706 & n6975 ;
  assign n8354 = ~n8349 & ~n8353 ;
  assign n8355 = ~\pi0299  & n8354 ;
  assign n8356 = n6975 & n7100 ;
  assign n8357 = ~n7094 & n7100 ;
  assign n8358 = ~n7138 & n8357 ;
  assign n8359 = ~n8356 & ~n8358 ;
  assign n8360 = n6706 & ~n8359 ;
  assign n8361 = n7551 & ~n8360 ;
  assign n8362 = n8355 & n8361 ;
  assign n8363 = ~n8352 & ~n8362 ;
  assign n8364 = ~\pi0039  & \pi0232  ;
  assign n8365 = ~n8363 & n8364 ;
  assign n8366 = \pi0232  & n7160 ;
  assign n8367 = \pi0299  & ~n8366 ;
  assign n8368 = ~\pi0232  & ~\pi0299  ;
  assign n8369 = ~n6975 & n8368 ;
  assign n8370 = ~n8367 & ~n8369 ;
  assign n8371 = n7151 & ~n8369 ;
  assign n8372 = ~n8370 & ~n8371 ;
  assign n8373 = ~n7146 & n8372 ;
  assign n8374 = ~\pi0039  & n8373 ;
  assign n8375 = n1638 & n4520 ;
  assign n8376 = \pi0038  & ~n8375 ;
  assign n8377 = \pi0299  & n6706 ;
  assign n8378 = ~n6732 & n8377 ;
  assign n8379 = \pi0299  & ~n6706 ;
  assign n8380 = ~n6713 & n8379 ;
  assign n8381 = ~n8378 & ~n8380 ;
  assign n8382 = ~n7599 & ~n8381 ;
  assign n8383 = ~\pi0299  & n6706 ;
  assign n8384 = ~n6761 & n8383 ;
  assign n8385 = ~\pi0299  & ~n6706 ;
  assign n8386 = ~n6713 & n8385 ;
  assign n8387 = ~n8384 & ~n8386 ;
  assign n8388 = ~n6957 & ~n8387 ;
  assign n8389 = \pi0039  & ~n8388 ;
  assign n8390 = ~n8382 & n8389 ;
  assign n8391 = ~n8376 & ~n8390 ;
  assign n8392 = ~n8374 & n8391 ;
  assign n8393 = ~n8365 & n8392 ;
  assign n8394 = \pi0038  & n4520 ;
  assign n8395 = n1638 & n8394 ;
  assign n8396 = ~\pi0100  & n2364 ;
  assign n8397 = ~n8395 & n8396 ;
  assign n8398 = ~n8393 & n8397 ;
  assign n8399 = ~n6798 & ~n6819 ;
  assign n8400 = n6789 & ~n8399 ;
  assign n8401 = ~\pi0038  & n6784 ;
  assign n8402 = n1266 & n8401 ;
  assign n8403 = n1354 & n8402 ;
  assign n8404 = n1358 & n8403 ;
  assign n8405 = \pi0100  & ~n8404 ;
  assign n8406 = ~\pi0087  & ~n8405 ;
  assign n8407 = ~n8400 & n8406 ;
  assign n8408 = n2364 & ~n8407 ;
  assign n8409 = n2324 & n2402 ;
  assign n8410 = n1281 & n8409 ;
  assign n8411 = n1260 & n8410 ;
  assign n8412 = \pi0054  & ~n8411 ;
  assign n8413 = n1266 & n6784 ;
  assign n8414 = n1354 & n2363 ;
  assign n8415 = n8413 & n8414 ;
  assign n8416 = n1358 & n8415 ;
  assign n8417 = \pi0075  & ~n8416 ;
  assign n8418 = n1281 & n2536 ;
  assign n8419 = n1260 & n8418 ;
  assign n8420 = \pi0092  & ~n8419 ;
  assign n8421 = ~n8417 & ~n8420 ;
  assign n8422 = ~n8412 & n8421 ;
  assign n8423 = ~n8408 & n8422 ;
  assign n8424 = ~n8398 & n8423 ;
  assign n8425 = \pi0054  & n8409 ;
  assign n8426 = n1281 & n8425 ;
  assign n8427 = n1260 & n8426 ;
  assign n8428 = n2404 & ~n8427 ;
  assign n8429 = ~n8424 & n8428 ;
  assign n8430 = n1638 & n6630 ;
  assign n8431 = ~\pi0055  & \pi0074  ;
  assign n8432 = ~n8430 & n8431 ;
  assign n8433 = ~\pi0056  & ~\pi0074  ;
  assign n8434 = n6630 & n8433 ;
  assign n8435 = n1638 & n8434 ;
  assign n8436 = ~n2423 & ~n8435 ;
  assign n8437 = ~\pi0055  & n6622 ;
  assign n8438 = n1291 & n8437 ;
  assign n8439 = n1281 & n8438 ;
  assign n8440 = n1260 & n8439 ;
  assign n8441 = ~n2467 & ~n8440 ;
  assign n8442 = ~\pi0062  & ~n8441 ;
  assign n8443 = ~n8436 & n8442 ;
  assign n8444 = ~n8432 & n8443 ;
  assign n8445 = ~n8429 & n8444 ;
  assign n8446 = ~n2467 & n8438 ;
  assign n8447 = n1281 & n8446 ;
  assign n8448 = n1260 & n8447 ;
  assign n8449 = ~\pi0954  & ~n8448 ;
  assign n8450 = ~n8445 & n8449 ;
  assign n8451 = \pi0024  & \pi0954  ;
  assign n8452 = ~n8450 & ~n8451 ;
  assign n8453 = ~\pi0100  & ~\pi0228  ;
  assign n8454 = ~n1639 & n8453 ;
  assign n8455 = ~n2591 & n8454 ;
  assign n8456 = ~n2581 & n8455 ;
  assign n8457 = \pi0299  & n2618 ;
  assign n8458 = \pi0299  & ~n2609 ;
  assign n8459 = n2614 & n8458 ;
  assign n8460 = ~n8457 & ~n8459 ;
  assign n8461 = n1281 & n7228 ;
  assign n8462 = n1260 & n8461 ;
  assign n8463 = ~\pi0299  & ~n8462 ;
  assign n8464 = \pi0100  & ~\pi0228  ;
  assign n8465 = n1281 & n8464 ;
  assign n8466 = n1260 & n8465 ;
  assign n8467 = ~n8463 & n8466 ;
  assign n8468 = n8460 & n8467 ;
  assign n8469 = ~\pi0039  & ~n1209 ;
  assign n8470 = ~n8468 & n8469 ;
  assign n8471 = ~n8456 & n8470 ;
  assign n8472 = \pi0038  & ~n1209 ;
  assign n8473 = n1281 & n8453 ;
  assign n8474 = n1260 & n8473 ;
  assign n8475 = \pi0039  & ~n1209 ;
  assign n8476 = ~n8474 & n8475 ;
  assign n8477 = ~n8472 & ~n8476 ;
  assign n8478 = \pi0075  & ~n1209 ;
  assign n8479 = n4539 & ~n8478 ;
  assign n8480 = n8477 & n8479 ;
  assign n8481 = ~n8471 & n8480 ;
  assign n8482 = ~\pi0228  & n2402 ;
  assign n8483 = n1281 & n8482 ;
  assign n8484 = n1260 & n8483 ;
  assign n8485 = ~\pi0075  & ~n1209 ;
  assign n8486 = ~n8484 & n8485 ;
  assign n8487 = ~\pi0092  & ~n8478 ;
  assign n8488 = ~n1286 & n8487 ;
  assign n8489 = ~n8486 & n8488 ;
  assign n8490 = ~\pi0056  & ~n1209 ;
  assign n8491 = ~n2423 & ~n8490 ;
  assign n8492 = ~\pi0075  & n2362 ;
  assign n8493 = n1259 & n8492 ;
  assign n8494 = n1249 & n8493 ;
  assign n8495 = n6858 & n8494 ;
  assign n8496 = ~\pi0074  & n1285 ;
  assign n8497 = ~n2423 & n8496 ;
  assign n8498 = n8495 & n8497 ;
  assign n8499 = ~n8491 & ~n8498 ;
  assign n8500 = ~\pi0092  & n2511 ;
  assign n8501 = ~n1209 & n2511 ;
  assign n8502 = ~n8495 & n8501 ;
  assign n8503 = ~n8500 & ~n8502 ;
  assign n8504 = n8499 & ~n8503 ;
  assign n8505 = ~n8489 & n8504 ;
  assign n8506 = ~n8481 & n8505 ;
  assign n8507 = ~n1209 & ~n2511 ;
  assign n8508 = ~\pi0055  & ~n8507 ;
  assign n8509 = n8499 & ~n8508 ;
  assign n8510 = ~\pi0228  & n2404 ;
  assign n8511 = n2403 & n8510 ;
  assign n8512 = n1281 & n8511 ;
  assign n8513 = n1260 & n8512 ;
  assign n8514 = \pi0056  & ~n1209 ;
  assign n8515 = ~n8513 & n8514 ;
  assign n8516 = ~\pi0062  & n2467 ;
  assign n8517 = ~n8515 & n8516 ;
  assign n8518 = ~n8509 & n8517 ;
  assign n8519 = ~n8506 & n8518 ;
  assign n8520 = ~\pi0228  & n2504 ;
  assign n8521 = n1281 & n8520 ;
  assign n8522 = n1260 & n8521 ;
  assign n8523 = ~n1209 & ~n8522 ;
  assign n8524 = \pi0062  & n2467 ;
  assign n8525 = ~n8523 & n8524 ;
  assign n8526 = n1209 & ~n2467 ;
  assign n8527 = ~n8525 & ~n8526 ;
  assign n8528 = ~n8519 & n8527 ;
  assign n8529 = ~\pi0228  & \pi0252  ;
  assign n8530 = ~\pi0119  & ~n8529 ;
  assign n8531 = \pi0119  & \pi1056  ;
  assign n8532 = ~\pi0468  & ~n8531 ;
  assign n8533 = ~n8530 & n8532 ;
  assign n8534 = \pi0119  & \pi1077  ;
  assign n8535 = ~\pi0468  & ~n8534 ;
  assign n8536 = ~n8530 & n8535 ;
  assign n8537 = \pi0119  & \pi1073  ;
  assign n8538 = ~\pi0468  & ~n8537 ;
  assign n8539 = ~n8530 & n8538 ;
  assign n8540 = \pi0119  & \pi1041  ;
  assign n8541 = ~\pi0468  & ~n8540 ;
  assign n8542 = ~n8530 & n8541 ;
  assign n8543 = ~\pi1091  & \pi1093  ;
  assign n8544 = ~\pi0122  & \pi0567  ;
  assign n8545 = n8543 & n8544 ;
  assign n8546 = ~\pi0098  & \pi0824  ;
  assign n8547 = n6809 & n8546 ;
  assign n8548 = n8545 & n8547 ;
  assign n8549 = ~n8496 & n8548 ;
  assign n8550 = ~\pi0841  & n6967 ;
  assign n8551 = n1354 & n8550 ;
  assign n8552 = n1358 & n8551 ;
  assign n8553 = \pi0096  & n2575 ;
  assign n8554 = n8552 & n8553 ;
  assign n8555 = ~\pi0093  & n1321 ;
  assign n8556 = ~\pi0841  & n1321 ;
  assign n8557 = n1829 & n8556 ;
  assign n8558 = n1358 & n8557 ;
  assign n8559 = ~n8555 & ~n8558 ;
  assign n8560 = ~\pi0109  & ~\pi0841  ;
  assign n8561 = \pi0090  & n8560 ;
  assign n8562 = n1327 & n8561 ;
  assign n8563 = n1319 & n8562 ;
  assign n8564 = ~\pi0093  & ~n8563 ;
  assign n8565 = ~n8559 & ~n8564 ;
  assign n8566 = n1269 & n1270 ;
  assign n8567 = ~\pi0047  & n1326 ;
  assign n8568 = n1322 & n8567 ;
  assign n8569 = n8566 & n8568 ;
  assign n8570 = \pi0097  & n8569 ;
  assign n8571 = ~\pi0088  & \pi0098  ;
  assign n8572 = n1252 & n8571 ;
  assign n8573 = n1276 & n8572 ;
  assign n8574 = n8569 & n8573 ;
  assign n8575 = n1542 & n8574 ;
  assign n8576 = ~n8570 & ~n8575 ;
  assign n8577 = ~\pi0051  & n8576 ;
  assign n8578 = ~n8565 & n8577 ;
  assign n8579 = n1321 & n1354 ;
  assign n8580 = n1358 & n8579 ;
  assign n8581 = \pi0051  & ~n8580 ;
  assign n8582 = \pi0096  & ~n8552 ;
  assign n8583 = n2575 & ~n8582 ;
  assign n8584 = ~n8581 & n8583 ;
  assign n8585 = ~n8578 & n8584 ;
  assign n8586 = ~n8554 & ~n8585 ;
  assign n8587 = ~\pi0122  & \pi0829  ;
  assign n8588 = n6809 & n8587 ;
  assign n8589 = ~\pi0072  & ~\pi1093  ;
  assign n8590 = n8588 & n8589 ;
  assign n8591 = ~n8586 & n8590 ;
  assign n8592 = n1263 & n1264 ;
  assign n8593 = ~n8581 & n8592 ;
  assign n8594 = n6811 & ~n8587 ;
  assign n8595 = ~\pi1093  & n8594 ;
  assign n8596 = n8593 & n8595 ;
  assign n8597 = ~n8578 & n8596 ;
  assign n8598 = ~\pi0087  & ~\pi0567  ;
  assign n8599 = ~n8597 & n8598 ;
  assign n8600 = ~n8591 & n8599 ;
  assign n8601 = ~\pi0075  & ~\pi0100  ;
  assign n8602 = n1288 & n8601 ;
  assign n8603 = ~\pi0567  & ~n8602 ;
  assign n8604 = ~\pi1093  & n6811 ;
  assign n8605 = n1281 & n8604 ;
  assign n8606 = n1260 & n8605 ;
  assign n8607 = \pi0087  & ~\pi0567  ;
  assign n8608 = ~n8606 & n8607 ;
  assign n8609 = ~n8603 & ~n8608 ;
  assign n8610 = n8496 & n8609 ;
  assign n8611 = ~n8600 & n8610 ;
  assign n8612 = ~n8549 & ~n8611 ;
  assign n8613 = \pi0592  & n8612 ;
  assign n8614 = \pi0122  & \pi0824  ;
  assign n8615 = n6809 & n8614 ;
  assign n8616 = n1281 & n8615 ;
  assign n8617 = n1260 & n8616 ;
  assign n8618 = ~\pi0122  & n8547 ;
  assign n8619 = ~n8617 & ~n8618 ;
  assign n8620 = \pi1093  & ~n8619 ;
  assign n8621 = ~\pi0122  & n8543 ;
  assign n8622 = n8547 & n8621 ;
  assign n8623 = ~\pi1091  & ~n8622 ;
  assign n8624 = ~n8606 & n8623 ;
  assign n8625 = ~n8620 & n8624 ;
  assign n8626 = ~n2328 & ~n8622 ;
  assign n8627 = \pi1093  & n1686 ;
  assign n8628 = n6811 & ~n8627 ;
  assign n8629 = n1281 & n8628 ;
  assign n8630 = n1260 & n8629 ;
  assign n8631 = \pi1091  & ~n8622 ;
  assign n8632 = ~n8630 & n8631 ;
  assign n8633 = ~n8626 & ~n8632 ;
  assign n8634 = \pi0087  & n8633 ;
  assign n8635 = ~n8625 & n8634 ;
  assign n8636 = ~\pi0075  & ~n8635 ;
  assign n8637 = ~\pi0299  & ~n2167 ;
  assign n8638 = \pi0299  & ~n1801 ;
  assign n8639 = ~n8637 & ~n8638 ;
  assign n8640 = \pi0232  & n6706 ;
  assign n8641 = n8639 & n8640 ;
  assign n8642 = ~\pi0122  & \pi1093  ;
  assign n8643 = n8547 & n8642 ;
  assign n8644 = ~\pi1091  & ~n8643 ;
  assign n8645 = n2342 & ~n8644 ;
  assign n8646 = ~n8641 & n8645 ;
  assign n8647 = ~\pi1091  & n8646 ;
  assign n8648 = \pi1093  & ~n1686 ;
  assign n8649 = ~\pi0024  & n8588 ;
  assign n8650 = n8648 & n8649 ;
  assign n8651 = ~n6808 & n8650 ;
  assign n8652 = n8646 & n8651 ;
  assign n8653 = n7207 & n8652 ;
  assign n8654 = ~n8647 & ~n8653 ;
  assign n8655 = n8622 & n8640 ;
  assign n8656 = n8639 & n8655 ;
  assign n8657 = ~n2342 & n8622 ;
  assign n8658 = \pi0075  & ~n8657 ;
  assign n8659 = ~n8656 & n8658 ;
  assign n8660 = n8654 & n8659 ;
  assign n8661 = ~n8636 & ~n8660 ;
  assign n8662 = n8588 & n8648 ;
  assign n8663 = ~n6808 & n8662 ;
  assign n8664 = n1281 & n8663 ;
  assign n8665 = n1260 & n8664 ;
  assign n8666 = \pi0228  & n1288 ;
  assign n8667 = \pi1091  & n8666 ;
  assign n8668 = ~n8641 & n8667 ;
  assign n8669 = n8665 & n8668 ;
  assign n8670 = \pi0100  & ~n8622 ;
  assign n8671 = ~n8669 & n8670 ;
  assign n8672 = ~\pi0087  & ~n8671 ;
  assign n8673 = ~n8660 & n8672 ;
  assign n8674 = ~n8661 & ~n8673 ;
  assign n8675 = \pi0829  & n6809 ;
  assign n8676 = n8648 & n8675 ;
  assign n8677 = n1259 & n8676 ;
  assign n8678 = n1249 & n8677 ;
  assign n8679 = n6920 & n8678 ;
  assign n8680 = \pi1091  & ~n8679 ;
  assign n8681 = \pi1091  & ~n6709 ;
  assign n8682 = n6735 & n8681 ;
  assign n8683 = ~n8644 & ~n8682 ;
  assign n8684 = ~\pi0216  & n6936 ;
  assign n8685 = ~n6732 & n8684 ;
  assign n8686 = n8683 & n8685 ;
  assign n8687 = ~n8680 & n8686 ;
  assign n8688 = \pi1091  & ~n6714 ;
  assign n8689 = n6732 & n8684 ;
  assign n8690 = ~n8644 & n8689 ;
  assign n8691 = ~n8688 & n8690 ;
  assign n8692 = ~n8680 & n8691 ;
  assign n8693 = ~n8687 & ~n8692 ;
  assign n8694 = ~\pi0122  & \pi0824  ;
  assign n8695 = n6809 & n8694 ;
  assign n8696 = n8543 & n8695 ;
  assign n8697 = ~\pi0098  & ~n8684 ;
  assign n8698 = n8696 & n8697 ;
  assign n8699 = \pi0299  & ~n8698 ;
  assign n8700 = n8693 & n8699 ;
  assign n8701 = ~\pi0223  & n6148 ;
  assign n8702 = ~n6761 & n8701 ;
  assign n8703 = n8683 & n8702 ;
  assign n8704 = ~n8680 & n8703 ;
  assign n8705 = n6761 & n8701 ;
  assign n8706 = ~n8644 & n8705 ;
  assign n8707 = ~n8688 & n8706 ;
  assign n8708 = ~n8680 & n8707 ;
  assign n8709 = ~n8704 & ~n8708 ;
  assign n8710 = ~\pi0098  & ~n8701 ;
  assign n8711 = n8696 & n8710 ;
  assign n8712 = ~\pi0299  & ~n8711 ;
  assign n8713 = n8709 & n8712 ;
  assign n8714 = ~n8700 & ~n8713 ;
  assign n8715 = \pi0039  & n8714 ;
  assign n8716 = ~\pi0038  & n8715 ;
  assign n8717 = ~n8591 & ~n8597 ;
  assign n8718 = ~\pi1091  & ~\pi1093  ;
  assign n8719 = ~\pi0051  & ~n8565 ;
  assign n8720 = n8593 & n8615 ;
  assign n8721 = ~n8719 & n8720 ;
  assign n8722 = ~\pi1091  & ~n8618 ;
  assign n8723 = ~n8721 & n8722 ;
  assign n8724 = ~n8718 & ~n8723 ;
  assign n8725 = n8717 & ~n8724 ;
  assign n8726 = ~\pi0039  & ~n8725 ;
  assign n8727 = ~\pi0024  & n1325 ;
  assign n8728 = n1398 & n8727 ;
  assign n8729 = n1319 & n8728 ;
  assign n8730 = ~\pi0046  & \pi0097  ;
  assign n8731 = n7114 & n8730 ;
  assign n8732 = n1675 & n8731 ;
  assign n8733 = n1542 & n8732 ;
  assign n8734 = ~\pi0091  & n8733 ;
  assign n8735 = ~n8729 & ~n8734 ;
  assign n8736 = n1277 & ~n8559 ;
  assign n8737 = ~n8735 & n8736 ;
  assign n8738 = n8719 & ~n8737 ;
  assign n8739 = \pi0829  & \pi1092  ;
  assign n8740 = \pi0950  & n1329 ;
  assign n8741 = n1264 & n8740 ;
  assign n8742 = ~n8582 & n8741 ;
  assign n8743 = n8739 & n8742 ;
  assign n8744 = ~n8581 & n8743 ;
  assign n8745 = ~n8738 & n8744 ;
  assign n8746 = \pi0096  & n8739 ;
  assign n8747 = n8742 & n8746 ;
  assign n8748 = \pi0122  & n6811 ;
  assign n8749 = n8592 & n8748 ;
  assign n8750 = ~n8581 & n8749 ;
  assign n8751 = \pi0824  & ~\pi0829  ;
  assign n8752 = n6809 & n8751 ;
  assign n8753 = n8592 & n8752 ;
  assign n8754 = ~n8581 & n8753 ;
  assign n8755 = ~n8750 & ~n8754 ;
  assign n8756 = ~n8719 & ~n8755 ;
  assign n8757 = ~n8747 & ~n8756 ;
  assign n8758 = ~n8745 & n8757 ;
  assign n8759 = \pi0122  & ~n8750 ;
  assign n8760 = ~\pi0051  & \pi0122  ;
  assign n8761 = ~n8565 & n8760 ;
  assign n8762 = ~n8759 & ~n8761 ;
  assign n8763 = n8648 & n8762 ;
  assign n8764 = ~n8758 & n8763 ;
  assign n8765 = \pi1091  & ~n8597 ;
  assign n8766 = ~n8591 & n8765 ;
  assign n8767 = ~n8764 & n8766 ;
  assign n8768 = ~\pi0038  & ~n8767 ;
  assign n8769 = n8726 & n8768 ;
  assign n8770 = ~n8716 & ~n8769 ;
  assign n8771 = \pi0038  & ~\pi0098  ;
  assign n8772 = n8543 & n8771 ;
  assign n8773 = n8695 & n8772 ;
  assign n8774 = ~\pi0100  & ~n8773 ;
  assign n8775 = ~n8661 & n8774 ;
  assign n8776 = n8770 & n8775 ;
  assign n8777 = ~n8674 & ~n8776 ;
  assign n8778 = \pi0567  & ~n8549 ;
  assign n8779 = \pi0592  & n8778 ;
  assign n8780 = ~n8777 & n8779 ;
  assign n8781 = ~n8613 & ~n8780 ;
  assign n8782 = ~n1686 & n6703 ;
  assign n8783 = n8762 & n8782 ;
  assign n8784 = ~n8758 & n8783 ;
  assign n8785 = n2320 & ~n8597 ;
  assign n8786 = ~n8591 & n8785 ;
  assign n8787 = ~n8784 & n8786 ;
  assign n8788 = n1259 & n1696 ;
  assign n8789 = n1249 & n8788 ;
  assign n8790 = n6920 & n8789 ;
  assign n8791 = ~n8381 & n8684 ;
  assign n8792 = ~n8387 & n8701 ;
  assign n8793 = ~n8791 & ~n8792 ;
  assign n8794 = ~\pi0038  & ~n8793 ;
  assign n8795 = n8790 & n8794 ;
  assign n8796 = n3688 & ~n8795 ;
  assign n8797 = n2342 & ~n8641 ;
  assign n8798 = ~\pi0024  & \pi1093  ;
  assign n8799 = \pi1091  & ~n1686 ;
  assign n8800 = n8588 & n8799 ;
  assign n8801 = ~n6808 & n8800 ;
  assign n8802 = n8798 & n8801 ;
  assign n8803 = n8797 & n8802 ;
  assign n8804 = n7207 & n8803 ;
  assign n8805 = \pi0075  & ~n8804 ;
  assign n8806 = ~\pi0087  & n8668 ;
  assign n8807 = n8665 & n8806 ;
  assign n8808 = ~n2362 & ~n8807 ;
  assign n8809 = ~n8805 & ~n8808 ;
  assign n8810 = ~n8796 & n8809 ;
  assign n8811 = ~n8787 & n8810 ;
  assign n8812 = ~\pi0039  & \pi0087  ;
  assign n8813 = n2327 & n8812 ;
  assign n8814 = ~\pi1091  & n8813 ;
  assign n8815 = n8604 & n8814 ;
  assign n8816 = n1281 & n8815 ;
  assign n8817 = n1260 & n8816 ;
  assign n8818 = \pi1091  & n8813 ;
  assign n8819 = n8628 & n8818 ;
  assign n8820 = n1281 & n8819 ;
  assign n8821 = n1260 & n8820 ;
  assign n8822 = ~\pi0075  & ~n8821 ;
  assign n8823 = ~n8817 & n8822 ;
  assign n8824 = ~n8805 & ~n8823 ;
  assign n8825 = \pi0567  & ~n8824 ;
  assign n8826 = ~n8811 & n8825 ;
  assign n8827 = n8611 & ~n8826 ;
  assign n8828 = ~\pi0592  & ~n8827 ;
  assign n8829 = n8781 & ~n8828 ;
  assign n8830 = \pi0351  & \pi1199  ;
  assign n8831 = \pi0461  & n8830 ;
  assign n8832 = ~n8829 & n8831 ;
  assign n8833 = ~\pi0323  & ~\pi0346  ;
  assign n8834 = \pi0323  & \pi0346  ;
  assign n8835 = ~n8833 & ~n8834 ;
  assign n8836 = \pi0450  & n8835 ;
  assign n8837 = ~\pi0450  & ~n8835 ;
  assign n8838 = ~n8836 & ~n8837 ;
  assign n8839 = \pi0345  & ~\pi0358  ;
  assign n8840 = ~\pi0345  & \pi0358  ;
  assign n8841 = ~n8839 & ~n8840 ;
  assign n8842 = n8838 & n8841 ;
  assign n8843 = ~n8838 & ~n8841 ;
  assign n8844 = ~n8842 & ~n8843 ;
  assign n8845 = ~\pi0327  & ~\pi0362  ;
  assign n8846 = \pi0327  & \pi0362  ;
  assign n8847 = ~n8845 & ~n8846 ;
  assign n8848 = \pi0343  & ~\pi0344  ;
  assign n8849 = ~\pi0343  & \pi0344  ;
  assign n8850 = ~n8848 & ~n8849 ;
  assign n8851 = n8847 & n8850 ;
  assign n8852 = ~n8847 & ~n8850 ;
  assign n8853 = ~n8851 & ~n8852 ;
  assign n8854 = n8844 & n8853 ;
  assign n8855 = \pi1197  & n8841 ;
  assign n8856 = ~n8838 & n8855 ;
  assign n8857 = \pi1197  & n8853 ;
  assign n8858 = \pi1197  & ~n8841 ;
  assign n8859 = n8838 & n8858 ;
  assign n8860 = ~n8857 & ~n8859 ;
  assign n8861 = ~n8856 & n8860 ;
  assign n8862 = ~n8854 & ~n8861 ;
  assign n8863 = ~\pi0342  & ~\pi0460  ;
  assign n8864 = \pi0342  & \pi0460  ;
  assign n8865 = ~n8863 & ~n8864 ;
  assign n8866 = \pi0361  & n8865 ;
  assign n8867 = ~\pi0361  & ~n8865 ;
  assign n8868 = ~n8866 & ~n8867 ;
  assign n8869 = \pi0320  & ~\pi0441  ;
  assign n8870 = ~\pi0320  & \pi0441  ;
  assign n8871 = ~n8869 & ~n8870 ;
  assign n8872 = \pi0355  & ~\pi0458  ;
  assign n8873 = ~\pi0355  & \pi0458  ;
  assign n8874 = ~n8872 & ~n8873 ;
  assign n8875 = \pi0452  & ~\pi0455  ;
  assign n8876 = ~\pi0452  & \pi0455  ;
  assign n8877 = ~n8875 & ~n8876 ;
  assign n8878 = ~n8874 & n8877 ;
  assign n8879 = ~n8871 & n8878 ;
  assign n8880 = ~n8868 & n8879 ;
  assign n8881 = ~n8874 & ~n8877 ;
  assign n8882 = n8871 & n8881 ;
  assign n8883 = ~n8868 & n8882 ;
  assign n8884 = ~n8880 & ~n8883 ;
  assign n8885 = ~n8871 & n8881 ;
  assign n8886 = n8868 & n8885 ;
  assign n8887 = n8871 & n8878 ;
  assign n8888 = n8868 & n8887 ;
  assign n8889 = ~n8886 & ~n8888 ;
  assign n8890 = n8884 & n8889 ;
  assign n8891 = n8874 & n8877 ;
  assign n8892 = ~n8871 & n8891 ;
  assign n8893 = n8868 & n8892 ;
  assign n8894 = n8874 & ~n8877 ;
  assign n8895 = n8871 & n8894 ;
  assign n8896 = n8868 & n8895 ;
  assign n8897 = ~n8893 & ~n8896 ;
  assign n8898 = ~n8871 & n8894 ;
  assign n8899 = ~n8868 & n8898 ;
  assign n8900 = n8871 & n8891 ;
  assign n8901 = ~n8868 & n8900 ;
  assign n8902 = ~n8899 & ~n8901 ;
  assign n8903 = n8897 & n8902 ;
  assign n8904 = n8890 & n8903 ;
  assign n8905 = \pi1196  & n8904 ;
  assign n8906 = ~n8862 & ~n8905 ;
  assign n8907 = \pi0592  & ~n8906 ;
  assign n8908 = n8611 & ~n8906 ;
  assign n8909 = ~n8826 & n8908 ;
  assign n8910 = ~n8907 & ~n8909 ;
  assign n8911 = n8781 & ~n8910 ;
  assign n8912 = ~\pi0347  & ~\pi0359  ;
  assign n8913 = \pi0347  & \pi0359  ;
  assign n8914 = ~n8912 & ~n8913 ;
  assign n8915 = \pi0315  & ~\pi0322  ;
  assign n8916 = ~\pi0315  & \pi0322  ;
  assign n8917 = ~n8915 & ~n8916 ;
  assign n8918 = ~\pi0321  & n8917 ;
  assign n8919 = \pi0321  & ~n8917 ;
  assign n8920 = ~n8918 & ~n8919 ;
  assign n8921 = ~n8914 & ~n8920 ;
  assign n8922 = n8914 & n8920 ;
  assign n8923 = ~n8921 & ~n8922 ;
  assign n8924 = \pi0316  & ~\pi0348  ;
  assign n8925 = ~\pi0316  & \pi0348  ;
  assign n8926 = ~n8924 & ~n8925 ;
  assign n8927 = ~\pi0349  & ~\pi0350  ;
  assign n8928 = \pi0349  & \pi0350  ;
  assign n8929 = ~n8927 & ~n8928 ;
  assign n8930 = ~n8926 & ~n8929 ;
  assign n8931 = n8926 & n8929 ;
  assign n8932 = ~n8930 & ~n8931 ;
  assign n8933 = ~\pi0592  & \pi1198  ;
  assign n8934 = ~n8932 & n8933 ;
  assign n8935 = ~n8923 & n8934 ;
  assign n8936 = n8932 & n8933 ;
  assign n8937 = n8923 & n8936 ;
  assign n8938 = ~n8935 & ~n8937 ;
  assign n8939 = n8906 & n8938 ;
  assign n8940 = n8611 & n8906 ;
  assign n8941 = ~n8826 & n8940 ;
  assign n8942 = ~n8939 & ~n8941 ;
  assign n8943 = n8612 & n8938 ;
  assign n8944 = n8778 & n8938 ;
  assign n8945 = ~n8777 & n8944 ;
  assign n8946 = ~n8943 & ~n8945 ;
  assign n8947 = ~n8942 & n8946 ;
  assign n8948 = ~n8911 & ~n8947 ;
  assign n8949 = \pi0461  & ~n8830 ;
  assign n8950 = n8948 & n8949 ;
  assign n8951 = ~n8832 & ~n8950 ;
  assign n8952 = ~\pi0351  & \pi1199  ;
  assign n8953 = ~\pi0461  & ~n8952 ;
  assign n8954 = n8948 & n8953 ;
  assign n8955 = ~\pi0461  & n8952 ;
  assign n8956 = ~n8829 & n8955 ;
  assign n8957 = ~\pi0352  & ~\pi0353  ;
  assign n8958 = \pi0352  & \pi0353  ;
  assign n8959 = ~n8957 & ~n8958 ;
  assign n8960 = ~\pi0360  & ~\pi0462  ;
  assign n8961 = \pi0360  & \pi0462  ;
  assign n8962 = ~n8960 & ~n8961 ;
  assign n8963 = ~n8959 & ~n8962 ;
  assign n8964 = n8959 & n8962 ;
  assign n8965 = ~n8963 & ~n8964 ;
  assign n8966 = \pi0354  & ~\pi0356  ;
  assign n8967 = ~\pi0354  & \pi0356  ;
  assign n8968 = ~n8966 & ~n8967 ;
  assign n8969 = \pi0357  & ~n8968 ;
  assign n8970 = n8965 & n8969 ;
  assign n8971 = \pi0357  & n8968 ;
  assign n8972 = ~n8965 & n8971 ;
  assign n8973 = ~n8970 & ~n8972 ;
  assign n8974 = ~n8956 & ~n8973 ;
  assign n8975 = ~n8954 & n8974 ;
  assign n8976 = n8951 & n8975 ;
  assign n8977 = ~\pi0357  & ~n8968 ;
  assign n8978 = ~n8965 & n8977 ;
  assign n8979 = ~\pi0357  & n8968 ;
  assign n8980 = n8965 & n8979 ;
  assign n8981 = ~n8978 & ~n8980 ;
  assign n8982 = ~n8956 & ~n8981 ;
  assign n8983 = ~n8954 & n8982 ;
  assign n8984 = n8951 & n8983 ;
  assign n8985 = ~\pi0591  & ~n8984 ;
  assign n8986 = ~\pi0461  & ~n8830 ;
  assign n8987 = n8948 & n8986 ;
  assign n8988 = ~\pi0461  & n8830 ;
  assign n8989 = ~n8829 & n8988 ;
  assign n8990 = \pi0461  & n8952 ;
  assign n8991 = ~n8829 & n8990 ;
  assign n8992 = ~n8989 & ~n8991 ;
  assign n8993 = ~n8987 & n8992 ;
  assign n8994 = \pi0461  & ~n8952 ;
  assign n8995 = n8948 & n8994 ;
  assign n8996 = n8965 & n8977 ;
  assign n8997 = ~n8965 & n8979 ;
  assign n8998 = ~n8996 & ~n8997 ;
  assign n8999 = ~n8995 & ~n8998 ;
  assign n9000 = n8993 & n8999 ;
  assign n9001 = ~n8965 & n8969 ;
  assign n9002 = n8965 & n8971 ;
  assign n9003 = ~n9001 & ~n9002 ;
  assign n9004 = ~n8995 & ~n9003 ;
  assign n9005 = n8993 & n9004 ;
  assign n9006 = ~n9000 & ~n9005 ;
  assign n9007 = n8985 & n9006 ;
  assign n9008 = ~n8976 & n9007 ;
  assign n9009 = \pi0075  & ~\pi1196  ;
  assign n9010 = ~\pi0087  & \pi0100  ;
  assign n9011 = ~n8669 & n9010 ;
  assign n9012 = \pi0824  & n6809 ;
  assign n9013 = n8592 & n9012 ;
  assign n9014 = ~n8581 & n9013 ;
  assign n9015 = ~n8719 & n9014 ;
  assign n9016 = \pi1093  & n1288 ;
  assign n9017 = \pi1093  & n8790 ;
  assign n9018 = n8794 & n9017 ;
  assign n9019 = ~n9016 & ~n9018 ;
  assign n9020 = n9015 & ~n9019 ;
  assign n9021 = n8763 & n9020 ;
  assign n9022 = ~n8758 & n9021 ;
  assign n9023 = ~\pi1091  & ~n9019 ;
  assign n9024 = n9015 & n9023 ;
  assign n9025 = ~\pi0087  & ~n9024 ;
  assign n9026 = ~n9022 & n9025 ;
  assign n9027 = ~n9011 & ~n9026 ;
  assign n9028 = ~n8796 & ~n9011 ;
  assign n9029 = ~n8787 & n9028 ;
  assign n9030 = ~n9027 & ~n9029 ;
  assign n9031 = ~n8543 & n8628 ;
  assign n9032 = n1281 & n9031 ;
  assign n9033 = n1260 & n9032 ;
  assign n9034 = n2328 & n9033 ;
  assign n9035 = n1281 & n9012 ;
  assign n9036 = n2328 & n8543 ;
  assign n9037 = n1259 & n9036 ;
  assign n9038 = n1249 & n9037 ;
  assign n9039 = n9035 & n9038 ;
  assign n9040 = \pi0087  & ~n9039 ;
  assign n9041 = ~n9034 & n9040 ;
  assign n9042 = ~\pi1196  & ~n9041 ;
  assign n9043 = ~n9030 & n9042 ;
  assign n9044 = ~n9009 & ~n9043 ;
  assign n9045 = ~\pi0075  & ~\pi0592  ;
  assign n9046 = ~n8543 & ~n8630 ;
  assign n9047 = n8813 & ~n9046 ;
  assign n9048 = n1260 & n9035 ;
  assign n9049 = n8543 & ~n9048 ;
  assign n9050 = ~\pi0324  & ~\pi0410  ;
  assign n9051 = \pi0324  & \pi0410  ;
  assign n9052 = ~n9050 & ~n9051 ;
  assign n9053 = \pi0319  & ~\pi0404  ;
  assign n9054 = ~\pi0319  & \pi0404  ;
  assign n9055 = ~n9053 & ~n9054 ;
  assign n9056 = ~\pi0390  & n9055 ;
  assign n9057 = \pi0390  & ~n9055 ;
  assign n9058 = ~n9056 & ~n9057 ;
  assign n9059 = ~n9052 & ~n9058 ;
  assign n9060 = n9052 & n9058 ;
  assign n9061 = ~n9059 & ~n9060 ;
  assign n9062 = \pi0411  & ~\pi0412  ;
  assign n9063 = ~\pi0411  & \pi0412  ;
  assign n9064 = ~n9062 & ~n9063 ;
  assign n9065 = ~\pi0397  & ~\pi0456  ;
  assign n9066 = \pi0397  & \pi0456  ;
  assign n9067 = ~n9065 & ~n9066 ;
  assign n9068 = ~n9064 & ~n9067 ;
  assign n9069 = n9064 & n9067 ;
  assign n9070 = ~n9068 & ~n9069 ;
  assign n9071 = n8543 & ~n9070 ;
  assign n9072 = ~n9061 & n9071 ;
  assign n9073 = n8543 & n9070 ;
  assign n9074 = n9061 & n9073 ;
  assign n9075 = ~n9072 & ~n9074 ;
  assign n9076 = ~n9049 & n9075 ;
  assign n9077 = n9047 & n9076 ;
  assign n9078 = n9045 & ~n9077 ;
  assign n9079 = \pi1196  & ~n9078 ;
  assign n9080 = ~n8787 & ~n8796 ;
  assign n9081 = n9061 & ~n9070 ;
  assign n9082 = ~n9061 & n9070 ;
  assign n9083 = ~n9081 & ~n9082 ;
  assign n9084 = ~n9022 & ~n9024 ;
  assign n9085 = ~n9083 & ~n9084 ;
  assign n9086 = ~n9080 & ~n9085 ;
  assign n9087 = \pi1196  & ~n8808 ;
  assign n9088 = ~n9086 & n9087 ;
  assign n9089 = ~n9079 & ~n9088 ;
  assign n9090 = n9044 & n9089 ;
  assign n9091 = ~\pi1199  & n9090 ;
  assign n9092 = ~\pi0318  & ~\pi0403  ;
  assign n9093 = \pi0318  & \pi0403  ;
  assign n9094 = ~n9092 & ~n9093 ;
  assign n9095 = \pi0402  & ~\pi0406  ;
  assign n9096 = ~\pi0402  & \pi0406  ;
  assign n9097 = ~n9095 & ~n9096 ;
  assign n9098 = ~\pi0401  & n9097 ;
  assign n9099 = \pi0401  & ~n9097 ;
  assign n9100 = ~n9098 & ~n9099 ;
  assign n9101 = ~n9094 & ~n9100 ;
  assign n9102 = n9094 & n9100 ;
  assign n9103 = ~n9101 & ~n9102 ;
  assign n9104 = \pi0325  & ~\pi0405  ;
  assign n9105 = ~\pi0325  & \pi0405  ;
  assign n9106 = ~n9104 & ~n9105 ;
  assign n9107 = ~\pi0326  & ~\pi0409  ;
  assign n9108 = \pi0326  & \pi0409  ;
  assign n9109 = ~n9107 & ~n9108 ;
  assign n9110 = ~n9106 & ~n9109 ;
  assign n9111 = n9106 & n9109 ;
  assign n9112 = ~n9110 & ~n9111 ;
  assign n9113 = n9103 & ~n9112 ;
  assign n9114 = ~n9103 & n9112 ;
  assign n9115 = ~n9113 & ~n9114 ;
  assign n9116 = ~\pi0075  & \pi1196  ;
  assign n9117 = ~n9070 & n9116 ;
  assign n9118 = ~n9061 & n9117 ;
  assign n9119 = n9070 & n9116 ;
  assign n9120 = n9061 & n9119 ;
  assign n9121 = ~n9118 & ~n9120 ;
  assign n9122 = ~n9115 & n9121 ;
  assign n9123 = ~n9084 & n9122 ;
  assign n9124 = \pi1199  & n9045 ;
  assign n9125 = ~n8813 & n9124 ;
  assign n9126 = ~n8543 & n9124 ;
  assign n9127 = ~n8630 & n9126 ;
  assign n9128 = ~n9125 & ~n9127 ;
  assign n9129 = \pi1196  & ~n9070 ;
  assign n9130 = ~n9061 & n9129 ;
  assign n9131 = \pi1196  & n9070 ;
  assign n9132 = n9061 & n9131 ;
  assign n9133 = ~n9130 & ~n9132 ;
  assign n9134 = ~n9115 & n9133 ;
  assign n9135 = n9048 & n9134 ;
  assign n9136 = n8543 & n9124 ;
  assign n9137 = ~n9135 & n9136 ;
  assign n9138 = n9128 & ~n9137 ;
  assign n9139 = ~n9080 & ~n9138 ;
  assign n9140 = ~n9123 & n9139 ;
  assign n9141 = n8808 & ~n9138 ;
  assign n9142 = ~n9140 & ~n9141 ;
  assign n9143 = ~n8805 & ~n9041 ;
  assign n9144 = ~n9030 & n9143 ;
  assign n9145 = \pi0075  & n8804 ;
  assign n9146 = ~n9045 & ~n9145 ;
  assign n9147 = ~n9144 & n9146 ;
  assign n9148 = n9142 & ~n9147 ;
  assign n9149 = ~n9091 & n9148 ;
  assign n9150 = n8611 & n9149 ;
  assign n9151 = ~\pi0394  & ~\pi0399  ;
  assign n9152 = \pi0394  & \pi0399  ;
  assign n9153 = ~n9151 & ~n9152 ;
  assign n9154 = \pi0328  & ~\pi0398  ;
  assign n9155 = ~\pi0328  & \pi0398  ;
  assign n9156 = ~n9154 & ~n9155 ;
  assign n9157 = ~\pi0395  & n9156 ;
  assign n9158 = \pi0395  & ~n9156 ;
  assign n9159 = ~n9157 & ~n9158 ;
  assign n9160 = ~n9153 & ~n9159 ;
  assign n9161 = n9153 & n9159 ;
  assign n9162 = ~n9160 & ~n9161 ;
  assign n9163 = \pi0396  & ~\pi0408  ;
  assign n9164 = ~\pi0396  & \pi0408  ;
  assign n9165 = ~n9163 & ~n9164 ;
  assign n9166 = ~\pi0329  & ~\pi0400  ;
  assign n9167 = \pi0329  & \pi0400  ;
  assign n9168 = ~n9166 & ~n9167 ;
  assign n9169 = ~n9165 & ~n9168 ;
  assign n9170 = n9165 & n9168 ;
  assign n9171 = ~n9169 & ~n9170 ;
  assign n9172 = \pi1198  & ~n9171 ;
  assign n9173 = ~n9162 & n9172 ;
  assign n9174 = \pi1198  & n9171 ;
  assign n9175 = n9162 & n9174 ;
  assign n9176 = ~n9173 & ~n9175 ;
  assign n9177 = ~\pi0391  & ~\pi0392  ;
  assign n9178 = \pi0391  & \pi0392  ;
  assign n9179 = ~n9177 & ~n9178 ;
  assign n9180 = \pi0334  & ~\pi0413  ;
  assign n9181 = ~n9179 & n9180 ;
  assign n9182 = \pi0334  & \pi0413  ;
  assign n9183 = n9179 & n9182 ;
  assign n9184 = ~n9181 & ~n9183 ;
  assign n9185 = ~\pi0334  & \pi0413  ;
  assign n9186 = ~n9179 & n9185 ;
  assign n9187 = ~\pi0334  & ~\pi0413  ;
  assign n9188 = n9179 & n9187 ;
  assign n9189 = ~n9186 & ~n9188 ;
  assign n9190 = n9184 & n9189 ;
  assign n9191 = \pi0335  & ~\pi0393  ;
  assign n9192 = ~\pi0335  & \pi0393  ;
  assign n9193 = ~n9191 & ~n9192 ;
  assign n9194 = ~\pi0333  & \pi1197  ;
  assign n9195 = \pi0407  & ~\pi0463  ;
  assign n9196 = ~\pi0407  & \pi0463  ;
  assign n9197 = ~n9195 & ~n9196 ;
  assign n9198 = n9194 & ~n9197 ;
  assign n9199 = ~n9193 & n9198 ;
  assign n9200 = ~n9190 & n9199 ;
  assign n9201 = n9193 & n9198 ;
  assign n9202 = n9190 & n9201 ;
  assign n9203 = ~n9200 & ~n9202 ;
  assign n9204 = \pi0333  & \pi1197  ;
  assign n9205 = ~n9197 & n9204 ;
  assign n9206 = n9193 & n9205 ;
  assign n9207 = ~n9190 & n9206 ;
  assign n9208 = ~n9193 & n9205 ;
  assign n9209 = n9190 & n9208 ;
  assign n9210 = ~n9207 & ~n9209 ;
  assign n9211 = n9203 & n9210 ;
  assign n9212 = n9197 & n9204 ;
  assign n9213 = ~n9193 & n9212 ;
  assign n9214 = ~n9190 & n9213 ;
  assign n9215 = n9193 & n9212 ;
  assign n9216 = n9190 & n9215 ;
  assign n9217 = ~n9214 & ~n9216 ;
  assign n9218 = n9194 & n9197 ;
  assign n9219 = n9193 & n9218 ;
  assign n9220 = ~n9190 & n9219 ;
  assign n9221 = ~n9193 & n9218 ;
  assign n9222 = n9190 & n9221 ;
  assign n9223 = ~n9220 & ~n9222 ;
  assign n9224 = n9217 & n9223 ;
  assign n9225 = n9211 & n9224 ;
  assign n9226 = n9176 & n9225 ;
  assign n9227 = \pi0087  & ~n8606 ;
  assign n9228 = n8602 & ~n9227 ;
  assign n9229 = ~\pi0567  & n8496 ;
  assign n9230 = n9228 & n9229 ;
  assign n9231 = ~n8600 & n9230 ;
  assign n9232 = n9226 & ~n9231 ;
  assign n9233 = ~n9150 & n9232 ;
  assign n9234 = \pi0591  & n9176 ;
  assign n9235 = n9225 & n9234 ;
  assign n9236 = \pi0592  & ~n8611 ;
  assign n9237 = \pi0567  & \pi0592  ;
  assign n9238 = ~n9145 & n9237 ;
  assign n9239 = ~n9144 & n9238 ;
  assign n9240 = ~n9236 & ~n9239 ;
  assign n9241 = \pi0591  & \pi0592  ;
  assign n9242 = \pi0591  & n8611 ;
  assign n9243 = ~n8826 & n9242 ;
  assign n9244 = ~n9241 & ~n9243 ;
  assign n9245 = n9240 & ~n9244 ;
  assign n9246 = ~n9235 & ~n9245 ;
  assign n9247 = ~n9233 & ~n9246 ;
  assign n9248 = ~\pi0285  & ~\pi0286  ;
  assign n9249 = ~\pi0288  & ~\pi0289  ;
  assign n9250 = n9248 & n9249 ;
  assign n9251 = \pi0376  & ~\pi0378  ;
  assign n9252 = ~\pi0376  & \pi0378  ;
  assign n9253 = ~n9251 & ~n9252 ;
  assign n9254 = \pi0381  & ~n9253 ;
  assign n9255 = ~\pi0381  & n9253 ;
  assign n9256 = ~n9254 & ~n9255 ;
  assign n9257 = \pi0317  & ~\pi0385  ;
  assign n9258 = ~\pi0317  & \pi0385  ;
  assign n9259 = ~n9257 & ~n9258 ;
  assign n9260 = ~\pi0377  & ~\pi0439  ;
  assign n9261 = \pi0377  & \pi0439  ;
  assign n9262 = ~n9260 & ~n9261 ;
  assign n9263 = ~\pi0379  & ~\pi0382  ;
  assign n9264 = \pi0379  & \pi0382  ;
  assign n9265 = ~n9263 & ~n9264 ;
  assign n9266 = ~n9262 & ~n9265 ;
  assign n9267 = n9262 & n9265 ;
  assign n9268 = ~n9266 & ~n9267 ;
  assign n9269 = n9259 & ~n9268 ;
  assign n9270 = ~n9259 & n9268 ;
  assign n9271 = ~n9269 & ~n9270 ;
  assign n9272 = n9256 & n9271 ;
  assign n9273 = ~\pi0381  & \pi1199  ;
  assign n9274 = ~n9253 & n9273 ;
  assign n9275 = \pi0381  & \pi1199  ;
  assign n9276 = n9253 & n9275 ;
  assign n9277 = ~n9274 & ~n9276 ;
  assign n9278 = \pi1199  & ~n9259 ;
  assign n9279 = ~n9268 & n9278 ;
  assign n9280 = \pi1199  & n9259 ;
  assign n9281 = n9268 & n9280 ;
  assign n9282 = ~n9279 & ~n9281 ;
  assign n9283 = n9277 & n9282 ;
  assign n9284 = ~n9272 & ~n9283 ;
  assign n9285 = ~\pi0369  & ~\pi0375  ;
  assign n9286 = \pi0369  & \pi0375  ;
  assign n9287 = ~n9285 & ~n9286 ;
  assign n9288 = \pi0374  & n9287 ;
  assign n9289 = ~\pi0374  & ~n9287 ;
  assign n9290 = ~n9288 & ~n9289 ;
  assign n9291 = \pi0370  & ~\pi0371  ;
  assign n9292 = ~\pi0370  & \pi0371  ;
  assign n9293 = ~n9291 & ~n9292 ;
  assign n9294 = n9290 & n9293 ;
  assign n9295 = ~n9290 & ~n9293 ;
  assign n9296 = ~n9294 & ~n9295 ;
  assign n9297 = \pi0373  & ~\pi0440  ;
  assign n9298 = ~\pi0373  & \pi0440  ;
  assign n9299 = ~n9297 & ~n9298 ;
  assign n9300 = \pi0384  & ~\pi0442  ;
  assign n9301 = ~\pi0384  & \pi0442  ;
  assign n9302 = ~n9300 & ~n9301 ;
  assign n9303 = n9299 & n9302 ;
  assign n9304 = ~n9299 & ~n9302 ;
  assign n9305 = ~n9303 & ~n9304 ;
  assign n9306 = ~n9296 & n9305 ;
  assign n9307 = \pi1198  & n9293 ;
  assign n9308 = n9290 & n9307 ;
  assign n9309 = \pi1198  & n9305 ;
  assign n9310 = \pi1198  & ~n9293 ;
  assign n9311 = ~n9290 & n9310 ;
  assign n9312 = ~n9309 & ~n9311 ;
  assign n9313 = ~n9308 & n9312 ;
  assign n9314 = ~n9306 & ~n9313 ;
  assign n9315 = ~n9284 & ~n9314 ;
  assign n9316 = \pi0336  & ~\pi0383  ;
  assign n9317 = ~\pi0336  & \pi0383  ;
  assign n9318 = ~n9316 & ~n9317 ;
  assign n9319 = \pi0367  & ~n9318 ;
  assign n9320 = ~\pi0367  & n9318 ;
  assign n9321 = ~n9319 & ~n9320 ;
  assign n9322 = \pi0368  & ~\pi0389  ;
  assign n9323 = ~\pi0368  & \pi0389  ;
  assign n9324 = ~n9322 & ~n9323 ;
  assign n9325 = ~\pi0365  & ~\pi0447  ;
  assign n9326 = \pi0365  & \pi0447  ;
  assign n9327 = ~n9325 & ~n9326 ;
  assign n9328 = ~\pi0364  & ~\pi0366  ;
  assign n9329 = \pi0364  & \pi0366  ;
  assign n9330 = ~n9328 & ~n9329 ;
  assign n9331 = ~n9327 & ~n9330 ;
  assign n9332 = n9327 & n9330 ;
  assign n9333 = ~n9331 & ~n9332 ;
  assign n9334 = n9324 & ~n9333 ;
  assign n9335 = ~n9324 & n9333 ;
  assign n9336 = ~n9334 & ~n9335 ;
  assign n9337 = n9321 & n9336 ;
  assign n9338 = ~\pi0367  & \pi1197  ;
  assign n9339 = ~n9318 & n9338 ;
  assign n9340 = \pi0367  & \pi1197  ;
  assign n9341 = n9318 & n9340 ;
  assign n9342 = ~n9339 & ~n9341 ;
  assign n9343 = \pi1197  & ~n9324 ;
  assign n9344 = ~n9333 & n9343 ;
  assign n9345 = \pi1197  & n9324 ;
  assign n9346 = n9333 & n9345 ;
  assign n9347 = ~n9344 & ~n9346 ;
  assign n9348 = n9342 & n9347 ;
  assign n9349 = ~n9337 & ~n9348 ;
  assign n9350 = \pi0338  & ~\pi0388  ;
  assign n9351 = ~\pi0338  & \pi0388  ;
  assign n9352 = ~n9350 & ~n9351 ;
  assign n9353 = \pi0337  & ~n9352 ;
  assign n9354 = ~\pi0337  & n9352 ;
  assign n9355 = ~n9353 & ~n9354 ;
  assign n9356 = \pi0380  & ~\pi0387  ;
  assign n9357 = ~\pi0380  & \pi0387  ;
  assign n9358 = ~n9356 & ~n9357 ;
  assign n9359 = ~\pi0363  & ~\pi0372  ;
  assign n9360 = \pi0363  & \pi0372  ;
  assign n9361 = ~n9359 & ~n9360 ;
  assign n9362 = ~\pi0339  & ~\pi0386  ;
  assign n9363 = \pi0339  & \pi0386  ;
  assign n9364 = ~n9362 & ~n9363 ;
  assign n9365 = ~n9361 & ~n9364 ;
  assign n9366 = n9361 & n9364 ;
  assign n9367 = ~n9365 & ~n9366 ;
  assign n9368 = n9358 & ~n9367 ;
  assign n9369 = ~n9358 & n9367 ;
  assign n9370 = ~n9368 & ~n9369 ;
  assign n9371 = n9355 & n9370 ;
  assign n9372 = ~\pi0337  & \pi1196  ;
  assign n9373 = ~n9352 & n9372 ;
  assign n9374 = \pi0337  & \pi1196  ;
  assign n9375 = n9352 & n9374 ;
  assign n9376 = ~n9373 & ~n9375 ;
  assign n9377 = \pi1196  & ~n9358 ;
  assign n9378 = ~n9367 & n9377 ;
  assign n9379 = \pi1196  & n9358 ;
  assign n9380 = n9367 & n9379 ;
  assign n9381 = ~n9378 & ~n9380 ;
  assign n9382 = n9376 & n9381 ;
  assign n9383 = ~n9371 & ~n9382 ;
  assign n9384 = ~n9349 & ~n9383 ;
  assign n9385 = n9315 & n9384 ;
  assign n9386 = \pi0592  & ~n9385 ;
  assign n9387 = ~n8611 & ~n9386 ;
  assign n9388 = \pi0567  & ~n9386 ;
  assign n9389 = ~n9145 & n9388 ;
  assign n9390 = ~n9144 & n9389 ;
  assign n9391 = ~\pi0591  & ~n9386 ;
  assign n9392 = ~\pi0591  & n8611 ;
  assign n9393 = ~n8826 & n9392 ;
  assign n9394 = ~n9391 & ~n9393 ;
  assign n9395 = ~n9390 & ~n9394 ;
  assign n9396 = ~n9387 & n9395 ;
  assign n9397 = ~\pi0590  & ~n9396 ;
  assign n9398 = n9250 & n9397 ;
  assign n9399 = ~n9247 & n9398 ;
  assign n9400 = ~n8828 & n9240 ;
  assign n9401 = ~\pi0357  & ~\pi0461  ;
  assign n9402 = \pi0357  & \pi0461  ;
  assign n9403 = ~n9401 & ~n9402 ;
  assign n9404 = ~n8968 & ~n9403 ;
  assign n9405 = n8965 & n9404 ;
  assign n9406 = n8968 & ~n9403 ;
  assign n9407 = ~n8965 & n9406 ;
  assign n9408 = ~n9405 & ~n9407 ;
  assign n9409 = ~n8968 & n9403 ;
  assign n9410 = ~n8965 & n9409 ;
  assign n9411 = n8968 & n9403 ;
  assign n9412 = n8965 & n9411 ;
  assign n9413 = ~n9410 & ~n9412 ;
  assign n9414 = n9408 & n9413 ;
  assign n9415 = n8830 & ~n9414 ;
  assign n9416 = ~n9400 & n9415 ;
  assign n9417 = ~n8910 & n9240 ;
  assign n9418 = ~n8611 & n8938 ;
  assign n9419 = \pi0567  & n8938 ;
  assign n9420 = ~n9145 & n9419 ;
  assign n9421 = ~n9144 & n9420 ;
  assign n9422 = ~n9418 & ~n9421 ;
  assign n9423 = ~n8942 & n9422 ;
  assign n9424 = ~n9417 & ~n9423 ;
  assign n9425 = ~n8830 & n9403 ;
  assign n9426 = ~n8968 & n9425 ;
  assign n9427 = ~n8965 & n9426 ;
  assign n9428 = ~n8830 & ~n9403 ;
  assign n9429 = n8968 & n9428 ;
  assign n9430 = ~n8965 & n9429 ;
  assign n9431 = ~n9427 & ~n9430 ;
  assign n9432 = ~n8968 & n9428 ;
  assign n9433 = n8965 & n9432 ;
  assign n9434 = n8968 & n9425 ;
  assign n9435 = n8965 & n9434 ;
  assign n9436 = ~n9433 & ~n9435 ;
  assign n9437 = n9431 & n9436 ;
  assign n9438 = n9424 & ~n9437 ;
  assign n9439 = ~n9416 & ~n9438 ;
  assign n9440 = ~n8952 & n9414 ;
  assign n9441 = n9424 & n9440 ;
  assign n9442 = n8952 & n9414 ;
  assign n9443 = ~n9400 & n9442 ;
  assign n9444 = ~\pi0591  & ~n9443 ;
  assign n9445 = ~n9441 & n9444 ;
  assign n9446 = n9439 & n9445 ;
  assign n9447 = \pi0567  & ~n9145 ;
  assign n9448 = ~n9144 & n9447 ;
  assign n9449 = \pi0591  & n8496 ;
  assign n9450 = n8609 & n9449 ;
  assign n9451 = ~n8600 & n9450 ;
  assign n9452 = ~n9448 & n9451 ;
  assign n9453 = \pi0590  & n9250 ;
  assign n9454 = ~n9452 & n9453 ;
  assign n9455 = ~n9446 & n9454 ;
  assign n9456 = ~n9399 & ~n9455 ;
  assign n9457 = \pi0591  & n8612 ;
  assign n9458 = \pi0591  & n8778 ;
  assign n9459 = ~n8777 & n9458 ;
  assign n9460 = ~n9457 & ~n9459 ;
  assign n9461 = \pi0590  & n9460 ;
  assign n9462 = n9456 & n9461 ;
  assign n9463 = ~n9008 & n9462 ;
  assign n9464 = \pi0038  & ~\pi0100  ;
  assign n9465 = n8773 & ~n9070 ;
  assign n9466 = n9061 & n9465 ;
  assign n9467 = n8773 & n9070 ;
  assign n9468 = ~n9061 & n9467 ;
  assign n9469 = ~n9466 & ~n9468 ;
  assign n9470 = n9464 & n9469 ;
  assign n9471 = ~\pi0100  & n9469 ;
  assign n9472 = \pi0039  & ~n8793 ;
  assign n9473 = n8790 & n9472 ;
  assign n9474 = \pi0039  & n8622 ;
  assign n9475 = ~n9070 & n9474 ;
  assign n9476 = n9061 & n9475 ;
  assign n9477 = n9070 & n9474 ;
  assign n9478 = ~n9061 & n9477 ;
  assign n9479 = ~n9476 & ~n9478 ;
  assign n9480 = ~n9473 & n9479 ;
  assign n9481 = n9471 & n9480 ;
  assign n9482 = ~n9470 & ~n9481 ;
  assign n9483 = ~\pi1091  & ~n9070 ;
  assign n9484 = ~n9061 & n9483 ;
  assign n9485 = ~\pi1091  & n9070 ;
  assign n9486 = n9061 & n9485 ;
  assign n9487 = ~n9484 & ~n9486 ;
  assign n9488 = ~n8597 & ~n9487 ;
  assign n9489 = ~n8591 & n9488 ;
  assign n9490 = ~\pi0039  & ~n9489 ;
  assign n9491 = ~n8725 & n9490 ;
  assign n9492 = ~n8767 & ~n9470 ;
  assign n9493 = n9491 & n9492 ;
  assign n9494 = ~n9482 & ~n9493 ;
  assign n9495 = ~n2328 & n8622 ;
  assign n9496 = ~n9070 & n9495 ;
  assign n9497 = n9061 & n9496 ;
  assign n9498 = n9070 & n9495 ;
  assign n9499 = ~n9061 & n9498 ;
  assign n9500 = ~n9497 & ~n9499 ;
  assign n9501 = \pi0087  & n9500 ;
  assign n9502 = ~\pi1091  & ~n8606 ;
  assign n9503 = ~n8620 & n9502 ;
  assign n9504 = \pi1091  & ~n8630 ;
  assign n9505 = n2328 & ~n9504 ;
  assign n9506 = n9083 & n9502 ;
  assign n9507 = n9505 & ~n9506 ;
  assign n9508 = ~n9503 & n9507 ;
  assign n9509 = n9501 & ~n9508 ;
  assign n9510 = \pi0100  & ~n8669 ;
  assign n9511 = n8622 & ~n9070 ;
  assign n9512 = n9061 & n9511 ;
  assign n9513 = n8622 & n9070 ;
  assign n9514 = ~n9061 & n9513 ;
  assign n9515 = ~n9512 & ~n9514 ;
  assign n9516 = n9510 & n9515 ;
  assign n9517 = ~n9509 & ~n9516 ;
  assign n9518 = ~n9494 & n9517 ;
  assign n9519 = \pi0087  & ~n9509 ;
  assign n9520 = ~\pi0075  & \pi0567  ;
  assign n9521 = ~n9519 & n9520 ;
  assign n9522 = ~n9518 & n9521 ;
  assign n9523 = n7207 & n8651 ;
  assign n9524 = \pi1091  & n8797 ;
  assign n9525 = n9523 & n9524 ;
  assign n9526 = ~\pi1091  & n8797 ;
  assign n9527 = n8643 & ~n9070 ;
  assign n9528 = n9061 & n9527 ;
  assign n9529 = n8643 & n9070 ;
  assign n9530 = ~n9061 & n9529 ;
  assign n9531 = ~n9528 & ~n9530 ;
  assign n9532 = n9526 & ~n9531 ;
  assign n9533 = ~n9525 & ~n9532 ;
  assign n9534 = ~n8797 & ~n9515 ;
  assign n9535 = \pi0075  & \pi0567  ;
  assign n9536 = ~n9534 & n9535 ;
  assign n9537 = n9533 & n9536 ;
  assign n9538 = n8611 & ~n9537 ;
  assign n9539 = ~n9522 & n9538 ;
  assign n9540 = ~\pi0592  & \pi1196  ;
  assign n9541 = n8549 & ~n9070 ;
  assign n9542 = n9061 & n9541 ;
  assign n9543 = n8549 & n9070 ;
  assign n9544 = ~n9061 & n9543 ;
  assign n9545 = ~n9542 & ~n9544 ;
  assign n9546 = n9540 & n9545 ;
  assign n9547 = ~n9539 & n9546 ;
  assign n9548 = ~\pi1196  & n8612 ;
  assign n9549 = ~\pi1196  & n8778 ;
  assign n9550 = ~n8777 & n9549 ;
  assign n9551 = ~n9548 & ~n9550 ;
  assign n9552 = ~\pi1199  & n9551 ;
  assign n9553 = ~n9547 & n9552 ;
  assign n9554 = n8773 & ~n9112 ;
  assign n9555 = n9103 & n9554 ;
  assign n9556 = n8773 & n9112 ;
  assign n9557 = ~n9103 & n9556 ;
  assign n9558 = ~n9555 & ~n9557 ;
  assign n9559 = n9464 & n9558 ;
  assign n9560 = ~\pi0100  & n9558 ;
  assign n9561 = ~n9112 & n9474 ;
  assign n9562 = n9103 & n9561 ;
  assign n9563 = n9112 & n9474 ;
  assign n9564 = ~n9103 & n9563 ;
  assign n9565 = ~n9562 & ~n9564 ;
  assign n9566 = ~n9473 & n9565 ;
  assign n9567 = n9560 & n9566 ;
  assign n9568 = ~n9559 & ~n9567 ;
  assign n9569 = ~n8618 & ~n8721 ;
  assign n9570 = \pi1093  & ~n9115 ;
  assign n9571 = ~n9569 & n9570 ;
  assign n9572 = ~\pi1091  & ~n9571 ;
  assign n9573 = n8717 & n9572 ;
  assign n9574 = ~\pi0039  & ~n9573 ;
  assign n9575 = ~n8767 & ~n9559 ;
  assign n9576 = n9574 & n9575 ;
  assign n9577 = ~n9568 & ~n9576 ;
  assign n9578 = ~n2402 & n8622 ;
  assign n9579 = ~n9112 & n9578 ;
  assign n9580 = n9103 & n9579 ;
  assign n9581 = n9112 & n9578 ;
  assign n9582 = ~n9103 & n9581 ;
  assign n9583 = ~n9580 & ~n9582 ;
  assign n9584 = \pi0087  & n9583 ;
  assign n9585 = n9115 & n9502 ;
  assign n9586 = n9505 & ~n9585 ;
  assign n9587 = ~n9503 & n9586 ;
  assign n9588 = n9584 & ~n9587 ;
  assign n9589 = n8622 & ~n9112 ;
  assign n9590 = n9103 & n9589 ;
  assign n9591 = n8622 & n9112 ;
  assign n9592 = ~n9103 & n9591 ;
  assign n9593 = ~n9590 & ~n9592 ;
  assign n9594 = n9510 & n9593 ;
  assign n9595 = ~n9588 & ~n9594 ;
  assign n9596 = ~n9577 & n9595 ;
  assign n9597 = \pi0087  & ~n9588 ;
  assign n9598 = n8549 & ~n9112 ;
  assign n9599 = n9103 & n9598 ;
  assign n9600 = n8549 & n9112 ;
  assign n9601 = ~n9103 & n9600 ;
  assign n9602 = ~n9599 & ~n9601 ;
  assign n9603 = ~\pi0592  & ~\pi1196  ;
  assign n9604 = n9602 & n9603 ;
  assign n9605 = ~\pi0075  & n9604 ;
  assign n9606 = ~n9597 & n9605 ;
  assign n9607 = ~n9596 & n9606 ;
  assign n9608 = ~n8797 & ~n9593 ;
  assign n9609 = \pi0075  & ~n9608 ;
  assign n9610 = n8643 & ~n9112 ;
  assign n9611 = n9103 & n9610 ;
  assign n9612 = n8643 & n9112 ;
  assign n9613 = ~n9103 & n9612 ;
  assign n9614 = ~n9611 & ~n9613 ;
  assign n9615 = n9526 & ~n9614 ;
  assign n9616 = ~n9525 & ~n9615 ;
  assign n9617 = n9609 & n9616 ;
  assign n9618 = n9604 & n9617 ;
  assign n9619 = ~n9607 & ~n9618 ;
  assign n9620 = \pi0567  & ~n9619 ;
  assign n9621 = ~n8767 & n9491 ;
  assign n9622 = ~\pi0038  & ~n9573 ;
  assign n9623 = n9621 & n9622 ;
  assign n9624 = ~n9083 & ~n9593 ;
  assign n9625 = n8790 & ~n8793 ;
  assign n9626 = ~n9624 & ~n9625 ;
  assign n9627 = ~\pi0038  & \pi0039  ;
  assign n9628 = ~n9626 & n9627 ;
  assign n9629 = n2362 & n9469 ;
  assign n9630 = n2362 & n9558 ;
  assign n9631 = ~n9629 & ~n9630 ;
  assign n9632 = ~n9628 & ~n9631 ;
  assign n9633 = ~n9623 & n9632 ;
  assign n9634 = n6706 & ~n8638 ;
  assign n9635 = ~\pi0039  & \pi0228  ;
  assign n9636 = ~\pi0038  & \pi0232  ;
  assign n9637 = \pi1091  & n9636 ;
  assign n9638 = n9635 & n9637 ;
  assign n9639 = ~n8637 & n9638 ;
  assign n9640 = ~n9634 & n9639 ;
  assign n9641 = n9624 & ~n9640 ;
  assign n9642 = \pi0100  & ~n9641 ;
  assign n9643 = ~\pi0087  & ~n8665 ;
  assign n9644 = ~\pi0087  & ~n8668 ;
  assign n9645 = ~n9624 & n9644 ;
  assign n9646 = ~n9643 & ~n9645 ;
  assign n9647 = n9642 & ~n9646 ;
  assign n9648 = \pi0075  & ~n9534 ;
  assign n9649 = ~n9609 & ~n9648 ;
  assign n9650 = \pi1091  & n8651 ;
  assign n9651 = n8797 & n9650 ;
  assign n9652 = n7207 & n9651 ;
  assign n9653 = ~\pi1091  & n2342 ;
  assign n9654 = ~n8641 & n9653 ;
  assign n9655 = n9624 & n9654 ;
  assign n9656 = ~n9652 & ~n9655 ;
  assign n9657 = ~n9649 & n9656 ;
  assign n9658 = ~n9501 & ~n9584 ;
  assign n9659 = ~n9506 & n9587 ;
  assign n9660 = ~n9658 & ~n9659 ;
  assign n9661 = ~n9657 & ~n9660 ;
  assign n9662 = ~n9647 & n9661 ;
  assign n9663 = ~n9633 & n9662 ;
  assign n9664 = \pi0075  & ~n9657 ;
  assign n9665 = n8547 & ~n9070 ;
  assign n9666 = n9061 & n9665 ;
  assign n9667 = n8547 & n9070 ;
  assign n9668 = ~n9061 & n9667 ;
  assign n9669 = ~n9666 & ~n9668 ;
  assign n9670 = ~n9602 & ~n9669 ;
  assign n9671 = \pi0567  & \pi1196  ;
  assign n9672 = ~\pi0592  & n9671 ;
  assign n9673 = ~n9670 & n9672 ;
  assign n9674 = ~n9664 & n9673 ;
  assign n9675 = ~n9663 & n9674 ;
  assign n9676 = n9540 & ~n9670 ;
  assign n9677 = \pi1199  & ~n9604 ;
  assign n9678 = ~n9676 & n9677 ;
  assign n9679 = ~\pi0074  & \pi1199  ;
  assign n9680 = n1285 & n9679 ;
  assign n9681 = n8609 & n9680 ;
  assign n9682 = ~n8600 & n9681 ;
  assign n9683 = ~n9678 & ~n9682 ;
  assign n9684 = ~n9675 & ~n9683 ;
  assign n9685 = ~n9620 & n9684 ;
  assign n9686 = n9176 & ~n9685 ;
  assign n9687 = ~n9553 & n9686 ;
  assign n9688 = ~\pi0592  & ~n9176 ;
  assign n9689 = ~n8827 & n9688 ;
  assign n9690 = ~n9194 & ~n9689 ;
  assign n9691 = n8781 & n9690 ;
  assign n9692 = ~n9687 & n9691 ;
  assign n9693 = n9193 & n9197 ;
  assign n9694 = ~n9190 & n9693 ;
  assign n9695 = ~n9193 & n9197 ;
  assign n9696 = n9190 & n9695 ;
  assign n9697 = ~n9694 & ~n9696 ;
  assign n9698 = ~n9193 & ~n9197 ;
  assign n9699 = ~n9190 & n9698 ;
  assign n9700 = n9193 & ~n9197 ;
  assign n9701 = n9190 & n9700 ;
  assign n9702 = ~n9699 & ~n9701 ;
  assign n9703 = n9697 & n9702 ;
  assign n9704 = ~n8828 & n9194 ;
  assign n9705 = n8781 & n9704 ;
  assign n9706 = ~n9703 & ~n9705 ;
  assign n9707 = ~n9692 & n9706 ;
  assign n9708 = ~n9204 & ~n9689 ;
  assign n9709 = n8781 & n9708 ;
  assign n9710 = ~n9687 & n9709 ;
  assign n9711 = ~n8828 & n9204 ;
  assign n9712 = n8781 & n9711 ;
  assign n9713 = n9703 & ~n9712 ;
  assign n9714 = ~n9710 & n9713 ;
  assign n9715 = ~n9707 & ~n9714 ;
  assign n9716 = \pi0591  & ~n9250 ;
  assign n9717 = ~n9715 & n9716 ;
  assign n9718 = n8612 & n9391 ;
  assign n9719 = n8778 & n9391 ;
  assign n9720 = ~n8777 & n9719 ;
  assign n9721 = ~n9718 & ~n9720 ;
  assign n9722 = ~\pi0591  & n9386 ;
  assign n9723 = ~n8827 & n9722 ;
  assign n9724 = ~\pi0590  & ~n9723 ;
  assign n9725 = n9721 & n9724 ;
  assign n9726 = ~n9250 & ~n9725 ;
  assign n9727 = n9456 & ~n9726 ;
  assign n9728 = ~n9717 & n9727 ;
  assign n9729 = ~\pi0217  & n9250 ;
  assign n9730 = ~\pi0057  & ~\pi0217  ;
  assign n9731 = n6848 & n9730 ;
  assign n9732 = ~n9729 & ~n9731 ;
  assign n9733 = n8923 & ~n8932 ;
  assign n9734 = ~n8923 & n8932 ;
  assign n9735 = ~n9733 & ~n9734 ;
  assign n9736 = ~n8905 & ~n9735 ;
  assign n9737 = n8548 & n8933 ;
  assign n9738 = ~n8862 & n9737 ;
  assign n9739 = n9736 & n9738 ;
  assign n9740 = n8904 & n9540 ;
  assign n9741 = \pi1196  & ~n8548 ;
  assign n9742 = ~\pi1198  & ~n9741 ;
  assign n9743 = ~n8862 & n9742 ;
  assign n9744 = ~n9740 & n9743 ;
  assign n9745 = ~\pi0592  & ~n8830 ;
  assign n9746 = ~n9744 & n9745 ;
  assign n9747 = ~n9739 & n9746 ;
  assign n9748 = ~n8548 & ~n8830 ;
  assign n9749 = \pi0592  & n8548 ;
  assign n9750 = n8830 & ~n9749 ;
  assign n9751 = ~n9414 & ~n9750 ;
  assign n9752 = ~n9748 & n9751 ;
  assign n9753 = ~n9747 & n9752 ;
  assign n9754 = ~\pi0592  & ~n8952 ;
  assign n9755 = ~n9744 & n9754 ;
  assign n9756 = ~n9739 & n9755 ;
  assign n9757 = ~n8548 & ~n8952 ;
  assign n9758 = n8952 & ~n9749 ;
  assign n9759 = n9414 & ~n9758 ;
  assign n9760 = ~n9757 & n9759 ;
  assign n9761 = ~n9756 & n9760 ;
  assign n9762 = ~n9753 & ~n9761 ;
  assign n9763 = ~\pi0588  & ~\pi0591  ;
  assign n9764 = ~\pi0588  & \pi0590  ;
  assign n9765 = n8548 & n9764 ;
  assign n9766 = ~n9763 & ~n9765 ;
  assign n9767 = \pi1199  & ~n9112 ;
  assign n9768 = ~n9103 & n9767 ;
  assign n9769 = \pi1199  & n9112 ;
  assign n9770 = n9103 & n9769 ;
  assign n9771 = ~n9768 & ~n9770 ;
  assign n9772 = n9133 & n9771 ;
  assign n9773 = n8548 & n9772 ;
  assign n9774 = ~n9171 & n9204 ;
  assign n9775 = n9162 & n9774 ;
  assign n9776 = n9171 & n9204 ;
  assign n9777 = ~n9162 & n9776 ;
  assign n9778 = ~n9775 & ~n9777 ;
  assign n9779 = n9703 & ~n9778 ;
  assign n9780 = ~n9749 & ~n9779 ;
  assign n9781 = ~n9773 & n9780 ;
  assign n9782 = ~\pi0588  & ~\pi0590  ;
  assign n9783 = n9749 & n9782 ;
  assign n9784 = n9176 & n9782 ;
  assign n9785 = n9225 & n9784 ;
  assign n9786 = ~n9783 & ~n9785 ;
  assign n9787 = ~n9781 & ~n9786 ;
  assign n9788 = n9766 & ~n9787 ;
  assign n9789 = \pi0590  & ~n9788 ;
  assign n9790 = ~n9762 & n9789 ;
  assign n9791 = ~\pi0590  & n8548 ;
  assign n9792 = ~\pi0591  & ~n9791 ;
  assign n9793 = ~\pi0591  & \pi0592  ;
  assign n9794 = ~n9385 & n9793 ;
  assign n9795 = ~n9792 & ~n9794 ;
  assign n9796 = ~n9788 & n9795 ;
  assign n9797 = ~\pi0423  & ~\pi0424  ;
  assign n9798 = \pi0423  & \pi0424  ;
  assign n9799 = ~n9797 & ~n9798 ;
  assign n9800 = \pi0459  & n9799 ;
  assign n9801 = ~\pi0459  & ~n9799 ;
  assign n9802 = ~n9800 & ~n9801 ;
  assign n9803 = \pi0419  & ~\pi0420  ;
  assign n9804 = ~\pi0419  & \pi0420  ;
  assign n9805 = ~n9803 & ~n9804 ;
  assign n9806 = \pi0432  & n9805 ;
  assign n9807 = ~\pi0432  & ~n9805 ;
  assign n9808 = ~n9806 & ~n9807 ;
  assign n9809 = n9802 & n9808 ;
  assign n9810 = ~n9802 & ~n9808 ;
  assign n9811 = ~n9809 & ~n9810 ;
  assign n9812 = \pi0421  & ~\pi0454  ;
  assign n9813 = ~\pi0421  & \pi0454  ;
  assign n9814 = ~n9812 & ~n9813 ;
  assign n9815 = ~\pi0425  & \pi1198  ;
  assign n9816 = ~n9814 & n9815 ;
  assign n9817 = n9811 & n9816 ;
  assign n9818 = \pi0425  & \pi1198  ;
  assign n9819 = ~n9814 & n9818 ;
  assign n9820 = ~n9811 & n9819 ;
  assign n9821 = ~n9817 & ~n9820 ;
  assign n9822 = n9814 & n9818 ;
  assign n9823 = n9811 & n9822 ;
  assign n9824 = n9814 & n9815 ;
  assign n9825 = ~n9811 & n9824 ;
  assign n9826 = ~n9823 & ~n9825 ;
  assign n9827 = n9821 & n9826 ;
  assign n9828 = ~\pi0417  & ~\pi0453  ;
  assign n9829 = \pi0417  & \pi0453  ;
  assign n9830 = ~n9828 & ~n9829 ;
  assign n9831 = \pi0464  & n9830 ;
  assign n9832 = ~\pi0464  & ~n9830 ;
  assign n9833 = ~n9831 & ~n9832 ;
  assign n9834 = \pi0418  & ~\pi0437  ;
  assign n9835 = ~\pi0418  & \pi0437  ;
  assign n9836 = ~n9834 & ~n9835 ;
  assign n9837 = n9833 & n9836 ;
  assign n9838 = ~n9833 & ~n9836 ;
  assign n9839 = ~n9837 & ~n9838 ;
  assign n9840 = \pi0415  & ~\pi0431  ;
  assign n9841 = ~\pi0415  & \pi0431  ;
  assign n9842 = ~n9840 & ~n9841 ;
  assign n9843 = \pi0416  & ~\pi0438  ;
  assign n9844 = ~\pi0416  & \pi0438  ;
  assign n9845 = ~n9843 & ~n9844 ;
  assign n9846 = n9842 & n9845 ;
  assign n9847 = ~n9842 & ~n9845 ;
  assign n9848 = ~n9846 & ~n9847 ;
  assign n9849 = ~n9839 & n9848 ;
  assign n9850 = \pi1197  & n9836 ;
  assign n9851 = n9833 & n9850 ;
  assign n9852 = \pi1197  & n9848 ;
  assign n9853 = \pi1197  & ~n9836 ;
  assign n9854 = ~n9833 & n9853 ;
  assign n9855 = ~n9852 & ~n9854 ;
  assign n9856 = ~n9851 & n9855 ;
  assign n9857 = ~n9849 & ~n9856 ;
  assign n9858 = ~\pi0433  & ~\pi0451  ;
  assign n9859 = \pi0433  & \pi0451  ;
  assign n9860 = ~n9858 & ~n9859 ;
  assign n9861 = \pi0448  & n9860 ;
  assign n9862 = ~\pi0448  & ~n9860 ;
  assign n9863 = ~n9861 & ~n9862 ;
  assign n9864 = \pi0445  & ~\pi0449  ;
  assign n9865 = ~\pi0445  & \pi0449  ;
  assign n9866 = ~n9864 & ~n9865 ;
  assign n9867 = n9863 & n9866 ;
  assign n9868 = ~n9863 & ~n9866 ;
  assign n9869 = ~n9867 & ~n9868 ;
  assign n9870 = \pi0427  & ~\pi0428  ;
  assign n9871 = ~\pi0427  & \pi0428  ;
  assign n9872 = ~n9870 & ~n9871 ;
  assign n9873 = \pi0426  & ~\pi0430  ;
  assign n9874 = ~\pi0426  & \pi0430  ;
  assign n9875 = ~n9873 & ~n9874 ;
  assign n9876 = n9872 & n9875 ;
  assign n9877 = ~n9872 & ~n9875 ;
  assign n9878 = ~n9876 & ~n9877 ;
  assign n9879 = ~n9869 & n9878 ;
  assign n9880 = \pi1199  & n9866 ;
  assign n9881 = n9863 & n9880 ;
  assign n9882 = \pi1199  & n9878 ;
  assign n9883 = \pi1199  & ~n9866 ;
  assign n9884 = ~n9863 & n9883 ;
  assign n9885 = ~n9882 & ~n9884 ;
  assign n9886 = ~n9881 & n9885 ;
  assign n9887 = ~n9879 & ~n9886 ;
  assign n9888 = ~n9857 & ~n9887 ;
  assign n9889 = n9827 & n9888 ;
  assign n9890 = \pi0588  & n8548 ;
  assign n9891 = \pi0436  & ~\pi0443  ;
  assign n9892 = ~\pi0436  & \pi0443  ;
  assign n9893 = ~n9891 & ~n9892 ;
  assign n9894 = ~\pi0444  & n9893 ;
  assign n9895 = \pi0444  & ~n9893 ;
  assign n9896 = ~n9894 & ~n9895 ;
  assign n9897 = ~\pi0434  & ~\pi0446  ;
  assign n9898 = \pi0434  & \pi0446  ;
  assign n9899 = ~n9897 & ~n9898 ;
  assign n9900 = ~\pi0414  & ~\pi0422  ;
  assign n9901 = \pi0414  & \pi0422  ;
  assign n9902 = ~n9900 & ~n9901 ;
  assign n9903 = ~n9899 & ~n9902 ;
  assign n9904 = n9899 & n9902 ;
  assign n9905 = ~n9903 & ~n9904 ;
  assign n9906 = \pi0429  & ~\pi0435  ;
  assign n9907 = ~\pi0429  & \pi0435  ;
  assign n9908 = ~n9906 & ~n9907 ;
  assign n9909 = ~n9905 & n9908 ;
  assign n9910 = n9905 & ~n9908 ;
  assign n9911 = ~n9909 & ~n9910 ;
  assign n9912 = n9896 & n9911 ;
  assign n9913 = \pi1196  & ~n9908 ;
  assign n9914 = ~n9905 & n9913 ;
  assign n9915 = ~\pi0444  & \pi1196  ;
  assign n9916 = ~n9893 & n9915 ;
  assign n9917 = \pi0444  & \pi1196  ;
  assign n9918 = n9893 & n9917 ;
  assign n9919 = ~n9916 & ~n9918 ;
  assign n9920 = \pi1196  & n9908 ;
  assign n9921 = n9905 & n9920 ;
  assign n9922 = n9919 & ~n9921 ;
  assign n9923 = ~n9914 & n9922 ;
  assign n9924 = ~n9912 & ~n9923 ;
  assign n9925 = n9890 & ~n9924 ;
  assign n9926 = n9889 & n9925 ;
  assign n9927 = ~\pi0590  & ~\pi0591  ;
  assign n9928 = ~\pi0592  & n9927 ;
  assign n9929 = \pi0588  & ~n9928 ;
  assign n9930 = n8548 & n9929 ;
  assign n9931 = ~\pi0217  & ~n9930 ;
  assign n9932 = ~n9926 & n9931 ;
  assign n9933 = ~n9796 & n9932 ;
  assign n9934 = ~n9790 & n9933 ;
  assign n9935 = n9732 & ~n9934 ;
  assign n9936 = ~\pi0588  & ~n9935 ;
  assign n9937 = ~n9728 & n9936 ;
  assign n9938 = ~n9463 & n9937 ;
  assign n9939 = n8612 & ~n9250 ;
  assign n9940 = n8778 & ~n9250 ;
  assign n9941 = ~n8777 & n9940 ;
  assign n9942 = ~n9939 & ~n9941 ;
  assign n9943 = ~n8611 & n9250 ;
  assign n9944 = \pi0567  & n9250 ;
  assign n9945 = ~n9145 & n9944 ;
  assign n9946 = ~n9144 & n9945 ;
  assign n9947 = ~n9943 & ~n9946 ;
  assign n9948 = ~\pi0057  & n6848 ;
  assign n9949 = ~n9928 & n9948 ;
  assign n9950 = \pi0443  & ~\pi0444  ;
  assign n9951 = ~\pi0443  & \pi0444  ;
  assign n9952 = ~n9950 & ~n9951 ;
  assign n9953 = ~\pi0436  & ~n9908 ;
  assign n9954 = n9952 & n9953 ;
  assign n9955 = n9905 & n9954 ;
  assign n9956 = \pi0436  & ~n9908 ;
  assign n9957 = n9952 & n9956 ;
  assign n9958 = ~n9905 & n9957 ;
  assign n9959 = ~n9955 & ~n9958 ;
  assign n9960 = ~\pi0436  & n9908 ;
  assign n9961 = n9952 & n9960 ;
  assign n9962 = ~n9905 & n9961 ;
  assign n9963 = \pi0436  & n9908 ;
  assign n9964 = n9952 & n9963 ;
  assign n9965 = n9905 & n9964 ;
  assign n9966 = ~n9962 & ~n9965 ;
  assign n9967 = n9959 & n9966 ;
  assign n9968 = ~n9952 & n9956 ;
  assign n9969 = n9905 & n9968 ;
  assign n9970 = ~n9952 & n9953 ;
  assign n9971 = ~n9905 & n9970 ;
  assign n9972 = ~n9969 & ~n9971 ;
  assign n9973 = ~n9952 & n9960 ;
  assign n9974 = n9905 & n9973 ;
  assign n9975 = ~n9952 & n9963 ;
  assign n9976 = ~n9905 & n9975 ;
  assign n9977 = ~n9974 & ~n9976 ;
  assign n9978 = \pi1196  & n9977 ;
  assign n9979 = n9972 & n9978 ;
  assign n9980 = n9967 & n9979 ;
  assign n9981 = n9948 & ~n9980 ;
  assign n9982 = n9889 & n9981 ;
  assign n9983 = ~n9949 & ~n9982 ;
  assign n9984 = n9947 & ~n9983 ;
  assign n9985 = n9942 & n9984 ;
  assign n9986 = ~\pi0588  & n9948 ;
  assign n9987 = n9889 & ~n9980 ;
  assign n9988 = n9928 & ~n9987 ;
  assign n9989 = n8610 & n9988 ;
  assign n9990 = ~n8600 & n9989 ;
  assign n9991 = n9948 & n9990 ;
  assign n9992 = ~n8826 & n9991 ;
  assign n9993 = ~n9986 & ~n9992 ;
  assign n9994 = ~n9935 & n9993 ;
  assign n9995 = ~n9985 & n9994 ;
  assign n9996 = ~\pi1161  & ~\pi1162  ;
  assign n9997 = ~\pi0217  & ~\pi1163  ;
  assign n9998 = ~n9250 & ~n9948 ;
  assign n9999 = ~\pi1163  & n8548 ;
  assign n10000 = n9998 & n9999 ;
  assign n10001 = ~n9997 & ~n10000 ;
  assign n10002 = n9996 & ~n10001 ;
  assign n10003 = ~\pi1163  & n9996 ;
  assign n10004 = n9948 & n10003 ;
  assign n10005 = n9947 & n10004 ;
  assign n10006 = n9942 & n10005 ;
  assign n10007 = ~n10002 & ~n10006 ;
  assign n10008 = ~n9995 & ~n10007 ;
  assign n10009 = ~n9938 & n10008 ;
  assign n10010 = \pi1161  & ~\pi1163  ;
  assign n10011 = n1689 & n10010 ;
  assign n10012 = ~\pi0031  & \pi1162  ;
  assign n10013 = n10011 & n10012 ;
  assign n10014 = ~n10009 & ~n10013 ;
  assign n10015 = n1292 & n2404 ;
  assign n10016 = n1285 & n2467 ;
  assign n10017 = n10015 & n10016 ;
  assign n10018 = ~\pi0024  & ~\pi0841  ;
  assign n10019 = ~n6684 & ~n10018 ;
  assign n10020 = n1627 & n10019 ;
  assign n10021 = n1319 & n10020 ;
  assign n10022 = n1952 & n10021 ;
  assign n10023 = n1354 & n1652 ;
  assign n10024 = \pi0032  & n6684 ;
  assign n10025 = n10023 & n10024 ;
  assign n10026 = n1358 & n10025 ;
  assign n10027 = ~n10022 & ~n10026 ;
  assign n10028 = \pi0076  & ~\pi0084  ;
  assign n10029 = n1231 & n10028 ;
  assign n10030 = ~\pi0049  & ~\pi0066  ;
  assign n10031 = ~\pi0068  & ~\pi0073  ;
  assign n10032 = n10030 & n10031 ;
  assign n10033 = n10029 & n10032 ;
  assign n10034 = ~\pi0089  & ~\pi0102  ;
  assign n10035 = n1252 & n10034 ;
  assign n10036 = n1531 & n10035 ;
  assign n10037 = n10033 & n10036 ;
  assign n10038 = n1257 & n1423 ;
  assign n10039 = ~\pi0045  & ~\pi0048  ;
  assign n10040 = ~\pi0061  & ~\pi0104  ;
  assign n10041 = n10039 & n10040 ;
  assign n10042 = n10038 & n10041 ;
  assign n10043 = n1253 & n1424 ;
  assign n10044 = ~\pi0103  & n1238 ;
  assign n10045 = n10043 & n10044 ;
  assign n10046 = n10042 & n10045 ;
  assign n10047 = n10037 & n10046 ;
  assign n10048 = ~\pi0137  & ~n6684 ;
  assign n10049 = \pi1092  & ~\pi1093  ;
  assign n10050 = n1687 & n10049 ;
  assign n10051 = ~n9250 & ~n10050 ;
  assign n10052 = ~n1696 & n10051 ;
  assign n10053 = n10048 & ~n10052 ;
  assign n10054 = n10047 & n10053 ;
  assign n10055 = n1618 & n1635 ;
  assign n10056 = n1270 & n1320 ;
  assign n10057 = n8567 & n10056 ;
  assign n10058 = n1315 & n10057 ;
  assign n10059 = n10055 & n10058 ;
  assign n10060 = n10054 & n10059 ;
  assign n10061 = \pi0050  & n1543 ;
  assign n10062 = n1542 & n10061 ;
  assign n10063 = ~\pi0024  & n10055 ;
  assign n10064 = n10058 & n10063 ;
  assign n10065 = n10062 & n10064 ;
  assign n10066 = ~n10060 & ~n10065 ;
  assign n10067 = n10027 & n10066 ;
  assign n10068 = n1286 & n6629 ;
  assign n10069 = ~n10067 & n10068 ;
  assign n10070 = ~n6795 & n6808 ;
  assign n10071 = ~n6814 & ~n6815 ;
  assign n10072 = n1281 & n10071 ;
  assign n10073 = n1260 & n10072 ;
  assign n10074 = n10070 & n10073 ;
  assign n10075 = \pi0129  & n1281 ;
  assign n10076 = n1260 & n10075 ;
  assign n10077 = \pi0252  & n6808 ;
  assign n10078 = \pi0252  & n8640 ;
  assign n10079 = n8639 & n10078 ;
  assign n10080 = ~n10077 & ~n10079 ;
  assign n10081 = n6795 & ~n10080 ;
  assign n10082 = n10076 & n10081 ;
  assign n10083 = ~n10074 & ~n10082 ;
  assign n10084 = ~\pi0038  & ~\pi0137  ;
  assign n10085 = n1286 & n10084 ;
  assign n10086 = n2851 & n10085 ;
  assign n10087 = ~n10083 & n10086 ;
  assign n10088 = ~\pi0024  & ~n10050 ;
  assign n10089 = ~n1696 & n10088 ;
  assign n10090 = n1281 & n10089 ;
  assign n10091 = n1260 & n10090 ;
  assign n10092 = ~n6795 & ~n6808 ;
  assign n10093 = ~\pi0087  & n1288 ;
  assign n10094 = \pi0075  & ~\pi0100  ;
  assign n10095 = ~\pi0137  & n10094 ;
  assign n10096 = n10093 & n10095 ;
  assign n10097 = ~n10092 & n10096 ;
  assign n10098 = n10080 & n10097 ;
  assign n10099 = n10091 & n10098 ;
  assign n10100 = ~n10087 & ~n10099 ;
  assign n10101 = ~n10069 & n10100 ;
  assign n10102 = n10017 & ~n10101 ;
  assign n10103 = ~\pi0186  & ~\pi0299  ;
  assign n10104 = ~\pi0164  & \pi0299  ;
  assign n10105 = ~n10103 & ~n10104 ;
  assign n10106 = n8640 & n10105 ;
  assign n10107 = n8601 & n10106 ;
  assign n10108 = \pi0054  & n10107 ;
  assign n10109 = \pi0178  & \pi0183  ;
  assign n10110 = ~\pi0178  & ~\pi0183  ;
  assign n10111 = n6706 & ~n10110 ;
  assign n10112 = ~n10109 & n10111 ;
  assign n10113 = ~\pi0299  & ~n10112 ;
  assign n10114 = ~\pi0149  & ~\pi0157  ;
  assign n10115 = \pi0149  & \pi0157  ;
  assign n10116 = ~n10114 & ~n10115 ;
  assign n10117 = n8640 & n10116 ;
  assign n10118 = \pi0232  & ~\pi0299  ;
  assign n10119 = ~n10117 & ~n10118 ;
  assign n10120 = ~n10113 & ~n10119 ;
  assign n10121 = \pi0054  & ~n8601 ;
  assign n10122 = ~n10120 & n10121 ;
  assign n10123 = ~n10108 & ~n10122 ;
  assign n10124 = ~\pi0074  & ~n10123 ;
  assign n10125 = n1292 & n2467 ;
  assign n10126 = \pi0164  & \pi0232  ;
  assign n10127 = n6706 & n10126 ;
  assign n10128 = ~\pi0074  & n8601 ;
  assign n10129 = n10127 & n10128 ;
  assign n10130 = ~\pi0074  & ~n8601 ;
  assign n10131 = ~n10117 & n10130 ;
  assign n10132 = ~n10129 & ~n10131 ;
  assign n10133 = ~n8601 & ~n10117 ;
  assign n10134 = ~\pi0038  & ~\pi0054  ;
  assign n10135 = ~n10133 & n10134 ;
  assign n10136 = ~n10132 & ~n10135 ;
  assign n10137 = \pi0169  & \pi0232  ;
  assign n10138 = n6706 & n10137 ;
  assign n10139 = \pi0074  & n8601 ;
  assign n10140 = n10138 & n10139 ;
  assign n10141 = \pi0074  & ~n8601 ;
  assign n10142 = ~n10117 & n10141 ;
  assign n10143 = ~n10140 & ~n10142 ;
  assign n10144 = n2467 & n10143 ;
  assign n10145 = ~n10136 & n10144 ;
  assign n10146 = ~n10125 & ~n10145 ;
  assign n10147 = n8601 & n8640 ;
  assign n10148 = \pi0191  & ~\pi0299  ;
  assign n10149 = \pi0169  & \pi0299  ;
  assign n10150 = ~n10148 & ~n10149 ;
  assign n10151 = n10147 & ~n10150 ;
  assign n10152 = \pi0074  & n10151 ;
  assign n10153 = ~n10120 & n10141 ;
  assign n10154 = ~n10152 & ~n10153 ;
  assign n10155 = ~\pi0038  & ~\pi0040  ;
  assign n10156 = n1256 & n10155 ;
  assign n10157 = n2511 & n8601 ;
  assign n10158 = n10156 & n10157 ;
  assign n10159 = ~n1292 & n10158 ;
  assign n10160 = ~\pi0055  & ~n10159 ;
  assign n10161 = n10154 & n10160 ;
  assign n10162 = ~n10146 & n10161 ;
  assign n10163 = ~n10124 & n10162 ;
  assign n10164 = ~n10146 & ~n10159 ;
  assign n10165 = \pi0055  & ~n10140 ;
  assign n10166 = ~n10142 & n10165 ;
  assign n10167 = n1292 & ~n10166 ;
  assign n10168 = ~\pi0035  & ~\pi0058  ;
  assign n10169 = n1320 & n10168 ;
  assign n10170 = n1344 & n10169 ;
  assign n10171 = n1273 & n10170 ;
  assign n10172 = n1355 & n10171 ;
  assign n10173 = n1249 & n10172 ;
  assign n10174 = ~\pi0032  & n1618 ;
  assign n10175 = ~\pi0095  & n2341 ;
  assign n10176 = n10174 & n10175 ;
  assign n10177 = \pi0149  & \pi0232  ;
  assign n10178 = n6706 & n10177 ;
  assign n10179 = ~\pi0092  & ~n10178 ;
  assign n10180 = n10176 & n10179 ;
  assign n10181 = n10173 & n10180 ;
  assign n10182 = ~\pi0040  & n1256 ;
  assign n10183 = n8601 & n10182 ;
  assign n10184 = n10134 & n10183 ;
  assign n10185 = ~n10181 & n10184 ;
  assign n10186 = \pi0164  & ~n10134 ;
  assign n10187 = n10147 & n10186 ;
  assign n10188 = ~n10133 & ~n10187 ;
  assign n10189 = ~n10185 & n10188 ;
  assign n10190 = ~\pi0074  & n1292 ;
  assign n10191 = ~n10189 & n10190 ;
  assign n10192 = ~n10167 & ~n10191 ;
  assign n10193 = n10164 & n10192 ;
  assign n10194 = ~n10163 & ~n10193 ;
  assign n10195 = n6706 & n10118 ;
  assign n10196 = ~\pi0164  & \pi0186  ;
  assign n10197 = n10195 & n10196 ;
  assign n10198 = \pi0038  & n10197 ;
  assign n10199 = ~n8375 & n10198 ;
  assign n10200 = \pi0299  & n8640 ;
  assign n10201 = ~n8375 & n10200 ;
  assign n10202 = ~\pi0186  & ~n10201 ;
  assign n10203 = \pi0186  & n6784 ;
  assign n10204 = n1266 & n10203 ;
  assign n10205 = n1354 & n10204 ;
  assign n10206 = n1358 & n10205 ;
  assign n10207 = \pi0164  & ~\pi0186  ;
  assign n10208 = ~n10127 & ~n10207 ;
  assign n10209 = ~n10206 & ~n10208 ;
  assign n10210 = \pi0038  & n10209 ;
  assign n10211 = ~n10202 & n10210 ;
  assign n10212 = ~n10199 & ~n10211 ;
  assign n10213 = ~\pi0100  & ~n10212 ;
  assign n10214 = ~\pi0176  & ~\pi0299  ;
  assign n10215 = ~n10182 & n10214 ;
  assign n10216 = n1696 & n6745 ;
  assign n10217 = n1264 & n1618 ;
  assign n10218 = n10216 & n10217 ;
  assign n10219 = n10173 & n10218 ;
  assign n10220 = ~n6955 & n10182 ;
  assign n10221 = n6769 & ~n10220 ;
  assign n10222 = n10214 & n10221 ;
  assign n10223 = n10219 & n10222 ;
  assign n10224 = ~n10215 & ~n10223 ;
  assign n10225 = ~\pi0040  & ~\pi0174  ;
  assign n10226 = n1256 & n10225 ;
  assign n10227 = ~n6955 & n10226 ;
  assign n10228 = n6922 & ~n6931 ;
  assign n10229 = n6722 & n10228 ;
  assign n10230 = ~n10216 & ~n10229 ;
  assign n10231 = n10173 & ~n10230 ;
  assign n10232 = n6714 & n10217 ;
  assign n10233 = n10231 & n10232 ;
  assign n10234 = n10226 & ~n10233 ;
  assign n10235 = ~n10227 & ~n10234 ;
  assign n10236 = n10224 & ~n10235 ;
  assign n10237 = n10182 & ~n10233 ;
  assign n10238 = ~\pi0299  & ~n10220 ;
  assign n10239 = ~n10237 & n10238 ;
  assign n10240 = ~n6761 & ~n10182 ;
  assign n10241 = n6706 & n6955 ;
  assign n10242 = ~n6761 & n10241 ;
  assign n10243 = n10217 & n10242 ;
  assign n10244 = n10229 & n10243 ;
  assign n10245 = n10173 & n10244 ;
  assign n10246 = ~n10240 & ~n10245 ;
  assign n10247 = ~\pi0299  & ~n10246 ;
  assign n10248 = n10224 & ~n10247 ;
  assign n10249 = ~n10239 & n10248 ;
  assign n10250 = ~n10236 & ~n10249 ;
  assign n10251 = \pi0232  & n10250 ;
  assign n10252 = ~n6732 & ~n10182 ;
  assign n10253 = n6743 & n10217 ;
  assign n10254 = n10231 & n10253 ;
  assign n10255 = ~n10252 & ~n10254 ;
  assign n10256 = n10237 & n10255 ;
  assign n10257 = ~n6736 & n10217 ;
  assign n10258 = n10216 & n10257 ;
  assign n10259 = n10173 & n10258 ;
  assign n10260 = ~\pi0152  & n6706 ;
  assign n10261 = n10182 & n10260 ;
  assign n10262 = ~n10259 & n10261 ;
  assign n10263 = ~\pi0154  & ~n10262 ;
  assign n10264 = ~n10256 & n10263 ;
  assign n10265 = n10217 & n10229 ;
  assign n10266 = n10173 & n10265 ;
  assign n10267 = n10182 & ~n10266 ;
  assign n10268 = \pi0152  & n6706 ;
  assign n10269 = ~n6732 & n10268 ;
  assign n10270 = ~n10267 & n10269 ;
  assign n10271 = n10237 & ~n10270 ;
  assign n10272 = \pi0154  & ~n10271 ;
  assign n10273 = ~n10264 & ~n10272 ;
  assign n10274 = n7597 & n10273 ;
  assign n10275 = ~n7597 & n10182 ;
  assign n10276 = \pi0232  & \pi0299  ;
  assign n10277 = ~n10275 & n10276 ;
  assign n10278 = ~n10274 & n10277 ;
  assign n10279 = ~n10251 & ~n10278 ;
  assign n10280 = \pi0299  & ~n10275 ;
  assign n10281 = ~n10256 & n10280 ;
  assign n10282 = n6769 & n10217 ;
  assign n10283 = n10231 & n10282 ;
  assign n10284 = ~n10240 & ~n10283 ;
  assign n10285 = n10238 & ~n10284 ;
  assign n10286 = ~n10239 & ~n10285 ;
  assign n10287 = ~n10281 & n10286 ;
  assign n10288 = ~\pi0232  & ~n10287 ;
  assign n10289 = \pi0039  & ~n10288 ;
  assign n10290 = n10279 & n10289 ;
  assign n10291 = n2327 & n10290 ;
  assign n10292 = n1256 & ~n10173 ;
  assign n10293 = ~\pi0051  & \pi0070  ;
  assign n10294 = ~n10292 & n10293 ;
  assign n10295 = \pi0051  & ~n1256 ;
  assign n10296 = ~\pi0040  & n1262 ;
  assign n10297 = ~n10295 & n10296 ;
  assign n10298 = ~n10294 & n10297 ;
  assign n10299 = n1256 & ~n1262 ;
  assign n10300 = ~\pi0040  & n10299 ;
  assign n10301 = n1264 & ~n10300 ;
  assign n10302 = ~n10298 & n10301 ;
  assign n10303 = \pi0050  & ~\pi0060  ;
  assign n10304 = n1543 & n10303 ;
  assign n10305 = n1542 & n10304 ;
  assign n10306 = ~\pi0053  & ~n1559 ;
  assign n10307 = ~\pi0111  & n1244 ;
  assign n10308 = ~\pi0036  & ~\pi0082  ;
  assign n10309 = ~\pi0084  & n10308 ;
  assign n10310 = n10307 & n10309 ;
  assign n10311 = ~\pi0068  & n1245 ;
  assign n10312 = ~\pi0066  & \pi0073  ;
  assign n10313 = n1243 & n10312 ;
  assign n10314 = n10311 & n10313 ;
  assign n10315 = n1242 & n10314 ;
  assign n10316 = n10310 & n10315 ;
  assign n10317 = n1257 & n1275 ;
  assign n10318 = n1255 & n10317 ;
  assign n10319 = n10316 & n10318 ;
  assign n10320 = n1256 & ~n10319 ;
  assign n10321 = n10306 & n10320 ;
  assign n10322 = ~n10305 & n10321 ;
  assign n10323 = n1249 & n1355 ;
  assign n10324 = \pi0053  & ~n10323 ;
  assign n10325 = n10320 & n10324 ;
  assign n10326 = n1256 & ~n1273 ;
  assign n10327 = ~\pi0058  & n1274 ;
  assign n10328 = ~n10326 & n10327 ;
  assign n10329 = ~n10325 & n10328 ;
  assign n10330 = ~n10322 & n10329 ;
  assign n10331 = ~\pi0058  & ~n1256 ;
  assign n10332 = ~n1274 & n10331 ;
  assign n10333 = ~n1273 & n10331 ;
  assign n10334 = ~n10332 & ~n10333 ;
  assign n10335 = ~\pi0090  & n7083 ;
  assign n10336 = n1256 & n7083 ;
  assign n10337 = ~n10335 & ~n10336 ;
  assign n10338 = ~\pi0058  & ~\pi0841  ;
  assign n10339 = ~n10335 & n10338 ;
  assign n10340 = n1358 & n10339 ;
  assign n10341 = ~n10337 & ~n10340 ;
  assign n10342 = n1256 & ~n1358 ;
  assign n10343 = \pi0058  & ~n10342 ;
  assign n10344 = n10341 & ~n10343 ;
  assign n10345 = n10334 & n10344 ;
  assign n10346 = ~n10330 & n10345 ;
  assign n10347 = n1358 & n10338 ;
  assign n10348 = \pi0090  & n10336 ;
  assign n10349 = ~n10347 & n10348 ;
  assign n10350 = n1256 & ~n7083 ;
  assign n10351 = n1364 & ~n10350 ;
  assign n10352 = ~n10349 & n10351 ;
  assign n10353 = n10301 & n10352 ;
  assign n10354 = ~n10346 & n10353 ;
  assign n10355 = ~n10302 & ~n10354 ;
  assign n10356 = ~\pi0040  & \pi0479  ;
  assign n10357 = n1256 & n10356 ;
  assign n10358 = \pi0095  & ~n10357 ;
  assign n10359 = n10173 & n10174 ;
  assign n10360 = ~\pi0040  & ~\pi0479  ;
  assign n10361 = n1256 & n10360 ;
  assign n10362 = ~n10359 & n10361 ;
  assign n10363 = n10358 & ~n10362 ;
  assign n10364 = n1739 & ~n10182 ;
  assign n10365 = ~n10363 & ~n10364 ;
  assign n10366 = n10355 & n10365 ;
  assign n10367 = ~\pi0232  & ~n10366 ;
  assign n10368 = \pi0032  & ~n10182 ;
  assign n10369 = n1618 & n1718 ;
  assign n10370 = \pi0032  & n10338 ;
  assign n10371 = n10369 & n10370 ;
  assign n10372 = n1358 & n10371 ;
  assign n10373 = ~n10368 & ~n10372 ;
  assign n10374 = ~\pi0095  & ~n10373 ;
  assign n10375 = n10355 & ~n10374 ;
  assign n10376 = ~\pi0232  & ~n6684 ;
  assign n10377 = ~n10375 & n10376 ;
  assign n10378 = ~n10367 & ~n10377 ;
  assign n10379 = n2328 & n10378 ;
  assign n10380 = ~n10291 & ~n10379 ;
  assign n10381 = ~n10213 & n10380 ;
  assign n10382 = ~\pi0174  & ~n10363 ;
  assign n10383 = \pi0095  & n10382 ;
  assign n10384 = \pi0095  & n6706 ;
  assign n10385 = n10182 & n10384 ;
  assign n10386 = n1262 & ~n10295 ;
  assign n10387 = ~\pi0032  & ~n10299 ;
  assign n10388 = ~n10386 & n10387 ;
  assign n10389 = ~n10305 & n10306 ;
  assign n10390 = ~\pi0053  & n1274 ;
  assign n10391 = n1274 & n1355 ;
  assign n10392 = n1249 & n10391 ;
  assign n10393 = ~n10390 & ~n10392 ;
  assign n10394 = n1273 & ~n10393 ;
  assign n10395 = ~n10389 & n10394 ;
  assign n10396 = ~\pi0058  & n1256 ;
  assign n10397 = ~n10342 & ~n10396 ;
  assign n10398 = ~n10395 & ~n10397 ;
  assign n10399 = ~n1358 & n6637 ;
  assign n10400 = ~\pi0070  & ~\pi0090  ;
  assign n10401 = ~n10350 & n10400 ;
  assign n10402 = ~n10399 & n10401 ;
  assign n10403 = ~n10398 & n10402 ;
  assign n10404 = \pi0070  & ~n10292 ;
  assign n10405 = ~\pi0070  & ~n10350 ;
  assign n10406 = ~n10341 & n10405 ;
  assign n10407 = ~n10404 & ~n10406 ;
  assign n10408 = ~n10403 & n10407 ;
  assign n10409 = ~\pi0051  & n10387 ;
  assign n10410 = ~n10408 & n10409 ;
  assign n10411 = ~n10388 & ~n10410 ;
  assign n10412 = ~\pi0032  & \pi0040  ;
  assign n10413 = n6706 & n10182 ;
  assign n10414 = n1264 & n6706 ;
  assign n10415 = ~n10413 & ~n10414 ;
  assign n10416 = ~n10412 & ~n10415 ;
  assign n10417 = n10411 & n10416 ;
  assign n10418 = ~n10385 & ~n10417 ;
  assign n10419 = n10373 & ~n10412 ;
  assign n10420 = n10411 & n10419 ;
  assign n10421 = ~\pi0095  & ~\pi0198  ;
  assign n10422 = ~n10420 & n10421 ;
  assign n10423 = ~n10418 & ~n10422 ;
  assign n10424 = ~n6706 & ~n10364 ;
  assign n10425 = ~n10363 & n10424 ;
  assign n10426 = n10355 & n10425 ;
  assign n10427 = ~\pi0198  & ~n10375 ;
  assign n10428 = n10426 & ~n10427 ;
  assign n10429 = ~\pi0183  & ~n10428 ;
  assign n10430 = ~n10423 & n10429 ;
  assign n10431 = \pi0095  & ~n10182 ;
  assign n10432 = n6706 & ~n10431 ;
  assign n10433 = n1256 & ~n10323 ;
  assign n10434 = \pi0058  & n1344 ;
  assign n10435 = n1273 & n10434 ;
  assign n10436 = n1256 & ~n10435 ;
  assign n10437 = n1320 & ~n10436 ;
  assign n10438 = ~n10433 & n10437 ;
  assign n10439 = ~n1256 & n7081 ;
  assign n10440 = n7081 & n10338 ;
  assign n10441 = n1358 & n10440 ;
  assign n10442 = ~n10439 & ~n10441 ;
  assign n10443 = ~n10438 & n10442 ;
  assign n10444 = ~n1634 & ~n10182 ;
  assign n10445 = ~\pi0035  & n1618 ;
  assign n10446 = \pi0093  & ~n1256 ;
  assign n10447 = n10445 & ~n10446 ;
  assign n10448 = ~n10444 & n10447 ;
  assign n10449 = n10443 & n10448 ;
  assign n10450 = ~\pi0032  & ~n1256 ;
  assign n10451 = ~\pi0032  & ~\pi0035  ;
  assign n10452 = n1618 & n10451 ;
  assign n10453 = ~n10450 & ~n10452 ;
  assign n10454 = ~n10444 & n10453 ;
  assign n10455 = ~\pi0095  & ~n10454 ;
  assign n10456 = ~n10449 & n10455 ;
  assign n10457 = n10432 & ~n10456 ;
  assign n10458 = ~n10426 & ~n10457 ;
  assign n10459 = ~\pi0198  & ~n10457 ;
  assign n10460 = ~n10375 & n10459 ;
  assign n10461 = ~n10458 & ~n10460 ;
  assign n10462 = \pi0183  & ~n10461 ;
  assign n10463 = n10382 & ~n10462 ;
  assign n10464 = ~n10430 & n10463 ;
  assign n10465 = ~n10383 & ~n10464 ;
  assign n10466 = \pi0090  & n1256 ;
  assign n10467 = ~n10347 & n10466 ;
  assign n10468 = n1273 & n10327 ;
  assign n10469 = n10318 & n10468 ;
  assign n10470 = n10316 & n10469 ;
  assign n10471 = ~\pi0090  & ~n10470 ;
  assign n10472 = ~\pi0093  & ~n10453 ;
  assign n10473 = ~n10471 & n10472 ;
  assign n10474 = ~n10436 & n10472 ;
  assign n10475 = ~n10433 & n10474 ;
  assign n10476 = ~n10473 & ~n10475 ;
  assign n10477 = ~n10467 & ~n10476 ;
  assign n10478 = ~n10447 & ~n10453 ;
  assign n10479 = ~n10444 & ~n10478 ;
  assign n10480 = ~n10363 & n10479 ;
  assign n10481 = ~n10477 & n10480 ;
  assign n10482 = \pi0095  & ~n10363 ;
  assign n10483 = \pi0183  & n6706 ;
  assign n10484 = ~n10482 & n10483 ;
  assign n10485 = ~n10481 & n10484 ;
  assign n10486 = \pi0174  & ~n10485 ;
  assign n10487 = ~\pi0180  & ~n10486 ;
  assign n10488 = ~\pi0180  & ~n10483 ;
  assign n10489 = ~n10366 & n10488 ;
  assign n10490 = ~\pi0198  & n10488 ;
  assign n10491 = ~n10375 & n10490 ;
  assign n10492 = ~n10489 & ~n10491 ;
  assign n10493 = ~n10487 & n10492 ;
  assign n10494 = n10465 & ~n10493 ;
  assign n10495 = n10355 & ~n10364 ;
  assign n10496 = ~\pi0040  & n6706 ;
  assign n10497 = ~n10431 & n10496 ;
  assign n10498 = \pi0198  & n10497 ;
  assign n10499 = ~n10374 & n10497 ;
  assign n10500 = n10355 & n10499 ;
  assign n10501 = ~n10498 & ~n10500 ;
  assign n10502 = n10495 & ~n10501 ;
  assign n10503 = ~n10428 & ~n10502 ;
  assign n10504 = ~\pi0183  & n10503 ;
  assign n10505 = n10432 & ~n10444 ;
  assign n10506 = ~n10478 & n10505 ;
  assign n10507 = ~n10477 & n10506 ;
  assign n10508 = \pi0183  & ~n10385 ;
  assign n10509 = ~n10507 & n10508 ;
  assign n10510 = ~n10426 & n10509 ;
  assign n10511 = ~\pi0198  & n10509 ;
  assign n10512 = ~n10375 & n10511 ;
  assign n10513 = ~n10510 & ~n10512 ;
  assign n10514 = \pi0174  & n10513 ;
  assign n10515 = ~n10504 & n10514 ;
  assign n10516 = ~\pi0174  & ~n10462 ;
  assign n10517 = ~n10430 & n10516 ;
  assign n10518 = \pi0180  & ~n10517 ;
  assign n10519 = ~n10515 & n10518 ;
  assign n10520 = ~n10494 & ~n10519 ;
  assign n10521 = ~\pi0193  & n10520 ;
  assign n10522 = ~\pi0183  & ~n10426 ;
  assign n10523 = ~\pi0183  & ~\pi0198  ;
  assign n10524 = ~n10375 & n10523 ;
  assign n10525 = ~n10522 & ~n10524 ;
  assign n10526 = ~\pi0040  & \pi0095  ;
  assign n10527 = n1256 & n10526 ;
  assign n10528 = n1320 & n1321 ;
  assign n10529 = ~\pi0070  & n10386 ;
  assign n10530 = n1256 & n10386 ;
  assign n10531 = ~n10173 & n10530 ;
  assign n10532 = ~n10529 & ~n10531 ;
  assign n10533 = n1277 & n7083 ;
  assign n10534 = ~\pi0070  & ~n1256 ;
  assign n10535 = ~n10533 & n10534 ;
  assign n10536 = ~n10532 & ~n10535 ;
  assign n10537 = ~n10528 & n10536 ;
  assign n10538 = n10334 & n10536 ;
  assign n10539 = ~n10330 & n10538 ;
  assign n10540 = ~n10537 & ~n10539 ;
  assign n10541 = \pi0051  & n1256 ;
  assign n10542 = n1262 & n10541 ;
  assign n10543 = ~\pi0040  & ~n1256 ;
  assign n10544 = n1262 & n1634 ;
  assign n10545 = ~n10543 & ~n10544 ;
  assign n10546 = ~n10542 & ~n10545 ;
  assign n10547 = n10540 & n10546 ;
  assign n10548 = \pi0032  & ~\pi0040  ;
  assign n10549 = ~n1256 & n10548 ;
  assign n10550 = ~n1263 & ~n10182 ;
  assign n10551 = ~n10431 & ~n10550 ;
  assign n10552 = ~n10549 & n10551 ;
  assign n10553 = ~n10547 & n10552 ;
  assign n10554 = ~n10527 & ~n10553 ;
  assign n10555 = \pi0095  & ~n10543 ;
  assign n10556 = \pi0032  & ~n10543 ;
  assign n10557 = ~\pi0040  & n10338 ;
  assign n10558 = n10369 & n10557 ;
  assign n10559 = n1358 & n10558 ;
  assign n10560 = n10556 & ~n10559 ;
  assign n10561 = ~\pi0040  & ~n10299 ;
  assign n10562 = ~n10542 & n10561 ;
  assign n10563 = ~n10560 & n10562 ;
  assign n10564 = n10540 & n10563 ;
  assign n10565 = \pi0032  & ~n10560 ;
  assign n10566 = ~\pi0095  & ~n10565 ;
  assign n10567 = ~n10564 & n10566 ;
  assign n10568 = ~n10555 & ~n10567 ;
  assign n10569 = ~n10554 & ~n10568 ;
  assign n10570 = ~\pi0198  & ~n6706 ;
  assign n10571 = ~\pi0040  & ~\pi0198  ;
  assign n10572 = n1256 & n10571 ;
  assign n10573 = ~n10570 & ~n10572 ;
  assign n10574 = ~n10569 & ~n10573 ;
  assign n10575 = ~n10363 & ~n10550 ;
  assign n10576 = ~n10549 & n10575 ;
  assign n10577 = ~n10547 & n10576 ;
  assign n10578 = ~n10482 & ~n10577 ;
  assign n10579 = n6706 & ~n10578 ;
  assign n10580 = ~n10574 & n10579 ;
  assign n10581 = ~n10525 & ~n10580 ;
  assign n10582 = n1314 & n10316 ;
  assign n10583 = ~\pi0095  & n10452 ;
  assign n10584 = n10058 & n10583 ;
  assign n10585 = n10582 & n10584 ;
  assign n10586 = ~\pi0095  & ~n10182 ;
  assign n10587 = n6706 & ~n10586 ;
  assign n10588 = ~n10585 & n10587 ;
  assign n10589 = \pi0183  & ~n10588 ;
  assign n10590 = \pi0183  & n10358 ;
  assign n10591 = ~n10362 & n10590 ;
  assign n10592 = ~n10589 & ~n10591 ;
  assign n10593 = ~n10426 & ~n10592 ;
  assign n10594 = ~\pi0198  & ~n10592 ;
  assign n10595 = ~n10375 & n10594 ;
  assign n10596 = ~n10593 & ~n10595 ;
  assign n10597 = ~\pi0180  & n10596 ;
  assign n10598 = ~n10581 & n10597 ;
  assign n10599 = n6706 & ~n10554 ;
  assign n10600 = ~\pi0198  & ~n10569 ;
  assign n10601 = n10599 & ~n10600 ;
  assign n10602 = ~n10525 & ~n10601 ;
  assign n10603 = n10432 & ~n10586 ;
  assign n10604 = ~n10585 & n10603 ;
  assign n10605 = ~n10426 & ~n10604 ;
  assign n10606 = ~\pi0198  & ~n10604 ;
  assign n10607 = ~n10375 & n10606 ;
  assign n10608 = ~n10605 & ~n10607 ;
  assign n10609 = \pi0183  & ~n10608 ;
  assign n10610 = \pi0180  & ~n10609 ;
  assign n10611 = ~n10602 & n10610 ;
  assign n10612 = ~n10598 & ~n10611 ;
  assign n10613 = \pi0174  & n10612 ;
  assign n10614 = \pi0183  & ~n10586 ;
  assign n10615 = ~n10363 & n10614 ;
  assign n10616 = ~n10373 & n10421 ;
  assign n10617 = ~n1256 & ~n10533 ;
  assign n10618 = ~\pi0070  & ~n10617 ;
  assign n10619 = n1256 & ~n10617 ;
  assign n10620 = ~n10173 & n10619 ;
  assign n10621 = ~n10618 & ~n10620 ;
  assign n10622 = ~n10169 & ~n10621 ;
  assign n10623 = n1256 & ~n10621 ;
  assign n10624 = ~n10395 & n10623 ;
  assign n10625 = ~n10622 & ~n10624 ;
  assign n10626 = \pi0070  & n1256 ;
  assign n10627 = ~n10173 & n10626 ;
  assign n10628 = ~\pi0051  & ~n10299 ;
  assign n10629 = ~n10627 & n10628 ;
  assign n10630 = n10625 & n10629 ;
  assign n10631 = ~n1256 & ~n1262 ;
  assign n10632 = ~n10295 & ~n10631 ;
  assign n10633 = ~\pi0040  & n10632 ;
  assign n10634 = ~n10630 & n10633 ;
  assign n10635 = ~\pi0032  & n10421 ;
  assign n10636 = ~n10634 & n10635 ;
  assign n10637 = ~n10616 & ~n10636 ;
  assign n10638 = ~n10444 & n10632 ;
  assign n10639 = ~n10630 & n10638 ;
  assign n10640 = n1256 & n10548 ;
  assign n10641 = ~\pi0095  & ~n10640 ;
  assign n10642 = ~n10639 & n10641 ;
  assign n10643 = \pi0183  & n10586 ;
  assign n10644 = ~n10591 & ~n10643 ;
  assign n10645 = ~n10363 & n10644 ;
  assign n10646 = ~n10642 & n10645 ;
  assign n10647 = n10637 & n10646 ;
  assign n10648 = ~n10615 & ~n10647 ;
  assign n10649 = ~\pi0180  & n6706 ;
  assign n10650 = ~n10648 & n10649 ;
  assign n10651 = ~\pi0180  & n10426 ;
  assign n10652 = ~n10427 & n10651 ;
  assign n10653 = ~\pi0174  & ~n10652 ;
  assign n10654 = ~n10650 & n10653 ;
  assign n10655 = \pi0193  & ~n10654 ;
  assign n10656 = \pi0193  & n10525 ;
  assign n10657 = ~\pi0040  & ~n10560 ;
  assign n10658 = ~n10565 & ~n10657 ;
  assign n10659 = ~n10565 & n10632 ;
  assign n10660 = ~n10630 & n10659 ;
  assign n10661 = ~n10658 & ~n10660 ;
  assign n10662 = n10421 & ~n10661 ;
  assign n10663 = ~n1634 & ~n10543 ;
  assign n10664 = ~n10549 & n10663 ;
  assign n10665 = ~n10549 & n10632 ;
  assign n10666 = ~n10630 & n10665 ;
  assign n10667 = ~n10664 & ~n10666 ;
  assign n10668 = ~\pi0095  & \pi0198  ;
  assign n10669 = ~n10667 & n10668 ;
  assign n10670 = ~n10555 & ~n10669 ;
  assign n10671 = ~n10662 & n10670 ;
  assign n10672 = \pi0193  & n10496 ;
  assign n10673 = ~n10671 & n10672 ;
  assign n10674 = ~n10656 & ~n10673 ;
  assign n10675 = ~n10182 & n10483 ;
  assign n10676 = \pi0183  & ~n6706 ;
  assign n10677 = ~n10366 & n10676 ;
  assign n10678 = ~\pi0198  & n10676 ;
  assign n10679 = ~n10375 & n10678 ;
  assign n10680 = ~n10677 & ~n10679 ;
  assign n10681 = ~n10675 & n10680 ;
  assign n10682 = \pi0180  & n10681 ;
  assign n10683 = ~n10674 & n10682 ;
  assign n10684 = ~n10655 & ~n10683 ;
  assign n10685 = ~n10613 & ~n10684 ;
  assign n10686 = ~n10521 & ~n10685 ;
  assign n10687 = ~\pi0299  & n10686 ;
  assign n10688 = ~\pi0210  & ~n10375 ;
  assign n10689 = \pi0152  & n10426 ;
  assign n10690 = ~n10688 & n10689 ;
  assign n10691 = ~n10364 & ~n10431 ;
  assign n10692 = n10355 & n10691 ;
  assign n10693 = n10268 & n10692 ;
  assign n10694 = ~n10688 & n10693 ;
  assign n10695 = ~n10690 & ~n10694 ;
  assign n10696 = \pi0158  & \pi0299  ;
  assign n10697 = \pi0152  & ~\pi0172  ;
  assign n10698 = n10696 & n10697 ;
  assign n10699 = ~\pi0095  & ~\pi0210  ;
  assign n10700 = ~n10420 & n10699 ;
  assign n10701 = ~n10418 & ~n10700 ;
  assign n10702 = ~\pi0172  & ~n10426 ;
  assign n10703 = ~\pi0172  & ~\pi0210  ;
  assign n10704 = ~n10375 & n10703 ;
  assign n10705 = ~n10702 & ~n10704 ;
  assign n10706 = n10696 & ~n10705 ;
  assign n10707 = ~n10701 & n10706 ;
  assign n10708 = ~n10698 & ~n10707 ;
  assign n10709 = n10695 & ~n10708 ;
  assign n10710 = n10426 & ~n10688 ;
  assign n10711 = \pi0152  & n10710 ;
  assign n10712 = ~\pi0210  & ~n10569 ;
  assign n10713 = \pi0152  & n10599 ;
  assign n10714 = ~n10712 & n10713 ;
  assign n10715 = ~n10711 & ~n10714 ;
  assign n10716 = \pi0152  & \pi0172  ;
  assign n10717 = ~n10373 & n10699 ;
  assign n10718 = ~\pi0032  & n10699 ;
  assign n10719 = ~n10634 & n10718 ;
  assign n10720 = ~n10717 & ~n10719 ;
  assign n10721 = \pi0095  & ~\pi0210  ;
  assign n10722 = ~n10182 & n10721 ;
  assign n10723 = n10432 & ~n10722 ;
  assign n10724 = ~n10642 & n10723 ;
  assign n10725 = n10720 & n10724 ;
  assign n10726 = ~n10710 & ~n10725 ;
  assign n10727 = \pi0172  & n10726 ;
  assign n10728 = ~n10716 & ~n10727 ;
  assign n10729 = n10715 & ~n10728 ;
  assign n10730 = n10696 & n10729 ;
  assign n10731 = ~n10368 & ~n10412 ;
  assign n10732 = ~n10363 & n10731 ;
  assign n10733 = n10411 & n10732 ;
  assign n10734 = ~n10482 & ~n10733 ;
  assign n10735 = ~n10700 & ~n10734 ;
  assign n10736 = n10260 & n10735 ;
  assign n10737 = \pi0152  & n10366 ;
  assign n10738 = ~n10688 & n10737 ;
  assign n10739 = ~\pi0172  & ~n10738 ;
  assign n10740 = ~n10736 & n10739 ;
  assign n10741 = n6706 & ~n10182 ;
  assign n10742 = ~\pi0210  & ~n10741 ;
  assign n10743 = ~n10569 & n10742 ;
  assign n10744 = \pi0152  & ~n10578 ;
  assign n10745 = n6706 & n10744 ;
  assign n10746 = ~n10743 & n10745 ;
  assign n10747 = ~\pi0152  & ~n10363 ;
  assign n10748 = ~n10642 & n10747 ;
  assign n10749 = \pi0172  & ~n10748 ;
  assign n10750 = n6706 & ~n10722 ;
  assign n10751 = n10720 & n10750 ;
  assign n10752 = \pi0172  & ~n10741 ;
  assign n10753 = ~n10751 & n10752 ;
  assign n10754 = ~n10749 & ~n10753 ;
  assign n10755 = ~n10746 & ~n10754 ;
  assign n10756 = ~n10740 & ~n10755 ;
  assign n10757 = ~\pi0158  & \pi0299  ;
  assign n10758 = ~n10710 & n10757 ;
  assign n10759 = ~n10756 & n10758 ;
  assign n10760 = ~n10730 & ~n10759 ;
  assign n10761 = ~n10709 & n10760 ;
  assign n10762 = ~\pi0149  & ~n10761 ;
  assign n10763 = ~\pi0152  & \pi0172  ;
  assign n10764 = \pi0172  & ~n10588 ;
  assign n10765 = \pi0172  & n10358 ;
  assign n10766 = ~n10362 & n10765 ;
  assign n10767 = ~n10764 & ~n10766 ;
  assign n10768 = ~n10426 & ~n10767 ;
  assign n10769 = ~\pi0210  & ~n10767 ;
  assign n10770 = ~n10375 & n10769 ;
  assign n10771 = ~n10768 & ~n10770 ;
  assign n10772 = ~n10763 & n10771 ;
  assign n10773 = ~n10363 & n10587 ;
  assign n10774 = ~n10426 & ~n10773 ;
  assign n10775 = ~\pi0210  & ~n10773 ;
  assign n10776 = ~n10375 & n10775 ;
  assign n10777 = ~n10774 & ~n10776 ;
  assign n10778 = ~\pi0152  & n10777 ;
  assign n10779 = n10757 & ~n10778 ;
  assign n10780 = ~n10772 & n10779 ;
  assign n10781 = ~n6706 & ~n10366 ;
  assign n10782 = ~\pi0210  & ~n6706 ;
  assign n10783 = ~n10375 & n10782 ;
  assign n10784 = ~n10781 & ~n10783 ;
  assign n10785 = ~\pi0172  & ~n10784 ;
  assign n10786 = n6706 & ~n10482 ;
  assign n10787 = ~n10481 & n10786 ;
  assign n10788 = \pi0152  & ~n10787 ;
  assign n10789 = ~\pi0152  & ~n6706 ;
  assign n10790 = ~n10456 & n10747 ;
  assign n10791 = ~n10789 & ~n10790 ;
  assign n10792 = ~\pi0172  & n10791 ;
  assign n10793 = ~n10788 & n10792 ;
  assign n10794 = ~n10785 & ~n10793 ;
  assign n10795 = n10757 & ~n10794 ;
  assign n10796 = ~n10780 & ~n10795 ;
  assign n10797 = ~n10385 & ~n10507 ;
  assign n10798 = ~n10426 & n10797 ;
  assign n10799 = ~\pi0210  & n10797 ;
  assign n10800 = ~n10375 & n10799 ;
  assign n10801 = ~n10798 & ~n10800 ;
  assign n10802 = n10697 & ~n10801 ;
  assign n10803 = ~\pi0210  & ~n10457 ;
  assign n10804 = ~n10375 & n10803 ;
  assign n10805 = ~n10458 & ~n10804 ;
  assign n10806 = ~\pi0152  & ~\pi0172  ;
  assign n10807 = ~n10805 & n10806 ;
  assign n10808 = ~n10802 & ~n10807 ;
  assign n10809 = ~\pi0040  & ~\pi0152  ;
  assign n10810 = n1256 & n10809 ;
  assign n10811 = ~n10789 & ~n10810 ;
  assign n10812 = n10784 & ~n10811 ;
  assign n10813 = \pi0172  & ~n10604 ;
  assign n10814 = ~n10426 & n10813 ;
  assign n10815 = ~\pi0210  & n10813 ;
  assign n10816 = ~n10375 & n10815 ;
  assign n10817 = ~n10814 & ~n10816 ;
  assign n10818 = ~n10763 & n10817 ;
  assign n10819 = ~n10812 & ~n10818 ;
  assign n10820 = n10808 & ~n10819 ;
  assign n10821 = n10696 & ~n10820 ;
  assign n10822 = n10796 & ~n10821 ;
  assign n10823 = \pi0149  & ~n10822 ;
  assign n10824 = ~n10762 & ~n10823 ;
  assign n10825 = ~n10687 & n10824 ;
  assign n10826 = \pi0232  & ~n10290 ;
  assign n10827 = ~n10213 & n10826 ;
  assign n10828 = ~n10825 & n10827 ;
  assign n10829 = ~n10381 & ~n10828 ;
  assign n10830 = \pi0100  & ~n10120 ;
  assign n10831 = ~\pi0087  & ~n10830 ;
  assign n10832 = \pi0075  & ~n10120 ;
  assign n10833 = \pi0038  & \pi0232  ;
  assign n10834 = n6706 & n10833 ;
  assign n10835 = n10105 & n10834 ;
  assign n10836 = ~\pi0100  & n10835 ;
  assign n10837 = ~n10830 & ~n10836 ;
  assign n10838 = ~n2619 & ~n10214 ;
  assign n10839 = n8640 & n10838 ;
  assign n10840 = n10175 & ~n10839 ;
  assign n10841 = n10174 & n10840 ;
  assign n10842 = n10173 & n10841 ;
  assign n10843 = n10837 & n10842 ;
  assign n10844 = n2327 & n10182 ;
  assign n10845 = ~n10836 & ~n10844 ;
  assign n10846 = ~n10830 & n10845 ;
  assign n10847 = n6895 & ~n10846 ;
  assign n10848 = ~n10843 & n10847 ;
  assign n10849 = ~n10832 & ~n10848 ;
  assign n10850 = n10831 & n10849 ;
  assign n10851 = ~n10829 & n10850 ;
  assign n10852 = \pi0087  & ~n10844 ;
  assign n10853 = ~n10836 & n10852 ;
  assign n10854 = ~n10830 & n10853 ;
  assign n10855 = n2364 & ~n10854 ;
  assign n10856 = ~n10832 & ~n10855 ;
  assign n10857 = ~n10848 & n10856 ;
  assign n10858 = n2511 & ~n10857 ;
  assign n10859 = ~n10193 & n10858 ;
  assign n10860 = ~n10851 & n10859 ;
  assign n10861 = ~n10194 & ~n10860 ;
  assign n10862 = ~\pi0055  & n10154 ;
  assign n10863 = ~n2467 & ~n10129 ;
  assign n10864 = ~n10131 & n10863 ;
  assign n10865 = n10143 & n10864 ;
  assign n10866 = n10147 & n10190 ;
  assign n10867 = ~n8601 & n10190 ;
  assign n10868 = ~n10117 & n10867 ;
  assign n10869 = ~n10866 & ~n10868 ;
  assign n10870 = ~n10167 & n10869 ;
  assign n10871 = \pi0149  & n1285 ;
  assign n10872 = n2855 & n10871 ;
  assign n10873 = n4520 & n10872 ;
  assign n10874 = n1638 & n10873 ;
  assign n10875 = ~n10133 & ~n10186 ;
  assign n10876 = ~n10167 & n10875 ;
  assign n10877 = ~n10874 & n10876 ;
  assign n10878 = ~n10870 & ~n10877 ;
  assign n10879 = ~n10865 & n10878 ;
  assign n10880 = ~n10862 & n10879 ;
  assign n10881 = ~n10199 & n10831 ;
  assign n10882 = ~n10211 & n10881 ;
  assign n10883 = \pi0038  & n10882 ;
  assign n10884 = n1256 & n1274 ;
  assign n10885 = n1273 & n10169 ;
  assign n10886 = ~\pi0053  & n10885 ;
  assign n10887 = n1340 & n10885 ;
  assign n10888 = n1249 & n10887 ;
  assign n10889 = ~n10886 & ~n10888 ;
  assign n10890 = n10884 & ~n10889 ;
  assign n10891 = ~n10325 & n10890 ;
  assign n10892 = ~n10322 & n10891 ;
  assign n10893 = n1327 & n8560 ;
  assign n10894 = \pi0090  & n7083 ;
  assign n10895 = n10893 & n10894 ;
  assign n10896 = n1319 & n10895 ;
  assign n10897 = n6637 & n10335 ;
  assign n10898 = n1358 & n10897 ;
  assign n10899 = ~n10896 & ~n10898 ;
  assign n10900 = ~\pi0070  & n10899 ;
  assign n10901 = ~n10892 & n10900 ;
  assign n10902 = ~\pi0051  & n1264 ;
  assign n10903 = n1263 & n10902 ;
  assign n10904 = ~n1864 & n10903 ;
  assign n10905 = n10483 & n10904 ;
  assign n10906 = ~n10901 & n10905 ;
  assign n10907 = n6967 & n6970 ;
  assign n10908 = n1354 & n10907 ;
  assign n10909 = n1358 & n10908 ;
  assign n10910 = \pi0032  & ~\pi0095  ;
  assign n10911 = n10909 & n10910 ;
  assign n10912 = ~\pi0070  & ~n10911 ;
  assign n10913 = ~n10892 & n10912 ;
  assign n10914 = ~n10904 & ~n10911 ;
  assign n10915 = \pi0183  & ~\pi0198  ;
  assign n10916 = n6706 & n10915 ;
  assign n10917 = ~n10914 & n10916 ;
  assign n10918 = ~n10913 & n10917 ;
  assign n10919 = ~n10906 & ~n10918 ;
  assign n10920 = n1319 & n10893 ;
  assign n10921 = \pi0090  & ~n10920 ;
  assign n10922 = n1618 & n7083 ;
  assign n10923 = ~n10921 & n10922 ;
  assign n10924 = n1256 & n10327 ;
  assign n10925 = n1273 & n10924 ;
  assign n10926 = n10318 & n10925 ;
  assign n10927 = n10316 & n10926 ;
  assign n10928 = ~\pi0090  & ~n10927 ;
  assign n10929 = ~n6638 & n10928 ;
  assign n10930 = ~\pi0040  & ~\pi0183  ;
  assign n10931 = n10414 & n10930 ;
  assign n10932 = ~n10929 & n10931 ;
  assign n10933 = n10923 & n10932 ;
  assign n10934 = \pi0193  & ~n10933 ;
  assign n10935 = n10919 & n10934 ;
  assign n10936 = n1256 & n10369 ;
  assign n10937 = n10468 & n10936 ;
  assign n10938 = n10931 & n10937 ;
  assign n10939 = n10319 & n10938 ;
  assign n10940 = ~\pi0193  & ~n10939 ;
  assign n10941 = ~\pi0174  & ~n10940 ;
  assign n10942 = ~\pi0070  & ~n6975 ;
  assign n10943 = ~n10892 & n10942 ;
  assign n10944 = ~n6975 & ~n10904 ;
  assign n10945 = ~\pi0174  & \pi0183  ;
  assign n10946 = n6706 & n10945 ;
  assign n10947 = ~n10944 & n10946 ;
  assign n10948 = ~n10943 & n10947 ;
  assign n10949 = ~n10941 & ~n10948 ;
  assign n10950 = ~n10935 & ~n10949 ;
  assign n10951 = n1274 & ~n10889 ;
  assign n10952 = ~n10389 & n10951 ;
  assign n10953 = n10899 & n10942 ;
  assign n10954 = ~n10952 & n10953 ;
  assign n10955 = ~n10944 & ~n10954 ;
  assign n10956 = n6706 & n10955 ;
  assign n10957 = \pi0183  & ~\pi0193  ;
  assign n10958 = n6706 & n10957 ;
  assign n10959 = n10903 & n10958 ;
  assign n10960 = ~n1864 & n10959 ;
  assign n10961 = n6975 & n10958 ;
  assign n10962 = ~n10960 & ~n10961 ;
  assign n10963 = ~\pi0070  & ~n10961 ;
  assign n10964 = ~n10952 & n10963 ;
  assign n10965 = ~n10962 & ~n10964 ;
  assign n10966 = \pi0183  & ~n10965 ;
  assign n10967 = ~n10956 & n10966 ;
  assign n10968 = ~\pi0070  & ~n10952 ;
  assign n10969 = n10960 & ~n10968 ;
  assign n10970 = ~\pi0193  & ~n10961 ;
  assign n10971 = ~\pi0040  & n10414 ;
  assign n10972 = n1618 & n10971 ;
  assign n10973 = ~n10899 & n10972 ;
  assign n10974 = ~\pi0183  & ~n10961 ;
  assign n10975 = ~n10973 & n10974 ;
  assign n10976 = ~n10970 & ~n10975 ;
  assign n10977 = ~n10969 & ~n10976 ;
  assign n10978 = \pi0174  & ~n10977 ;
  assign n10979 = ~n10967 & n10978 ;
  assign n10980 = n1979 & n6706 ;
  assign n10981 = ~\pi0035  & n1354 ;
  assign n10982 = n10980 & n10981 ;
  assign n10983 = n1358 & n10982 ;
  assign n10984 = ~\pi0040  & \pi0180  ;
  assign n10985 = n10983 & n10984 ;
  assign n10986 = ~\pi0299  & ~n10985 ;
  assign n10987 = ~n10979 & n10986 ;
  assign n10988 = ~n10950 & n10987 ;
  assign n10989 = ~\pi0040  & \pi0158  ;
  assign n10990 = n10983 & n10989 ;
  assign n10991 = \pi0299  & ~n10990 ;
  assign n10992 = n8364 & ~n10991 ;
  assign n10993 = ~\pi0152  & n10971 ;
  assign n10994 = ~n10929 & n10993 ;
  assign n10995 = n10923 & n10994 ;
  assign n10996 = \pi0172  & ~n10973 ;
  assign n10997 = ~n10995 & n10996 ;
  assign n10998 = n10414 & n10809 ;
  assign n10999 = n10937 & n10998 ;
  assign n11000 = n10319 & n10999 ;
  assign n11001 = ~\pi0172  & ~n11000 ;
  assign n11002 = ~\pi0149  & ~n11001 ;
  assign n11003 = n8364 & n11002 ;
  assign n11004 = ~n10997 & n11003 ;
  assign n11005 = ~n10992 & ~n11004 ;
  assign n11006 = \pi0172  & n10903 ;
  assign n11007 = ~n1864 & n11006 ;
  assign n11008 = ~n10901 & n11007 ;
  assign n11009 = ~n7151 & ~n10904 ;
  assign n11010 = ~\pi0070  & ~n7151 ;
  assign n11011 = ~n10892 & n11010 ;
  assign n11012 = ~n11009 & ~n11011 ;
  assign n11013 = ~n11008 & ~n11012 ;
  assign n11014 = ~\pi0152  & n11013 ;
  assign n11015 = n10900 & ~n10952 ;
  assign n11016 = n11007 & ~n11015 ;
  assign n11017 = \pi0152  & ~n7151 ;
  assign n11018 = ~n10904 & n11017 ;
  assign n11019 = ~\pi0070  & n11017 ;
  assign n11020 = ~n10952 & n11019 ;
  assign n11021 = ~n11018 & ~n11020 ;
  assign n11022 = ~n11016 & ~n11021 ;
  assign n11023 = \pi0149  & n8364 ;
  assign n11024 = n6706 & n11023 ;
  assign n11025 = ~n11022 & n11024 ;
  assign n11026 = ~n11014 & n11025 ;
  assign n11027 = n11005 & ~n11026 ;
  assign n11028 = ~n10988 & ~n11027 ;
  assign n11029 = ~\pi0174  & n6706 ;
  assign n11030 = n6955 & n11029 ;
  assign n11031 = ~n6761 & n11030 ;
  assign n11032 = n6954 & n11031 ;
  assign n11033 = \pi0174  & \pi1091  ;
  assign n11034 = n1689 & n11033 ;
  assign n11035 = n1688 & n11034 ;
  assign n11036 = n10242 & n11035 ;
  assign n11037 = n6921 & n11036 ;
  assign n11038 = \pi0176  & ~n11037 ;
  assign n11039 = ~n11032 & n11038 ;
  assign n11040 = \pi0039  & \pi0232  ;
  assign n11041 = ~n10214 & n11040 ;
  assign n11042 = ~\pi0174  & n11040 ;
  assign n11043 = n10242 & n11042 ;
  assign n11044 = n6948 & n11043 ;
  assign n11045 = ~n11041 & ~n11044 ;
  assign n11046 = ~\pi0299  & ~n11045 ;
  assign n11047 = ~n11039 & n11046 ;
  assign n11048 = n6743 & n6954 ;
  assign n11049 = \pi0154  & ~n11048 ;
  assign n11050 = ~\pi0152  & \pi0154  ;
  assign n11051 = ~\pi0152  & n6743 ;
  assign n11052 = n6948 & n11051 ;
  assign n11053 = ~n11050 & ~n11052 ;
  assign n11054 = ~n11049 & ~n11053 ;
  assign n11055 = n1696 & n6743 ;
  assign n11056 = \pi0152  & \pi0154  ;
  assign n11057 = n1259 & n11056 ;
  assign n11058 = n1249 & n11057 ;
  assign n11059 = n6920 & n11058 ;
  assign n11060 = n11055 & n11059 ;
  assign n11061 = ~n11054 & ~n11060 ;
  assign n11062 = n2256 & n6746 ;
  assign n11063 = ~n11045 & n11062 ;
  assign n11064 = ~n11061 & n11063 ;
  assign n11065 = ~n11047 & ~n11064 ;
  assign n11066 = n10882 & n11065 ;
  assign n11067 = ~n11028 & n11066 ;
  assign n11068 = ~n10883 & ~n11067 ;
  assign n11069 = \pi0087  & ~n10835 ;
  assign n11070 = ~\pi0100  & ~n11069 ;
  assign n11071 = n7265 & n11070 ;
  assign n11072 = \pi0100  & n7265 ;
  assign n11073 = ~n10120 & n11072 ;
  assign n11074 = ~n11071 & ~n11073 ;
  assign n11075 = n11068 & ~n11074 ;
  assign n11076 = n2363 & n10839 ;
  assign n11077 = n4520 & n11076 ;
  assign n11078 = n1638 & n11077 ;
  assign n11079 = ~n10832 & n10837 ;
  assign n11080 = ~n11078 & n11079 ;
  assign n11081 = ~\pi0054  & n6895 ;
  assign n11082 = ~\pi0054  & \pi0075  ;
  assign n11083 = ~n10120 & n11082 ;
  assign n11084 = ~n11081 & ~n11083 ;
  assign n11085 = ~n11080 & ~n11084 ;
  assign n11086 = n10123 & ~n11085 ;
  assign n11087 = ~n11075 & n11086 ;
  assign n11088 = ~\pi0074  & n10879 ;
  assign n11089 = ~n11087 & n11088 ;
  assign n11090 = ~n10880 & ~n11089 ;
  assign n11091 = n10146 & ~n10865 ;
  assign n11092 = \pi0033  & ~n11091 ;
  assign n11093 = n11090 & n11092 ;
  assign n11094 = \pi0954  & ~n10865 ;
  assign n11095 = ~n11093 & n11094 ;
  assign n11096 = ~n10861 & n11095 ;
  assign n11097 = ~\pi0034  & ~\pi0118  ;
  assign n11098 = ~\pi0079  & n11097 ;
  assign n11099 = ~\pi0195  & ~\pi0196  ;
  assign n11100 = ~\pi0138  & ~\pi0139  ;
  assign n11101 = n11099 & n11100 ;
  assign n11102 = n11098 & n11101 ;
  assign n11103 = ~\pi0033  & ~n11102 ;
  assign n11104 = ~n11091 & n11103 ;
  assign n11105 = n11090 & n11104 ;
  assign n11106 = ~\pi0954  & ~n10865 ;
  assign n11107 = ~n11105 & n11106 ;
  assign n11108 = ~n10861 & n11107 ;
  assign n11109 = n11090 & ~n11091 ;
  assign n11110 = ~\pi0954  & n11103 ;
  assign n11111 = ~n11109 & n11110 ;
  assign n11112 = \pi0033  & \pi0954  ;
  assign n11113 = ~n11109 & n11112 ;
  assign n11114 = ~n11111 & ~n11113 ;
  assign n11115 = ~n11108 & n11114 ;
  assign n11116 = ~n11096 & n11115 ;
  assign n11117 = \pi0197  & n10114 ;
  assign n11118 = ~\pi0197  & ~n10114 ;
  assign n11119 = ~n11117 & ~n11118 ;
  assign n11120 = \pi0162  & n6706 ;
  assign n11121 = n11117 & n11120 ;
  assign n11122 = n6706 & n10114 ;
  assign n11123 = ~\pi0162  & ~\pi0197  ;
  assign n11124 = n6706 & n11123 ;
  assign n11125 = ~n11122 & ~n11124 ;
  assign n11126 = ~n11121 & ~n11125 ;
  assign n11127 = ~n11119 & ~n11126 ;
  assign n11128 = n11119 & ~n11120 ;
  assign n11129 = \pi0232  & ~n8601 ;
  assign n11130 = ~n11128 & n11129 ;
  assign n11131 = ~n11127 & n11130 ;
  assign n11132 = ~\pi0074  & \pi0167  ;
  assign n11133 = n8601 & n11132 ;
  assign n11134 = n8640 & n11133 ;
  assign n11135 = \pi0148  & \pi0232  ;
  assign n11136 = n6706 & n11135 ;
  assign n11137 = n10139 & n11136 ;
  assign n11138 = ~n11134 & ~n11137 ;
  assign n11139 = \pi0167  & \pi0232  ;
  assign n11140 = n6706 & n11139 ;
  assign n11141 = \pi0038  & n8601 ;
  assign n11142 = n11140 & n11141 ;
  assign n11143 = ~n11138 & n11142 ;
  assign n11144 = ~n2511 & ~n11138 ;
  assign n11145 = ~n11143 & ~n11144 ;
  assign n11146 = ~n11131 & n11145 ;
  assign n11147 = ~n1292 & n11146 ;
  assign n11148 = n2467 & ~n11147 ;
  assign n11149 = ~n1292 & ~n10158 ;
  assign n11150 = n2467 & ~n11149 ;
  assign n11151 = ~n11148 & ~n11150 ;
  assign n11152 = \pi0299  & n11128 ;
  assign n11153 = \pi0299  & ~n11119 ;
  assign n11154 = ~n11126 & n11153 ;
  assign n11155 = ~n11152 & ~n11154 ;
  assign n11156 = \pi0140  & \pi0145  ;
  assign n11157 = ~\pi0140  & ~\pi0145  ;
  assign n11158 = ~n11156 & ~n11157 ;
  assign n11159 = n10111 & ~n11158 ;
  assign n11160 = n10110 & ~n11156 ;
  assign n11161 = n6706 & ~n11157 ;
  assign n11162 = n11160 & n11161 ;
  assign n11163 = ~n11159 & ~n11162 ;
  assign n11164 = ~\pi0299  & n11163 ;
  assign n11165 = n11129 & ~n11164 ;
  assign n11166 = n11155 & n11165 ;
  assign n11167 = \pi0141  & ~\pi0299  ;
  assign n11168 = \pi0148  & \pi0299  ;
  assign n11169 = ~n11167 & ~n11168 ;
  assign n11170 = n8640 & ~n11169 ;
  assign n11171 = n8601 & n11170 ;
  assign n11172 = \pi0074  & ~n11171 ;
  assign n11173 = ~n11166 & n11172 ;
  assign n11174 = ~\pi0055  & ~n11173 ;
  assign n11175 = n8601 & n11136 ;
  assign n11176 = \pi0074  & ~n11175 ;
  assign n11177 = n1292 & n11176 ;
  assign n11178 = ~n11131 & n11177 ;
  assign n11179 = ~n1293 & ~n11178 ;
  assign n11180 = \pi0162  & \pi0232  ;
  assign n11181 = n6706 & n11180 ;
  assign n11182 = ~\pi0092  & ~n11181 ;
  assign n11183 = n10176 & n11182 ;
  assign n11184 = n10173 & n11183 ;
  assign n11185 = \pi0054  & ~n11140 ;
  assign n11186 = n8601 & ~n11185 ;
  assign n11187 = n10156 & n11186 ;
  assign n11188 = ~n11184 & n11187 ;
  assign n11189 = \pi0054  & n8601 ;
  assign n11190 = n11140 & n11189 ;
  assign n11191 = ~n11142 & ~n11190 ;
  assign n11192 = n10190 & n11191 ;
  assign n11193 = ~n11131 & n11192 ;
  assign n11194 = ~n11188 & n11193 ;
  assign n11195 = n11179 & ~n11194 ;
  assign n11196 = ~n11174 & ~n11195 ;
  assign n11197 = ~\pi0142  & n10428 ;
  assign n11198 = ~\pi0142  & n10496 ;
  assign n11199 = ~n10671 & n11198 ;
  assign n11200 = ~n11197 & ~n11199 ;
  assign n11201 = ~\pi0140  & ~\pi0142  ;
  assign n11202 = ~\pi0140  & ~n10428 ;
  assign n11203 = ~n10423 & n11202 ;
  assign n11204 = ~n11201 & ~n11203 ;
  assign n11205 = n11200 & ~n11204 ;
  assign n11206 = ~n10375 & n10570 ;
  assign n11207 = ~n10781 & ~n11206 ;
  assign n11208 = ~\pi0142  & ~n6706 ;
  assign n11209 = ~\pi0040  & ~\pi0142  ;
  assign n11210 = n1256 & n11209 ;
  assign n11211 = ~n11208 & ~n11210 ;
  assign n11212 = n11207 & ~n11211 ;
  assign n11213 = \pi0140  & ~\pi0142  ;
  assign n11214 = \pi0140  & ~n10457 ;
  assign n11215 = ~n10426 & n11214 ;
  assign n11216 = ~\pi0198  & n11214 ;
  assign n11217 = ~n10375 & n11216 ;
  assign n11218 = ~n11215 & ~n11217 ;
  assign n11219 = ~n11213 & n11218 ;
  assign n11220 = ~n11212 & ~n11219 ;
  assign n11221 = \pi0181  & ~n11220 ;
  assign n11222 = ~n11205 & n11221 ;
  assign n11223 = \pi0095  & \pi0140  ;
  assign n11224 = ~n10357 & n11223 ;
  assign n11225 = ~n10362 & n11224 ;
  assign n11226 = ~\pi0095  & \pi0140  ;
  assign n11227 = ~n10182 & n11226 ;
  assign n11228 = ~\pi0142  & ~n11227 ;
  assign n11229 = ~n11225 & n11228 ;
  assign n11230 = ~n10363 & n11229 ;
  assign n11231 = ~n10642 & n11230 ;
  assign n11232 = n10637 & n11231 ;
  assign n11233 = ~n10586 & n11213 ;
  assign n11234 = ~n11225 & n11233 ;
  assign n11235 = n6706 & ~n11234 ;
  assign n11236 = ~n11232 & n11235 ;
  assign n11237 = ~\pi0181  & n11207 ;
  assign n11238 = ~n11236 & n11237 ;
  assign n11239 = ~n10422 & ~n10734 ;
  assign n11240 = ~\pi0140  & ~n11239 ;
  assign n11241 = ~n10454 & n11226 ;
  assign n11242 = ~n10449 & n11241 ;
  assign n11243 = \pi0140  & n10358 ;
  assign n11244 = ~n10362 & n11243 ;
  assign n11245 = \pi0142  & ~n11244 ;
  assign n11246 = ~n11242 & n11245 ;
  assign n11247 = n11237 & n11246 ;
  assign n11248 = ~n11240 & n11247 ;
  assign n11249 = ~n11238 & ~n11248 ;
  assign n11250 = ~\pi0144  & ~\pi0299  ;
  assign n11251 = n11249 & n11250 ;
  assign n11252 = ~n11222 & n11251 ;
  assign n11253 = ~\pi0142  & n10599 ;
  assign n11254 = ~n10600 & n11253 ;
  assign n11255 = ~n11197 & ~n11254 ;
  assign n11256 = \pi0142  & ~n10503 ;
  assign n11257 = ~\pi0140  & ~n11256 ;
  assign n11258 = n11255 & n11257 ;
  assign n11259 = ~\pi0198  & n10797 ;
  assign n11260 = ~n10375 & n11259 ;
  assign n11261 = ~n10798 & ~n11260 ;
  assign n11262 = \pi0140  & \pi0142  ;
  assign n11263 = ~n11261 & n11262 ;
  assign n11264 = ~n10608 & n11213 ;
  assign n11265 = ~n11263 & ~n11264 ;
  assign n11266 = \pi0181  & n11265 ;
  assign n11267 = ~n11258 & n11266 ;
  assign n11268 = \pi0144  & ~n11267 ;
  assign n11269 = \pi0142  & ~n10364 ;
  assign n11270 = ~n10363 & n11269 ;
  assign n11271 = n10355 & n11270 ;
  assign n11272 = ~\pi0140  & ~n11271 ;
  assign n11273 = ~\pi0140  & ~\pi0198  ;
  assign n11274 = ~n10375 & n11273 ;
  assign n11275 = ~n11272 & ~n11274 ;
  assign n11276 = \pi0142  & ~n11275 ;
  assign n11277 = ~n10428 & ~n11275 ;
  assign n11278 = ~n10580 & n11277 ;
  assign n11279 = ~n11276 & ~n11278 ;
  assign n11280 = ~n10363 & n10588 ;
  assign n11281 = ~n10426 & ~n11280 ;
  assign n11282 = ~\pi0198  & ~n11280 ;
  assign n11283 = ~n10375 & n11282 ;
  assign n11284 = ~n11281 & ~n11283 ;
  assign n11285 = ~\pi0142  & n11284 ;
  assign n11286 = \pi0142  & ~n10787 ;
  assign n11287 = n11207 & n11286 ;
  assign n11288 = \pi0140  & ~n11287 ;
  assign n11289 = ~n11285 & n11288 ;
  assign n11290 = ~\pi0181  & ~n11289 ;
  assign n11291 = n11279 & n11290 ;
  assign n11292 = ~\pi0299  & ~n11291 ;
  assign n11293 = n11268 & n11292 ;
  assign n11294 = ~n11252 & ~n11293 ;
  assign n11295 = \pi0146  & ~\pi0161  ;
  assign n11296 = ~\pi0161  & ~n10773 ;
  assign n11297 = ~n10426 & n11296 ;
  assign n11298 = ~\pi0210  & n11296 ;
  assign n11299 = ~n10375 & n11298 ;
  assign n11300 = ~n11297 & ~n11299 ;
  assign n11301 = ~n11295 & n11300 ;
  assign n11302 = ~\pi0159  & \pi0299  ;
  assign n11303 = \pi0146  & ~n6706 ;
  assign n11304 = \pi0146  & ~n10363 ;
  assign n11305 = ~n10456 & n11304 ;
  assign n11306 = ~n11303 & ~n11305 ;
  assign n11307 = n10784 & ~n11306 ;
  assign n11308 = n11302 & ~n11307 ;
  assign n11309 = ~n11301 & n11308 ;
  assign n11310 = \pi0146  & ~n10787 ;
  assign n11311 = n10784 & n11310 ;
  assign n11312 = \pi0161  & ~n11311 ;
  assign n11313 = ~\pi0210  & ~n11280 ;
  assign n11314 = ~n10375 & n11313 ;
  assign n11315 = ~n11281 & ~n11314 ;
  assign n11316 = ~\pi0146  & n11315 ;
  assign n11317 = n11302 & ~n11316 ;
  assign n11318 = n11312 & n11317 ;
  assign n11319 = ~n11309 & ~n11318 ;
  assign n11320 = \pi0146  & \pi0161  ;
  assign n11321 = \pi0161  & ~n10604 ;
  assign n11322 = ~n10426 & n11321 ;
  assign n11323 = ~\pi0210  & n11321 ;
  assign n11324 = ~n10375 & n11323 ;
  assign n11325 = ~n11322 & ~n11324 ;
  assign n11326 = ~n11320 & n11325 ;
  assign n11327 = \pi0159  & \pi0299  ;
  assign n11328 = \pi0146  & n10801 ;
  assign n11329 = n11327 & ~n11328 ;
  assign n11330 = ~n11326 & n11329 ;
  assign n11331 = ~\pi0146  & ~n6706 ;
  assign n11332 = ~\pi0040  & ~\pi0146  ;
  assign n11333 = n1256 & n11332 ;
  assign n11334 = ~n11331 & ~n11333 ;
  assign n11335 = n10784 & ~n11334 ;
  assign n11336 = ~\pi0161  & ~n11335 ;
  assign n11337 = \pi0146  & n10805 ;
  assign n11338 = n11327 & ~n11337 ;
  assign n11339 = n11336 & n11338 ;
  assign n11340 = ~n11330 & ~n11339 ;
  assign n11341 = n11319 & n11340 ;
  assign n11342 = \pi0162  & ~n11341 ;
  assign n11343 = n6706 & n11295 ;
  assign n11344 = n10735 & n11343 ;
  assign n11345 = n10366 & n11320 ;
  assign n11346 = ~n10688 & n11345 ;
  assign n11347 = ~n10710 & n11302 ;
  assign n11348 = ~n11346 & n11347 ;
  assign n11349 = ~n11344 & n11348 ;
  assign n11350 = ~\pi0161  & ~n10741 ;
  assign n11351 = ~n10751 & n11350 ;
  assign n11352 = ~\pi0161  & n10363 ;
  assign n11353 = ~\pi0161  & n10641 ;
  assign n11354 = ~n10639 & n11353 ;
  assign n11355 = ~n11352 & ~n11354 ;
  assign n11356 = ~\pi0146  & n11355 ;
  assign n11357 = ~n11351 & n11356 ;
  assign n11358 = ~\pi0162  & ~n11357 ;
  assign n11359 = n10579 & ~n10743 ;
  assign n11360 = \pi0161  & ~\pi0162  ;
  assign n11361 = ~n11359 & n11360 ;
  assign n11362 = ~n11358 & ~n11361 ;
  assign n11363 = n11349 & ~n11362 ;
  assign n11364 = ~\pi0146  & ~n10726 ;
  assign n11365 = ~\pi0146  & ~\pi0161  ;
  assign n11366 = ~\pi0161  & ~n10710 ;
  assign n11367 = ~n10701 & n11366 ;
  assign n11368 = ~n11365 & ~n11367 ;
  assign n11369 = ~n11364 & ~n11368 ;
  assign n11370 = ~\pi0146  & n10710 ;
  assign n11371 = ~\pi0146  & n10599 ;
  assign n11372 = ~n10712 & n11371 ;
  assign n11373 = ~n11370 & ~n11372 ;
  assign n11374 = \pi0146  & n10426 ;
  assign n11375 = ~n10688 & n11374 ;
  assign n11376 = \pi0146  & n6706 ;
  assign n11377 = n10692 & n11376 ;
  assign n11378 = ~n10688 & n11377 ;
  assign n11379 = \pi0161  & ~n11378 ;
  assign n11380 = ~n11375 & n11379 ;
  assign n11381 = n11373 & n11380 ;
  assign n11382 = ~n11369 & ~n11381 ;
  assign n11383 = ~\pi0162  & n11327 ;
  assign n11384 = ~n11382 & n11383 ;
  assign n11385 = ~n11363 & ~n11384 ;
  assign n11386 = ~n11342 & n11385 ;
  assign n11387 = n11294 & n11386 ;
  assign n11388 = \pi0232  & n1288 ;
  assign n11389 = ~n11387 & n11388 ;
  assign n11390 = ~\pi0167  & ~n10195 ;
  assign n11391 = ~\pi0167  & n4520 ;
  assign n11392 = n1638 & n11391 ;
  assign n11393 = ~n11390 & ~n11392 ;
  assign n11394 = \pi0167  & n6784 ;
  assign n11395 = n1266 & n11394 ;
  assign n11396 = n1354 & n11395 ;
  assign n11397 = n1358 & n11396 ;
  assign n11398 = \pi0167  & ~n8640 ;
  assign n11399 = \pi0188  & ~n11398 ;
  assign n11400 = ~n11397 & n11399 ;
  assign n11401 = n11393 & n11400 ;
  assign n11402 = ~\pi0188  & n11140 ;
  assign n11403 = \pi0299  & n11402 ;
  assign n11404 = ~n8375 & n11403 ;
  assign n11405 = \pi0038  & ~n11404 ;
  assign n11406 = ~n11401 & n11405 ;
  assign n11407 = ~\pi0039  & ~\pi0087  ;
  assign n11408 = ~n11406 & n11407 ;
  assign n11409 = ~\pi0038  & ~\pi0155  ;
  assign n11410 = ~n7597 & n11409 ;
  assign n11411 = ~\pi0161  & n6706 ;
  assign n11412 = n10182 & n11411 ;
  assign n11413 = ~n10259 & n11412 ;
  assign n11414 = n11409 & ~n11413 ;
  assign n11415 = ~n10256 & n11414 ;
  assign n11416 = ~n11410 & ~n11415 ;
  assign n11417 = ~\pi0038  & \pi0155  ;
  assign n11418 = \pi0161  & n6706 ;
  assign n11419 = ~n6732 & n11418 ;
  assign n11420 = ~n10267 & n11419 ;
  assign n11421 = n7597 & n10182 ;
  assign n11422 = ~n10233 & n11421 ;
  assign n11423 = ~n11420 & n11422 ;
  assign n11424 = n11417 & ~n11423 ;
  assign n11425 = n11416 & ~n11424 ;
  assign n11426 = \pi0232  & n10280 ;
  assign n11427 = ~n11425 & n11426 ;
  assign n11428 = ~n10239 & ~n10247 ;
  assign n11429 = ~\pi0144  & n10220 ;
  assign n11430 = ~\pi0144  & n10182 ;
  assign n11431 = ~n10233 & n11430 ;
  assign n11432 = ~n11429 & ~n11431 ;
  assign n11433 = \pi0177  & n11432 ;
  assign n11434 = ~n11428 & n11433 ;
  assign n11435 = n9636 & n11434 ;
  assign n11436 = ~n10220 & ~n10284 ;
  assign n11437 = \pi0144  & n10220 ;
  assign n11438 = \pi0144  & n10182 ;
  assign n11439 = ~n10233 & n11438 ;
  assign n11440 = ~n11437 & ~n11439 ;
  assign n11441 = ~n11436 & ~n11440 ;
  assign n11442 = n10219 & n10221 ;
  assign n11443 = n10182 & ~n11442 ;
  assign n11444 = ~n11432 & n11443 ;
  assign n11445 = ~n11441 & ~n11444 ;
  assign n11446 = ~\pi0177  & ~\pi0299  ;
  assign n11447 = n9636 & n11446 ;
  assign n11448 = n11445 & n11447 ;
  assign n11449 = ~n11435 & ~n11448 ;
  assign n11450 = ~n11427 & n11449 ;
  assign n11451 = ~\pi0087  & ~n11406 ;
  assign n11452 = ~\pi0038  & ~\pi0232  ;
  assign n11453 = ~n10287 & n11452 ;
  assign n11454 = n11451 & ~n11453 ;
  assign n11455 = n11450 & n11454 ;
  assign n11456 = ~n11408 & ~n11455 ;
  assign n11457 = n1288 & ~n10378 ;
  assign n11458 = ~\pi0100  & ~n11457 ;
  assign n11459 = ~n11456 & n11458 ;
  assign n11460 = ~n11389 & n11459 ;
  assign n11461 = \pi0100  & \pi0232  ;
  assign n11462 = ~n11164 & n11461 ;
  assign n11463 = n11155 & n11462 ;
  assign n11464 = n2364 & ~n11463 ;
  assign n11465 = \pi0188  & ~\pi0299  ;
  assign n11466 = \pi0167  & \pi0299  ;
  assign n11467 = ~n11465 & ~n11466 ;
  assign n11468 = n10834 & ~n11467 ;
  assign n11469 = ~n10156 & ~n11468 ;
  assign n11470 = \pi0087  & ~\pi0100  ;
  assign n11471 = ~n11469 & n11470 ;
  assign n11472 = ~\pi0054  & ~n11471 ;
  assign n11473 = n11464 & n11472 ;
  assign n11474 = ~n11460 & n11473 ;
  assign n11475 = \pi0232  & ~n11164 ;
  assign n11476 = n11155 & n11475 ;
  assign n11477 = \pi0075  & ~n11476 ;
  assign n11478 = \pi0177  & ~\pi0299  ;
  assign n11479 = \pi0155  & \pi0299  ;
  assign n11480 = ~n11478 & ~n11479 ;
  assign n11481 = ~\pi0038  & n11480 ;
  assign n11482 = n8640 & ~n11481 ;
  assign n11483 = n10176 & ~n11482 ;
  assign n11484 = n10173 & n11483 ;
  assign n11485 = ~\pi0100  & ~n11469 ;
  assign n11486 = ~n11484 & n11485 ;
  assign n11487 = ~n11477 & n11486 ;
  assign n11488 = n6895 & ~n11463 ;
  assign n11489 = ~n11477 & ~n11488 ;
  assign n11490 = ~\pi0054  & ~n11489 ;
  assign n11491 = ~n11487 & n11490 ;
  assign n11492 = n8640 & ~n11467 ;
  assign n11493 = n8601 & n11492 ;
  assign n11494 = \pi0054  & ~n11493 ;
  assign n11495 = ~n11166 & n11494 ;
  assign n11496 = ~n11491 & ~n11495 ;
  assign n11497 = ~n11474 & n11496 ;
  assign n11498 = ~\pi0074  & ~n11195 ;
  assign n11499 = ~n11497 & n11498 ;
  assign n11500 = ~n11196 & ~n11499 ;
  assign n11501 = ~n11151 & n11500 ;
  assign n11502 = ~n11131 & n11138 ;
  assign n11503 = ~n2467 & ~n11502 ;
  assign n11504 = ~\pi0034  & ~n11503 ;
  assign n11505 = ~n11501 & n11504 ;
  assign n11506 = ~\pi0033  & ~\pi0954  ;
  assign n11507 = ~\pi0040  & \pi0181  ;
  assign n11508 = n10983 & n11507 ;
  assign n11509 = ~\pi0299  & ~n11508 ;
  assign n11510 = \pi0144  & ~n6975 ;
  assign n11511 = n10904 & ~n10968 ;
  assign n11512 = ~\pi0142  & n10903 ;
  assign n11513 = ~n1864 & n11512 ;
  assign n11514 = ~n11015 & n11513 ;
  assign n11515 = ~n11511 & ~n11514 ;
  assign n11516 = n11510 & n11515 ;
  assign n11517 = n6706 & ~n11516 ;
  assign n11518 = \pi0140  & ~n11517 ;
  assign n11519 = ~\pi0144  & n10944 ;
  assign n11520 = ~\pi0144  & n10942 ;
  assign n11521 = ~n10892 & n11520 ;
  assign n11522 = ~n11519 & ~n11521 ;
  assign n11523 = ~\pi0142  & n10904 ;
  assign n11524 = ~n10901 & n11523 ;
  assign n11525 = \pi0140  & ~n11524 ;
  assign n11526 = ~n11522 & n11525 ;
  assign n11527 = ~n10929 & n10971 ;
  assign n11528 = n10923 & n11527 ;
  assign n11529 = ~\pi0142  & ~n11528 ;
  assign n11530 = n1264 & n10496 ;
  assign n11531 = n10937 & n11530 ;
  assign n11532 = n10319 & n11531 ;
  assign n11533 = \pi0142  & ~n11532 ;
  assign n11534 = ~\pi0144  & ~n11533 ;
  assign n11535 = ~n11529 & n11534 ;
  assign n11536 = ~\pi0142  & \pi0144  ;
  assign n11537 = n1618 & n11536 ;
  assign n11538 = n10971 & n11537 ;
  assign n11539 = ~n10899 & n11538 ;
  assign n11540 = ~\pi0140  & ~n11539 ;
  assign n11541 = ~n11535 & n11540 ;
  assign n11542 = ~n11526 & ~n11541 ;
  assign n11543 = ~n11518 & n11542 ;
  assign n11544 = n11509 & ~n11543 ;
  assign n11545 = \pi0159  & n1983 ;
  assign n11546 = ~\pi0162  & ~n11545 ;
  assign n11547 = ~\pi0146  & n10903 ;
  assign n11548 = ~n1864 & n11547 ;
  assign n11549 = ~n11015 & n11548 ;
  assign n11550 = ~n11511 & ~n11549 ;
  assign n11551 = \pi0161  & ~n7151 ;
  assign n11552 = ~n11545 & n11551 ;
  assign n11553 = n11550 & n11552 ;
  assign n11554 = ~n11546 & ~n11553 ;
  assign n11555 = ~\pi0161  & n11009 ;
  assign n11556 = ~\pi0161  & n11010 ;
  assign n11557 = ~n10892 & n11556 ;
  assign n11558 = ~n11555 & ~n11557 ;
  assign n11559 = ~n11545 & ~n11548 ;
  assign n11560 = n10900 & ~n11545 ;
  assign n11561 = ~n10892 & n11560 ;
  assign n11562 = ~n11559 & ~n11561 ;
  assign n11563 = ~n11558 & ~n11562 ;
  assign n11564 = n6706 & ~n11563 ;
  assign n11565 = n11554 & n11564 ;
  assign n11566 = ~\pi0146  & \pi0161  ;
  assign n11567 = n1618 & n11566 ;
  assign n11568 = n10971 & n11567 ;
  assign n11569 = ~n10899 & n11568 ;
  assign n11570 = ~\pi0146  & ~n11569 ;
  assign n11571 = ~n11528 & n11570 ;
  assign n11572 = \pi0146  & ~n11532 ;
  assign n11573 = ~\pi0161  & ~n11572 ;
  assign n11574 = ~n11569 & ~n11573 ;
  assign n11575 = ~\pi0162  & ~n11574 ;
  assign n11576 = ~n11571 & n11575 ;
  assign n11577 = \pi0299  & ~n11576 ;
  assign n11578 = ~n11565 & n11577 ;
  assign n11579 = \pi0232  & ~n11578 ;
  assign n11580 = ~n11544 & n11579 ;
  assign n11581 = \pi0087  & n11468 ;
  assign n11582 = n1288 & ~n11581 ;
  assign n11583 = ~n11580 & n11582 ;
  assign n11584 = ~n11451 & ~n11581 ;
  assign n11585 = ~\pi0161  & n7597 ;
  assign n11586 = n6743 & n11585 ;
  assign n11587 = n6948 & n11586 ;
  assign n11588 = \pi0299  & n11409 ;
  assign n11589 = ~n11587 & n11588 ;
  assign n11590 = n1259 & n6743 ;
  assign n11591 = n1249 & n11590 ;
  assign n11592 = n6920 & n11591 ;
  assign n11593 = n1696 & n11592 ;
  assign n11594 = \pi0161  & n7597 ;
  assign n11595 = n11593 & n11594 ;
  assign n11596 = n11048 & n11585 ;
  assign n11597 = ~n11595 & ~n11596 ;
  assign n11598 = \pi0299  & n11417 ;
  assign n11599 = n11597 & n11598 ;
  assign n11600 = ~n11589 & ~n11599 ;
  assign n11601 = \pi0232  & ~n11446 ;
  assign n11602 = ~\pi0144  & \pi0232  ;
  assign n11603 = n10242 & n11602 ;
  assign n11604 = n6948 & n11603 ;
  assign n11605 = ~n11601 & ~n11604 ;
  assign n11606 = ~\pi0038  & n11605 ;
  assign n11607 = \pi0144  & \pi1091  ;
  assign n11608 = n1689 & n11607 ;
  assign n11609 = n1688 & n11608 ;
  assign n11610 = n1259 & n10242 ;
  assign n11611 = n1249 & n11610 ;
  assign n11612 = n6920 & n11611 ;
  assign n11613 = n11609 & n11612 ;
  assign n11614 = n11478 & ~n11613 ;
  assign n11615 = ~\pi0144  & n6706 ;
  assign n11616 = n6955 & n11615 ;
  assign n11617 = ~n6761 & n11616 ;
  assign n11618 = n6954 & n11617 ;
  assign n11619 = ~\pi0038  & ~n11618 ;
  assign n11620 = n11614 & n11619 ;
  assign n11621 = ~n11606 & ~n11620 ;
  assign n11622 = n11600 & n11621 ;
  assign n11623 = \pi0039  & ~n11581 ;
  assign n11624 = ~n11622 & n11623 ;
  assign n11625 = ~n11584 & ~n11624 ;
  assign n11626 = n2855 & ~n11480 ;
  assign n11627 = n1354 & n11626 ;
  assign n11628 = n8413 & n11627 ;
  assign n11629 = n1358 & n11628 ;
  assign n11630 = \pi0038  & ~n11467 ;
  assign n11631 = \pi0092  & ~n11630 ;
  assign n11632 = ~n11629 & n11631 ;
  assign n11633 = ~\pi0100  & \pi0232  ;
  assign n11634 = n6706 & n11633 ;
  assign n11635 = \pi0092  & ~n11634 ;
  assign n11636 = ~\pi0075  & ~n11635 ;
  assign n11637 = ~n11632 & n11636 ;
  assign n11638 = ~n11166 & ~n11637 ;
  assign n11639 = ~\pi0100  & ~n11638 ;
  assign n11640 = n11625 & n11639 ;
  assign n11641 = ~n11583 & n11640 ;
  assign n11642 = n2511 & n11464 ;
  assign n11643 = n2511 & ~n11166 ;
  assign n11644 = ~n11637 & n11643 ;
  assign n11645 = ~n11642 & ~n11644 ;
  assign n11646 = ~n11641 & ~n11645 ;
  assign n11647 = ~\pi0074  & n11494 ;
  assign n11648 = ~n11166 & n11647 ;
  assign n11649 = n11148 & ~n11648 ;
  assign n11650 = n11174 & n11649 ;
  assign n11651 = ~n11646 & n11650 ;
  assign n11652 = n10190 & ~n11131 ;
  assign n11653 = \pi0038  & n11140 ;
  assign n11654 = ~\pi0054  & ~n11653 ;
  assign n11655 = n11186 & ~n11654 ;
  assign n11656 = ~\pi0092  & \pi0162  ;
  assign n11657 = n2855 & n11656 ;
  assign n11658 = n6706 & n8364 ;
  assign n11659 = n11657 & n11658 ;
  assign n11660 = n1259 & n11659 ;
  assign n11661 = n1249 & n11660 ;
  assign n11662 = n1281 & n11186 ;
  assign n11663 = n11661 & n11662 ;
  assign n11664 = ~n11655 & ~n11663 ;
  assign n11665 = n11652 & n11664 ;
  assign n11666 = n11148 & n11179 ;
  assign n11667 = ~n11665 & n11666 ;
  assign n11668 = \pi0034  & n2467 ;
  assign n11669 = \pi0034  & n11138 ;
  assign n11670 = ~n11131 & n11669 ;
  assign n11671 = ~n11668 & ~n11670 ;
  assign n11672 = ~n11667 & ~n11671 ;
  assign n11673 = ~n11651 & n11672 ;
  assign n11674 = ~n11506 & ~n11673 ;
  assign n11675 = ~n11505 & n11674 ;
  assign n11676 = ~\pi0079  & ~\pi0118  ;
  assign n11677 = n11101 & n11676 ;
  assign n11678 = ~\pi0034  & ~n11677 ;
  assign n11679 = ~n11503 & ~n11678 ;
  assign n11680 = ~n11501 & n11679 ;
  assign n11681 = ~n11503 & n11678 ;
  assign n11682 = ~n11667 & n11681 ;
  assign n11683 = ~n11651 & n11682 ;
  assign n11684 = n11506 & ~n11683 ;
  assign n11685 = ~n11680 & n11684 ;
  assign n11686 = ~n11675 & ~n11685 ;
  assign n11687 = \pi0137  & n6807 ;
  assign n11688 = n6804 & n11687 ;
  assign n11689 = ~n6795 & n11688 ;
  assign n11690 = ~\pi0038  & n2851 ;
  assign n11691 = n10071 & n11690 ;
  assign n11692 = n1281 & n11691 ;
  assign n11693 = n1260 & n11692 ;
  assign n11694 = n11689 & n11693 ;
  assign n11695 = ~\pi0137  & \pi0252  ;
  assign n11696 = \pi0146  & \pi0299  ;
  assign n11697 = ~n1801 & n11696 ;
  assign n11698 = \pi0142  & ~\pi0299  ;
  assign n11699 = ~n2167 & n11698 ;
  assign n11700 = ~n11697 & ~n11699 ;
  assign n11701 = ~n8639 & n11700 ;
  assign n11702 = \pi0683  & \pi0824  ;
  assign n11703 = n6809 & n11702 ;
  assign n11704 = ~n6704 & n11703 ;
  assign n11705 = \pi0252  & ~n11704 ;
  assign n11706 = ~n6808 & n11705 ;
  assign n11707 = ~n11701 & ~n11706 ;
  assign n11708 = ~n8641 & ~n11707 ;
  assign n11709 = ~n11695 & ~n11708 ;
  assign n11710 = n6795 & ~n6808 ;
  assign n11711 = ~n8641 & ~n11706 ;
  assign n11712 = n11710 & n11711 ;
  assign n11713 = ~n11709 & ~n11712 ;
  assign n11714 = n10076 & n11690 ;
  assign n11715 = ~n11713 & n11714 ;
  assign n11716 = ~n11694 & ~n11715 ;
  assign n11717 = ~\pi0024  & n1281 ;
  assign n11718 = n1260 & n11717 ;
  assign n11719 = \pi0038  & ~n11718 ;
  assign n11720 = n2320 & ~n11719 ;
  assign n11721 = n11716 & ~n11720 ;
  assign n11722 = \pi1082  & n1264 ;
  assign n11723 = n1621 & n11722 ;
  assign n11724 = ~\pi0090  & n6637 ;
  assign n11725 = n1358 & n11724 ;
  assign n11726 = n7083 & ~n11725 ;
  assign n11727 = n1896 & ~n6642 ;
  assign n11728 = ~n11726 & ~n11727 ;
  assign n11729 = ~\pi0035  & n1364 ;
  assign n11730 = n1263 & n11729 ;
  assign n11731 = \pi0841  & n1364 ;
  assign n11732 = n1263 & n11731 ;
  assign n11733 = n1354 & n11732 ;
  assign n11734 = n1358 & n11733 ;
  assign n11735 = ~n11730 & ~n11734 ;
  assign n11736 = n11722 & ~n11735 ;
  assign n11737 = n11728 & n11736 ;
  assign n11738 = ~n11723 & ~n11737 ;
  assign n11739 = n1264 & ~n10048 ;
  assign n11740 = ~\pi0038  & ~n11739 ;
  assign n11741 = ~\pi0038  & ~n11730 ;
  assign n11742 = ~n11734 & n11741 ;
  assign n11743 = ~n11740 & ~n11742 ;
  assign n11744 = ~\pi0122  & ~n8604 ;
  assign n11745 = ~n6684 & n9250 ;
  assign n11746 = ~n11744 & n11745 ;
  assign n11747 = ~\pi0122  & \pi1091  ;
  assign n11748 = n1689 & n11747 ;
  assign n11749 = n1688 & n11748 ;
  assign n11750 = ~n6684 & ~n9250 ;
  assign n11751 = ~n11749 & n11750 ;
  assign n11752 = ~n11746 & ~n11751 ;
  assign n11753 = n11728 & n11752 ;
  assign n11754 = n10047 & n10058 ;
  assign n11755 = ~n9250 & ~n11749 ;
  assign n11756 = n9250 & ~n11744 ;
  assign n11757 = ~n11755 & ~n11756 ;
  assign n11758 = n11754 & n11757 ;
  assign n11759 = ~\pi0038  & ~n11758 ;
  assign n11760 = ~n11753 & n11759 ;
  assign n11761 = n11743 & ~n11760 ;
  assign n11762 = n11738 & ~n11761 ;
  assign n11763 = ~\pi0032  & ~n11735 ;
  assign n11764 = n11728 & n11763 ;
  assign n11765 = \pi0032  & n10018 ;
  assign n11766 = n1329 & n11765 ;
  assign n11767 = n1627 & n11766 ;
  assign n11768 = n1319 & n11767 ;
  assign n11769 = ~n11764 & ~n11768 ;
  assign n11770 = ~\pi0095  & ~n6684 ;
  assign n11771 = ~n11769 & n11770 ;
  assign n11772 = n11716 & ~n11771 ;
  assign n11773 = n11762 & n11772 ;
  assign n11774 = ~n11721 & ~n11773 ;
  assign n11775 = n1287 & n11774 ;
  assign n11776 = \pi0137  & ~n10050 ;
  assign n11777 = ~n1696 & n11776 ;
  assign n11778 = ~n10092 & n11777 ;
  assign n11779 = n10080 & ~n11778 ;
  assign n11780 = ~\pi0024  & n10094 ;
  assign n11781 = n10093 & n11780 ;
  assign n11782 = n1259 & n11781 ;
  assign n11783 = n1249 & n11782 ;
  assign n11784 = n1281 & n1285 ;
  assign n11785 = n11783 & n11784 ;
  assign n11786 = ~n11779 & n11785 ;
  assign n11787 = ~\pi0024  & \pi0054  ;
  assign n11788 = n1259 & n11787 ;
  assign n11789 = n1249 & n11788 ;
  assign n11790 = n8410 & n11789 ;
  assign n11791 = ~\pi0059  & ~n11790 ;
  assign n11792 = ~n11786 & n11791 ;
  assign n11793 = ~n11775 & n11792 ;
  assign n11794 = ~\pi0059  & ~n10015 ;
  assign n11795 = ~\pi0024  & n1293 ;
  assign n11796 = n1291 & n11795 ;
  assign n11797 = n1281 & n11796 ;
  assign n11798 = n1260 & n11797 ;
  assign n11799 = \pi0059  & ~n11798 ;
  assign n11800 = ~\pi0057  & ~n11799 ;
  assign n11801 = ~n11794 & n11800 ;
  assign n11802 = ~n11793 & n11801 ;
  assign n11803 = n1504 & n6988 ;
  assign n11804 = n1253 & n1256 ;
  assign n11805 = n11803 & n11804 ;
  assign n11806 = \pi0036  & ~\pi0103  ;
  assign n11807 = n1252 & n11806 ;
  assign n11808 = n1275 & n11807 ;
  assign n11809 = ~\pi0067  & ~\pi0071  ;
  assign n11810 = ~\pi0083  & n11809 ;
  assign n11811 = ~\pi0069  & n11810 ;
  assign n11812 = n11808 & n11811 ;
  assign n11813 = n11805 & n11812 ;
  assign n11814 = n1468 & n10468 ;
  assign n11815 = n11813 & n11814 ;
  assign n11816 = ~\pi0024  & ~\pi0058  ;
  assign n11817 = n1325 & n1398 ;
  assign n11818 = n11816 & n11817 ;
  assign n11819 = n1319 & n11818 ;
  assign n11820 = ~n11815 & ~n11819 ;
  assign n11821 = n1293 & n2467 ;
  assign n11822 = n1291 & n11821 ;
  assign n11823 = n1322 & n10903 ;
  assign n11824 = n11822 & n11823 ;
  assign n11825 = n8604 & n11824 ;
  assign n11826 = ~n11820 & n11825 ;
  assign n11827 = ~n8445 & ~n8448 ;
  assign n11828 = \pi0024  & ~\pi0039  ;
  assign n11829 = n1264 & n11828 ;
  assign n11830 = n1329 & n11829 ;
  assign n11831 = n1627 & n11830 ;
  assign n11832 = n1319 & n11831 ;
  assign n11833 = \pi0038  & ~n11832 ;
  assign n11834 = n6861 & n9948 ;
  assign n11835 = \pi0038  & n11834 ;
  assign n11836 = ~\pi0045  & ~\pi0073  ;
  assign n11837 = n10030 & n11836 ;
  assign n11838 = ~\pi0048  & ~\pi0065  ;
  assign n11839 = \pi0089  & n11838 ;
  assign n11840 = n11837 & n11839 ;
  assign n11841 = ~\pi0071  & ~\pi0104  ;
  assign n11842 = n1256 & n11841 ;
  assign n11843 = n1239 & n11842 ;
  assign n11844 = n11840 & n11843 ;
  assign n11845 = \pi0332  & n10311 ;
  assign n11846 = n10310 & n11845 ;
  assign n11847 = n11844 & n11846 ;
  assign n11848 = ~\pi0064  & ~n11847 ;
  assign n11849 = ~\pi0039  & ~\pi0841  ;
  assign n11850 = n1504 & n11849 ;
  assign n11851 = n1254 & n11850 ;
  assign n11852 = n1281 & n11851 ;
  assign n11853 = ~n11848 & n11852 ;
  assign n11854 = ~n1497 & n11834 ;
  assign n11855 = n11853 & n11854 ;
  assign n11856 = ~n11835 & ~n11855 ;
  assign n11857 = ~n11833 & ~n11856 ;
  assign n11858 = n2467 & n10015 ;
  assign n11859 = \pi0786  & ~\pi1082  ;
  assign n11860 = ~\pi0223  & ~\pi1093  ;
  assign n11861 = n11859 & n11860 ;
  assign n11862 = n6811 & n11861 ;
  assign n11863 = ~n8387 & n11862 ;
  assign n11864 = ~\pi1093  & n11859 ;
  assign n11865 = n6811 & n11864 ;
  assign n11866 = n2256 & n6706 ;
  assign n11867 = ~n6732 & n11866 ;
  assign n11868 = n2256 & ~n6706 ;
  assign n11869 = ~n6713 & n11868 ;
  assign n11870 = ~n11867 & ~n11869 ;
  assign n11871 = n11865 & ~n11870 ;
  assign n11872 = ~n11863 & ~n11871 ;
  assign n11873 = n6921 & ~n11872 ;
  assign n11874 = \pi0039  & n11873 ;
  assign n11875 = n6716 & n6718 ;
  assign n11876 = n1281 & n11875 ;
  assign n11877 = n1260 & n11876 ;
  assign n11878 = ~\pi0299  & ~n11877 ;
  assign n11879 = ~\pi0984  & ~n6809 ;
  assign n11880 = \pi0835  & ~n11879 ;
  assign n11881 = n6716 & ~n11880 ;
  assign n11882 = n6705 & ~n11881 ;
  assign n11883 = ~n6770 & n11882 ;
  assign n11884 = \pi1093  & ~n6716 ;
  assign n11885 = \pi0835  & \pi1093  ;
  assign n11886 = ~n11879 & n11885 ;
  assign n11887 = ~n11884 & ~n11886 ;
  assign n11888 = n6705 & ~n11887 ;
  assign n11889 = ~\pi0223  & ~n11888 ;
  assign n11890 = ~\pi0299  & ~n11889 ;
  assign n11891 = n11883 & n11890 ;
  assign n11892 = ~n11878 & ~n11891 ;
  assign n11893 = ~n11859 & n11892 ;
  assign n11894 = \pi0299  & ~n11877 ;
  assign n11895 = ~n6744 & n11882 ;
  assign n11896 = ~\pi0215  & ~n11888 ;
  assign n11897 = \pi0299  & ~n11896 ;
  assign n11898 = n11895 & n11897 ;
  assign n11899 = ~n11894 & ~n11898 ;
  assign n11900 = \pi0039  & n11899 ;
  assign n11901 = n11893 & n11900 ;
  assign n11902 = ~n11874 & ~n11901 ;
  assign n11903 = n2363 & n7265 ;
  assign n11904 = ~n11902 & n11903 ;
  assign n11905 = ~\pi0841  & n1618 ;
  assign n11906 = n1354 & n11905 ;
  assign n11907 = n1358 & n11906 ;
  assign n11908 = ~n2582 & ~n11907 ;
  assign n11909 = n1634 & ~n11908 ;
  assign n11910 = n10024 & n10909 ;
  assign n11911 = ~n11909 & ~n11910 ;
  assign n11912 = \pi0252  & ~\pi1093  ;
  assign n11913 = n6811 & n11912 ;
  assign n11914 = \pi0252  & \pi0986  ;
  assign n11915 = \pi0314  & ~n11914 ;
  assign n11916 = ~n11913 & n11915 ;
  assign n11917 = n1270 & n1326 ;
  assign n11918 = n1315 & n11917 ;
  assign n11919 = ~n11916 & n11918 ;
  assign n11920 = n1249 & n1388 ;
  assign n11921 = ~\pi0065  & ~\pi0069  ;
  assign n11922 = ~\pi0068  & ~\pi0082  ;
  assign n11923 = \pi0048  & n11922 ;
  assign n11924 = ~\pi0049  & n11836 ;
  assign n11925 = n11923 & n11924 ;
  assign n11926 = n11921 & n11925 ;
  assign n11927 = n10035 & n10043 ;
  assign n11928 = ~\pi0066  & ~\pi0084  ;
  assign n11929 = n1530 & n11928 ;
  assign n11930 = n10307 & n11929 ;
  assign n11931 = n11927 & n11930 ;
  assign n11932 = n11926 & n11931 ;
  assign n11933 = ~\pi0047  & ~\pi0841  ;
  assign n11934 = n11843 & n11933 ;
  assign n11935 = n11932 & n11934 ;
  assign n11936 = ~n11920 & ~n11935 ;
  assign n11937 = n11919 & ~n11936 ;
  assign n11938 = n1320 & n11937 ;
  assign n11939 = ~\pi0046  & n1270 ;
  assign n11940 = ~\pi0097  & ~\pi0841  ;
  assign n11941 = n1276 & n11940 ;
  assign n11942 = n11939 & n11941 ;
  assign n11943 = n11843 & n11942 ;
  assign n11944 = n11932 & n11943 ;
  assign n11945 = ~n1595 & n11944 ;
  assign n11946 = ~\pi0046  & \pi0108  ;
  assign n11947 = n1270 & n11946 ;
  assign n11948 = n1592 & n11947 ;
  assign n11949 = n1568 & n11948 ;
  assign n11950 = n1542 & n11949 ;
  assign n11951 = ~\pi0047  & ~n11950 ;
  assign n11952 = ~n11945 & n11951 ;
  assign n11953 = n1326 & n11916 ;
  assign n11954 = ~n1392 & n11953 ;
  assign n11955 = n1320 & n11954 ;
  assign n11956 = ~n11952 & n11955 ;
  assign n11957 = ~n11938 & ~n11956 ;
  assign n11958 = ~\pi0035  & ~n11910 ;
  assign n11959 = n11957 & n11958 ;
  assign n11960 = ~n11911 & ~n11959 ;
  assign n11961 = n4520 & n11903 ;
  assign n11962 = n11960 & n11961 ;
  assign n11963 = ~n11904 & ~n11962 ;
  assign n11964 = n11858 & ~n11963 ;
  assign n11965 = \pi0102  & n1276 ;
  assign n11966 = ~\pi0035  & n1252 ;
  assign n11967 = n1618 & n11966 ;
  assign n11968 = n11965 & n11967 ;
  assign n11969 = n1253 & n1278 ;
  assign n11970 = n1273 & n11969 ;
  assign n11971 = n11968 & n11970 ;
  assign n11972 = n1534 & n11971 ;
  assign n11973 = ~\pi0040  & ~n11972 ;
  assign n11974 = n1264 & ~n11973 ;
  assign n11975 = ~n2585 & n11974 ;
  assign n11976 = ~\pi1082  & ~n11975 ;
  assign n11977 = n1253 & n2575 ;
  assign n11978 = n11968 & n11977 ;
  assign n11979 = n1351 & n11978 ;
  assign n11980 = n1534 & n11979 ;
  assign n11981 = \pi1082  & ~n11980 ;
  assign n11982 = n11822 & ~n11981 ;
  assign n11983 = ~n11976 & n11982 ;
  assign n11984 = ~\pi0166  & n6706 ;
  assign n11985 = ~\pi0152  & \pi0161  ;
  assign n11986 = n11984 & n11985 ;
  assign n11987 = ~n8637 & ~n11986 ;
  assign n11988 = \pi0232  & ~n11987 ;
  assign n11989 = \pi0144  & ~\pi0189  ;
  assign n11990 = n6706 & n11989 ;
  assign n11991 = \pi0039  & ~\pi0174  ;
  assign n11992 = n11990 & n11991 ;
  assign n11993 = ~n2297 & ~n11992 ;
  assign n11994 = n11988 & ~n11993 ;
  assign n11995 = \pi0039  & \pi0072  ;
  assign n11996 = ~\pi0041  & ~\pi0072  ;
  assign n11997 = ~\pi0039  & ~n11996 ;
  assign n11998 = n9948 & ~n11997 ;
  assign n11999 = ~n11995 & n11998 ;
  assign n12000 = ~n11994 & n11999 ;
  assign n12001 = ~\pi0057  & ~\pi0074  ;
  assign n12002 = n1285 & n12001 ;
  assign n12003 = n6848 & n12002 ;
  assign n12004 = n11040 & n11985 ;
  assign n12005 = n11984 & n12004 ;
  assign n12006 = \pi0039  & ~\pi0072  ;
  assign n12007 = ~n11996 & ~n12006 ;
  assign n12008 = ~n9948 & ~n12007 ;
  assign n12009 = ~n12005 & n12008 ;
  assign n12010 = ~n12003 & ~n12009 ;
  assign n12011 = ~n12000 & n12010 ;
  assign n12012 = ~\pi0072  & \pi0101  ;
  assign n12013 = ~\pi0041  & ~n12012 ;
  assign n12014 = ~\pi0110  & n1682 ;
  assign n12015 = \pi0097  & n12014 ;
  assign n12016 = n8573 & n12014 ;
  assign n12017 = n1542 & n12016 ;
  assign n12018 = ~n12015 & ~n12017 ;
  assign n12019 = ~n1678 & ~n12018 ;
  assign n12020 = n8564 & ~n8729 ;
  assign n12021 = ~n12019 & n12020 ;
  assign n12022 = ~\pi0093  & ~n1277 ;
  assign n12023 = ~n8563 & n12022 ;
  assign n12024 = ~\pi0035  & ~\pi0070  ;
  assign n12025 = n1354 & n12024 ;
  assign n12026 = n1358 & n12025 ;
  assign n12027 = \pi0051  & ~n12026 ;
  assign n12028 = ~n8559 & ~n12027 ;
  assign n12029 = ~n12023 & n12028 ;
  assign n12030 = ~n12021 & n12029 ;
  assign n12031 = \pi0051  & n12026 ;
  assign n12032 = ~\pi0096  & ~n12031 ;
  assign n12033 = ~n12030 & n12032 ;
  assign n12034 = ~\pi0122  & n8743 ;
  assign n12035 = ~n12033 & n12034 ;
  assign n12036 = ~n8588 & n8592 ;
  assign n12037 = ~n8581 & n12036 ;
  assign n12038 = ~n8578 & n12037 ;
  assign n12039 = ~\pi0072  & ~n12038 ;
  assign n12040 = ~n12035 & n12039 ;
  assign n12041 = ~\pi0044  & \pi1093  ;
  assign n12042 = ~n12040 & n12041 ;
  assign n12043 = \pi0044  & \pi0072  ;
  assign n12044 = ~\pi0101  & ~n12043 ;
  assign n12045 = ~\pi0072  & n8588 ;
  assign n12046 = ~n8554 & n12045 ;
  assign n12047 = ~n8585 & n12046 ;
  assign n12048 = ~n8578 & n8593 ;
  assign n12049 = ~\pi0072  & ~n8588 ;
  assign n12050 = ~n12048 & n12049 ;
  assign n12051 = ~n12047 & ~n12050 ;
  assign n12052 = ~\pi0044  & ~\pi1093  ;
  assign n12053 = n12051 & n12052 ;
  assign n12054 = n12044 & ~n12053 ;
  assign n12055 = ~n12042 & n12054 ;
  assign n12056 = n12013 & ~n12055 ;
  assign n12057 = \pi1093  & ~n12038 ;
  assign n12058 = ~n12035 & n12057 ;
  assign n12059 = ~\pi0044  & n12037 ;
  assign n12060 = ~n8578 & n12059 ;
  assign n12061 = ~n12041 & ~n12060 ;
  assign n12062 = ~\pi0044  & n12045 ;
  assign n12063 = ~n8586 & n12062 ;
  assign n12064 = n12061 & ~n12063 ;
  assign n12065 = ~\pi0101  & ~n12064 ;
  assign n12066 = ~n12058 & n12065 ;
  assign n12067 = \pi0041  & ~n12066 ;
  assign n12068 = ~n12056 & ~n12067 ;
  assign n12069 = n8799 & n12068 ;
  assign n12070 = ~\pi0174  & n11990 ;
  assign n12071 = ~\pi0299  & ~n12070 ;
  assign n12072 = n11988 & ~n12071 ;
  assign n12073 = \pi0039  & \pi0287  ;
  assign n12074 = n1281 & n12073 ;
  assign n12075 = n1260 & n12074 ;
  assign n12076 = n12072 & n12075 ;
  assign n12077 = n12006 & ~n12072 ;
  assign n12078 = n2327 & ~n12077 ;
  assign n12079 = ~n12076 & n12078 ;
  assign n12080 = \pi1093  & ~n12048 ;
  assign n12081 = ~\pi0101  & ~n12080 ;
  assign n12082 = ~n12064 & n12081 ;
  assign n12083 = \pi0041  & ~n12082 ;
  assign n12084 = n12079 & n12083 ;
  assign n12085 = n12047 & ~n12048 ;
  assign n12086 = ~n12050 & ~n12080 ;
  assign n12087 = ~n12085 & n12086 ;
  assign n12088 = ~\pi0044  & n12087 ;
  assign n12089 = ~\pi0101  & ~n8799 ;
  assign n12090 = ~\pi0072  & n12089 ;
  assign n12091 = ~n12088 & n12090 ;
  assign n12092 = ~n8799 & ~n12013 ;
  assign n12093 = n12079 & ~n12092 ;
  assign n12094 = ~n12091 & n12093 ;
  assign n12095 = ~n12084 & ~n12094 ;
  assign n12096 = \pi0228  & ~n12095 ;
  assign n12097 = ~n12069 & n12096 ;
  assign n12098 = n12013 & ~n12044 ;
  assign n12099 = ~\pi0047  & ~\pi0109  ;
  assign n12100 = n1326 & n12099 ;
  assign n12101 = n1324 & n12100 ;
  assign n12102 = ~\pi0480  & \pi0949  ;
  assign n12103 = \pi0110  & n12102 ;
  assign n12104 = ~\pi0250  & \pi0252  ;
  assign n12105 = n12103 & ~n12104 ;
  assign n12106 = n2575 & n12105 ;
  assign n12107 = n12101 & n12106 ;
  assign n12108 = n1319 & n12107 ;
  assign n12109 = ~\pi0072  & ~n12108 ;
  assign n12110 = \pi0901  & ~\pi0959  ;
  assign n12111 = n1270 & n12110 ;
  assign n12112 = n1269 & n12111 ;
  assign n12113 = n1579 & n12112 ;
  assign n12114 = n1542 & n12113 ;
  assign n12115 = ~\pi0047  & ~\pi0250  ;
  assign n12116 = n1326 & n12115 ;
  assign n12117 = n7203 & n12116 ;
  assign n12118 = n1324 & n12117 ;
  assign n12119 = n12114 & n12118 ;
  assign n12120 = ~\pi0109  & \pi0110  ;
  assign n12121 = n12102 & n12120 ;
  assign n12122 = n12118 & n12121 ;
  assign n12123 = n1319 & n12122 ;
  assign n12124 = ~n12119 & ~n12123 ;
  assign n12125 = n12109 & n12124 ;
  assign n12126 = ~\pi0044  & n12013 ;
  assign n12127 = ~n12125 & n12126 ;
  assign n12128 = ~n12098 & ~n12127 ;
  assign n12129 = \pi0041  & ~n6806 ;
  assign n12130 = ~\pi0072  & n1323 ;
  assign n12131 = n1322 & n12130 ;
  assign n12132 = n12117 & n12131 ;
  assign n12133 = n12114 & n12132 ;
  assign n12134 = n12121 & n12132 ;
  assign n12135 = n1319 & n12134 ;
  assign n12136 = ~n12133 & ~n12135 ;
  assign n12137 = n8567 & n12120 ;
  assign n12138 = n1261 & n1320 ;
  assign n12139 = n12102 & ~n12104 ;
  assign n12140 = n12138 & n12139 ;
  assign n12141 = n1266 & n12140 ;
  assign n12142 = n12137 & n12141 ;
  assign n12143 = n1319 & n12142 ;
  assign n12144 = \pi0041  & ~n12143 ;
  assign n12145 = n12136 & n12144 ;
  assign n12146 = ~n12129 & ~n12145 ;
  assign n12147 = ~\pi0039  & n12146 ;
  assign n12148 = n12128 & n12147 ;
  assign n12149 = ~n9635 & ~n12148 ;
  assign n12150 = n12079 & n12149 ;
  assign n12151 = ~\pi0228  & ~n11996 ;
  assign n12152 = \pi0299  & ~n11996 ;
  assign n12153 = n1801 & n12152 ;
  assign n12154 = ~\pi0299  & ~n11996 ;
  assign n12155 = n2167 & n12154 ;
  assign n12156 = ~n12153 & ~n12155 ;
  assign n12157 = n8640 & ~n12156 ;
  assign n12158 = ~n12151 & ~n12157 ;
  assign n12159 = \pi0100  & ~n12158 ;
  assign n12160 = ~\pi0041  & \pi0072  ;
  assign n12161 = ~\pi0041  & ~\pi0044  ;
  assign n12162 = ~n12012 & n12161 ;
  assign n12163 = n2575 & n12162 ;
  assign n12164 = n1627 & n12163 ;
  assign n12165 = n1319 & n12164 ;
  assign n12166 = ~n12160 & ~n12165 ;
  assign n12167 = ~\pi0052  & ~\pi0099  ;
  assign n12168 = n6799 & n12167 ;
  assign n12169 = n6803 & n12168 ;
  assign n12170 = \pi1093  & n8588 ;
  assign n12171 = ~\pi0072  & ~n12170 ;
  assign n12172 = ~n12169 & ~n12171 ;
  assign n12173 = ~n12166 & n12172 ;
  assign n12174 = n8799 & ~n12160 ;
  assign n12175 = ~\pi0041  & n12174 ;
  assign n12176 = ~\pi0041  & n8799 ;
  assign n12177 = ~n12169 & n12176 ;
  assign n12178 = ~n12175 & ~n12177 ;
  assign n12179 = n1281 & n6806 ;
  assign n12180 = n1260 & n12179 ;
  assign n12181 = n8799 & ~n12169 ;
  assign n12182 = ~n12174 & ~n12181 ;
  assign n12183 = n12170 & ~n12182 ;
  assign n12184 = n12180 & n12183 ;
  assign n12185 = n12178 & ~n12184 ;
  assign n12186 = ~n12173 & ~n12185 ;
  assign n12187 = ~n8799 & n11996 ;
  assign n12188 = \pi0228  & ~n12187 ;
  assign n12189 = ~n8641 & n12188 ;
  assign n12190 = \pi0100  & n12189 ;
  assign n12191 = ~n12186 & n12190 ;
  assign n12192 = ~n12159 & ~n12191 ;
  assign n12193 = n1288 & ~n12192 ;
  assign n12194 = ~n11995 & ~n11997 ;
  assign n12195 = ~n11994 & n12194 ;
  assign n12196 = \pi0038  & ~n12195 ;
  assign n12197 = ~\pi0087  & ~n12196 ;
  assign n12198 = ~n12193 & n12197 ;
  assign n12199 = ~n2363 & ~n11995 ;
  assign n12200 = ~n11997 & n12199 ;
  assign n12201 = ~n11994 & n12200 ;
  assign n12202 = \pi0075  & ~n12201 ;
  assign n12203 = n8588 & n8798 ;
  assign n12204 = n6806 & n12203 ;
  assign n12205 = n1281 & n12204 ;
  assign n12206 = n1260 & n12205 ;
  assign n12207 = n7207 & n12206 ;
  assign n12208 = \pi0041  & ~n12207 ;
  assign n12209 = n7203 & n12203 ;
  assign n12210 = n1627 & n12209 ;
  assign n12211 = n1319 & n12210 ;
  assign n12212 = n12162 & ~n12169 ;
  assign n12213 = n12211 & n12212 ;
  assign n12214 = n12174 & ~n12213 ;
  assign n12215 = ~n12208 & n12214 ;
  assign n12216 = n9635 & ~n12187 ;
  assign n12217 = ~n8641 & n12216 ;
  assign n12218 = ~n12215 & n12217 ;
  assign n12219 = ~\pi0039  & n12151 ;
  assign n12220 = ~\pi0039  & n8640 ;
  assign n12221 = ~n12156 & n12220 ;
  assign n12222 = ~n12219 & ~n12221 ;
  assign n12223 = n2363 & ~n11995 ;
  assign n12224 = ~n11994 & n12223 ;
  assign n12225 = n12222 & n12224 ;
  assign n12226 = ~n12218 & n12225 ;
  assign n12227 = n12202 & ~n12226 ;
  assign n12228 = n6785 & n11995 ;
  assign n12229 = n6785 & ~n11993 ;
  assign n12230 = n11988 & n12229 ;
  assign n12231 = ~n12228 & ~n12230 ;
  assign n12232 = ~n12227 & n12231 ;
  assign n12233 = n12198 & n12232 ;
  assign n12234 = ~n12150 & n12233 ;
  assign n12235 = ~n12097 & n12234 ;
  assign n12236 = \pi0041  & ~n12180 ;
  assign n12237 = \pi0228  & ~n12160 ;
  assign n12238 = ~n12165 & n12237 ;
  assign n12239 = ~n12236 & n12238 ;
  assign n12240 = ~\pi0228  & n11996 ;
  assign n12241 = ~\pi0075  & ~n12240 ;
  assign n12242 = n2328 & n12241 ;
  assign n12243 = ~n12239 & n12242 ;
  assign n12244 = ~n2327 & n11997 ;
  assign n12245 = \pi0087  & ~n12244 ;
  assign n12246 = ~n11995 & n12245 ;
  assign n12247 = ~n11994 & n12246 ;
  assign n12248 = ~\pi0075  & ~n12247 ;
  assign n12249 = ~n12243 & ~n12248 ;
  assign n12250 = ~n12227 & n12249 ;
  assign n12251 = n8496 & ~n12009 ;
  assign n12252 = ~n12250 & n12251 ;
  assign n12253 = ~n12235 & n12252 ;
  assign n12254 = ~n12011 & ~n12253 ;
  assign n12255 = \pi0212  & \pi0214  ;
  assign n12256 = \pi0211  & n12255 ;
  assign n12257 = ~\pi0219  & ~n12256 ;
  assign n12258 = \pi0042  & ~\pi0072  ;
  assign n12259 = \pi0042  & ~\pi0114  ;
  assign n12260 = ~n12258 & ~n12259 ;
  assign n12261 = ~\pi0072  & \pi0113  ;
  assign n12262 = ~\pi0072  & \pi0116  ;
  assign n12263 = ~n12261 & ~n12262 ;
  assign n12264 = \pi0072  & ~n6805 ;
  assign n12265 = n6799 & ~n12264 ;
  assign n12266 = n12263 & ~n12265 ;
  assign n12267 = n6805 & ~n12012 ;
  assign n12268 = n12263 & n12267 ;
  assign n12269 = ~\pi0072  & ~\pi0101  ;
  assign n12270 = ~n12088 & n12269 ;
  assign n12271 = n12268 & ~n12270 ;
  assign n12272 = ~n12266 & ~n12271 ;
  assign n12273 = ~n12260 & n12272 ;
  assign n12274 = \pi0114  & ~n12258 ;
  assign n12275 = ~\pi0101  & n6805 ;
  assign n12276 = ~\pi1093  & n12275 ;
  assign n12277 = n8593 & n12275 ;
  assign n12278 = ~n8578 & n12277 ;
  assign n12279 = ~n12276 & ~n12278 ;
  assign n12280 = ~\pi0042  & n6799 ;
  assign n12281 = ~n12279 & n12280 ;
  assign n12282 = ~n12064 & n12281 ;
  assign n12283 = ~\pi0114  & ~n12282 ;
  assign n12284 = ~n12274 & ~n12283 ;
  assign n12285 = ~\pi0115  & ~n8799 ;
  assign n12286 = ~n12284 & n12285 ;
  assign n12287 = ~n12273 & n12286 ;
  assign n12288 = ~n12055 & n12268 ;
  assign n12289 = ~n12266 & ~n12288 ;
  assign n12290 = ~\pi0115  & \pi1091  ;
  assign n12291 = ~n1686 & n12290 ;
  assign n12292 = n12259 & n12291 ;
  assign n12293 = ~n12289 & n12292 ;
  assign n12294 = \pi0115  & ~n12258 ;
  assign n12295 = \pi0228  & ~n12294 ;
  assign n12296 = n6799 & ~n12274 ;
  assign n12297 = n6805 & n12296 ;
  assign n12298 = ~n12058 & n12297 ;
  assign n12299 = n12065 & n12298 ;
  assign n12300 = n12260 & n12291 ;
  assign n12301 = ~n12299 & n12300 ;
  assign n12302 = n12295 & ~n12301 ;
  assign n12303 = ~n12293 & n12302 ;
  assign n12304 = ~n12287 & n12303 ;
  assign n12305 = ~n12044 & n12267 ;
  assign n12306 = ~\pi0044  & n12267 ;
  assign n12307 = ~n12125 & n12306 ;
  assign n12308 = ~n12305 & ~n12307 ;
  assign n12309 = n12265 & n12308 ;
  assign n12310 = ~\pi0115  & n12259 ;
  assign n12311 = n12263 & n12310 ;
  assign n12312 = ~n12309 & n12311 ;
  assign n12313 = n12136 & ~n12143 ;
  assign n12314 = n6807 & n12296 ;
  assign n12315 = ~n12313 & n12314 ;
  assign n12316 = ~\pi0115  & n12260 ;
  assign n12317 = ~n12315 & n12316 ;
  assign n12318 = ~\pi0228  & ~n12294 ;
  assign n12319 = ~n12317 & n12318 ;
  assign n12320 = ~n12312 & n12319 ;
  assign n12321 = n2328 & ~n12320 ;
  assign n12322 = ~n12304 & n12321 ;
  assign n12323 = ~\pi0072  & \pi0199  ;
  assign n12324 = ~\pi0232  & ~n12323 ;
  assign n12325 = ~\pi0299  & ~n12324 ;
  assign n12326 = ~\pi0072  & \pi0200  ;
  assign n12327 = ~\pi0232  & ~n12326 ;
  assign n12328 = ~\pi0299  & ~n12327 ;
  assign n12329 = ~n12325 & ~n12328 ;
  assign n12330 = ~\pi0189  & n6706 ;
  assign n12331 = ~\pi0072  & ~n12330 ;
  assign n12332 = \pi0287  & n12330 ;
  assign n12333 = n1281 & n12332 ;
  assign n12334 = n1260 & n12333 ;
  assign n12335 = ~n12331 & ~n12334 ;
  assign n12336 = \pi0200  & ~n12335 ;
  assign n12337 = ~\pi0199  & \pi0232  ;
  assign n12338 = \pi0232  & ~n12331 ;
  assign n12339 = ~n12334 & n12338 ;
  assign n12340 = ~n12337 & ~n12339 ;
  assign n12341 = ~n12336 & ~n12340 ;
  assign n12342 = ~n12329 & ~n12341 ;
  assign n12343 = \pi0039  & n2327 ;
  assign n12344 = ~n12342 & n12343 ;
  assign n12345 = ~\pi0228  & ~n12258 ;
  assign n12346 = \pi0299  & ~n12258 ;
  assign n12347 = n1801 & n12346 ;
  assign n12348 = ~\pi0299  & ~n12258 ;
  assign n12349 = n2167 & n12348 ;
  assign n12350 = ~n12347 & ~n12349 ;
  assign n12351 = n8640 & ~n12350 ;
  assign n12352 = ~n12345 & ~n12351 ;
  assign n12353 = n12258 & ~n12291 ;
  assign n12354 = \pi0228  & ~n12353 ;
  assign n12355 = ~n8641 & n12354 ;
  assign n12356 = n12352 & ~n12355 ;
  assign n12357 = ~\pi0044  & ~\pi0095  ;
  assign n12358 = n1634 & n12357 ;
  assign n12359 = n12170 & n12358 ;
  assign n12360 = n1627 & n12359 ;
  assign n12361 = n1319 & n12360 ;
  assign n12362 = n6799 & n12275 ;
  assign n12363 = n12361 & n12362 ;
  assign n12364 = n12258 & ~n12363 ;
  assign n12365 = n6799 & n6806 ;
  assign n12366 = n1281 & n12365 ;
  assign n12367 = n1260 & n12366 ;
  assign n12368 = \pi1093  & n6805 ;
  assign n12369 = n8588 & n12368 ;
  assign n12370 = ~\pi0042  & ~\pi0043  ;
  assign n12371 = ~\pi0052  & n12370 ;
  assign n12372 = n6801 & ~n12371 ;
  assign n12373 = n12369 & n12372 ;
  assign n12374 = n12367 & n12373 ;
  assign n12375 = ~\pi0114  & ~n12374 ;
  assign n12376 = ~n12364 & n12375 ;
  assign n12377 = ~n12274 & n12291 ;
  assign n12378 = n12352 & n12377 ;
  assign n12379 = ~n12376 & n12378 ;
  assign n12380 = ~n12356 & ~n12379 ;
  assign n12381 = ~\pi0039  & n6785 ;
  assign n12382 = n12380 & n12381 ;
  assign n12383 = \pi0039  & ~\pi0232  ;
  assign n12384 = ~n12326 & n12383 ;
  assign n12385 = ~n2297 & ~n12384 ;
  assign n12386 = n12326 & ~n12330 ;
  assign n12387 = n11040 & ~n12386 ;
  assign n12388 = n12385 & ~n12387 ;
  assign n12389 = \pi0232  & ~n12323 ;
  assign n12390 = ~\pi0189  & \pi0232  ;
  assign n12391 = n6706 & n12390 ;
  assign n12392 = ~n12389 & ~n12391 ;
  assign n12393 = n12325 & n12392 ;
  assign n12394 = n6785 & ~n12393 ;
  assign n12395 = ~n12388 & n12394 ;
  assign n12396 = ~\pi0039  & ~n12258 ;
  assign n12397 = n1286 & ~n12396 ;
  assign n12398 = n12393 & n12397 ;
  assign n12399 = n12385 & n12397 ;
  assign n12400 = ~n12387 & n12399 ;
  assign n12401 = ~n12398 & ~n12400 ;
  assign n12402 = ~\pi0038  & n1286 ;
  assign n12403 = n12401 & ~n12402 ;
  assign n12404 = n8496 & ~n12403 ;
  assign n12405 = ~n12395 & n12404 ;
  assign n12406 = ~n12382 & n12405 ;
  assign n12407 = ~n12344 & n12406 ;
  assign n12408 = ~n12322 & n12407 ;
  assign n12409 = \pi0207  & \pi0208  ;
  assign n12410 = ~n8496 & ~n12396 ;
  assign n12411 = n12393 & n12410 ;
  assign n12412 = n12385 & n12410 ;
  assign n12413 = ~n12387 & n12412 ;
  assign n12414 = ~n12411 & ~n12413 ;
  assign n12415 = n12409 & n12414 ;
  assign n12416 = ~n12388 & ~n12393 ;
  assign n12417 = ~\pi0101  & \pi0228  ;
  assign n12418 = n6805 & n12417 ;
  assign n12419 = n12358 & n12418 ;
  assign n12420 = n1627 & n12419 ;
  assign n12421 = n1319 & n12420 ;
  assign n12422 = ~\pi0115  & n6799 ;
  assign n12423 = ~\pi0114  & n12422 ;
  assign n12424 = n12421 & n12423 ;
  assign n12425 = ~n2327 & n12396 ;
  assign n12426 = \pi0087  & ~n12425 ;
  assign n12427 = n12258 & n12426 ;
  assign n12428 = ~n12424 & n12427 ;
  assign n12429 = ~\pi0075  & ~n12426 ;
  assign n12430 = ~\pi0044  & n12418 ;
  assign n12431 = ~\pi0115  & n6801 ;
  assign n12432 = n6799 & n12431 ;
  assign n12433 = n12430 & n12432 ;
  assign n12434 = n1281 & n12433 ;
  assign n12435 = n1260 & n12434 ;
  assign n12436 = ~\pi0075  & n2328 ;
  assign n12437 = ~n12435 & n12436 ;
  assign n12438 = ~n12429 & ~n12437 ;
  assign n12439 = ~n12428 & ~n12438 ;
  assign n12440 = ~n12416 & ~n12439 ;
  assign n12441 = ~n2363 & n12258 ;
  assign n12442 = ~\pi0039  & \pi0075  ;
  assign n12443 = ~n12441 & n12442 ;
  assign n12444 = n8496 & ~n12443 ;
  assign n12445 = n12355 & ~n12377 ;
  assign n12446 = ~\pi0044  & ~\pi0113  ;
  assign n12447 = ~\pi0116  & n12446 ;
  assign n12448 = n12275 & n12447 ;
  assign n12449 = n12211 & n12448 ;
  assign n12450 = n12258 & ~n12449 ;
  assign n12451 = ~\pi0024  & n7207 ;
  assign n12452 = n12374 & n12451 ;
  assign n12453 = ~n12450 & ~n12452 ;
  assign n12454 = ~\pi0114  & n12355 ;
  assign n12455 = n12453 & n12454 ;
  assign n12456 = ~n12445 & ~n12455 ;
  assign n12457 = n2363 & ~n12345 ;
  assign n12458 = ~n12351 & n12457 ;
  assign n12459 = n8496 & n12458 ;
  assign n12460 = n12456 & n12459 ;
  assign n12461 = ~n12444 & ~n12460 ;
  assign n12462 = n12440 & ~n12461 ;
  assign n12463 = n12415 & ~n12462 ;
  assign n12464 = ~n12408 & n12463 ;
  assign n12465 = n12325 & n12340 ;
  assign n12466 = n12343 & ~n12465 ;
  assign n12467 = \pi0039  & n6785 ;
  assign n12468 = ~n12393 & n12467 ;
  assign n12469 = ~n12397 & ~n12402 ;
  assign n12470 = \pi0039  & ~n12402 ;
  assign n12471 = ~n12393 & n12470 ;
  assign n12472 = ~n12469 & ~n12471 ;
  assign n12473 = n8496 & n12472 ;
  assign n12474 = ~n12468 & n12473 ;
  assign n12475 = ~n12382 & n12474 ;
  assign n12476 = ~n12466 & n12475 ;
  assign n12477 = ~n12322 & n12476 ;
  assign n12478 = \pi0039  & ~n12393 ;
  assign n12479 = ~n12439 & ~n12478 ;
  assign n12480 = ~n12461 & n12479 ;
  assign n12481 = ~n12409 & ~n12410 ;
  assign n12482 = \pi0039  & ~n12409 ;
  assign n12483 = ~n12393 & n12482 ;
  assign n12484 = ~n12481 & ~n12483 ;
  assign n12485 = ~n12480 & ~n12484 ;
  assign n12486 = ~n12477 & n12485 ;
  assign n12487 = ~n12464 & ~n12486 ;
  assign n12488 = n12257 & ~n12487 ;
  assign n12489 = \pi0199  & ~n12335 ;
  assign n12490 = ~\pi0200  & n10118 ;
  assign n12491 = n10118 & ~n12331 ;
  assign n12492 = ~n12334 & n12491 ;
  assign n12493 = ~n12490 & ~n12492 ;
  assign n12494 = ~n12489 & ~n12493 ;
  assign n12495 = \pi0287  & n11984 ;
  assign n12496 = n1281 & n12495 ;
  assign n12497 = n1260 & n12496 ;
  assign n12498 = ~\pi0166  & \pi0232  ;
  assign n12499 = n6706 & n12498 ;
  assign n12500 = ~\pi0072  & ~n12499 ;
  assign n12501 = n10276 & ~n12500 ;
  assign n12502 = ~n12497 & n12501 ;
  assign n12503 = \pi0072  & ~\pi0232  ;
  assign n12504 = \pi0299  & ~n12503 ;
  assign n12505 = n12324 & ~n12504 ;
  assign n12506 = ~n12326 & n12505 ;
  assign n12507 = ~n12502 & ~n12506 ;
  assign n12508 = ~n12494 & n12507 ;
  assign n12509 = n12343 & ~n12508 ;
  assign n12510 = n12393 & ~n12396 ;
  assign n12511 = ~\pi0039  & n12258 ;
  assign n12512 = ~\pi0072  & \pi0299  ;
  assign n12513 = \pi0039  & n12512 ;
  assign n12514 = ~n12499 & n12513 ;
  assign n12515 = ~n12511 & ~n12514 ;
  assign n12516 = \pi0038  & n12515 ;
  assign n12517 = ~n12510 & n12516 ;
  assign n12518 = n12385 & ~n12396 ;
  assign n12519 = ~n12387 & n12518 ;
  assign n12520 = ~n12510 & ~n12519 ;
  assign n12521 = n12517 & n12520 ;
  assign n12522 = n1286 & ~n12521 ;
  assign n12523 = ~n12499 & n12512 ;
  assign n12524 = \pi0039  & ~n12523 ;
  assign n12525 = \pi0232  & ~n12326 ;
  assign n12526 = ~n12391 & ~n12525 ;
  assign n12527 = n12328 & n12526 ;
  assign n12528 = n12524 & ~n12527 ;
  assign n12529 = n12468 & n12528 ;
  assign n12530 = n8496 & ~n12529 ;
  assign n12531 = n12522 & n12530 ;
  assign n12532 = ~n12382 & n12531 ;
  assign n12533 = ~n12509 & n12532 ;
  assign n12534 = ~n12322 & n12533 ;
  assign n12535 = n12478 & n12528 ;
  assign n12536 = ~n12439 & ~n12535 ;
  assign n12537 = ~n12461 & n12536 ;
  assign n12538 = ~n8496 & ~n12515 ;
  assign n12539 = ~n12411 & ~n12538 ;
  assign n12540 = ~n12257 & n12539 ;
  assign n12541 = n12415 & n12540 ;
  assign n12542 = ~n12537 & n12541 ;
  assign n12543 = ~n12534 & n12542 ;
  assign n12544 = ~\pi0199  & n10118 ;
  assign n12545 = ~n12492 & ~n12544 ;
  assign n12546 = ~n12502 & ~n12505 ;
  assign n12547 = n12545 & n12546 ;
  assign n12548 = n12343 & ~n12547 ;
  assign n12549 = ~n8496 & ~n12409 ;
  assign n12550 = n12467 & ~n12523 ;
  assign n12551 = ~n12393 & n12550 ;
  assign n12552 = n1286 & ~n12551 ;
  assign n12553 = ~n12517 & n12552 ;
  assign n12554 = ~n12382 & n12553 ;
  assign n12555 = ~n12549 & n12554 ;
  assign n12556 = ~n12548 & n12555 ;
  assign n12557 = ~n12322 & n12556 ;
  assign n12558 = ~n12393 & n12524 ;
  assign n12559 = ~n12439 & ~n12558 ;
  assign n12560 = ~n12443 & n12559 ;
  assign n12561 = n12458 & n12559 ;
  assign n12562 = n12456 & n12561 ;
  assign n12563 = ~n12560 & ~n12562 ;
  assign n12564 = n8496 & ~n12563 ;
  assign n12565 = ~n12409 & ~n12564 ;
  assign n12566 = n12540 & n12565 ;
  assign n12567 = ~n12557 & n12566 ;
  assign n12568 = n9948 & ~n12567 ;
  assign n12569 = ~n12543 & n12568 ;
  assign n12570 = ~n12488 & n12569 ;
  assign n12571 = ~n12257 & n12500 ;
  assign n12572 = \pi0039  & ~n12571 ;
  assign n12573 = ~n9948 & ~n12396 ;
  assign n12574 = ~n12572 & n12573 ;
  assign n12575 = ~n12570 & ~n12574 ;
  assign n12576 = \pi0211  & ~n12255 ;
  assign n12577 = ~\pi0211  & ~\pi0219  ;
  assign n12578 = n12255 & n12577 ;
  assign n12579 = ~n12576 & ~n12578 ;
  assign n12580 = \pi0228  & ~n8799 ;
  assign n12581 = ~n12272 & n12580 ;
  assign n12582 = \pi0228  & \pi1091  ;
  assign n12583 = ~n1686 & n12582 ;
  assign n12584 = ~n12289 & n12583 ;
  assign n12585 = ~n12581 & ~n12584 ;
  assign n12586 = n6805 & ~n12058 ;
  assign n12587 = n12065 & n12586 ;
  assign n12588 = n12583 & ~n12587 ;
  assign n12589 = ~n8799 & n12279 ;
  assign n12590 = ~n8799 & n12061 ;
  assign n12591 = ~n12063 & n12590 ;
  assign n12592 = ~n12589 & ~n12591 ;
  assign n12593 = \pi0228  & ~n12592 ;
  assign n12594 = n6807 & ~n12313 ;
  assign n12595 = ~\pi0228  & ~n12594 ;
  assign n12596 = n12432 & ~n12595 ;
  assign n12597 = ~n12593 & n12596 ;
  assign n12598 = ~n12588 & n12597 ;
  assign n12599 = \pi0043  & ~\pi0072  ;
  assign n12600 = \pi0043  & ~\pi0115  ;
  assign n12601 = n6801 & n12600 ;
  assign n12602 = ~n12599 & ~n12601 ;
  assign n12603 = ~n12598 & n12602 ;
  assign n12604 = ~\pi0228  & n12263 ;
  assign n12605 = ~n12309 & n12604 ;
  assign n12606 = ~n12603 & ~n12605 ;
  assign n12607 = n12585 & n12606 ;
  assign n12608 = ~n12601 & ~n12603 ;
  assign n12609 = n2328 & ~n12608 ;
  assign n12610 = ~n12607 & n12609 ;
  assign n12611 = ~\pi0200  & \pi0232  ;
  assign n12612 = ~n12339 & ~n12611 ;
  assign n12613 = n12328 & n12612 ;
  assign n12614 = n12343 & ~n12613 ;
  assign n12615 = n8799 & n12431 ;
  assign n12616 = ~\pi0043  & \pi0052  ;
  assign n12617 = n12615 & n12616 ;
  assign n12618 = n12369 & n12617 ;
  assign n12619 = n12367 & n12618 ;
  assign n12620 = n12451 & n12619 ;
  assign n12621 = n12599 & n12615 ;
  assign n12622 = ~n12449 & n12621 ;
  assign n12623 = ~n12620 & ~n12622 ;
  assign n12624 = n12599 & ~n12615 ;
  assign n12625 = ~\pi0039  & ~n12599 ;
  assign n12626 = ~n6901 & ~n12625 ;
  assign n12627 = \pi0228  & ~n12626 ;
  assign n12628 = ~n12624 & n12627 ;
  assign n12629 = ~n8641 & n12628 ;
  assign n12630 = n12623 & n12629 ;
  assign n12631 = \pi0299  & ~n12599 ;
  assign n12632 = n1801 & n12631 ;
  assign n12633 = ~\pi0299  & ~n12599 ;
  assign n12634 = n2167 & n12633 ;
  assign n12635 = ~n12632 & ~n12634 ;
  assign n12636 = n8640 & ~n12635 ;
  assign n12637 = ~\pi0228  & ~n12599 ;
  assign n12638 = n2363 & ~n12637 ;
  assign n12639 = ~n12636 & n12638 ;
  assign n12640 = ~n12626 & ~n12639 ;
  assign n12641 = n12388 & ~n12640 ;
  assign n12642 = ~n12630 & n12641 ;
  assign n12643 = \pi0075  & ~n12642 ;
  assign n12644 = n8496 & ~n12643 ;
  assign n12645 = \pi0228  & ~n12624 ;
  assign n12646 = ~n8641 & n12645 ;
  assign n12647 = n12369 & n12616 ;
  assign n12648 = n12367 & n12647 ;
  assign n12649 = n12615 & n12648 ;
  assign n12650 = ~n12363 & n12621 ;
  assign n12651 = ~n12649 & ~n12650 ;
  assign n12652 = n12646 & n12651 ;
  assign n12653 = ~n12636 & ~n12637 ;
  assign n12654 = n12388 & n12653 ;
  assign n12655 = ~n12652 & n12654 ;
  assign n12656 = \pi0039  & n12328 ;
  assign n12657 = ~n12387 & n12656 ;
  assign n12658 = n6785 & ~n12657 ;
  assign n12659 = ~n12655 & n12658 ;
  assign n12660 = ~\pi0087  & ~n12625 ;
  assign n12661 = n12385 & n12660 ;
  assign n12662 = ~n12387 & n12661 ;
  assign n12663 = ~n2855 & ~n12662 ;
  assign n12664 = ~n12659 & ~n12663 ;
  assign n12665 = n12644 & n12664 ;
  assign n12666 = ~n12614 & n12665 ;
  assign n12667 = ~n12610 & n12666 ;
  assign n12668 = n6799 & n6803 ;
  assign n12669 = n12430 & n12668 ;
  assign n12670 = n1281 & n12669 ;
  assign n12671 = n1260 & n12670 ;
  assign n12672 = n2328 & ~n12671 ;
  assign n12673 = ~n2327 & n12625 ;
  assign n12674 = \pi0087  & ~n12673 ;
  assign n12675 = ~n12672 & n12674 ;
  assign n12676 = n12421 & n12432 ;
  assign n12677 = n12599 & n12674 ;
  assign n12678 = ~n12676 & n12677 ;
  assign n12679 = ~n12675 & ~n12678 ;
  assign n12680 = n12388 & ~n12679 ;
  assign n12681 = ~\pi0075  & ~n12680 ;
  assign n12682 = n8496 & ~n12681 ;
  assign n12683 = ~n12643 & n12682 ;
  assign n12684 = ~n8496 & ~n12625 ;
  assign n12685 = n12385 & n12684 ;
  assign n12686 = ~n12387 & n12685 ;
  assign n12687 = ~n12409 & ~n12686 ;
  assign n12688 = ~n12683 & n12687 ;
  assign n12689 = ~n12667 & n12688 ;
  assign n12690 = n12579 & n12689 ;
  assign n12691 = ~\pi0199  & ~\pi0200  ;
  assign n12692 = ~\pi0072  & ~\pi0299  ;
  assign n12693 = n12691 & n12692 ;
  assign n12694 = ~n10118 & ~n12693 ;
  assign n12695 = \pi0232  & ~n12691 ;
  assign n12696 = ~n12339 & ~n12695 ;
  assign n12697 = ~n12694 & n12696 ;
  assign n12698 = n12343 & ~n12697 ;
  assign n12699 = ~\pi0072  & n12691 ;
  assign n12700 = ~n12330 & n12699 ;
  assign n12701 = n11040 & ~n12700 ;
  assign n12702 = \pi0039  & ~n10118 ;
  assign n12703 = ~n12693 & n12702 ;
  assign n12704 = ~n12637 & ~n12703 ;
  assign n12705 = ~n12701 & n12704 ;
  assign n12706 = ~n12636 & n12705 ;
  assign n12707 = \pi0039  & ~n12694 ;
  assign n12708 = ~n12701 & n12707 ;
  assign n12709 = n6785 & ~n12708 ;
  assign n12710 = ~n12706 & n12709 ;
  assign n12711 = n12646 & n12709 ;
  assign n12712 = n12651 & n12711 ;
  assign n12713 = ~n12710 & ~n12712 ;
  assign n12714 = n12660 & ~n12703 ;
  assign n12715 = ~n12701 & n12714 ;
  assign n12716 = ~n2855 & ~n12715 ;
  assign n12717 = ~\pi0075  & ~n12716 ;
  assign n12718 = n12713 & n12717 ;
  assign n12719 = ~n12698 & n12718 ;
  assign n12720 = ~n12610 & n12719 ;
  assign n12721 = ~n12625 & ~n12703 ;
  assign n12722 = ~n12701 & n12721 ;
  assign n12723 = ~n2402 & ~n12722 ;
  assign n12724 = ~\pi0075  & ~n12723 ;
  assign n12725 = ~n12679 & n12724 ;
  assign n12726 = \pi0075  & ~n12703 ;
  assign n12727 = ~n12701 & n12726 ;
  assign n12728 = ~n12640 & n12727 ;
  assign n12729 = ~n12630 & n12728 ;
  assign n12730 = ~n12725 & ~n12729 ;
  assign n12731 = ~n12720 & n12730 ;
  assign n12732 = n8496 & ~n12731 ;
  assign n12733 = n12684 & ~n12703 ;
  assign n12734 = ~n12701 & n12733 ;
  assign n12735 = n12409 & ~n12734 ;
  assign n12736 = n12579 & n12735 ;
  assign n12737 = ~n12732 & n12736 ;
  assign n12738 = ~n12690 & ~n12737 ;
  assign n12739 = n12327 & ~n12504 ;
  assign n12740 = ~n12502 & ~n12739 ;
  assign n12741 = n12493 & n12740 ;
  assign n12742 = n12343 & ~n12741 ;
  assign n12743 = ~n12528 & ~n12640 ;
  assign n12744 = ~n12630 & n12743 ;
  assign n12745 = \pi0075  & ~n12744 ;
  assign n12746 = n8496 & ~n12745 ;
  assign n12747 = ~n12528 & n12653 ;
  assign n12748 = n6785 & ~n12523 ;
  assign n12749 = ~n12527 & n12748 ;
  assign n12750 = ~n12381 & ~n12749 ;
  assign n12751 = ~n12747 & ~n12750 ;
  assign n12752 = n12646 & ~n12750 ;
  assign n12753 = n12651 & n12752 ;
  assign n12754 = ~n12751 & ~n12753 ;
  assign n12755 = n12526 & ~n12625 ;
  assign n12756 = n12328 & n12755 ;
  assign n12757 = ~\pi0039  & n12599 ;
  assign n12758 = ~n12514 & ~n12757 ;
  assign n12759 = \pi0038  & n12758 ;
  assign n12760 = ~n12756 & n12759 ;
  assign n12761 = ~\pi0087  & ~n12760 ;
  assign n12762 = n12754 & n12761 ;
  assign n12763 = n12746 & n12762 ;
  assign n12764 = ~n12742 & n12763 ;
  assign n12765 = ~n12610 & n12764 ;
  assign n12766 = ~n12528 & ~n12679 ;
  assign n12767 = ~\pi0075  & ~n12766 ;
  assign n12768 = n8496 & ~n12767 ;
  assign n12769 = ~n12745 & n12768 ;
  assign n12770 = ~n8496 & ~n12758 ;
  assign n12771 = ~n8496 & n12328 ;
  assign n12772 = n12755 & n12771 ;
  assign n12773 = ~n12770 & ~n12772 ;
  assign n12774 = ~n12409 & n12773 ;
  assign n12775 = ~n12769 & n12774 ;
  assign n12776 = ~n12765 & n12775 ;
  assign n12777 = n10118 & ~n12691 ;
  assign n12778 = ~n12492 & ~n12777 ;
  assign n12779 = n8368 & ~n12691 ;
  assign n12780 = ~n12503 & ~n12779 ;
  assign n12781 = ~n12502 & n12780 ;
  assign n12782 = n12778 & n12781 ;
  assign n12783 = n12343 & ~n12782 ;
  assign n12784 = ~\pi0074  & ~\pi0075  ;
  assign n12785 = n1285 & n12784 ;
  assign n12786 = ~n12701 & ~n12703 ;
  assign n12787 = ~n12523 & ~n12786 ;
  assign n12788 = n8496 & ~n12787 ;
  assign n12789 = ~n12640 & n12788 ;
  assign n12790 = ~n12630 & n12789 ;
  assign n12791 = ~n12785 & ~n12790 ;
  assign n12792 = n12653 & ~n12787 ;
  assign n12793 = ~n12652 & n12792 ;
  assign n12794 = \pi0039  & n12523 ;
  assign n12795 = ~n12708 & ~n12794 ;
  assign n12796 = n6785 & n12795 ;
  assign n12797 = ~n12793 & n12796 ;
  assign n12798 = \pi0038  & ~n12523 ;
  assign n12799 = ~n12786 & n12798 ;
  assign n12800 = \pi0038  & ~\pi0039  ;
  assign n12801 = ~n12599 & n12800 ;
  assign n12802 = ~\pi0087  & ~n12801 ;
  assign n12803 = ~n12799 & n12802 ;
  assign n12804 = ~n12797 & n12803 ;
  assign n12805 = ~n12791 & n12804 ;
  assign n12806 = ~n12783 & n12805 ;
  assign n12807 = ~n12610 & n12806 ;
  assign n12808 = ~n12679 & ~n12787 ;
  assign n12809 = ~\pi0075  & ~n12808 ;
  assign n12810 = ~n12791 & ~n12809 ;
  assign n12811 = n12523 & n12684 ;
  assign n12812 = ~n12734 & ~n12811 ;
  assign n12813 = n12409 & n12812 ;
  assign n12814 = ~n12810 & n12813 ;
  assign n12815 = ~n12807 & n12814 ;
  assign n12816 = ~n12776 & ~n12815 ;
  assign n12817 = ~n12579 & ~n12816 ;
  assign n12818 = n9948 & ~n12817 ;
  assign n12819 = n12738 & n12818 ;
  assign n12820 = n12500 & ~n12579 ;
  assign n12821 = \pi0039  & ~n12820 ;
  assign n12822 = ~n9948 & ~n12625 ;
  assign n12823 = ~n12821 & n12822 ;
  assign n12824 = ~n12819 & ~n12823 ;
  assign n12825 = \pi0228  & n2327 ;
  assign n12826 = n1328 & n2575 ;
  assign n12827 = n1324 & n12826 ;
  assign n12828 = n1319 & n12827 ;
  assign n12829 = n12825 & n12828 ;
  assign n12830 = \pi0044  & ~\pi0072  ;
  assign n12831 = n1801 & n12512 ;
  assign n12832 = n2167 & n12692 ;
  assign n12833 = ~n12831 & ~n12832 ;
  assign n12834 = \pi0087  & n8640 ;
  assign n12835 = ~n12833 & n12834 ;
  assign n12836 = ~n8812 & ~n12835 ;
  assign n12837 = n12830 & ~n12836 ;
  assign n12838 = ~n12829 & n12837 ;
  assign n12839 = ~\pi0075  & n12836 ;
  assign n12840 = ~\pi0044  & \pi0228  ;
  assign n12841 = n2327 & n12840 ;
  assign n12842 = n1281 & n12841 ;
  assign n12843 = n1260 & n12842 ;
  assign n12844 = ~\pi0039  & ~\pi0075  ;
  assign n12845 = ~n12843 & n12844 ;
  assign n12846 = ~n12839 & ~n12845 ;
  assign n12847 = ~n12838 & ~n12846 ;
  assign n12848 = \pi0039  & n8640 ;
  assign n12849 = ~n12833 & n12848 ;
  assign n12850 = n6785 & ~n12849 ;
  assign n12851 = \pi0299  & ~n12830 ;
  assign n12852 = n1801 & n12851 ;
  assign n12853 = ~\pi0299  & ~n12830 ;
  assign n12854 = n2167 & n12853 ;
  assign n12855 = ~n12852 & ~n12854 ;
  assign n12856 = n8640 & ~n12855 ;
  assign n12857 = ~\pi0228  & ~n12830 ;
  assign n12858 = ~\pi0039  & ~n12857 ;
  assign n12859 = ~n12856 & n12858 ;
  assign n12860 = n12850 & ~n12859 ;
  assign n12861 = n8799 & ~n12043 ;
  assign n12862 = ~n6808 & n12861 ;
  assign n12863 = n8588 & n12041 ;
  assign n12864 = n1281 & n12863 ;
  assign n12865 = n1260 & n12864 ;
  assign n12866 = n12862 & n12865 ;
  assign n12867 = ~\pi0095  & \pi1093  ;
  assign n12868 = n1634 & n12867 ;
  assign n12869 = n8588 & n12868 ;
  assign n12870 = n1627 & n12869 ;
  assign n12871 = n1319 & n12870 ;
  assign n12872 = n8799 & n12830 ;
  assign n12873 = ~n6808 & n12872 ;
  assign n12874 = ~n12871 & n12873 ;
  assign n12875 = ~n12866 & ~n12874 ;
  assign n12876 = ~n8799 & n12830 ;
  assign n12877 = \pi0228  & ~n12876 ;
  assign n12878 = ~n8641 & n12877 ;
  assign n12879 = n12850 & n12878 ;
  assign n12880 = n12875 & n12879 ;
  assign n12881 = ~n12860 & ~n12880 ;
  assign n12882 = n12800 & ~n12830 ;
  assign n12883 = \pi0038  & \pi0039  ;
  assign n12884 = ~n12882 & ~n12883 ;
  assign n12885 = n8640 & ~n12882 ;
  assign n12886 = ~n12833 & n12885 ;
  assign n12887 = ~n12884 & ~n12886 ;
  assign n12888 = ~\pi0087  & ~n12887 ;
  assign n12889 = n12881 & n12888 ;
  assign n12890 = n12847 & ~n12889 ;
  assign n12891 = ~\pi0044  & ~n12313 ;
  assign n12892 = ~n12108 & n12830 ;
  assign n12893 = n12124 & n12892 ;
  assign n12894 = ~\pi0228  & ~n12893 ;
  assign n12895 = ~n12891 & n12894 ;
  assign n12896 = ~\pi0039  & ~n12895 ;
  assign n12897 = ~\pi0228  & n12896 ;
  assign n12898 = \pi1093  & ~n12040 ;
  assign n12899 = ~\pi1093  & n12051 ;
  assign n12900 = \pi0044  & ~n12899 ;
  assign n12901 = ~n12898 & n12900 ;
  assign n12902 = ~n12058 & ~n12064 ;
  assign n12903 = n8799 & ~n12902 ;
  assign n12904 = ~n12901 & n12903 ;
  assign n12905 = ~\pi0072  & ~n12048 ;
  assign n12906 = \pi0044  & n12905 ;
  assign n12907 = ~n12899 & n12906 ;
  assign n12908 = ~n8799 & n12080 ;
  assign n12909 = ~n12591 & ~n12908 ;
  assign n12910 = ~n12907 & ~n12909 ;
  assign n12911 = n12896 & ~n12910 ;
  assign n12912 = ~n12904 & n12911 ;
  assign n12913 = ~n12897 & ~n12912 ;
  assign n12914 = ~\pi0095  & \pi0287  ;
  assign n12915 = n1634 & n12914 ;
  assign n12916 = n1328 & n12915 ;
  assign n12917 = n1324 & n12916 ;
  assign n12918 = n1319 & n12917 ;
  assign n12919 = n12849 & ~n12918 ;
  assign n12920 = n2327 & ~n12919 ;
  assign n12921 = n12847 & n12920 ;
  assign n12922 = n12913 & n12921 ;
  assign n12923 = ~n12890 & ~n12922 ;
  assign n12924 = n8640 & ~n12833 ;
  assign n12925 = \pi0039  & ~n8496 ;
  assign n12926 = ~n12924 & n12925 ;
  assign n12927 = ~\pi0039  & ~n12830 ;
  assign n12928 = ~n8496 & n12927 ;
  assign n12929 = n9948 & ~n12928 ;
  assign n12930 = ~n12926 & n12929 ;
  assign n12931 = ~n2363 & ~n12927 ;
  assign n12932 = ~\pi0039  & n12931 ;
  assign n12933 = n8640 & n12931 ;
  assign n12934 = ~n12833 & n12933 ;
  assign n12935 = ~n12932 & ~n12934 ;
  assign n12936 = \pi0075  & ~n2363 ;
  assign n12937 = n12935 & n12936 ;
  assign n12938 = n12859 & ~n12878 ;
  assign n12939 = \pi0075  & ~n12849 ;
  assign n12940 = n12935 & n12939 ;
  assign n12941 = ~n12938 & n12940 ;
  assign n12942 = ~n12937 & ~n12941 ;
  assign n12943 = ~\pi0024  & n12863 ;
  assign n12944 = n1281 & n12943 ;
  assign n12945 = n1260 & n12944 ;
  assign n12946 = n7207 & n12945 ;
  assign n12947 = \pi0044  & ~n12211 ;
  assign n12948 = ~n12946 & ~n12947 ;
  assign n12949 = n12859 & n12862 ;
  assign n12950 = ~n12937 & n12949 ;
  assign n12951 = ~n12948 & n12950 ;
  assign n12952 = ~n12942 & ~n12951 ;
  assign n12953 = n12930 & ~n12952 ;
  assign n12954 = n12923 & n12953 ;
  assign n12955 = ~n8496 & n12929 ;
  assign n12956 = ~n12926 & n12955 ;
  assign n12957 = ~\pi0072  & ~\pi0166  ;
  assign n12958 = n1800 & n12957 ;
  assign n12959 = n8640 & n12958 ;
  assign n12960 = \pi0039  & ~n12959 ;
  assign n12961 = ~n9948 & ~n12927 ;
  assign n12962 = ~n12960 & n12961 ;
  assign n12963 = ~n12956 & ~n12962 ;
  assign n12964 = ~n12954 & n12963 ;
  assign n12965 = ~\pi0287  & n1281 ;
  assign n12966 = n1260 & n12965 ;
  assign n12967 = ~\pi0100  & n9627 ;
  assign n12968 = n2324 & n12967 ;
  assign n12969 = ~\pi0057  & n2511 ;
  assign n12970 = n6848 & n12969 ;
  assign n12971 = n12968 & n12970 ;
  assign n12972 = \pi0979  & n12971 ;
  assign n12973 = n12966 & n12972 ;
  assign n12974 = ~\pi0049  & ~\pi0076  ;
  assign n12975 = n10031 & n12974 ;
  assign n12976 = ~\pi0102  & ~\pi0104  ;
  assign n12977 = ~\pi0111  & n12976 ;
  assign n12978 = n12975 & n12977 ;
  assign n12979 = ~\pi0071  & n1256 ;
  assign n12980 = n8567 & n12979 ;
  assign n12981 = n12978 & n12980 ;
  assign n12982 = n1270 & n11929 ;
  assign n12983 = n1315 & n12982 ;
  assign n12984 = n12981 & n12983 ;
  assign n12985 = ~\pi0083  & ~\pi0089  ;
  assign n12986 = \pi0061  & ~\pi0082  ;
  assign n12987 = n12985 & n12986 ;
  assign n12988 = n1252 & n10039 ;
  assign n12989 = n12987 & n12988 ;
  assign n12990 = n10045 & n12989 ;
  assign n12991 = ~\pi0841  & n11921 ;
  assign n12992 = n12990 & n12991 ;
  assign n12993 = n12984 & n12992 ;
  assign n12994 = \pi0024  & n1270 ;
  assign n12995 = n8567 & n12994 ;
  assign n12996 = ~\pi0097  & n12995 ;
  assign n12997 = n1586 & n12996 ;
  assign n12998 = ~n12993 & ~n12997 ;
  assign n12999 = n11824 & ~n12998 ;
  assign n13000 = ~n6930 & ~n8543 ;
  assign n13001 = n1264 & n1329 ;
  assign n13002 = n9012 & n13001 ;
  assign n13003 = n1324 & n13002 ;
  assign n13004 = ~n13000 & ~n13003 ;
  assign n13005 = ~n11815 & ~n13000 ;
  assign n13006 = ~n11819 & n13005 ;
  assign n13007 = ~n13004 & ~n13006 ;
  assign n13008 = n11822 & n13007 ;
  assign n13009 = ~\pi0047  & \pi0088  ;
  assign n13010 = ~\pi0048  & ~\pi0089  ;
  assign n13011 = ~\pi0082  & n13010 ;
  assign n13012 = n1239 & n13011 ;
  assign n13013 = ~\pi0084  & \pi0104  ;
  assign n13014 = n1420 & n13013 ;
  assign n13015 = n11837 & n13014 ;
  assign n13016 = n13012 & n13015 ;
  assign n13017 = ~\pi0036  & ~n13016 ;
  assign n13018 = ~n1469 & ~n13017 ;
  assign n13019 = ~\pi0071  & n1423 ;
  assign n13020 = n11803 & n13019 ;
  assign n13021 = ~\pi0067  & ~\pi0103  ;
  assign n13022 = n1256 & n13021 ;
  assign n13023 = ~\pi0098  & n13022 ;
  assign n13024 = n13020 & n13023 ;
  assign n13025 = ~\pi0047  & n13024 ;
  assign n13026 = n13018 & n13025 ;
  assign n13027 = ~n13009 & ~n13026 ;
  assign n13028 = ~\pi0088  & n1252 ;
  assign n13029 = n1326 & n13028 ;
  assign n13030 = ~\pi0098  & n1252 ;
  assign n13031 = n1326 & n13030 ;
  assign n13032 = n1542 & n13031 ;
  assign n13033 = ~n13029 & ~n13032 ;
  assign n13034 = n1389 & ~n13033 ;
  assign n13035 = ~n13027 & n13034 ;
  assign n13036 = ~n11819 & ~n13035 ;
  assign n13037 = ~n9012 & n12138 ;
  assign n13038 = n1266 & n13037 ;
  assign n13039 = n11822 & n13038 ;
  assign n13040 = ~n13036 & n13039 ;
  assign n13041 = ~n13008 & ~n13040 ;
  assign n13042 = n1266 & n12138 ;
  assign n13043 = n8627 & ~n13042 ;
  assign n13044 = n8627 & ~n11819 ;
  assign n13045 = ~n13035 & n13044 ;
  assign n13046 = ~n13043 & ~n13045 ;
  assign n13047 = \pi1091  & ~n13046 ;
  assign n13048 = ~n6809 & n12138 ;
  assign n13049 = n1266 & n13048 ;
  assign n13050 = ~n13036 & n13049 ;
  assign n13051 = n1542 & n13030 ;
  assign n13052 = ~n13028 & ~n13051 ;
  assign n13053 = ~\pi0824  & n6809 ;
  assign n13054 = n1281 & n13053 ;
  assign n13055 = ~\pi0036  & ~\pi0098  ;
  assign n13056 = n13022 & n13055 ;
  assign n13057 = n13020 & n13056 ;
  assign n13058 = n13016 & n13057 ;
  assign n13059 = ~\pi0088  & ~n13058 ;
  assign n13060 = n13054 & ~n13059 ;
  assign n13061 = ~n13052 & n13060 ;
  assign n13062 = \pi0829  & ~n1686 ;
  assign n13063 = ~n13061 & n13062 ;
  assign n13064 = \pi1091  & n13063 ;
  assign n13065 = ~n13050 & n13064 ;
  assign n13066 = ~n13047 & ~n13065 ;
  assign n13067 = ~\pi0829  & ~n13038 ;
  assign n13068 = ~\pi0829  & ~n11819 ;
  assign n13069 = ~n13035 & n13068 ;
  assign n13070 = ~n13067 & ~n13069 ;
  assign n13071 = ~\pi1093  & ~n13070 ;
  assign n13072 = \pi0829  & ~n13061 ;
  assign n13073 = ~\pi1093  & n13072 ;
  assign n13074 = ~n13050 & n13073 ;
  assign n13075 = ~n13071 & ~n13074 ;
  assign n13076 = n13066 & n13075 ;
  assign n13077 = ~n13041 & n13076 ;
  assign n13078 = n11843 & n11932 ;
  assign n13079 = \pi0841  & n11822 ;
  assign n13080 = n1281 & n13079 ;
  assign n13081 = n13078 & n13080 ;
  assign n13082 = ~\pi0024  & \pi0074  ;
  assign n13083 = n1281 & n13082 ;
  assign n13084 = n1260 & n13083 ;
  assign n13085 = ~\pi0036  & n13021 ;
  assign n13086 = n11929 & n13085 ;
  assign n13087 = n10031 & n10038 ;
  assign n13088 = n13086 & n13087 ;
  assign n13089 = n1254 & n1256 ;
  assign n13090 = ~\pi0045  & ~\pi0111  ;
  assign n13091 = n12976 & n13090 ;
  assign n13092 = \pi0049  & n13091 ;
  assign n13093 = n13089 & n13092 ;
  assign n13094 = n13088 & n13093 ;
  assign n13095 = ~\pi0110  & n1261 ;
  assign n13096 = n12100 & n13095 ;
  assign n13097 = n1315 & n13012 ;
  assign n13098 = n13096 & n13097 ;
  assign n13099 = n13094 & n13098 ;
  assign n13100 = n1266 & n1320 ;
  assign n13101 = ~\pi0074  & \pi0841  ;
  assign n13102 = n13100 & n13101 ;
  assign n13103 = n13099 & n13102 ;
  assign n13104 = ~n13084 & ~n13103 ;
  assign n13105 = n2403 & n9948 ;
  assign n13106 = ~n13104 & n13105 ;
  assign n13107 = \pi0252  & ~n10050 ;
  assign n13108 = ~n1696 & n13107 ;
  assign n13109 = ~\pi0252  & n6808 ;
  assign n13110 = ~\pi0252  & n8640 ;
  assign n13111 = n8639 & n13110 ;
  assign n13112 = ~n13109 & ~n13111 ;
  assign n13113 = ~n13108 & n13112 ;
  assign n13114 = n1270 & n8567 ;
  assign n13115 = n1315 & n13114 ;
  assign n13116 = \pi0024  & n12138 ;
  assign n13117 = n1266 & n13116 ;
  assign n13118 = n13115 & n13117 ;
  assign n13119 = ~\pi0100  & n13118 ;
  assign n13120 = n10062 & n13119 ;
  assign n13121 = ~n13113 & n13120 ;
  assign n13122 = ~\pi0100  & n1261 ;
  assign n13123 = n1266 & n13122 ;
  assign n13124 = n1351 & n13123 ;
  assign n13125 = ~n13108 & n13124 ;
  assign n13126 = n13112 & n13125 ;
  assign n13127 = ~\pi0060  & n1274 ;
  assign n13128 = \pi0024  & ~\pi0053  ;
  assign n13129 = \pi0050  & n13128 ;
  assign n13130 = n1543 & n13129 ;
  assign n13131 = n1542 & n13130 ;
  assign n13132 = n13127 & n13131 ;
  assign n13133 = ~n1580 & ~n13132 ;
  assign n13134 = n13126 & ~n13133 ;
  assign n13135 = ~n13121 & ~n13134 ;
  assign n13136 = n10093 & n10094 ;
  assign n13137 = n10092 & n13136 ;
  assign n13138 = n10091 & n13137 ;
  assign n13139 = \pi0100  & n10092 ;
  assign n13140 = n7217 & n13139 ;
  assign n13141 = ~n13138 & ~n13140 ;
  assign n13142 = n13135 & n13141 ;
  assign n13143 = n1286 & n1288 ;
  assign n13144 = n10017 & n13143 ;
  assign n13145 = n10017 & n13137 ;
  assign n13146 = n10091 & n13145 ;
  assign n13147 = ~n13144 & ~n13146 ;
  assign n13148 = ~n13142 & ~n13147 ;
  assign n13149 = n11824 & n13115 ;
  assign n13150 = ~\pi0071  & n1244 ;
  assign n13151 = n11803 & n13150 ;
  assign n13152 = n13089 & n13151 ;
  assign n13153 = ~\pi0069  & n1424 ;
  assign n13154 = n13152 & n13153 ;
  assign n13155 = n1422 & n13154 ;
  assign n13156 = n13149 & n13155 ;
  assign n13157 = \pi0052  & ~\pi0072  ;
  assign n13158 = ~n6803 & ~n13157 ;
  assign n13159 = \pi0052  & ~\pi0228  ;
  assign n13160 = ~n13158 & n13159 ;
  assign n13161 = ~n12263 & n13160 ;
  assign n13162 = n12265 & n13160 ;
  assign n13163 = n12308 & n13162 ;
  assign n13164 = ~n13161 & ~n13163 ;
  assign n13165 = \pi0228  & ~n13158 ;
  assign n13166 = ~\pi0228  & ~n13158 ;
  assign n13167 = ~\pi0039  & ~n13166 ;
  assign n13168 = n6800 & n6807 ;
  assign n13169 = ~n12313 & n13168 ;
  assign n13170 = ~\pi0039  & n6803 ;
  assign n13171 = ~n13169 & n13170 ;
  assign n13172 = ~n13167 & ~n13171 ;
  assign n13173 = ~n13165 & ~n13172 ;
  assign n13174 = n13164 & n13173 ;
  assign n13175 = n2327 & n13174 ;
  assign n13176 = \pi0052  & ~n8799 ;
  assign n13177 = n12272 & n13176 ;
  assign n13178 = \pi0052  & n8799 ;
  assign n13179 = n12289 & n13178 ;
  assign n13180 = ~n13177 & ~n13179 ;
  assign n13181 = n13164 & ~n13172 ;
  assign n13182 = n6800 & n12592 ;
  assign n13183 = n13181 & ~n13182 ;
  assign n13184 = n8799 & n13181 ;
  assign n13185 = ~n12587 & n13184 ;
  assign n13186 = ~n13183 & ~n13185 ;
  assign n13187 = n6803 & ~n13186 ;
  assign n13188 = n2327 & n13187 ;
  assign n13189 = n13180 & n13188 ;
  assign n13190 = ~n13175 & ~n13189 ;
  assign n13191 = \pi0100  & n6803 ;
  assign n13192 = n12583 & n13191 ;
  assign n13193 = ~n8641 & n13192 ;
  assign n13194 = n12362 & n13193 ;
  assign n13195 = n12361 & n13194 ;
  assign n13196 = \pi0100  & ~n13157 ;
  assign n13197 = ~\pi0039  & ~n13196 ;
  assign n13198 = ~n13195 & n13197 ;
  assign n13199 = ~\pi0038  & ~n13198 ;
  assign n13200 = n11407 & n13157 ;
  assign n13201 = ~n2855 & ~n13200 ;
  assign n13202 = ~\pi0075  & ~n13201 ;
  assign n13203 = ~n13199 & n13202 ;
  assign n13204 = n13190 & n13203 ;
  assign n13205 = ~\pi0039  & n13157 ;
  assign n13206 = \pi0087  & \pi0100  ;
  assign n13207 = n13205 & n13206 ;
  assign n13208 = ~\pi0075  & n13207 ;
  assign n13209 = n6804 & n12430 ;
  assign n13210 = n1281 & n13209 ;
  assign n13211 = n1260 & n13210 ;
  assign n13212 = ~\pi0038  & ~n13211 ;
  assign n13213 = \pi0038  & ~n13205 ;
  assign n13214 = ~n13212 & ~n13213 ;
  assign n13215 = n12421 & n12668 ;
  assign n13216 = n13157 & ~n13213 ;
  assign n13217 = ~n13215 & n13216 ;
  assign n13218 = ~n13214 & ~n13217 ;
  assign n13219 = \pi0100  & ~n13205 ;
  assign n13220 = \pi0087  & ~n12967 ;
  assign n13221 = ~n13219 & n13220 ;
  assign n13222 = ~\pi0075  & n13221 ;
  assign n13223 = ~n13218 & n13222 ;
  assign n13224 = ~n13208 & ~n13223 ;
  assign n13225 = n12275 & n12446 ;
  assign n13226 = n6803 & n12583 ;
  assign n13227 = ~n8641 & n13226 ;
  assign n13228 = n13225 & n13227 ;
  assign n13229 = n12211 & n13228 ;
  assign n13230 = ~\pi0116  & n2363 ;
  assign n13231 = n13229 & n13230 ;
  assign n13232 = n12442 & n13157 ;
  assign n13233 = ~n13231 & n13232 ;
  assign n13234 = n8496 & ~n13233 ;
  assign n13235 = n13224 & n13234 ;
  assign n13236 = ~n13204 & n13235 ;
  assign n13237 = ~n8496 & ~n13205 ;
  assign n13238 = ~n12255 & n12577 ;
  assign n13239 = n12409 & ~n13238 ;
  assign n13240 = ~n13237 & n13239 ;
  assign n13241 = ~n13236 & n13240 ;
  assign n13242 = n13180 & n13187 ;
  assign n13243 = \pi0039  & n10276 ;
  assign n13244 = ~n12500 & n13243 ;
  assign n13245 = ~n12497 & n13244 ;
  assign n13246 = \pi0039  & ~n12504 ;
  assign n13247 = n2327 & ~n13246 ;
  assign n13248 = ~n13245 & n13247 ;
  assign n13249 = n6803 & n11690 ;
  assign n13250 = n12583 & n13249 ;
  assign n13251 = ~n8641 & n13250 ;
  assign n13252 = n12362 & n13251 ;
  assign n13253 = n12361 & n13252 ;
  assign n13254 = n13248 & ~n13253 ;
  assign n13255 = ~n13174 & n13254 ;
  assign n13256 = ~n13242 & n13255 ;
  assign n13257 = ~\pi0039  & ~n13157 ;
  assign n13258 = ~n2327 & ~n13257 ;
  assign n13259 = ~n12524 & n13258 ;
  assign n13260 = ~n13253 & n13259 ;
  assign n13261 = ~\pi0087  & ~n13260 ;
  assign n13262 = ~n13256 & n13261 ;
  assign n13263 = \pi0087  & ~n13258 ;
  assign n13264 = \pi0039  & \pi0087  ;
  assign n13265 = ~n12523 & n13264 ;
  assign n13266 = ~n13263 & ~n13265 ;
  assign n13267 = ~\pi0039  & ~n13211 ;
  assign n13268 = ~\pi0039  & n2327 ;
  assign n13269 = n2327 & n12512 ;
  assign n13270 = ~n12499 & n13269 ;
  assign n13271 = ~n13268 & ~n13270 ;
  assign n13272 = ~n13267 & ~n13271 ;
  assign n13273 = n13157 & ~n13271 ;
  assign n13274 = ~n13215 & n13273 ;
  assign n13275 = ~n13272 & ~n13274 ;
  assign n13276 = ~n13266 & n13275 ;
  assign n13277 = n12409 & ~n13276 ;
  assign n13278 = ~n13262 & n13277 ;
  assign n13279 = \pi0039  & ~n12782 ;
  assign n13280 = ~n12703 & ~n13257 ;
  assign n13281 = ~n12701 & n13280 ;
  assign n13282 = ~n12514 & n13213 ;
  assign n13283 = ~n13281 & n13282 ;
  assign n13284 = ~n6785 & ~n13283 ;
  assign n13285 = n12583 & n13170 ;
  assign n13286 = ~n8641 & n13285 ;
  assign n13287 = n12362 & n13286 ;
  assign n13288 = n12361 & n13287 ;
  assign n13289 = ~n12787 & ~n13283 ;
  assign n13290 = ~n13257 & n13289 ;
  assign n13291 = ~n13288 & n13290 ;
  assign n13292 = ~n13284 & ~n13291 ;
  assign n13293 = ~n13279 & ~n13292 ;
  assign n13294 = ~n13174 & n13293 ;
  assign n13295 = ~n13242 & n13294 ;
  assign n13296 = ~\pi0087  & n2327 ;
  assign n13297 = ~\pi0087  & ~n13284 ;
  assign n13298 = ~n13291 & n13297 ;
  assign n13299 = ~n13296 & ~n13298 ;
  assign n13300 = ~n13295 & ~n13299 ;
  assign n13301 = ~n12703 & n13258 ;
  assign n13302 = ~n12701 & n13301 ;
  assign n13303 = ~n13266 & ~n13302 ;
  assign n13304 = ~n12409 & ~n13303 ;
  assign n13305 = ~n12409 & n12523 ;
  assign n13306 = ~n12409 & ~n12703 ;
  assign n13307 = ~n12701 & n13306 ;
  assign n13308 = ~n13305 & ~n13307 ;
  assign n13309 = n2327 & ~n13267 ;
  assign n13310 = n2327 & n13157 ;
  assign n13311 = ~n13215 & n13310 ;
  assign n13312 = ~n13309 & ~n13311 ;
  assign n13313 = ~n13308 & ~n13312 ;
  assign n13314 = ~n13304 & ~n13313 ;
  assign n13315 = ~n13300 & ~n13314 ;
  assign n13316 = ~n13278 & ~n13315 ;
  assign n13317 = ~n12523 & n12925 ;
  assign n13318 = ~n8496 & n13257 ;
  assign n13319 = ~\pi0075  & n13238 ;
  assign n13320 = ~n13318 & n13319 ;
  assign n13321 = ~n13317 & n13320 ;
  assign n13322 = ~n13316 & n13321 ;
  assign n13323 = \pi0039  & ~n12697 ;
  assign n13324 = \pi0038  & ~n13281 ;
  assign n13325 = ~\pi0087  & ~n13324 ;
  assign n13326 = n13281 & n13325 ;
  assign n13327 = ~n13288 & n13326 ;
  assign n13328 = ~\pi0087  & ~n6785 ;
  assign n13329 = ~n13324 & n13328 ;
  assign n13330 = ~n13327 & ~n13329 ;
  assign n13331 = ~n13323 & ~n13330 ;
  assign n13332 = ~n13174 & n13331 ;
  assign n13333 = ~n13242 & n13332 ;
  assign n13334 = ~n2327 & ~n13330 ;
  assign n13335 = \pi0087  & n2327 ;
  assign n13336 = ~n12703 & n13335 ;
  assign n13337 = ~n12701 & n13336 ;
  assign n13338 = ~n13267 & n13337 ;
  assign n13339 = n13157 & n13337 ;
  assign n13340 = ~n13215 & n13339 ;
  assign n13341 = ~n13338 & ~n13340 ;
  assign n13342 = \pi0075  & n13157 ;
  assign n13343 = ~n12703 & n13342 ;
  assign n13344 = ~n12701 & n13343 ;
  assign n13345 = ~n13231 & n13344 ;
  assign n13346 = \pi0039  & \pi0075  ;
  assign n13347 = ~n12694 & n13346 ;
  assign n13348 = ~n12701 & n13347 ;
  assign n13349 = \pi0087  & n13302 ;
  assign n13350 = ~n13348 & ~n13349 ;
  assign n13351 = ~n13345 & n13350 ;
  assign n13352 = n13341 & n13351 ;
  assign n13353 = ~n13334 & n13352 ;
  assign n13354 = ~n13333 & n13353 ;
  assign n13355 = \pi0075  & ~n13348 ;
  assign n13356 = ~n13345 & n13355 ;
  assign n13357 = n8496 & ~n12409 ;
  assign n13358 = ~n13356 & n13357 ;
  assign n13359 = ~n13354 & n13358 ;
  assign n13360 = ~n13238 & n13359 ;
  assign n13361 = n13238 & ~n13318 ;
  assign n13362 = ~n13317 & n13361 ;
  assign n13363 = n12549 & n13281 ;
  assign n13364 = n9948 & ~n13363 ;
  assign n13365 = ~n13362 & n13364 ;
  assign n13366 = \pi0232  & ~n12700 ;
  assign n13367 = ~n12409 & ~n12694 ;
  assign n13368 = ~n13366 & n13367 ;
  assign n13369 = n12524 & ~n13368 ;
  assign n13370 = \pi0075  & ~n13369 ;
  assign n13371 = n13157 & n13370 ;
  assign n13372 = ~n13231 & n13371 ;
  assign n13373 = n13346 & ~n13369 ;
  assign n13374 = n8496 & ~n13373 ;
  assign n13375 = n13364 & n13374 ;
  assign n13376 = ~n13372 & n13375 ;
  assign n13377 = ~n13365 & ~n13376 ;
  assign n13378 = ~n13360 & ~n13377 ;
  assign n13379 = ~n13322 & n13378 ;
  assign n13380 = ~n13241 & n13379 ;
  assign n13381 = \pi0039  & n13238 ;
  assign n13382 = n12500 & n13381 ;
  assign n13383 = ~n9948 & ~n13205 ;
  assign n13384 = ~n13382 & n13383 ;
  assign n13385 = ~n13380 & ~n13384 ;
  assign n13386 = n11858 & n11903 ;
  assign n13387 = n1261 & n11828 ;
  assign n13388 = n1320 & n13387 ;
  assign n13389 = n1266 & n13388 ;
  assign n13390 = \pi0053  & ~\pi0058  ;
  assign n13391 = n1274 & n13390 ;
  assign n13392 = n1273 & n13391 ;
  assign n13393 = n13389 & n13392 ;
  assign n13394 = n1564 & n13393 ;
  assign n13395 = ~\pi0287  & ~\pi0979  ;
  assign n13396 = n6717 & n13395 ;
  assign n13397 = \pi0039  & n13396 ;
  assign n13398 = n1281 & n13397 ;
  assign n13399 = n1260 & n13398 ;
  assign n13400 = ~n13394 & ~n13399 ;
  assign n13401 = n13386 & ~n13400 ;
  assign n13402 = n10042 & n13086 ;
  assign n13403 = ~\pi0060  & ~\pi0085  ;
  assign n13404 = \pi0106  & n13403 ;
  assign n13405 = n1231 & n10034 ;
  assign n13406 = n13404 & n13405 ;
  assign n13407 = n12975 & n13406 ;
  assign n13408 = n13402 & n13407 ;
  assign n13409 = n13089 & n13408 ;
  assign n13410 = ~\pi0058  & ~\pi0094  ;
  assign n13411 = n1344 & n13410 ;
  assign n13412 = n1273 & n13411 ;
  assign n13413 = ~\pi0841  & n1320 ;
  assign n13414 = n1266 & n13413 ;
  assign n13415 = n2342 & n7265 ;
  assign n13416 = n1261 & n13415 ;
  assign n13417 = n13414 & n13416 ;
  assign n13418 = n13412 & n13417 ;
  assign n13419 = n13409 & n13418 ;
  assign n13420 = n2363 & n8322 ;
  assign n13421 = n11830 & n13420 ;
  assign n13422 = n1627 & n13421 ;
  assign n13423 = n1319 & n13422 ;
  assign n13424 = ~n13419 & ~n13423 ;
  assign n13425 = n11858 & ~n13424 ;
  assign n13426 = n13042 & n13115 ;
  assign n13427 = \pi0045  & n1256 ;
  assign n13428 = n1231 & n13427 ;
  assign n13429 = n1444 & n13428 ;
  assign n13430 = n13088 & n13429 ;
  assign n13431 = ~\pi0102  & n2404 ;
  assign n13432 = n1254 & n13431 ;
  assign n13433 = n2403 & n13432 ;
  assign n13434 = n10125 & n13433 ;
  assign n13435 = n13430 & n13434 ;
  assign n13436 = n13426 & n13435 ;
  assign n13437 = n1328 & n11829 ;
  assign n13438 = n1324 & n13437 ;
  assign n13439 = n1319 & n13438 ;
  assign n13440 = n1329 & n2363 ;
  assign n13441 = n2364 & n2511 ;
  assign n13442 = \pi0055  & n13441 ;
  assign n13443 = n10125 & n13442 ;
  assign n13444 = n13440 & n13443 ;
  assign n13445 = n13439 & n13444 ;
  assign n13446 = ~n13436 & ~n13445 ;
  assign n13447 = n1264 & n2404 ;
  assign n13448 = n2403 & n13447 ;
  assign n13449 = n10023 & n13448 ;
  assign n13450 = n1358 & n13449 ;
  assign n13451 = \pi0056  & ~n13450 ;
  assign n13452 = \pi0056  & ~\pi0062  ;
  assign n13453 = n2467 & n13452 ;
  assign n13454 = ~\pi0024  & n1292 ;
  assign n13455 = n1291 & n13454 ;
  assign n13456 = \pi0055  & n2467 ;
  assign n13457 = n13455 & n13456 ;
  assign n13458 = n1281 & n13457 ;
  assign n13459 = n1260 & n13458 ;
  assign n13460 = ~n13453 & ~n13459 ;
  assign n13461 = ~n13451 & ~n13460 ;
  assign n13462 = n7265 & n10015 ;
  assign n13463 = n13440 & n13462 ;
  assign n13464 = n13439 & n13463 ;
  assign n13465 = n7672 & n13464 ;
  assign n13466 = ~\pi0056  & \pi0062  ;
  assign n13467 = ~\pi0924  & n13466 ;
  assign n13468 = ~n13452 & ~n13467 ;
  assign n13469 = n2467 & ~n13468 ;
  assign n13470 = n13448 & n13469 ;
  assign n13471 = n10909 & n13470 ;
  assign n13472 = ~n13465 & ~n13471 ;
  assign n13473 = \pi0090  & n8555 ;
  assign n13474 = n10903 & n13473 ;
  assign n13475 = n11822 & n13474 ;
  assign n13476 = n10893 & n13475 ;
  assign n13477 = n1319 & n13476 ;
  assign n13478 = \pi0924  & n13466 ;
  assign n13479 = n13447 & n13478 ;
  assign n13480 = n2403 & n13479 ;
  assign n13481 = n2467 & n13480 ;
  assign n13482 = n10909 & n13481 ;
  assign n13483 = ~\pi0057  & \pi0059  ;
  assign n13484 = n13464 & n13483 ;
  assign n13485 = ~n13482 & ~n13484 ;
  assign n13486 = n13389 & n13412 ;
  assign n13487 = n1559 & n13486 ;
  assign n13488 = \pi0039  & ~\pi0979  ;
  assign n13489 = n6715 & ~n6717 ;
  assign n13490 = n13488 & n13489 ;
  assign n13491 = ~\pi0287  & n13490 ;
  assign n13492 = n1281 & n13491 ;
  assign n13493 = n1260 & n13492 ;
  assign n13494 = ~n13487 & ~n13493 ;
  assign n13495 = n13386 & ~n13494 ;
  assign n13496 = \pi0841  & n11921 ;
  assign n13497 = n12990 & n13496 ;
  assign n13498 = n12984 & n13497 ;
  assign n13499 = ~\pi0024  & n13410 ;
  assign n13500 = n1344 & n13499 ;
  assign n13501 = n1273 & n13500 ;
  assign n13502 = n1347 & n13501 ;
  assign n13503 = n1249 & n13502 ;
  assign n13504 = ~n13498 & ~n13503 ;
  assign n13505 = n11824 & ~n13504 ;
  assign n13506 = n13447 & n13466 ;
  assign n13507 = n2403 & n13506 ;
  assign n13508 = n10023 & n13507 ;
  assign n13509 = n1358 & n13508 ;
  assign n13510 = n2467 & n13509 ;
  assign n13511 = n7672 & n11798 ;
  assign n13512 = ~n13510 & ~n13511 ;
  assign n13513 = \pi0999  & n1255 ;
  assign n13514 = n13115 & n13513 ;
  assign n13515 = n1513 & n13514 ;
  assign n13516 = ~\pi0024  & n1270 ;
  assign n13517 = n8567 & n13516 ;
  assign n13518 = ~\pi0097  & n13517 ;
  assign n13519 = n1586 & n13518 ;
  assign n13520 = ~n13515 & ~n13519 ;
  assign n13521 = n11824 & ~n13520 ;
  assign n13522 = ~\pi0064  & ~\pi0107  ;
  assign n13523 = ~\pi0063  & ~\pi0081  ;
  assign n13524 = ~n13522 & n13523 ;
  assign n13525 = n1236 & n13524 ;
  assign n13526 = n1248 & n13525 ;
  assign n13527 = ~\pi0102  & n1254 ;
  assign n13528 = ~\pi0107  & \pi0841  ;
  assign n13529 = \pi0064  & ~n13528 ;
  assign n13530 = n1257 & ~n13529 ;
  assign n13531 = n13527 & n13530 ;
  assign n13532 = n13526 & n13531 ;
  assign n13533 = n13149 & n13532 ;
  assign n13534 = \pi0299  & n11859 ;
  assign n13535 = n12971 & n13534 ;
  assign n13536 = ~n11895 & n13535 ;
  assign n13537 = n11877 & n13536 ;
  assign n13538 = ~\pi0299  & n11859 ;
  assign n13539 = n12971 & n13538 ;
  assign n13540 = ~n11883 & n13539 ;
  assign n13541 = n11877 & n13540 ;
  assign n13542 = ~n13537 & ~n13541 ;
  assign n13543 = ~\pi0102  & \pi0314  ;
  assign n13544 = n1254 & n13543 ;
  assign n13545 = n13426 & n13544 ;
  assign n13546 = \pi0081  & n1257 ;
  assign n13547 = n1525 & n13546 ;
  assign n13548 = n1236 & n13547 ;
  assign n13549 = n1248 & n13548 ;
  assign n13550 = ~\pi0199  & ~\pi0299  ;
  assign n13551 = n1291 & ~n13550 ;
  assign n13552 = n13549 & n13551 ;
  assign n13553 = n13545 & n13552 ;
  assign n13554 = \pi0219  & ~n13553 ;
  assign n13555 = ~\pi0057  & \pi0219  ;
  assign n13556 = n6848 & n13555 ;
  assign n13557 = n2327 & n13441 ;
  assign n13558 = \pi0199  & ~\pi0299  ;
  assign n13559 = n2341 & n13558 ;
  assign n13560 = n13557 & n13559 ;
  assign n13561 = n9948 & n13560 ;
  assign n13562 = n13549 & n13561 ;
  assign n13563 = n13545 & n13562 ;
  assign n13564 = ~n13556 & ~n13563 ;
  assign n13565 = ~n13554 & ~n13564 ;
  assign n13566 = \pi0083  & ~\pi0103  ;
  assign n13567 = ~\pi0071  & n13566 ;
  assign n13568 = n11803 & n13567 ;
  assign n13569 = n13089 & n13568 ;
  assign n13570 = n11822 & n13569 ;
  assign n13571 = n1236 & n1245 ;
  assign n13572 = n1471 & n13571 ;
  assign n13573 = n13570 & n13572 ;
  assign n13574 = \pi0314  & n1254 ;
  assign n13575 = n13426 & n13574 ;
  assign n13576 = n13573 & n13575 ;
  assign n13577 = ~n6744 & n6932 ;
  assign n13578 = n2256 & n2291 ;
  assign n13579 = n13577 & n13578 ;
  assign n13580 = n6921 & n13579 ;
  assign n13581 = ~n6770 & n6932 ;
  assign n13582 = n2522 & n3058 ;
  assign n13583 = n13581 & n13582 ;
  assign n13584 = n6921 & n13583 ;
  assign n13585 = ~n13580 & ~n13584 ;
  assign n13586 = n12971 & ~n13585 ;
  assign n13587 = n1252 & n11805 ;
  assign n13588 = \pi0071  & \pi0314  ;
  assign n13589 = n1236 & n13588 ;
  assign n13590 = n1248 & n13589 ;
  assign n13591 = n13587 & n13590 ;
  assign n13592 = n13149 & n13591 ;
  assign n13593 = ~\pi0081  & ~\pi0314  ;
  assign n13594 = ~\pi0102  & n13593 ;
  assign n13595 = n1254 & n13594 ;
  assign n13596 = ~\pi0071  & n13595 ;
  assign n13597 = n1236 & n13595 ;
  assign n13598 = n1248 & n13597 ;
  assign n13599 = ~n13596 & ~n13598 ;
  assign n13600 = n6989 & ~n13599 ;
  assign n13601 = \pi0069  & ~\pi0103  ;
  assign n13602 = ~\pi0036  & ~\pi0083  ;
  assign n13603 = n13601 & n13602 ;
  assign n13604 = ~\pi0067  & n13603 ;
  assign n13605 = n1466 & n13604 ;
  assign n13606 = n1459 & n13605 ;
  assign n13607 = ~\pi0071  & ~n13606 ;
  assign n13608 = n13149 & ~n13607 ;
  assign n13609 = n13600 & n13608 ;
  assign n13610 = ~n13592 & ~n13609 ;
  assign n13611 = \pi0070  & ~\pi0096  ;
  assign n13612 = n1261 & n13611 ;
  assign n13613 = n1354 & n13612 ;
  assign n13614 = n1358 & n13613 ;
  assign n13615 = n11830 & n13386 ;
  assign n13616 = n13614 & n13615 ;
  assign n13617 = \pi0198  & \pi0589  ;
  assign n13618 = n2214 & n13617 ;
  assign n13619 = ~n8387 & n13618 ;
  assign n13620 = \pi0210  & \pi0589  ;
  assign n13621 = ~\pi0216  & \pi0299  ;
  assign n13622 = n1295 & n13621 ;
  assign n13623 = n6706 & n13622 ;
  assign n13624 = ~n6732 & n13623 ;
  assign n13625 = ~n6706 & n13622 ;
  assign n13626 = ~n6713 & n13625 ;
  assign n13627 = ~n13624 & ~n13626 ;
  assign n13628 = n13620 & ~n13627 ;
  assign n13629 = ~n13619 & ~n13628 ;
  assign n13630 = ~n1696 & ~n6925 ;
  assign n13631 = ~\pi0593  & \pi0835  ;
  assign n13632 = ~n6717 & n13631 ;
  assign n13633 = n6716 & n13632 ;
  assign n13634 = ~n13630 & n13633 ;
  assign n13635 = ~n13629 & n13634 ;
  assign n13636 = ~\pi0287  & ~n13635 ;
  assign n13637 = n1259 & n13386 ;
  assign n13638 = n1249 & n13637 ;
  assign n13639 = n2595 & n13638 ;
  assign n13640 = ~n13636 & n13639 ;
  assign n13641 = ~n13616 & ~n13640 ;
  assign n13642 = ~n1448 & ~n1449 ;
  assign n13643 = \pi0085  & n13022 ;
  assign n13644 = n1236 & n13643 ;
  assign n13645 = ~\pi0199  & \pi0200  ;
  assign n13646 = ~\pi0299  & n13645 ;
  assign n13647 = \pi0211  & ~\pi0219  ;
  assign n13648 = \pi0299  & n13647 ;
  assign n13649 = ~n13646 & ~n13648 ;
  assign n13650 = n13574 & n13649 ;
  assign n13651 = n13020 & n13650 ;
  assign n13652 = n13644 & n13651 ;
  assign n13653 = n13426 & n13652 ;
  assign n13654 = ~n13642 & n13653 ;
  assign n13655 = \pi0299  & \pi0314  ;
  assign n13656 = n13647 & n13655 ;
  assign n13657 = ~\pi0299  & \pi0314  ;
  assign n13658 = n13645 & n13657 ;
  assign n13659 = ~n13656 & ~n13658 ;
  assign n13660 = \pi0081  & ~n13659 ;
  assign n13661 = n13042 & n13660 ;
  assign n13662 = ~\pi0102  & n1253 ;
  assign n13663 = n1252 & n1270 ;
  assign n13664 = n8567 & n13663 ;
  assign n13665 = n1315 & n13664 ;
  assign n13666 = n13662 & n13665 ;
  assign n13667 = ~n1529 & n13666 ;
  assign n13668 = n13661 & n13667 ;
  assign n13669 = n1449 & n13644 ;
  assign n13670 = ~n1434 & n13644 ;
  assign n13671 = n1447 & n13670 ;
  assign n13672 = ~n13669 & ~n13671 ;
  assign n13673 = ~\pi0064  & n10038 ;
  assign n13674 = ~n13659 & n13673 ;
  assign n13675 = n13042 & n13674 ;
  assign n13676 = n13667 & n13675 ;
  assign n13677 = ~n13672 & n13676 ;
  assign n13678 = ~n13668 & ~n13677 ;
  assign n13679 = ~n13654 & n13678 ;
  assign n13680 = n11822 & ~n13679 ;
  assign n13681 = ~\pi0039  & ~n2575 ;
  assign n13682 = \pi0024  & \pi0072  ;
  assign n13683 = n1328 & n13682 ;
  assign n13684 = n1324 & n13683 ;
  assign n13685 = n1319 & n13684 ;
  assign n13686 = \pi0088  & n13665 ;
  assign n13687 = n6925 & n10369 ;
  assign n13688 = ~\pi0098  & n13687 ;
  assign n13689 = n13686 & n13688 ;
  assign n13690 = n1542 & n13689 ;
  assign n13691 = ~\pi0039  & ~n13690 ;
  assign n13692 = ~n13685 & n13691 ;
  assign n13693 = ~n13681 & ~n13692 ;
  assign n13694 = ~\pi0039  & n2467 ;
  assign n13695 = n10015 & n13694 ;
  assign n13696 = n11903 & n13695 ;
  assign n13697 = ~n8793 & n13386 ;
  assign n13698 = n6948 & n13697 ;
  assign n13699 = ~n13696 & ~n13698 ;
  assign n13700 = n13693 & ~n13699 ;
  assign n13701 = n2297 & n7597 ;
  assign n13702 = n13577 & n13701 ;
  assign n13703 = n6921 & n13702 ;
  assign n13704 = n6205 & n6955 ;
  assign n13705 = n13581 & n13704 ;
  assign n13706 = n6921 & n13705 ;
  assign n13707 = ~n13703 & ~n13706 ;
  assign n13708 = ~\pi0040  & n1264 ;
  assign n13709 = ~\pi0314  & \pi1050  ;
  assign n13710 = ~\pi0039  & n13709 ;
  assign n13711 = n13708 & n13710 ;
  assign n13712 = n10937 & n13711 ;
  assign n13713 = n10319 & n13712 ;
  assign n13714 = n13707 & ~n13713 ;
  assign n13715 = n13386 & ~n13714 ;
  assign n13716 = n1329 & n7267 ;
  assign n13717 = n2363 & n13716 ;
  assign n13718 = n13439 & n13717 ;
  assign n13719 = n9948 & n13718 ;
  assign n13720 = ~n1696 & ~n10050 ;
  assign n13721 = ~\pi0096  & ~\pi1093  ;
  assign n13722 = n9012 & n13721 ;
  assign n13723 = n1291 & ~n13722 ;
  assign n13724 = ~\pi0096  & ~n6684 ;
  assign n13725 = \pi0479  & ~n13724 ;
  assign n13726 = n13723 & ~n13725 ;
  assign n13727 = n13720 & n13726 ;
  assign n13728 = n13001 & n13727 ;
  assign n13729 = ~n8582 & n13728 ;
  assign n13730 = n1720 & n8733 ;
  assign n13731 = ~\pi0096  & ~n13730 ;
  assign n13732 = n9948 & ~n13731 ;
  assign n13733 = n13729 & n13732 ;
  assign n13734 = ~n13719 & ~n13733 ;
  assign n13735 = n13439 & n13440 ;
  assign n13736 = \pi0075  & ~n13735 ;
  assign n13737 = n10017 & ~n13736 ;
  assign n13738 = \pi1093  & ~n8799 ;
  assign n13739 = n2342 & ~n13738 ;
  assign n13740 = n8739 & n13739 ;
  assign n13741 = \pi1093  & n1720 ;
  assign n13742 = n8733 & n13741 ;
  assign n13743 = ~\pi0096  & ~n13742 ;
  assign n13744 = n13740 & ~n13743 ;
  assign n13745 = n8742 & n13744 ;
  assign n13746 = ~\pi0075  & ~n13745 ;
  assign n13747 = n13737 & ~n13746 ;
  assign n13748 = n1281 & n10047 ;
  assign n13749 = \pi0122  & \pi0137  ;
  assign n13750 = \pi0137  & ~\pi1093  ;
  assign n13751 = n6811 & n13750 ;
  assign n13752 = ~n13749 & ~n13751 ;
  assign n13753 = n13748 & ~n13752 ;
  assign n13754 = ~\pi0210  & ~n6808 ;
  assign n13755 = ~n13753 & n13754 ;
  assign n13756 = ~\pi0210  & n6807 ;
  assign n13757 = n6804 & n13756 ;
  assign n13758 = ~n13755 & ~n13757 ;
  assign n13759 = \pi0252  & \pi0829  ;
  assign n13760 = n6809 & n13759 ;
  assign n13761 = n1261 & ~n13760 ;
  assign n13762 = n1266 & n13761 ;
  assign n13763 = n1351 & n13762 ;
  assign n13764 = ~\pi0137  & n13763 ;
  assign n13765 = n1580 & n13764 ;
  assign n13766 = ~\pi0137  & \pi1091  ;
  assign n13767 = ~n1686 & n13766 ;
  assign n13768 = ~n13765 & n13767 ;
  assign n13769 = n8799 & ~n13765 ;
  assign n13770 = ~n13768 & ~n13769 ;
  assign n13771 = n1267 & n1351 ;
  assign n13772 = n1276 & n10047 ;
  assign n13773 = ~n1580 & ~n13772 ;
  assign n13774 = n13771 & ~n13773 ;
  assign n13775 = \pi0122  & ~n8675 ;
  assign n13776 = ~n13774 & n13775 ;
  assign n13777 = ~\pi0252  & n13771 ;
  assign n13778 = ~n13773 & n13777 ;
  assign n13779 = \pi0252  & n13748 ;
  assign n13780 = \pi0122  & n8675 ;
  assign n13781 = ~n13779 & n13780 ;
  assign n13782 = ~n13778 & n13781 ;
  assign n13783 = ~n13776 & ~n13782 ;
  assign n13784 = ~\pi1093  & ~n13783 ;
  assign n13785 = n8675 & ~n13779 ;
  assign n13786 = ~n13778 & n13785 ;
  assign n13787 = n8752 & ~n13774 ;
  assign n13788 = n1542 & n1568 ;
  assign n13789 = n1261 & n1578 ;
  assign n13790 = n1266 & n13789 ;
  assign n13791 = n1351 & n13790 ;
  assign n13792 = n13788 & n13791 ;
  assign n13793 = ~n6811 & ~n13792 ;
  assign n13794 = ~n13787 & ~n13793 ;
  assign n13795 = ~n13786 & n13794 ;
  assign n13796 = ~\pi0122  & ~\pi1093  ;
  assign n13797 = ~n13795 & n13796 ;
  assign n13798 = ~n13784 & ~n13797 ;
  assign n13799 = n1580 & n13763 ;
  assign n13800 = ~\pi0122  & ~n13799 ;
  assign n13801 = n13783 & ~n13800 ;
  assign n13802 = \pi1093  & ~n13801 ;
  assign n13803 = ~n13768 & ~n13802 ;
  assign n13804 = n13798 & n13803 ;
  assign n13805 = ~n13770 & ~n13804 ;
  assign n13806 = ~\pi0122  & n13791 ;
  assign n13807 = n13788 & n13806 ;
  assign n13808 = \pi1093  & ~n13807 ;
  assign n13809 = \pi0122  & n13771 ;
  assign n13810 = ~n13773 & n13809 ;
  assign n13811 = n13808 & ~n13810 ;
  assign n13812 = \pi0137  & ~n13811 ;
  assign n13813 = ~n13784 & n13812 ;
  assign n13814 = ~n13797 & n13813 ;
  assign n13815 = \pi0252  & \pi1092  ;
  assign n13816 = ~\pi1093  & n13815 ;
  assign n13817 = n1687 & n13816 ;
  assign n13818 = ~\pi0137  & ~n13817 ;
  assign n13819 = n13791 & n13818 ;
  assign n13820 = n13788 & n13819 ;
  assign n13821 = ~n8799 & ~n13820 ;
  assign n13822 = ~n13814 & n13821 ;
  assign n13823 = ~n13755 & ~n13822 ;
  assign n13824 = ~n13805 & n13823 ;
  assign n13825 = ~n13758 & ~n13824 ;
  assign n13826 = n13798 & ~n13802 ;
  assign n13827 = n6807 & n8799 ;
  assign n13828 = n6804 & n13827 ;
  assign n13829 = ~n13826 & n13828 ;
  assign n13830 = ~n11744 & n13748 ;
  assign n13831 = ~n6808 & ~n13830 ;
  assign n13832 = ~n13784 & ~n13811 ;
  assign n13833 = ~n13797 & n13832 ;
  assign n13834 = n6807 & ~n8799 ;
  assign n13835 = n6804 & n13834 ;
  assign n13836 = ~n13833 & n13835 ;
  assign n13837 = ~n13831 & ~n13836 ;
  assign n13838 = ~n13829 & n13837 ;
  assign n13839 = \pi0210  & ~n13838 ;
  assign n13840 = ~\pi0232  & ~n13839 ;
  assign n13841 = ~n13825 & n13840 ;
  assign n13842 = ~n8368 & ~n13841 ;
  assign n13843 = \pi0299  & n9250 ;
  assign n13844 = ~\pi0198  & ~n6808 ;
  assign n13845 = ~n13753 & n13844 ;
  assign n13846 = \pi0198  & ~n13838 ;
  assign n13847 = ~n13845 & ~n13846 ;
  assign n13848 = ~n13805 & ~n13822 ;
  assign n13849 = ~\pi0198  & n6807 ;
  assign n13850 = n6804 & n13849 ;
  assign n13851 = ~n13848 & n13850 ;
  assign n13852 = n9250 & ~n13851 ;
  assign n13853 = n13847 & n13852 ;
  assign n13854 = ~n13843 & ~n13853 ;
  assign n13855 = ~n13842 & ~n13854 ;
  assign n13856 = ~n13825 & ~n13839 ;
  assign n13857 = n1800 & n11984 ;
  assign n13858 = ~n13856 & ~n13857 ;
  assign n13859 = ~\pi0210  & n13857 ;
  assign n13860 = ~n13848 & n13859 ;
  assign n13861 = \pi0299  & ~n13857 ;
  assign n13862 = \pi0210  & n8799 ;
  assign n13863 = ~n13826 & n13862 ;
  assign n13864 = \pi0210  & ~n8799 ;
  assign n13865 = ~n13833 & n13864 ;
  assign n13866 = \pi0299  & ~n13865 ;
  assign n13867 = ~n13863 & n13866 ;
  assign n13868 = ~n13861 & ~n13867 ;
  assign n13869 = ~n13860 & ~n13868 ;
  assign n13870 = ~n13858 & n13869 ;
  assign n13871 = \pi0232  & n9250 ;
  assign n13872 = n13870 & n13871 ;
  assign n13873 = n13847 & ~n13851 ;
  assign n13874 = n2167 & n6706 ;
  assign n13875 = ~n13873 & ~n13874 ;
  assign n13876 = ~\pi0198  & n13874 ;
  assign n13877 = ~n13848 & n13876 ;
  assign n13878 = \pi0198  & ~n8799 ;
  assign n13879 = ~n13833 & n13878 ;
  assign n13880 = n13874 & n13879 ;
  assign n13881 = \pi0198  & \pi1091  ;
  assign n13882 = ~n1686 & n13881 ;
  assign n13883 = n13874 & n13882 ;
  assign n13884 = ~n13826 & n13883 ;
  assign n13885 = ~n13880 & ~n13884 ;
  assign n13886 = ~\pi0299  & n13885 ;
  assign n13887 = ~n13877 & n13886 ;
  assign n13888 = n13871 & n13887 ;
  assign n13889 = ~n13875 & n13888 ;
  assign n13890 = ~n13872 & ~n13889 ;
  assign n13891 = ~n13855 & n13890 ;
  assign n13892 = ~n8675 & ~n13760 ;
  assign n13893 = ~n13760 & n13791 ;
  assign n13894 = n13788 & n13893 ;
  assign n13895 = ~n13892 & ~n13894 ;
  assign n13896 = n8642 & n13895 ;
  assign n13897 = n8642 & ~n8675 ;
  assign n13898 = ~n13774 & n13897 ;
  assign n13899 = ~n13896 & ~n13898 ;
  assign n13900 = n13783 & n13899 ;
  assign n13901 = \pi0137  & ~n13900 ;
  assign n13902 = ~n8675 & ~n13774 ;
  assign n13903 = ~n13786 & ~n13902 ;
  assign n13904 = n13750 & ~n13903 ;
  assign n13905 = ~\pi0137  & n13895 ;
  assign n13906 = ~\pi0137  & ~n8675 ;
  assign n13907 = ~n13774 & n13906 ;
  assign n13908 = ~n13905 & ~n13907 ;
  assign n13909 = ~n13904 & n13908 ;
  assign n13910 = ~n13901 & n13909 ;
  assign n13911 = n6808 & ~n13910 ;
  assign n13912 = \pi0137  & ~n8642 ;
  assign n13913 = n8675 & ~n13912 ;
  assign n13914 = n8799 & ~n13913 ;
  assign n13915 = n13748 & n13914 ;
  assign n13916 = ~n13828 & ~n13915 ;
  assign n13917 = ~\pi0210  & ~n13916 ;
  assign n13918 = ~n13911 & n13917 ;
  assign n13919 = n8799 & ~n13900 ;
  assign n13920 = ~\pi1093  & ~n13903 ;
  assign n13921 = n13738 & ~n13774 ;
  assign n13922 = n6808 & ~n13921 ;
  assign n13923 = ~n13920 & n13922 ;
  assign n13924 = ~n13919 & n13923 ;
  assign n13925 = ~n6808 & ~n11749 ;
  assign n13926 = n13748 & n13925 ;
  assign n13927 = ~n13924 & ~n13926 ;
  assign n13928 = \pi0210  & ~n13927 ;
  assign n13929 = ~n6808 & n13748 ;
  assign n13930 = ~\pi1093  & n6808 ;
  assign n13931 = n6808 & n13771 ;
  assign n13932 = ~n13773 & n13931 ;
  assign n13933 = ~n13930 & ~n13932 ;
  assign n13934 = ~\pi0137  & ~\pi1093  ;
  assign n13935 = n13895 & n13934 ;
  assign n13936 = ~n8675 & n13934 ;
  assign n13937 = ~n13774 & n13936 ;
  assign n13938 = ~n13935 & ~n13937 ;
  assign n13939 = ~n13933 & n13938 ;
  assign n13940 = ~n13904 & n13939 ;
  assign n13941 = ~n13929 & ~n13940 ;
  assign n13942 = ~\pi0137  & n10050 ;
  assign n13943 = ~n8799 & ~n13942 ;
  assign n13944 = ~n13835 & ~n13943 ;
  assign n13945 = ~\pi0210  & ~n13944 ;
  assign n13946 = ~n13941 & n13945 ;
  assign n13947 = ~n13928 & ~n13946 ;
  assign n13948 = ~n13918 & n13947 ;
  assign n13949 = ~n13857 & ~n13948 ;
  assign n13950 = n8799 & n13908 ;
  assign n13951 = ~n13904 & n13950 ;
  assign n13952 = ~n13901 & n13951 ;
  assign n13953 = ~\pi1093  & ~n8799 ;
  assign n13954 = ~n8799 & n13771 ;
  assign n13955 = ~n13773 & n13954 ;
  assign n13956 = ~n13953 & ~n13955 ;
  assign n13957 = n13938 & ~n13956 ;
  assign n13958 = ~n13904 & n13957 ;
  assign n13959 = ~\pi0210  & ~n13958 ;
  assign n13960 = ~n13952 & n13959 ;
  assign n13961 = ~n13920 & ~n13921 ;
  assign n13962 = ~n13919 & n13961 ;
  assign n13963 = \pi0210  & ~n13962 ;
  assign n13964 = n13857 & ~n13963 ;
  assign n13965 = ~n13960 & n13964 ;
  assign n13966 = \pi0299  & ~n13965 ;
  assign n13967 = ~n13949 & n13966 ;
  assign n13968 = ~\pi0198  & ~n13958 ;
  assign n13969 = ~n13952 & n13968 ;
  assign n13970 = n13882 & ~n13900 ;
  assign n13971 = \pi0198  & n13921 ;
  assign n13972 = \pi0198  & ~\pi1093  ;
  assign n13973 = ~n13903 & n13972 ;
  assign n13974 = ~n13971 & ~n13973 ;
  assign n13975 = n13874 & n13974 ;
  assign n13976 = ~n13970 & n13975 ;
  assign n13977 = ~n13969 & n13976 ;
  assign n13978 = n13874 & ~n13977 ;
  assign n13979 = ~\pi0198  & ~n13944 ;
  assign n13980 = ~n13941 & n13979 ;
  assign n13981 = ~\pi0198  & ~n13916 ;
  assign n13982 = ~n13911 & n13981 ;
  assign n13983 = ~n13980 & ~n13982 ;
  assign n13984 = \pi0198  & ~n13927 ;
  assign n13985 = ~n13977 & ~n13984 ;
  assign n13986 = n13983 & n13985 ;
  assign n13987 = ~n13978 & ~n13986 ;
  assign n13988 = ~\pi0299  & ~n13987 ;
  assign n13989 = ~n13967 & ~n13988 ;
  assign n13990 = \pi0232  & ~n13989 ;
  assign n13991 = \pi0299  & ~n13948 ;
  assign n13992 = ~\pi0232  & \pi0299  ;
  assign n13993 = ~\pi0232  & ~n13984 ;
  assign n13994 = n13983 & n13993 ;
  assign n13995 = ~n13992 & ~n13994 ;
  assign n13996 = ~n13991 & ~n13995 ;
  assign n13997 = ~n9250 & ~n13996 ;
  assign n13998 = ~n13990 & n13997 ;
  assign n13999 = n13891 & ~n13998 ;
  assign n14000 = n11822 & ~n13999 ;
  assign n14001 = \pi0086  & n13114 ;
  assign n14002 = n1555 & n1567 ;
  assign n14003 = n13114 & n14002 ;
  assign n14004 = n1542 & n14003 ;
  assign n14005 = ~n14001 & ~n14004 ;
  assign n14006 = ~n7038 & ~n14005 ;
  assign n14007 = ~\pi0314  & ~n14006 ;
  assign n14008 = ~\pi0314  & n1322 ;
  assign n14009 = n10903 & n14008 ;
  assign n14010 = n11822 & n14009 ;
  assign n14011 = \pi0086  & n13410 ;
  assign n14012 = n1273 & n14011 ;
  assign n14013 = n11824 & n14012 ;
  assign n14014 = n13788 & n14013 ;
  assign n14015 = ~n14010 & ~n14014 ;
  assign n14016 = ~n14007 & ~n14015 ;
  assign n14017 = \pi0119  & \pi0232  ;
  assign n14018 = ~\pi0468  & n14017 ;
  assign n14019 = \pi0147  & \pi0232  ;
  assign n14020 = n6706 & n14019 ;
  assign n14021 = \pi0038  & ~n14020 ;
  assign n14022 = ~\pi0100  & ~n10155 ;
  assign n14023 = ~n14021 & n14022 ;
  assign n14024 = ~\pi0100  & ~n14023 ;
  assign n14025 = \pi0163  & ~n11126 ;
  assign n14026 = n6706 & ~n10114 ;
  assign n14027 = ~n11123 & n14026 ;
  assign n14028 = ~\pi0163  & ~n11121 ;
  assign n14029 = ~n14027 & n14028 ;
  assign n14030 = ~n14025 & ~n14029 ;
  assign n14031 = \pi0232  & ~n14023 ;
  assign n14032 = n14030 & n14031 ;
  assign n14033 = ~n14024 & ~n14032 ;
  assign n14034 = n8248 & n14033 ;
  assign n14035 = \pi0232  & n14030 ;
  assign n14036 = n11082 & ~n14035 ;
  assign n14037 = n11129 & n14030 ;
  assign n14038 = n8601 & ~n14020 ;
  assign n14039 = \pi0054  & ~n14038 ;
  assign n14040 = ~\pi0074  & ~n14039 ;
  assign n14041 = ~n14037 & ~n14040 ;
  assign n14042 = ~n14036 & ~n14041 ;
  assign n14043 = ~n14034 & n14042 ;
  assign n14044 = \pi0074  & n11129 ;
  assign n14045 = n14030 & n14044 ;
  assign n14046 = ~n1292 & ~n14045 ;
  assign n14047 = ~n14043 & n14046 ;
  assign n14048 = n2467 & ~n10159 ;
  assign n14049 = ~n14047 & n14048 ;
  assign n14050 = ~n11160 & n11161 ;
  assign n14051 = \pi0184  & n6706 ;
  assign n14052 = ~\pi0299  & ~n14051 ;
  assign n14053 = ~n14050 & n14052 ;
  assign n14054 = \pi0232  & ~n14053 ;
  assign n14055 = \pi0184  & ~\pi0299  ;
  assign n14056 = n14050 & n14055 ;
  assign n14057 = ~n8601 & ~n14056 ;
  assign n14058 = n14054 & n14057 ;
  assign n14059 = \pi0074  & ~n14058 ;
  assign n14060 = \pi0074  & \pi0299  ;
  assign n14061 = ~n14030 & n14060 ;
  assign n14062 = ~n14059 & ~n14061 ;
  assign n14063 = ~\pi0055  & n14062 ;
  assign n14064 = \pi0055  & ~\pi0074  ;
  assign n14065 = \pi0055  & n11129 ;
  assign n14066 = n14030 & n14065 ;
  assign n14067 = ~n14064 & ~n14066 ;
  assign n14068 = n1292 & n14067 ;
  assign n14069 = \pi0039  & ~n10543 ;
  assign n14070 = n2855 & ~n14069 ;
  assign n14071 = \pi0039  & n14070 ;
  assign n14072 = n10173 & n10217 ;
  assign n14073 = ~\pi0063  & ~\pi0107  ;
  assign n14074 = ~n14072 & n14073 ;
  assign n14075 = ~\pi0040  & ~n14074 ;
  assign n14076 = ~\pi0095  & ~n6706 ;
  assign n14077 = n10174 & n14076 ;
  assign n14078 = n10173 & n14077 ;
  assign n14079 = \pi0163  & \pi0232  ;
  assign n14080 = n10182 & n14079 ;
  assign n14081 = ~n14078 & n14080 ;
  assign n14082 = n14070 & ~n14081 ;
  assign n14083 = n14075 & n14082 ;
  assign n14084 = ~n14071 & ~n14083 ;
  assign n14085 = \pi0087  & ~n1256 ;
  assign n14086 = n10155 & n14085 ;
  assign n14087 = n2364 & ~n14086 ;
  assign n14088 = ~\pi0100  & ~n14021 ;
  assign n14089 = n14087 & n14088 ;
  assign n14090 = n14084 & n14089 ;
  assign n14091 = \pi0100  & n2364 ;
  assign n14092 = ~n14035 & n14091 ;
  assign n14093 = ~n10844 & ~n14033 ;
  assign n14094 = n6895 & ~n14093 ;
  assign n14095 = \pi0075  & ~n14035 ;
  assign n14096 = ~n14037 & n14039 ;
  assign n14097 = ~n14095 & ~n14096 ;
  assign n14098 = ~n14094 & n14097 ;
  assign n14099 = ~n14092 & n14098 ;
  assign n14100 = ~n14090 & n14099 ;
  assign n14101 = \pi0054  & n14038 ;
  assign n14102 = \pi0054  & n11129 ;
  assign n14103 = n14030 & n14102 ;
  assign n14104 = ~n14101 & ~n14103 ;
  assign n14105 = n10190 & n14104 ;
  assign n14106 = ~n14100 & n14105 ;
  assign n14107 = ~n14068 & ~n14106 ;
  assign n14108 = ~n14063 & ~n14107 ;
  assign n14109 = n14054 & ~n14056 ;
  assign n14110 = \pi0100  & ~n14109 ;
  assign n14111 = \pi0100  & \pi0299  ;
  assign n14112 = ~n14030 & n14111 ;
  assign n14113 = ~n14110 & ~n14112 ;
  assign n14114 = ~\pi0187  & ~\pi0299  ;
  assign n14115 = ~\pi0147  & \pi0299  ;
  assign n14116 = ~n14114 & ~n14115 ;
  assign n14117 = n8640 & n14116 ;
  assign n14118 = \pi0038  & ~n14117 ;
  assign n14119 = n11470 & ~n14086 ;
  assign n14120 = ~n14118 & n14119 ;
  assign n14121 = n14113 & ~n14120 ;
  assign n14122 = ~\pi0092  & ~n14121 ;
  assign n14123 = ~\pi0040  & ~n10454 ;
  assign n14124 = ~n10449 & n14123 ;
  assign n14125 = ~\pi0095  & ~n14124 ;
  assign n14126 = ~n10477 & n10479 ;
  assign n14127 = ~\pi0040  & \pi0166  ;
  assign n14128 = ~n14126 & n14127 ;
  assign n14129 = n14125 & ~n14128 ;
  assign n14130 = n6706 & ~n10555 ;
  assign n14131 = n10543 & n11984 ;
  assign n14132 = \pi0153  & ~n14131 ;
  assign n14133 = \pi0160  & ~n14132 ;
  assign n14134 = ~\pi0040  & n10452 ;
  assign n14135 = n10058 & n14134 ;
  assign n14136 = n10582 & n14135 ;
  assign n14137 = ~\pi0095  & ~n10543 ;
  assign n14138 = ~n14136 & n14137 ;
  assign n14139 = \pi0166  & n6706 ;
  assign n14140 = ~n10555 & n14139 ;
  assign n14141 = \pi0160  & n14140 ;
  assign n14142 = ~n14138 & n14141 ;
  assign n14143 = ~n14133 & ~n14142 ;
  assign n14144 = n14130 & ~n14143 ;
  assign n14145 = ~n14129 & n14144 ;
  assign n14146 = ~\pi0095  & ~\pi0153  ;
  assign n14147 = ~n14124 & n14146 ;
  assign n14148 = ~n14128 & n14147 ;
  assign n14149 = ~\pi0032  & n10360 ;
  assign n14150 = n1618 & n14149 ;
  assign n14151 = n10173 & n14150 ;
  assign n14152 = ~n1256 & n10356 ;
  assign n14153 = \pi0095  & ~n14152 ;
  assign n14154 = ~n1256 & n10360 ;
  assign n14155 = n14153 & ~n14154 ;
  assign n14156 = ~n14151 & n14155 ;
  assign n14157 = ~\pi0160  & n6706 ;
  assign n14158 = ~n14156 & n14157 ;
  assign n14159 = \pi0153  & n14138 ;
  assign n14160 = n10937 & n13708 ;
  assign n14161 = n10319 & n14160 ;
  assign n14162 = \pi0153  & ~\pi0166  ;
  assign n14163 = n14161 & n14162 ;
  assign n14164 = ~n14159 & ~n14163 ;
  assign n14165 = n14158 & n14164 ;
  assign n14166 = ~n14148 & n14165 ;
  assign n14167 = \pi0153  & ~n14143 ;
  assign n14168 = \pi0163  & ~n14167 ;
  assign n14169 = ~n14166 & n14168 ;
  assign n14170 = ~n14145 & n14169 ;
  assign n14171 = ~n10386 & n10561 ;
  assign n14172 = ~\pi0051  & n10561 ;
  assign n14173 = ~n10408 & n14172 ;
  assign n14174 = ~n14171 & ~n14173 ;
  assign n14175 = n1264 & n14174 ;
  assign n14176 = \pi0032  & ~\pi0095  ;
  assign n14177 = ~n10543 & n14176 ;
  assign n14178 = ~n10555 & ~n14177 ;
  assign n14179 = ~n14175 & n14178 ;
  assign n14180 = \pi0210  & ~n14179 ;
  assign n14181 = ~\pi0166  & \pi0210  ;
  assign n14182 = n6706 & n14181 ;
  assign n14183 = ~\pi0095  & n10556 ;
  assign n14184 = ~n10559 & n14183 ;
  assign n14185 = ~n10555 & n11984 ;
  assign n14186 = ~n14184 & n14185 ;
  assign n14187 = ~n14175 & n14186 ;
  assign n14188 = ~n14182 & ~n14187 ;
  assign n14189 = ~n14180 & ~n14188 ;
  assign n14190 = ~\pi0040  & ~n10692 ;
  assign n14191 = ~\pi0040  & ~\pi0210  ;
  assign n14192 = ~n10375 & n14191 ;
  assign n14193 = ~n14190 & ~n14192 ;
  assign n14194 = n14139 & ~n14193 ;
  assign n14195 = ~\pi0153  & ~n14194 ;
  assign n14196 = ~n14189 & n14195 ;
  assign n14197 = ~\pi0153  & \pi0160  ;
  assign n14198 = ~n10565 & n10699 ;
  assign n14199 = ~n10564 & n14198 ;
  assign n14200 = ~\pi0095  & \pi0210  ;
  assign n14201 = ~n10549 & n14200 ;
  assign n14202 = ~n10547 & n14201 ;
  assign n14203 = ~n14199 & ~n14202 ;
  assign n14204 = n14139 & n14203 ;
  assign n14205 = ~\pi0095  & \pi0160  ;
  assign n14206 = ~\pi0040  & \pi0160  ;
  assign n14207 = ~n1256 & n14206 ;
  assign n14208 = ~n14205 & ~n14207 ;
  assign n14209 = n14204 & ~n14208 ;
  assign n14210 = ~n10661 & n10699 ;
  assign n14211 = ~n10667 & n14200 ;
  assign n14212 = ~n14210 & ~n14211 ;
  assign n14213 = n11984 & ~n14208 ;
  assign n14214 = n14212 & n14213 ;
  assign n14215 = ~n14209 & ~n14214 ;
  assign n14216 = ~n14197 & n14215 ;
  assign n14217 = ~n14196 & ~n14216 ;
  assign n14218 = ~\pi0163  & ~n14217 ;
  assign n14219 = \pi0095  & ~n14156 ;
  assign n14220 = ~\pi0040  & ~n14156 ;
  assign n14221 = ~n10692 & n14220 ;
  assign n14222 = ~\pi0210  & n14220 ;
  assign n14223 = ~n10375 & n14222 ;
  assign n14224 = ~n14221 & ~n14223 ;
  assign n14225 = ~n14219 & n14224 ;
  assign n14226 = \pi0166  & ~n14225 ;
  assign n14227 = ~n14156 & ~n14184 ;
  assign n14228 = ~n14175 & n14227 ;
  assign n14229 = ~\pi0210  & ~n14228 ;
  assign n14230 = ~\pi0166  & ~\pi0210  ;
  assign n14231 = n6706 & n14230 ;
  assign n14232 = n11984 & ~n14156 ;
  assign n14233 = ~n14177 & n14232 ;
  assign n14234 = ~n14175 & n14233 ;
  assign n14235 = ~n14231 & ~n14234 ;
  assign n14236 = ~n14229 & ~n14235 ;
  assign n14237 = ~n14226 & ~n14236 ;
  assign n14238 = ~\pi0153  & n14237 ;
  assign n14239 = ~\pi0153  & ~\pi0160  ;
  assign n14240 = ~\pi0160  & ~n14156 ;
  assign n14241 = n14204 & n14240 ;
  assign n14242 = n11984 & n14240 ;
  assign n14243 = n14212 & n14242 ;
  assign n14244 = ~n14241 & ~n14243 ;
  assign n14245 = ~n14239 & n14244 ;
  assign n14246 = ~n14238 & ~n14245 ;
  assign n14247 = n14218 & ~n14246 ;
  assign n14248 = ~n14170 & ~n14247 ;
  assign n14249 = \pi0299  & ~n14219 ;
  assign n14250 = n14224 & n14249 ;
  assign n14251 = ~n8377 & ~n14250 ;
  assign n14252 = ~n14248 & ~n14251 ;
  assign n14253 = ~\pi0198  & n14220 ;
  assign n14254 = ~n10375 & n14253 ;
  assign n14255 = ~n14221 & ~n14254 ;
  assign n14256 = ~n14219 & n14255 ;
  assign n14257 = ~n12330 & ~n14256 ;
  assign n14258 = ~\pi0198  & ~n14228 ;
  assign n14259 = ~\pi0189  & ~\pi0198  ;
  assign n14260 = n6706 & n14259 ;
  assign n14261 = n12330 & ~n14156 ;
  assign n14262 = ~n14177 & n14261 ;
  assign n14263 = ~n14175 & n14262 ;
  assign n14264 = ~n14260 & ~n14263 ;
  assign n14265 = ~n14258 & ~n14264 ;
  assign n14266 = ~\pi0175  & ~\pi0299  ;
  assign n14267 = ~\pi0184  & n14266 ;
  assign n14268 = ~\pi0182  & n14267 ;
  assign n14269 = ~n14265 & n14268 ;
  assign n14270 = ~n14257 & n14269 ;
  assign n14271 = ~n6706 & ~n14256 ;
  assign n14272 = \pi0095  & ~\pi0182  ;
  assign n14273 = ~\pi0095  & \pi0189  ;
  assign n14274 = n1256 & ~n14273 ;
  assign n14275 = n10543 & ~n14274 ;
  assign n14276 = n14135 & ~n14274 ;
  assign n14277 = n10582 & n14276 ;
  assign n14278 = ~n14275 & ~n14277 ;
  assign n14279 = ~n14272 & n14278 ;
  assign n14280 = ~n14152 & n14272 ;
  assign n14281 = ~n14154 & n14280 ;
  assign n14282 = ~n14151 & n14281 ;
  assign n14283 = n14051 & ~n14282 ;
  assign n14284 = ~n14279 & n14283 ;
  assign n14285 = \pi0175  & ~\pi0299  ;
  assign n14286 = ~n14284 & n14285 ;
  assign n14287 = n12330 & ~n14282 ;
  assign n14288 = ~n10662 & n14287 ;
  assign n14289 = n10670 & n14288 ;
  assign n14290 = n12330 & n14272 ;
  assign n14291 = ~n14282 & n14290 ;
  assign n14292 = n10421 & ~n10565 ;
  assign n14293 = ~n10564 & n14292 ;
  assign n14294 = ~n10549 & n10668 ;
  assign n14295 = ~n10547 & n14294 ;
  assign n14296 = ~n14293 & ~n14295 ;
  assign n14297 = \pi0189  & n6706 ;
  assign n14298 = \pi0095  & \pi0182  ;
  assign n14299 = ~n10543 & n14298 ;
  assign n14300 = ~n14282 & ~n14299 ;
  assign n14301 = n14297 & n14300 ;
  assign n14302 = n14296 & n14301 ;
  assign n14303 = ~n14291 & ~n14302 ;
  assign n14304 = ~n14289 & n14303 ;
  assign n14305 = ~\pi0184  & ~n14304 ;
  assign n14306 = n14286 & ~n14305 ;
  assign n14307 = ~n14271 & n14306 ;
  assign n14308 = ~\pi0040  & \pi0189  ;
  assign n14309 = ~n14126 & n14308 ;
  assign n14310 = n14125 & ~n14309 ;
  assign n14311 = n6706 & ~n14299 ;
  assign n14312 = ~n14282 & n14311 ;
  assign n14313 = ~n14310 & n14312 ;
  assign n14314 = \pi0184  & ~n14313 ;
  assign n14315 = ~n10555 & ~n14184 ;
  assign n14316 = ~n14175 & n14315 ;
  assign n14317 = ~\pi0198  & n12330 ;
  assign n14318 = n14316 & n14317 ;
  assign n14319 = \pi0198  & n12330 ;
  assign n14320 = n14179 & n14319 ;
  assign n14321 = ~n14318 & ~n14320 ;
  assign n14322 = \pi0182  & ~\pi0184  ;
  assign n14323 = ~n10375 & n10571 ;
  assign n14324 = ~n14190 & ~n14323 ;
  assign n14325 = n14297 & ~n14324 ;
  assign n14326 = n14322 & ~n14325 ;
  assign n14327 = n14321 & n14326 ;
  assign n14328 = ~n14314 & ~n14327 ;
  assign n14329 = n14266 & ~n14271 ;
  assign n14330 = ~n14328 & n14329 ;
  assign n14331 = ~n14307 & ~n14330 ;
  assign n14332 = ~n14270 & n14331 ;
  assign n14333 = ~n14252 & n14332 ;
  assign n14334 = ~\pi0040  & ~n6706 ;
  assign n14335 = ~n6713 & n14334 ;
  assign n14336 = n10217 & n14335 ;
  assign n14337 = n10231 & n14336 ;
  assign n14338 = ~\pi0189  & ~n10543 ;
  assign n14339 = ~n14337 & n14338 ;
  assign n14340 = ~n6709 & n10543 ;
  assign n14341 = n6735 & n14340 ;
  assign n14342 = ~n1256 & n14335 ;
  assign n14343 = ~n14337 & ~n14342 ;
  assign n14344 = ~n14341 & n14343 ;
  assign n14345 = \pi0189  & ~n6761 ;
  assign n14346 = n1256 & ~n10266 ;
  assign n14347 = n10496 & ~n14346 ;
  assign n14348 = n14345 & ~n14347 ;
  assign n14349 = n14344 & n14348 ;
  assign n14350 = ~n14339 & ~n14349 ;
  assign n14351 = \pi0179  & ~n14350 ;
  assign n14352 = ~\pi0040  & ~n1256 ;
  assign n14353 = ~\pi0040  & n10217 ;
  assign n14354 = n10231 & n14353 ;
  assign n14355 = ~n14352 & ~n14354 ;
  assign n14356 = ~n6736 & ~n14355 ;
  assign n14357 = ~\pi0179  & ~n6761 ;
  assign n14358 = ~n14341 & n14357 ;
  assign n14359 = ~n14356 & n14358 ;
  assign n14360 = n6761 & ~n10543 ;
  assign n14361 = ~n14337 & n14360 ;
  assign n14362 = ~\pi0179  & ~\pi0189  ;
  assign n14363 = ~n6761 & n14362 ;
  assign n14364 = ~n14361 & ~n14363 ;
  assign n14365 = ~n14359 & n14364 ;
  assign n14366 = n1256 & ~n10219 ;
  assign n14367 = n10496 & ~n14366 ;
  assign n14368 = n14344 & ~n14367 ;
  assign n14369 = ~\pi0189  & ~n14361 ;
  assign n14370 = ~n14368 & n14369 ;
  assign n14371 = ~n14365 & ~n14370 ;
  assign n14372 = ~n14351 & ~n14371 ;
  assign n14373 = \pi0224  & ~\pi0299  ;
  assign n14374 = n6949 & n14373 ;
  assign n14375 = ~n14372 & n14374 ;
  assign n14376 = ~n6955 & ~n10543 ;
  assign n14377 = ~\pi0299  & n14376 ;
  assign n14378 = ~n7597 & n10543 ;
  assign n14379 = \pi0299  & ~n14378 ;
  assign n14380 = \pi0166  & ~n6732 ;
  assign n14381 = ~n14347 & n14380 ;
  assign n14382 = n14344 & n14381 ;
  assign n14383 = ~n10543 & ~n14380 ;
  assign n14384 = ~n14337 & n14383 ;
  assign n14385 = n7597 & ~n14384 ;
  assign n14386 = ~n14382 & n14385 ;
  assign n14387 = n14379 & ~n14386 ;
  assign n14388 = ~n14377 & ~n14387 ;
  assign n14389 = ~n14375 & n14388 ;
  assign n14390 = \pi0156  & \pi0232  ;
  assign n14391 = ~n14389 & n14390 ;
  assign n14392 = n6955 & n14361 ;
  assign n14393 = ~n6761 & ~n14341 ;
  assign n14394 = n6955 & n14393 ;
  assign n14395 = ~n14356 & n14394 ;
  assign n14396 = ~n14392 & ~n14395 ;
  assign n14397 = ~\pi0299  & ~n14376 ;
  assign n14398 = n14396 & n14397 ;
  assign n14399 = ~n6732 & ~n14341 ;
  assign n14400 = ~n14356 & n14399 ;
  assign n14401 = n6732 & ~n10543 ;
  assign n14402 = ~n14337 & n14401 ;
  assign n14403 = n10280 & ~n14402 ;
  assign n14404 = ~n14400 & n14403 ;
  assign n14405 = ~\pi0232  & ~n14404 ;
  assign n14406 = ~n14398 & n14405 ;
  assign n14407 = \pi0039  & ~n14406 ;
  assign n14408 = ~\pi0156  & \pi0232  ;
  assign n14409 = ~\pi0166  & ~n6732 ;
  assign n14410 = n14402 & ~n14409 ;
  assign n14411 = n14399 & ~n14409 ;
  assign n14412 = ~n14356 & n14411 ;
  assign n14413 = ~n14410 & ~n14412 ;
  assign n14414 = ~n14367 & n14409 ;
  assign n14415 = n14344 & n14414 ;
  assign n14416 = n7597 & ~n14415 ;
  assign n14417 = n14413 & n14416 ;
  assign n14418 = n14379 & ~n14417 ;
  assign n14419 = ~n14377 & ~n14418 ;
  assign n14420 = ~n14375 & n14419 ;
  assign n14421 = n14408 & ~n14420 ;
  assign n14422 = n14407 & ~n14421 ;
  assign n14423 = ~n14391 & n14422 ;
  assign n14424 = n9636 & ~n14423 ;
  assign n14425 = ~n14333 & n14424 ;
  assign n14426 = n8368 & ~n14219 ;
  assign n14427 = n14255 & n14426 ;
  assign n14428 = n13992 & ~n14219 ;
  assign n14429 = n14224 & n14428 ;
  assign n14430 = ~\pi0039  & ~n14429 ;
  assign n14431 = ~n14427 & n14430 ;
  assign n14432 = ~n14423 & ~n14431 ;
  assign n14433 = ~\pi0038  & n14432 ;
  assign n14434 = ~\pi0147  & \pi0187  ;
  assign n14435 = \pi0038  & n14434 ;
  assign n14436 = n10195 & n14435 ;
  assign n14437 = ~n8375 & n14436 ;
  assign n14438 = ~\pi0187  & ~n10201 ;
  assign n14439 = \pi0187  & n6784 ;
  assign n14440 = n1266 & n14439 ;
  assign n14441 = n1354 & n14440 ;
  assign n14442 = n1358 & n14441 ;
  assign n14443 = \pi0147  & ~\pi0187  ;
  assign n14444 = ~n14020 & ~n14443 ;
  assign n14445 = ~n14442 & ~n14444 ;
  assign n14446 = \pi0038  & n14445 ;
  assign n14447 = ~n14438 & n14446 ;
  assign n14448 = ~n14437 & ~n14447 ;
  assign n14449 = ~n14433 & n14448 ;
  assign n14450 = ~n14425 & n14449 ;
  assign n14451 = ~\pi0092  & n2362 ;
  assign n14452 = ~n14450 & n14451 ;
  assign n14453 = ~n14122 & ~n14452 ;
  assign n14454 = ~\pi0054  & ~\pi0075  ;
  assign n14455 = ~n14453 & n14454 ;
  assign n14456 = ~\pi0179  & ~\pi0299  ;
  assign n14457 = ~\pi0156  & \pi0299  ;
  assign n14458 = ~n14456 & ~n14457 ;
  assign n14459 = n8640 & n14458 ;
  assign n14460 = n1256 & n14459 ;
  assign n14461 = ~\pi0040  & ~n14460 ;
  assign n14462 = ~n14074 & n14461 ;
  assign n14463 = ~\pi0100  & ~n14086 ;
  assign n14464 = ~n14118 & n14463 ;
  assign n14465 = ~\pi0039  & n14464 ;
  assign n14466 = ~n14462 & n14465 ;
  assign n14467 = ~n14070 & n14464 ;
  assign n14468 = \pi0075  & ~n14109 ;
  assign n14469 = \pi0075  & \pi0299  ;
  assign n14470 = ~n14030 & n14469 ;
  assign n14471 = ~n14468 & ~n14470 ;
  assign n14472 = n14113 & n14471 ;
  assign n14473 = ~n14467 & n14472 ;
  assign n14474 = ~n14466 & n14473 ;
  assign n14475 = ~n6895 & n14471 ;
  assign n14476 = ~\pi0054  & ~n14475 ;
  assign n14477 = ~n14474 & n14476 ;
  assign n14478 = n8601 & ~n14117 ;
  assign n14479 = \pi0054  & ~n14478 ;
  assign n14480 = ~n14058 & n14479 ;
  assign n14481 = \pi0299  & n14479 ;
  assign n14482 = ~n14030 & n14481 ;
  assign n14483 = ~n14480 & ~n14482 ;
  assign n14484 = ~n14477 & n14483 ;
  assign n14485 = ~n14455 & n14484 ;
  assign n14486 = ~\pi0074  & ~n14107 ;
  assign n14487 = ~n14485 & n14486 ;
  assign n14488 = ~n14108 & ~n14487 ;
  assign n14489 = n14049 & n14488 ;
  assign n14490 = ~n2467 & n11129 ;
  assign n14491 = n14030 & n14490 ;
  assign n14492 = ~\pi0074  & ~n2467 ;
  assign n14493 = n14038 & n14492 ;
  assign n14494 = ~n14491 & ~n14493 ;
  assign n14495 = ~\pi0079  & n14494 ;
  assign n14496 = ~n14489 & n14495 ;
  assign n14497 = ~\pi0034  & n11506 ;
  assign n14498 = ~n10155 & n11470 ;
  assign n14499 = ~n14118 & n14498 ;
  assign n14500 = ~n2362 & ~n14499 ;
  assign n14501 = n2582 & n10414 ;
  assign n14502 = n1354 & n14501 ;
  assign n14503 = n1358 & n14502 ;
  assign n14504 = ~n6732 & n7597 ;
  assign n14505 = \pi0156  & \pi1091  ;
  assign n14506 = n1689 & n14505 ;
  assign n14507 = n1688 & n14506 ;
  assign n14508 = n6745 & n14507 ;
  assign n14509 = ~\pi0166  & n6922 ;
  assign n14510 = ~n6931 & n14509 ;
  assign n14511 = n6722 & n14510 ;
  assign n14512 = ~n14508 & ~n14511 ;
  assign n14513 = n14504 & ~n14512 ;
  assign n14514 = n14503 & n14513 ;
  assign n14515 = ~\pi0040  & \pi0299  ;
  assign n14516 = ~n14514 & n14515 ;
  assign n14517 = ~\pi0040  & ~\pi0299  ;
  assign n14518 = \pi0039  & ~n14517 ;
  assign n14519 = ~\pi0189  & n6922 ;
  assign n14520 = ~n6931 & n14519 ;
  assign n14521 = n6722 & n14520 ;
  assign n14522 = \pi0179  & \pi1091  ;
  assign n14523 = n1689 & n14522 ;
  assign n14524 = n1688 & n14523 ;
  assign n14525 = n6745 & n14524 ;
  assign n14526 = ~n14521 & ~n14525 ;
  assign n14527 = ~n6761 & n6955 ;
  assign n14528 = \pi0039  & n14527 ;
  assign n14529 = ~n14526 & n14528 ;
  assign n14530 = n14503 & n14529 ;
  assign n14531 = ~n14518 & ~n14530 ;
  assign n14532 = ~n14516 & ~n14531 ;
  assign n14533 = \pi0232  & ~n14532 ;
  assign n14534 = ~\pi0040  & ~\pi0232  ;
  assign n14535 = ~\pi0038  & ~n14534 ;
  assign n14536 = ~n14533 & n14535 ;
  assign n14537 = ~\pi0210  & ~n10914 ;
  assign n14538 = ~n10913 & n14537 ;
  assign n14539 = \pi0153  & \pi0160  ;
  assign n14540 = ~n10904 & ~n10983 ;
  assign n14541 = n10900 & ~n10983 ;
  assign n14542 = ~n10892 & n14541 ;
  assign n14543 = ~n14540 & ~n14542 ;
  assign n14544 = n14539 & ~n14543 ;
  assign n14545 = ~n14538 & n14544 ;
  assign n14546 = ~n10901 & n10904 ;
  assign n14547 = ~\pi0160  & n11009 ;
  assign n14548 = ~\pi0160  & n11010 ;
  assign n14549 = ~n10892 & n14548 ;
  assign n14550 = ~n14547 & ~n14549 ;
  assign n14551 = ~n14546 & ~n14550 ;
  assign n14552 = \pi0160  & n10983 ;
  assign n14553 = ~\pi0153  & ~n14552 ;
  assign n14554 = n11009 & n14553 ;
  assign n14555 = n11010 & n14553 ;
  assign n14556 = ~n10892 & n14555 ;
  assign n14557 = ~n14554 & ~n14556 ;
  assign n14558 = \pi0153  & n10414 ;
  assign n14559 = n1618 & n14558 ;
  assign n14560 = ~n10899 & n14559 ;
  assign n14561 = n1264 & n11984 ;
  assign n14562 = n10937 & n14561 ;
  assign n14563 = n10319 & n14562 ;
  assign n14564 = ~\pi0040  & ~\pi0163  ;
  assign n14565 = ~n14563 & n14564 ;
  assign n14566 = ~n14552 & n14565 ;
  assign n14567 = ~n14560 & n14566 ;
  assign n14568 = ~n11984 & ~n14552 ;
  assign n14569 = ~n14567 & ~n14568 ;
  assign n14570 = n14557 & n14569 ;
  assign n14571 = ~n14551 & n14570 ;
  assign n14572 = ~n14545 & n14571 ;
  assign n14573 = ~\pi0040  & \pi0163  ;
  assign n14574 = ~n14567 & ~n14573 ;
  assign n14575 = ~n10952 & n11010 ;
  assign n14576 = ~n11009 & ~n14575 ;
  assign n14577 = \pi0153  & n10903 ;
  assign n14578 = ~n1864 & n14577 ;
  assign n14579 = ~n11015 & n14578 ;
  assign n14580 = ~n14576 & ~n14579 ;
  assign n14581 = n14139 & ~n14567 ;
  assign n14582 = ~n14580 & n14581 ;
  assign n14583 = ~n14574 & ~n14582 ;
  assign n14584 = \pi0299  & n14583 ;
  assign n14585 = ~n14572 & n14584 ;
  assign n14586 = n6706 & n14266 ;
  assign n14587 = ~\pi0035  & \pi0182  ;
  assign n14588 = n1979 & n14587 ;
  assign n14589 = n1354 & n14588 ;
  assign n14590 = n1358 & n14589 ;
  assign n14591 = \pi0184  & \pi0189  ;
  assign n14592 = n10942 & ~n10952 ;
  assign n14593 = ~n10944 & ~n14592 ;
  assign n14594 = n14591 & n14593 ;
  assign n14595 = ~n14590 & ~n14594 ;
  assign n14596 = \pi0184  & n10944 ;
  assign n14597 = \pi0184  & n10942 ;
  assign n14598 = ~n10892 & n14597 ;
  assign n14599 = ~n14596 & ~n14598 ;
  assign n14600 = \pi0184  & ~\pi0189  ;
  assign n14601 = ~\pi0189  & n1264 ;
  assign n14602 = n10937 & n14601 ;
  assign n14603 = n10319 & n14602 ;
  assign n14604 = ~n14600 & ~n14603 ;
  assign n14605 = n14599 & ~n14604 ;
  assign n14606 = n14595 & ~n14605 ;
  assign n14607 = n14586 & ~n14606 ;
  assign n14608 = n14585 & ~n14607 ;
  assign n14609 = \pi0175  & n6706 ;
  assign n14610 = n14590 & n14609 ;
  assign n14611 = ~\pi0189  & n10904 ;
  assign n14612 = ~n10901 & n14611 ;
  assign n14613 = n2265 & ~n10914 ;
  assign n14614 = ~n10913 & n14613 ;
  assign n14615 = ~n14612 & ~n14614 ;
  assign n14616 = \pi0189  & n10955 ;
  assign n14617 = \pi0184  & ~n14616 ;
  assign n14618 = n14615 & n14617 ;
  assign n14619 = ~n10929 & n14601 ;
  assign n14620 = n10923 & n14619 ;
  assign n14621 = \pi0189  & n1264 ;
  assign n14622 = n1618 & n14621 ;
  assign n14623 = ~n10899 & n14622 ;
  assign n14624 = ~\pi0184  & ~n14623 ;
  assign n14625 = ~n14620 & n14624 ;
  assign n14626 = n14609 & ~n14625 ;
  assign n14627 = ~n14618 & n14626 ;
  assign n14628 = ~n14610 & ~n14627 ;
  assign n14629 = n14517 & ~n14607 ;
  assign n14630 = n14628 & n14629 ;
  assign n14631 = ~n14608 & ~n14630 ;
  assign n14632 = ~\pi0039  & n14535 ;
  assign n14633 = n14631 & n14632 ;
  assign n14634 = ~n14536 & ~n14633 ;
  assign n14635 = n14448 & ~n14499 ;
  assign n14636 = n14634 & n14635 ;
  assign n14637 = ~n14500 & ~n14636 ;
  assign n14638 = ~\pi0035  & n1264 ;
  assign n14639 = n1618 & n14638 ;
  assign n14640 = n14459 & n14639 ;
  assign n14641 = n2341 & n14640 ;
  assign n14642 = n1354 & n14641 ;
  assign n14643 = n1358 & n14642 ;
  assign n14644 = ~\pi0038  & ~\pi0040  ;
  assign n14645 = ~n14643 & n14644 ;
  assign n14646 = n6895 & ~n14118 ;
  assign n14647 = ~\pi0100  & n14646 ;
  assign n14648 = ~n14645 & n14647 ;
  assign n14649 = \pi0299  & ~n14030 ;
  assign n14650 = n14109 & ~n14649 ;
  assign n14651 = ~n2364 & ~n8601 ;
  assign n14652 = ~n14650 & n14651 ;
  assign n14653 = ~n14648 & ~n14652 ;
  assign n14654 = n14113 & n14653 ;
  assign n14655 = ~n14637 & n14654 ;
  assign n14656 = ~n2364 & n14653 ;
  assign n14657 = n2511 & ~n14656 ;
  assign n14658 = ~n14655 & n14657 ;
  assign n14659 = n2467 & ~n14047 ;
  assign n14660 = ~\pi0074  & ~n14483 ;
  assign n14661 = n14063 & ~n14660 ;
  assign n14662 = n14659 & n14661 ;
  assign n14663 = ~n14658 & n14662 ;
  assign n14664 = n8601 & ~n14021 ;
  assign n14665 = ~\pi0092  & n14079 ;
  assign n14666 = n11407 & n14665 ;
  assign n14667 = n1354 & n14666 ;
  assign n14668 = n14501 & n14667 ;
  assign n14669 = n1358 & n14668 ;
  assign n14670 = n10155 & ~n14669 ;
  assign n14671 = n14664 & ~n14670 ;
  assign n14672 = n8601 & ~n14039 ;
  assign n14673 = ~n14037 & ~n14672 ;
  assign n14674 = ~n14671 & ~n14673 ;
  assign n14675 = n14105 & ~n14674 ;
  assign n14676 = ~n14068 & ~n14675 ;
  assign n14677 = n14659 & n14676 ;
  assign n14678 = \pi0079  & ~n14493 ;
  assign n14679 = ~n14491 & n14678 ;
  assign n14680 = ~n14677 & n14679 ;
  assign n14681 = ~n14663 & n14680 ;
  assign n14682 = ~n14497 & ~n14681 ;
  assign n14683 = ~n14496 & n14682 ;
  assign n14684 = ~\pi0118  & n11101 ;
  assign n14685 = ~\pi0079  & ~n14684 ;
  assign n14686 = n14494 & ~n14685 ;
  assign n14687 = ~n14489 & n14686 ;
  assign n14688 = n14494 & n14685 ;
  assign n14689 = ~n14677 & n14688 ;
  assign n14690 = ~n14663 & n14689 ;
  assign n14691 = n14497 & ~n14690 ;
  assign n14692 = ~n14687 & n14691 ;
  assign n14693 = ~n14683 & ~n14692 ;
  assign n14694 = ~\pi0088  & n1252 ;
  assign n14695 = n13115 & n14694 ;
  assign n14696 = n1542 & n14695 ;
  assign n14697 = \pi0090  & \pi0093  ;
  assign n14698 = ~\pi0841  & ~n1320 ;
  assign n14699 = ~n14697 & n14698 ;
  assign n14700 = n6967 & n14699 ;
  assign n14701 = ~n1322 & ~n14700 ;
  assign n14702 = ~\pi0051  & ~n14698 ;
  assign n14703 = ~\pi0051  & ~n1321 ;
  assign n14704 = ~\pi0051  & n14697 ;
  assign n14705 = ~n14703 & ~n14704 ;
  assign n14706 = ~n14702 & n14705 ;
  assign n14707 = \pi0824  & \pi0950  ;
  assign n14708 = n1264 & n14707 ;
  assign n14709 = n1263 & n14708 ;
  assign n14710 = n14706 & n14709 ;
  assign n14711 = ~n14701 & n14710 ;
  assign n14712 = n14696 & n14711 ;
  assign n14713 = ~\pi0098  & ~n14712 ;
  assign n14714 = ~\pi0098  & ~n9112 ;
  assign n14715 = n9103 & n14714 ;
  assign n14716 = ~\pi0098  & n9112 ;
  assign n14717 = ~n9103 & n14716 ;
  assign n14718 = ~n14715 & ~n14717 ;
  assign n14719 = \pi1092  & n14718 ;
  assign n14720 = ~n14713 & n14719 ;
  assign n14721 = \pi0098  & \pi1092  ;
  assign n14722 = \pi1092  & n14709 ;
  assign n14723 = n14706 & n14722 ;
  assign n14724 = ~n14701 & n14723 ;
  assign n14725 = n14696 & n14724 ;
  assign n14726 = ~n14721 & ~n14725 ;
  assign n14727 = \pi1092  & \pi1093  ;
  assign n14728 = \pi0098  & \pi1091  ;
  assign n14729 = n14727 & n14728 ;
  assign n14730 = ~n8543 & ~n14729 ;
  assign n14731 = n2342 & ~n14730 ;
  assign n14732 = ~n14726 & n14731 ;
  assign n14733 = n14720 & n14732 ;
  assign n14734 = \pi1093  & n14721 ;
  assign n14735 = ~n2328 & n14734 ;
  assign n14736 = ~n14733 & ~n14735 ;
  assign n14737 = n1322 & n13028 ;
  assign n14738 = n13115 & n14737 ;
  assign n14739 = n1542 & n14738 ;
  assign n14740 = ~\pi0040  & \pi1092  ;
  assign n14741 = n1262 & n14740 ;
  assign n14742 = n10902 & n14741 ;
  assign n14743 = n14707 & n14742 ;
  assign n14744 = n14739 & n14743 ;
  assign n14745 = ~n14721 & ~n14744 ;
  assign n14746 = n9115 & ~n14745 ;
  assign n14747 = ~n9112 & n14721 ;
  assign n14748 = n9103 & n14747 ;
  assign n14749 = n9112 & n14721 ;
  assign n14750 = ~n9103 & n14749 ;
  assign n14751 = ~n14748 & ~n14750 ;
  assign n14752 = ~n14746 & n14751 ;
  assign n14753 = n8813 & ~n14730 ;
  assign n14754 = n14721 & n14753 ;
  assign n14755 = n14743 & n14753 ;
  assign n14756 = n14739 & n14755 ;
  assign n14757 = ~n14754 & ~n14756 ;
  assign n14758 = ~n14752 & ~n14757 ;
  assign n14759 = n14736 & ~n14758 ;
  assign n14760 = ~\pi0098  & \pi0567  ;
  assign n14761 = n14727 & ~n14760 ;
  assign n14762 = ~n8496 & ~n14761 ;
  assign n14763 = n9603 & ~n14762 ;
  assign n14764 = n9520 & n14763 ;
  assign n14765 = ~n14759 & n14764 ;
  assign n14766 = n14729 & n14731 ;
  assign n14767 = n9083 & n14726 ;
  assign n14768 = ~n9070 & ~n14721 ;
  assign n14769 = n9061 & n14768 ;
  assign n14770 = n9070 & ~n14721 ;
  assign n14771 = ~n9061 & n14770 ;
  assign n14772 = ~n14769 & ~n14771 ;
  assign n14773 = n14731 & n14772 ;
  assign n14774 = ~n14767 & n14773 ;
  assign n14775 = ~n14766 & ~n14774 ;
  assign n14776 = ~n9070 & ~n14729 ;
  assign n14777 = ~n9061 & n14776 ;
  assign n14778 = n9070 & ~n14729 ;
  assign n14779 = n9061 & n14778 ;
  assign n14780 = ~n14777 & ~n14779 ;
  assign n14781 = n14745 & ~n14780 ;
  assign n14782 = ~n14721 & ~n14729 ;
  assign n14783 = ~n9070 & n14782 ;
  assign n14784 = n9061 & n14783 ;
  assign n14785 = n9070 & n14782 ;
  assign n14786 = ~n9061 & n14785 ;
  assign n14787 = ~n14784 & ~n14786 ;
  assign n14788 = n14753 & n14787 ;
  assign n14789 = ~n14781 & n14788 ;
  assign n14790 = n9115 & ~n14757 ;
  assign n14791 = ~n14789 & ~n14790 ;
  assign n14792 = n14775 & n14791 ;
  assign n14793 = n14736 & n14792 ;
  assign n14794 = n9540 & ~n14762 ;
  assign n14795 = n9520 & n14794 ;
  assign n14796 = ~n14793 & n14795 ;
  assign n14797 = ~n14765 & ~n14796 ;
  assign n14798 = \pi1199  & ~n14761 ;
  assign n14799 = ~\pi0567  & n1689 ;
  assign n14800 = n8496 & ~n14799 ;
  assign n14801 = n9124 & n14800 ;
  assign n14802 = ~n14798 & ~n14801 ;
  assign n14803 = n14797 & ~n14802 ;
  assign n14804 = n9226 & ~n14803 ;
  assign n14805 = ~\pi0591  & ~n14761 ;
  assign n14806 = ~n9794 & ~n14805 ;
  assign n14807 = ~\pi0567  & n14800 ;
  assign n14808 = ~\pi0075  & ~n14757 ;
  assign n14809 = ~\pi0075  & n2342 ;
  assign n14810 = ~n14730 & n14809 ;
  assign n14811 = ~n14726 & n14810 ;
  assign n14812 = ~n14808 & ~n14811 ;
  assign n14813 = ~n8602 & n14734 ;
  assign n14814 = n14800 & ~n14813 ;
  assign n14815 = n14812 & n14814 ;
  assign n14816 = ~n14807 & ~n14815 ;
  assign n14817 = \pi0592  & ~n14762 ;
  assign n14818 = ~n9385 & n14817 ;
  assign n14819 = n14816 & n14818 ;
  assign n14820 = ~n14806 & ~n14819 ;
  assign n14821 = ~n9540 & n14761 ;
  assign n14822 = ~\pi1199  & ~n14821 ;
  assign n14823 = n14794 & ~n14800 ;
  assign n14824 = \pi0075  & ~n14813 ;
  assign n14825 = ~n14789 & ~n14813 ;
  assign n14826 = n14775 & n14825 ;
  assign n14827 = ~n14824 & ~n14826 ;
  assign n14828 = \pi0567  & n14794 ;
  assign n14829 = n14827 & n14828 ;
  assign n14830 = ~n14823 & ~n14829 ;
  assign n14831 = n14822 & n14830 ;
  assign n14832 = ~n14820 & ~n14831 ;
  assign n14833 = n14804 & n14832 ;
  assign n14834 = \pi0592  & n14761 ;
  assign n14835 = \pi0591  & ~n14834 ;
  assign n14836 = ~n9235 & ~n14835 ;
  assign n14837 = ~\pi0592  & ~n14762 ;
  assign n14838 = ~n9235 & n14837 ;
  assign n14839 = n14816 & n14838 ;
  assign n14840 = ~n14836 & ~n14839 ;
  assign n14841 = ~n14820 & ~n14840 ;
  assign n14842 = ~\pi0590  & ~n14841 ;
  assign n14843 = ~n14833 & n14842 ;
  assign n14844 = ~\pi0588  & ~n14843 ;
  assign n14845 = \pi0588  & ~n9927 ;
  assign n14846 = n14761 & n14845 ;
  assign n14847 = n14816 & n14837 ;
  assign n14848 = ~n9987 & ~n14834 ;
  assign n14849 = ~n14847 & n14848 ;
  assign n14850 = ~n9927 & ~n14761 ;
  assign n14851 = \pi0588  & ~n14850 ;
  assign n14852 = ~n9980 & ~n14761 ;
  assign n14853 = n9889 & n14852 ;
  assign n14854 = n14851 & ~n14853 ;
  assign n14855 = ~n14849 & n14854 ;
  assign n14856 = ~n14846 & ~n14855 ;
  assign n14857 = ~n14844 & n14856 ;
  assign n14858 = n8862 & ~n14834 ;
  assign n14859 = ~n14847 & n14858 ;
  assign n14860 = ~n8830 & ~n14859 ;
  assign n14861 = n8830 & n14834 ;
  assign n14862 = n8830 & n14837 ;
  assign n14863 = n14816 & n14862 ;
  assign n14864 = ~n14861 & ~n14863 ;
  assign n14865 = ~n14860 & n14864 ;
  assign n14866 = ~\pi0455  & n14761 ;
  assign n14867 = ~n14834 & ~n14866 ;
  assign n14868 = ~n14847 & n14867 ;
  assign n14869 = ~\pi0455  & ~n14761 ;
  assign n14870 = ~n14868 & ~n14869 ;
  assign n14871 = \pi0355  & \pi0452  ;
  assign n14872 = ~n14870 & n14871 ;
  assign n14873 = \pi0455  & n14761 ;
  assign n14874 = ~n14834 & ~n14873 ;
  assign n14875 = ~n14847 & n14874 ;
  assign n14876 = \pi0455  & ~n14761 ;
  assign n14877 = ~n14875 & ~n14876 ;
  assign n14878 = \pi0355  & ~\pi0452  ;
  assign n14879 = ~n14877 & n14878 ;
  assign n14880 = ~n14872 & ~n14879 ;
  assign n14881 = \pi0355  & \pi0458  ;
  assign n14882 = ~n8877 & ~n14834 ;
  assign n14883 = ~n14847 & n14882 ;
  assign n14884 = n8877 & ~n14761 ;
  assign n14885 = \pi0458  & ~n14884 ;
  assign n14886 = ~n14883 & n14885 ;
  assign n14887 = ~n14881 & ~n14886 ;
  assign n14888 = n14880 & ~n14887 ;
  assign n14889 = ~n8868 & ~n8871 ;
  assign n14890 = n8868 & n8871 ;
  assign n14891 = ~n14889 & ~n14890 ;
  assign n14892 = ~\pi0355  & \pi0452  ;
  assign n14893 = ~n14870 & n14892 ;
  assign n14894 = ~\pi0355  & ~\pi0452  ;
  assign n14895 = ~n14877 & n14894 ;
  assign n14896 = ~n14893 & ~n14895 ;
  assign n14897 = ~\pi0355  & ~\pi0458  ;
  assign n14898 = ~\pi0458  & ~n14884 ;
  assign n14899 = ~n14883 & n14898 ;
  assign n14900 = ~n14897 & ~n14899 ;
  assign n14901 = n14896 & ~n14900 ;
  assign n14902 = ~n14891 & ~n14901 ;
  assign n14903 = ~n14888 & n14902 ;
  assign n14904 = \pi1196  & ~n14903 ;
  assign n14905 = n8932 & ~n14761 ;
  assign n14906 = ~n8923 & n14905 ;
  assign n14907 = ~n8932 & ~n14761 ;
  assign n14908 = n8923 & n14907 ;
  assign n14909 = ~n14906 & ~n14908 ;
  assign n14910 = ~n8905 & ~n14909 ;
  assign n14911 = ~n9736 & ~n14834 ;
  assign n14912 = ~n14847 & n14911 ;
  assign n14913 = ~n14910 & ~n14912 ;
  assign n14914 = \pi1198  & ~n14913 ;
  assign n14915 = ~n8873 & ~n14886 ;
  assign n14916 = n14896 & ~n14915 ;
  assign n14917 = \pi0355  & ~\pi0458  ;
  assign n14918 = ~n14899 & ~n14917 ;
  assign n14919 = n14880 & ~n14918 ;
  assign n14920 = n14891 & ~n14919 ;
  assign n14921 = ~n14916 & n14920 ;
  assign n14922 = ~n14914 & ~n14921 ;
  assign n14923 = n14904 & n14922 ;
  assign n14924 = ~\pi1196  & n14761 ;
  assign n14925 = ~\pi1198  & ~n14924 ;
  assign n14926 = ~\pi1198  & ~n14925 ;
  assign n14927 = ~n14910 & ~n14925 ;
  assign n14928 = ~n14912 & n14927 ;
  assign n14929 = ~n14926 & ~n14928 ;
  assign n14930 = ~n8862 & n14929 ;
  assign n14931 = n14864 & n14930 ;
  assign n14932 = ~n14923 & n14931 ;
  assign n14933 = ~n14865 & ~n14932 ;
  assign n14934 = ~n9414 & ~n14933 ;
  assign n14935 = ~\pi0351  & \pi1199  ;
  assign n14936 = ~n14859 & ~n14935 ;
  assign n14937 = n14834 & n14935 ;
  assign n14938 = n14837 & n14935 ;
  assign n14939 = n14816 & n14938 ;
  assign n14940 = ~n14937 & ~n14939 ;
  assign n14941 = n9414 & n14940 ;
  assign n14942 = ~n14936 & n14941 ;
  assign n14943 = n14930 & n14941 ;
  assign n14944 = ~n14923 & n14943 ;
  assign n14945 = ~n14942 & ~n14944 ;
  assign n14946 = ~\pi0591  & n14945 ;
  assign n14947 = ~n14934 & n14946 ;
  assign n14948 = \pi0591  & n14761 ;
  assign n14949 = \pi0590  & ~n14948 ;
  assign n14950 = n14856 & n14949 ;
  assign n14951 = ~n14947 & n14950 ;
  assign n14952 = ~n14857 & ~n14951 ;
  assign n14953 = n9250 & ~n14952 ;
  assign n14954 = n2342 & ~n14729 ;
  assign n14955 = ~n14720 & n14954 ;
  assign n14956 = \pi0411  & \pi0412  ;
  assign n14957 = ~n9067 & n14956 ;
  assign n14958 = n9062 & n9067 ;
  assign n14959 = ~n14957 & ~n14958 ;
  assign n14960 = ~n9061 & ~n14959 ;
  assign n14961 = n9062 & ~n9067 ;
  assign n14962 = n9067 & n14956 ;
  assign n14963 = ~n14961 & ~n14962 ;
  assign n14964 = n9061 & ~n14963 ;
  assign n14965 = ~n14960 & ~n14964 ;
  assign n14966 = n14772 & n14965 ;
  assign n14967 = ~n14767 & n14966 ;
  assign n14968 = n14955 & ~n14967 ;
  assign n14969 = ~\pi0122  & n14721 ;
  assign n14970 = ~\pi0122  & \pi0824  ;
  assign n14971 = n6809 & n14970 ;
  assign n14972 = ~n14969 & ~n14971 ;
  assign n14973 = ~n14721 & n14972 ;
  assign n14974 = ~n14769 & ~n14973 ;
  assign n14975 = ~n14771 & n14974 ;
  assign n14976 = n8543 & n14975 ;
  assign n14977 = n9012 & n9112 ;
  assign n14978 = ~\pi0122  & ~n14721 ;
  assign n14979 = ~n14977 & n14978 ;
  assign n14980 = n9103 & n14979 ;
  assign n14981 = n9012 & ~n9112 ;
  assign n14982 = n14978 & ~n14981 ;
  assign n14983 = ~n9103 & n14982 ;
  assign n14984 = ~n14980 & ~n14983 ;
  assign n14985 = ~n14730 & n14984 ;
  assign n14986 = n2328 & ~n14985 ;
  assign n14987 = ~n14976 & n14986 ;
  assign n14988 = ~n14781 & n14787 ;
  assign n14989 = n8813 & ~n14746 ;
  assign n14990 = ~n14988 & n14989 ;
  assign n14991 = ~n14987 & ~n14990 ;
  assign n14992 = ~n14968 & n14991 ;
  assign n14993 = n14772 & ~n14972 ;
  assign n14994 = n9112 & n14971 ;
  assign n14995 = n9103 & n14994 ;
  assign n14996 = ~n9112 & n14971 ;
  assign n14997 = ~n9103 & n14996 ;
  assign n14998 = ~n14995 & ~n14997 ;
  assign n14999 = ~n14993 & n14998 ;
  assign n15000 = ~n14987 & ~n14999 ;
  assign n15001 = n14799 & ~n14800 ;
  assign n15002 = ~n8695 & ~n14721 ;
  assign n15003 = \pi0567  & ~n14730 ;
  assign n15004 = ~n15002 & n15003 ;
  assign n15005 = ~n14800 & n15004 ;
  assign n15006 = n14984 & n15005 ;
  assign n15007 = ~n15001 & ~n15006 ;
  assign n15008 = \pi0567  & ~n8496 ;
  assign n15009 = ~n14730 & n15008 ;
  assign n15010 = n14975 & n15009 ;
  assign n15011 = n15007 & ~n15010 ;
  assign n15012 = ~\pi0075  & n15011 ;
  assign n15013 = ~n15000 & n15012 ;
  assign n15014 = ~n14992 & n15013 ;
  assign n15015 = n9540 & ~n15011 ;
  assign n15016 = ~n14730 & ~n15002 ;
  assign n15017 = n14984 & n15016 ;
  assign n15018 = ~n8602 & ~n15017 ;
  assign n15019 = ~n14976 & n15018 ;
  assign n15020 = ~\pi0092  & \pi0567  ;
  assign n15021 = n2511 & n15020 ;
  assign n15022 = n9540 & n15021 ;
  assign n15023 = ~n15019 & n15022 ;
  assign n15024 = ~n15015 & ~n15023 ;
  assign n15025 = ~n15014 & ~n15024 ;
  assign n15026 = \pi1199  & ~n9603 ;
  assign n15027 = n8602 & n15021 ;
  assign n15028 = n15016 & n15021 ;
  assign n15029 = n14984 & n15028 ;
  assign n15030 = ~n15027 & ~n15029 ;
  assign n15031 = \pi1199  & n15007 ;
  assign n15032 = n15030 & n15031 ;
  assign n15033 = \pi0122  & n14954 ;
  assign n15034 = ~n14720 & n15033 ;
  assign n15035 = n8813 & ~n14729 ;
  assign n15036 = \pi0122  & n15035 ;
  assign n15037 = n14751 & n15036 ;
  assign n15038 = ~n14746 & n15037 ;
  assign n15039 = ~n14986 & ~n15038 ;
  assign n15040 = ~n15034 & n15039 ;
  assign n15041 = ~\pi0075  & n15031 ;
  assign n15042 = ~n15040 & n15041 ;
  assign n15043 = ~n15032 & ~n15042 ;
  assign n15044 = ~n15026 & n15043 ;
  assign n15045 = ~n15025 & ~n15044 ;
  assign n15046 = n8813 & ~n14988 ;
  assign n15047 = ~n14767 & n14772 ;
  assign n15048 = n14954 & ~n15047 ;
  assign n15049 = ~n15046 & ~n15048 ;
  assign n15050 = ~\pi0075  & ~n14993 ;
  assign n15051 = ~n15049 & n15050 ;
  assign n15052 = ~n9012 & ~n14721 ;
  assign n15053 = ~n14730 & ~n15052 ;
  assign n15054 = n14772 & n15053 ;
  assign n15055 = \pi0122  & ~n14730 ;
  assign n15056 = n2328 & ~n15055 ;
  assign n15057 = ~\pi0075  & n15056 ;
  assign n15058 = ~n15054 & n15057 ;
  assign n15059 = ~n14730 & n15021 ;
  assign n15060 = n14975 & n15059 ;
  assign n15061 = ~n15027 & ~n15060 ;
  assign n15062 = n9540 & ~n15061 ;
  assign n15063 = ~n15058 & n15062 ;
  assign n15064 = ~n15051 & n15063 ;
  assign n15065 = ~\pi1199  & ~n14924 ;
  assign n15066 = ~n9540 & n15065 ;
  assign n15067 = ~n14799 & n15065 ;
  assign n15068 = ~n15010 & n15067 ;
  assign n15069 = ~n15066 & ~n15068 ;
  assign n15070 = ~n15064 & ~n15069 ;
  assign n15071 = n9226 & ~n15070 ;
  assign n15072 = ~n15045 & n15071 ;
  assign n15073 = ~n8602 & ~n14734 ;
  assign n15074 = ~n8696 & n15073 ;
  assign n15075 = n15021 & ~n15074 ;
  assign n15076 = ~\pi0075  & ~n14729 ;
  assign n15077 = n15075 & ~n15076 ;
  assign n15078 = \pi0122  & ~n14721 ;
  assign n15079 = n8813 & n15078 ;
  assign n15080 = ~n14744 & n15079 ;
  assign n15081 = \pi0122  & n2342 ;
  assign n15082 = ~n14721 & n15081 ;
  assign n15083 = ~n14725 & n15082 ;
  assign n15084 = ~n15080 & ~n15083 ;
  assign n15085 = n2328 & ~n8543 ;
  assign n15086 = ~\pi0122  & ~n14734 ;
  assign n15087 = n2328 & ~n8695 ;
  assign n15088 = n15086 & n15087 ;
  assign n15089 = ~n15085 & ~n15088 ;
  assign n15090 = n15075 & n15089 ;
  assign n15091 = n15084 & n15090 ;
  assign n15092 = ~n15077 & ~n15091 ;
  assign n15093 = ~n14734 & ~n14799 ;
  assign n15094 = ~n8696 & n15093 ;
  assign n15095 = ~n14800 & ~n15094 ;
  assign n15096 = n15092 & ~n15095 ;
  assign n15097 = ~\pi0592  & ~n9226 ;
  assign n15098 = ~n15096 & n15097 ;
  assign n15099 = ~\pi0590  & n14835 ;
  assign n15100 = ~n15098 & n15099 ;
  assign n15101 = ~n15072 & n15100 ;
  assign n15102 = n9385 & n14805 ;
  assign n15103 = ~\pi0592  & n14805 ;
  assign n15104 = ~n15102 & ~n15103 ;
  assign n15105 = ~\pi0590  & ~n15104 ;
  assign n15106 = n14805 & ~n15095 ;
  assign n15107 = n9793 & ~n15095 ;
  assign n15108 = ~n9385 & n15107 ;
  assign n15109 = ~n15106 & ~n15108 ;
  assign n15110 = ~\pi0590  & n15092 ;
  assign n15111 = ~n15109 & n15110 ;
  assign n15112 = ~n15105 & ~n15111 ;
  assign n15113 = ~\pi0588  & n15112 ;
  assign n15114 = ~n15101 & n15113 ;
  assign n15115 = ~n14949 & n15114 ;
  assign n15116 = ~n8830 & ~n8862 ;
  assign n15117 = ~n14834 & ~n15095 ;
  assign n15118 = n15092 & n15117 ;
  assign n15119 = \pi0592  & ~n14761 ;
  assign n15120 = ~n8830 & ~n15119 ;
  assign n15121 = ~n15118 & n15120 ;
  assign n15122 = ~n15116 & ~n15121 ;
  assign n15123 = n8830 & ~n15119 ;
  assign n15124 = ~n15118 & n15123 ;
  assign n15125 = ~n9414 & ~n15124 ;
  assign n15126 = n15122 & n15125 ;
  assign n15127 = \pi1198  & ~n14909 ;
  assign n15128 = ~n8905 & n15127 ;
  assign n15129 = \pi1198  & n9735 ;
  assign n15130 = \pi1196  & \pi1198  ;
  assign n15131 = n8904 & n15130 ;
  assign n15132 = ~n15129 & ~n15131 ;
  assign n15133 = ~n15128 & n15132 ;
  assign n15134 = ~n15119 & ~n15128 ;
  assign n15135 = ~n15118 & n15134 ;
  assign n15136 = ~n15133 & ~n15135 ;
  assign n15137 = ~n14925 & ~n15136 ;
  assign n15138 = ~\pi0452  & ~\pi0455  ;
  assign n15139 = ~n15119 & n15138 ;
  assign n15140 = ~n15118 & n15139 ;
  assign n15141 = ~\pi0452  & \pi0455  ;
  assign n15142 = n14761 & n15141 ;
  assign n15143 = \pi0452  & ~\pi0455  ;
  assign n15144 = n14761 & n15143 ;
  assign n15145 = ~n15142 & ~n15144 ;
  assign n15146 = ~n15140 & n15145 ;
  assign n15147 = \pi0452  & \pi0455  ;
  assign n15148 = ~n15119 & n15147 ;
  assign n15149 = ~n15118 & n15148 ;
  assign n15150 = \pi0355  & ~n15149 ;
  assign n15151 = n15146 & n15150 ;
  assign n15152 = ~\pi0355  & n14884 ;
  assign n15153 = ~\pi0355  & ~n8877 ;
  assign n15154 = ~n15152 & ~n15153 ;
  assign n15155 = ~n15119 & ~n15152 ;
  assign n15156 = ~n15118 & n15155 ;
  assign n15157 = ~n15154 & ~n15156 ;
  assign n15158 = ~\pi0458  & ~n15157 ;
  assign n15159 = ~n15151 & n15158 ;
  assign n15160 = ~\pi0355  & ~n15149 ;
  assign n15161 = n15146 & n15160 ;
  assign n15162 = \pi0355  & n14884 ;
  assign n15163 = \pi0355  & ~n8877 ;
  assign n15164 = ~n15162 & ~n15163 ;
  assign n15165 = ~n15119 & ~n15162 ;
  assign n15166 = ~n15118 & n15165 ;
  assign n15167 = ~n15164 & ~n15166 ;
  assign n15168 = \pi0458  & ~n15167 ;
  assign n15169 = ~n15161 & n15168 ;
  assign n15170 = n14891 & ~n15169 ;
  assign n15171 = ~n15159 & n15170 ;
  assign n15172 = \pi1196  & ~n15171 ;
  assign n15173 = ~\pi0458  & ~n15167 ;
  assign n15174 = ~n15161 & n15173 ;
  assign n15175 = \pi0458  & ~n15157 ;
  assign n15176 = ~n15151 & n15175 ;
  assign n15177 = ~n14891 & ~n15176 ;
  assign n15178 = ~n15174 & n15177 ;
  assign n15179 = ~n15136 & ~n15178 ;
  assign n15180 = n15172 & n15179 ;
  assign n15181 = ~n15137 & ~n15180 ;
  assign n15182 = ~n8854 & ~n8861 ;
  assign n15183 = n15125 & ~n15182 ;
  assign n15184 = n15181 & n15183 ;
  assign n15185 = ~n15126 & ~n15184 ;
  assign n15186 = ~\pi0591  & n15185 ;
  assign n15187 = ~n8862 & ~n8952 ;
  assign n15188 = ~n8952 & ~n15119 ;
  assign n15189 = ~n15118 & n15188 ;
  assign n15190 = ~n15187 & ~n15189 ;
  assign n15191 = n14935 & ~n15119 ;
  assign n15192 = ~n15118 & n15191 ;
  assign n15193 = n9414 & ~n15192 ;
  assign n15194 = n15190 & n15193 ;
  assign n15195 = ~n15182 & n15193 ;
  assign n15196 = n15181 & n15195 ;
  assign n15197 = ~n15194 & ~n15196 ;
  assign n15198 = n15114 & n15197 ;
  assign n15199 = n15186 & n15198 ;
  assign n15200 = ~n15115 & ~n15199 ;
  assign n15201 = n9927 & ~n14761 ;
  assign n15202 = ~n9980 & n15201 ;
  assign n15203 = n9889 & n15202 ;
  assign n15204 = n14851 & ~n15203 ;
  assign n15205 = ~n9250 & ~n15204 ;
  assign n15206 = ~n15118 & ~n15119 ;
  assign n15207 = n9927 & ~n9987 ;
  assign n15208 = ~n9250 & n15207 ;
  assign n15209 = ~n15206 & n15208 ;
  assign n15210 = ~n15205 & ~n15209 ;
  assign n15211 = n15200 & ~n15210 ;
  assign n15212 = ~\pi0057  & ~\pi0080  ;
  assign n15213 = n6848 & n15212 ;
  assign n15214 = ~n15211 & n15213 ;
  assign n15215 = ~n14953 & n15214 ;
  assign n15216 = ~\pi0592  & \pi1199  ;
  assign n15217 = ~n9540 & ~n15216 ;
  assign n15218 = n14761 & n15217 ;
  assign n15219 = n9176 & ~n15218 ;
  assign n15220 = n9225 & n15219 ;
  assign n15221 = \pi0592  & n15220 ;
  assign n15222 = ~\pi0567  & \pi1196  ;
  assign n15223 = n1689 & n15222 ;
  assign n15224 = n9671 & ~n14730 ;
  assign n15225 = n14975 & n15224 ;
  assign n15226 = ~n15223 & ~n15225 ;
  assign n15227 = n14799 & ~n14822 ;
  assign n15228 = ~n14822 & n15004 ;
  assign n15229 = n14984 & n15228 ;
  assign n15230 = ~n15227 & ~n15229 ;
  assign n15231 = n15220 & n15230 ;
  assign n15232 = n15226 & n15231 ;
  assign n15233 = ~n15221 & ~n15232 ;
  assign n15234 = \pi0591  & ~\pi0592  ;
  assign n15235 = n8548 & n15234 ;
  assign n15236 = ~n14948 & ~n15235 ;
  assign n15237 = ~n9235 & n15236 ;
  assign n15238 = n15233 & ~n15237 ;
  assign n15239 = ~\pi0592  & n8548 ;
  assign n15240 = n15201 & ~n15239 ;
  assign n15241 = n14851 & ~n15240 ;
  assign n15242 = ~n9250 & ~n15241 ;
  assign n15243 = ~n9924 & n15201 ;
  assign n15244 = ~n9250 & n15243 ;
  assign n15245 = n9889 & n15244 ;
  assign n15246 = ~n15242 & ~n15245 ;
  assign n15247 = ~\pi0590  & \pi0591  ;
  assign n15248 = ~\pi0590  & ~n14761 ;
  assign n15249 = ~n15247 & ~n15248 ;
  assign n15250 = n9749 & ~n15247 ;
  assign n15251 = ~n9385 & n15250 ;
  assign n15252 = ~n15249 & ~n15251 ;
  assign n15253 = ~n15246 & n15252 ;
  assign n15254 = ~n15238 & n15253 ;
  assign n15255 = n8952 & n9403 ;
  assign n15256 = ~n8968 & n15255 ;
  assign n15257 = n8965 & n15256 ;
  assign n15258 = n8952 & ~n9403 ;
  assign n15259 = ~n8968 & n15258 ;
  assign n15260 = ~n8965 & n15259 ;
  assign n15261 = ~n15257 & ~n15260 ;
  assign n15262 = n8968 & n15258 ;
  assign n15263 = n8965 & n15262 ;
  assign n15264 = n8968 & n15255 ;
  assign n15265 = ~n8965 & n15264 ;
  assign n15266 = ~n15263 & ~n15265 ;
  assign n15267 = n15261 & n15266 ;
  assign n15268 = n8830 & n9403 ;
  assign n15269 = ~n8968 & n15268 ;
  assign n15270 = ~n8965 & n15269 ;
  assign n15271 = n8830 & ~n9403 ;
  assign n15272 = ~n8968 & n15271 ;
  assign n15273 = n8965 & n15272 ;
  assign n15274 = ~n15270 & ~n15273 ;
  assign n15275 = n8830 & n8968 ;
  assign n15276 = ~n9403 & n15275 ;
  assign n15277 = ~n8965 & n15276 ;
  assign n15278 = n9403 & n15275 ;
  assign n15279 = n8965 & n15278 ;
  assign n15280 = ~n15277 & ~n15279 ;
  assign n15281 = n15274 & n15280 ;
  assign n15282 = n15267 & n15281 ;
  assign n15283 = \pi0590  & ~n14761 ;
  assign n15284 = ~n9749 & n15283 ;
  assign n15285 = n15282 & n15284 ;
  assign n15286 = n9744 & n15285 ;
  assign n15287 = ~n9735 & n9737 ;
  assign n15288 = ~n8905 & n15287 ;
  assign n15289 = ~n8862 & n15285 ;
  assign n15290 = n15288 & n15289 ;
  assign n15291 = ~n15286 & ~n15290 ;
  assign n15292 = ~\pi0591  & ~\pi0592  ;
  assign n15293 = n8548 & n15292 ;
  assign n15294 = n15283 & ~n15293 ;
  assign n15295 = ~\pi0588  & ~n15294 ;
  assign n15296 = n15291 & n15295 ;
  assign n15297 = ~n15246 & ~n15296 ;
  assign n15298 = ~\pi0080  & ~n9948 ;
  assign n15299 = n9250 & ~n14761 ;
  assign n15300 = n15298 & ~n15299 ;
  assign n15301 = ~n15297 & n15300 ;
  assign n15302 = ~n15254 & n15301 ;
  assign n15303 = ~\pi0217  & ~n15302 ;
  assign n15304 = ~n15215 & n15303 ;
  assign n15305 = ~\pi0080  & n14761 ;
  assign n15306 = \pi0217  & ~n15305 ;
  assign n15307 = n10003 & ~n15306 ;
  assign n15308 = ~n15304 & n15307 ;
  assign n15309 = ~\pi0314  & n13549 ;
  assign n15310 = \pi0068  & ~\pi0081  ;
  assign n15311 = n1232 & n13022 ;
  assign n15312 = n15310 & n15311 ;
  assign n15313 = n1417 & n13673 ;
  assign n15314 = n15312 & n15313 ;
  assign n15315 = ~n15309 & ~n15314 ;
  assign n15316 = n13149 & n13527 ;
  assign n15317 = ~n15315 & n15316 ;
  assign n15318 = \pi0069  & \pi0314  ;
  assign n15319 = ~\pi0067  & n15318 ;
  assign n15320 = n1236 & n15319 ;
  assign n15321 = n1471 & n15320 ;
  assign n15322 = \pi0066  & ~\pi0073  ;
  assign n15323 = n1233 & n1245 ;
  assign n15324 = n1232 & n15323 ;
  assign n15325 = n15322 & n15324 ;
  assign n15326 = n1242 & n1243 ;
  assign n15327 = n15325 & n15326 ;
  assign n15328 = ~n15321 & ~n15327 ;
  assign n15329 = n13115 & n13152 ;
  assign n15330 = n11824 & n15329 ;
  assign n15331 = ~n15328 & n15330 ;
  assign n15332 = ~\pi0071  & n11803 ;
  assign n15333 = n13089 & n15332 ;
  assign n15334 = n13115 & n15333 ;
  assign n15335 = ~\pi0068  & \pi0084  ;
  assign n15336 = n1245 & n15335 ;
  assign n15337 = n1458 & n15336 ;
  assign n15338 = n1242 & n15337 ;
  assign n15339 = n1232 & n1244 ;
  assign n15340 = n15338 & n15339 ;
  assign n15341 = n15334 & n15340 ;
  assign n15342 = \pi0314  & n15341 ;
  assign n15343 = n1232 & n15338 ;
  assign n15344 = ~\pi0083  & ~n15343 ;
  assign n15345 = ~\pi0103  & n15334 ;
  assign n15346 = ~n15344 & n15345 ;
  assign n15347 = ~\pi0314  & ~n1482 ;
  assign n15348 = n15346 & n15347 ;
  assign n15349 = ~n15342 & ~n15348 ;
  assign n15350 = n11824 & ~n15349 ;
  assign n15351 = ~\pi0299  & n12691 ;
  assign n15352 = \pi0299  & n12577 ;
  assign n15353 = ~n15351 & ~n15352 ;
  assign n15354 = n9948 & ~n15353 ;
  assign n15355 = n1291 & n15354 ;
  assign n15356 = n13549 & n15355 ;
  assign n15357 = n13545 & n15356 ;
  assign n15358 = ~\pi0069  & n13152 ;
  assign n15359 = n6985 & n15358 ;
  assign n15360 = n13149 & n15359 ;
  assign n15361 = ~\pi0069  & ~\pi0314  ;
  assign n15362 = n1424 & n15361 ;
  assign n15363 = n13152 & n15362 ;
  assign n15364 = n1449 & n15363 ;
  assign n15365 = ~n1434 & n15363 ;
  assign n15366 = n1447 & n15365 ;
  assign n15367 = ~n15364 & ~n15366 ;
  assign n15368 = ~\pi0036  & \pi0085  ;
  assign n15369 = n1231 & n15368 ;
  assign n15370 = n1235 & n15369 ;
  assign n15371 = n13149 & n15370 ;
  assign n15372 = ~n15367 & n15371 ;
  assign n15373 = ~n15360 & ~n15372 ;
  assign n15374 = n1696 & ~n6744 ;
  assign n15375 = n1259 & n13578 ;
  assign n15376 = n1249 & n15375 ;
  assign n15377 = n6920 & n15376 ;
  assign n15378 = n15374 & n15377 ;
  assign n15379 = n1696 & n13582 ;
  assign n15380 = ~n6770 & n15379 ;
  assign n15381 = n6921 & n15380 ;
  assign n15382 = ~n15378 & ~n15381 ;
  assign n15383 = n12971 & ~n15382 ;
  assign n15384 = \pi0314  & n15333 ;
  assign n15385 = n1490 & n15384 ;
  assign n15386 = n13149 & n15385 ;
  assign n15387 = ~\pi0088  & ~\pi0109  ;
  assign n15388 = n1252 & n15387 ;
  assign n15389 = n1315 & n15388 ;
  assign n15390 = n13016 & n15389 ;
  assign n15391 = ~\pi0036  & n13023 ;
  assign n15392 = n13020 & n15391 ;
  assign n15393 = n15390 & n15392 ;
  assign n15394 = n1325 & n1326 ;
  assign n15395 = ~n6704 & n15394 ;
  assign n15396 = n1291 & n15395 ;
  assign n15397 = n13003 & n15396 ;
  assign n15398 = n15393 & n15397 ;
  assign n15399 = ~\pi1093  & n1291 ;
  assign n15400 = n9250 & ~n15399 ;
  assign n15401 = ~n15398 & n15400 ;
  assign n15402 = n9035 & ~n13059 ;
  assign n15403 = ~n13052 & n15402 ;
  assign n15404 = ~\pi1093  & n9250 ;
  assign n15405 = ~n15403 & n15404 ;
  assign n15406 = ~n15401 & ~n15405 ;
  assign n15407 = n9250 & n9948 ;
  assign n15408 = n1324 & n9012 ;
  assign n15409 = ~\pi0038  & n1289 ;
  assign n15410 = n1287 & n15409 ;
  assign n15411 = ~\pi0032  & n4520 ;
  assign n15412 = ~\pi1093  & n1329 ;
  assign n15413 = n15411 & n15412 ;
  assign n15414 = n15410 & n15413 ;
  assign n15415 = n9948 & n15414 ;
  assign n15416 = n15408 & n15415 ;
  assign n15417 = ~\pi0098  & n13686 ;
  assign n15418 = n15416 & n15417 ;
  assign n15419 = n1542 & n15418 ;
  assign n15420 = ~n15407 & ~n15419 ;
  assign n15421 = n15406 & ~n15420 ;
  assign n15422 = n10310 & n10311 ;
  assign n15423 = n11844 & n15422 ;
  assign n15424 = \pi0841  & n1322 ;
  assign n15425 = n1255 & n15424 ;
  assign n15426 = n13115 & n15425 ;
  assign n15427 = n15423 & n15426 ;
  assign n15428 = ~\pi0024  & \pi0070  ;
  assign n15429 = ~\pi0035  & n15428 ;
  assign n15430 = n1354 & n15429 ;
  assign n15431 = n1358 & n15430 ;
  assign n15432 = ~n15427 & ~n15431 ;
  assign n15433 = n10903 & n11822 ;
  assign n15434 = ~n15432 & n15433 ;
  assign n15435 = ~\pi0090  & n1256 ;
  assign n15436 = n10327 & n15435 ;
  assign n15437 = n1273 & n15436 ;
  assign n15438 = ~\pi1050  & n15437 ;
  assign n15439 = n10319 & n15438 ;
  assign n15440 = ~\pi0093  & n1321 ;
  assign n15441 = n10903 & n15440 ;
  assign n15442 = n11822 & n15441 ;
  assign n15443 = n15439 & n15442 ;
  assign n15444 = \pi0090  & n15442 ;
  assign n15445 = ~n10920 & n15444 ;
  assign n15446 = ~n15443 & ~n15445 ;
  assign n15447 = ~n1857 & ~n15446 ;
  assign n15448 = ~n1288 & ~n8795 ;
  assign n15449 = ~\pi0058  & n1696 ;
  assign n15450 = n13042 & n15449 ;
  assign n15451 = n11817 & n15450 ;
  assign n15452 = n1319 & n15451 ;
  assign n15453 = \pi0024  & ~\pi0093  ;
  assign n15454 = n1277 & n15453 ;
  assign n15455 = ~n1696 & n15454 ;
  assign n15456 = n11817 & n15455 ;
  assign n15457 = n1319 & n15456 ;
  assign n15458 = n1267 & n15457 ;
  assign n15459 = n1696 & n13042 ;
  assign n15460 = n11815 & n15459 ;
  assign n15461 = ~\pi0039  & ~n15460 ;
  assign n15462 = ~n15458 & n15461 ;
  assign n15463 = ~n15452 & n15462 ;
  assign n15464 = ~n15448 & ~n15463 ;
  assign n15465 = n11834 & n15464 ;
  assign n15466 = n1286 & n13709 ;
  assign n15467 = n2402 & n15466 ;
  assign n15468 = \pi0092  & n15467 ;
  assign n15469 = n1281 & n15468 ;
  assign n15470 = n1260 & n15469 ;
  assign n15471 = n12970 & n15470 ;
  assign n15472 = n7597 & ~n8381 ;
  assign n15473 = ~\pi0223  & n6771 ;
  assign n15474 = ~n8387 & n15473 ;
  assign n15475 = ~n15472 & ~n15474 ;
  assign n15476 = n12968 & ~n15475 ;
  assign n15477 = n8790 & n12970 ;
  assign n15478 = n15476 & n15477 ;
  assign n15479 = ~n15471 & ~n15478 ;
  assign n15480 = ~\pi1050  & n1259 ;
  assign n15481 = n1281 & n15480 ;
  assign n15482 = n1249 & n15481 ;
  assign n15483 = \pi0092  & n15482 ;
  assign n15484 = \pi0093  & n1261 ;
  assign n15485 = n1266 & n15484 ;
  assign n15486 = n1256 & n1277 ;
  assign n15487 = n15485 & n15486 ;
  assign n15488 = n1358 & n15487 ;
  assign n15489 = ~\pi0092  & \pi0841  ;
  assign n15490 = n15488 & n15489 ;
  assign n15491 = ~n15483 & ~n15490 ;
  assign n15492 = n2536 & n12970 ;
  assign n15493 = ~n15491 & n15492 ;
  assign n15494 = ~\pi0841  & n1276 ;
  assign n15495 = n13012 & n15494 ;
  assign n15496 = n13094 & n15495 ;
  assign n15497 = ~n1580 & ~n15496 ;
  assign n15498 = ~n6808 & n13108 ;
  assign n15499 = ~n8641 & n15498 ;
  assign n15500 = n13771 & n15499 ;
  assign n15501 = n1261 & n13413 ;
  assign n15502 = n1266 & n15501 ;
  assign n15503 = n1351 & n15502 ;
  assign n15504 = n13099 & n15503 ;
  assign n15505 = ~n15500 & ~n15504 ;
  assign n15506 = ~n15497 & ~n15505 ;
  assign n15507 = n13099 & n13414 ;
  assign n15508 = \pi0252  & ~n6808 ;
  assign n15509 = ~n8641 & n15508 ;
  assign n15510 = n15507 & ~n15509 ;
  assign n15511 = ~\pi1093  & ~n10050 ;
  assign n15512 = ~n1696 & n15511 ;
  assign n15513 = n13414 & ~n13738 ;
  assign n15514 = n13099 & n15513 ;
  assign n15515 = ~n15512 & ~n15514 ;
  assign n15516 = ~n6808 & n8675 ;
  assign n15517 = ~n8641 & n15516 ;
  assign n15518 = ~n15515 & n15517 ;
  assign n15519 = ~n15510 & ~n15518 ;
  assign n15520 = ~n15506 & n15519 ;
  assign n15521 = n11822 & ~n15520 ;
  assign n15522 = ~n13620 & ~n13627 ;
  assign n15523 = n2214 & ~n13617 ;
  assign n15524 = ~n8387 & n15523 ;
  assign n15525 = ~n15522 & ~n15524 ;
  assign n15526 = n6954 & ~n15525 ;
  assign n15527 = \pi0039  & ~n15526 ;
  assign n15528 = ~\pi0072  & \pi0095  ;
  assign n15529 = n1634 & n15528 ;
  assign n15530 = \pi0024  & n15529 ;
  assign n15531 = n1627 & n15530 ;
  assign n15532 = n1319 & n15531 ;
  assign n15533 = n1255 & n13115 ;
  assign n15534 = n15423 & n15533 ;
  assign n15535 = ~\pi0332  & n1261 ;
  assign n15536 = n13413 & n15535 ;
  assign n15537 = n1266 & n15536 ;
  assign n15538 = n15534 & n15537 ;
  assign n15539 = ~\pi0039  & ~n15538 ;
  assign n15540 = ~n15532 & n15539 ;
  assign n15541 = ~n15527 & ~n15540 ;
  assign n15542 = n13386 & n15541 ;
  assign n15543 = ~\pi0024  & n15529 ;
  assign n15544 = n11822 & n15543 ;
  assign n15545 = n1627 & n15544 ;
  assign n15546 = n1319 & n15545 ;
  assign n15547 = \pi0479  & ~n10050 ;
  assign n15548 = ~n1696 & n15547 ;
  assign n15549 = n1732 & n15548 ;
  assign n15550 = n1721 & n15549 ;
  assign n15551 = n1319 & n15550 ;
  assign n15552 = ~\pi0051  & \pi0096  ;
  assign n15553 = n1650 & n15552 ;
  assign n15554 = n1321 & n15553 ;
  assign n15555 = ~n15548 & n15554 ;
  assign n15556 = n1354 & n15555 ;
  assign n15557 = n1358 & n15556 ;
  assign n15558 = ~n15551 & ~n15557 ;
  assign n15559 = n1264 & n11822 ;
  assign n15560 = ~n15558 & n15559 ;
  assign n15561 = ~n15546 & ~n15560 ;
  assign n15562 = ~\pi0039  & n1264 ;
  assign n15563 = n1263 & n15562 ;
  assign n15564 = n8604 & n15563 ;
  assign n15565 = n6684 & n15563 ;
  assign n15566 = n15548 & n15565 ;
  assign n15567 = ~n15564 & ~n15566 ;
  assign n15568 = n8733 & ~n15567 ;
  assign n15569 = n1720 & n15568 ;
  assign n15570 = n11903 & n15569 ;
  assign n15571 = n6954 & ~n13629 ;
  assign n15572 = \pi0039  & \pi0593  ;
  assign n15573 = n11903 & n15572 ;
  assign n15574 = n15571 & n15573 ;
  assign n15575 = ~n15570 & ~n15574 ;
  assign n15576 = n11858 & ~n15575 ;
  assign n15577 = \pi0092  & n1281 ;
  assign n15578 = n1260 & n15577 ;
  assign n15579 = ~\pi0040  & ~\pi0092  ;
  assign n15580 = n1264 & n15579 ;
  assign n15581 = n10937 & n15580 ;
  assign n15582 = n10319 & n15581 ;
  assign n15583 = ~n15578 & ~n15582 ;
  assign n15584 = \pi0314  & \pi1050  ;
  assign n15585 = n1286 & n15584 ;
  assign n15586 = n2402 & n15585 ;
  assign n15587 = n12970 & n15586 ;
  assign n15588 = ~n15583 & n15587 ;
  assign n15589 = \pi0152  & ~\pi0166  ;
  assign n15590 = n6706 & n15589 ;
  assign n15591 = ~\pi0072  & \pi0161  ;
  assign n15592 = \pi0299  & n15591 ;
  assign n15593 = n15590 & n15592 ;
  assign n15594 = ~\pi0072  & \pi0174  ;
  assign n15595 = ~\pi0299  & n15594 ;
  assign n15596 = n11990 & n15595 ;
  assign n15597 = ~n15593 & ~n15596 ;
  assign n15598 = ~\pi0072  & \pi0099  ;
  assign n15599 = ~\pi0039  & ~n15598 ;
  assign n15600 = \pi0232  & ~n15599 ;
  assign n15601 = ~n15597 & n15600 ;
  assign n15602 = ~\pi0039  & n15598 ;
  assign n15603 = ~n8496 & ~n15602 ;
  assign n15604 = ~n15601 & n15603 ;
  assign n15605 = n9948 & ~n15604 ;
  assign n15606 = \pi0228  & n12165 ;
  assign n15607 = ~n2402 & ~n15602 ;
  assign n15608 = ~n15601 & n15607 ;
  assign n15609 = \pi0087  & ~n15608 ;
  assign n15610 = n15598 & n15609 ;
  assign n15611 = ~n15606 & n15610 ;
  assign n15612 = ~\pi0075  & ~n15609 ;
  assign n15613 = n1281 & n12430 ;
  assign n15614 = n1260 & n15613 ;
  assign n15615 = ~\pi0075  & n2402 ;
  assign n15616 = ~n15614 & n15615 ;
  assign n15617 = ~n15612 & ~n15616 ;
  assign n15618 = ~n15611 & ~n15617 ;
  assign n15619 = \pi0232  & n2363 ;
  assign n15620 = ~n15597 & n15619 ;
  assign n15621 = ~n6901 & ~n15620 ;
  assign n15622 = ~n2363 & n15602 ;
  assign n15623 = ~n2363 & n15600 ;
  assign n15624 = ~n15597 & n15623 ;
  assign n15625 = ~n15622 & ~n15624 ;
  assign n15626 = \pi0075  & n15625 ;
  assign n15627 = n15621 & n15626 ;
  assign n15628 = ~n8799 & n15598 ;
  assign n15629 = \pi0228  & ~n15628 ;
  assign n15630 = ~n8641 & n15629 ;
  assign n15631 = ~\pi0228  & ~n15598 ;
  assign n15632 = n8640 & ~n15598 ;
  assign n15633 = n8639 & n15632 ;
  assign n15634 = ~n15631 & ~n15633 ;
  assign n15635 = ~n15630 & n15634 ;
  assign n15636 = ~\pi0024  & ~\pi0101  ;
  assign n15637 = n6805 & n15636 ;
  assign n15638 = n7207 & n12865 ;
  assign n15639 = n15637 & n15638 ;
  assign n15640 = n12162 & n12211 ;
  assign n15641 = n15598 & ~n15640 ;
  assign n15642 = ~n15639 & ~n15641 ;
  assign n15643 = n12181 & n15634 ;
  assign n15644 = ~n15642 & n15643 ;
  assign n15645 = ~n15635 & ~n15644 ;
  assign n15646 = ~\pi0039  & n15626 ;
  assign n15647 = n15645 & n15646 ;
  assign n15648 = ~n15627 & ~n15647 ;
  assign n15649 = ~n15618 & n15648 ;
  assign n15650 = \pi0041  & \pi0072  ;
  assign n15651 = \pi0099  & ~n15650 ;
  assign n15652 = n8799 & ~n15651 ;
  assign n15653 = ~n12587 & n15652 ;
  assign n15654 = n8799 & n12013 ;
  assign n15655 = ~n12587 & n15654 ;
  assign n15656 = ~n12055 & n15655 ;
  assign n15657 = ~n15653 & ~n15656 ;
  assign n15658 = ~\pi0039  & ~n12595 ;
  assign n15659 = ~\pi0039  & \pi0099  ;
  assign n15660 = ~n15650 & n15659 ;
  assign n15661 = n12128 & n15660 ;
  assign n15662 = ~n15658 & ~n15661 ;
  assign n15663 = n12269 & n15651 ;
  assign n15664 = ~n12088 & n15663 ;
  assign n15665 = ~n12013 & n15651 ;
  assign n15666 = ~n12592 & ~n15665 ;
  assign n15667 = ~n15664 & n15666 ;
  assign n15668 = ~n15662 & ~n15667 ;
  assign n15669 = n15657 & n15668 ;
  assign n15670 = ~\pi0228  & ~n15662 ;
  assign n15671 = n11040 & ~n15597 ;
  assign n15672 = ~n12918 & n15671 ;
  assign n15673 = n2327 & ~n15672 ;
  assign n15674 = ~n15670 & n15673 ;
  assign n15675 = ~n15669 & n15674 ;
  assign n15676 = \pi0232  & ~n15597 ;
  assign n15677 = \pi0039  & ~n15676 ;
  assign n15678 = n15634 & ~n15677 ;
  assign n15679 = ~n15630 & n15678 ;
  assign n15680 = ~n12165 & n15598 ;
  assign n15681 = ~n12170 & n15598 ;
  assign n15682 = n6806 & n12369 ;
  assign n15683 = n1281 & n15682 ;
  assign n15684 = n1260 & n15683 ;
  assign n15685 = ~n15681 & ~n15684 ;
  assign n15686 = ~n15680 & n15685 ;
  assign n15687 = n12181 & n15678 ;
  assign n15688 = ~n15686 & n15687 ;
  assign n15689 = ~n15679 & ~n15688 ;
  assign n15690 = n6785 & ~n15671 ;
  assign n15691 = n15689 & n15690 ;
  assign n15692 = \pi0038  & ~n15602 ;
  assign n15693 = ~n15601 & n15692 ;
  assign n15694 = ~\pi0087  & ~n15693 ;
  assign n15695 = ~n15691 & n15694 ;
  assign n15696 = n15648 & n15695 ;
  assign n15697 = ~n15675 & n15696 ;
  assign n15698 = ~n15649 & ~n15697 ;
  assign n15699 = n15605 & ~n15698 ;
  assign n15700 = ~n15601 & ~n15602 ;
  assign n15701 = ~n8496 & n9948 ;
  assign n15702 = ~n15700 & n15701 ;
  assign n15703 = \pi0232  & n15591 ;
  assign n15704 = n15590 & n15703 ;
  assign n15705 = \pi0039  & ~n15704 ;
  assign n15706 = ~n9948 & ~n15599 ;
  assign n15707 = ~n15705 & n15706 ;
  assign n15708 = ~n15702 & ~n15707 ;
  assign n15709 = ~n15699 & n15708 ;
  assign n15710 = n8640 & n11700 ;
  assign n15711 = n11706 & ~n15710 ;
  assign n15712 = \pi0129  & ~n15711 ;
  assign n15713 = ~\pi0075  & n2341 ;
  assign n15714 = n6785 & n15713 ;
  assign n15715 = ~n11701 & n15714 ;
  assign n15716 = ~n15712 & n15715 ;
  assign n15717 = ~\pi0683  & ~n6808 ;
  assign n15718 = n10071 & ~n15717 ;
  assign n15719 = ~n6795 & n15714 ;
  assign n15720 = ~n15718 & n15719 ;
  assign n15721 = n11781 & ~n13720 ;
  assign n15722 = n10080 & n15721 ;
  assign n15723 = ~n15720 & ~n15722 ;
  assign n15724 = ~n15716 & n15723 ;
  assign n15725 = n1281 & n10017 ;
  assign n15726 = n1260 & n15725 ;
  assign n15727 = ~n15724 & n15726 ;
  assign n15728 = n6804 & n12275 ;
  assign n15729 = n8799 & n12012 ;
  assign n15730 = ~n15728 & n15729 ;
  assign n15731 = ~\pi0044  & n12211 ;
  assign n15732 = n15730 & ~n15731 ;
  assign n15733 = \pi0228  & ~n12012 ;
  assign n15734 = ~n12583 & ~n15733 ;
  assign n15735 = ~\pi0039  & ~n15734 ;
  assign n15736 = ~n8641 & n15735 ;
  assign n15737 = n8799 & ~n15728 ;
  assign n15738 = n12207 & n15737 ;
  assign n15739 = n15736 & ~n15738 ;
  assign n15740 = ~n15732 & n15739 ;
  assign n15741 = ~\pi0228  & ~n12012 ;
  assign n15742 = ~\pi0039  & n15741 ;
  assign n15743 = n8640 & ~n12012 ;
  assign n15744 = ~\pi0039  & n15743 ;
  assign n15745 = n8639 & n15744 ;
  assign n15746 = ~n15742 & ~n15745 ;
  assign n15747 = ~\pi0144  & \pi0174  ;
  assign n15748 = ~\pi0072  & n15747 ;
  assign n15749 = n12330 & n15748 ;
  assign n15750 = n10118 & n15749 ;
  assign n15751 = ~\pi0072  & ~\pi0161  ;
  assign n15752 = n10276 & n15751 ;
  assign n15753 = n15590 & n15752 ;
  assign n15754 = \pi0039  & ~n15753 ;
  assign n15755 = ~n15750 & n15754 ;
  assign n15756 = n2363 & ~n15755 ;
  assign n15757 = n15746 & n15756 ;
  assign n15758 = ~n15740 & n15757 ;
  assign n15759 = ~\pi0039  & ~n12012 ;
  assign n15760 = ~n2363 & ~n15759 ;
  assign n15761 = ~n15755 & n15760 ;
  assign n15762 = \pi0075  & ~n15761 ;
  assign n15763 = n8496 & n15762 ;
  assign n15764 = ~n15758 & n15763 ;
  assign n15765 = n12925 & ~n15753 ;
  assign n15766 = ~n15750 & n15765 ;
  assign n15767 = ~n8496 & n15759 ;
  assign n15768 = n9948 & ~n15767 ;
  assign n15769 = ~n15766 & n15768 ;
  assign n15770 = ~n15764 & n15769 ;
  assign n15771 = ~\pi0072  & \pi0232  ;
  assign n15772 = ~\pi0161  & n15771 ;
  assign n15773 = n15590 & n15772 ;
  assign n15774 = \pi0039  & ~n15773 ;
  assign n15775 = ~n9948 & ~n15759 ;
  assign n15776 = ~n15774 & n15775 ;
  assign n15777 = ~n15770 & ~n15776 ;
  assign n15778 = \pi0101  & ~n12043 ;
  assign n15779 = ~n12053 & n15778 ;
  assign n15780 = ~n12042 & n15779 ;
  assign n15781 = \pi0228  & n8799 ;
  assign n15782 = ~n12066 & n15781 ;
  assign n15783 = ~n15780 & n15782 ;
  assign n15784 = n12012 & ~n12088 ;
  assign n15785 = ~n12082 & n12580 ;
  assign n15786 = ~n15784 & n15785 ;
  assign n15787 = n12883 & ~n15753 ;
  assign n15788 = ~n15750 & n15787 ;
  assign n15789 = ~n12012 & n12800 ;
  assign n15790 = ~\pi0087  & ~n15789 ;
  assign n15791 = ~n15788 & n15790 ;
  assign n15792 = n12170 & n15737 ;
  assign n15793 = n12180 & n15792 ;
  assign n15794 = ~n12361 & n15730 ;
  assign n15795 = ~n15793 & ~n15794 ;
  assign n15796 = n15736 & n15795 ;
  assign n15797 = n15746 & ~n15755 ;
  assign n15798 = ~n15796 & n15797 ;
  assign n15799 = n6785 & ~n15798 ;
  assign n15800 = n15791 & ~n15799 ;
  assign n15801 = ~\pi0044  & ~n12125 ;
  assign n15802 = n15778 & ~n15801 ;
  assign n15803 = ~\pi0228  & ~n6806 ;
  assign n15804 = ~\pi0228  & ~n12143 ;
  assign n15805 = n12136 & n15804 ;
  assign n15806 = ~n15803 & ~n15805 ;
  assign n15807 = ~n15802 & ~n15806 ;
  assign n15808 = ~\pi0039  & ~n15807 ;
  assign n15809 = n15800 & n15808 ;
  assign n15810 = ~n15786 & n15809 ;
  assign n15811 = ~n15783 & n15810 ;
  assign n15812 = ~\pi0299  & n11040 ;
  assign n15813 = n15749 & n15812 ;
  assign n15814 = ~\pi0161  & n15590 ;
  assign n15815 = n11040 & n12512 ;
  assign n15816 = n15814 & n15815 ;
  assign n15817 = ~n15813 & ~n15816 ;
  assign n15818 = ~n12918 & ~n15817 ;
  assign n15819 = n2327 & ~n15818 ;
  assign n15820 = n15791 & ~n15819 ;
  assign n15821 = ~n15799 & n15820 ;
  assign n15822 = ~\pi0101  & n12841 ;
  assign n15823 = n1281 & n15822 ;
  assign n15824 = n1260 & n15823 ;
  assign n15825 = ~\pi0039  & ~n15824 ;
  assign n15826 = \pi0087  & ~n15755 ;
  assign n15827 = ~n15825 & n15826 ;
  assign n15828 = n1328 & n12825 ;
  assign n15829 = n1324 & n15828 ;
  assign n15830 = n1319 & n15829 ;
  assign n15831 = n12358 & n15830 ;
  assign n15832 = n12012 & n15826 ;
  assign n15833 = ~n15831 & n15832 ;
  assign n15834 = ~n15827 & ~n15833 ;
  assign n15835 = ~\pi0075  & n8496 ;
  assign n15836 = n15834 & n15835 ;
  assign n15837 = ~n15821 & n15836 ;
  assign n15838 = ~n15776 & n15837 ;
  assign n15839 = ~n15811 & n15838 ;
  assign n15840 = ~n15777 & ~n15839 ;
  assign n15841 = n13115 & n13527 ;
  assign n15842 = n11824 & n15841 ;
  assign n15843 = n1406 & n1531 ;
  assign n15844 = n1236 & n15843 ;
  assign n15845 = n1248 & n15844 ;
  assign n15846 = n15842 & n15845 ;
  assign n15847 = \pi0109  & n1256 ;
  assign n15848 = n1255 & n15847 ;
  assign n15849 = n1257 & n15848 ;
  assign n15850 = n1249 & n15849 ;
  assign n15851 = ~\pi0109  & ~\pi0314  ;
  assign n15852 = n15333 & n15851 ;
  assign n15853 = n1490 & n15852 ;
  assign n15854 = ~n15850 & ~n15853 ;
  assign n15855 = n1315 & n1327 ;
  assign n15856 = n11824 & n15855 ;
  assign n15857 = ~n15854 & n15856 ;
  assign n15858 = n12137 & n13042 ;
  assign n15859 = n1319 & n15858 ;
  assign n15860 = ~n6704 & n9012 ;
  assign n15861 = n6808 & n9250 ;
  assign n15862 = n8640 & n9250 ;
  assign n15863 = n8639 & n15862 ;
  assign n15864 = ~n15861 & ~n15863 ;
  assign n15865 = n15860 & n15864 ;
  assign n15866 = n15859 & ~n15865 ;
  assign n15867 = n11822 & n15866 ;
  assign n15868 = ~\pi0110  & ~n15393 ;
  assign n15869 = ~n6808 & ~n8641 ;
  assign n15870 = n8567 & n13003 ;
  assign n15871 = ~n15869 & n15870 ;
  assign n15872 = ~n15868 & n15871 ;
  assign n15873 = ~n6647 & n15872 ;
  assign n15874 = n13003 & n15394 ;
  assign n15875 = n15393 & n15874 ;
  assign n15876 = n15869 & n15875 ;
  assign n15877 = ~n15873 & ~n15876 ;
  assign n15878 = ~n6704 & ~n9250 ;
  assign n15879 = n11822 & n15878 ;
  assign n15880 = ~n15877 & n15879 ;
  assign n15881 = ~n15867 & ~n15880 ;
  assign n15882 = n10390 & n13089 ;
  assign n15883 = n13408 & n15882 ;
  assign n15884 = n1340 & n1341 ;
  assign n15885 = n1249 & n15884 ;
  assign n15886 = ~n15883 & ~n15885 ;
  assign n15887 = ~\pi0108  & \pi0841  ;
  assign n15888 = n1268 & n15887 ;
  assign n15889 = n1272 & n15888 ;
  assign n15890 = n11816 & n15889 ;
  assign n15891 = ~n15886 & n15890 ;
  assign n15892 = \pi0024  & n13410 ;
  assign n15893 = n1344 & n15892 ;
  assign n15894 = n1273 & n15893 ;
  assign n15895 = \pi0841  & n13089 ;
  assign n15896 = n15894 & n15895 ;
  assign n15897 = n13408 & n15896 ;
  assign n15898 = n1274 & n10018 ;
  assign n15899 = n13390 & n15898 ;
  assign n15900 = n1273 & n15899 ;
  assign n15901 = n1340 & n15900 ;
  assign n15902 = n1249 & n15901 ;
  assign n15903 = ~n15897 & ~n15902 ;
  assign n15904 = ~n15891 & n15903 ;
  assign n15905 = n11824 & ~n15904 ;
  assign n15906 = ~\pi0999  & n1255 ;
  assign n15907 = n13115 & n15906 ;
  assign n15908 = n11824 & n15907 ;
  assign n15909 = n1513 & n15908 ;
  assign n15910 = ~n1595 & n11939 ;
  assign n15911 = \pi0108  & ~n11916 ;
  assign n15912 = \pi0098  & n1276 ;
  assign n15913 = ~\pi0088  & ~\pi0097  ;
  assign n15914 = n1252 & n15913 ;
  assign n15915 = n15912 & n15914 ;
  assign n15916 = ~n11916 & n15915 ;
  assign n15917 = n1542 & n15916 ;
  assign n15918 = ~n15911 & ~n15917 ;
  assign n15919 = n8568 & ~n15918 ;
  assign n15920 = n15910 & n15919 ;
  assign n15921 = \pi0097  & n11916 ;
  assign n15922 = n8573 & n11916 ;
  assign n15923 = n1542 & n15922 ;
  assign n15924 = ~n15921 & ~n15923 ;
  assign n15925 = n8569 & ~n15924 ;
  assign n15926 = ~\pi0051  & ~\pi0087  ;
  assign n15927 = ~n15925 & n15926 ;
  assign n15928 = ~n15920 & n15927 ;
  assign n15929 = n2402 & n8592 ;
  assign n15930 = ~n8581 & n15929 ;
  assign n15931 = ~\pi0087  & ~n15930 ;
  assign n15932 = ~\pi0075  & n10017 ;
  assign n15933 = ~\pi0087  & n15932 ;
  assign n15934 = n6629 & n15932 ;
  assign n15935 = n1638 & n15934 ;
  assign n15936 = ~n15933 & ~n15935 ;
  assign n15937 = ~n15931 & ~n15936 ;
  assign n15938 = ~n15928 & n15937 ;
  assign n15939 = n1542 & n14002 ;
  assign n15940 = ~\pi0058  & \pi0314  ;
  assign n15941 = n1274 & n15940 ;
  assign n15942 = n1273 & n15941 ;
  assign n15943 = n11824 & n15942 ;
  assign n15944 = n15939 & n15943 ;
  assign n15945 = ~\pi0082  & \pi0111  ;
  assign n15946 = n1270 & n15945 ;
  assign n15947 = n8567 & n15946 ;
  assign n15948 = n1315 & n15947 ;
  assign n15949 = n13152 & n15948 ;
  assign n15950 = n13153 & n15949 ;
  assign n15951 = \pi0314  & n1412 ;
  assign n15952 = n11824 & n15951 ;
  assign n15953 = n15950 & n15952 ;
  assign n15954 = n1319 & n12137 ;
  assign n15955 = ~n6808 & n15860 ;
  assign n15956 = ~n8641 & n15955 ;
  assign n15957 = n11824 & n15956 ;
  assign n15958 = n15954 & n15957 ;
  assign n15959 = ~n15953 & ~n15958 ;
  assign n15960 = ~\pi0024  & \pi0072  ;
  assign n15961 = n1328 & n15960 ;
  assign n15962 = n1324 & n15961 ;
  assign n15963 = n1319 & n15962 ;
  assign n15964 = ~\pi0035  & ~\pi0314  ;
  assign n15965 = n1320 & n15964 ;
  assign n15966 = n1618 & n15965 ;
  assign n15967 = n13153 & n15966 ;
  assign n15968 = n1412 & n15967 ;
  assign n15969 = n15949 & n15968 ;
  assign n15970 = ~n15963 & ~n15969 ;
  assign n15971 = ~\pi0095  & n1634 ;
  assign n15972 = n11822 & n15971 ;
  assign n15973 = ~n15970 & n15972 ;
  assign n15974 = \pi0124  & ~\pi0468  ;
  assign n15975 = ~\pi0113  & n12592 ;
  assign n15976 = n2327 & ~n15975 ;
  assign n15977 = n2327 & n8799 ;
  assign n15978 = ~n12587 & n15977 ;
  assign n15979 = ~n15976 & ~n15978 ;
  assign n15980 = \pi0228  & ~n15979 ;
  assign n15981 = \pi0113  & ~n12264 ;
  assign n15982 = n8799 & n15981 ;
  assign n15983 = ~n12056 & n15982 ;
  assign n15984 = ~\pi0099  & ~n12092 ;
  assign n15985 = ~n12091 & n15984 ;
  assign n15986 = n15981 & ~n15985 ;
  assign n15987 = ~n15983 & ~n15986 ;
  assign n15988 = n15980 & n15987 ;
  assign n15989 = ~\pi0113  & n6806 ;
  assign n15990 = n6805 & n15989 ;
  assign n15991 = ~n12313 & n15990 ;
  assign n15992 = ~\pi0228  & ~n15991 ;
  assign n15993 = ~\pi0039  & ~n15992 ;
  assign n15994 = ~\pi0039  & n15981 ;
  assign n15995 = n12308 & n15994 ;
  assign n15996 = ~n15993 & ~n15995 ;
  assign n15997 = n2327 & n15996 ;
  assign n15998 = ~\pi0113  & n12430 ;
  assign n15999 = n1281 & n15998 ;
  assign n16000 = n1260 & n15999 ;
  assign n16001 = n2402 & n16000 ;
  assign n16002 = n2402 & n12261 ;
  assign n16003 = ~n12421 & n16002 ;
  assign n16004 = ~n16001 & ~n16003 ;
  assign n16005 = ~\pi0039  & n12261 ;
  assign n16006 = ~n2327 & n16005 ;
  assign n16007 = \pi0087  & ~n16006 ;
  assign n16008 = n16004 & n16007 ;
  assign n16009 = \pi0038  & ~n16005 ;
  assign n16010 = n12275 & n12583 ;
  assign n16011 = ~n8641 & n16010 ;
  assign n16012 = n12361 & n16011 ;
  assign n16013 = n6804 & n12583 ;
  assign n16014 = ~n8641 & n16013 ;
  assign n16015 = n16005 & ~n16014 ;
  assign n16016 = ~n16012 & n16015 ;
  assign n16017 = ~\pi0113  & n12583 ;
  assign n16018 = ~n6804 & n16017 ;
  assign n16019 = ~n8641 & n16018 ;
  assign n16020 = ~\pi0039  & n16019 ;
  assign n16021 = n15684 & n16020 ;
  assign n16022 = n6785 & ~n16021 ;
  assign n16023 = ~n16016 & n16022 ;
  assign n16024 = ~n16009 & ~n16023 ;
  assign n16025 = ~n16008 & n16024 ;
  assign n16026 = ~n15997 & n16025 ;
  assign n16027 = ~n15988 & n16026 ;
  assign n16028 = n15932 & n16007 ;
  assign n16029 = n16004 & n16028 ;
  assign n16030 = ~n15933 & ~n16029 ;
  assign n16031 = ~n16027 & ~n16030 ;
  assign n16032 = ~n2363 & n16005 ;
  assign n16033 = \pi0075  & ~n2342 ;
  assign n16034 = ~n16032 & n16033 ;
  assign n16035 = ~n8641 & n12583 ;
  assign n16036 = n6804 & n16035 ;
  assign n16037 = n6807 & n16035 ;
  assign n16038 = n12211 & n16037 ;
  assign n16039 = ~n16036 & ~n16038 ;
  assign n16040 = n12261 & n16039 ;
  assign n16041 = \pi0075  & ~n16032 ;
  assign n16042 = n15684 & n16019 ;
  assign n16043 = n12451 & n16042 ;
  assign n16044 = n16041 & ~n16043 ;
  assign n16045 = ~n16040 & n16044 ;
  assign n16046 = ~n16034 & ~n16045 ;
  assign n16047 = n10017 & ~n16046 ;
  assign n16048 = ~n10017 & ~n16005 ;
  assign n16049 = ~n16047 & ~n16048 ;
  assign n16050 = ~n16031 & n16049 ;
  assign n16051 = n6799 & ~n12595 ;
  assign n16052 = ~n12593 & n16051 ;
  assign n16053 = ~n12588 & n16052 ;
  assign n16054 = ~\pi0114  & ~n16053 ;
  assign n16055 = ~n12605 & ~n16054 ;
  assign n16056 = n12585 & n16055 ;
  assign n16057 = ~\pi0114  & n16051 ;
  assign n16058 = ~n12593 & n16057 ;
  assign n16059 = ~n12588 & n16058 ;
  assign n16060 = ~\pi0115  & n2327 ;
  assign n16061 = ~n16059 & n16060 ;
  assign n16062 = ~n16056 & n16061 ;
  assign n16063 = ~\pi0072  & \pi0114  ;
  assign n16064 = \pi0115  & ~n16063 ;
  assign n16065 = ~\pi0039  & ~n16064 ;
  assign n16066 = n2327 & ~n16065 ;
  assign n16067 = ~\pi0115  & n12583 ;
  assign n16068 = ~n8641 & n16067 ;
  assign n16069 = n13225 & n16068 ;
  assign n16070 = n12211 & n16069 ;
  assign n16071 = ~\pi0116  & n16070 ;
  assign n16072 = n2342 & n16063 ;
  assign n16073 = ~n16071 & n16072 ;
  assign n16074 = ~\pi0024  & n12583 ;
  assign n16075 = ~n8641 & n16074 ;
  assign n16076 = ~\pi0114  & ~\pi0115  ;
  assign n16077 = ~n12371 & n16076 ;
  assign n16078 = n12369 & n16077 ;
  assign n16079 = n16075 & n16078 ;
  assign n16080 = n12367 & n16079 ;
  assign n16081 = n2342 & n7207 ;
  assign n16082 = n16080 & n16081 ;
  assign n16083 = ~\pi0039  & n16063 ;
  assign n16084 = ~n2363 & n16083 ;
  assign n16085 = \pi0075  & ~n16084 ;
  assign n16086 = ~n16082 & n16085 ;
  assign n16087 = ~n16073 & n16086 ;
  assign n16088 = n11407 & n16063 ;
  assign n16089 = ~n2855 & ~n16088 ;
  assign n16090 = ~n6785 & ~n16089 ;
  assign n16091 = ~n12363 & n16063 ;
  assign n16092 = ~\pi0114  & ~n12371 ;
  assign n16093 = n12369 & n16092 ;
  assign n16094 = n12367 & n16093 ;
  assign n16095 = \pi0228  & n12291 ;
  assign n16096 = ~n8641 & n16095 ;
  assign n16097 = ~n16094 & n16096 ;
  assign n16098 = ~n16091 & n16097 ;
  assign n16099 = ~n16063 & ~n16096 ;
  assign n16100 = ~\pi0039  & ~n16089 ;
  assign n16101 = ~n16099 & n16100 ;
  assign n16102 = ~n16098 & n16101 ;
  assign n16103 = ~n16090 & ~n16102 ;
  assign n16104 = ~n16087 & ~n16103 ;
  assign n16105 = ~n16066 & n16104 ;
  assign n16106 = ~n16062 & n16105 ;
  assign n16107 = n10017 & n16087 ;
  assign n16108 = n12421 & n12422 ;
  assign n16109 = n16063 & ~n16108 ;
  assign n16110 = n12422 & n12430 ;
  assign n16111 = n1281 & n16110 ;
  assign n16112 = n1260 & n16111 ;
  assign n16113 = ~\pi0114  & n16112 ;
  assign n16114 = n2327 & ~n16113 ;
  assign n16115 = ~n16109 & n16114 ;
  assign n16116 = ~n2327 & ~n16083 ;
  assign n16117 = n13220 & ~n16116 ;
  assign n16118 = ~n16115 & n16117 ;
  assign n16119 = n15932 & ~n16118 ;
  assign n16120 = ~n16107 & ~n16119 ;
  assign n16121 = ~n16106 & ~n16120 ;
  assign n16122 = ~n10017 & ~n16083 ;
  assign n16123 = ~n16121 & ~n16122 ;
  assign n16124 = ~\pi0115  & ~n16053 ;
  assign n16125 = ~\pi0039  & ~n12605 ;
  assign n16126 = ~n16124 & n16125 ;
  assign n16127 = n12585 & n16126 ;
  assign n16128 = ~\pi0039  & ~\pi0115  ;
  assign n16129 = n16053 & n16128 ;
  assign n16130 = n2327 & n6799 ;
  assign n16131 = n12421 & n16130 ;
  assign n16132 = ~\pi0072  & \pi0115  ;
  assign n16133 = ~\pi0039  & n16132 ;
  assign n16134 = ~n2327 & ~n16133 ;
  assign n16135 = n13220 & ~n16134 ;
  assign n16136 = n16132 & n16135 ;
  assign n16137 = ~n16131 & n16136 ;
  assign n16138 = n16112 & n16135 ;
  assign n16139 = ~\pi0075  & n2327 ;
  assign n16140 = ~n16138 & n16139 ;
  assign n16141 = ~n16137 & n16140 ;
  assign n16142 = ~n16129 & n16141 ;
  assign n16143 = ~n16127 & n16142 ;
  assign n16144 = ~\pi0024  & n16035 ;
  assign n16145 = n7207 & n16144 ;
  assign n16146 = ~\pi0052  & ~\pi0114  ;
  assign n16147 = n12370 & n16146 ;
  assign n16148 = ~\pi0115  & ~n16147 ;
  assign n16149 = n12369 & n16148 ;
  assign n16150 = n12367 & n16149 ;
  assign n16151 = n16145 & n16150 ;
  assign n16152 = n2342 & n16151 ;
  assign n16153 = ~\pi0116  & n12583 ;
  assign n16154 = ~n8641 & n16153 ;
  assign n16155 = n13225 & n16154 ;
  assign n16156 = n12211 & n16155 ;
  assign n16157 = n2342 & n16132 ;
  assign n16158 = ~n16156 & n16157 ;
  assign n16159 = ~n2363 & n16133 ;
  assign n16160 = \pi0075  & ~n16159 ;
  assign n16161 = ~n16158 & n16160 ;
  assign n16162 = ~n16152 & n16161 ;
  assign n16163 = ~n12363 & n16132 ;
  assign n16164 = n16035 & ~n16150 ;
  assign n16165 = ~n16163 & n16164 ;
  assign n16166 = ~n12583 & ~n16132 ;
  assign n16167 = n8640 & ~n16132 ;
  assign n16168 = n8639 & n16167 ;
  assign n16169 = ~n16166 & ~n16168 ;
  assign n16170 = n11407 & n16132 ;
  assign n16171 = ~n2855 & ~n16170 ;
  assign n16172 = ~\pi0039  & ~n16171 ;
  assign n16173 = n16169 & n16172 ;
  assign n16174 = ~n16165 & n16173 ;
  assign n16175 = ~n6785 & ~n16171 ;
  assign n16176 = ~\pi0075  & ~n16175 ;
  assign n16177 = ~n16138 & n16176 ;
  assign n16178 = ~n16137 & n16177 ;
  assign n16179 = ~n16174 & n16178 ;
  assign n16180 = ~n16162 & ~n16179 ;
  assign n16181 = ~n16143 & n16180 ;
  assign n16182 = n10017 & ~n16181 ;
  assign n16183 = ~n10017 & ~n16133 ;
  assign n16184 = ~n16182 & ~n16183 ;
  assign n16185 = n12211 & n13225 ;
  assign n16186 = n12262 & ~n16185 ;
  assign n16187 = n6799 & n15637 ;
  assign n16188 = n15638 & n16187 ;
  assign n16189 = ~n16186 & ~n16188 ;
  assign n16190 = n2342 & n12583 ;
  assign n16191 = ~n6804 & n16190 ;
  assign n16192 = ~n8641 & n16191 ;
  assign n16193 = ~n16189 & n16192 ;
  assign n16194 = n12262 & ~n12583 ;
  assign n16195 = n8640 & n12262 ;
  assign n16196 = n8639 & n16195 ;
  assign n16197 = ~n16194 & ~n16196 ;
  assign n16198 = n2342 & ~n16197 ;
  assign n16199 = ~\pi0039  & n12262 ;
  assign n16200 = ~n2363 & n16199 ;
  assign n16201 = \pi0075  & ~n16200 ;
  assign n16202 = ~n16198 & n16201 ;
  assign n16203 = ~n16193 & n16202 ;
  assign n16204 = n11407 & n12262 ;
  assign n16205 = ~n2855 & ~n16204 ;
  assign n16206 = ~n6785 & ~n16205 ;
  assign n16207 = ~\pi0101  & ~\pi0113  ;
  assign n16208 = n6805 & n16207 ;
  assign n16209 = n12361 & n16208 ;
  assign n16210 = n12262 & n12583 ;
  assign n16211 = ~n6804 & n16210 ;
  assign n16212 = ~n8641 & n16211 ;
  assign n16213 = ~n16209 & n16212 ;
  assign n16214 = ~n6804 & n12583 ;
  assign n16215 = ~n8641 & n16214 ;
  assign n16216 = n12369 & n16215 ;
  assign n16217 = n12367 & n16216 ;
  assign n16218 = n16197 & ~n16217 ;
  assign n16219 = ~n16213 & n16218 ;
  assign n16220 = ~\pi0039  & ~n16205 ;
  assign n16221 = ~n16219 & n16220 ;
  assign n16222 = ~n16206 & ~n16221 ;
  assign n16223 = \pi0100  & ~n16199 ;
  assign n16224 = n13220 & ~n16223 ;
  assign n16225 = ~\pi0075  & ~n16224 ;
  assign n16226 = ~\pi0038  & ~\pi0113  ;
  assign n16227 = n12421 & n16226 ;
  assign n16228 = ~\pi0038  & n12262 ;
  assign n16229 = ~n16199 & ~n16228 ;
  assign n16230 = ~n16227 & ~n16229 ;
  assign n16231 = \pi0038  & ~n16199 ;
  assign n16232 = n6799 & n12430 ;
  assign n16233 = n1281 & n16232 ;
  assign n16234 = n1260 & n16233 ;
  assign n16235 = ~n16231 & n16234 ;
  assign n16236 = n8601 & ~n16235 ;
  assign n16237 = ~n16230 & n16236 ;
  assign n16238 = ~n16225 & ~n16237 ;
  assign n16239 = n16222 & ~n16238 ;
  assign n16240 = \pi0072  & \pi0113  ;
  assign n16241 = ~n12264 & ~n16240 ;
  assign n16242 = ~n8799 & ~n12261 ;
  assign n16243 = ~n16241 & n16242 ;
  assign n16244 = n12267 & n16242 ;
  assign n16245 = ~n12270 & n16244 ;
  assign n16246 = ~n16243 & ~n16245 ;
  assign n16247 = \pi0116  & n16246 ;
  assign n16248 = n6805 & n8799 ;
  assign n16249 = ~n12058 & n16248 ;
  assign n16250 = n12065 & n16249 ;
  assign n16251 = n6799 & n16250 ;
  assign n16252 = n6799 & ~n8799 ;
  assign n16253 = ~n12279 & n16252 ;
  assign n16254 = ~n12064 & n16253 ;
  assign n16255 = \pi0228  & ~n16254 ;
  assign n16256 = ~n16251 & n16255 ;
  assign n16257 = ~n16247 & n16256 ;
  assign n16258 = ~n12261 & ~n16241 ;
  assign n16259 = ~n12261 & n12267 ;
  assign n16260 = ~n12055 & n16259 ;
  assign n16261 = ~n16258 & ~n16260 ;
  assign n16262 = n8799 & n16255 ;
  assign n16263 = ~n16251 & n16262 ;
  assign n16264 = ~n16261 & n16263 ;
  assign n16265 = n6805 & n12365 ;
  assign n16266 = ~n12313 & n16265 ;
  assign n16267 = ~\pi0228  & ~n16266 ;
  assign n16268 = ~\pi0039  & ~n16267 ;
  assign n16269 = ~\pi0039  & \pi0116  ;
  assign n16270 = n12261 & n16269 ;
  assign n16271 = n16241 & n16269 ;
  assign n16272 = n12308 & n16271 ;
  assign n16273 = ~n16270 & ~n16272 ;
  assign n16274 = ~n16268 & n16273 ;
  assign n16275 = ~n16264 & ~n16274 ;
  assign n16276 = ~n16257 & n16275 ;
  assign n16277 = n2327 & ~n16238 ;
  assign n16278 = ~n16276 & n16277 ;
  assign n16279 = ~n16239 & ~n16278 ;
  assign n16280 = ~n16203 & n16279 ;
  assign n16281 = n10017 & ~n16280 ;
  assign n16282 = ~n10017 & ~n16199 ;
  assign n16283 = ~n16281 & ~n16282 ;
  assign n16284 = \pi0062  & ~n6633 ;
  assign n16285 = n2467 & ~n16284 ;
  assign n16286 = ~\pi0074  & n6630 ;
  assign n16287 = n1638 & n16286 ;
  assign n16288 = \pi0055  & ~n16287 ;
  assign n16289 = ~n6834 & ~n16288 ;
  assign n16290 = ~n2423 & n16289 ;
  assign n16291 = ~\pi0075  & ~\pi0087  ;
  assign n16292 = ~\pi0075  & n6629 ;
  assign n16293 = n1638 & n16292 ;
  assign n16294 = ~n16291 & ~n16293 ;
  assign n16295 = ~\pi0092  & n16294 ;
  assign n16296 = n2851 & ~n8463 ;
  assign n16297 = n8460 & n16296 ;
  assign n16298 = ~n2596 & ~n16297 ;
  assign n16299 = ~n2594 & n16298 ;
  assign n16300 = \pi0100  & ~n16297 ;
  assign n16301 = ~\pi0038  & ~n16300 ;
  assign n16302 = ~n16299 & n16301 ;
  assign n16303 = n4539 & ~n16302 ;
  assign n16304 = ~n16295 & ~n16303 ;
  assign n16305 = n2511 & ~n8420 ;
  assign n16306 = n16289 & n16305 ;
  assign n16307 = n16304 & n16306 ;
  assign n16308 = ~n16290 & ~n16307 ;
  assign n16309 = ~\pi0062  & n16308 ;
  assign n16310 = n16285 & ~n16309 ;
  assign n16311 = \pi0163  & ~n6706 ;
  assign n16312 = ~\pi0150  & \pi0232  ;
  assign n16313 = ~n8601 & n16312 ;
  assign n16314 = ~n16311 & n16313 ;
  assign n16315 = ~n14029 & n16314 ;
  assign n16316 = \pi0150  & ~\pi0163  ;
  assign n16317 = n11129 & n16316 ;
  assign n16318 = n11126 & n16317 ;
  assign n16319 = \pi0165  & \pi0232  ;
  assign n16320 = n6706 & n16319 ;
  assign n16321 = n8601 & ~n10134 ;
  assign n16322 = ~n16320 & n16321 ;
  assign n16323 = ~\pi0074  & n16322 ;
  assign n16324 = ~n16318 & ~n16323 ;
  assign n16325 = ~n16315 & n16324 ;
  assign n16326 = ~n1292 & ~n2467 ;
  assign n16327 = ~n11149 & ~n16326 ;
  assign n16328 = n16325 & ~n16327 ;
  assign n16329 = n2467 & ~n16328 ;
  assign n16330 = n10128 & ~n16320 ;
  assign n16331 = ~n16318 & ~n16330 ;
  assign n16332 = ~n16315 & n16331 ;
  assign n16333 = ~n2467 & ~n16332 ;
  assign n16334 = \pi0118  & ~n16333 ;
  assign n16335 = ~n16329 & n16334 ;
  assign n16336 = n6706 & n10735 ;
  assign n16337 = \pi0151  & ~\pi0168  ;
  assign n16338 = ~n16336 & n16337 ;
  assign n16339 = \pi0168  & ~n10578 ;
  assign n16340 = n6706 & n16339 ;
  assign n16341 = ~n10743 & n16340 ;
  assign n16342 = ~\pi0168  & ~n10363 ;
  assign n16343 = ~n10642 & n16342 ;
  assign n16344 = ~\pi0151  & ~n16343 ;
  assign n16345 = ~\pi0151  & ~n10741 ;
  assign n16346 = ~n10751 & n16345 ;
  assign n16347 = ~n16344 & ~n16346 ;
  assign n16348 = ~n16341 & ~n16347 ;
  assign n16349 = ~n16338 & ~n16348 ;
  assign n16350 = \pi0168  & n10588 ;
  assign n16351 = ~n10363 & n16350 ;
  assign n16352 = \pi0168  & n6706 ;
  assign n16353 = ~n10586 & ~n16352 ;
  assign n16354 = ~n10363 & n16353 ;
  assign n16355 = ~\pi0151  & ~n16354 ;
  assign n16356 = ~n16351 & n16355 ;
  assign n16357 = ~\pi0150  & ~n16356 ;
  assign n16358 = \pi0299  & ~n16357 ;
  assign n16359 = ~n6706 & n10586 ;
  assign n16360 = ~n6706 & n10358 ;
  assign n16361 = ~n10362 & n16360 ;
  assign n16362 = ~n16359 & ~n16361 ;
  assign n16363 = ~\pi0168  & n16362 ;
  assign n16364 = \pi0151  & ~n16363 ;
  assign n16365 = ~n10363 & ~n10456 ;
  assign n16366 = \pi0151  & n6706 ;
  assign n16367 = ~n16365 & n16366 ;
  assign n16368 = ~n16364 & ~n16367 ;
  assign n16369 = \pi0168  & n16362 ;
  assign n16370 = ~n10787 & n16369 ;
  assign n16371 = \pi0299  & ~n16370 ;
  assign n16372 = ~n16368 & n16371 ;
  assign n16373 = ~n16358 & ~n16372 ;
  assign n16374 = ~n6706 & ~n10586 ;
  assign n16375 = ~n10363 & n16374 ;
  assign n16376 = ~n16373 & ~n16375 ;
  assign n16377 = ~n16349 & n16376 ;
  assign n16378 = \pi0151  & \pi0168  ;
  assign n16379 = n6706 & ~n10366 ;
  assign n16380 = ~\pi0210  & n6706 ;
  assign n16381 = ~n10375 & n16380 ;
  assign n16382 = ~n16379 & ~n16381 ;
  assign n16383 = n16378 & ~n16382 ;
  assign n16384 = ~n16362 & n16378 ;
  assign n16385 = \pi0150  & ~n16384 ;
  assign n16386 = ~n16383 & n16385 ;
  assign n16387 = ~n16373 & ~n16386 ;
  assign n16388 = \pi0173  & n6706 ;
  assign n16389 = n11239 & n16388 ;
  assign n16390 = ~\pi0173  & ~n10363 ;
  assign n16391 = ~n10642 & n16390 ;
  assign n16392 = n10637 & n16391 ;
  assign n16393 = n6706 & n16392 ;
  assign n16394 = \pi0185  & ~\pi0299  ;
  assign n16395 = ~n16375 & n16394 ;
  assign n16396 = ~n16393 & n16395 ;
  assign n16397 = ~n16389 & n16396 ;
  assign n16398 = \pi0173  & n16362 ;
  assign n16399 = \pi0095  & ~\pi0173  ;
  assign n16400 = ~\pi0040  & ~\pi0173  ;
  assign n16401 = n1256 & n16400 ;
  assign n16402 = ~n16399 & ~n16401 ;
  assign n16403 = ~\pi0185  & n16402 ;
  assign n16404 = ~\pi0185  & n10358 ;
  assign n16405 = ~n10362 & n16404 ;
  assign n16406 = ~n16403 & ~n16405 ;
  assign n16407 = ~n16398 & ~n16406 ;
  assign n16408 = n6706 & ~n16406 ;
  assign n16409 = ~n16365 & n16408 ;
  assign n16410 = ~n16407 & ~n16409 ;
  assign n16411 = ~\pi0190  & \pi0232  ;
  assign n16412 = n16410 & n16411 ;
  assign n16413 = ~n10276 & ~n16412 ;
  assign n16414 = ~n16397 & ~n16413 ;
  assign n16415 = ~\pi0173  & ~n10578 ;
  assign n16416 = n6706 & n16415 ;
  assign n16417 = ~n10574 & n16416 ;
  assign n16418 = ~\pi0173  & ~n6706 ;
  assign n16419 = ~n10586 & n16418 ;
  assign n16420 = ~n10363 & n16419 ;
  assign n16421 = \pi0185  & ~n16398 ;
  assign n16422 = \pi0185  & n6706 ;
  assign n16423 = ~n10366 & n16422 ;
  assign n16424 = ~\pi0198  & n16422 ;
  assign n16425 = ~n10375 & n16424 ;
  assign n16426 = ~n16423 & ~n16425 ;
  assign n16427 = ~n16421 & n16426 ;
  assign n16428 = ~n16420 & ~n16427 ;
  assign n16429 = ~n16417 & n16428 ;
  assign n16430 = \pi0185  & \pi0190  ;
  assign n16431 = ~n10482 & n16388 ;
  assign n16432 = ~n10481 & n16431 ;
  assign n16433 = \pi0173  & ~n16362 ;
  assign n16434 = ~\pi0173  & ~n10588 ;
  assign n16435 = ~\pi0173  & n10358 ;
  assign n16436 = ~n10362 & n16435 ;
  assign n16437 = ~n16434 & ~n16436 ;
  assign n16438 = ~n16375 & ~n16437 ;
  assign n16439 = \pi0190  & ~n16438 ;
  assign n16440 = ~n16433 & n16439 ;
  assign n16441 = ~n16432 & n16440 ;
  assign n16442 = ~n16430 & ~n16441 ;
  assign n16443 = \pi0232  & ~n16442 ;
  assign n16444 = ~n16429 & n16443 ;
  assign n16445 = ~n16414 & ~n16444 ;
  assign n16446 = ~n16387 & ~n16445 ;
  assign n16447 = ~n16377 & n16446 ;
  assign n16448 = ~\pi0087  & ~\pi0100  ;
  assign n16449 = \pi0143  & ~\pi0165  ;
  assign n16450 = n10195 & n16449 ;
  assign n16451 = ~n8375 & n16450 ;
  assign n16452 = \pi0038  & ~n16451 ;
  assign n16453 = n16448 & ~n16452 ;
  assign n16454 = ~\pi0143  & ~n10201 ;
  assign n16455 = \pi0143  & n6784 ;
  assign n16456 = n1266 & n16455 ;
  assign n16457 = n1354 & n16456 ;
  assign n16458 = n1358 & n16457 ;
  assign n16459 = ~\pi0143  & \pi0165  ;
  assign n16460 = ~n16320 & ~n16459 ;
  assign n16461 = ~n16458 & ~n16460 ;
  assign n16462 = n2362 & n16461 ;
  assign n16463 = ~n16454 & n16462 ;
  assign n16464 = ~n16453 & ~n16463 ;
  assign n16465 = ~\pi0039  & ~n16464 ;
  assign n16466 = ~\pi0232  & ~n10586 ;
  assign n16467 = ~n10363 & n16466 ;
  assign n16468 = n16465 & ~n16467 ;
  assign n16469 = ~n16447 & n16468 ;
  assign n16470 = \pi0178  & \pi0190  ;
  assign n16471 = n10217 & n16470 ;
  assign n16472 = n10231 & n16471 ;
  assign n16473 = ~\pi0178  & \pi0190  ;
  assign n16474 = n10217 & n16473 ;
  assign n16475 = n10229 & n16474 ;
  assign n16476 = n10173 & n16475 ;
  assign n16477 = \pi0178  & ~\pi0190  ;
  assign n16478 = n10217 & n16477 ;
  assign n16479 = n10216 & n16478 ;
  assign n16480 = n10173 & n16479 ;
  assign n16481 = ~n16476 & ~n16480 ;
  assign n16482 = ~n16472 & n16481 ;
  assign n16483 = n3058 & n6771 ;
  assign n16484 = n6706 & n16483 ;
  assign n16485 = ~n6761 & n16484 ;
  assign n16486 = ~n16482 & n16485 ;
  assign n16487 = \pi0168  & n10217 ;
  assign n16488 = n10229 & n16487 ;
  assign n16489 = n10173 & n16488 ;
  assign n16490 = \pi0157  & n10217 ;
  assign n16491 = n10216 & n16490 ;
  assign n16492 = n10173 & n16491 ;
  assign n16493 = ~n16489 & ~n16492 ;
  assign n16494 = ~n6732 & n11062 ;
  assign n16495 = n6706 & n16494 ;
  assign n16496 = ~n16493 & n16495 ;
  assign n16497 = ~\pi0040  & \pi0232  ;
  assign n16498 = n1256 & n16497 ;
  assign n16499 = ~n16496 & n16498 ;
  assign n16500 = ~n16486 & n16499 ;
  assign n16501 = n1256 & n14534 ;
  assign n16502 = \pi0039  & ~n16501 ;
  assign n16503 = ~n16500 & n16502 ;
  assign n16504 = ~\pi0038  & ~n16503 ;
  assign n16505 = ~n16464 & ~n16504 ;
  assign n16506 = ~\pi0150  & ~n16311 ;
  assign n16507 = ~n14029 & n16506 ;
  assign n16508 = n11126 & n16316 ;
  assign n16509 = \pi0299  & ~n16508 ;
  assign n16510 = ~n16507 & n16509 ;
  assign n16511 = ~\pi0185  & n6706 ;
  assign n16512 = ~\pi0184  & n6706 ;
  assign n16513 = ~n14050 & n16512 ;
  assign n16514 = ~n16511 & ~n16513 ;
  assign n16515 = ~\pi0184  & ~\pi0185  ;
  assign n16516 = ~n14050 & n16515 ;
  assign n16517 = \pi0232  & ~n16516 ;
  assign n16518 = ~n16514 & n16517 ;
  assign n16519 = ~n10276 & ~n16518 ;
  assign n16520 = ~n16510 & ~n16519 ;
  assign n16521 = \pi0100  & ~n16520 ;
  assign n16522 = ~\pi0143  & ~\pi0299  ;
  assign n16523 = ~\pi0165  & \pi0299  ;
  assign n16524 = ~n16522 & ~n16523 ;
  assign n16525 = n8640 & n16524 ;
  assign n16526 = \pi0038  & ~n16525 ;
  assign n16527 = ~\pi0178  & ~\pi0299  ;
  assign n16528 = ~\pi0157  & \pi0299  ;
  assign n16529 = ~n16527 & ~n16528 ;
  assign n16530 = n8640 & n16529 ;
  assign n16531 = ~\pi0100  & n16530 ;
  assign n16532 = ~n16526 & n16531 ;
  assign n16533 = n10176 & n16532 ;
  assign n16534 = n10173 & n16533 ;
  assign n16535 = ~\pi0100  & ~n10156 ;
  assign n16536 = ~n16526 & n16535 ;
  assign n16537 = ~n16534 & ~n16536 ;
  assign n16538 = ~n16521 & n16537 ;
  assign n16539 = n6895 & ~n16538 ;
  assign n16540 = \pi0075  & ~n16520 ;
  assign n16541 = ~n10156 & n11470 ;
  assign n16542 = ~n16526 & n16541 ;
  assign n16543 = ~\pi0100  & ~n16542 ;
  assign n16544 = n16520 & ~n16542 ;
  assign n16545 = ~n16543 & ~n16544 ;
  assign n16546 = ~n16540 & ~n16545 ;
  assign n16547 = ~n16539 & n16546 ;
  assign n16548 = ~n16505 & n16547 ;
  assign n16549 = ~n16469 & n16548 ;
  assign n16550 = ~n2364 & ~n16540 ;
  assign n16551 = ~n16539 & n16550 ;
  assign n16552 = n2511 & ~n16551 ;
  assign n16553 = ~n16549 & n16552 ;
  assign n16554 = ~\pi0055  & ~\pi0074  ;
  assign n16555 = ~n8601 & ~n16519 ;
  assign n16556 = ~\pi0055  & ~n16510 ;
  assign n16557 = n16555 & n16556 ;
  assign n16558 = ~n16554 & ~n16557 ;
  assign n16559 = ~n16510 & n16555 ;
  assign n16560 = n8601 & ~n16525 ;
  assign n16561 = \pi0054  & ~n16560 ;
  assign n16562 = ~\pi0074  & n16561 ;
  assign n16563 = ~n16559 & n16562 ;
  assign n16564 = ~n16558 & ~n16563 ;
  assign n16565 = ~n16553 & n16564 ;
  assign n16566 = \pi0074  & ~n16318 ;
  assign n16567 = ~n16315 & n16566 ;
  assign n16568 = \pi0055  & ~n16567 ;
  assign n16569 = n8601 & n10134 ;
  assign n16570 = n10182 & n16569 ;
  assign n16571 = \pi0150  & \pi0232  ;
  assign n16572 = n6706 & n16571 ;
  assign n16573 = ~\pi0092  & n16572 ;
  assign n16574 = n10176 & n16573 ;
  assign n16575 = n10173 & n16574 ;
  assign n16576 = n16570 & ~n16575 ;
  assign n16577 = ~\pi0074  & ~n16318 ;
  assign n16578 = ~n16315 & n16577 ;
  assign n16579 = ~n16322 & n16578 ;
  assign n16580 = ~n16576 & n16579 ;
  assign n16581 = n16568 & ~n16580 ;
  assign n16582 = n1292 & ~n16581 ;
  assign n16583 = n16334 & n16582 ;
  assign n16584 = ~n16565 & n16583 ;
  assign n16585 = ~n16335 & ~n16584 ;
  assign n16586 = ~n1292 & ~n16323 ;
  assign n16587 = ~n16318 & n16586 ;
  assign n16588 = ~n16315 & n16587 ;
  assign n16589 = n2467 & ~n16588 ;
  assign n16590 = ~\pi0074  & ~n16322 ;
  assign n16591 = ~n16318 & n16590 ;
  assign n16592 = ~n16315 & n16591 ;
  assign n16593 = ~\pi0150  & ~\pi0165  ;
  assign n16594 = ~\pi0054  & ~\pi0150  ;
  assign n16595 = ~n16593 & ~n16594 ;
  assign n16596 = n8640 & n16595 ;
  assign n16597 = n1259 & ~n16596 ;
  assign n16598 = n1249 & n16597 ;
  assign n16599 = n8410 & n16598 ;
  assign n16600 = n16592 & ~n16599 ;
  assign n16601 = n16568 & ~n16600 ;
  assign n16602 = n1292 & ~n16601 ;
  assign n16603 = n16589 & ~n16602 ;
  assign n16604 = ~\pi0173  & \pi0190  ;
  assign n16605 = ~\pi0040  & n16604 ;
  assign n16606 = n10414 & n16605 ;
  assign n16607 = n1618 & n16606 ;
  assign n16608 = ~n10899 & n16607 ;
  assign n16609 = ~\pi0190  & n6706 ;
  assign n16610 = ~\pi0173  & n2575 ;
  assign n16611 = n2575 & n10937 ;
  assign n16612 = n10319 & n16611 ;
  assign n16613 = ~n16610 & ~n16612 ;
  assign n16614 = n16609 & ~n16613 ;
  assign n16615 = \pi0185  & ~n16614 ;
  assign n16616 = ~n16608 & n16615 ;
  assign n16617 = n10923 & ~n10929 ;
  assign n16618 = ~\pi0173  & \pi0185  ;
  assign n16619 = ~n16608 & n16618 ;
  assign n16620 = ~n16617 & n16619 ;
  assign n16621 = ~n16616 & ~n16620 ;
  assign n16622 = ~n10943 & ~n10944 ;
  assign n16623 = ~\pi0173  & n10903 ;
  assign n16624 = ~n1864 & n16623 ;
  assign n16625 = ~n10901 & n16624 ;
  assign n16626 = ~n16622 & ~n16625 ;
  assign n16627 = ~\pi0190  & ~n16626 ;
  assign n16628 = \pi0173  & ~n6975 ;
  assign n16629 = ~n10904 & n16628 ;
  assign n16630 = ~\pi0070  & n16628 ;
  assign n16631 = ~n10952 & n16630 ;
  assign n16632 = ~n16629 & ~n16631 ;
  assign n16633 = \pi0190  & n16632 ;
  assign n16634 = n10956 & n16633 ;
  assign n16635 = ~\pi0185  & ~n16634 ;
  assign n16636 = ~n16627 & n16635 ;
  assign n16637 = n16621 & ~n16636 ;
  assign n16638 = ~n6706 & n10904 ;
  assign n16639 = ~n10901 & n16638 ;
  assign n16640 = ~\pi0299  & ~n16639 ;
  assign n16641 = n10570 & ~n10914 ;
  assign n16642 = ~n10913 & n16641 ;
  assign n16643 = \pi0232  & ~n16642 ;
  assign n16644 = n16640 & n16643 ;
  assign n16645 = ~n16637 & n16644 ;
  assign n16646 = ~\pi0151  & n10903 ;
  assign n16647 = ~n1864 & n16646 ;
  assign n16648 = ~n11015 & n16647 ;
  assign n16649 = ~n14576 & ~n16648 ;
  assign n16650 = ~\pi0150  & n16352 ;
  assign n16651 = ~n16649 & n16650 ;
  assign n16652 = ~n10901 & n16647 ;
  assign n16653 = ~n11012 & ~n16652 ;
  assign n16654 = ~\pi0150  & ~\pi0168  ;
  assign n16655 = ~n16653 & n16654 ;
  assign n16656 = ~n16651 & ~n16655 ;
  assign n16657 = ~n14538 & ~n14546 ;
  assign n16658 = ~n6706 & ~n16657 ;
  assign n16659 = ~\pi0040  & \pi0150  ;
  assign n16660 = n10414 & n16659 ;
  assign n16661 = \pi0299  & ~n16660 ;
  assign n16662 = ~\pi0151  & ~\pi0168  ;
  assign n16663 = ~n10929 & n16662 ;
  assign n16664 = n10923 & n16663 ;
  assign n16665 = ~\pi0151  & \pi0168  ;
  assign n16666 = n1618 & n16665 ;
  assign n16667 = ~n10899 & n16666 ;
  assign n16668 = n10937 & n16337 ;
  assign n16669 = n10319 & n16668 ;
  assign n16670 = \pi0299  & ~n16669 ;
  assign n16671 = ~n16667 & n16670 ;
  assign n16672 = ~n16664 & n16671 ;
  assign n16673 = ~n16661 & ~n16672 ;
  assign n16674 = \pi0232  & ~n16673 ;
  assign n16675 = ~n16658 & n16674 ;
  assign n16676 = n16656 & n16675 ;
  assign n16677 = ~n6684 & ~n10914 ;
  assign n16678 = ~n10913 & n16677 ;
  assign n16679 = ~\pi0232  & ~n10904 ;
  assign n16680 = ~\pi0232  & n10900 ;
  assign n16681 = ~n10892 & n16680 ;
  assign n16682 = ~n16679 & ~n16681 ;
  assign n16683 = ~n16678 & ~n16682 ;
  assign n16684 = n1288 & ~n16683 ;
  assign n16685 = ~n16676 & n16684 ;
  assign n16686 = ~n16645 & n16685 ;
  assign n16687 = n6954 & ~n15475 ;
  assign n16688 = \pi0039  & n16687 ;
  assign n16689 = ~n11040 & ~n16688 ;
  assign n16690 = n6948 & n16477 ;
  assign n16691 = ~\pi0178  & ~\pi0190  ;
  assign n16692 = n6954 & n16691 ;
  assign n16693 = ~n16690 & ~n16692 ;
  assign n16694 = n6714 & n6954 ;
  assign n16695 = n8790 & n16473 ;
  assign n16696 = ~n16694 & ~n16695 ;
  assign n16697 = n16693 & n16696 ;
  assign n16698 = n6769 & n16483 ;
  assign n16699 = n6714 & n16483 ;
  assign n16700 = n6954 & n16699 ;
  assign n16701 = ~n16698 & ~n16700 ;
  assign n16702 = ~n16697 & ~n16701 ;
  assign n16703 = ~\pi0038  & n16702 ;
  assign n16704 = ~\pi0168  & ~n11048 ;
  assign n16705 = ~\pi0157  & ~\pi0168  ;
  assign n16706 = ~\pi0157  & n1696 ;
  assign n16707 = n11592 & n16706 ;
  assign n16708 = ~n16705 & ~n16707 ;
  assign n16709 = ~n16704 & ~n16708 ;
  assign n16710 = \pi0232  & ~n16694 ;
  assign n16711 = \pi0157  & ~\pi0168  ;
  assign n16712 = n6743 & n16711 ;
  assign n16713 = n6948 & n16712 ;
  assign n16714 = n16710 & ~n16713 ;
  assign n16715 = ~n16709 & n16714 ;
  assign n16716 = \pi0232  & ~n11062 ;
  assign n16717 = ~\pi0038  & ~n16716 ;
  assign n16718 = ~n16715 & n16717 ;
  assign n16719 = ~n16703 & ~n16718 ;
  assign n16720 = ~n16689 & ~n16719 ;
  assign n16721 = n2364 & ~n16464 ;
  assign n16722 = ~n16720 & n16721 ;
  assign n16723 = ~n16686 & n16722 ;
  assign n16724 = n11470 & ~n16526 ;
  assign n16725 = n16520 & ~n16724 ;
  assign n16726 = \pi0038  & ~\pi0100  ;
  assign n16727 = ~n16525 & n16726 ;
  assign n16728 = ~n16448 & ~n16727 ;
  assign n16729 = n2364 & n16728 ;
  assign n16730 = ~n16725 & n16729 ;
  assign n16731 = ~\pi0100  & ~n16526 ;
  assign n16732 = n10093 & ~n16530 ;
  assign n16733 = n1259 & n16732 ;
  assign n16734 = n1249 & n16733 ;
  assign n16735 = n1281 & n16734 ;
  assign n16736 = n16731 & ~n16735 ;
  assign n16737 = n6895 & n16736 ;
  assign n16738 = \pi0100  & n6895 ;
  assign n16739 = ~n16520 & n16738 ;
  assign n16740 = ~n16737 & ~n16739 ;
  assign n16741 = ~n16559 & n16561 ;
  assign n16742 = ~n16540 & ~n16741 ;
  assign n16743 = n16740 & n16742 ;
  assign n16744 = ~n16730 & n16743 ;
  assign n16745 = ~n16723 & n16744 ;
  assign n16746 = \pi0054  & n16560 ;
  assign n16747 = \pi0054  & ~n16510 ;
  assign n16748 = n16555 & n16747 ;
  assign n16749 = ~n16746 & ~n16748 ;
  assign n16750 = ~\pi0074  & n16749 ;
  assign n16751 = ~n16745 & n16750 ;
  assign n16752 = ~n16558 & n16589 ;
  assign n16753 = ~n16751 & n16752 ;
  assign n16754 = ~n16603 & ~n16753 ;
  assign n16755 = ~\pi0118  & ~n16333 ;
  assign n16756 = n16754 & n16755 ;
  assign n16757 = ~\pi0034  & ~\pi0079  ;
  assign n16758 = n11506 & n16757 ;
  assign n16759 = ~n16756 & ~n16758 ;
  assign n16760 = n16585 & n16759 ;
  assign n16761 = ~\pi0118  & ~n11101 ;
  assign n16762 = ~n16329 & ~n16333 ;
  assign n16763 = ~n16333 & n16582 ;
  assign n16764 = ~n16565 & n16763 ;
  assign n16765 = ~n16762 & ~n16764 ;
  assign n16766 = n16761 & ~n16765 ;
  assign n16767 = ~n16333 & ~n16761 ;
  assign n16768 = n16754 & n16767 ;
  assign n16769 = n16758 & ~n16768 ;
  assign n16770 = ~n16766 & n16769 ;
  assign n16771 = ~n16760 & ~n16770 ;
  assign n16772 = \pi0128  & \pi0228  ;
  assign n16773 = ~n12970 & n16772 ;
  assign n16774 = ~\pi0087  & ~n16772 ;
  assign n16775 = ~n6859 & n16774 ;
  assign n16776 = ~n16448 & ~n16775 ;
  assign n16777 = \pi0075  & n2362 ;
  assign n16778 = n1259 & n16777 ;
  assign n16779 = n1249 & n16778 ;
  assign n16780 = n6858 & n16779 ;
  assign n16781 = ~\pi0100  & n16772 ;
  assign n16782 = \pi0075  & n16772 ;
  assign n16783 = ~\pi0092  & ~n16782 ;
  assign n16784 = ~n16781 & n16783 ;
  assign n16785 = ~n16780 & n16784 ;
  assign n16786 = ~n16776 & n16785 ;
  assign n16787 = \pi0087  & ~n16772 ;
  assign n16788 = ~\pi0075  & ~n16787 ;
  assign n16789 = n16783 & ~n16788 ;
  assign n16790 = ~n16780 & n16789 ;
  assign n16791 = \pi0092  & ~n16772 ;
  assign n16792 = ~n8495 & n16791 ;
  assign n16793 = n12970 & ~n16792 ;
  assign n16794 = ~n16790 & n16793 ;
  assign n16795 = ~n16786 & n16794 ;
  assign n16796 = n1696 & ~n6770 ;
  assign n16797 = ~n2165 & n3058 ;
  assign n16798 = n1259 & n16797 ;
  assign n16799 = n1249 & n16798 ;
  assign n16800 = n6920 & n16799 ;
  assign n16801 = n16796 & n16800 ;
  assign n16802 = n2256 & ~n2352 ;
  assign n16803 = n1259 & n16802 ;
  assign n16804 = n1249 & n16803 ;
  assign n16805 = n6920 & n16804 ;
  assign n16806 = n15374 & n16805 ;
  assign n16807 = ~n16801 & ~n16806 ;
  assign n16808 = n9627 & ~n16807 ;
  assign n16809 = n1383 & n8402 ;
  assign n16810 = n1278 & n8402 ;
  assign n16811 = ~n7069 & n16810 ;
  assign n16812 = ~n16809 & ~n16811 ;
  assign n16813 = ~n16808 & n16812 ;
  assign n16814 = ~\pi0299  & n7100 ;
  assign n16815 = \pi0299  & n7162 ;
  assign n16816 = ~n16814 & ~n16815 ;
  assign n16817 = n8640 & ~n16816 ;
  assign n16818 = \pi0109  & ~n16817 ;
  assign n16819 = \pi0086  & ~n1696 ;
  assign n16820 = ~n1696 & n14002 ;
  assign n16821 = n1542 & n16820 ;
  assign n16822 = ~n16819 & ~n16821 ;
  assign n16823 = ~n7038 & ~n16822 ;
  assign n16824 = ~n16818 & ~n16823 ;
  assign n16825 = ~n7114 & n8640 ;
  assign n16826 = ~n16816 & n16825 ;
  assign n16827 = ~n1325 & ~n16817 ;
  assign n16828 = ~n1319 & n16818 ;
  assign n16829 = ~n16827 & ~n16828 ;
  assign n16830 = ~n16826 & n16829 ;
  assign n16831 = ~n16824 & n16830 ;
  assign n16832 = ~\pi0097  & n1574 ;
  assign n16833 = n1468 & n11813 ;
  assign n16834 = ~\pi0086  & ~n16833 ;
  assign n16835 = ~\pi0097  & ~n15939 ;
  assign n16836 = n16834 & n16835 ;
  assign n16837 = ~n16832 & ~n16836 ;
  assign n16838 = ~\pi0046  & \pi1091  ;
  assign n16839 = n1689 & n16838 ;
  assign n16840 = n1688 & n16839 ;
  assign n16841 = ~n16826 & n16840 ;
  assign n16842 = ~n1678 & n16841 ;
  assign n16843 = n16829 & n16842 ;
  assign n16844 = n16837 & n16843 ;
  assign n16845 = ~n16831 & ~n16844 ;
  assign n16846 = ~\pi0091  & ~n1383 ;
  assign n16847 = ~n16808 & n16846 ;
  assign n16848 = n16845 & n16847 ;
  assign n16849 = ~n16813 & ~n16848 ;
  assign n16850 = n8453 & n16794 ;
  assign n16851 = n16849 & n16850 ;
  assign n16852 = ~n16795 & ~n16851 ;
  assign n16853 = ~n16773 & n16852 ;
  assign n16854 = ~n8496 & n8696 ;
  assign n16855 = ~\pi0120  & ~\pi1093  ;
  assign n16856 = ~n8496 & n16855 ;
  assign n16857 = ~n9250 & ~n16856 ;
  assign n16858 = ~n16854 & n16857 ;
  assign n16859 = \pi0950  & n1281 ;
  assign n16860 = n1260 & n16859 ;
  assign n16861 = \pi0951  & \pi0982  ;
  assign n16862 = n14727 & n16861 ;
  assign n16863 = ~\pi1091  & n16862 ;
  assign n16864 = ~n1686 & n8587 ;
  assign n16865 = ~\pi0120  & n16864 ;
  assign n16866 = ~n16863 & n16865 ;
  assign n16867 = ~n6808 & n16866 ;
  assign n16868 = n16860 & n16867 ;
  assign n16869 = \pi0120  & \pi1091  ;
  assign n16870 = n1259 & n16869 ;
  assign n16871 = n1249 & n16870 ;
  assign n16872 = n8664 & n16871 ;
  assign n16873 = \pi1092  & n16861 ;
  assign n16874 = n6703 & n16873 ;
  assign n16875 = ~\pi0120  & ~n16863 ;
  assign n16876 = ~n16874 & n16875 ;
  assign n16877 = \pi0100  & ~n16876 ;
  assign n16878 = ~n16872 & n16877 ;
  assign n16879 = ~n16868 & n16878 ;
  assign n16880 = \pi0100  & ~n9635 ;
  assign n16881 = \pi0100  & n8640 ;
  assign n16882 = n8639 & n16881 ;
  assign n16883 = ~n16880 & ~n16882 ;
  assign n16884 = ~\pi0038  & n16883 ;
  assign n16885 = ~n16879 & n16884 ;
  assign n16886 = ~\pi0120  & ~n16862 ;
  assign n16887 = n8640 & n16886 ;
  assign n16888 = n8639 & n16887 ;
  assign n16889 = ~n8666 & n16886 ;
  assign n16890 = ~n16888 & ~n16889 ;
  assign n16891 = ~n16885 & n16890 ;
  assign n16892 = ~n2327 & ~n16891 ;
  assign n16893 = \pi0075  & n2342 ;
  assign n16894 = \pi0075  & ~\pi0120  ;
  assign n16895 = ~n16862 & n16894 ;
  assign n16896 = ~n16893 & ~n16895 ;
  assign n16897 = n2342 & ~n16888 ;
  assign n16898 = ~n16896 & ~n16897 ;
  assign n16899 = ~n8641 & ~n16896 ;
  assign n16900 = ~n16898 & ~n16899 ;
  assign n16901 = ~\pi0024  & n7203 ;
  assign n16902 = ~\pi0072  & ~\pi0122  ;
  assign n16903 = n1688 & n16902 ;
  assign n16904 = n16901 & n16903 ;
  assign n16905 = n1627 & n16904 ;
  assign n16906 = n1319 & n16905 ;
  assign n16907 = ~n6808 & n16875 ;
  assign n16908 = n16906 & n16907 ;
  assign n16909 = ~n16876 & ~n16908 ;
  assign n16910 = \pi0120  & n8798 ;
  assign n16911 = n8801 & n16910 ;
  assign n16912 = n7207 & n16911 ;
  assign n16913 = ~n16898 & ~n16912 ;
  assign n16914 = n16909 & n16913 ;
  assign n16915 = ~n16900 & ~n16914 ;
  assign n16916 = ~\pi0087  & ~n16915 ;
  assign n16917 = ~n16892 & n16916 ;
  assign n16918 = n8496 & n16915 ;
  assign n16919 = ~n2328 & n16886 ;
  assign n16920 = \pi0087  & ~n16919 ;
  assign n16921 = \pi0120  & ~n8543 ;
  assign n16922 = ~n8630 & n16921 ;
  assign n16923 = \pi0120  & n8543 ;
  assign n16924 = ~n9048 & n16923 ;
  assign n16925 = n2328 & ~n16924 ;
  assign n16926 = ~n16922 & n16925 ;
  assign n16927 = ~n1686 & ~n6810 ;
  assign n16928 = \pi0950  & n16927 ;
  assign n16929 = n1281 & n16928 ;
  assign n16930 = n1260 & n16929 ;
  assign n16931 = n16874 & ~n16930 ;
  assign n16932 = n1281 & n14707 ;
  assign n16933 = n1260 & n16932 ;
  assign n16934 = n16863 & ~n16933 ;
  assign n16935 = ~n16931 & ~n16934 ;
  assign n16936 = ~\pi0120  & ~n16935 ;
  assign n16937 = n16926 & ~n16936 ;
  assign n16938 = n16920 & ~n16937 ;
  assign n16939 = n15835 & ~n16938 ;
  assign n16940 = ~n16918 & ~n16939 ;
  assign n16941 = ~n16917 & ~n16940 ;
  assign n16942 = n8587 & n16873 ;
  assign n16943 = n8742 & ~n12033 ;
  assign n16944 = n16942 & ~n16943 ;
  assign n16945 = \pi0122  & \pi1092  ;
  assign n16946 = n16861 & n16945 ;
  assign n16947 = \pi0829  & n16946 ;
  assign n16948 = \pi0950  & n8592 ;
  assign n16949 = ~n8581 & n16948 ;
  assign n16950 = n16947 & ~n16949 ;
  assign n16951 = n1273 & n13028 ;
  assign n16952 = n1277 & n15912 ;
  assign n16953 = n16951 & n16952 ;
  assign n16954 = n1542 & n16953 ;
  assign n16955 = ~n8559 & n16954 ;
  assign n16956 = n16947 & ~n16955 ;
  assign n16957 = n8719 & n16956 ;
  assign n16958 = ~n16950 & ~n16957 ;
  assign n16959 = n8719 & ~n16955 ;
  assign n16960 = \pi0824  & n16949 ;
  assign n16961 = ~n16959 & n16960 ;
  assign n16962 = ~\pi0829  & \pi1092  ;
  assign n16963 = n16861 & n16962 ;
  assign n16964 = ~n16961 & n16963 ;
  assign n16965 = n16958 & ~n16964 ;
  assign n16966 = ~n16944 & n16965 ;
  assign n16967 = n8782 & ~n16966 ;
  assign n16968 = \pi1091  & n1686 ;
  assign n16969 = n16862 & n16968 ;
  assign n16970 = n16863 & ~n16961 ;
  assign n16971 = ~\pi0120  & ~n16970 ;
  assign n16972 = ~n16969 & n16971 ;
  assign n16973 = ~n16967 & n16972 ;
  assign n16974 = ~n8586 & n12045 ;
  assign n16975 = n8593 & n8594 ;
  assign n16976 = ~n8578 & n16975 ;
  assign n16977 = ~\pi1093  & ~n16976 ;
  assign n16978 = ~n16974 & n16977 ;
  assign n16979 = \pi0120  & ~n16978 ;
  assign n16980 = ~\pi0039  & ~n16979 ;
  assign n16981 = n8743 & ~n12033 ;
  assign n16982 = n8593 & n8752 ;
  assign n16983 = ~n8578 & n16982 ;
  assign n16984 = ~\pi0122  & ~n16983 ;
  assign n16985 = ~n16981 & n16984 ;
  assign n16986 = n6811 & n8593 ;
  assign n16987 = ~n8578 & n16986 ;
  assign n16988 = \pi0122  & ~n16987 ;
  assign n16989 = ~\pi0833  & \pi0957  ;
  assign n16990 = ~n16988 & ~n16989 ;
  assign n16991 = ~n8578 & n9014 ;
  assign n16992 = n8543 & ~n16991 ;
  assign n16993 = n16990 & ~n16992 ;
  assign n16994 = ~n16985 & n16993 ;
  assign n16995 = ~\pi1091  & n9014 ;
  assign n16996 = ~n8578 & n16995 ;
  assign n16997 = \pi1093  & ~n16996 ;
  assign n16998 = ~\pi0039  & n16997 ;
  assign n16999 = ~n16994 & n16998 ;
  assign n17000 = ~n16980 & ~n16999 ;
  assign n17001 = ~n16973 & ~n17000 ;
  assign n17002 = \pi0039  & ~n16886 ;
  assign n17003 = ~n9625 & n17002 ;
  assign n17004 = ~n16891 & ~n17003 ;
  assign n17005 = ~n16940 & n17004 ;
  assign n17006 = ~n17001 & n17005 ;
  assign n17007 = ~n16941 & ~n17006 ;
  assign n17008 = n9250 & n17007 ;
  assign n17009 = ~n16858 & ~n17008 ;
  assign n17010 = n8543 & ~n8695 ;
  assign n17011 = ~n8617 & n17010 ;
  assign n17012 = n2328 & ~n17011 ;
  assign n17013 = ~n9046 & n17012 ;
  assign n17014 = ~n16926 & ~n17013 ;
  assign n17015 = ~\pi0120  & n16874 ;
  assign n17016 = ~n16930 & n17015 ;
  assign n17017 = ~\pi0120  & ~n8695 ;
  assign n17018 = n16863 & n17017 ;
  assign n17019 = n16863 & n17018 ;
  assign n17020 = ~n16933 & n17019 ;
  assign n17021 = ~n17016 & ~n17020 ;
  assign n17022 = ~n17014 & n17021 ;
  assign n17023 = ~n2328 & n8696 ;
  assign n17024 = n16920 & ~n17023 ;
  assign n17025 = ~n17022 & n17024 ;
  assign n17026 = ~\pi0075  & n17025 ;
  assign n17027 = n16873 & n17010 ;
  assign n17028 = ~n16961 & n17027 ;
  assign n17029 = ~\pi0039  & ~n16969 ;
  assign n17030 = ~n17028 & n17029 ;
  assign n17031 = ~n16967 & n17030 ;
  assign n17032 = ~\pi0120  & n17031 ;
  assign n17033 = ~n6703 & ~n17010 ;
  assign n17034 = ~n6703 & n9014 ;
  assign n17035 = ~n8578 & n17034 ;
  assign n17036 = ~n17033 & ~n17035 ;
  assign n17037 = ~n16991 & n17010 ;
  assign n17038 = n16990 & ~n17037 ;
  assign n17039 = ~n16985 & n17038 ;
  assign n17040 = n17036 & ~n17039 ;
  assign n17041 = ~\pi0039  & n16979 ;
  assign n17042 = ~n17040 & n17041 ;
  assign n17043 = ~n8696 & ~n16855 ;
  assign n17044 = ~\pi0100  & ~n16886 ;
  assign n17045 = n17043 & n17044 ;
  assign n17046 = ~n2327 & ~n17045 ;
  assign n17047 = ~n8695 & n16863 ;
  assign n17048 = n1259 & ~n17047 ;
  assign n17049 = n1249 & n17048 ;
  assign n17050 = n6920 & n17049 ;
  assign n17051 = n1688 & n17050 ;
  assign n17052 = ~n16874 & ~n17047 ;
  assign n17053 = ~\pi0120  & ~n6736 ;
  assign n17054 = ~n17052 & n17053 ;
  assign n17055 = ~n17051 & n17054 ;
  assign n17056 = \pi0120  & ~n8696 ;
  assign n17057 = ~n6736 & n17056 ;
  assign n17058 = ~n8790 & n17057 ;
  assign n17059 = n6736 & n17043 ;
  assign n17060 = ~n16886 & n17059 ;
  assign n17061 = ~n17058 & ~n17060 ;
  assign n17062 = ~n17055 & n17061 ;
  assign n17063 = ~n6732 & ~n17062 ;
  assign n17064 = ~\pi0120  & ~n6706 ;
  assign n17065 = ~n6713 & n17064 ;
  assign n17066 = ~n17052 & n17065 ;
  assign n17067 = ~n17051 & n17066 ;
  assign n17068 = n6714 & n17056 ;
  assign n17069 = ~n8790 & n17068 ;
  assign n17070 = ~n16886 & n17043 ;
  assign n17071 = ~n6714 & n17070 ;
  assign n17072 = n8684 & ~n17071 ;
  assign n17073 = ~n17069 & n17072 ;
  assign n17074 = ~n17067 & n17073 ;
  assign n17075 = ~n8685 & ~n17074 ;
  assign n17076 = ~n17063 & ~n17075 ;
  assign n17077 = ~n8684 & n8696 ;
  assign n17078 = \pi0299  & ~n17077 ;
  assign n17079 = ~n8684 & n16886 ;
  assign n17080 = n17078 & ~n17079 ;
  assign n17081 = ~n17076 & n17080 ;
  assign n17082 = ~n6761 & ~n17062 ;
  assign n17083 = ~n6761 & n8701 ;
  assign n17084 = n8701 & ~n17071 ;
  assign n17085 = ~n17069 & n17084 ;
  assign n17086 = ~n17067 & n17085 ;
  assign n17087 = ~n17083 & ~n17086 ;
  assign n17088 = ~n17082 & ~n17087 ;
  assign n17089 = ~\pi0299  & n8701 ;
  assign n17090 = ~\pi0299  & ~n16886 ;
  assign n17091 = n17043 & n17090 ;
  assign n17092 = ~n17089 & ~n17091 ;
  assign n17093 = ~n17088 & ~n17092 ;
  assign n17094 = \pi0039  & ~n17093 ;
  assign n17095 = ~n17081 & n17094 ;
  assign n17096 = ~n17046 & ~n17095 ;
  assign n17097 = ~n17042 & n17096 ;
  assign n17098 = ~n17032 & n17097 ;
  assign n17099 = n16726 & ~n16886 ;
  assign n17100 = n17043 & n17099 ;
  assign n17101 = \pi0228  & ~n8641 ;
  assign n17102 = ~n8641 & n8666 ;
  assign n17103 = n1288 & ~n17070 ;
  assign n17104 = ~n17102 & ~n17103 ;
  assign n17105 = ~n17101 & ~n17104 ;
  assign n17106 = ~n6808 & n16864 ;
  assign n17107 = ~n17047 & n17106 ;
  assign n17108 = n16860 & n17107 ;
  assign n17109 = ~\pi0120  & ~n17052 ;
  assign n17110 = ~n17108 & n17109 ;
  assign n17111 = \pi1091  & n1259 ;
  assign n17112 = n1249 & n17111 ;
  assign n17113 = n8664 & n17112 ;
  assign n17114 = n17056 & ~n17113 ;
  assign n17115 = ~n17104 & ~n17114 ;
  assign n17116 = ~n17110 & n17115 ;
  assign n17117 = ~n17105 & ~n17116 ;
  assign n17118 = \pi0100  & n1288 ;
  assign n17119 = \pi0100  & ~n16886 ;
  assign n17120 = n17043 & n17119 ;
  assign n17121 = ~n17118 & ~n17120 ;
  assign n17122 = n17117 & ~n17121 ;
  assign n17123 = ~n17100 & ~n17122 ;
  assign n17124 = ~n17098 & n17123 ;
  assign n17125 = n16291 & ~n17124 ;
  assign n17126 = ~n17026 & ~n17125 ;
  assign n17127 = \pi0075  & ~n16886 ;
  assign n17128 = n17043 & n17127 ;
  assign n17129 = ~n2347 & ~n17128 ;
  assign n17130 = n8641 & ~n17070 ;
  assign n17131 = ~n17129 & ~n17130 ;
  assign n17132 = n16033 & ~n16886 ;
  assign n17133 = n17043 & n17132 ;
  assign n17134 = n8496 & ~n17133 ;
  assign n17135 = ~n17131 & n17134 ;
  assign n17136 = ~n6808 & n16906 ;
  assign n17137 = n17015 & ~n17136 ;
  assign n17138 = ~n8641 & ~n17018 ;
  assign n17139 = ~n17137 & n17138 ;
  assign n17140 = \pi1093  & n8695 ;
  assign n17141 = \pi0120  & ~\pi1091  ;
  assign n17142 = ~n17140 & n17141 ;
  assign n17143 = ~n16869 & ~n17142 ;
  assign n17144 = n8651 & ~n17142 ;
  assign n17145 = n7207 & n17144 ;
  assign n17146 = ~n17143 & ~n17145 ;
  assign n17147 = n17134 & ~n17146 ;
  assign n17148 = n17139 & n17147 ;
  assign n17149 = ~n17135 & ~n17148 ;
  assign n17150 = ~n17008 & ~n17149 ;
  assign n17151 = n17126 & n17150 ;
  assign n17152 = ~n17009 & ~n17151 ;
  assign n17153 = ~\pi0031  & ~\pi0080  ;
  assign n17154 = \pi0818  & n17153 ;
  assign n17155 = n9250 & ~n16855 ;
  assign n17156 = n17154 & n17155 ;
  assign n17157 = ~n16855 & n17154 ;
  assign n17158 = ~n8696 & n17157 ;
  assign n17159 = ~n17156 & ~n17158 ;
  assign n17160 = ~n9948 & n17159 ;
  assign n17161 = ~n9250 & ~n17043 ;
  assign n17162 = ~n16886 & ~n17161 ;
  assign n17163 = n17160 & ~n17162 ;
  assign n17164 = ~\pi0120  & ~n8496 ;
  assign n17165 = ~n16862 & n17164 ;
  assign n17166 = n10003 & ~n17165 ;
  assign n17167 = ~n17154 & n17166 ;
  assign n17168 = ~n17163 & n17167 ;
  assign n17169 = n17152 & n17168 ;
  assign n17170 = ~\pi1091  & n8695 ;
  assign n17171 = ~\pi0120  & \pi1093  ;
  assign n17172 = ~n17170 & n17171 ;
  assign n17173 = ~n8641 & ~n17172 ;
  assign n17174 = n8649 & n8799 ;
  assign n17175 = ~n6808 & n17174 ;
  assign n17176 = ~n8641 & n17175 ;
  assign n17177 = n7207 & n17176 ;
  assign n17178 = ~n17173 & ~n17177 ;
  assign n17179 = ~n17146 & ~n17178 ;
  assign n17180 = \pi0075  & ~n16855 ;
  assign n17181 = ~n8696 & n17180 ;
  assign n17182 = ~n16893 & ~n17181 ;
  assign n17183 = n8641 & ~n17043 ;
  assign n17184 = ~n17182 & ~n17183 ;
  assign n17185 = ~n17179 & n17184 ;
  assign n17186 = ~n2342 & n17180 ;
  assign n17187 = ~n8696 & n17186 ;
  assign n17188 = n8496 & ~n17187 ;
  assign n17189 = ~n17185 & n17188 ;
  assign n17190 = ~n16854 & ~n17189 ;
  assign n17191 = \pi0299  & n8684 ;
  assign n17192 = \pi0299  & ~n16855 ;
  assign n17193 = ~n8696 & n17192 ;
  assign n17194 = ~n17191 & ~n17193 ;
  assign n17195 = \pi0039  & n17194 ;
  assign n17196 = ~n8790 & n17056 ;
  assign n17197 = ~n6732 & ~n6736 ;
  assign n17198 = n17196 & n17197 ;
  assign n17199 = n1259 & n8675 ;
  assign n17200 = n1249 & n17199 ;
  assign n17201 = n6920 & n17200 ;
  assign n17202 = n8799 & n17201 ;
  assign n17203 = n17172 & n17197 ;
  assign n17204 = ~n17202 & n17203 ;
  assign n17205 = ~n17198 & ~n17204 ;
  assign n17206 = ~n6732 & n17059 ;
  assign n17207 = \pi0039  & ~n17206 ;
  assign n17208 = n17205 & n17207 ;
  assign n17209 = ~n6714 & n17043 ;
  assign n17210 = n6732 & n17209 ;
  assign n17211 = n8684 & ~n17210 ;
  assign n17212 = n6714 & n6732 ;
  assign n17213 = n17196 & n17212 ;
  assign n17214 = n17172 & n17212 ;
  assign n17215 = ~n17202 & n17214 ;
  assign n17216 = ~n17213 & ~n17215 ;
  assign n17217 = n17211 & n17216 ;
  assign n17218 = n17208 & n17217 ;
  assign n17219 = ~n17195 & ~n17218 ;
  assign n17220 = ~\pi0299  & ~n16855 ;
  assign n17221 = ~n8696 & n17220 ;
  assign n17222 = ~n17089 & ~n17221 ;
  assign n17223 = ~\pi0038  & n17222 ;
  assign n17224 = n6714 & n6761 ;
  assign n17225 = n17196 & n17224 ;
  assign n17226 = n17172 & n17224 ;
  assign n17227 = ~n17202 & n17226 ;
  assign n17228 = ~n17225 & ~n17227 ;
  assign n17229 = ~n6761 & n17059 ;
  assign n17230 = n6761 & n17209 ;
  assign n17231 = n8701 & ~n17230 ;
  assign n17232 = ~n17229 & n17231 ;
  assign n17233 = n17228 & n17232 ;
  assign n17234 = ~n6736 & ~n6761 ;
  assign n17235 = n17196 & n17234 ;
  assign n17236 = n17172 & n17234 ;
  assign n17237 = ~n17202 & n17236 ;
  assign n17238 = ~n17235 & ~n17237 ;
  assign n17239 = ~\pi0038  & n17238 ;
  assign n17240 = n17233 & n17239 ;
  assign n17241 = ~n17223 & ~n17240 ;
  assign n17242 = ~n17219 & ~n17241 ;
  assign n17243 = \pi0120  & ~\pi1093  ;
  assign n17244 = ~n16976 & n17243 ;
  assign n17245 = ~\pi0039  & ~n17244 ;
  assign n17246 = ~\pi0039  & n12045 ;
  assign n17247 = ~n8586 & n17246 ;
  assign n17248 = ~n17245 & ~n17247 ;
  assign n17249 = ~\pi0038  & ~n17248 ;
  assign n17250 = ~n17242 & ~n17249 ;
  assign n17251 = n17036 & ~n17242 ;
  assign n17252 = ~n17039 & n17251 ;
  assign n17253 = ~n17250 & ~n17252 ;
  assign n17254 = \pi0038  & n8543 ;
  assign n17255 = n8695 & n17254 ;
  assign n17256 = \pi0038  & n16855 ;
  assign n17257 = n16448 & ~n17256 ;
  assign n17258 = ~n17255 & n17257 ;
  assign n17259 = ~n17253 & n17258 ;
  assign n17260 = n1281 & n8801 ;
  assign n17261 = n1260 & n17260 ;
  assign n17262 = \pi1093  & n8666 ;
  assign n17263 = ~n8641 & n17262 ;
  assign n17264 = n17261 & n17263 ;
  assign n17265 = \pi0100  & ~n16855 ;
  assign n17266 = ~\pi0087  & n17265 ;
  assign n17267 = ~n8696 & n17266 ;
  assign n17268 = ~n17264 & n17267 ;
  assign n17269 = \pi0087  & ~n16855 ;
  assign n17270 = ~n9039 & n17269 ;
  assign n17271 = ~n9034 & n17270 ;
  assign n17272 = \pi0087  & ~n17023 ;
  assign n17273 = n17271 & n17272 ;
  assign n17274 = ~n17013 & n17273 ;
  assign n17275 = ~n17268 & ~n17274 ;
  assign n17276 = ~n17259 & n17275 ;
  assign n17277 = ~\pi0075  & ~n16854 ;
  assign n17278 = ~n17276 & n17277 ;
  assign n17279 = ~n17190 & ~n17278 ;
  assign n17280 = n16857 & ~n17279 ;
  assign n17281 = ~n8804 & n17180 ;
  assign n17282 = n8496 & ~n17281 ;
  assign n17283 = ~n16856 & ~n17282 ;
  assign n17284 = n6736 & ~n6761 ;
  assign n17285 = n8701 & ~n17284 ;
  assign n17286 = \pi1093  & n6761 ;
  assign n17287 = ~n6714 & n17286 ;
  assign n17288 = n1696 & ~n17287 ;
  assign n17289 = n17285 & n17288 ;
  assign n17290 = n6921 & n17289 ;
  assign n17291 = n17220 & ~n17290 ;
  assign n17292 = ~n6732 & n6736 ;
  assign n17293 = n8684 & ~n17292 ;
  assign n17294 = \pi1093  & n6732 ;
  assign n17295 = ~n6714 & n17294 ;
  assign n17296 = n1696 & ~n17295 ;
  assign n17297 = n17293 & n17296 ;
  assign n17298 = n6921 & n17297 ;
  assign n17299 = n17192 & ~n17298 ;
  assign n17300 = ~n17291 & ~n17299 ;
  assign n17301 = n9627 & n17300 ;
  assign n17302 = ~n17249 & ~n17301 ;
  assign n17303 = n16997 & ~n17301 ;
  assign n17304 = ~n16994 & n17303 ;
  assign n17305 = ~n17302 & ~n17304 ;
  assign n17306 = n17257 & ~n17305 ;
  assign n17307 = ~\pi0120  & n1259 ;
  assign n17308 = n1249 & n17307 ;
  assign n17309 = n17260 & n17308 ;
  assign n17310 = ~n16872 & ~n17309 ;
  assign n17311 = n17102 & ~n17310 ;
  assign n17312 = n17266 & ~n17311 ;
  assign n17313 = ~n17271 & ~n17312 ;
  assign n17314 = ~n17306 & n17313 ;
  assign n17315 = ~\pi0075  & ~n16856 ;
  assign n17316 = ~n17314 & n17315 ;
  assign n17317 = ~n17283 & ~n17316 ;
  assign n17318 = n9250 & ~n17317 ;
  assign n17319 = ~n17280 & ~n17318 ;
  assign n17320 = \pi0120  & n9250 ;
  assign n17321 = ~n17056 & ~n17320 ;
  assign n17322 = n17160 & n17321 ;
  assign n17323 = ~n10003 & ~n17322 ;
  assign n17324 = n10003 & ~n17163 ;
  assign n17325 = ~n17323 & ~n17324 ;
  assign n17326 = n17154 & ~n17325 ;
  assign n17327 = ~n17319 & n17326 ;
  assign n17328 = ~n9948 & ~n10003 ;
  assign n17329 = ~n17322 & n17328 ;
  assign n17330 = ~n9948 & n10003 ;
  assign n17331 = ~n17163 & n17330 ;
  assign n17332 = ~n17329 & ~n17331 ;
  assign n17333 = ~n9250 & ~n16854 ;
  assign n17334 = ~\pi1091  & ~n17140 ;
  assign n17335 = n2342 & ~n17334 ;
  assign n17336 = ~n8641 & n17335 ;
  assign n17337 = ~\pi1091  & n17336 ;
  assign n17338 = n8651 & n17336 ;
  assign n17339 = n7207 & n17338 ;
  assign n17340 = ~n17337 & ~n17339 ;
  assign n17341 = n8640 & n8696 ;
  assign n17342 = n8639 & n17341 ;
  assign n17343 = ~n2342 & n8696 ;
  assign n17344 = \pi0075  & ~n17343 ;
  assign n17345 = ~n17342 & n17344 ;
  assign n17346 = n17340 & n17345 ;
  assign n17347 = n17333 & n17346 ;
  assign n17348 = ~\pi1091  & n17140 ;
  assign n17349 = \pi1091  & ~n6706 ;
  assign n17350 = ~n6713 & n17349 ;
  assign n17351 = ~n17348 & ~n17350 ;
  assign n17352 = n8689 & ~n17351 ;
  assign n17353 = ~n8680 & n17352 ;
  assign n17354 = ~n8682 & ~n17334 ;
  assign n17355 = n8685 & n17354 ;
  assign n17356 = ~n8680 & n17355 ;
  assign n17357 = n17078 & ~n17356 ;
  assign n17358 = ~n17353 & n17357 ;
  assign n17359 = n8705 & ~n17351 ;
  assign n17360 = ~n8680 & n17359 ;
  assign n17361 = n17083 & n17354 ;
  assign n17362 = ~n8680 & n17361 ;
  assign n17363 = n8696 & ~n8701 ;
  assign n17364 = ~\pi0299  & ~n17363 ;
  assign n17365 = ~n17362 & n17364 ;
  assign n17366 = ~n17360 & n17365 ;
  assign n17367 = ~n17358 & ~n17366 ;
  assign n17368 = n9627 & n17367 ;
  assign n17369 = \pi0039  & ~n17367 ;
  assign n17370 = ~\pi0038  & ~n17369 ;
  assign n17371 = ~n16978 & n17370 ;
  assign n17372 = ~n17368 & ~n17371 ;
  assign n17373 = n17036 & ~n17368 ;
  assign n17374 = ~n17039 & n17373 ;
  assign n17375 = ~n17372 & ~n17374 ;
  assign n17376 = ~\pi0100  & ~n17255 ;
  assign n17377 = ~\pi0087  & n17376 ;
  assign n17378 = ~n17375 & n17377 ;
  assign n17379 = ~n17013 & n17272 ;
  assign n17380 = ~n8696 & n9010 ;
  assign n17381 = ~n8669 & n17380 ;
  assign n17382 = ~n17379 & ~n17381 ;
  assign n17383 = ~n17378 & n17382 ;
  assign n17384 = ~\pi0075  & n17333 ;
  assign n17385 = ~n17383 & n17384 ;
  assign n17386 = ~n17347 & ~n17385 ;
  assign n17387 = \pi0039  & n8790 ;
  assign n17388 = n8794 & n17387 ;
  assign n17389 = ~n15448 & ~n16978 ;
  assign n17390 = ~n17388 & ~n17389 ;
  assign n17391 = n16997 & ~n17388 ;
  assign n17392 = ~n16994 & n17391 ;
  assign n17393 = ~n17390 & ~n17392 ;
  assign n17394 = n2362 & ~n17393 ;
  assign n17395 = ~n8805 & ~n9041 ;
  assign n17396 = ~n9011 & n17395 ;
  assign n17397 = ~n17394 & n17396 ;
  assign n17398 = ~n8641 & n16893 ;
  assign n17399 = n8802 & n17398 ;
  assign n17400 = n7207 & n17399 ;
  assign n17401 = n9250 & ~n17164 ;
  assign n17402 = ~n17400 & n17401 ;
  assign n17403 = ~n17397 & n17402 ;
  assign n17404 = ~n8496 & n9250 ;
  assign n17405 = ~n8496 & ~n16855 ;
  assign n17406 = ~n8696 & n17405 ;
  assign n17407 = ~n17404 & ~n17406 ;
  assign n17408 = ~n17403 & n17407 ;
  assign n17409 = n17386 & n17408 ;
  assign n17410 = \pi0120  & ~n17154 ;
  assign n17411 = n17323 & n17410 ;
  assign n17412 = ~n17409 & n17411 ;
  assign n17413 = n17332 & ~n17412 ;
  assign n17414 = ~n17327 & n17413 ;
  assign n17415 = ~n17169 & n17414 ;
  assign n17416 = \pi0163  & n6706 ;
  assign n17417 = \pi0087  & \pi0232  ;
  assign n17418 = n17416 & n17417 ;
  assign n17419 = n1233 & n11809 ;
  assign n17420 = ~\pi0051  & n17419 ;
  assign n17421 = n6706 & ~n17420 ;
  assign n17422 = ~\pi0087  & \pi0232  ;
  assign n17423 = n6706 & n14079 ;
  assign n17424 = ~n17422 & ~n17423 ;
  assign n17425 = \pi0051  & ~\pi0146  ;
  assign n17426 = n6706 & n17425 ;
  assign n17427 = ~\pi0051  & ~\pi0161  ;
  assign n17428 = ~n11365 & ~n17427 ;
  assign n17429 = ~n17426 & n17428 ;
  assign n17430 = ~n17424 & ~n17429 ;
  assign n17431 = n17421 & n17430 ;
  assign n17432 = ~n17418 & ~n17431 ;
  assign n17433 = ~\pi0121  & ~\pi0132  ;
  assign n17434 = ~\pi0126  & n17433 ;
  assign n17435 = ~\pi0134  & ~\pi0135  ;
  assign n17436 = ~\pi0130  & ~\pi0136  ;
  assign n17437 = n17435 & n17436 ;
  assign n17438 = n17434 & n17437 ;
  assign n17439 = ~\pi0125  & ~\pi0133  ;
  assign n17440 = \pi0121  & ~n17439 ;
  assign n17441 = ~\pi0121  & n17439 ;
  assign n17442 = ~n17440 & ~n17441 ;
  assign n17443 = ~n17438 & ~n17442 ;
  assign n17444 = n15926 & n17419 ;
  assign n17445 = ~n17443 & n17444 ;
  assign n17446 = ~n9948 & ~n17445 ;
  assign n17447 = n17432 & n17446 ;
  assign n17448 = \pi0051  & \pi0142  ;
  assign n17449 = n6706 & ~n17448 ;
  assign n17450 = \pi0144  & ~n17449 ;
  assign n17451 = n1568 & n14012 ;
  assign n17452 = n1542 & n17451 ;
  assign n17453 = ~\pi0024  & ~n17452 ;
  assign n17454 = ~\pi0314  & n17453 ;
  assign n17455 = \pi0024  & ~\pi0314  ;
  assign n17456 = ~n14006 & n17455 ;
  assign n17457 = ~n17454 & ~n17456 ;
  assign n17458 = \pi0314  & ~n14006 ;
  assign n17459 = ~\pi0096  & n1322 ;
  assign n17460 = n13001 & n17459 ;
  assign n17461 = ~n17458 & n17460 ;
  assign n17462 = n17457 & n17461 ;
  assign n17463 = ~\pi0051  & \pi0144  ;
  assign n17464 = ~n17462 & n17463 ;
  assign n17465 = ~n17450 & ~n17464 ;
  assign n17466 = n1232 & n1458 ;
  assign n17467 = n1242 & n17466 ;
  assign n17468 = ~\pi0069  & n1244 ;
  assign n17469 = n1567 & n17468 ;
  assign n17470 = n11805 & n17469 ;
  assign n17471 = ~\pi0024  & ~\pi0108  ;
  assign n17472 = n1268 & n17471 ;
  assign n17473 = n1272 & n17472 ;
  assign n17474 = ~\pi0077  & \pi0086  ;
  assign n17475 = n13410 & n17474 ;
  assign n17476 = n17473 & n17475 ;
  assign n17477 = n17470 & n17476 ;
  assign n17478 = n17467 & n17477 ;
  assign n17479 = n17419 & ~n17478 ;
  assign n17480 = n17467 & n17470 ;
  assign n17481 = \pi0024  & ~\pi0108  ;
  assign n17482 = n1268 & n17481 ;
  assign n17483 = n1272 & n17482 ;
  assign n17484 = ~\pi0077  & ~\pi0086  ;
  assign n17485 = \pi0077  & \pi0086  ;
  assign n17486 = ~n17484 & ~n17485 ;
  assign n17487 = n13410 & n17486 ;
  assign n17488 = n17483 & n17487 ;
  assign n17489 = n17480 & n17488 ;
  assign n17490 = n17479 & ~n17489 ;
  assign n17491 = \pi0077  & ~\pi0086  ;
  assign n17492 = ~\pi0096  & \pi0314  ;
  assign n17493 = n13410 & n17492 ;
  assign n17494 = n1322 & n17493 ;
  assign n17495 = n17473 & n17494 ;
  assign n17496 = n17491 & n17495 ;
  assign n17497 = n17480 & n17496 ;
  assign n17498 = n13001 & n17419 ;
  assign n17499 = n17459 & n17498 ;
  assign n17500 = ~n17497 & n17499 ;
  assign n17501 = n17490 & n17500 ;
  assign n17502 = n1329 & n10414 ;
  assign n17503 = ~\pi0051  & n6706 ;
  assign n17504 = ~n17419 & n17503 ;
  assign n17505 = ~n17502 & ~n17504 ;
  assign n17506 = \pi0142  & ~n17505 ;
  assign n17507 = ~\pi0051  & ~n17419 ;
  assign n17508 = ~n1324 & ~n17507 ;
  assign n17509 = n13001 & n17508 ;
  assign n17510 = n17506 & ~n17509 ;
  assign n17511 = ~n17501 & n17510 ;
  assign n17512 = n13001 & n17491 ;
  assign n17513 = n17495 & n17512 ;
  assign n17514 = n17480 & n17513 ;
  assign n17515 = n17420 & ~n17514 ;
  assign n17516 = ~\pi0142  & n6706 ;
  assign n17517 = ~n17515 & n17516 ;
  assign n17518 = n13001 & ~n17508 ;
  assign n17519 = n17516 & n17518 ;
  assign n17520 = ~n17490 & n17519 ;
  assign n17521 = ~n17517 & ~n17520 ;
  assign n17522 = ~\pi0144  & n17521 ;
  assign n17523 = ~n17511 & n17522 ;
  assign n17524 = ~\pi0051  & n17491 ;
  assign n17525 = n17495 & n17524 ;
  assign n17526 = n17480 & n17525 ;
  assign n17527 = n13001 & ~n17507 ;
  assign n17528 = ~n17526 & n17527 ;
  assign n17529 = n17506 & ~n17528 ;
  assign n17530 = ~\pi0144  & ~n17516 ;
  assign n17531 = ~\pi0144  & n17420 ;
  assign n17532 = ~n17514 & n17531 ;
  assign n17533 = ~n17530 & ~n17532 ;
  assign n17534 = ~n17529 & ~n17533 ;
  assign n17535 = \pi0051  & ~\pi0142  ;
  assign n17536 = n6706 & n17535 ;
  assign n17537 = \pi0144  & ~n17536 ;
  assign n17538 = \pi0180  & ~n17537 ;
  assign n17539 = ~\pi0024  & ~\pi0096  ;
  assign n17540 = ~\pi0051  & n17539 ;
  assign n17541 = n1322 & n17540 ;
  assign n17542 = n17502 & n17541 ;
  assign n17543 = n14002 & n17542 ;
  assign n17544 = n1542 & n17543 ;
  assign n17545 = \pi0180  & n15942 ;
  assign n17546 = n17544 & n17545 ;
  assign n17547 = ~n17538 & ~n17546 ;
  assign n17548 = ~n17534 & ~n17547 ;
  assign n17549 = ~n17420 & n17449 ;
  assign n17550 = ~\pi0180  & ~n17537 ;
  assign n17551 = n17549 & n17550 ;
  assign n17552 = ~\pi0179  & ~n17551 ;
  assign n17553 = ~n17548 & n17552 ;
  assign n17554 = \pi0180  & ~n17553 ;
  assign n17555 = ~n17523 & n17554 ;
  assign n17556 = n17465 & n17555 ;
  assign n17557 = n1324 & n17502 ;
  assign n17558 = ~n17453 & n17557 ;
  assign n17559 = n17537 & ~n17558 ;
  assign n17560 = \pi0024  & n17537 ;
  assign n17561 = ~n14006 & n17560 ;
  assign n17562 = ~n17559 & ~n17561 ;
  assign n17563 = ~\pi0180  & n17562 ;
  assign n17564 = \pi0179  & ~n17563 ;
  assign n17565 = n13001 & ~n17489 ;
  assign n17566 = n17479 & n17565 ;
  assign n17567 = ~n17505 & ~n17509 ;
  assign n17568 = ~n17566 & n17567 ;
  assign n17569 = \pi0142  & ~n17568 ;
  assign n17570 = ~\pi0142  & ~n6706 ;
  assign n17571 = ~\pi0051  & ~\pi0142  ;
  assign n17572 = n17419 & n17571 ;
  assign n17573 = ~n17518 & n17572 ;
  assign n17574 = ~n17489 & n17572 ;
  assign n17575 = n17479 & n17574 ;
  assign n17576 = ~n17573 & ~n17575 ;
  assign n17577 = ~n17570 & n17576 ;
  assign n17578 = ~n17569 & n17577 ;
  assign n17579 = ~\pi0144  & \pi0179  ;
  assign n17580 = ~n17578 & n17579 ;
  assign n17581 = ~n17564 & ~n17580 ;
  assign n17582 = ~n17553 & n17581 ;
  assign n17583 = ~\pi0299  & ~n17582 ;
  assign n17584 = ~n17556 & n17583 ;
  assign n17585 = ~\pi0039  & ~\pi0156  ;
  assign n17586 = ~\pi0051  & ~n17462 ;
  assign n17587 = \pi0051  & \pi0146  ;
  assign n17588 = n6706 & ~n17587 ;
  assign n17589 = ~n17586 & n17588 ;
  assign n17590 = \pi0161  & n10696 ;
  assign n17591 = ~n17589 & n17590 ;
  assign n17592 = \pi0146  & ~n17505 ;
  assign n17593 = ~n17509 & n17592 ;
  assign n17594 = ~n17501 & n17593 ;
  assign n17595 = ~\pi0161  & ~n17594 ;
  assign n17596 = ~\pi0146  & n6706 ;
  assign n17597 = ~n17515 & n17596 ;
  assign n17598 = n17518 & n17596 ;
  assign n17599 = ~n17490 & n17598 ;
  assign n17600 = ~n17597 & ~n17599 ;
  assign n17601 = n10696 & n17600 ;
  assign n17602 = n17595 & n17601 ;
  assign n17603 = \pi0146  & ~n17568 ;
  assign n17604 = ~\pi0051  & ~\pi0146  ;
  assign n17605 = n17419 & n17604 ;
  assign n17606 = ~n17518 & n17605 ;
  assign n17607 = ~n17489 & n17605 ;
  assign n17608 = n17479 & n17607 ;
  assign n17609 = ~n17606 & ~n17608 ;
  assign n17610 = ~n11331 & n17609 ;
  assign n17611 = ~n17603 & n17610 ;
  assign n17612 = ~\pi0161  & n10757 ;
  assign n17613 = ~n17611 & n17612 ;
  assign n17614 = \pi0161  & ~n17426 ;
  assign n17615 = ~n17558 & n17614 ;
  assign n17616 = \pi0024  & n17614 ;
  assign n17617 = ~n14006 & n17616 ;
  assign n17618 = ~n17615 & ~n17617 ;
  assign n17619 = n10757 & ~n17618 ;
  assign n17620 = ~\pi0039  & \pi0232  ;
  assign n17621 = ~n17619 & n17620 ;
  assign n17622 = ~n17613 & n17621 ;
  assign n17623 = ~n17602 & n17622 ;
  assign n17624 = ~n17591 & n17623 ;
  assign n17625 = ~n17585 & ~n17624 ;
  assign n17626 = ~n17584 & ~n17625 ;
  assign n17627 = ~\pi0287  & n6706 ;
  assign n17628 = n1281 & n17627 ;
  assign n17629 = n1260 & n17628 ;
  assign n17630 = n17614 & ~n17629 ;
  assign n17631 = n1274 & n1376 ;
  assign n17632 = n10533 & n17631 ;
  assign n17633 = n1273 & n17632 ;
  assign n17634 = ~\pi0077  & n13001 ;
  assign n17635 = n17633 & n17634 ;
  assign n17636 = n17480 & n17635 ;
  assign n17637 = ~\pi0051  & ~\pi0287  ;
  assign n17638 = n17419 & n17637 ;
  assign n17639 = ~n17636 & n17638 ;
  assign n17640 = \pi0051  & ~\pi0287  ;
  assign n17641 = ~n17504 & ~n17627 ;
  assign n17642 = ~n17640 & ~n17641 ;
  assign n17643 = ~n17639 & n17642 ;
  assign n17644 = ~n17630 & n17643 ;
  assign n17645 = \pi0159  & \pi0216  ;
  assign n17646 = n6936 & n17645 ;
  assign n17647 = ~\pi0161  & ~n17426 ;
  assign n17648 = n17646 & n17647 ;
  assign n17649 = n17614 & n17646 ;
  assign n17650 = ~n17629 & n17649 ;
  assign n17651 = ~n17648 & ~n17650 ;
  assign n17652 = ~n17644 & ~n17651 ;
  assign n17653 = \pi0299  & n17646 ;
  assign n17654 = \pi0299  & ~n17429 ;
  assign n17655 = n17421 & n17654 ;
  assign n17656 = ~n17653 & ~n17655 ;
  assign n17657 = n11040 & ~n17656 ;
  assign n17658 = ~n17652 & n17657 ;
  assign n17659 = ~\pi0038  & ~n17658 ;
  assign n17660 = ~\pi0074  & n1287 ;
  assign n17661 = n17421 & ~n17429 ;
  assign n17662 = \pi0299  & ~n17661 ;
  assign n17663 = \pi0232  & ~n17537 ;
  assign n17664 = n17549 & n17663 ;
  assign n17665 = ~n10276 & ~n17664 ;
  assign n17666 = ~n17662 & ~n17665 ;
  assign n17667 = \pi0100  & n17666 ;
  assign n17668 = n17660 & ~n17667 ;
  assign n17669 = n1321 & n17627 ;
  assign n17670 = n1354 & n8592 ;
  assign n17671 = n17669 & n17670 ;
  assign n17672 = n1358 & n17671 ;
  assign n17673 = n6949 & ~n17448 ;
  assign n17674 = \pi0224  & n17673 ;
  assign n17675 = n17672 & n17674 ;
  assign n17676 = \pi0181  & n17537 ;
  assign n17677 = ~n17675 & n17676 ;
  assign n17678 = n6955 & ~n17641 ;
  assign n17679 = ~n17640 & n17678 ;
  assign n17680 = ~n17639 & n17679 ;
  assign n17681 = \pi0181  & ~n17449 ;
  assign n17682 = ~\pi0051  & \pi0181  ;
  assign n17683 = n17419 & n17682 ;
  assign n17684 = ~n17681 & ~n17683 ;
  assign n17685 = n6955 & n17449 ;
  assign n17686 = ~n17420 & n17685 ;
  assign n17687 = ~\pi0144  & ~n17686 ;
  assign n17688 = ~n17684 & n17687 ;
  assign n17689 = ~n17680 & n17688 ;
  assign n17690 = ~n17677 & ~n17689 ;
  assign n17691 = \pi0181  & ~\pi0299  ;
  assign n17692 = ~\pi0299  & ~n17537 ;
  assign n17693 = n17549 & n17692 ;
  assign n17694 = ~n17691 & ~n17693 ;
  assign n17695 = n11040 & ~n17694 ;
  assign n17696 = n17690 & n17695 ;
  assign n17697 = n17668 & ~n17696 ;
  assign n17698 = n17659 & n17697 ;
  assign n17699 = ~n17626 & n17698 ;
  assign n17700 = \pi0232  & ~n10757 ;
  assign n17701 = \pi0232  & ~n17429 ;
  assign n17702 = n17421 & n17701 ;
  assign n17703 = ~n17700 & ~n17702 ;
  assign n17704 = n15942 & n17544 ;
  assign n17705 = n17614 & ~n17704 ;
  assign n17706 = n10696 & n17705 ;
  assign n17707 = ~n17528 & n17592 ;
  assign n17708 = ~n17597 & ~n17707 ;
  assign n17709 = ~\pi0161  & n10696 ;
  assign n17710 = n17708 & n17709 ;
  assign n17711 = ~n17706 & ~n17710 ;
  assign n17712 = ~n17703 & n17711 ;
  assign n17713 = ~\pi0038  & ~\pi0156  ;
  assign n17714 = ~\pi0039  & n17713 ;
  assign n17715 = ~n17712 & n17714 ;
  assign n17716 = \pi0038  & ~n17666 ;
  assign n17717 = ~\pi0100  & ~n17716 ;
  assign n17718 = ~n17715 & n17717 ;
  assign n17719 = n17668 & ~n17718 ;
  assign n17720 = ~\pi0087  & ~n13441 ;
  assign n17721 = ~n17666 & n17720 ;
  assign n17722 = ~\pi0184  & ~\pi0299  ;
  assign n17723 = ~\pi0163  & \pi0299  ;
  assign n17724 = ~n17722 & ~n17723 ;
  assign n17725 = n8640 & n17724 ;
  assign n17726 = \pi0087  & ~n17725 ;
  assign n17727 = n17443 & ~n17726 ;
  assign n17728 = ~n17721 & n17727 ;
  assign n17729 = ~n17719 & n17728 ;
  assign n17730 = ~n17699 & n17729 ;
  assign n17731 = n9948 & ~n17730 ;
  assign n17732 = ~n17420 & n17720 ;
  assign n17733 = ~n17666 & n17732 ;
  assign n17734 = ~n17443 & ~n17726 ;
  assign n17735 = ~n17733 & n17734 ;
  assign n17736 = n17731 & ~n17735 ;
  assign n17737 = \pi0038  & ~n17420 ;
  assign n17738 = ~n17666 & n17737 ;
  assign n17739 = ~\pi0100  & ~n17738 ;
  assign n17740 = \pi0038  & n17739 ;
  assign n17741 = \pi0051  & n6706 ;
  assign n17742 = \pi0072  & ~\pi0095  ;
  assign n17743 = n1634 & n17742 ;
  assign n17744 = n1328 & n17743 ;
  assign n17745 = n1324 & n17744 ;
  assign n17746 = n1319 & n17745 ;
  assign n17747 = ~n17741 & ~n17746 ;
  assign n17748 = n6706 & n17647 ;
  assign n17749 = ~n17747 & n17748 ;
  assign n17750 = ~n17490 & n17518 ;
  assign n17751 = ~\pi0077  & n17480 ;
  assign n17752 = n17633 & n17743 ;
  assign n17753 = n17751 & n17752 ;
  assign n17754 = n17515 & ~n17753 ;
  assign n17755 = ~n17750 & n17754 ;
  assign n17756 = ~\pi0161  & ~n6706 ;
  assign n17757 = ~n17755 & n17756 ;
  assign n17758 = ~n17749 & ~n17757 ;
  assign n17759 = n17419 & n17503 ;
  assign n17760 = ~n17421 & n17515 ;
  assign n17761 = ~n17750 & n17760 ;
  assign n17762 = ~n17759 & ~n17761 ;
  assign n17763 = \pi0146  & ~n17753 ;
  assign n17764 = ~n17762 & n17763 ;
  assign n17765 = ~\pi0146  & n17419 ;
  assign n17766 = ~n17753 & n17765 ;
  assign n17767 = ~\pi0051  & \pi0161  ;
  assign n17768 = n6706 & n17767 ;
  assign n17769 = ~n11320 & ~n17768 ;
  assign n17770 = ~n17766 & ~n17769 ;
  assign n17771 = \pi0161  & ~n6706 ;
  assign n17772 = ~n17755 & n17771 ;
  assign n17773 = ~n17770 & ~n17772 ;
  assign n17774 = ~n17764 & ~n17773 ;
  assign n17775 = n17758 & ~n17774 ;
  assign n17776 = n10696 & ~n17775 ;
  assign n17777 = ~n6706 & n17515 ;
  assign n17778 = ~n17753 & n17777 ;
  assign n17779 = ~n17750 & n17778 ;
  assign n17780 = ~n17753 & n17759 ;
  assign n17781 = \pi0146  & ~n17420 ;
  assign n17782 = ~n17514 & ~n17781 ;
  assign n17783 = n17780 & n17782 ;
  assign n17784 = n17614 & ~n17783 ;
  assign n17785 = ~n17779 & n17784 ;
  assign n17786 = n11331 & n17515 ;
  assign n17787 = ~n17753 & n17786 ;
  assign n17788 = ~n17750 & n17787 ;
  assign n17789 = n14002 & n17541 ;
  assign n17790 = n15942 & n17789 ;
  assign n17791 = n1542 & n17790 ;
  assign n17792 = ~\pi0072  & ~n17791 ;
  assign n17793 = n2575 & ~n17792 ;
  assign n17794 = ~n1629 & n17793 ;
  assign n17795 = n17596 & ~n17794 ;
  assign n17796 = ~\pi0161  & ~n17795 ;
  assign n17797 = ~n17788 & n17796 ;
  assign n17798 = ~n6706 & ~n17755 ;
  assign n17799 = n6706 & ~n17747 ;
  assign n17800 = \pi0146  & ~n17704 ;
  assign n17801 = ~n17799 & n17800 ;
  assign n17802 = ~n17798 & n17801 ;
  assign n17803 = n17797 & ~n17802 ;
  assign n17804 = ~n17785 & ~n17803 ;
  assign n17805 = n10757 & ~n17804 ;
  assign n17806 = ~n17776 & ~n17805 ;
  assign n17807 = \pi0156  & ~n17806 ;
  assign n17808 = ~\pi0051  & ~n17746 ;
  assign n17809 = ~n17462 & n17808 ;
  assign n17810 = n6706 & ~n17809 ;
  assign n17811 = \pi0146  & ~n17798 ;
  assign n17812 = ~n17810 & n17811 ;
  assign n17813 = \pi0146  & n10757 ;
  assign n17814 = n1324 & ~n17458 ;
  assign n17815 = n17457 & n17814 ;
  assign n17816 = ~\pi0072  & n6706 ;
  assign n17817 = ~n17815 & n17816 ;
  assign n17818 = ~n2575 & n6706 ;
  assign n17819 = \pi0072  & n6706 ;
  assign n17820 = ~n1628 & n17819 ;
  assign n17821 = ~n17818 & ~n17820 ;
  assign n17822 = n10757 & ~n17779 ;
  assign n17823 = n17821 & n17822 ;
  assign n17824 = ~n17817 & n17823 ;
  assign n17825 = ~n17813 & ~n17824 ;
  assign n17826 = ~n17812 & ~n17825 ;
  assign n17827 = \pi0024  & ~n14006 ;
  assign n17828 = n17558 & ~n17827 ;
  assign n17829 = \pi0146  & ~n17799 ;
  assign n17830 = ~n17828 & n17829 ;
  assign n17831 = ~n17798 & n17830 ;
  assign n17832 = n10696 & ~n17831 ;
  assign n17833 = ~\pi0161  & ~n17832 ;
  assign n17834 = n1324 & ~n17453 ;
  assign n17835 = ~n17827 & n17834 ;
  assign n17836 = n17816 & ~n17835 ;
  assign n17837 = ~n17779 & n17821 ;
  assign n17838 = ~n17836 & n17837 ;
  assign n17839 = n11365 & ~n17838 ;
  assign n17840 = ~n17833 & ~n17839 ;
  assign n17841 = ~n17826 & ~n17840 ;
  assign n17842 = n17420 & ~n17753 ;
  assign n17843 = n17503 & ~n17842 ;
  assign n17844 = n17503 & n17518 ;
  assign n17845 = ~n17490 & n17844 ;
  assign n17846 = ~n17843 & ~n17845 ;
  assign n17847 = n10696 & ~n17846 ;
  assign n17848 = ~n6706 & n10696 ;
  assign n17849 = ~n17755 & n17848 ;
  assign n17850 = ~n17847 & ~n17849 ;
  assign n17851 = n10696 & ~n17759 ;
  assign n17852 = ~n17761 & n17851 ;
  assign n17853 = ~n17611 & n17852 ;
  assign n17854 = n17850 & ~n17853 ;
  assign n17855 = n10757 & ~n17426 ;
  assign n17856 = ~n17755 & n17855 ;
  assign n17857 = \pi0161  & ~n17856 ;
  assign n17858 = n17854 & n17857 ;
  assign n17859 = ~\pi0156  & ~n17858 ;
  assign n17860 = ~n17841 & n17859 ;
  assign n17861 = ~n17807 & ~n17860 ;
  assign n17862 = n8364 & ~n17861 ;
  assign n17863 = ~\pi0180  & n17537 ;
  assign n17864 = ~n17755 & n17863 ;
  assign n17865 = \pi0142  & ~\pi0144  ;
  assign n17866 = ~\pi0144  & ~n17779 ;
  assign n17867 = n17821 & n17866 ;
  assign n17868 = ~n17817 & n17867 ;
  assign n17869 = ~n17865 & ~n17868 ;
  assign n17870 = \pi0142  & ~n17798 ;
  assign n17871 = ~\pi0180  & ~n17870 ;
  assign n17872 = ~\pi0180  & n6706 ;
  assign n17873 = ~n17809 & n17872 ;
  assign n17874 = ~n17871 & ~n17873 ;
  assign n17875 = ~n17869 & ~n17874 ;
  assign n17876 = ~n17864 & ~n17875 ;
  assign n17877 = \pi0142  & ~n17704 ;
  assign n17878 = ~n17799 & n17877 ;
  assign n17879 = ~n17798 & n17878 ;
  assign n17880 = n17516 & ~n17794 ;
  assign n17881 = n17515 & n17570 ;
  assign n17882 = ~n17753 & n17881 ;
  assign n17883 = ~n17750 & n17882 ;
  assign n17884 = ~\pi0144  & ~n17883 ;
  assign n17885 = ~n17880 & n17884 ;
  assign n17886 = ~n17879 & n17885 ;
  assign n17887 = ~n17514 & ~n17753 ;
  assign n17888 = ~n17762 & n17887 ;
  assign n17889 = n17537 & ~n17888 ;
  assign n17890 = ~\pi0180  & ~n17889 ;
  assign n17891 = ~n17886 & n17890 ;
  assign n17892 = \pi0179  & ~\pi0180  ;
  assign n17893 = \pi0144  & ~n17753 ;
  assign n17894 = ~n17762 & n17893 ;
  assign n17895 = ~n17536 & ~n17894 ;
  assign n17896 = ~\pi0144  & ~n6706 ;
  assign n17897 = ~\pi0144  & ~n17741 ;
  assign n17898 = ~n17746 & n17897 ;
  assign n17899 = ~n17896 & ~n17898 ;
  assign n17900 = \pi0179  & n17899 ;
  assign n17901 = \pi0179  & ~n6706 ;
  assign n17902 = ~n17755 & n17901 ;
  assign n17903 = ~n17900 & ~n17902 ;
  assign n17904 = n17895 & ~n17903 ;
  assign n17905 = ~n17892 & ~n17904 ;
  assign n17906 = ~n17891 & ~n17905 ;
  assign n17907 = ~\pi0142  & n17821 ;
  assign n17908 = ~n17779 & n17907 ;
  assign n17909 = ~n17836 & n17908 ;
  assign n17910 = ~\pi0142  & ~\pi0144  ;
  assign n17911 = ~\pi0144  & ~n17799 ;
  assign n17912 = ~n17828 & n17911 ;
  assign n17913 = ~n17798 & n17912 ;
  assign n17914 = ~n17910 & ~n17913 ;
  assign n17915 = ~n17909 & ~n17914 ;
  assign n17916 = ~n17578 & n17762 ;
  assign n17917 = \pi0144  & n17846 ;
  assign n17918 = ~n17798 & n17917 ;
  assign n17919 = ~n17916 & n17918 ;
  assign n17920 = \pi0180  & ~n17919 ;
  assign n17921 = ~n17915 & n17920 ;
  assign n17922 = ~n17906 & ~n17921 ;
  assign n17923 = n17876 & n17922 ;
  assign n17924 = \pi0179  & ~n17906 ;
  assign n17925 = ~\pi0299  & n8364 ;
  assign n17926 = ~n17924 & n17925 ;
  assign n17927 = ~n17923 & n17926 ;
  assign n17928 = ~n17862 & ~n17927 ;
  assign n17929 = ~\pi0299  & n6949 ;
  assign n17930 = ~n7412 & ~n17929 ;
  assign n17931 = n13001 & ~n17930 ;
  assign n17932 = n17633 & n17931 ;
  assign n17933 = n17751 & n17932 ;
  assign n17934 = ~\pi0051  & ~\pi0232  ;
  assign n17935 = n17419 & n17934 ;
  assign n17936 = ~n17933 & n17935 ;
  assign n17937 = \pi0039  & ~n17936 ;
  assign n17938 = ~\pi0039  & ~\pi0232  ;
  assign n17939 = ~n17755 & n17938 ;
  assign n17940 = ~n17937 & ~n17939 ;
  assign n17941 = n1264 & n1321 ;
  assign n17942 = n1263 & n17941 ;
  assign n17943 = n1354 & n17942 ;
  assign n17944 = n1358 & n17943 ;
  assign n17945 = ~\pi0051  & ~n17944 ;
  assign n17946 = n6706 & ~n17945 ;
  assign n17947 = \pi0142  & n6706 ;
  assign n17948 = \pi0142  & n17420 ;
  assign n17949 = ~n17636 & n17948 ;
  assign n17950 = ~n17947 & ~n17949 ;
  assign n17951 = ~n17946 & ~n17950 ;
  assign n17952 = \pi0181  & \pi0224  ;
  assign n17953 = n17420 & ~n17636 ;
  assign n17954 = ~n6706 & ~n17953 ;
  assign n17955 = n1281 & n6706 ;
  assign n17956 = n1260 & n17955 ;
  assign n17957 = ~\pi0142  & ~n17956 ;
  assign n17958 = ~n17954 & n17957 ;
  assign n17959 = ~n17952 & ~n17958 ;
  assign n17960 = ~n17951 & n17959 ;
  assign n17961 = n6706 & ~n17637 ;
  assign n17962 = ~n17945 & n17961 ;
  assign n17963 = ~n17954 & ~n17962 ;
  assign n17964 = ~n17536 & n17952 ;
  assign n17965 = ~n17963 & n17964 ;
  assign n17966 = ~n17960 & ~n17965 ;
  assign n17967 = n6949 & n17966 ;
  assign n17968 = ~n6949 & n17504 ;
  assign n17969 = ~n6949 & n17536 ;
  assign n17970 = ~\pi0051  & ~n6949 ;
  assign n17971 = n17419 & n17970 ;
  assign n17972 = ~n17969 & ~n17971 ;
  assign n17973 = n11250 & n17972 ;
  assign n17974 = ~n17968 & n17973 ;
  assign n17975 = ~n17967 & n17974 ;
  assign n17976 = ~n17680 & ~n17686 ;
  assign n17977 = \pi0181  & n17419 ;
  assign n17978 = ~n17976 & n17977 ;
  assign n17979 = ~n17741 & ~n17953 ;
  assign n17980 = n17673 & ~n17979 ;
  assign n17981 = \pi0144  & n17972 ;
  assign n17982 = ~\pi0299  & n17981 ;
  assign n17983 = ~n17980 & n17982 ;
  assign n17984 = ~n17978 & n17983 ;
  assign n17985 = n6706 & ~n6936 ;
  assign n17986 = ~n17429 & n17985 ;
  assign n17987 = ~\pi0051  & ~n6936 ;
  assign n17988 = n17419 & n17987 ;
  assign n17989 = n11302 & ~n17988 ;
  assign n17990 = ~n17986 & n17989 ;
  assign n17991 = \pi0161  & n17426 ;
  assign n17992 = \pi0161  & n17420 ;
  assign n17993 = ~n17636 & n17992 ;
  assign n17994 = ~n17991 & ~n17993 ;
  assign n17995 = n17990 & n17994 ;
  assign n17996 = ~n6936 & n11302 ;
  assign n17997 = ~n17420 & n17996 ;
  assign n17998 = ~n17986 & n17997 ;
  assign n17999 = \pi0232  & ~n17998 ;
  assign n18000 = ~n17995 & n17999 ;
  assign n18001 = \pi0146  & n17954 ;
  assign n18002 = n11376 & ~n17945 ;
  assign n18003 = ~n18001 & ~n18002 ;
  assign n18004 = n11331 & ~n17953 ;
  assign n18005 = ~\pi0146  & n1259 ;
  assign n18006 = n1249 & n18005 ;
  assign n18007 = n17955 & n18006 ;
  assign n18008 = ~\pi0161  & ~n18007 ;
  assign n18009 = ~n18004 & n18008 ;
  assign n18010 = n17999 & n18009 ;
  assign n18011 = n18003 & n18010 ;
  assign n18012 = ~n18000 & ~n18011 ;
  assign n18013 = ~n17984 & ~n18012 ;
  assign n18014 = ~n17975 & n18013 ;
  assign n18015 = ~\pi0216  & n17994 ;
  assign n18016 = n6936 & ~n18015 ;
  assign n18017 = n6936 & n18009 ;
  assign n18018 = n18003 & n18017 ;
  assign n18019 = ~n18016 & ~n18018 ;
  assign n18020 = \pi0216  & ~n17420 ;
  assign n18021 = \pi0216  & ~n17627 ;
  assign n18022 = n17636 & n18021 ;
  assign n18023 = ~n18020 & ~n18022 ;
  assign n18024 = n17614 & ~n18023 ;
  assign n18025 = ~\pi0161  & \pi0216  ;
  assign n18026 = ~n17426 & n18025 ;
  assign n18027 = ~n17963 & n18026 ;
  assign n18028 = ~n18024 & ~n18027 ;
  assign n18029 = ~n18019 & n18028 ;
  assign n18030 = ~n17986 & ~n17988 ;
  assign n18031 = n11327 & n18030 ;
  assign n18032 = ~n18029 & n18031 ;
  assign n18033 = ~n17939 & ~n18032 ;
  assign n18034 = n18014 & n18033 ;
  assign n18035 = ~n17940 & ~n18034 ;
  assign n18036 = n17739 & ~n18035 ;
  assign n18037 = n17928 & n18036 ;
  assign n18038 = ~n17740 & ~n18037 ;
  assign n18039 = ~\pi0051  & \pi0100  ;
  assign n18040 = n17419 & n18039 ;
  assign n18041 = n17660 & ~n18040 ;
  assign n18042 = ~n17667 & n18041 ;
  assign n18043 = n17731 & n18042 ;
  assign n18044 = n18038 & n18043 ;
  assign n18045 = ~n17736 & ~n18044 ;
  assign n18046 = ~n17447 & n18045 ;
  assign n18047 = n8696 & n9998 ;
  assign n18048 = n9250 & ~n17400 ;
  assign n18049 = ~n17397 & n18048 ;
  assign n18050 = ~n17404 & ~n18049 ;
  assign n18051 = ~n18047 & ~n18050 ;
  assign n18052 = ~\pi0075  & ~n17383 ;
  assign n18053 = n12003 & ~n17346 ;
  assign n18054 = ~n18052 & n18053 ;
  assign n18055 = n9948 & ~n17333 ;
  assign n18056 = ~n18047 & ~n18055 ;
  assign n18057 = ~n18054 & n18056 ;
  assign n18058 = ~n18051 & ~n18057 ;
  assign n18059 = ~\pi0072  & n2575 ;
  assign n18060 = n2575 & n12101 ;
  assign n18061 = n1319 & n18060 ;
  assign n18062 = ~n18059 & ~n18061 ;
  assign n18063 = ~\pi0110  & n18062 ;
  assign n18064 = ~\pi0072  & ~\pi0110  ;
  assign n18065 = ~n18063 & ~n18064 ;
  assign n18066 = ~\pi0090  & ~n13666 ;
  assign n18067 = \pi0081  & ~\pi0090  ;
  assign n18068 = ~n1528 & n18067 ;
  assign n18069 = ~n18066 & ~n18068 ;
  assign n18070 = \pi0071  & n6989 ;
  assign n18071 = n1236 & n18070 ;
  assign n18072 = n1248 & n18071 ;
  assign n18073 = ~\pi0081  & ~\pi0090  ;
  assign n18074 = ~n18072 & n18073 ;
  assign n18075 = n18069 & ~n18074 ;
  assign n18076 = ~\pi0111  & ~n7015 ;
  assign n18077 = ~n1413 & n10308 ;
  assign n18078 = ~n18076 & n18077 ;
  assign n18079 = ~\pi0083  & ~n18078 ;
  assign n18080 = ~\pi0111  & n1233 ;
  assign n18081 = ~\pi0083  & n18080 ;
  assign n18082 = ~n7013 & n18081 ;
  assign n18083 = ~n18079 & ~n18082 ;
  assign n18084 = ~\pi0067  & ~\pi0069  ;
  assign n18085 = ~n18083 & n18084 ;
  assign n18086 = \pi0067  & ~n1472 ;
  assign n18087 = ~n1479 & ~n18086 ;
  assign n18088 = ~\pi0083  & ~n18087 ;
  assign n18089 = n1483 & ~n6993 ;
  assign n18090 = ~n18088 & n18089 ;
  assign n18091 = n18069 & n18090 ;
  assign n18092 = ~n18085 & n18091 ;
  assign n18093 = ~n18075 & ~n18092 ;
  assign n18094 = ~\pi0090  & n1651 ;
  assign n18095 = n1651 & n12100 ;
  assign n18096 = n1319 & n18095 ;
  assign n18097 = ~n18094 & ~n18096 ;
  assign n18098 = ~\pi0093  & ~n18097 ;
  assign n18099 = ~n18063 & n18098 ;
  assign n18100 = ~n18093 & n18099 ;
  assign n18101 = ~n18065 & ~n18100 ;
  assign n18102 = ~\pi0110  & n6922 ;
  assign n18103 = ~n6931 & n18102 ;
  assign n18104 = n6722 & n18103 ;
  assign n18105 = ~n6744 & n18104 ;
  assign n18106 = n7412 & n18105 ;
  assign n18107 = n6706 & n17929 ;
  assign n18108 = ~n6761 & n18107 ;
  assign n18109 = ~n6706 & n17929 ;
  assign n18110 = ~n6713 & n18109 ;
  assign n18111 = ~n18108 & ~n18110 ;
  assign n18112 = n18104 & ~n18111 ;
  assign n18113 = \pi0039  & ~n18112 ;
  assign n18114 = ~n18106 & n18113 ;
  assign n18115 = \pi0110  & \pi0824  ;
  assign n18116 = n6809 & n18115 ;
  assign n18117 = ~n6704 & n18116 ;
  assign n18118 = ~n6808 & n18117 ;
  assign n18119 = ~n8641 & n18118 ;
  assign n18120 = ~\pi0039  & ~n15410 ;
  assign n18121 = ~n18119 & n18120 ;
  assign n18122 = ~n18114 & ~n18121 ;
  assign n18123 = n15956 & n18122 ;
  assign n18124 = ~n18101 & n18123 ;
  assign n18125 = n2575 & ~n15956 ;
  assign n18126 = n1291 & ~n18125 ;
  assign n18127 = \pi0072  & n1291 ;
  assign n18128 = ~n1628 & n18127 ;
  assign n18129 = ~n18126 & ~n18128 ;
  assign n18130 = ~\pi0072  & n1291 ;
  assign n18131 = n18129 & ~n18130 ;
  assign n18132 = ~n1609 & n1651 ;
  assign n18133 = n18129 & n18132 ;
  assign n18134 = ~n18093 & n18133 ;
  assign n18135 = ~n18131 & ~n18134 ;
  assign n18136 = n18122 & ~n18135 ;
  assign n18137 = n9948 & ~n18136 ;
  assign n18138 = ~n18124 & n18137 ;
  assign n18139 = \pi0039  & n6936 ;
  assign n18140 = n18105 & n18139 ;
  assign n18141 = n1801 & n8640 ;
  assign n18142 = ~\pi0039  & \pi0110  ;
  assign n18143 = ~n18141 & n18142 ;
  assign n18144 = n15860 & n18143 ;
  assign n18145 = ~n6808 & n18144 ;
  assign n18146 = ~n9948 & ~n18145 ;
  assign n18147 = ~n18140 & n18146 ;
  assign n18148 = ~n18138 & ~n18147 ;
  assign n18149 = ~\pi0125  & n17438 ;
  assign n18150 = \pi0125  & \pi0133  ;
  assign n18151 = ~n17439 & ~n18150 ;
  assign n18152 = ~n18149 & ~n18151 ;
  assign n18153 = n17444 & ~n18152 ;
  assign n18154 = \pi0051  & \pi0172  ;
  assign n18155 = n6706 & n18154 ;
  assign n18156 = ~\pi0051  & ~\pi0152  ;
  assign n18157 = n6706 & n18156 ;
  assign n18158 = ~n17419 & n18157 ;
  assign n18159 = ~n18155 & ~n18158 ;
  assign n18160 = n17422 & ~n18159 ;
  assign n18161 = \pi0087  & n11181 ;
  assign n18162 = ~n9948 & ~n18161 ;
  assign n18163 = ~n18160 & n18162 ;
  assign n18164 = ~n18153 & n18163 ;
  assign n18165 = ~\pi0051  & ~\pi0174  ;
  assign n18166 = n6706 & n18165 ;
  assign n18167 = ~n17419 & n18166 ;
  assign n18168 = \pi0051  & \pi0193  ;
  assign n18169 = n6706 & n18168 ;
  assign n18170 = ~\pi0299  & ~n18169 ;
  assign n18171 = ~n18167 & n18170 ;
  assign n18172 = \pi0232  & ~n18171 ;
  assign n18173 = \pi0299  & ~n18155 ;
  assign n18174 = ~n18158 & n18173 ;
  assign n18175 = \pi0100  & ~n18174 ;
  assign n18176 = n18172 & n18175 ;
  assign n18177 = n18041 & ~n18176 ;
  assign n18178 = \pi0216  & n6936 ;
  assign n18179 = n13001 & n18178 ;
  assign n18180 = n17633 & n18179 ;
  assign n18181 = n17751 & n18180 ;
  assign n18182 = ~\pi0051  & \pi0299  ;
  assign n18183 = n17419 & n18182 ;
  assign n18184 = ~n18181 & n18183 ;
  assign n18185 = \pi0224  & n6949 ;
  assign n18186 = n13001 & n18185 ;
  assign n18187 = n17633 & n18186 ;
  assign n18188 = n17751 & n18187 ;
  assign n18189 = ~\pi0051  & ~\pi0299  ;
  assign n18190 = n17419 & n18189 ;
  assign n18191 = ~n18188 & n18190 ;
  assign n18192 = ~n18184 & ~n18191 ;
  assign n18193 = ~\pi0232  & n18192 ;
  assign n18194 = \pi0039  & ~n18193 ;
  assign n18195 = ~\pi0039  & n17515 ;
  assign n18196 = ~n17750 & n18195 ;
  assign n18197 = ~n18194 & ~n18196 ;
  assign n18198 = ~\pi0152  & \pi0216  ;
  assign n18199 = n6936 & n18198 ;
  assign n18200 = ~n17954 & n18199 ;
  assign n18201 = ~n17962 & n18200 ;
  assign n18202 = n10696 & ~n18201 ;
  assign n18203 = ~n17420 & n18159 ;
  assign n18204 = ~n7597 & ~n18203 ;
  assign n18205 = ~n17627 & n17636 ;
  assign n18206 = ~\pi0051  & \pi0152  ;
  assign n18207 = n17419 & n18206 ;
  assign n18208 = ~n18205 & n18207 ;
  assign n18209 = ~n18155 & ~n18208 ;
  assign n18210 = n7597 & ~n18209 ;
  assign n18211 = ~n18204 & ~n18210 ;
  assign n18212 = n18202 & n18211 ;
  assign n18213 = \pi0152  & ~n17979 ;
  assign n18214 = ~\pi0152  & ~n17956 ;
  assign n18215 = ~n17954 & n18214 ;
  assign n18216 = \pi0172  & ~n18215 ;
  assign n18217 = ~n18213 & n18216 ;
  assign n18218 = ~n10260 & ~n17953 ;
  assign n18219 = ~\pi0172  & n18218 ;
  assign n18220 = ~\pi0172  & n10260 ;
  assign n18221 = ~n17945 & n18220 ;
  assign n18222 = ~n18219 & ~n18221 ;
  assign n18223 = n7597 & n18222 ;
  assign n18224 = ~n18217 & n18223 ;
  assign n18225 = n7597 & n10757 ;
  assign n18226 = n10757 & ~n17420 ;
  assign n18227 = n18159 & n18226 ;
  assign n18228 = ~n18225 & ~n18227 ;
  assign n18229 = ~n18224 & ~n18228 ;
  assign n18230 = ~n18212 & ~n18229 ;
  assign n18231 = ~\pi0174  & n6955 ;
  assign n18232 = ~\pi0174  & ~n6706 ;
  assign n18233 = ~n17420 & n18232 ;
  assign n18234 = ~n18231 & ~n18233 ;
  assign n18235 = \pi0287  & n6706 ;
  assign n18236 = n1281 & n18235 ;
  assign n18237 = n1260 & n18236 ;
  assign n18238 = n6955 & n17420 ;
  assign n18239 = ~n17636 & n18238 ;
  assign n18240 = ~n10241 & ~n18239 ;
  assign n18241 = ~n18237 & ~n18240 ;
  assign n18242 = ~n18234 & ~n18241 ;
  assign n18243 = \pi0174  & ~n17420 ;
  assign n18244 = \pi0174  & n18187 ;
  assign n18245 = n17751 & n18244 ;
  assign n18246 = ~n18243 & ~n18245 ;
  assign n18247 = ~n17741 & ~n17759 ;
  assign n18248 = ~n17627 & ~n17741 ;
  assign n18249 = n17636 & n18248 ;
  assign n18250 = ~n18247 & ~n18249 ;
  assign n18251 = ~n18246 & ~n18250 ;
  assign n18252 = \pi0180  & ~n18251 ;
  assign n18253 = ~n18242 & n18252 ;
  assign n18254 = n6955 & ~n17956 ;
  assign n18255 = ~n17954 & n18254 ;
  assign n18256 = ~n18234 & ~n18255 ;
  assign n18257 = \pi0174  & ~n17741 ;
  assign n18258 = ~n17420 & n18257 ;
  assign n18259 = n18187 & n18257 ;
  assign n18260 = n17751 & n18259 ;
  assign n18261 = ~n18258 & ~n18260 ;
  assign n18262 = ~\pi0180  & n18261 ;
  assign n18263 = ~n18256 & n18262 ;
  assign n18264 = ~n18253 & ~n18263 ;
  assign n18265 = \pi0193  & ~n18264 ;
  assign n18266 = n6955 & ~n17954 ;
  assign n18267 = ~n17946 & n18266 ;
  assign n18268 = n6706 & n17637 ;
  assign n18269 = \pi0180  & n18268 ;
  assign n18270 = ~\pi0174  & ~n18269 ;
  assign n18271 = ~n6706 & ~n17419 ;
  assign n18272 = ~\pi0051  & ~n6955 ;
  assign n18273 = ~n18271 & n18272 ;
  assign n18274 = n18270 & ~n18273 ;
  assign n18275 = ~n18267 & n18274 ;
  assign n18276 = ~\pi0051  & \pi0180  ;
  assign n18277 = n17419 & n18276 ;
  assign n18278 = ~n18205 & n18277 ;
  assign n18279 = ~n18246 & ~n18278 ;
  assign n18280 = ~\pi0193  & ~n18279 ;
  assign n18281 = ~n18275 & n18280 ;
  assign n18282 = ~\pi0299  & ~n18281 ;
  assign n18283 = ~n18265 & n18282 ;
  assign n18284 = n18230 & ~n18283 ;
  assign n18285 = \pi0232  & ~n18196 ;
  assign n18286 = ~n18284 & n18285 ;
  assign n18287 = ~n18197 & ~n18286 ;
  assign n18288 = ~\pi0038  & ~n8364 ;
  assign n18289 = ~n18287 & n18288 ;
  assign n18290 = ~\pi0100  & ~n18174 ;
  assign n18291 = n18172 & n18290 ;
  assign n18292 = ~\pi0051  & ~\pi0100  ;
  assign n18293 = n17419 & n18292 ;
  assign n18294 = ~n2327 & ~n18293 ;
  assign n18295 = ~n18291 & n18294 ;
  assign n18296 = ~n18289 & ~n18295 ;
  assign n18297 = n18177 & ~n18296 ;
  assign n18298 = \pi0174  & n6706 ;
  assign n18299 = n17420 & n18298 ;
  assign n18300 = ~n17514 & n18299 ;
  assign n18301 = \pi0174  & n17515 ;
  assign n18302 = ~n17750 & n18301 ;
  assign n18303 = ~n18300 & ~n18302 ;
  assign n18304 = ~\pi0193  & ~n18303 ;
  assign n18305 = n17515 & ~n17741 ;
  assign n18306 = ~n17750 & n18305 ;
  assign n18307 = ~n17503 & ~n18306 ;
  assign n18308 = ~\pi0145  & n15942 ;
  assign n18309 = n17544 & n18308 ;
  assign n18310 = ~\pi0174  & ~\pi0193  ;
  assign n18311 = \pi0145  & ~\pi0193  ;
  assign n18312 = n17419 & n18311 ;
  assign n18313 = ~n18310 & ~n18312 ;
  assign n18314 = ~n18309 & ~n18313 ;
  assign n18315 = ~n18307 & n18314 ;
  assign n18316 = ~n18304 & ~n18315 ;
  assign n18317 = ~\pi0174  & ~n18309 ;
  assign n18318 = \pi0145  & ~n17504 ;
  assign n18319 = ~\pi0145  & \pi0174  ;
  assign n18320 = ~n18318 & ~n18319 ;
  assign n18321 = ~n17505 & ~n18318 ;
  assign n18322 = ~n17528 & n18321 ;
  assign n18323 = ~n18320 & ~n18322 ;
  assign n18324 = ~n18317 & ~n18323 ;
  assign n18325 = ~n6706 & ~n17515 ;
  assign n18326 = ~n6706 & n17518 ;
  assign n18327 = ~n17490 & n18326 ;
  assign n18328 = ~n18325 & ~n18327 ;
  assign n18329 = \pi0193  & n18328 ;
  assign n18330 = ~n18324 & n18329 ;
  assign n18331 = n11478 & ~n18330 ;
  assign n18332 = n18316 & n18331 ;
  assign n18333 = ~\pi0038  & n18332 ;
  assign n18334 = ~n17501 & n17567 ;
  assign n18335 = n18328 & ~n18334 ;
  assign n18336 = ~n17515 & ~n17759 ;
  assign n18337 = ~\pi0145  & ~n17515 ;
  assign n18338 = ~n18336 & ~n18337 ;
  assign n18339 = ~n17750 & n18338 ;
  assign n18340 = n13001 & n18339 ;
  assign n18341 = \pi0174  & ~n18340 ;
  assign n18342 = ~n18335 & n18341 ;
  assign n18343 = \pi0193  & ~n18342 ;
  assign n18344 = ~n17828 & n18328 ;
  assign n18345 = \pi0145  & n18344 ;
  assign n18346 = ~\pi0174  & ~n18345 ;
  assign n18347 = ~n17458 & n17557 ;
  assign n18348 = n17457 & n18347 ;
  assign n18349 = ~\pi0145  & n18328 ;
  assign n18350 = ~n18348 & n18349 ;
  assign n18351 = n18346 & ~n18350 ;
  assign n18352 = n18343 & ~n18351 ;
  assign n18353 = n11446 & ~n18352 ;
  assign n18354 = ~\pi0145  & ~n6706 ;
  assign n18355 = n17515 & n18354 ;
  assign n18356 = ~n17750 & n18355 ;
  assign n18357 = ~\pi0051  & ~\pi0145  ;
  assign n18358 = n18328 & n18357 ;
  assign n18359 = ~n17462 & n18358 ;
  assign n18360 = ~n18356 & ~n18359 ;
  assign n18361 = ~\pi0051  & \pi0145  ;
  assign n18362 = n18344 & n18361 ;
  assign n18363 = ~\pi0174  & ~n18362 ;
  assign n18364 = n18360 & n18363 ;
  assign n18365 = \pi0174  & ~n18339 ;
  assign n18366 = ~\pi0193  & ~n18365 ;
  assign n18367 = ~n18364 & n18366 ;
  assign n18368 = ~\pi0038  & ~n18367 ;
  assign n18369 = n18353 & n18368 ;
  assign n18370 = ~n18333 & ~n18369 ;
  assign n18371 = n18328 & ~n18348 ;
  assign n18372 = ~\pi0152  & ~n18371 ;
  assign n18373 = \pi0152  & ~n18335 ;
  assign n18374 = \pi0172  & ~n18373 ;
  assign n18375 = ~n18372 & n18374 ;
  assign n18376 = n10260 & ~n17586 ;
  assign n18377 = ~n10260 & ~n17515 ;
  assign n18378 = ~n10260 & n17518 ;
  assign n18379 = ~n17490 & n18378 ;
  assign n18380 = ~n18377 & ~n18379 ;
  assign n18381 = ~\pi0172  & n18380 ;
  assign n18382 = ~n18376 & n18381 ;
  assign n18383 = ~n18375 & ~n18382 ;
  assign n18384 = ~\pi0197  & ~n18383 ;
  assign n18385 = ~n17750 & ~n18336 ;
  assign n18386 = ~\pi0172  & n18385 ;
  assign n18387 = \pi0172  & ~n17568 ;
  assign n18388 = n18328 & n18387 ;
  assign n18389 = ~n18386 & ~n18388 ;
  assign n18390 = \pi0152  & n18389 ;
  assign n18391 = ~\pi0152  & ~n18344 ;
  assign n18392 = \pi0051  & ~\pi0172  ;
  assign n18393 = n6706 & n18392 ;
  assign n18394 = \pi0197  & ~n18393 ;
  assign n18395 = ~n18391 & n18394 ;
  assign n18396 = ~n18390 & n18395 ;
  assign n18397 = n11588 & ~n18396 ;
  assign n18398 = ~n18384 & n18397 ;
  assign n18399 = ~\pi0152  & ~n18393 ;
  assign n18400 = ~n17704 & n18399 ;
  assign n18401 = n18328 & n18400 ;
  assign n18402 = ~\pi0197  & n18401 ;
  assign n18403 = ~n17505 & ~n17528 ;
  assign n18404 = n18328 & ~n18403 ;
  assign n18405 = \pi0172  & ~n18404 ;
  assign n18406 = ~\pi0172  & ~n6706 ;
  assign n18407 = n17518 & n18406 ;
  assign n18408 = ~n17490 & n18407 ;
  assign n18409 = ~\pi0172  & ~n17515 ;
  assign n18410 = \pi0152  & ~n18409 ;
  assign n18411 = ~n18408 & n18410 ;
  assign n18412 = ~\pi0197  & n18411 ;
  assign n18413 = ~n18405 & n18412 ;
  assign n18414 = ~n18402 & ~n18413 ;
  assign n18415 = n6706 & n18206 ;
  assign n18416 = ~n17419 & n18415 ;
  assign n18417 = n17515 & ~n18416 ;
  assign n18418 = ~n17750 & n18417 ;
  assign n18419 = n6706 & ~n18416 ;
  assign n18420 = \pi0172  & ~n18419 ;
  assign n18421 = ~n18418 & n18420 ;
  assign n18422 = ~\pi0172  & ~n18158 ;
  assign n18423 = ~n17759 & n18422 ;
  assign n18424 = ~n17761 & n18423 ;
  assign n18425 = \pi0197  & ~n18424 ;
  assign n18426 = ~n18421 & n18425 ;
  assign n18427 = n11598 & ~n18426 ;
  assign n18428 = n18414 & n18427 ;
  assign n18429 = ~n18398 & ~n18428 ;
  assign n18430 = n18370 & n18429 ;
  assign n18431 = n8364 & n18177 ;
  assign n18432 = ~n18430 & n18431 ;
  assign n18433 = ~n18297 & ~n18432 ;
  assign n18434 = \pi0140  & ~\pi0299  ;
  assign n18435 = \pi0162  & \pi0299  ;
  assign n18436 = ~n18434 & ~n18435 ;
  assign n18437 = n8640 & ~n18436 ;
  assign n18438 = \pi0087  & ~n18437 ;
  assign n18439 = n18172 & ~n18174 ;
  assign n18440 = n17732 & ~n18439 ;
  assign n18441 = ~n18152 & ~n18440 ;
  assign n18442 = ~n18438 & n18441 ;
  assign n18443 = n18433 & n18442 ;
  assign n18444 = ~n17720 & ~n18438 ;
  assign n18445 = ~n18174 & ~n18438 ;
  assign n18446 = n18172 & n18445 ;
  assign n18447 = ~n18444 & ~n18446 ;
  assign n18448 = n18152 & ~n18447 ;
  assign n18449 = n9948 & ~n18448 ;
  assign n18450 = \pi0232  & n9627 ;
  assign n18451 = ~n2327 & ~n18291 ;
  assign n18452 = n11452 & ~n17746 ;
  assign n18453 = ~n9627 & ~n18452 ;
  assign n18454 = n6936 & n13621 ;
  assign n18455 = n3058 & n6148 ;
  assign n18456 = ~n18454 & ~n18455 ;
  assign n18457 = n1281 & ~n18456 ;
  assign n18458 = n1260 & n18457 ;
  assign n18459 = ~\pi0232  & ~n18458 ;
  assign n18460 = \pi0039  & ~n18459 ;
  assign n18461 = ~n18453 & ~n18460 ;
  assign n18462 = ~n18451 & ~n18461 ;
  assign n18463 = ~n18450 & n18462 ;
  assign n18464 = ~\pi0224  & n6949 ;
  assign n18465 = n6949 & ~n17641 ;
  assign n18466 = ~n17640 & n18465 ;
  assign n18467 = ~n17639 & n18466 ;
  assign n18468 = ~n18464 & ~n18467 ;
  assign n18469 = n17503 & ~n17953 ;
  assign n18470 = n1281 & ~n6706 ;
  assign n18471 = n1260 & n18470 ;
  assign n18472 = ~\pi0224  & ~n18471 ;
  assign n18473 = ~n18469 & n18472 ;
  assign n18474 = ~\pi0193  & ~n18473 ;
  assign n18475 = ~n18468 & n18474 ;
  assign n18476 = n6706 & ~n17953 ;
  assign n18477 = n8701 & ~n18471 ;
  assign n18478 = ~n18476 & n18477 ;
  assign n18479 = ~n6706 & ~n6949 ;
  assign n18480 = ~n17971 & ~n18479 ;
  assign n18481 = \pi0224  & ~n6706 ;
  assign n18482 = ~\pi0051  & \pi0224  ;
  assign n18483 = n17419 & n18482 ;
  assign n18484 = ~n18481 & ~n18483 ;
  assign n18485 = n18480 & n18484 ;
  assign n18486 = n17627 & n18480 ;
  assign n18487 = n17636 & n18486 ;
  assign n18488 = ~n18485 & ~n18487 ;
  assign n18489 = \pi0193  & ~n18488 ;
  assign n18490 = ~n18478 & n18489 ;
  assign n18491 = ~\pi0193  & ~n6949 ;
  assign n18492 = n17504 & n18491 ;
  assign n18493 = ~\pi0174  & ~n18492 ;
  assign n18494 = ~n18490 & n18493 ;
  assign n18495 = ~n18475 & n18494 ;
  assign n18496 = \pi0224  & ~n17741 ;
  assign n18497 = ~n17672 & n18496 ;
  assign n18498 = n6949 & ~n18497 ;
  assign n18499 = \pi0051  & ~n6706 ;
  assign n18500 = n8701 & n18499 ;
  assign n18501 = ~\pi0051  & n8701 ;
  assign n18502 = ~n17944 & n18501 ;
  assign n18503 = ~n18500 & ~n18502 ;
  assign n18504 = n18498 & n18503 ;
  assign n18505 = n6955 & n17627 ;
  assign n18506 = ~n8701 & ~n18505 ;
  assign n18507 = ~\pi0193  & ~n18506 ;
  assign n18508 = n1281 & n18507 ;
  assign n18509 = n1260 & n18508 ;
  assign n18510 = n18257 & ~n18509 ;
  assign n18511 = ~n18504 & n18510 ;
  assign n18512 = \pi0174  & ~\pi0193  ;
  assign n18513 = ~n18509 & n18512 ;
  assign n18514 = \pi0180  & ~n18513 ;
  assign n18515 = ~n18511 & n18514 ;
  assign n18516 = ~n18495 & n18515 ;
  assign n18517 = ~\pi0174  & n8701 ;
  assign n18518 = n11029 & ~n17420 ;
  assign n18519 = ~n18517 & ~n18518 ;
  assign n18520 = n18471 & ~n18519 ;
  assign n18521 = n17503 & ~n18519 ;
  assign n18522 = ~n17953 & n18521 ;
  assign n18523 = ~n18520 & ~n18522 ;
  assign n18524 = n1321 & n8701 ;
  assign n18525 = n17670 & n18524 ;
  assign n18526 = n1358 & n18525 ;
  assign n18527 = ~\pi0051  & \pi0174  ;
  assign n18528 = n18526 & n18527 ;
  assign n18529 = ~n18169 & ~n18528 ;
  assign n18530 = n18523 & n18529 ;
  assign n18531 = ~\pi0180  & ~n18530 ;
  assign n18532 = ~\pi0299  & ~n18531 ;
  assign n18533 = ~n18516 & n18532 ;
  assign n18534 = ~n8684 & ~n18155 ;
  assign n18535 = ~n18158 & n18534 ;
  assign n18536 = ~n8684 & ~n18535 ;
  assign n18537 = ~\pi0152  & ~n18471 ;
  assign n18538 = ~n18476 & n18537 ;
  assign n18539 = ~n18392 & ~n18538 ;
  assign n18540 = \pi0152  & n18499 ;
  assign n18541 = ~n17944 & n18206 ;
  assign n18542 = ~n18540 & ~n18541 ;
  assign n18543 = ~n18535 & n18542 ;
  assign n18544 = n18539 & n18543 ;
  assign n18545 = ~n18536 & ~n18544 ;
  assign n18546 = n10757 & n18545 ;
  assign n18547 = ~n18533 & ~n18546 ;
  assign n18548 = ~\pi0152  & ~n17641 ;
  assign n18549 = ~n17640 & n18548 ;
  assign n18550 = ~n17639 & n18549 ;
  assign n18551 = \pi0152  & ~\pi0287  ;
  assign n18552 = n6706 & n18551 ;
  assign n18553 = n1281 & n18552 ;
  assign n18554 = n1260 & n18553 ;
  assign n18555 = ~\pi0172  & ~n18554 ;
  assign n18556 = ~n18550 & n18555 ;
  assign n18557 = \pi0216  & n18556 ;
  assign n18558 = ~n17672 & ~n17741 ;
  assign n18559 = \pi0152  & ~n18558 ;
  assign n18560 = \pi0172  & ~n6706 ;
  assign n18561 = ~\pi0051  & \pi0172  ;
  assign n18562 = n17419 & n18561 ;
  assign n18563 = ~n18560 & ~n18562 ;
  assign n18564 = ~n10716 & n18563 ;
  assign n18565 = ~n10716 & n17627 ;
  assign n18566 = n17636 & n18565 ;
  assign n18567 = ~n18564 & ~n18566 ;
  assign n18568 = \pi0216  & n18567 ;
  assign n18569 = ~n18559 & n18568 ;
  assign n18570 = ~n18557 & ~n18569 ;
  assign n18571 = n6936 & n18542 ;
  assign n18572 = n18539 & n18571 ;
  assign n18573 = ~n18178 & ~n18572 ;
  assign n18574 = n18570 & ~n18573 ;
  assign n18575 = n6936 & n10696 ;
  assign n18576 = n10696 & ~n18155 ;
  assign n18577 = ~n18158 & n18576 ;
  assign n18578 = ~n18575 & ~n18577 ;
  assign n18579 = ~n18574 & ~n18578 ;
  assign n18580 = n18462 & ~n18579 ;
  assign n18581 = n18547 & n18580 ;
  assign n18582 = ~n18463 & ~n18581 ;
  assign n18583 = ~n8364 & ~n18582 ;
  assign n18584 = ~n6706 & ~n17746 ;
  assign n18585 = \pi0152  & ~n18584 ;
  assign n18586 = ~n17809 & n18585 ;
  assign n18587 = ~n17753 & ~n18154 ;
  assign n18588 = n17515 & n18587 ;
  assign n18589 = ~n17750 & n18588 ;
  assign n18590 = n6706 & n18589 ;
  assign n18591 = \pi0072  & ~n6706 ;
  assign n18592 = n2575 & n18591 ;
  assign n18593 = n1627 & n18592 ;
  assign n18594 = n1319 & n18593 ;
  assign n18595 = ~n17503 & ~n18155 ;
  assign n18596 = ~n18594 & n18595 ;
  assign n18597 = ~\pi0152  & ~n18596 ;
  assign n18598 = ~n18590 & n18597 ;
  assign n18599 = ~n10697 & ~n18598 ;
  assign n18600 = ~n18586 & n18599 ;
  assign n18601 = n17821 & ~n18584 ;
  assign n18602 = ~n17817 & n18601 ;
  assign n18603 = ~\pi0172  & ~n18597 ;
  assign n18604 = ~\pi0172  & n6706 ;
  assign n18605 = n18589 & n18604 ;
  assign n18606 = ~n18603 & ~n18605 ;
  assign n18607 = ~n18602 & ~n18606 ;
  assign n18608 = ~n18600 & ~n18607 ;
  assign n18609 = n17752 & n18157 ;
  assign n18610 = n17751 & n18609 ;
  assign n18611 = ~n18158 & ~n18610 ;
  assign n18612 = ~n10260 & n17743 ;
  assign n18613 = n1627 & n18612 ;
  assign n18614 = n1319 & n18613 ;
  assign n18615 = ~\pi0197  & ~n18155 ;
  assign n18616 = ~n18614 & n18615 ;
  assign n18617 = n18611 & n18616 ;
  assign n18618 = n11409 & n18617 ;
  assign n18619 = ~n17503 & ~n18594 ;
  assign n18620 = ~n17514 & n17759 ;
  assign n18621 = ~n17753 & n18620 ;
  assign n18622 = ~n18619 & ~n18621 ;
  assign n18623 = ~\pi0152  & \pi0197  ;
  assign n18624 = ~n18155 & n18623 ;
  assign n18625 = n11409 & n18624 ;
  assign n18626 = ~n18622 & n18625 ;
  assign n18627 = ~n18618 & ~n18626 ;
  assign n18628 = n6706 & ~n17794 ;
  assign n18629 = ~\pi0172  & ~n18584 ;
  assign n18630 = ~n18628 & n18629 ;
  assign n18631 = \pi0152  & \pi0197  ;
  assign n18632 = ~\pi0172  & n18631 ;
  assign n18633 = ~n17704 & n18631 ;
  assign n18634 = n17747 & n18633 ;
  assign n18635 = ~n18632 & ~n18634 ;
  assign n18636 = n11409 & ~n18635 ;
  assign n18637 = ~n18630 & n18636 ;
  assign n18638 = n18627 & ~n18637 ;
  assign n18639 = \pi0197  & n18638 ;
  assign n18640 = n18608 & n18639 ;
  assign n18641 = ~\pi0172  & ~\pi0197  ;
  assign n18642 = n17420 & n17780 ;
  assign n18643 = ~n17750 & n18642 ;
  assign n18644 = ~\pi0152  & ~n18584 ;
  assign n18645 = ~\pi0197  & n18644 ;
  assign n18646 = ~n18643 & n18645 ;
  assign n18647 = ~n18641 & ~n18646 ;
  assign n18648 = \pi0152  & ~\pi0197  ;
  assign n18649 = ~n17747 & n18648 ;
  assign n18650 = n17558 & n18648 ;
  assign n18651 = ~n17827 & n18650 ;
  assign n18652 = ~n18649 & ~n18651 ;
  assign n18653 = n11417 & n18652 ;
  assign n18654 = n18647 & n18653 ;
  assign n18655 = n17821 & n18585 ;
  assign n18656 = ~n17836 & n18655 ;
  assign n18657 = ~n17842 & n18157 ;
  assign n18658 = n17518 & n18157 ;
  assign n18659 = ~n17490 & n18658 ;
  assign n18660 = ~n18657 & ~n18659 ;
  assign n18661 = ~\pi0152  & n18594 ;
  assign n18662 = ~\pi0172  & n11417 ;
  assign n18663 = ~n18661 & n18662 ;
  assign n18664 = n18660 & n18663 ;
  assign n18665 = ~n18656 & n18664 ;
  assign n18666 = ~n18654 & ~n18665 ;
  assign n18667 = n18638 & n18666 ;
  assign n18668 = \pi0299  & ~n18667 ;
  assign n18669 = ~n18640 & n18668 ;
  assign n18670 = \pi0145  & n18622 ;
  assign n18671 = ~\pi0145  & n18594 ;
  assign n18672 = ~\pi0174  & ~n18671 ;
  assign n18673 = n6706 & n18357 ;
  assign n18674 = ~n17419 & n18673 ;
  assign n18675 = n17752 & n18673 ;
  assign n18676 = n17751 & n18675 ;
  assign n18677 = ~n18674 & ~n18676 ;
  assign n18678 = ~\pi0193  & n18677 ;
  assign n18679 = n18672 & n18678 ;
  assign n18680 = ~n18670 & n18679 ;
  assign n18681 = \pi0145  & ~n18584 ;
  assign n18682 = \pi0072  & ~\pi0145  ;
  assign n18683 = n2575 & n18682 ;
  assign n18684 = n1627 & n18683 ;
  assign n18685 = n1319 & n18684 ;
  assign n18686 = n18512 & ~n18685 ;
  assign n18687 = ~n18681 & n18686 ;
  assign n18688 = n6706 & n18686 ;
  assign n18689 = ~n17794 & n18688 ;
  assign n18690 = ~n18687 & ~n18689 ;
  assign n18691 = ~n18680 & n18690 ;
  assign n18692 = ~n17704 & n17747 ;
  assign n18693 = ~n17746 & n18309 ;
  assign n18694 = \pi0174  & ~n18693 ;
  assign n18695 = ~n18692 & n18694 ;
  assign n18696 = \pi0193  & n18584 ;
  assign n18697 = ~\pi0174  & ~n17780 ;
  assign n18698 = ~n17514 & ~n17741 ;
  assign n18699 = \pi0145  & ~\pi0174  ;
  assign n18700 = ~n18698 & n18699 ;
  assign n18701 = \pi0193  & ~n18700 ;
  assign n18702 = ~n18697 & n18701 ;
  assign n18703 = ~n18696 & ~n18702 ;
  assign n18704 = ~n18695 & ~n18703 ;
  assign n18705 = n18691 & ~n18704 ;
  assign n18706 = ~\pi0038  & n11446 ;
  assign n18707 = ~n18705 & n18706 ;
  assign n18708 = ~n18669 & ~n18707 ;
  assign n18709 = ~\pi0145  & ~n17741 ;
  assign n18710 = ~n17746 & n18709 ;
  assign n18711 = \pi0193  & ~n18710 ;
  assign n18712 = \pi0193  & n17558 ;
  assign n18713 = ~n17827 & n18712 ;
  assign n18714 = ~n18711 & ~n18713 ;
  assign n18715 = \pi0174  & ~n18584 ;
  assign n18716 = ~n17809 & n18715 ;
  assign n18717 = ~n18319 & ~n18716 ;
  assign n18718 = ~n18714 & ~n18717 ;
  assign n18719 = \pi0145  & ~n18602 ;
  assign n18720 = ~\pi0193  & ~n18584 ;
  assign n18721 = n17821 & n18720 ;
  assign n18722 = ~n17836 & n18721 ;
  assign n18723 = ~n18311 & ~n18722 ;
  assign n18724 = \pi0174  & ~n18723 ;
  assign n18725 = ~n18719 & n18724 ;
  assign n18726 = ~n18718 & ~n18725 ;
  assign n18727 = n17846 & ~n18594 ;
  assign n18728 = ~\pi0193  & ~n18727 ;
  assign n18729 = \pi0193  & ~n18584 ;
  assign n18730 = ~n18643 & n18729 ;
  assign n18731 = ~\pi0145  & ~n18730 ;
  assign n18732 = ~n18728 & n18731 ;
  assign n18733 = \pi0145  & ~n18169 ;
  assign n18734 = ~n17753 & n18733 ;
  assign n18735 = n17515 & n18734 ;
  assign n18736 = ~n17750 & n18735 ;
  assign n18737 = n6706 & n18736 ;
  assign n18738 = ~n17503 & n18733 ;
  assign n18739 = ~n18594 & n18738 ;
  assign n18740 = ~\pi0174  & ~n18739 ;
  assign n18741 = ~n18737 & n18740 ;
  assign n18742 = ~n18732 & n18741 ;
  assign n18743 = ~\pi0038  & n11478 ;
  assign n18744 = ~n18742 & n18743 ;
  assign n18745 = n18726 & n18744 ;
  assign n18746 = ~n18582 & ~n18745 ;
  assign n18747 = n18708 & n18746 ;
  assign n18748 = ~n18583 & ~n18747 ;
  assign n18749 = n17660 & ~n18176 ;
  assign n18750 = n9948 & n18749 ;
  assign n18751 = n18748 & n18750 ;
  assign n18752 = ~n18449 & ~n18751 ;
  assign n18753 = ~n18443 & ~n18752 ;
  assign n18754 = ~n18164 & ~n18753 ;
  assign n18755 = ~\pi0232  & ~n17746 ;
  assign n18756 = ~\pi0039  & ~n18755 ;
  assign n18757 = ~\pi0232  & n18756 ;
  assign n18758 = ~\pi0153  & ~n18584 ;
  assign n18759 = n17821 & n18758 ;
  assign n18760 = ~n17817 & n18759 ;
  assign n18761 = \pi0153  & ~n18584 ;
  assign n18762 = ~n17809 & n18761 ;
  assign n18763 = \pi0157  & ~n18762 ;
  assign n18764 = ~n18760 & n18763 ;
  assign n18765 = n6706 & n17515 ;
  assign n18766 = ~n17753 & n18765 ;
  assign n18767 = ~n17750 & n18766 ;
  assign n18768 = \pi0157  & ~n18619 ;
  assign n18769 = ~n18767 & n18768 ;
  assign n18770 = ~\pi0157  & n18622 ;
  assign n18771 = \pi0051  & \pi0153  ;
  assign n18772 = n6706 & n18771 ;
  assign n18773 = ~\pi0166  & ~n18772 ;
  assign n18774 = ~n18770 & n18773 ;
  assign n18775 = ~n18769 & n18774 ;
  assign n18776 = ~n18628 & n18758 ;
  assign n18777 = ~\pi0153  & ~\pi0157  ;
  assign n18778 = ~\pi0157  & ~n17704 ;
  assign n18779 = n17747 & n18778 ;
  assign n18780 = ~n18777 & ~n18779 ;
  assign n18781 = ~n18776 & ~n18780 ;
  assign n18782 = ~n18775 & ~n18781 ;
  assign n18783 = ~n18764 & n18782 ;
  assign n18784 = ~\pi0166  & ~n18775 ;
  assign n18785 = n11327 & ~n18784 ;
  assign n18786 = ~n18783 & n18785 ;
  assign n18787 = ~\pi0189  & ~n18619 ;
  assign n18788 = ~n18767 & n18787 ;
  assign n18789 = \pi0178  & ~n18788 ;
  assign n18790 = \pi0178  & \pi0181  ;
  assign n18791 = ~\pi0189  & ~n17741 ;
  assign n18792 = ~n18622 & n18791 ;
  assign n18793 = \pi0189  & ~n17704 ;
  assign n18794 = n17747 & n18793 ;
  assign n18795 = \pi0181  & ~n18794 ;
  assign n18796 = ~n18792 & n18795 ;
  assign n18797 = ~n18790 & ~n18796 ;
  assign n18798 = ~n18789 & ~n18797 ;
  assign n18799 = ~n17809 & ~n18584 ;
  assign n18800 = ~\pi0189  & ~n18307 ;
  assign n18801 = ~n18797 & ~n18800 ;
  assign n18802 = n18799 & n18801 ;
  assign n18803 = ~n18798 & ~n18802 ;
  assign n18804 = n17747 & ~n17828 ;
  assign n18805 = ~\pi0189  & n18594 ;
  assign n18806 = ~\pi0051  & ~\pi0189  ;
  assign n18807 = n6706 & n18806 ;
  assign n18808 = ~n17419 & n18807 ;
  assign n18809 = n17752 & n18807 ;
  assign n18810 = n17751 & n18809 ;
  assign n18811 = ~n18808 & ~n18810 ;
  assign n18812 = ~n18805 & n18811 ;
  assign n18813 = ~\pi0178  & ~n17741 ;
  assign n18814 = \pi0189  & n17746 ;
  assign n18815 = n18813 & ~n18814 ;
  assign n18816 = n18812 & n18815 ;
  assign n18817 = ~\pi0181  & \pi0189  ;
  assign n18818 = ~n18816 & n18817 ;
  assign n18819 = ~n18804 & n18818 ;
  assign n18820 = ~\pi0181  & ~n18816 ;
  assign n18821 = n14285 & ~n18820 ;
  assign n18822 = ~\pi0189  & ~n18584 ;
  assign n18823 = ~n18643 & n18822 ;
  assign n18824 = \pi0178  & n14285 ;
  assign n18825 = ~n18823 & n18824 ;
  assign n18826 = ~n18821 & ~n18825 ;
  assign n18827 = ~n18819 & ~n18826 ;
  assign n18828 = n18803 & n18827 ;
  assign n18829 = \pi0166  & ~n18584 ;
  assign n18830 = n17821 & n18829 ;
  assign n18831 = ~n17836 & n18830 ;
  assign n18832 = ~\pi0153  & \pi0166  ;
  assign n18833 = ~\pi0153  & ~n18594 ;
  assign n18834 = n17846 & n18833 ;
  assign n18835 = ~n18832 & ~n18834 ;
  assign n18836 = ~n18831 & ~n18835 ;
  assign n18837 = \pi0157  & n18836 ;
  assign n18838 = ~\pi0166  & ~n18584 ;
  assign n18839 = ~n18643 & n18838 ;
  assign n18840 = \pi0153  & ~n18839 ;
  assign n18841 = \pi0166  & ~n17747 ;
  assign n18842 = \pi0166  & n17558 ;
  assign n18843 = ~n17827 & n18842 ;
  assign n18844 = ~n18841 & ~n18843 ;
  assign n18845 = \pi0157  & n18844 ;
  assign n18846 = n18840 & n18845 ;
  assign n18847 = ~\pi0166  & n18594 ;
  assign n18848 = ~\pi0051  & ~\pi0166  ;
  assign n18849 = n6706 & n18848 ;
  assign n18850 = ~n17419 & n18849 ;
  assign n18851 = n17752 & n18849 ;
  assign n18852 = n17751 & n18851 ;
  assign n18853 = ~n18850 & ~n18852 ;
  assign n18854 = ~n18847 & n18853 ;
  assign n18855 = ~\pi0157  & ~n18772 ;
  assign n18856 = \pi0166  & n17746 ;
  assign n18857 = n18855 & ~n18856 ;
  assign n18858 = n18854 & n18857 ;
  assign n18859 = ~n18846 & ~n18858 ;
  assign n18860 = ~n18837 & n18859 ;
  assign n18861 = n11302 & ~n18860 ;
  assign n18862 = ~n18828 & ~n18861 ;
  assign n18863 = ~n18786 & n18862 ;
  assign n18864 = \pi0189  & ~n18584 ;
  assign n18865 = n17821 & n18864 ;
  assign n18866 = ~n17817 & n18865 ;
  assign n18867 = \pi0189  & n18584 ;
  assign n18868 = n14297 & ~n17794 ;
  assign n18869 = ~n18867 & ~n18868 ;
  assign n18870 = ~\pi0189  & ~n18622 ;
  assign n18871 = ~\pi0178  & ~n18870 ;
  assign n18872 = n18869 & n18871 ;
  assign n18873 = ~n18788 & ~n18872 ;
  assign n18874 = ~n18866 & n18873 ;
  assign n18875 = \pi0181  & ~n18870 ;
  assign n18876 = n18869 & n18875 ;
  assign n18877 = ~n18790 & ~n18876 ;
  assign n18878 = ~n18874 & ~n18877 ;
  assign n18879 = n17503 & n17752 ;
  assign n18880 = n17751 & n18879 ;
  assign n18881 = ~n17504 & ~n18880 ;
  assign n18882 = ~\pi0178  & ~n18594 ;
  assign n18883 = ~n18814 & n18882 ;
  assign n18884 = n18881 & n18883 ;
  assign n18885 = n18820 & ~n18884 ;
  assign n18886 = n14266 & ~n18885 ;
  assign n18887 = ~n17836 & n18865 ;
  assign n18888 = ~n17842 & n18807 ;
  assign n18889 = n17518 & n18807 ;
  assign n18890 = ~n17490 & n18889 ;
  assign n18891 = ~n18888 & ~n18890 ;
  assign n18892 = \pi0178  & n14266 ;
  assign n18893 = ~n18805 & n18892 ;
  assign n18894 = n18891 & n18893 ;
  assign n18895 = ~n18887 & n18894 ;
  assign n18896 = ~n18886 & ~n18895 ;
  assign n18897 = ~n18878 & ~n18896 ;
  assign n18898 = n18756 & ~n18897 ;
  assign n18899 = n18863 & n18898 ;
  assign n18900 = ~n18757 & ~n18899 ;
  assign n18901 = ~\pi0126  & ~\pi0132  ;
  assign n18902 = n17437 & n18901 ;
  assign n18903 = ~\pi0121  & ~\pi0126  ;
  assign n18904 = n17439 & n18903 ;
  assign n18905 = \pi0126  & ~n17441 ;
  assign n18906 = ~n18904 & ~n18905 ;
  assign n18907 = ~n18902 & ~n18906 ;
  assign n18908 = \pi0189  & ~n18506 ;
  assign n18909 = n1281 & n18908 ;
  assign n18910 = n1260 & n18909 ;
  assign n18911 = \pi0182  & ~n18910 ;
  assign n18912 = \pi0189  & n18911 ;
  assign n18913 = ~n18468 & ~n18473 ;
  assign n18914 = ~n17968 & n18911 ;
  assign n18915 = ~n18913 & n18914 ;
  assign n18916 = ~n18912 & ~n18915 ;
  assign n18917 = n14266 & ~n18916 ;
  assign n18918 = \pi0166  & ~n17741 ;
  assign n18919 = ~n17672 & n18918 ;
  assign n18920 = ~\pi0166  & ~n6706 ;
  assign n18921 = n17419 & n18848 ;
  assign n18922 = ~n18920 & ~n18921 ;
  assign n18923 = \pi0153  & n18922 ;
  assign n18924 = \pi0153  & n17627 ;
  assign n18925 = n17636 & n18924 ;
  assign n18926 = ~n18923 & ~n18925 ;
  assign n18927 = ~n18919 & ~n18926 ;
  assign n18928 = \pi0160  & n18927 ;
  assign n18929 = ~\pi0166  & ~n17641 ;
  assign n18930 = ~n17640 & n18929 ;
  assign n18931 = ~n17639 & n18930 ;
  assign n18932 = ~\pi0287  & n14139 ;
  assign n18933 = n1281 & n18932 ;
  assign n18934 = n1260 & n18933 ;
  assign n18935 = ~n18931 & ~n18934 ;
  assign n18936 = n14197 & ~n18935 ;
  assign n18937 = ~n18928 & ~n18936 ;
  assign n18938 = ~n11984 & ~n17419 ;
  assign n18939 = ~\pi0051  & ~n18938 ;
  assign n18940 = ~n18772 & ~n18939 ;
  assign n18941 = ~\pi0051  & ~n17504 ;
  assign n18942 = ~\pi0160  & \pi0216  ;
  assign n18943 = n6936 & ~n18942 ;
  assign n18944 = ~n18941 & ~n18943 ;
  assign n18945 = ~n18940 & n18944 ;
  assign n18946 = \pi0299  & ~n18945 ;
  assign n18947 = \pi0216  & n18946 ;
  assign n18948 = n18937 & n18947 ;
  assign n18949 = ~\pi0189  & n8701 ;
  assign n18950 = n12330 & ~n17420 ;
  assign n18951 = ~n18949 & ~n18950 ;
  assign n18952 = n18471 & ~n18951 ;
  assign n18953 = n17503 & ~n18951 ;
  assign n18954 = ~n17953 & n18953 ;
  assign n18955 = ~n18952 & ~n18954 ;
  assign n18956 = ~\pi0051  & \pi0189  ;
  assign n18957 = n18526 & n18956 ;
  assign n18958 = ~\pi0182  & n14266 ;
  assign n18959 = ~n18957 & n18958 ;
  assign n18960 = n18955 & n18959 ;
  assign n18961 = ~\pi0166  & ~n18471 ;
  assign n18962 = ~n18476 & n18961 ;
  assign n18963 = ~\pi0051  & \pi0166  ;
  assign n18964 = ~n17944 & n18963 ;
  assign n18965 = \pi0051  & ~\pi0153  ;
  assign n18966 = \pi0051  & \pi0166  ;
  assign n18967 = ~n6706 & n18966 ;
  assign n18968 = n6936 & ~n18967 ;
  assign n18969 = ~n18965 & n18968 ;
  assign n18970 = ~n18964 & n18969 ;
  assign n18971 = ~n18962 & n18970 ;
  assign n18972 = ~n7597 & n18946 ;
  assign n18973 = ~n18971 & n18972 ;
  assign n18974 = ~n18960 & ~n18973 ;
  assign n18975 = ~n18948 & n18974 ;
  assign n18976 = ~n18917 & n18975 ;
  assign n18977 = ~\pi0182  & ~n17741 ;
  assign n18978 = ~n18957 & n18977 ;
  assign n18979 = n14285 & n18955 ;
  assign n18980 = n18978 & n18979 ;
  assign n18981 = ~n17741 & ~n18504 ;
  assign n18982 = \pi0189  & ~n18981 ;
  assign n18983 = ~\pi0189  & ~n18488 ;
  assign n18984 = ~n18478 & n18983 ;
  assign n18985 = \pi0182  & n14285 ;
  assign n18986 = ~n18984 & n18985 ;
  assign n18987 = ~n18982 & n18986 ;
  assign n18988 = ~n18980 & ~n18987 ;
  assign n18989 = n18976 & n18988 ;
  assign n18990 = \pi0232  & ~n18989 ;
  assign n18991 = n18460 & ~n18990 ;
  assign n18992 = n18907 & ~n18991 ;
  assign n18993 = n18900 & n18992 ;
  assign n18994 = ~n17568 & n18328 ;
  assign n18995 = \pi0153  & \pi0166  ;
  assign n18996 = ~n18994 & n18995 ;
  assign n18997 = \pi0051  & ~\pi0166  ;
  assign n18998 = n6706 & n18997 ;
  assign n18999 = \pi0166  & n18336 ;
  assign n19000 = \pi0166  & n17518 ;
  assign n19001 = ~n17490 & n19000 ;
  assign n19002 = ~n18999 & ~n19001 ;
  assign n19003 = ~n18998 & n19002 ;
  assign n19004 = ~\pi0153  & ~n19003 ;
  assign n19005 = ~n18996 & ~n19004 ;
  assign n19006 = ~\pi0166  & ~n18344 ;
  assign n19007 = ~\pi0157  & ~n19006 ;
  assign n19008 = n19005 & n19007 ;
  assign n19009 = n6706 & n18963 ;
  assign n19010 = ~n17419 & n19009 ;
  assign n19011 = n17515 & ~n19010 ;
  assign n19012 = ~n17750 & n19011 ;
  assign n19013 = n6706 & ~n19010 ;
  assign n19014 = \pi0153  & ~n19013 ;
  assign n19015 = ~n19012 & n19014 ;
  assign n19016 = \pi0157  & ~n19015 ;
  assign n19017 = ~\pi0153  & ~n18850 ;
  assign n19018 = ~n17759 & n19017 ;
  assign n19019 = ~n17761 & n19018 ;
  assign n19020 = n19016 & ~n19019 ;
  assign n19021 = n11327 & ~n19020 ;
  assign n19022 = ~n19008 & n19021 ;
  assign n19023 = ~n12330 & ~n17515 ;
  assign n19024 = ~n12330 & n17518 ;
  assign n19025 = ~n17490 & n19024 ;
  assign n19026 = ~n19023 & ~n19025 ;
  assign n19027 = ~n12330 & n19026 ;
  assign n19028 = ~\pi0051  & n19026 ;
  assign n19029 = ~n17462 & n19028 ;
  assign n19030 = ~n19027 & ~n19029 ;
  assign n19031 = ~\pi0178  & n19030 ;
  assign n19032 = \pi0189  & n17515 ;
  assign n19033 = ~n17750 & n19032 ;
  assign n19034 = n14297 & n17420 ;
  assign n19035 = ~n17514 & n19034 ;
  assign n19036 = \pi0178  & ~n19035 ;
  assign n19037 = ~n19033 & n19036 ;
  assign n19038 = ~\pi0189  & ~n17704 ;
  assign n19039 = n18328 & n19038 ;
  assign n19040 = ~n18307 & n19039 ;
  assign n19041 = n19037 & ~n19040 ;
  assign n19042 = ~\pi0181  & ~n19041 ;
  assign n19043 = ~n19031 & n19042 ;
  assign n19044 = ~\pi0189  & ~n17828 ;
  assign n19045 = ~n18307 & n19044 ;
  assign n19046 = \pi0189  & ~n18336 ;
  assign n19047 = ~n17750 & n19046 ;
  assign n19048 = ~\pi0178  & ~n19047 ;
  assign n19049 = ~n19045 & n19048 ;
  assign n19050 = \pi0178  & \pi0189  ;
  assign n19051 = ~n17759 & n19050 ;
  assign n19052 = ~n17761 & n19051 ;
  assign n19053 = \pi0178  & ~\pi0189  ;
  assign n19054 = ~n17503 & n19053 ;
  assign n19055 = ~n18306 & n19054 ;
  assign n19056 = \pi0181  & ~n19055 ;
  assign n19057 = ~n19052 & n19056 ;
  assign n19058 = ~n19049 & n19057 ;
  assign n19059 = n14266 & ~n19058 ;
  assign n19060 = ~n19043 & n19059 ;
  assign n19061 = ~\pi0189  & n18328 ;
  assign n19062 = ~n18348 & n19061 ;
  assign n19063 = \pi0189  & n18335 ;
  assign n19064 = ~\pi0178  & ~n19063 ;
  assign n19065 = ~n19062 & n19064 ;
  assign n19066 = \pi0178  & ~n19039 ;
  assign n19067 = \pi0189  & ~n18403 ;
  assign n19068 = n18328 & n19067 ;
  assign n19069 = n19066 & ~n19068 ;
  assign n19070 = ~\pi0181  & ~n19069 ;
  assign n19071 = ~n19065 & n19070 ;
  assign n19072 = n6706 & n19050 ;
  assign n19073 = n17507 & n19072 ;
  assign n19074 = \pi0181  & ~n19073 ;
  assign n19075 = n17515 & n19074 ;
  assign n19076 = ~n17750 & n19075 ;
  assign n19077 = \pi0181  & n6706 ;
  assign n19078 = ~n19073 & n19077 ;
  assign n19079 = n14285 & ~n19078 ;
  assign n19080 = ~n19076 & n19079 ;
  assign n19081 = ~\pi0189  & ~n17558 ;
  assign n19082 = \pi0024  & ~\pi0189  ;
  assign n19083 = ~n14006 & n19082 ;
  assign n19084 = ~n19081 & ~n19083 ;
  assign n19085 = ~\pi0178  & ~\pi0189  ;
  assign n19086 = ~\pi0178  & ~n17505 ;
  assign n19087 = ~n17509 & n19086 ;
  assign n19088 = ~n17566 & n19087 ;
  assign n19089 = ~n19085 & ~n19088 ;
  assign n19090 = n19084 & ~n19089 ;
  assign n19091 = n14285 & n19090 ;
  assign n19092 = ~n19080 & ~n19091 ;
  assign n19093 = ~n19071 & ~n19092 ;
  assign n19094 = ~n19060 & ~n19093 ;
  assign n19095 = ~n19022 & n19094 ;
  assign n19096 = ~\pi0232  & ~n17515 ;
  assign n19097 = ~\pi0232  & n17518 ;
  assign n19098 = ~n17490 & n19097 ;
  assign n19099 = ~n19096 & ~n19098 ;
  assign n19100 = ~\pi0039  & n19099 ;
  assign n19101 = ~n11984 & ~n17515 ;
  assign n19102 = ~n11984 & n17518 ;
  assign n19103 = ~n17490 & n19102 ;
  assign n19104 = ~n19101 & ~n19103 ;
  assign n19105 = ~n11984 & n19104 ;
  assign n19106 = ~\pi0051  & n19104 ;
  assign n19107 = ~n17462 & n19106 ;
  assign n19108 = ~n19105 & ~n19107 ;
  assign n19109 = ~\pi0153  & n19108 ;
  assign n19110 = ~\pi0166  & n18328 ;
  assign n19111 = ~n18348 & n19110 ;
  assign n19112 = \pi0166  & n18335 ;
  assign n19113 = \pi0153  & ~n19112 ;
  assign n19114 = ~n19111 & n19113 ;
  assign n19115 = ~n19109 & ~n19114 ;
  assign n19116 = ~\pi0157  & n19115 ;
  assign n19117 = \pi0166  & ~n6706 ;
  assign n19118 = n17518 & n19117 ;
  assign n19119 = ~n17490 & n19118 ;
  assign n19120 = \pi0166  & ~n17515 ;
  assign n19121 = ~n18998 & ~n19120 ;
  assign n19122 = ~n19119 & n19121 ;
  assign n19123 = ~\pi0153  & ~n19122 ;
  assign n19124 = ~n18404 & n18995 ;
  assign n19125 = \pi0157  & \pi0166  ;
  assign n19126 = \pi0157  & ~n17704 ;
  assign n19127 = n18328 & n19126 ;
  assign n19128 = ~n19125 & ~n19127 ;
  assign n19129 = ~n19124 & ~n19128 ;
  assign n19130 = ~n19123 & n19129 ;
  assign n19131 = n11302 & ~n19130 ;
  assign n19132 = ~n19116 & n19131 ;
  assign n19133 = n19100 & ~n19132 ;
  assign n19134 = n19095 & n19133 ;
  assign n19135 = ~n6706 & ~n17420 ;
  assign n19136 = ~n6955 & ~n19135 ;
  assign n19137 = ~\pi0189  & n19136 ;
  assign n19138 = ~\pi0189  & ~n18237 ;
  assign n19139 = ~n18240 & n19138 ;
  assign n19140 = ~n19137 & ~n19139 ;
  assign n19141 = \pi0182  & ~\pi0189  ;
  assign n19142 = \pi0182  & ~n17420 ;
  assign n19143 = \pi0182  & n18187 ;
  assign n19144 = n17751 & n19143 ;
  assign n19145 = ~n19142 & ~n19144 ;
  assign n19146 = ~n18250 & ~n19145 ;
  assign n19147 = ~n19141 & ~n19146 ;
  assign n19148 = n19140 & ~n19147 ;
  assign n19149 = n14285 & n19148 ;
  assign n19150 = ~n18255 & ~n19136 ;
  assign n19151 = ~\pi0189  & ~n19150 ;
  assign n19152 = \pi0189  & n17420 ;
  assign n19153 = ~n18188 & n19152 ;
  assign n19154 = \pi0051  & \pi0189  ;
  assign n19155 = n6706 & n19154 ;
  assign n19156 = ~\pi0182  & n14285 ;
  assign n19157 = ~n19155 & n19156 ;
  assign n19158 = ~n19153 & n19157 ;
  assign n19159 = ~n19151 & n19158 ;
  assign n19160 = ~n19149 & ~n19159 ;
  assign n19161 = ~\pi0051  & \pi0182  ;
  assign n19162 = n17419 & n19161 ;
  assign n19163 = ~n18205 & n19162 ;
  assign n19164 = \pi0189  & ~n17420 ;
  assign n19165 = \pi0189  & n18187 ;
  assign n19166 = n17751 & n19165 ;
  assign n19167 = ~n19164 & ~n19166 ;
  assign n19168 = ~n19163 & ~n19167 ;
  assign n19169 = \pi0182  & n18268 ;
  assign n19170 = ~\pi0189  & ~n19169 ;
  assign n19171 = ~n18273 & n19170 ;
  assign n19172 = ~n18267 & n19171 ;
  assign n19173 = ~n19168 & ~n19172 ;
  assign n19174 = n14266 & ~n19173 ;
  assign n19175 = n19160 & ~n19174 ;
  assign n19176 = \pi0232  & ~n19175 ;
  assign n19177 = ~\pi0166  & ~n17954 ;
  assign n19178 = ~n17962 & n19177 ;
  assign n19179 = \pi0160  & ~n18772 ;
  assign n19180 = n17419 & n18963 ;
  assign n19181 = ~n18205 & n19180 ;
  assign n19182 = n19179 & ~n19181 ;
  assign n19183 = ~n19178 & n19182 ;
  assign n19184 = ~n17953 & n18918 ;
  assign n19185 = ~n17953 & n18920 ;
  assign n19186 = ~\pi0166  & n1259 ;
  assign n19187 = n1249 & n19186 ;
  assign n19188 = n17955 & n19187 ;
  assign n19189 = \pi0153  & ~n19188 ;
  assign n19190 = ~n19185 & n19189 ;
  assign n19191 = ~n19184 & n19190 ;
  assign n19192 = ~\pi0153  & n11984 ;
  assign n19193 = ~\pi0153  & n17420 ;
  assign n19194 = ~n17636 & n19193 ;
  assign n19195 = ~n19192 & ~n19194 ;
  assign n19196 = ~\pi0160  & n19195 ;
  assign n19197 = ~\pi0160  & n11984 ;
  assign n19198 = ~n17945 & n19197 ;
  assign n19199 = ~n19196 & ~n19198 ;
  assign n19200 = ~n19191 & ~n19199 ;
  assign n19201 = ~n19183 & ~n19200 ;
  assign n19202 = n7597 & n19201 ;
  assign n19203 = ~n7597 & n18772 ;
  assign n19204 = ~\pi0051  & ~n7597 ;
  assign n19205 = ~n18938 & n19204 ;
  assign n19206 = ~n19203 & ~n19205 ;
  assign n19207 = n10276 & n19206 ;
  assign n19208 = ~n19202 & n19207 ;
  assign n19209 = n18194 & ~n19208 ;
  assign n19210 = ~n19176 & n19209 ;
  assign n19211 = n17515 & n17938 ;
  assign n19212 = ~n17750 & n19211 ;
  assign n19213 = ~n18907 & ~n19212 ;
  assign n19214 = ~n19210 & n19213 ;
  assign n19215 = ~n19134 & n19214 ;
  assign n19216 = n2327 & ~n19215 ;
  assign n19217 = ~n18993 & n19216 ;
  assign n19218 = ~n17504 & n18182 ;
  assign n19219 = \pi0299  & ~n18772 ;
  assign n19220 = ~n18939 & n19219 ;
  assign n19221 = ~n19218 & ~n19220 ;
  assign n19222 = \pi0051  & \pi0175  ;
  assign n19223 = n6706 & n19222 ;
  assign n19224 = ~\pi0299  & ~n19223 ;
  assign n19225 = ~n18808 & n19224 ;
  assign n19226 = \pi0232  & ~n19225 ;
  assign n19227 = ~n2327 & n19226 ;
  assign n19228 = n19221 & n19227 ;
  assign n19229 = ~n2327 & n17420 ;
  assign n19230 = ~n18907 & n19229 ;
  assign n19231 = n17660 & ~n19230 ;
  assign n19232 = ~n19228 & n19231 ;
  assign n19233 = n9948 & n19232 ;
  assign n19234 = ~n19217 & n19233 ;
  assign n19235 = n19221 & n19226 ;
  assign n19236 = n17420 & ~n18907 ;
  assign n19237 = n17720 & ~n19236 ;
  assign n19238 = ~n19235 & n19237 ;
  assign n19239 = ~\pi0185  & ~\pi0299  ;
  assign n19240 = ~\pi0150  & \pi0299  ;
  assign n19241 = ~n19239 & ~n19240 ;
  assign n19242 = n8640 & n19241 ;
  assign n19243 = \pi0087  & ~n19242 ;
  assign n19244 = ~n19238 & ~n19243 ;
  assign n19245 = n9948 & ~n19244 ;
  assign n19246 = ~\pi0232  & ~n17420 ;
  assign n19247 = ~\pi0232  & ~n18902 ;
  assign n19248 = ~n18906 & n19247 ;
  assign n19249 = ~n19246 & ~n19248 ;
  assign n19250 = n18907 & n18941 ;
  assign n19251 = ~\pi0087  & n18772 ;
  assign n19252 = n15926 & ~n18938 ;
  assign n19253 = ~n19251 & ~n19252 ;
  assign n19254 = ~n19250 & ~n19253 ;
  assign n19255 = n19249 & n19254 ;
  assign n19256 = \pi0087  & n16572 ;
  assign n19257 = ~n9948 & ~n19256 ;
  assign n19258 = ~n19255 & n19257 ;
  assign n19259 = ~n19245 & ~n19258 ;
  assign n19260 = ~n19234 & n19259 ;
  assign n19261 = \pi0129  & n2404 ;
  assign n19262 = n2403 & n19261 ;
  assign n19263 = n1281 & n19262 ;
  assign n19264 = n1260 & n19263 ;
  assign n19265 = ~n1292 & ~n19264 ;
  assign n19266 = n2467 & ~n19265 ;
  assign n19267 = \pi0129  & ~n2467 ;
  assign n19268 = n8438 & n19267 ;
  assign n19269 = n1281 & n19268 ;
  assign n19270 = n1260 & n19269 ;
  assign n19271 = ~n19266 & ~n19270 ;
  assign n19272 = \pi0054  & \pi0129  ;
  assign n19273 = n2364 & n19272 ;
  assign n19274 = n2342 & n19273 ;
  assign n19275 = n1281 & n19274 ;
  assign n19276 = n1260 & n19275 ;
  assign n19277 = ~\pi0074  & ~n19276 ;
  assign n19278 = ~\pi0056  & n2404 ;
  assign n19279 = ~\pi0038  & \pi0129  ;
  assign n19280 = n2362 & n19279 ;
  assign n19281 = n1354 & n19280 ;
  assign n19282 = n8413 & n19281 ;
  assign n19283 = n1358 & n19282 ;
  assign n19284 = ~\pi0054  & ~\pi0055  ;
  assign n19285 = n2364 & n19284 ;
  assign n19286 = ~\pi0056  & n19285 ;
  assign n19287 = n19283 & n19286 ;
  assign n19288 = ~n19278 & ~n19287 ;
  assign n19289 = ~n19277 & ~n19288 ;
  assign n19290 = \pi0039  & \pi0129  ;
  assign n19291 = n1281 & n19290 ;
  assign n19292 = n1260 & n19291 ;
  assign n19293 = ~n2590 & ~n19292 ;
  assign n19294 = ~n1629 & ~n1963 ;
  assign n19295 = ~n1571 & ~n1574 ;
  assign n19296 = \pi0086  & n19295 ;
  assign n19297 = n1546 & n10306 ;
  assign n19298 = n1253 & n1504 ;
  assign n19299 = ~n1507 & n19298 ;
  assign n19300 = ~n1503 & n19299 ;
  assign n19301 = ~n1537 & n1551 ;
  assign n19302 = ~n19300 & n19301 ;
  assign n19303 = n1557 & n10306 ;
  assign n19304 = ~n19302 & n19303 ;
  assign n19305 = ~n19297 & ~n19304 ;
  assign n19306 = ~n7055 & n19295 ;
  assign n19307 = n19305 & n19306 ;
  assign n19308 = ~n19296 & ~n19307 ;
  assign n19309 = \pi0097  & ~n1571 ;
  assign n19310 = \pi0250  & \pi0252  ;
  assign n19311 = ~n6808 & n19310 ;
  assign n19312 = ~n8641 & n19311 ;
  assign n19313 = ~\pi0127  & ~n19312 ;
  assign n19314 = n8604 & n19312 ;
  assign n19315 = ~n19313 & ~n19314 ;
  assign n19316 = ~n1571 & n1580 ;
  assign n19317 = n19315 & n19316 ;
  assign n19318 = ~n19309 & ~n19317 ;
  assign n19319 = ~n1587 & n1588 ;
  assign n19320 = n19318 & n19319 ;
  assign n19321 = n19308 & n19320 ;
  assign n19322 = ~n1598 & n2034 ;
  assign n19323 = ~n19321 & n19322 ;
  assign n19324 = ~n1400 & n10533 ;
  assign n19325 = ~n2043 & n19324 ;
  assign n19326 = ~n19323 & n19325 ;
  assign n19327 = ~n1858 & n7083 ;
  assign n19328 = ~n1360 & ~n1831 ;
  assign n19329 = ~n1864 & n19328 ;
  assign n19330 = ~n19327 & n19329 ;
  assign n19331 = ~n19326 & n19330 ;
  assign n19332 = ~\pi0035  & \pi0070  ;
  assign n19333 = n1354 & n19332 ;
  assign n19334 = n1358 & n19333 ;
  assign n19335 = ~\pi0051  & ~n19334 ;
  assign n19336 = ~n19331 & n19335 ;
  assign n19337 = n2569 & ~n19336 ;
  assign n19338 = ~n19294 & ~n19337 ;
  assign n19339 = n1634 & ~n19292 ;
  assign n19340 = n19338 & n19339 ;
  assign n19341 = ~n19293 & ~n19340 ;
  assign n19342 = ~\pi0038  & ~\pi0095  ;
  assign n19343 = ~n19341 & n19342 ;
  assign n19344 = ~\pi0039  & \pi0129  ;
  assign n19345 = ~n1639 & n19344 ;
  assign n19346 = ~\pi0038  & ~n19292 ;
  assign n19347 = ~n19345 & n19346 ;
  assign n19348 = n1288 & ~n13206 ;
  assign n19349 = \pi0129  & n19348 ;
  assign n19350 = n1281 & n19349 ;
  assign n19351 = n1260 & n19350 ;
  assign n19352 = ~n2362 & ~n19351 ;
  assign n19353 = ~\pi0075  & ~n19352 ;
  assign n19354 = \pi0129  & n4520 ;
  assign n19355 = n1638 & n19354 ;
  assign n19356 = \pi0038  & ~n19355 ;
  assign n19357 = n19353 & ~n19356 ;
  assign n19358 = ~n19347 & n19357 ;
  assign n19359 = ~n19343 & n19358 ;
  assign n19360 = ~\pi0075  & ~n2362 ;
  assign n19361 = n19351 & n19360 ;
  assign n19362 = \pi0075  & n19283 ;
  assign n19363 = ~\pi0092  & ~n19362 ;
  assign n19364 = ~n19361 & n19363 ;
  assign n19365 = ~n19359 & n19364 ;
  assign n19366 = \pi0092  & ~\pi0129  ;
  assign n19367 = ~\pi0054  & ~n19366 ;
  assign n19368 = ~n8420 & n19367 ;
  assign n19369 = ~n19288 & n19368 ;
  assign n19370 = ~n19365 & n19369 ;
  assign n19371 = ~n19289 & ~n19370 ;
  assign n19372 = ~\pi0056  & n13442 ;
  assign n19373 = n19283 & n19372 ;
  assign n19374 = ~n13452 & ~n13466 ;
  assign n19375 = ~n19270 & n19374 ;
  assign n19376 = ~n19373 & n19375 ;
  assign n19377 = n19371 & n19376 ;
  assign n19378 = ~n19271 & ~n19377 ;
  assign n19379 = n6787 & n10071 ;
  assign n19380 = n1354 & n19379 ;
  assign n19381 = n1358 & n19380 ;
  assign n19382 = ~\pi0087  & ~n19381 ;
  assign n19383 = n6693 & n19382 ;
  assign n19384 = ~\pi0038  & ~n2596 ;
  assign n19385 = n19382 & n19384 ;
  assign n19386 = ~n2594 & n19385 ;
  assign n19387 = ~n19383 & ~n19386 ;
  assign n19388 = ~n16294 & n19387 ;
  assign n19389 = ~n6808 & n12104 ;
  assign n19390 = ~n8641 & n19389 ;
  assign n19391 = \pi0129  & n10094 ;
  assign n19392 = n10093 & n19391 ;
  assign n19393 = ~n19390 & n19392 ;
  assign n19394 = ~n8604 & n13136 ;
  assign n19395 = n19390 & n19394 ;
  assign n19396 = ~n19393 & ~n19395 ;
  assign n19397 = n2280 & ~n19396 ;
  assign n19398 = n1285 & ~n19397 ;
  assign n19399 = n2404 & n19398 ;
  assign n19400 = ~n19388 & n19399 ;
  assign n19401 = \pi0074  & ~n8430 ;
  assign n19402 = ~n16288 & ~n19401 ;
  assign n19403 = ~n6834 & ~n16284 ;
  assign n19404 = ~n8412 & ~n8420 ;
  assign n19405 = n2404 & ~n19404 ;
  assign n19406 = n19403 & ~n19405 ;
  assign n19407 = n19402 & n19406 ;
  assign n19408 = ~n19400 & n19407 ;
  assign n19409 = ~n1292 & n19403 ;
  assign n19410 = n2467 & ~n19409 ;
  assign n19411 = ~n19408 & n19410 ;
  assign n19412 = ~n8441 & ~n19411 ;
  assign n19413 = ~\pi0132  & n18904 ;
  assign n19414 = \pi0130  & ~n19413 ;
  assign n19415 = ~\pi0136  & n17435 ;
  assign n19416 = ~\pi0130  & ~n19415 ;
  assign n19417 = n19413 & n19416 ;
  assign n19418 = ~n19414 & ~n19417 ;
  assign n19419 = ~\pi0087  & n17419 ;
  assign n19420 = n19418 & n19419 ;
  assign n19421 = n10138 & ~n17419 ;
  assign n19422 = ~\pi0051  & ~n19421 ;
  assign n19423 = ~\pi0087  & ~n19422 ;
  assign n19424 = \pi0087  & n11140 ;
  assign n19425 = ~n9948 & ~n19424 ;
  assign n19426 = ~n19423 & n19425 ;
  assign n19427 = ~n19420 & n19426 ;
  assign n19428 = \pi0087  & ~n11492 ;
  assign n19429 = ~n17444 & n19428 ;
  assign n19430 = n8640 & ~n10150 ;
  assign n19431 = n17507 & ~n19430 ;
  assign n19432 = ~n18941 & ~n19431 ;
  assign n19433 = ~n17444 & n17720 ;
  assign n19434 = ~n19432 & n19433 ;
  assign n19435 = ~n19429 & ~n19434 ;
  assign n19436 = n19418 & n19435 ;
  assign n19437 = n9948 & ~n19436 ;
  assign n19438 = ~\pi0038  & n11040 ;
  assign n19439 = \pi0039  & ~\pi0051  ;
  assign n19440 = ~\pi0038  & n19439 ;
  assign n19441 = n18192 & n19440 ;
  assign n19442 = ~n19438 & ~n19441 ;
  assign n19443 = ~\pi0051  & ~n9627 ;
  assign n19444 = ~n17419 & n19443 ;
  assign n19445 = ~n19430 & n19444 ;
  assign n19446 = ~\pi0100  & ~n19445 ;
  assign n19447 = n19442 & n19446 ;
  assign n19448 = n11633 & ~n19445 ;
  assign n19449 = ~n19447 & ~n19448 ;
  assign n19450 = ~\pi0191  & ~\pi0299  ;
  assign n19451 = ~\pi0051  & n18187 ;
  assign n19452 = n17751 & n19451 ;
  assign n19453 = ~n17507 & ~n19452 ;
  assign n19454 = n19450 & n19453 ;
  assign n19455 = \pi0140  & n19450 ;
  assign n19456 = n18250 & n19455 ;
  assign n19457 = ~n19454 & ~n19456 ;
  assign n19458 = \pi0140  & ~\pi0287  ;
  assign n19459 = n6706 & n19458 ;
  assign n19460 = ~\pi0051  & ~n19459 ;
  assign n19461 = ~n18273 & n19460 ;
  assign n19462 = ~n18267 & n19461 ;
  assign n19463 = n10148 & ~n19462 ;
  assign n19464 = n19457 & ~n19463 ;
  assign n19465 = ~\pi0051  & ~n6706 ;
  assign n19466 = ~n17953 & n19465 ;
  assign n19467 = n1354 & n17503 ;
  assign n19468 = n17942 & n19467 ;
  assign n19469 = n1358 & n19468 ;
  assign n19470 = ~n19466 & ~n19469 ;
  assign n19471 = ~\pi0051  & ~n17627 ;
  assign n19472 = n17636 & n19471 ;
  assign n19473 = ~n17507 & ~n19472 ;
  assign n19474 = ~\pi0169  & n19473 ;
  assign n19475 = \pi0162  & \pi0216  ;
  assign n19476 = n6936 & n19475 ;
  assign n19477 = ~n17627 & n19476 ;
  assign n19478 = ~n19474 & n19477 ;
  assign n19479 = ~n19470 & n19478 ;
  assign n19480 = ~\pi0169  & n19475 ;
  assign n19481 = n6936 & n19480 ;
  assign n19482 = ~n19473 & n19481 ;
  assign n19483 = \pi0169  & n6706 ;
  assign n19484 = \pi0051  & ~n19483 ;
  assign n19485 = n17420 & ~n19483 ;
  assign n19486 = ~n17636 & n19485 ;
  assign n19487 = ~n19484 & ~n19486 ;
  assign n19488 = ~\pi0162  & \pi0216  ;
  assign n19489 = n6936 & n19488 ;
  assign n19490 = ~n19483 & n19489 ;
  assign n19491 = n1281 & n19489 ;
  assign n19492 = n1260 & n19491 ;
  assign n19493 = ~n19490 & ~n19492 ;
  assign n19494 = n19487 & ~n19493 ;
  assign n19495 = ~n7597 & ~n19483 ;
  assign n19496 = n17507 & n19495 ;
  assign n19497 = \pi0299  & ~n19496 ;
  assign n19498 = ~n19494 & n19497 ;
  assign n19499 = ~n19482 & n19498 ;
  assign n19500 = ~n19479 & n19499 ;
  assign n19501 = ~n19447 & ~n19500 ;
  assign n19502 = n19464 & n19501 ;
  assign n19503 = ~n19449 & ~n19502 ;
  assign n19504 = \pi0100  & n19432 ;
  assign n19505 = n18041 & ~n19504 ;
  assign n19506 = n9948 & n19505 ;
  assign n19507 = ~n19503 & n19506 ;
  assign n19508 = ~n19437 & ~n19507 ;
  assign n19509 = ~n19427 & n19508 ;
  assign n19510 = n17660 & ~n19504 ;
  assign n19511 = n17943 & ~n18456 ;
  assign n19512 = n1358 & n19511 ;
  assign n19513 = ~\pi0232  & n19439 ;
  assign n19514 = ~n19512 & n19513 ;
  assign n19515 = ~\pi0051  & ~\pi0169  ;
  assign n19516 = ~n17672 & n19515 ;
  assign n19517 = ~\pi0051  & \pi0169  ;
  assign n19518 = n17419 & n19517 ;
  assign n19519 = ~n6706 & n19517 ;
  assign n19520 = ~n19518 & ~n19519 ;
  assign n19521 = \pi0216  & n19520 ;
  assign n19522 = \pi0216  & n17627 ;
  assign n19523 = n17636 & n19522 ;
  assign n19524 = ~n19521 & ~n19523 ;
  assign n19525 = \pi0162  & ~n19524 ;
  assign n19526 = ~n19516 & n19525 ;
  assign n19527 = ~\pi0216  & ~n19483 ;
  assign n19528 = ~n17945 & n19527 ;
  assign n19529 = ~\pi0216  & n19483 ;
  assign n19530 = ~n17953 & n19529 ;
  assign n19531 = ~n17419 & n19483 ;
  assign n19532 = ~\pi0051  & ~n19531 ;
  assign n19533 = n6936 & ~n19488 ;
  assign n19534 = ~n19532 & ~n19533 ;
  assign n19535 = ~n19530 & ~n19534 ;
  assign n19536 = ~n19528 & n19535 ;
  assign n19537 = ~n19526 & n19536 ;
  assign n19538 = n17987 & ~n19531 ;
  assign n19539 = \pi0299  & ~n19538 ;
  assign n19540 = ~n19537 & n19539 ;
  assign n19541 = n1354 & n6949 ;
  assign n19542 = n17942 & n19541 ;
  assign n19543 = n1358 & n19542 ;
  assign n19544 = ~\pi0051  & \pi0140  ;
  assign n19545 = ~n19543 & n19544 ;
  assign n19546 = n18496 & n19544 ;
  assign n19547 = ~n17672 & n19546 ;
  assign n19548 = ~n19545 & ~n19547 ;
  assign n19549 = ~\pi0051  & ~\pi0140  ;
  assign n19550 = ~n18526 & n19549 ;
  assign n19551 = n19450 & ~n19550 ;
  assign n19552 = n19548 & n19551 ;
  assign n19553 = ~n19540 & ~n19552 ;
  assign n19554 = n19439 & ~n19512 ;
  assign n19555 = ~n11040 & ~n19554 ;
  assign n19556 = n6706 & n8701 ;
  assign n19557 = ~n17953 & n19556 ;
  assign n19558 = ~n6706 & n8701 ;
  assign n19559 = ~n17945 & n19558 ;
  assign n19560 = ~n19557 & ~n19559 ;
  assign n19561 = n17627 & n17636 ;
  assign n19562 = ~n17421 & ~n18499 ;
  assign n19563 = ~n19561 & n19562 ;
  assign n19564 = n18185 & ~n19563 ;
  assign n19565 = \pi0051  & ~n6949 ;
  assign n19566 = n6706 & ~n6949 ;
  assign n19567 = ~n17419 & n19566 ;
  assign n19568 = ~n19565 & ~n19567 ;
  assign n19569 = \pi0140  & n19568 ;
  assign n19570 = ~n19564 & n19569 ;
  assign n19571 = n19560 & n19570 ;
  assign n19572 = ~\pi0140  & n8701 ;
  assign n19573 = ~n17504 & n19549 ;
  assign n19574 = ~n19572 & ~n19573 ;
  assign n19575 = ~n19557 & ~n19574 ;
  assign n19576 = ~n19559 & n19575 ;
  assign n19577 = n10148 & ~n19576 ;
  assign n19578 = ~n19571 & n19577 ;
  assign n19579 = ~n19555 & ~n19578 ;
  assign n19580 = n19553 & n19579 ;
  assign n19581 = ~n19514 & ~n19580 ;
  assign n19582 = ~\pi0038  & ~n19581 ;
  assign n19583 = ~n10150 & n18767 ;
  assign n19584 = ~n17746 & n19465 ;
  assign n19585 = ~n10150 & n19584 ;
  assign n19586 = ~n17462 & n19585 ;
  assign n19587 = ~n19583 & ~n19586 ;
  assign n19588 = ~\pi0051  & n10150 ;
  assign n19589 = ~n17746 & n19588 ;
  assign n19590 = ~n17462 & n19589 ;
  assign n19591 = \pi0232  & ~n19590 ;
  assign n19592 = n19587 & n19591 ;
  assign n19593 = ~\pi0039  & n17808 ;
  assign n19594 = ~n17462 & n19593 ;
  assign n19595 = ~n17620 & ~n19594 ;
  assign n19596 = ~\pi0038  & ~n19595 ;
  assign n19597 = ~n19592 & n19596 ;
  assign n19598 = \pi0038  & ~n19432 ;
  assign n19599 = ~\pi0100  & ~n19598 ;
  assign n19600 = ~n19597 & n19599 ;
  assign n19601 = ~n19582 & n19600 ;
  assign n19602 = n19510 & ~n19601 ;
  assign n19603 = n17720 & ~n19432 ;
  assign n19604 = ~n19418 & ~n19428 ;
  assign n19605 = ~n19603 & n19604 ;
  assign n19606 = ~n19427 & n19605 ;
  assign n19607 = ~n19602 & n19606 ;
  assign n19608 = ~n19509 & ~n19607 ;
  assign n19609 = ~n8420 & n12970 ;
  assign n19610 = n8601 & ~n16849 ;
  assign n19611 = ~\pi0075  & \pi0087  ;
  assign n19612 = ~\pi0075  & \pi0100  ;
  assign n19613 = ~n8404 & n19612 ;
  assign n19614 = ~n19611 & ~n19613 ;
  assign n19615 = ~n8417 & n19614 ;
  assign n19616 = ~n19610 & n19615 ;
  assign n19617 = ~\pi0092  & ~n19616 ;
  assign n19618 = n19609 & ~n19617 ;
  assign n19619 = ~\pi0051  & ~\pi0168  ;
  assign n19620 = \pi0051  & ~\pi0151  ;
  assign n19621 = n6706 & ~n19620 ;
  assign n19622 = ~n19619 & n19621 ;
  assign n19623 = ~n17420 & n19622 ;
  assign n19624 = \pi0299  & ~n19623 ;
  assign n19625 = ~\pi0051  & \pi0190  ;
  assign n19626 = n6706 & n19625 ;
  assign n19627 = ~n17419 & n19626 ;
  assign n19628 = \pi0051  & \pi0173  ;
  assign n19629 = n6706 & n19628 ;
  assign n19630 = ~\pi0299  & ~n19629 ;
  assign n19631 = ~n19627 & n19630 ;
  assign n19632 = \pi0232  & ~n2327 ;
  assign n19633 = ~n19631 & n19632 ;
  assign n19634 = ~n19624 & n19633 ;
  assign n19635 = ~\pi0132  & n17437 ;
  assign n19636 = \pi0132  & ~n18904 ;
  assign n19637 = ~n19413 & ~n19636 ;
  assign n19638 = ~n19635 & ~n19637 ;
  assign n19639 = \pi0087  & ~n10106 ;
  assign n19640 = ~n19638 & ~n19639 ;
  assign n19641 = n9948 & ~n19640 ;
  assign n19642 = \pi0232  & ~n19631 ;
  assign n19643 = ~n19624 & n19642 ;
  assign n19644 = n9948 & n17732 ;
  assign n19645 = ~n19643 & n19644 ;
  assign n19646 = ~n19641 & ~n19645 ;
  assign n19647 = ~\pi0168  & ~n6706 ;
  assign n19648 = ~n16662 & ~n19619 ;
  assign n19649 = ~n19647 & n19648 ;
  assign n19650 = \pi0149  & ~n17420 ;
  assign n19651 = \pi0149  & ~n17627 ;
  assign n19652 = n17636 & n19651 ;
  assign n19653 = ~n19650 & ~n19652 ;
  assign n19654 = ~n19649 & ~n19653 ;
  assign n19655 = \pi0168  & n17954 ;
  assign n19656 = n16352 & ~n17945 ;
  assign n19657 = ~n19655 & ~n19656 ;
  assign n19658 = \pi0149  & n19620 ;
  assign n19659 = \pi0149  & ~n17741 ;
  assign n19660 = ~n17672 & n19659 ;
  assign n19661 = ~n19658 & ~n19660 ;
  assign n19662 = ~n19657 & ~n19661 ;
  assign n19663 = ~n19654 & ~n19662 ;
  assign n19664 = \pi0168  & ~n6706 ;
  assign n19665 = ~n17953 & n19664 ;
  assign n19666 = \pi0168  & n17956 ;
  assign n19667 = ~n19665 & ~n19666 ;
  assign n19668 = ~\pi0168  & ~n17741 ;
  assign n19669 = ~n17953 & n19668 ;
  assign n19670 = \pi0151  & ~n19669 ;
  assign n19671 = n19667 & n19670 ;
  assign n19672 = ~\pi0151  & n16352 ;
  assign n19673 = ~\pi0151  & n17420 ;
  assign n19674 = ~n17636 & n19673 ;
  assign n19675 = ~n19672 & ~n19674 ;
  assign n19676 = ~\pi0149  & n19675 ;
  assign n19677 = ~\pi0149  & n16352 ;
  assign n19678 = ~n17945 & n19677 ;
  assign n19679 = ~n19676 & ~n19678 ;
  assign n19680 = ~n19671 & ~n19679 ;
  assign n19681 = n7597 & ~n19680 ;
  assign n19682 = n19663 & n19681 ;
  assign n19683 = \pi0299  & ~n17420 ;
  assign n19684 = ~n19623 & n19683 ;
  assign n19685 = ~n11062 & ~n19684 ;
  assign n19686 = \pi0232  & ~n19685 ;
  assign n19687 = ~n19682 & n19686 ;
  assign n19688 = \pi0173  & \pi0183  ;
  assign n19689 = \pi0173  & ~n19136 ;
  assign n19690 = ~n18255 & n19689 ;
  assign n19691 = ~n19688 & ~n19690 ;
  assign n19692 = \pi0183  & ~n18237 ;
  assign n19693 = ~n18240 & n19692 ;
  assign n19694 = \pi0190  & ~\pi0299  ;
  assign n19695 = \pi0183  & ~n6955 ;
  assign n19696 = ~n19135 & n19695 ;
  assign n19697 = n19694 & ~n19696 ;
  assign n19698 = ~n19693 & n19697 ;
  assign n19699 = ~n19691 & n19698 ;
  assign n19700 = \pi0183  & n18268 ;
  assign n19701 = ~\pi0173  & ~n19700 ;
  assign n19702 = ~n18273 & n19694 ;
  assign n19703 = n19701 & n19702 ;
  assign n19704 = ~n18267 & n19703 ;
  assign n19705 = ~\pi0190  & ~\pi0299  ;
  assign n19706 = ~n19629 & n19705 ;
  assign n19707 = n17420 & ~n18188 ;
  assign n19708 = ~\pi0051  & \pi0183  ;
  assign n19709 = n17419 & n19708 ;
  assign n19710 = ~n18205 & n19709 ;
  assign n19711 = ~n19707 & ~n19710 ;
  assign n19712 = n19706 & n19711 ;
  assign n19713 = ~n19704 & ~n19712 ;
  assign n19714 = ~n19699 & n19713 ;
  assign n19715 = \pi0232  & ~n19714 ;
  assign n19716 = n12343 & ~n18193 ;
  assign n19717 = ~n19715 & n19716 ;
  assign n19718 = ~n19687 & n19717 ;
  assign n19719 = n17420 & n17938 ;
  assign n19720 = ~n17514 & n19719 ;
  assign n19721 = \pi0182  & n6706 ;
  assign n19722 = n19162 & n19721 ;
  assign n19723 = n17420 & n19162 ;
  assign n19724 = ~n17514 & n19723 ;
  assign n19725 = ~n19722 & ~n19724 ;
  assign n19726 = ~n17515 & n19706 ;
  assign n19727 = n19725 & n19726 ;
  assign n19728 = \pi0232  & ~n19727 ;
  assign n19729 = ~\pi0182  & n15942 ;
  assign n19730 = n17544 & n19729 ;
  assign n19731 = n19694 & n19730 ;
  assign n19732 = \pi0051  & ~\pi0173  ;
  assign n19733 = n6706 & ~n19732 ;
  assign n19734 = n19694 & ~n19733 ;
  assign n19735 = ~n17515 & n19734 ;
  assign n19736 = ~n19731 & ~n19735 ;
  assign n19737 = ~\pi0039  & n19736 ;
  assign n19738 = n19728 & n19737 ;
  assign n19739 = ~n19720 & ~n19738 ;
  assign n19740 = n6706 & n19620 ;
  assign n19741 = \pi0168  & ~n19740 ;
  assign n19742 = ~n17704 & n19741 ;
  assign n19743 = ~\pi0160  & n17420 ;
  assign n19744 = ~n17514 & n19743 ;
  assign n19745 = ~n14157 & ~n19744 ;
  assign n19746 = n19742 & ~n19745 ;
  assign n19747 = \pi0151  & ~n17505 ;
  assign n19748 = ~n17528 & n19747 ;
  assign n19749 = ~\pi0168  & n17420 ;
  assign n19750 = ~n17514 & n19749 ;
  assign n19751 = ~n16337 & ~n19750 ;
  assign n19752 = ~n19745 & ~n19751 ;
  assign n19753 = ~n19748 & n19752 ;
  assign n19754 = ~n19746 & ~n19753 ;
  assign n19755 = ~\pi0151  & ~n19623 ;
  assign n19756 = ~n6706 & n19755 ;
  assign n19757 = n17514 & n19756 ;
  assign n19758 = ~\pi0151  & ~n17420 ;
  assign n19759 = ~n19622 & n19758 ;
  assign n19760 = \pi0160  & ~n19759 ;
  assign n19761 = ~n19757 & n19760 ;
  assign n19762 = n6706 & n19619 ;
  assign n19763 = ~n17419 & n19762 ;
  assign n19764 = n17420 & ~n19763 ;
  assign n19765 = ~n17514 & n19764 ;
  assign n19766 = n6706 & ~n19763 ;
  assign n19767 = \pi0151  & ~n19766 ;
  assign n19768 = ~n19765 & n19767 ;
  assign n19769 = n19761 & ~n19768 ;
  assign n19770 = \pi0299  & ~n19769 ;
  assign n19771 = ~n19720 & n19770 ;
  assign n19772 = n19754 & n19771 ;
  assign n19773 = ~n19739 & ~n19772 ;
  assign n19774 = n2327 & n19773 ;
  assign n19775 = ~\pi0051  & ~n2327 ;
  assign n19776 = n17419 & n19775 ;
  assign n19777 = n17660 & ~n19776 ;
  assign n19778 = n9948 & n19777 ;
  assign n19779 = ~n19634 & n19778 ;
  assign n19780 = ~n19774 & n19779 ;
  assign n19781 = ~n19718 & n19780 ;
  assign n19782 = n19646 & ~n19781 ;
  assign n19783 = ~n19634 & ~n19782 ;
  assign n19784 = ~\pi0151  & n2575 ;
  assign n19785 = ~n1629 & n19784 ;
  assign n19786 = ~\pi0168  & ~n19785 ;
  assign n19787 = ~\pi0072  & ~\pi0168  ;
  assign n19788 = ~n17815 & n19787 ;
  assign n19789 = ~n19786 & ~n19788 ;
  assign n19790 = n2575 & ~n6706 ;
  assign n19791 = ~n1629 & n19790 ;
  assign n19792 = \pi0160  & ~n19791 ;
  assign n19793 = ~\pi0072  & \pi0160  ;
  assign n19794 = ~n17835 & n19793 ;
  assign n19795 = ~n19792 & ~n19794 ;
  assign n19796 = \pi0151  & ~n17809 ;
  assign n19797 = ~n19795 & ~n19796 ;
  assign n19798 = ~n19789 & n19797 ;
  assign n19799 = ~\pi0072  & ~n6706 ;
  assign n19800 = ~n17835 & n19799 ;
  assign n19801 = ~n2575 & ~n6706 ;
  assign n19802 = ~n1628 & n18591 ;
  assign n19803 = ~n19801 & ~n19802 ;
  assign n19804 = ~n18643 & n19803 ;
  assign n19805 = ~n19800 & n19804 ;
  assign n19806 = \pi0168  & ~n19805 ;
  assign n19807 = ~\pi0168  & ~n17799 ;
  assign n19808 = ~n17828 & n19807 ;
  assign n19809 = \pi0151  & ~n19808 ;
  assign n19810 = ~\pi0072  & ~n17835 ;
  assign n19811 = \pi0151  & n19791 ;
  assign n19812 = ~n19810 & n19811 ;
  assign n19813 = ~n19809 & ~n19812 ;
  assign n19814 = ~n19806 & ~n19813 ;
  assign n19815 = \pi0151  & ~\pi0160  ;
  assign n19816 = \pi0168  & ~n17846 ;
  assign n19817 = ~\pi0160  & ~n19816 ;
  assign n19818 = n2575 & ~n16352 ;
  assign n19819 = ~n1629 & n19818 ;
  assign n19820 = ~n19810 & n19819 ;
  assign n19821 = n19817 & ~n19820 ;
  assign n19822 = ~n19815 & ~n19821 ;
  assign n19823 = ~n19814 & ~n19822 ;
  assign n19824 = ~\pi0168  & n6706 ;
  assign n19825 = ~n17755 & n19621 ;
  assign n19826 = ~n19824 & ~n19825 ;
  assign n19827 = ~n19795 & n19826 ;
  assign n19828 = ~n19823 & ~n19827 ;
  assign n19829 = ~n19798 & n19828 ;
  assign n19830 = n10276 & ~n19829 ;
  assign n19831 = \pi0182  & n13001 ;
  assign n19832 = n17491 & n19831 ;
  assign n19833 = n17495 & n19832 ;
  assign n19834 = n17480 & n19833 ;
  assign n19835 = n17842 & ~n19834 ;
  assign n19836 = ~n17750 & n19835 ;
  assign n19837 = n19733 & ~n19836 ;
  assign n19838 = n19694 & ~n19837 ;
  assign n19839 = ~\pi0173  & ~n2575 ;
  assign n19840 = \pi0072  & ~\pi0173  ;
  assign n19841 = ~n1628 & n19840 ;
  assign n19842 = ~n19839 & ~n19841 ;
  assign n19843 = ~\pi0072  & ~\pi0173  ;
  assign n19844 = ~n17815 & n19843 ;
  assign n19845 = n19842 & ~n19844 ;
  assign n19846 = ~\pi0051  & \pi0173  ;
  assign n19847 = ~n17746 & n19846 ;
  assign n19848 = ~n17462 & n19847 ;
  assign n19849 = n19721 & ~n19848 ;
  assign n19850 = n19845 & n19849 ;
  assign n19851 = ~n17835 & n19843 ;
  assign n19852 = n19842 & ~n19851 ;
  assign n19853 = \pi0173  & ~n6706 ;
  assign n19854 = \pi0173  & ~n17741 ;
  assign n19855 = ~n17746 & n19854 ;
  assign n19856 = ~n19853 & ~n19855 ;
  assign n19857 = ~\pi0182  & n19856 ;
  assign n19858 = ~\pi0182  & n17558 ;
  assign n19859 = ~n17827 & n19858 ;
  assign n19860 = ~n19857 & ~n19859 ;
  assign n19861 = n19852 & ~n19860 ;
  assign n19862 = n19705 & ~n19861 ;
  assign n19863 = ~n19850 & n19862 ;
  assign n19864 = ~n19838 & ~n19863 ;
  assign n19865 = \pi0232  & ~n19791 ;
  assign n19866 = n15771 & ~n17835 ;
  assign n19867 = ~n19865 & ~n19866 ;
  assign n19868 = ~n19864 & ~n19867 ;
  assign n19869 = ~\pi0072  & ~\pi0232  ;
  assign n19870 = ~n17835 & n19869 ;
  assign n19871 = ~\pi0232  & ~n2575 ;
  assign n19872 = ~n1628 & n12503 ;
  assign n19873 = ~n19871 & ~n19872 ;
  assign n19874 = n13268 & n19873 ;
  assign n19875 = ~n19870 & n19874 ;
  assign n19876 = ~n19868 & n19875 ;
  assign n19877 = ~n19830 & n19876 ;
  assign n19878 = n12383 & n18458 ;
  assign n19879 = ~\pi0183  & ~n8701 ;
  assign n19880 = ~n17421 & n19879 ;
  assign n19881 = \pi0173  & n8701 ;
  assign n19882 = ~n18471 & n19881 ;
  assign n19883 = ~n18476 & n19882 ;
  assign n19884 = n18488 & n19688 ;
  assign n19885 = ~n19883 & ~n19884 ;
  assign n19886 = ~n19880 & n19885 ;
  assign n19887 = n19694 & ~n19886 ;
  assign n19888 = ~\pi0149  & \pi0216  ;
  assign n19889 = n6936 & ~n19888 ;
  assign n19890 = n19623 & ~n19889 ;
  assign n19891 = \pi0299  & ~n19890 ;
  assign n19892 = \pi0168  & ~n18471 ;
  assign n19893 = ~n18476 & n19892 ;
  assign n19894 = ~n17944 & n19619 ;
  assign n19895 = \pi0051  & ~\pi0168  ;
  assign n19896 = ~n6706 & n19895 ;
  assign n19897 = n6936 & ~n19896 ;
  assign n19898 = ~n19620 & n19897 ;
  assign n19899 = ~n19894 & n19898 ;
  assign n19900 = ~n19893 & n19899 ;
  assign n19901 = ~n7597 & ~n19900 ;
  assign n19902 = n19891 & n19901 ;
  assign n19903 = ~\pi0168  & ~n18558 ;
  assign n19904 = \pi0168  & n17421 ;
  assign n19905 = \pi0168  & n17627 ;
  assign n19906 = n17636 & n19905 ;
  assign n19907 = ~n19904 & ~n19906 ;
  assign n19908 = \pi0151  & n19907 ;
  assign n19909 = ~n19903 & n19908 ;
  assign n19910 = \pi0168  & ~n17641 ;
  assign n19911 = ~n17640 & n19910 ;
  assign n19912 = ~n17639 & n19911 ;
  assign n19913 = ~\pi0168  & ~\pi0287  ;
  assign n19914 = n6706 & n19913 ;
  assign n19915 = n1281 & n19914 ;
  assign n19916 = n1260 & n19915 ;
  assign n19917 = ~\pi0151  & ~n19916 ;
  assign n19918 = ~n19912 & n19917 ;
  assign n19919 = \pi0149  & ~n19918 ;
  assign n19920 = ~n19909 & n19919 ;
  assign n19921 = \pi0216  & n19891 ;
  assign n19922 = ~n19920 & n19921 ;
  assign n19923 = ~n19902 & ~n19922 ;
  assign n19924 = ~n19887 & n19923 ;
  assign n19925 = ~n17968 & ~n18913 ;
  assign n19926 = \pi0183  & ~n19925 ;
  assign n19927 = ~\pi0173  & \pi0183  ;
  assign n19928 = ~\pi0173  & ~n18471 ;
  assign n19929 = ~n18469 & n19928 ;
  assign n19930 = ~n19927 & ~n19929 ;
  assign n19931 = n19694 & ~n19930 ;
  assign n19932 = ~n19926 & n19931 ;
  assign n19933 = ~\pi0173  & ~\pi0223  ;
  assign n19934 = n6148 & n19933 ;
  assign n19935 = ~n19927 & ~n19934 ;
  assign n19936 = ~n18506 & ~n19935 ;
  assign n19937 = n1281 & n19936 ;
  assign n19938 = n1260 & n19937 ;
  assign n19939 = n19705 & ~n19938 ;
  assign n19940 = ~\pi0173  & n19939 ;
  assign n19941 = \pi0183  & n6949 ;
  assign n19942 = ~n18497 & n19941 ;
  assign n19943 = n18503 & n19942 ;
  assign n19944 = ~\pi0051  & ~\pi0183  ;
  assign n19945 = n18526 & n19944 ;
  assign n19946 = ~n17741 & ~n19945 ;
  assign n19947 = n19939 & n19946 ;
  assign n19948 = ~n19943 & n19947 ;
  assign n19949 = ~n19940 & ~n19948 ;
  assign n19950 = n18460 & n19949 ;
  assign n19951 = ~n19932 & n19950 ;
  assign n19952 = n19924 & n19951 ;
  assign n19953 = ~n19878 & ~n19952 ;
  assign n19954 = n2327 & ~n19953 ;
  assign n19955 = n17660 & ~n19954 ;
  assign n19956 = ~n19877 & n19955 ;
  assign n19957 = n19783 & n19956 ;
  assign n19958 = n17444 & ~n19638 ;
  assign n19959 = \pi0232  & ~n19619 ;
  assign n19960 = n19621 & n19959 ;
  assign n19961 = ~n17420 & n19960 ;
  assign n19962 = ~\pi0087  & n19961 ;
  assign n19963 = \pi0087  & \pi0164  ;
  assign n19964 = n8640 & n19963 ;
  assign n19965 = ~n9948 & ~n19964 ;
  assign n19966 = ~n19962 & n19965 ;
  assign n19967 = ~n19958 & n19966 ;
  assign n19968 = n17720 & ~n19643 ;
  assign n19969 = n19638 & ~n19639 ;
  assign n19970 = ~n19968 & n19969 ;
  assign n19971 = ~n19967 & n19970 ;
  assign n19972 = n19646 & ~n19967 ;
  assign n19973 = ~n19781 & n19972 ;
  assign n19974 = ~n19971 & ~n19973 ;
  assign n19975 = ~n19957 & ~n19974 ;
  assign n19976 = ~n10839 & n17518 ;
  assign n19977 = ~n17490 & n19976 ;
  assign n19978 = ~\pi0039  & ~\pi0051  ;
  assign n19979 = n17419 & n19978 ;
  assign n19980 = ~n19977 & n19979 ;
  assign n19981 = ~\pi0038  & ~n19980 ;
  assign n19982 = ~n17732 & ~n18294 ;
  assign n19983 = ~n19981 & n19982 ;
  assign n19984 = \pi0197  & ~\pi0287  ;
  assign n19985 = n6706 & n19984 ;
  assign n19986 = \pi0299  & ~n19985 ;
  assign n19987 = n18180 & n19986 ;
  assign n19988 = n17751 & n19987 ;
  assign n19989 = ~n19683 & ~n19988 ;
  assign n19990 = \pi0232  & ~n19989 ;
  assign n19991 = \pi0039  & ~n19990 ;
  assign n19992 = ~n18193 & n19991 ;
  assign n19993 = ~\pi0299  & ~n17420 ;
  assign n19994 = ~\pi0299  & n18187 ;
  assign n19995 = n17751 & n19994 ;
  assign n19996 = ~n19993 & ~n19995 ;
  assign n19997 = \pi0145  & n17420 ;
  assign n19998 = ~n18205 & n19997 ;
  assign n19999 = \pi0232  & ~n19998 ;
  assign n20000 = ~n19996 & n19999 ;
  assign n20001 = n19982 & ~n20000 ;
  assign n20002 = n19992 & n20001 ;
  assign n20003 = ~n19983 & ~n20002 ;
  assign n20004 = ~\pi0133  & ~n18149 ;
  assign n20005 = ~n17732 & ~n18041 ;
  assign n20006 = ~n20004 & ~n20005 ;
  assign n20007 = n20003 & n20006 ;
  assign n20008 = ~\pi0183  & ~\pi0299  ;
  assign n20009 = ~\pi0149  & \pi0299  ;
  assign n20010 = ~n20008 & ~n20009 ;
  assign n20011 = n8640 & n20010 ;
  assign n20012 = \pi0087  & ~n20011 ;
  assign n20013 = ~n20007 & ~n20012 ;
  assign n20014 = n9948 & ~n20013 ;
  assign n20015 = ~n6103 & ~n19985 ;
  assign n20016 = n7412 & ~n20015 ;
  assign n20017 = \pi0145  & ~\pi0299  ;
  assign n20018 = ~n18455 & ~n20017 ;
  assign n20019 = ~n18506 & ~n20018 ;
  assign n20020 = ~n20016 & ~n20019 ;
  assign n20021 = n2280 & ~n20020 ;
  assign n20022 = \pi0232  & ~n20021 ;
  assign n20023 = n18460 & ~n20022 ;
  assign n20024 = n13557 & n20023 ;
  assign n20025 = ~n7093 & n10839 ;
  assign n20026 = ~\pi0072  & n10839 ;
  assign n20027 = ~n17815 & n20026 ;
  assign n20028 = ~n20025 & ~n20027 ;
  assign n20029 = ~n10839 & ~n17794 ;
  assign n20030 = ~\pi0039  & ~n20029 ;
  assign n20031 = n13557 & n20030 ;
  assign n20032 = n20028 & n20031 ;
  assign n20033 = ~n20024 & ~n20032 ;
  assign n20034 = n9948 & ~n18149 ;
  assign n20035 = ~\pi0087  & ~\pi0133  ;
  assign n20036 = n20034 & n20035 ;
  assign n20037 = n20033 & n20036 ;
  assign n20038 = ~n20014 & ~n20037 ;
  assign n20039 = n17444 & ~n20004 ;
  assign n20040 = \pi0087  & n10178 ;
  assign n20041 = ~n9948 & ~n20040 ;
  assign n20042 = ~n20039 & n20041 ;
  assign n20043 = n20038 & ~n20042 ;
  assign n20044 = ~\pi0134  & n17419 ;
  assign n20045 = ~\pi0132  & n17436 ;
  assign n20046 = n18904 & n20045 ;
  assign n20047 = ~\pi0135  & n17419 ;
  assign n20048 = n20046 & n20047 ;
  assign n20049 = ~n20044 & ~n20048 ;
  assign n20050 = \pi0171  & \pi0232  ;
  assign n20051 = n6706 & n20050 ;
  assign n20052 = ~n17419 & n20051 ;
  assign n20053 = ~n9948 & ~n20052 ;
  assign n20054 = n15926 & n20053 ;
  assign n20055 = n20049 & n20054 ;
  assign n20056 = ~\pi0132  & ~\pi0135  ;
  assign n20057 = n17436 & n20056 ;
  assign n20058 = n18904 & n20057 ;
  assign n20059 = \pi0134  & ~n20058 ;
  assign n20060 = n9948 & n20059 ;
  assign n20061 = \pi0192  & ~\pi0299  ;
  assign n20062 = \pi0171  & \pi0299  ;
  assign n20063 = ~n20061 & ~n20062 ;
  assign n20064 = n8640 & ~n20063 ;
  assign n20065 = n17507 & ~n20064 ;
  assign n20066 = n9948 & n17720 ;
  assign n20067 = n20065 & n20066 ;
  assign n20068 = ~n20060 & ~n20067 ;
  assign n20069 = ~n17419 & n19978 ;
  assign n20070 = ~n20064 & n20069 ;
  assign n20071 = \pi0232  & n2327 ;
  assign n20072 = ~n20070 & n20071 ;
  assign n20073 = n18192 & n19439 ;
  assign n20074 = n2327 & ~n20070 ;
  assign n20075 = ~n11040 & n20074 ;
  assign n20076 = ~n20073 & n20075 ;
  assign n20077 = ~n18941 & ~n20065 ;
  assign n20078 = ~n2327 & n20077 ;
  assign n20079 = n19778 & ~n20078 ;
  assign n20080 = ~n20076 & n20079 ;
  assign n20081 = ~n20072 & n20080 ;
  assign n20082 = ~\pi0171  & n19473 ;
  assign n20083 = \pi0164  & \pi0216  ;
  assign n20084 = n6936 & n20083 ;
  assign n20085 = ~n17627 & n20084 ;
  assign n20086 = ~n20082 & n20085 ;
  assign n20087 = ~n19470 & n20086 ;
  assign n20088 = ~\pi0171  & n6936 ;
  assign n20089 = n20083 & n20088 ;
  assign n20090 = ~n19473 & n20089 ;
  assign n20091 = \pi0171  & n6706 ;
  assign n20092 = ~n7597 & ~n20091 ;
  assign n20093 = n17507 & n20092 ;
  assign n20094 = \pi0299  & ~n20093 ;
  assign n20095 = ~\pi0164  & \pi0216  ;
  assign n20096 = n6936 & n20095 ;
  assign n20097 = n20094 & ~n20096 ;
  assign n20098 = ~\pi0051  & ~n20091 ;
  assign n20099 = ~n17953 & n20098 ;
  assign n20100 = n1281 & n20091 ;
  assign n20101 = n1260 & n20100 ;
  assign n20102 = n20094 & ~n20101 ;
  assign n20103 = ~n20099 & n20102 ;
  assign n20104 = ~n20097 & ~n20103 ;
  assign n20105 = ~n20090 & ~n20104 ;
  assign n20106 = ~n20087 & n20105 ;
  assign n20107 = \pi0186  & ~\pi0287  ;
  assign n20108 = n6706 & n20107 ;
  assign n20109 = ~\pi0051  & ~n20108 ;
  assign n20110 = ~n18273 & n20109 ;
  assign n20111 = ~n18267 & n20110 ;
  assign n20112 = n20061 & ~n20111 ;
  assign n20113 = ~n20106 & ~n20112 ;
  assign n20114 = ~\pi0192  & ~\pi0299  ;
  assign n20115 = n19453 & n20114 ;
  assign n20116 = \pi0186  & n20114 ;
  assign n20117 = n18250 & n20116 ;
  assign n20118 = ~n20115 & ~n20117 ;
  assign n20119 = n20080 & n20118 ;
  assign n20120 = n20113 & n20119 ;
  assign n20121 = ~n20081 & ~n20120 ;
  assign n20122 = n20068 & n20121 ;
  assign n20123 = ~n20055 & n20122 ;
  assign n20124 = n17660 & ~n20078 ;
  assign n20125 = ~\pi0051  & ~n19543 ;
  assign n20126 = ~\pi0051  & n18496 ;
  assign n20127 = ~n17672 & n20126 ;
  assign n20128 = ~n20125 & ~n20127 ;
  assign n20129 = n20114 & n20128 ;
  assign n20130 = \pi0186  & ~n20061 ;
  assign n20131 = \pi0186  & n19568 ;
  assign n20132 = ~n19564 & n20131 ;
  assign n20133 = n19560 & n20132 ;
  assign n20134 = ~n20130 & ~n20133 ;
  assign n20135 = ~n20129 & ~n20134 ;
  assign n20136 = ~n8701 & ~n18941 ;
  assign n20137 = \pi0039  & \pi0186  ;
  assign n20138 = ~n20114 & ~n20137 ;
  assign n20139 = ~n20136 & n20138 ;
  assign n20140 = ~\pi0051  & ~n20137 ;
  assign n20141 = ~n20136 & n20140 ;
  assign n20142 = ~n18526 & n20141 ;
  assign n20143 = ~n20139 & ~n20142 ;
  assign n20144 = n19560 & ~n20143 ;
  assign n20145 = ~n20061 & n20138 ;
  assign n20146 = ~n20061 & n20140 ;
  assign n20147 = ~n18526 & n20146 ;
  assign n20148 = ~n20145 & ~n20147 ;
  assign n20149 = \pi0232  & n20148 ;
  assign n20150 = ~n20144 & n20149 ;
  assign n20151 = ~n20135 & n20150 ;
  assign n20152 = ~\pi0051  & ~\pi0171  ;
  assign n20153 = ~n17672 & n20152 ;
  assign n20154 = \pi0171  & ~n18499 ;
  assign n20155 = ~n17421 & n20154 ;
  assign n20156 = ~n19561 & n20155 ;
  assign n20157 = ~n20153 & ~n20156 ;
  assign n20158 = n20083 & n20157 ;
  assign n20159 = ~\pi0216  & ~n20091 ;
  assign n20160 = ~n17945 & n20159 ;
  assign n20161 = ~n17419 & n20091 ;
  assign n20162 = ~\pi0051  & ~n20161 ;
  assign n20163 = n6936 & ~n20095 ;
  assign n20164 = ~n20162 & ~n20163 ;
  assign n20165 = ~\pi0216  & n20091 ;
  assign n20166 = ~n17953 & n20165 ;
  assign n20167 = ~n20164 & ~n20166 ;
  assign n20168 = ~n20160 & n20167 ;
  assign n20169 = ~n20158 & n20168 ;
  assign n20170 = n17987 & ~n20161 ;
  assign n20171 = \pi0299  & ~n20170 ;
  assign n20172 = \pi0232  & n20171 ;
  assign n20173 = ~n20169 & n20172 ;
  assign n20174 = ~n19555 & ~n20173 ;
  assign n20175 = ~n20151 & n20174 ;
  assign n20176 = ~n17462 & n19584 ;
  assign n20177 = \pi0232  & ~n20063 ;
  assign n20178 = ~n18767 & n20177 ;
  assign n20179 = ~n20176 & n20178 ;
  assign n20180 = ~\pi0039  & n20177 ;
  assign n20181 = ~n19594 & ~n20180 ;
  assign n20182 = ~n20179 & ~n20181 ;
  assign n20183 = n2327 & ~n20182 ;
  assign n20184 = ~n20175 & n20183 ;
  assign n20185 = n20124 & ~n20184 ;
  assign n20186 = n17720 & ~n20077 ;
  assign n20187 = n20059 & ~n20186 ;
  assign n20188 = ~n20055 & n20187 ;
  assign n20189 = ~n20185 & n20188 ;
  assign n20190 = ~n20123 & ~n20189 ;
  assign n20191 = \pi0170  & n6706 ;
  assign n20192 = n10276 & n20191 ;
  assign n20193 = n19444 & ~n20192 ;
  assign n20194 = ~\pi0194  & ~n20193 ;
  assign n20195 = \pi0170  & \pi0232  ;
  assign n20196 = n6706 & n20195 ;
  assign n20197 = ~n10195 & ~n20196 ;
  assign n20198 = n19444 & n20197 ;
  assign n20199 = \pi0194  & ~n20198 ;
  assign n20200 = ~n20194 & ~n20199 ;
  assign n20201 = n19442 & ~n20200 ;
  assign n20202 = n19453 & n20194 ;
  assign n20203 = \pi0185  & ~\pi0194  ;
  assign n20204 = ~n20193 & n20203 ;
  assign n20205 = n18250 & n20204 ;
  assign n20206 = ~n20202 & ~n20205 ;
  assign n20207 = ~\pi0299  & ~n20206 ;
  assign n20208 = ~n20201 & ~n20207 ;
  assign n20209 = \pi0185  & ~\pi0287  ;
  assign n20210 = n6706 & n20209 ;
  assign n20211 = ~\pi0051  & ~n20210 ;
  assign n20212 = ~n18273 & n20211 ;
  assign n20213 = ~n18267 & n20212 ;
  assign n20214 = \pi0194  & ~\pi0299  ;
  assign n20215 = ~n20198 & n20214 ;
  assign n20216 = ~n20213 & n20215 ;
  assign n20217 = ~\pi0051  & ~\pi0170  ;
  assign n20218 = n17419 & n20217 ;
  assign n20219 = ~n18205 & n20218 ;
  assign n20220 = \pi0051  & ~\pi0170  ;
  assign n20221 = n7597 & ~n20220 ;
  assign n20222 = ~n17627 & n20221 ;
  assign n20223 = ~n20219 & n20222 ;
  assign n20224 = ~n19470 & n20223 ;
  assign n20225 = n17420 & ~n18205 ;
  assign n20226 = ~\pi0170  & ~n20220 ;
  assign n20227 = n7597 & n20226 ;
  assign n20228 = ~n20225 & n20227 ;
  assign n20229 = \pi0150  & \pi0299  ;
  assign n20230 = ~n7597 & ~n20191 ;
  assign n20231 = n17507 & n20230 ;
  assign n20232 = ~n20200 & ~n20231 ;
  assign n20233 = n20229 & n20232 ;
  assign n20234 = ~n20228 & n20233 ;
  assign n20235 = ~n20224 & n20234 ;
  assign n20236 = \pi0051  & ~n20191 ;
  assign n20237 = n17420 & ~n20191 ;
  assign n20238 = ~n17636 & n20237 ;
  assign n20239 = ~n20236 & ~n20238 ;
  assign n20240 = n7597 & ~n20191 ;
  assign n20241 = n1281 & n7597 ;
  assign n20242 = n1260 & n20241 ;
  assign n20243 = ~n20240 & ~n20242 ;
  assign n20244 = n20239 & ~n20243 ;
  assign n20245 = n19240 & n20232 ;
  assign n20246 = ~n20244 & n20245 ;
  assign n20247 = ~n20235 & ~n20246 ;
  assign n20248 = ~n20216 & n20247 ;
  assign n20249 = n20208 & n20248 ;
  assign n20250 = ~\pi0232  & ~n20201 ;
  assign n20251 = \pi0135  & ~n20046 ;
  assign n20252 = \pi0134  & ~\pi0135  ;
  assign n20253 = n20046 & n20252 ;
  assign n20254 = ~n20251 & ~n20253 ;
  assign n20255 = n17507 & ~n20192 ;
  assign n20256 = \pi0194  & n10195 ;
  assign n20257 = n17720 & ~n20256 ;
  assign n20258 = n20255 & n20257 ;
  assign n20259 = n20254 & ~n20258 ;
  assign n20260 = ~\pi0100  & n20259 ;
  assign n20261 = ~n20250 & n20260 ;
  assign n20262 = ~n20249 & n20261 ;
  assign n20263 = n20255 & ~n20256 ;
  assign n20264 = \pi0051  & \pi0100  ;
  assign n20265 = \pi0100  & n6706 ;
  assign n20266 = ~n17419 & n20265 ;
  assign n20267 = ~n20264 & ~n20266 ;
  assign n20268 = ~n20263 & ~n20267 ;
  assign n20269 = n18041 & ~n20268 ;
  assign n20270 = n20259 & ~n20269 ;
  assign n20271 = n9948 & ~n20270 ;
  assign n20272 = ~n20262 & n20271 ;
  assign n20273 = n17419 & ~n20252 ;
  assign n20274 = n20046 & n20273 ;
  assign n20275 = ~n20046 & n20047 ;
  assign n20276 = ~n20274 & ~n20275 ;
  assign n20277 = ~n9948 & n15926 ;
  assign n20278 = ~n17419 & n20196 ;
  assign n20279 = n20277 & ~n20278 ;
  assign n20280 = n20276 & n20279 ;
  assign n20281 = ~n20272 & ~n20280 ;
  assign n20282 = n17660 & n20267 ;
  assign n20283 = n17660 & ~n20256 ;
  assign n20284 = n20255 & n20283 ;
  assign n20285 = ~n20282 & ~n20284 ;
  assign n20286 = \pi0100  & ~n20285 ;
  assign n20287 = ~n18941 & ~n20255 ;
  assign n20288 = \pi0038  & ~n20287 ;
  assign n20289 = ~\pi0194  & ~n20288 ;
  assign n20290 = n17507 & n20197 ;
  assign n20291 = ~n18941 & ~n20290 ;
  assign n20292 = \pi0038  & \pi0194  ;
  assign n20293 = n20291 & n20292 ;
  assign n20294 = ~n20289 & ~n20293 ;
  assign n20295 = \pi0170  & n18767 ;
  assign n20296 = \pi0170  & n19584 ;
  assign n20297 = ~n17462 & n20296 ;
  assign n20298 = ~n20295 & ~n20297 ;
  assign n20299 = ~n17746 & n20217 ;
  assign n20300 = ~n17462 & n20299 ;
  assign n20301 = n10276 & ~n20300 ;
  assign n20302 = n20298 & n20301 ;
  assign n20303 = ~\pi0299  & ~n17809 ;
  assign n20304 = ~n19595 & ~n20303 ;
  assign n20305 = ~n20302 & n20304 ;
  assign n20306 = \pi0170  & ~n18499 ;
  assign n20307 = ~n17421 & n20306 ;
  assign n20308 = ~n19561 & n20307 ;
  assign n20309 = \pi0216  & ~n20308 ;
  assign n20310 = ~n17672 & n20217 ;
  assign n20311 = ~n17419 & n20191 ;
  assign n20312 = n17987 & ~n20311 ;
  assign n20313 = n20229 & ~n20312 ;
  assign n20314 = ~n20310 & n20313 ;
  assign n20315 = n20309 & n20314 ;
  assign n20316 = n17953 & n20191 ;
  assign n20317 = ~\pi0051  & ~n20191 ;
  assign n20318 = ~n17944 & n20317 ;
  assign n20319 = ~n20316 & ~n20318 ;
  assign n20320 = n8684 & ~n20319 ;
  assign n20321 = ~n7597 & n20229 ;
  assign n20322 = ~n20312 & n20321 ;
  assign n20323 = ~n20320 & n20322 ;
  assign n20324 = ~n20315 & ~n20323 ;
  assign n20325 = ~\pi0051  & ~n8684 ;
  assign n20326 = ~n20311 & n20325 ;
  assign n20327 = n19240 & ~n20326 ;
  assign n20328 = ~n20320 & n20327 ;
  assign n20329 = \pi0185  & ~n20128 ;
  assign n20330 = ~\pi0051  & ~\pi0185  ;
  assign n20331 = ~n18526 & n20330 ;
  assign n20332 = ~\pi0299  & ~n20331 ;
  assign n20333 = ~n20329 & n20332 ;
  assign n20334 = ~n20328 & ~n20333 ;
  assign n20335 = n20324 & n20334 ;
  assign n20336 = \pi0232  & ~n20335 ;
  assign n20337 = ~n19555 & ~n20336 ;
  assign n20338 = ~n20305 & ~n20337 ;
  assign n20339 = ~\pi0038  & ~n20293 ;
  assign n20340 = ~n20338 & n20339 ;
  assign n20341 = ~n20294 & ~n20340 ;
  assign n20342 = \pi0038  & ~n20291 ;
  assign n20343 = \pi0194  & ~n20342 ;
  assign n20344 = n10118 & ~n18767 ;
  assign n20345 = ~n20176 & n20344 ;
  assign n20346 = ~n19595 & ~n20345 ;
  assign n20347 = ~n20302 & n20346 ;
  assign n20348 = ~\pi0232  & ~n19555 ;
  assign n20349 = n20324 & ~n20328 ;
  assign n20350 = \pi0185  & n19568 ;
  assign n20351 = ~n19564 & n20350 ;
  assign n20352 = n19560 & n20351 ;
  assign n20353 = ~\pi0185  & n8701 ;
  assign n20354 = ~n17504 & n20330 ;
  assign n20355 = ~n20353 & ~n20354 ;
  assign n20356 = ~n19557 & ~n20355 ;
  assign n20357 = ~n19559 & n20356 ;
  assign n20358 = ~\pi0299  & ~n20357 ;
  assign n20359 = ~n20352 & n20358 ;
  assign n20360 = ~n19555 & ~n20359 ;
  assign n20361 = n20349 & n20360 ;
  assign n20362 = ~n20348 & ~n20361 ;
  assign n20363 = ~n20347 & n20362 ;
  assign n20364 = n20343 & n20363 ;
  assign n20365 = ~n20285 & ~n20364 ;
  assign n20366 = ~n20341 & n20365 ;
  assign n20367 = ~n20286 & ~n20366 ;
  assign n20368 = n17720 & n18941 ;
  assign n20369 = ~n20258 & ~n20368 ;
  assign n20370 = ~n20254 & n20369 ;
  assign n20371 = ~n20280 & n20370 ;
  assign n20372 = n20367 & n20371 ;
  assign n20373 = ~n20281 & ~n20372 ;
  assign n20374 = ~n2327 & ~n17419 ;
  assign n20375 = n11170 & n20374 ;
  assign n20376 = \pi0051  & ~n2327 ;
  assign n20377 = n17660 & ~n20376 ;
  assign n20378 = ~n20375 & n20377 ;
  assign n20379 = n2327 & ~n11040 ;
  assign n20380 = ~n19554 & n20379 ;
  assign n20381 = ~n20071 & ~n20380 ;
  assign n20382 = n6706 & n8684 ;
  assign n20383 = ~n17953 & n20382 ;
  assign n20384 = ~n6706 & n8684 ;
  assign n20385 = ~n17945 & n20384 ;
  assign n20386 = ~n20383 & ~n20385 ;
  assign n20387 = ~\pi0163  & \pi0216  ;
  assign n20388 = n6936 & ~n20387 ;
  assign n20389 = \pi0148  & n20388 ;
  assign n20390 = ~\pi0051  & \pi0148  ;
  assign n20391 = ~n17504 & n20390 ;
  assign n20392 = ~n20389 & ~n20391 ;
  assign n20393 = \pi0163  & n6936 ;
  assign n20394 = ~n19563 & n20393 ;
  assign n20395 = ~n20392 & ~n20394 ;
  assign n20396 = n20386 & n20395 ;
  assign n20397 = ~\pi0051  & ~\pi0148  ;
  assign n20398 = \pi0163  & ~\pi0287  ;
  assign n20399 = n6706 & n20398 ;
  assign n20400 = \pi0216  & ~n20399 ;
  assign n20401 = n6936 & ~n20400 ;
  assign n20402 = n17943 & n20401 ;
  assign n20403 = n1358 & n20402 ;
  assign n20404 = n20397 & ~n20403 ;
  assign n20405 = \pi0299  & ~n20404 ;
  assign n20406 = ~n20396 & n20405 ;
  assign n20407 = \pi0184  & ~n20128 ;
  assign n20408 = ~\pi0141  & ~\pi0299  ;
  assign n20409 = ~\pi0051  & ~\pi0184  ;
  assign n20410 = ~n18526 & n20409 ;
  assign n20411 = n20408 & ~n20410 ;
  assign n20412 = ~n20407 & n20411 ;
  assign n20413 = ~n20406 & ~n20412 ;
  assign n20414 = \pi0184  & n19568 ;
  assign n20415 = ~n19564 & n20414 ;
  assign n20416 = n19560 & n20415 ;
  assign n20417 = ~\pi0184  & n8701 ;
  assign n20418 = ~n17504 & n20409 ;
  assign n20419 = ~n20417 & ~n20418 ;
  assign n20420 = ~n19557 & ~n20419 ;
  assign n20421 = ~n19559 & n20420 ;
  assign n20422 = n11167 & ~n20421 ;
  assign n20423 = ~n20416 & n20422 ;
  assign n20424 = ~n20380 & ~n20423 ;
  assign n20425 = n20413 & n20424 ;
  assign n20426 = ~n20381 & ~n20425 ;
  assign n20427 = n20378 & ~n20426 ;
  assign n20428 = ~n11169 & n18767 ;
  assign n20429 = ~n11169 & n19584 ;
  assign n20430 = ~n17462 & n20429 ;
  assign n20431 = ~n20428 & ~n20430 ;
  assign n20432 = ~\pi0051  & n11169 ;
  assign n20433 = ~n17746 & n20432 ;
  assign n20434 = ~n17462 & n20433 ;
  assign n20435 = \pi0232  & ~n20434 ;
  assign n20436 = n20431 & n20435 ;
  assign n20437 = ~n19595 & n20378 ;
  assign n20438 = ~n20436 & n20437 ;
  assign n20439 = ~n11136 & ~n17419 ;
  assign n20440 = n20277 & n20439 ;
  assign n20441 = n11170 & ~n17419 ;
  assign n20442 = ~n13441 & n15926 ;
  assign n20443 = ~n20441 & n20442 ;
  assign n20444 = ~n20440 & ~n20443 ;
  assign n20445 = ~\pi0130  & ~\pi0132  ;
  assign n20446 = ~n17435 & n20445 ;
  assign n20447 = n18904 & n20446 ;
  assign n20448 = ~\pi0136  & n20447 ;
  assign n20449 = n18904 & n20445 ;
  assign n20450 = \pi0136  & ~n20449 ;
  assign n20451 = ~n20448 & ~n20450 ;
  assign n20452 = ~n9948 & n17444 ;
  assign n20453 = ~n20451 & ~n20452 ;
  assign n20454 = n20444 & n20453 ;
  assign n20455 = ~n20438 & n20454 ;
  assign n20456 = ~n20427 & n20455 ;
  assign n20457 = ~n20451 & n20452 ;
  assign n20458 = ~n20440 & ~n20457 ;
  assign n20459 = ~n9948 & n20458 ;
  assign n20460 = \pi0184  & ~\pi0287  ;
  assign n20461 = n6706 & n20460 ;
  assign n20462 = ~\pi0051  & ~n20461 ;
  assign n20463 = ~n18273 & n20462 ;
  assign n20464 = ~n18267 & n20463 ;
  assign n20465 = n11167 & ~n20464 ;
  assign n20466 = ~\pi0051  & ~n20399 ;
  assign n20467 = n18180 & n20466 ;
  assign n20468 = n17751 & n20467 ;
  assign n20469 = \pi0148  & ~n20399 ;
  assign n20470 = ~n17419 & n20397 ;
  assign n20471 = ~n20469 & ~n20470 ;
  assign n20472 = ~n20468 & n20471 ;
  assign n20473 = n7597 & ~n20472 ;
  assign n20474 = ~n19470 & n20473 ;
  assign n20475 = ~n6706 & ~n7597 ;
  assign n20476 = n17507 & n20475 ;
  assign n20477 = \pi0148  & ~n20476 ;
  assign n20478 = ~n20472 & ~n20477 ;
  assign n20479 = \pi0299  & ~n20478 ;
  assign n20480 = ~n20474 & n20479 ;
  assign n20481 = \pi0184  & n20408 ;
  assign n20482 = n18250 & n20481 ;
  assign n20483 = n19453 & n20408 ;
  assign n20484 = ~n20482 & ~n20483 ;
  assign n20485 = ~n20480 & n20484 ;
  assign n20486 = ~n20465 & n20485 ;
  assign n20487 = ~n12967 & ~n17419 ;
  assign n20488 = ~\pi0051  & n20487 ;
  assign n20489 = ~n11170 & n20488 ;
  assign n20490 = \pi0232  & ~n20489 ;
  assign n20491 = ~n20486 & n20490 ;
  assign n20492 = n2327 & n11040 ;
  assign n20493 = n2327 & n19439 ;
  assign n20494 = n18192 & n20493 ;
  assign n20495 = ~n20492 & ~n20494 ;
  assign n20496 = ~n20489 & n20495 ;
  assign n20497 = n17660 & ~n20496 ;
  assign n20498 = ~n20491 & n20497 ;
  assign n20499 = ~n11170 & n17720 ;
  assign n20500 = n17507 & n20499 ;
  assign n20501 = n20451 & ~n20500 ;
  assign n20502 = n20458 & n20501 ;
  assign n20503 = ~n20498 & n20502 ;
  assign n20504 = ~n20459 & ~n20503 ;
  assign n20505 = ~n20456 & n20504 ;
  assign n20506 = ~\pi0038  & \pi0287  ;
  assign n20507 = n1289 & n20506 ;
  assign n20508 = n1287 & n20507 ;
  assign n20509 = n1281 & n20508 ;
  assign n20510 = n1260 & n20509 ;
  assign n20511 = n1800 & n6683 ;
  assign n20512 = n11984 & n20511 ;
  assign n20513 = n2166 & n6706 ;
  assign n20514 = n2265 & n20513 ;
  assign n20515 = ~\pi0057  & ~\pi0299  ;
  assign n20516 = n6848 & n20515 ;
  assign n20517 = n20514 & n20516 ;
  assign n20518 = ~n20512 & ~n20517 ;
  assign n20519 = n11040 & ~n20518 ;
  assign n20520 = ~n20510 & n20519 ;
  assign n20521 = ~\pi0039  & \pi0137  ;
  assign n20522 = ~\pi0210  & n1800 ;
  assign n20523 = n11984 & n20522 ;
  assign n20524 = ~n9948 & n20523 ;
  assign n20525 = n11040 & n20524 ;
  assign n20526 = ~n20521 & ~n20525 ;
  assign n20527 = ~n20520 & n20526 ;
  assign n20528 = n10173 & n10176 ;
  assign n20529 = n8601 & n10156 ;
  assign n20530 = n2511 & n20529 ;
  assign n20531 = ~n20528 & n20530 ;
  assign n20532 = ~n8500 & ~n20531 ;
  assign n20533 = \pi0092  & ~n20532 ;
  assign n20534 = n10182 & ~n10259 ;
  assign n20535 = n10182 & ~n14078 ;
  assign n20536 = ~n10275 & ~n20535 ;
  assign n20537 = ~n20534 & n20536 ;
  assign n20538 = \pi0148  & n10275 ;
  assign n20539 = \pi0148  & ~n10252 ;
  assign n20540 = ~n10254 & n20539 ;
  assign n20541 = ~n20538 & ~n20540 ;
  assign n20542 = ~n20537 & ~n20541 ;
  assign n20543 = ~n10280 & ~n11168 ;
  assign n20544 = n7597 & n10182 ;
  assign n20545 = ~n14078 & n20544 ;
  assign n20546 = ~n10259 & n20544 ;
  assign n20547 = ~n20545 & ~n20546 ;
  assign n20548 = n10219 & n17197 ;
  assign n20549 = ~n10252 & ~n11168 ;
  assign n20550 = ~n20548 & n20549 ;
  assign n20551 = ~n20547 & n20550 ;
  assign n20552 = ~n20543 & ~n20551 ;
  assign n20553 = ~n20542 & n20552 ;
  assign n20554 = \pi0141  & ~n10284 ;
  assign n20555 = n6955 & n10182 ;
  assign n20556 = n10216 & n10282 ;
  assign n20557 = n10173 & n20556 ;
  assign n20558 = n20555 & ~n20557 ;
  assign n20559 = ~n20534 & ~n20535 ;
  assign n20560 = n20558 & ~n20559 ;
  assign n20561 = ~n20554 & n20560 ;
  assign n20562 = n10238 & ~n20561 ;
  assign n20563 = ~n20553 & ~n20562 ;
  assign n20564 = n11040 & ~n20563 ;
  assign n20565 = n10238 & ~n20558 ;
  assign n20566 = ~\pi0232  & n20565 ;
  assign n20567 = n10238 & ~n20535 ;
  assign n20568 = ~\pi0232  & ~n20534 ;
  assign n20569 = n20567 & n20568 ;
  assign n20570 = ~n20566 & ~n20569 ;
  assign n20571 = ~n10252 & ~n20548 ;
  assign n20572 = ~n20547 & n20571 ;
  assign n20573 = ~n10275 & n13992 ;
  assign n20574 = ~n20572 & n20573 ;
  assign n20575 = n20570 & ~n20574 ;
  assign n20576 = \pi0039  & ~n20575 ;
  assign n20577 = n2327 & ~n20576 ;
  assign n20578 = ~n20564 & n20577 ;
  assign n20579 = ~\pi0087  & ~n20578 ;
  assign n20580 = n8368 & n11239 ;
  assign n20581 = ~\pi0039  & ~n20580 ;
  assign n20582 = n10735 & n13992 ;
  assign n20583 = ~\pi0087  & ~n20582 ;
  assign n20584 = n20581 & n20583 ;
  assign n20585 = ~n20579 & ~n20584 ;
  assign n20586 = ~n6706 & n11167 ;
  assign n20587 = ~n11239 & n20586 ;
  assign n20588 = n6706 & n11167 ;
  assign n20589 = ~n10366 & n20588 ;
  assign n20590 = ~\pi0198  & n20588 ;
  assign n20591 = ~n10375 & n20590 ;
  assign n20592 = ~n20589 & ~n20591 ;
  assign n20593 = ~n20587 & n20592 ;
  assign n20594 = ~n11239 & n20408 ;
  assign n20595 = \pi0232  & ~n20594 ;
  assign n20596 = n20593 & n20595 ;
  assign n20597 = \pi0148  & n6706 ;
  assign n20598 = ~n10366 & n20597 ;
  assign n20599 = ~\pi0210  & n20597 ;
  assign n20600 = ~n10375 & n20599 ;
  assign n20601 = ~n20598 & ~n20600 ;
  assign n20602 = \pi0299  & ~n20601 ;
  assign n20603 = \pi0299  & ~n20597 ;
  assign n20604 = ~n10735 & n20603 ;
  assign n20605 = ~n20602 & ~n20604 ;
  assign n20606 = ~n20579 & n20605 ;
  assign n20607 = n20596 & n20606 ;
  assign n20608 = ~n20585 & ~n20607 ;
  assign n20609 = n10182 & n16139 ;
  assign n20610 = ~n1286 & ~n20609 ;
  assign n20611 = ~n20532 & ~n20610 ;
  assign n20612 = ~n20608 & n20611 ;
  assign n20613 = ~n20533 & ~n20612 ;
  assign n20614 = ~\pi0055  & ~\pi0062  ;
  assign n20615 = ~\pi0056  & n20614 ;
  assign n20616 = n20613 & n20615 ;
  assign n20617 = \pi0055  & ~n10158 ;
  assign n20618 = \pi0055  & ~\pi0092  ;
  assign n20619 = n10175 & n20618 ;
  assign n20620 = n10174 & n20619 ;
  assign n20621 = n10173 & n20620 ;
  assign n20622 = ~n20617 & ~n20621 ;
  assign n20623 = n1292 & ~n20622 ;
  assign n20624 = \pi0138  & n2467 ;
  assign n20625 = ~n11149 & n20624 ;
  assign n20626 = ~n20623 & n20625 ;
  assign n20627 = ~n20616 & n20626 ;
  assign n20628 = ~\pi0118  & ~\pi0139  ;
  assign n20629 = n16758 & n20628 ;
  assign n20630 = ~n11170 & n13708 ;
  assign n20631 = n10937 & n20630 ;
  assign n20632 = n10319 & n20631 ;
  assign n20633 = ~\pi0039  & ~n20632 ;
  assign n20634 = ~\pi0138  & n13386 ;
  assign n20635 = ~n20633 & n20634 ;
  assign n20636 = ~\pi0039  & n20635 ;
  assign n20637 = n7597 & n13577 ;
  assign n20638 = n6921 & n20637 ;
  assign n20639 = \pi0299  & ~n20638 ;
  assign n20640 = n6955 & n13581 ;
  assign n20641 = n6921 & n20640 ;
  assign n20642 = ~\pi0232  & ~\pi0299  ;
  assign n20643 = ~n20408 & ~n20642 ;
  assign n20644 = ~n20641 & ~n20643 ;
  assign n20645 = ~n20639 & ~n20644 ;
  assign n20646 = n6714 & n6932 ;
  assign n20647 = n6955 & ~n11168 ;
  assign n20648 = ~n6706 & n6955 ;
  assign n20649 = ~n6713 & n20648 ;
  assign n20650 = ~n20647 & ~n20649 ;
  assign n20651 = n20646 & ~n20650 ;
  assign n20652 = n6921 & n20651 ;
  assign n20653 = ~n6706 & ~n11167 ;
  assign n20654 = ~n6713 & n20653 ;
  assign n20655 = ~n11169 & ~n20654 ;
  assign n20656 = \pi0232  & n20655 ;
  assign n20657 = ~n20652 & n20656 ;
  assign n20658 = n20635 & ~n20657 ;
  assign n20659 = n20645 & n20658 ;
  assign n20660 = ~n20636 & ~n20659 ;
  assign n20661 = ~n20629 & n20660 ;
  assign n20662 = ~n20627 & n20661 ;
  assign n20663 = ~\pi0138  & ~n11099 ;
  assign n20664 = n11150 & n20663 ;
  assign n20665 = ~n20623 & n20664 ;
  assign n20666 = ~n20616 & n20665 ;
  assign n20667 = n13386 & ~n20663 ;
  assign n20668 = ~n20633 & n20667 ;
  assign n20669 = ~\pi0039  & n20668 ;
  assign n20670 = ~n20657 & n20668 ;
  assign n20671 = n20645 & n20670 ;
  assign n20672 = ~n20669 & ~n20671 ;
  assign n20673 = n20629 & n20672 ;
  assign n20674 = ~n20666 & n20673 ;
  assign n20675 = ~n20662 & ~n20674 ;
  assign n20676 = \pi0087  & n20611 ;
  assign n20677 = ~n10240 & n20555 ;
  assign n20678 = ~n20557 & n20677 ;
  assign n20679 = ~n10283 & n20678 ;
  assign n20680 = ~n20559 & n20679 ;
  assign n20681 = n10148 & ~n10220 ;
  assign n20682 = \pi0232  & n20681 ;
  assign n20683 = ~n20680 & n20682 ;
  assign n20684 = n7597 & ~n10252 ;
  assign n20685 = ~n10254 & n20684 ;
  assign n20686 = ~n20559 & n20685 ;
  assign n20687 = ~\pi0169  & n10182 ;
  assign n20688 = n7597 & n20687 ;
  assign n20689 = ~n10259 & n20688 ;
  assign n20690 = n10277 & ~n20689 ;
  assign n20691 = ~n20686 & n20690 ;
  assign n20692 = ~n20683 & ~n20691 ;
  assign n20693 = ~\pi0191  & n20565 ;
  assign n20694 = ~\pi0191  & ~n20534 ;
  assign n20695 = n20567 & n20694 ;
  assign n20696 = ~n20693 & ~n20695 ;
  assign n20697 = n20692 & n20696 ;
  assign n20698 = ~\pi0038  & n20575 ;
  assign n20699 = n20697 & n20698 ;
  assign n20700 = ~n1288 & ~n20699 ;
  assign n20701 = ~\pi0100  & n20611 ;
  assign n20702 = ~n20700 & n20701 ;
  assign n20703 = ~n20676 & ~n20702 ;
  assign n20704 = ~n20584 & ~n20703 ;
  assign n20705 = ~\pi0198  & n6706 ;
  assign n20706 = ~n10375 & n20705 ;
  assign n20707 = ~n16379 & ~n20706 ;
  assign n20708 = n10148 & ~n20707 ;
  assign n20709 = ~n6706 & n10148 ;
  assign n20710 = ~n11239 & n20709 ;
  assign n20711 = ~n20708 & ~n20710 ;
  assign n20712 = ~n11239 & n19450 ;
  assign n20713 = \pi0232  & ~n20712 ;
  assign n20714 = n20711 & n20713 ;
  assign n20715 = ~n10366 & n19483 ;
  assign n20716 = ~\pi0210  & n19483 ;
  assign n20717 = ~n10375 & n20716 ;
  assign n20718 = ~n20715 & ~n20717 ;
  assign n20719 = \pi0299  & ~n20718 ;
  assign n20720 = \pi0299  & ~n19483 ;
  assign n20721 = ~n10735 & n20720 ;
  assign n20722 = ~n20719 & ~n20721 ;
  assign n20723 = ~n20703 & n20722 ;
  assign n20724 = n20714 & n20723 ;
  assign n20725 = ~n20704 & ~n20724 ;
  assign n20726 = ~\pi0055  & n1292 ;
  assign n20727 = \pi0092  & n2511 ;
  assign n20728 = n20529 & n20727 ;
  assign n20729 = ~n20528 & n20728 ;
  assign n20730 = n20726 & ~n20729 ;
  assign n20731 = n20725 & n20730 ;
  assign n20732 = \pi0139  & n2467 ;
  assign n20733 = ~n11149 & n20732 ;
  assign n20734 = ~n20623 & n20733 ;
  assign n20735 = ~n20731 & n20734 ;
  assign n20736 = ~\pi0118  & n16758 ;
  assign n20737 = n19450 & ~n20641 ;
  assign n20738 = n6955 & n20646 ;
  assign n20739 = n6921 & n20738 ;
  assign n20740 = n10148 & ~n20739 ;
  assign n20741 = ~n20737 & ~n20740 ;
  assign n20742 = n7597 & ~n10149 ;
  assign n20743 = ~n6706 & n7597 ;
  assign n20744 = ~n6713 & n20743 ;
  assign n20745 = ~n20742 & ~n20744 ;
  assign n20746 = n13577 & ~n20745 ;
  assign n20747 = n6921 & n20746 ;
  assign n20748 = \pi0299  & ~n20747 ;
  assign n20749 = \pi0232  & ~n20748 ;
  assign n20750 = n20741 & n20749 ;
  assign n20751 = n20641 & n20642 ;
  assign n20752 = n13992 & n20638 ;
  assign n20753 = ~n20751 & ~n20752 ;
  assign n20754 = \pi0039  & n20753 ;
  assign n20755 = ~n20750 & n20754 ;
  assign n20756 = n13708 & ~n19430 ;
  assign n20757 = n10937 & n20756 ;
  assign n20758 = n10319 & n20757 ;
  assign n20759 = ~\pi0039  & ~n20758 ;
  assign n20760 = ~\pi0139  & n13386 ;
  assign n20761 = ~n20759 & n20760 ;
  assign n20762 = ~n20755 & n20761 ;
  assign n20763 = ~n20736 & ~n20762 ;
  assign n20764 = ~n20735 & n20763 ;
  assign n20765 = ~\pi0138  & n11099 ;
  assign n20766 = ~\pi0139  & ~n20765 ;
  assign n20767 = n11150 & n20766 ;
  assign n20768 = ~n20623 & n20767 ;
  assign n20769 = ~n20731 & n20768 ;
  assign n20770 = n13386 & ~n20766 ;
  assign n20771 = ~n20759 & n20770 ;
  assign n20772 = ~n20755 & n20771 ;
  assign n20773 = n20736 & ~n20772 ;
  assign n20774 = ~n20769 & n20773 ;
  assign n20775 = ~n20764 & ~n20774 ;
  assign n20776 = ~\pi0626  & \pi1158  ;
  assign n20777 = \pi0626  & ~\pi1158  ;
  assign n20778 = ~n20776 & ~n20777 ;
  assign n20779 = ~\pi0140  & \pi0788  ;
  assign n20780 = ~n1689 & n20779 ;
  assign n20781 = ~n20778 & n20780 ;
  assign n20782 = ~\pi0140  & ~n1689 ;
  assign n20783 = \pi0621  & \pi1091  ;
  assign n20784 = \pi0603  & ~n20783 ;
  assign n20785 = ~\pi0761  & n1689 ;
  assign n20786 = n20784 & n20785 ;
  assign n20787 = ~n20782 & ~n20786 ;
  assign n20788 = \pi0608  & \pi1153  ;
  assign n20789 = \pi0778  & ~n20788 ;
  assign n20790 = ~\pi0608  & ~\pi1153  ;
  assign n20791 = n1689 & ~n20790 ;
  assign n20792 = n20789 & n20791 ;
  assign n20793 = \pi0609  & n1689 ;
  assign n20794 = ~n20792 & ~n20793 ;
  assign n20795 = ~n20787 & n20794 ;
  assign n20796 = \pi0785  & ~\pi1155  ;
  assign n20797 = ~n20795 & n20796 ;
  assign n20798 = ~\pi0609  & n1689 ;
  assign n20799 = ~n20792 & ~n20798 ;
  assign n20800 = ~n20787 & n20799 ;
  assign n20801 = \pi0785  & \pi1155  ;
  assign n20802 = ~n20800 & n20801 ;
  assign n20803 = ~n20797 & ~n20802 ;
  assign n20804 = ~\pi0785  & n20792 ;
  assign n20805 = ~\pi0785  & ~n20782 ;
  assign n20806 = ~n20786 & n20805 ;
  assign n20807 = ~n20804 & ~n20806 ;
  assign n20808 = \pi0781  & n1689 ;
  assign n20809 = ~\pi0618  & \pi1154  ;
  assign n20810 = \pi0618  & ~\pi1154  ;
  assign n20811 = ~n20809 & ~n20810 ;
  assign n20812 = n20808 & ~n20811 ;
  assign n20813 = n20807 & ~n20812 ;
  assign n20814 = ~\pi0789  & n20813 ;
  assign n20815 = n20803 & n20814 ;
  assign n20816 = \pi0788  & n20778 ;
  assign n20817 = n20815 & n20816 ;
  assign n20818 = n20803 & n20813 ;
  assign n20819 = ~\pi0789  & ~n20818 ;
  assign n20820 = ~\pi0619  & ~n20812 ;
  assign n20821 = n20807 & n20820 ;
  assign n20822 = n20803 & n20821 ;
  assign n20823 = ~\pi0140  & \pi0619  ;
  assign n20824 = ~n1689 & n20823 ;
  assign n20825 = ~\pi1159  & ~n20824 ;
  assign n20826 = ~n20822 & n20825 ;
  assign n20827 = ~n20819 & ~n20826 ;
  assign n20828 = ~\pi0619  & \pi1159  ;
  assign n20829 = ~n20782 & n20828 ;
  assign n20830 = \pi0619  & \pi1159  ;
  assign n20831 = ~n20829 & ~n20830 ;
  assign n20832 = n20813 & ~n20829 ;
  assign n20833 = n20803 & n20832 ;
  assign n20834 = ~n20831 & ~n20833 ;
  assign n20835 = n20816 & ~n20834 ;
  assign n20836 = n20827 & n20835 ;
  assign n20837 = ~n20817 & ~n20836 ;
  assign n20838 = ~n20781 & n20837 ;
  assign n20839 = ~\pi0788  & n20815 ;
  assign n20840 = ~\pi0788  & ~n20834 ;
  assign n20841 = n20827 & n20840 ;
  assign n20842 = ~n20839 & ~n20841 ;
  assign n20843 = ~\pi0629  & \pi1156  ;
  assign n20844 = \pi0629  & ~\pi1156  ;
  assign n20845 = ~n20843 & ~n20844 ;
  assign n20846 = \pi0792  & ~n20845 ;
  assign n20847 = n20842 & ~n20846 ;
  assign n20848 = n20838 & n20847 ;
  assign n20849 = ~\pi0630  & \pi1157  ;
  assign n20850 = ~\pi0647  & n20849 ;
  assign n20851 = ~n20782 & n20850 ;
  assign n20852 = \pi0647  & n20849 ;
  assign n20853 = ~n20851 & ~n20852 ;
  assign n20854 = \pi0665  & \pi1091  ;
  assign n20855 = \pi0680  & ~n20854 ;
  assign n20856 = ~\pi0738  & n1689 ;
  assign n20857 = n20855 & n20856 ;
  assign n20858 = \pi0625  & ~\pi1153  ;
  assign n20859 = ~\pi0625  & \pi1153  ;
  assign n20860 = ~n20858 & ~n20859 ;
  assign n20861 = \pi0778  & ~n20860 ;
  assign n20862 = n20857 & ~n20861 ;
  assign n20863 = ~n20782 & ~n20862 ;
  assign n20864 = ~\pi0660  & \pi1155  ;
  assign n20865 = \pi0660  & ~\pi1155  ;
  assign n20866 = ~n20864 & ~n20865 ;
  assign n20867 = \pi0785  & n1689 ;
  assign n20868 = ~n20866 & n20867 ;
  assign n20869 = ~\pi0627  & ~\pi1154  ;
  assign n20870 = \pi0627  & \pi1154  ;
  assign n20871 = ~n20869 & ~n20870 ;
  assign n20872 = n20808 & n20871 ;
  assign n20873 = ~n20868 & ~n20872 ;
  assign n20874 = \pi0648  & ~\pi1159  ;
  assign n20875 = ~\pi0648  & \pi1159  ;
  assign n20876 = ~n20874 & ~n20875 ;
  assign n20877 = \pi0789  & n1689 ;
  assign n20878 = ~n20876 & n20877 ;
  assign n20879 = n20873 & ~n20878 ;
  assign n20880 = ~n20863 & n20879 ;
  assign n20881 = ~\pi0641  & \pi1158  ;
  assign n20882 = \pi0641  & ~\pi1158  ;
  assign n20883 = ~n20881 & ~n20882 ;
  assign n20884 = \pi0788  & n1689 ;
  assign n20885 = ~n20883 & n20884 ;
  assign n20886 = ~\pi0628  & \pi1156  ;
  assign n20887 = \pi0628  & ~\pi1156  ;
  assign n20888 = ~n20886 & ~n20887 ;
  assign n20889 = \pi0792  & n1689 ;
  assign n20890 = ~n20888 & n20889 ;
  assign n20891 = ~n20885 & ~n20890 ;
  assign n20892 = ~n20851 & n20891 ;
  assign n20893 = n20880 & n20892 ;
  assign n20894 = ~n20853 & ~n20893 ;
  assign n20895 = ~\pi0647  & n20891 ;
  assign n20896 = n20880 & n20895 ;
  assign n20897 = \pi0630  & ~\pi1157  ;
  assign n20898 = ~\pi0140  & \pi0647  ;
  assign n20899 = ~n1689 & n20898 ;
  assign n20900 = n20897 & ~n20899 ;
  assign n20901 = ~n20896 & n20900 ;
  assign n20902 = ~n20894 & ~n20901 ;
  assign n20903 = ~n20782 & n20846 ;
  assign n20904 = n20902 & ~n20903 ;
  assign n20905 = ~n20848 & n20904 ;
  assign n20906 = \pi0630  & ~\pi0647  ;
  assign n20907 = \pi1157  & n20906 ;
  assign n20908 = ~\pi0630  & \pi0647  ;
  assign n20909 = ~\pi1157  & n20908 ;
  assign n20910 = ~n20907 & ~n20909 ;
  assign n20911 = n20902 & n20910 ;
  assign n20912 = \pi0787  & ~n20911 ;
  assign n20913 = ~n20905 & n20912 ;
  assign n20914 = ~\pi0644  & ~n20913 ;
  assign n20915 = ~\pi0787  & n20891 ;
  assign n20916 = n20880 & n20915 ;
  assign n20917 = \pi0644  & n20916 ;
  assign n20918 = n20880 & n20891 ;
  assign n20919 = ~\pi0787  & ~n20918 ;
  assign n20920 = ~\pi1157  & ~n20899 ;
  assign n20921 = ~n20896 & n20920 ;
  assign n20922 = ~n20919 & ~n20921 ;
  assign n20923 = ~\pi0647  & \pi1157  ;
  assign n20924 = ~n20782 & n20923 ;
  assign n20925 = \pi0647  & \pi1157  ;
  assign n20926 = ~n20924 & ~n20925 ;
  assign n20927 = n20891 & ~n20924 ;
  assign n20928 = n20880 & n20927 ;
  assign n20929 = ~n20926 & ~n20928 ;
  assign n20930 = \pi0644  & ~n20929 ;
  assign n20931 = n20922 & n20930 ;
  assign n20932 = ~n20917 & ~n20931 ;
  assign n20933 = ~\pi0715  & n20932 ;
  assign n20934 = ~n20914 & n20933 ;
  assign n20935 = ~\pi0629  & \pi0792  ;
  assign n20936 = \pi0628  & n1689 ;
  assign n20937 = ~\pi1156  & ~n20936 ;
  assign n20938 = ~n20885 & n20937 ;
  assign n20939 = \pi0792  & n20938 ;
  assign n20940 = n20880 & n20939 ;
  assign n20941 = ~n20935 & ~n20940 ;
  assign n20942 = ~\pi0628  & n20842 ;
  assign n20943 = n20838 & n20942 ;
  assign n20944 = \pi0792  & \pi1156  ;
  assign n20945 = ~n20943 & n20944 ;
  assign n20946 = n20941 & ~n20945 ;
  assign n20947 = n20778 & ~n20883 ;
  assign n20948 = ~\pi0626  & \pi0641  ;
  assign n20949 = \pi0626  & ~\pi0641  ;
  assign n20950 = ~n20948 & ~n20949 ;
  assign n20951 = ~n20778 & ~n20950 ;
  assign n20952 = n20880 & n20951 ;
  assign n20953 = ~n20778 & n20782 ;
  assign n20954 = ~n20883 & n20953 ;
  assign n20955 = ~n20952 & ~n20954 ;
  assign n20956 = ~n20947 & n20955 ;
  assign n20957 = n20827 & ~n20834 ;
  assign n20958 = ~n20815 & n20955 ;
  assign n20959 = ~n20957 & n20958 ;
  assign n20960 = ~n20956 & ~n20959 ;
  assign n20961 = \pi0788  & n20960 ;
  assign n20962 = \pi0628  & ~n20961 ;
  assign n20963 = \pi0618  & n1689 ;
  assign n20964 = ~\pi1154  & ~n20963 ;
  assign n20965 = n20807 & n20964 ;
  assign n20966 = n20803 & n20965 ;
  assign n20967 = n20809 & ~n20868 ;
  assign n20968 = \pi0627  & ~n20967 ;
  assign n20969 = \pi0627  & ~n20782 ;
  assign n20970 = ~n20862 & n20969 ;
  assign n20971 = ~n20968 & ~n20970 ;
  assign n20972 = ~n20966 & ~n20971 ;
  assign n20973 = ~\pi0618  & n1689 ;
  assign n20974 = \pi1154  & ~n20973 ;
  assign n20975 = n20807 & n20974 ;
  assign n20976 = n20803 & n20975 ;
  assign n20977 = n20810 & ~n20868 ;
  assign n20978 = ~\pi0627  & ~n20977 ;
  assign n20979 = ~\pi0627  & ~n20782 ;
  assign n20980 = ~n20862 & n20979 ;
  assign n20981 = ~n20978 & ~n20980 ;
  assign n20982 = ~n20976 & ~n20981 ;
  assign n20983 = ~n20972 & ~n20982 ;
  assign n20984 = \pi0781  & n20983 ;
  assign n20985 = n20789 & ~n20790 ;
  assign n20986 = n20784 & ~n20985 ;
  assign n20987 = \pi0680  & ~\pi0738  ;
  assign n20988 = ~n20854 & n20987 ;
  assign n20989 = ~n20861 & n20988 ;
  assign n20990 = ~n20986 & n20989 ;
  assign n20991 = \pi0603  & ~\pi0761  ;
  assign n20992 = ~n20783 & n20991 ;
  assign n20993 = ~n20985 & n20992 ;
  assign n20994 = ~n20782 & ~n20993 ;
  assign n20995 = ~n20990 & n20994 ;
  assign n20996 = \pi0140  & ~n1689 ;
  assign n20997 = ~\pi0609  & ~n20996 ;
  assign n20998 = ~n20995 & n20997 ;
  assign n20999 = ~\pi0609  & ~\pi1155  ;
  assign n21000 = ~\pi1155  & ~n20782 ;
  assign n21001 = ~n20862 & n21000 ;
  assign n21002 = ~n20999 & ~n21001 ;
  assign n21003 = ~n20998 & ~n21002 ;
  assign n21004 = \pi1155  & ~n20800 ;
  assign n21005 = ~\pi0660  & ~n21004 ;
  assign n21006 = ~n21003 & n21005 ;
  assign n21007 = ~\pi0660  & \pi0785  ;
  assign n21008 = ~n20797 & ~n21007 ;
  assign n21009 = \pi0609  & ~n20996 ;
  assign n21010 = ~n20995 & n21009 ;
  assign n21011 = ~\pi0609  & ~n20863 ;
  assign n21012 = n20801 & ~n21011 ;
  assign n21013 = ~n21010 & n21012 ;
  assign n21014 = n21008 & ~n21013 ;
  assign n21015 = ~n21006 & ~n21014 ;
  assign n21016 = ~\pi0618  & ~\pi0627  ;
  assign n21017 = \pi0781  & ~\pi1154  ;
  assign n21018 = ~n21016 & n21017 ;
  assign n21019 = \pi0618  & \pi0627  ;
  assign n21020 = \pi0781  & \pi1154  ;
  assign n21021 = ~n21019 & n21020 ;
  assign n21022 = ~n21018 & ~n21021 ;
  assign n21023 = \pi0785  & n21022 ;
  assign n21024 = ~n20996 & n21022 ;
  assign n21025 = ~n20995 & n21024 ;
  assign n21026 = ~n21023 & ~n21025 ;
  assign n21027 = ~n21015 & ~n21026 ;
  assign n21028 = ~\pi0619  & \pi0648  ;
  assign n21029 = \pi0619  & ~\pi0648  ;
  assign n21030 = ~n21028 & ~n21029 ;
  assign n21031 = \pi0619  & ~\pi1159  ;
  assign n21032 = ~n20828 & ~n21031 ;
  assign n21033 = n21030 & n21032 ;
  assign n21034 = \pi0789  & ~n21033 ;
  assign n21035 = ~n21027 & ~n21034 ;
  assign n21036 = ~n20984 & n21035 ;
  assign n21037 = n20778 & n20950 ;
  assign n21038 = \pi0788  & ~n21037 ;
  assign n21039 = ~\pi0619  & n20875 ;
  assign n21040 = ~n20782 & n21039 ;
  assign n21041 = \pi0619  & n20875 ;
  assign n21042 = ~n21040 & ~n21041 ;
  assign n21043 = n20813 & ~n21040 ;
  assign n21044 = n20803 & n21043 ;
  assign n21045 = ~n21042 & ~n21044 ;
  assign n21046 = ~n20824 & n20874 ;
  assign n21047 = ~n20822 & n21046 ;
  assign n21048 = \pi1159  & ~n21028 ;
  assign n21049 = ~\pi1159  & ~n21029 ;
  assign n21050 = ~n21048 & ~n21049 ;
  assign n21051 = ~n20873 & n21050 ;
  assign n21052 = ~n20782 & n21050 ;
  assign n21053 = ~n20862 & n21052 ;
  assign n21054 = ~n21051 & ~n21053 ;
  assign n21055 = ~n21047 & n21054 ;
  assign n21056 = ~n21045 & n21055 ;
  assign n21057 = \pi0789  & ~n21056 ;
  assign n21058 = ~n21038 & ~n21057 ;
  assign n21059 = ~n21036 & n21058 ;
  assign n21060 = n20941 & ~n21059 ;
  assign n21061 = n20962 & n21060 ;
  assign n21062 = ~n20946 & ~n21061 ;
  assign n21063 = ~n20849 & ~n20897 ;
  assign n21064 = \pi0647  & ~\pi1157  ;
  assign n21065 = ~n20923 & ~n21064 ;
  assign n21066 = n21063 & n21065 ;
  assign n21067 = \pi0787  & ~n21066 ;
  assign n21068 = ~n21062 & ~n21067 ;
  assign n21069 = ~\pi0628  & ~n21059 ;
  assign n21070 = ~n20961 & n21069 ;
  assign n21071 = \pi0628  & n20842 ;
  assign n21072 = n20838 & n21071 ;
  assign n21073 = ~\pi1156  & ~n21072 ;
  assign n21074 = ~n21070 & n21073 ;
  assign n21075 = ~\pi0628  & n1689 ;
  assign n21076 = \pi1156  & ~n21075 ;
  assign n21077 = ~n20885 & n21076 ;
  assign n21078 = n20880 & n21077 ;
  assign n21079 = ~\pi0629  & ~n21078 ;
  assign n21080 = ~n21067 & n21079 ;
  assign n21081 = ~n21074 & n21080 ;
  assign n21082 = ~n21068 & ~n21081 ;
  assign n21083 = ~n20961 & ~n21059 ;
  assign n21084 = ~\pi0792  & ~n21083 ;
  assign n21085 = n20933 & ~n21084 ;
  assign n21086 = ~n21082 & n21085 ;
  assign n21087 = ~n20934 & ~n21086 ;
  assign n21088 = \pi0787  & ~n21063 ;
  assign n21089 = ~n20781 & ~n21088 ;
  assign n21090 = n20837 & n21089 ;
  assign n21091 = n20847 & n21090 ;
  assign n21092 = ~n20846 & ~n21088 ;
  assign n21093 = ~n20782 & ~n21092 ;
  assign n21094 = ~\pi0644  & ~n21093 ;
  assign n21095 = ~n21091 & n21094 ;
  assign n21096 = ~\pi0140  & \pi0644  ;
  assign n21097 = ~n1689 & n21096 ;
  assign n21098 = \pi0715  & ~n21097 ;
  assign n21099 = ~n21095 & n21098 ;
  assign n21100 = ~\pi1160  & ~n21099 ;
  assign n21101 = n21087 & n21100 ;
  assign n21102 = \pi0790  & n21101 ;
  assign n21103 = \pi0644  & ~n20913 ;
  assign n21104 = ~\pi0644  & n20916 ;
  assign n21105 = ~\pi0644  & ~n20929 ;
  assign n21106 = n20922 & n21105 ;
  assign n21107 = ~n21104 & ~n21106 ;
  assign n21108 = ~n21103 & n21107 ;
  assign n21109 = ~n21084 & n21107 ;
  assign n21110 = ~n21082 & n21109 ;
  assign n21111 = ~n21108 & ~n21110 ;
  assign n21112 = \pi0715  & ~n21111 ;
  assign n21113 = ~\pi0140  & ~\pi0644  ;
  assign n21114 = ~n1689 & n21113 ;
  assign n21115 = ~\pi0715  & ~n21114 ;
  assign n21116 = \pi1160  & ~n21115 ;
  assign n21117 = \pi0644  & ~n21093 ;
  assign n21118 = \pi1160  & n21117 ;
  assign n21119 = ~n21091 & n21118 ;
  assign n21120 = ~n21116 & ~n21119 ;
  assign n21121 = \pi0790  & ~n21120 ;
  assign n21122 = ~n21112 & n21121 ;
  assign n21123 = ~n21102 & ~n21122 ;
  assign n21124 = ~\pi0790  & ~n20913 ;
  assign n21125 = \pi0832  & ~n21124 ;
  assign n21126 = \pi0832  & ~n21084 ;
  assign n21127 = ~n21082 & n21126 ;
  assign n21128 = ~n21125 & ~n21127 ;
  assign n21129 = n21123 & ~n21128 ;
  assign n21130 = \pi0140  & ~\pi0832  ;
  assign n21131 = ~\pi0057  & ~\pi0832  ;
  assign n21132 = n6848 & n21131 ;
  assign n21133 = ~n21130 & ~n21132 ;
  assign n21134 = n1264 & n9012 ;
  assign n21135 = ~n2585 & n21134 ;
  assign n21136 = ~\pi0098  & ~\pi0102  ;
  assign n21137 = n13430 & n21136 ;
  assign n21138 = ~\pi0098  & \pi0102  ;
  assign n21139 = n1534 & n21138 ;
  assign n21140 = ~n21137 & ~n21139 ;
  assign n21141 = ~\pi0088  & n21140 ;
  assign n21142 = ~\pi0035  & ~\pi0252  ;
  assign n21143 = n1618 & n21142 ;
  assign n21144 = n10058 & n13028 ;
  assign n21145 = n10058 & n13030 ;
  assign n21146 = n1542 & n21145 ;
  assign n21147 = ~n21144 & ~n21146 ;
  assign n21148 = n21143 & ~n21147 ;
  assign n21149 = ~n21141 & n21148 ;
  assign n21150 = ~\pi0040  & ~n21149 ;
  assign n21151 = \pi1093  & ~n21150 ;
  assign n21152 = n1320 & n1326 ;
  assign n21153 = ~n1392 & n21152 ;
  assign n21154 = ~\pi0035  & ~n21153 ;
  assign n21155 = n1389 & n13028 ;
  assign n21156 = n1389 & n13030 ;
  assign n21157 = n1542 & n21156 ;
  assign n21158 = ~n21155 & ~n21157 ;
  assign n21159 = ~n21141 & ~n21158 ;
  assign n21160 = \pi0314  & n1568 ;
  assign n21161 = n11948 & n21160 ;
  assign n21162 = n1542 & n21161 ;
  assign n21163 = ~\pi0047  & ~n21162 ;
  assign n21164 = ~\pi0035  & n21163 ;
  assign n21165 = ~n21159 & n21164 ;
  assign n21166 = ~n21154 & ~n21165 ;
  assign n21167 = \pi0252  & ~n11908 ;
  assign n21168 = \pi1093  & n21167 ;
  assign n21169 = n21166 & n21168 ;
  assign n21170 = ~n21151 & ~n21169 ;
  assign n21171 = n21135 & ~n21170 ;
  assign n21172 = n1270 & n13028 ;
  assign n21173 = n1315 & n21172 ;
  assign n21174 = ~n21140 & n21173 ;
  assign n21175 = n21164 & ~n21174 ;
  assign n21176 = ~\pi0040  & ~n11908 ;
  assign n21177 = ~n21154 & n21176 ;
  assign n21178 = ~n21175 & n21177 ;
  assign n21179 = \pi0252  & ~n1621 ;
  assign n21180 = ~n21178 & n21179 ;
  assign n21181 = n1264 & ~n2585 ;
  assign n21182 = n2582 & n13028 ;
  assign n21183 = n10058 & n21182 ;
  assign n21184 = ~n21140 & n21183 ;
  assign n21185 = ~\pi0040  & ~n21184 ;
  assign n21186 = n21181 & ~n21185 ;
  assign n21187 = ~\pi0252  & ~n21186 ;
  assign n21188 = \pi1092  & n1264 ;
  assign n21189 = \pi1093  & ~n14707 ;
  assign n21190 = n21188 & n21189 ;
  assign n21191 = ~n21187 & n21190 ;
  assign n21192 = ~n21180 & n21191 ;
  assign n21193 = ~n1686 & ~n21192 ;
  assign n21194 = ~n21171 & n21193 ;
  assign n21195 = n6704 & n21188 ;
  assign n21196 = ~n21187 & n21195 ;
  assign n21197 = ~n21180 & n21196 ;
  assign n21198 = ~n8799 & ~n21197 ;
  assign n21199 = ~n21194 & ~n21198 ;
  assign n21200 = ~\pi1091  & n21192 ;
  assign n21201 = ~\pi1091  & n21135 ;
  assign n21202 = ~n21170 & n21201 ;
  assign n21203 = ~n21200 & ~n21202 ;
  assign n21204 = ~\pi0210  & n21203 ;
  assign n21205 = ~n21199 & n21204 ;
  assign n21206 = n1686 & ~n21198 ;
  assign n21207 = ~n2585 & ~n21150 ;
  assign n21208 = ~n2585 & n21167 ;
  assign n21209 = n21166 & n21208 ;
  assign n21210 = ~n21207 & ~n21209 ;
  assign n21211 = ~\pi0032  & n21210 ;
  assign n21212 = \pi0032  & ~n10909 ;
  assign n21213 = ~\pi0095  & \pi0824  ;
  assign n21214 = n6809 & n21213 ;
  assign n21215 = ~n21212 & n21214 ;
  assign n21216 = ~n21211 & n21215 ;
  assign n21217 = ~n14707 & n21188 ;
  assign n21218 = ~n21187 & n21217 ;
  assign n21219 = ~n21180 & n21218 ;
  assign n21220 = ~\pi0032  & n21187 ;
  assign n21221 = ~\pi0032  & n21179 ;
  assign n21222 = ~n21178 & n21221 ;
  assign n21223 = ~n21220 & ~n21222 ;
  assign n21224 = ~\pi0095  & \pi0829  ;
  assign n21225 = n13053 & n21224 ;
  assign n21226 = ~n21212 & n21225 ;
  assign n21227 = n21223 & n21226 ;
  assign n21228 = ~n21219 & ~n21227 ;
  assign n21229 = ~n21216 & n21228 ;
  assign n21230 = \pi1093  & ~n21198 ;
  assign n21231 = ~n21229 & n21230 ;
  assign n21232 = ~n21206 & ~n21231 ;
  assign n21233 = n8543 & n21219 ;
  assign n21234 = n8543 & n21215 ;
  assign n21235 = ~n21211 & n21234 ;
  assign n21236 = ~n21233 & ~n21235 ;
  assign n21237 = \pi0210  & n21236 ;
  assign n21238 = n21232 & n21237 ;
  assign n21239 = ~n21205 & ~n21238 ;
  assign n21240 = \pi0621  & ~n21198 ;
  assign n21241 = ~n21194 & n21240 ;
  assign n21242 = ~\pi0210  & \pi0603  ;
  assign n21243 = ~n21241 & n21242 ;
  assign n21244 = n1686 & n21240 ;
  assign n21245 = \pi1093  & n21240 ;
  assign n21246 = ~n21229 & n21245 ;
  assign n21247 = ~n21244 & ~n21246 ;
  assign n21248 = \pi0210  & \pi0603  ;
  assign n21249 = n21247 & n21248 ;
  assign n21250 = ~n21243 & ~n21249 ;
  assign n21251 = n21239 & n21250 ;
  assign n21252 = \pi0299  & ~n21251 ;
  assign n21253 = ~\pi0621  & ~n21198 ;
  assign n21254 = ~n21194 & n21253 ;
  assign n21255 = n21203 & ~n21254 ;
  assign n21256 = ~\pi0198  & ~\pi0603  ;
  assign n21257 = ~n21255 & n21256 ;
  assign n21258 = \pi0198  & ~\pi0603  ;
  assign n21259 = n1686 & n21253 ;
  assign n21260 = \pi1093  & n21253 ;
  assign n21261 = ~n21229 & n21260 ;
  assign n21262 = ~n21259 & ~n21261 ;
  assign n21263 = n21236 & n21262 ;
  assign n21264 = n21258 & ~n21263 ;
  assign n21265 = ~n21257 & ~n21264 ;
  assign n21266 = ~\pi0198  & ~n21241 ;
  assign n21267 = ~\pi0299  & n21266 ;
  assign n21268 = \pi0198  & ~\pi0299  ;
  assign n21269 = n21247 & n21268 ;
  assign n21270 = ~n21267 & ~n21269 ;
  assign n21271 = n21265 & ~n21270 ;
  assign n21272 = ~n21252 & ~n21271 ;
  assign n21273 = ~\pi0039  & ~\pi0761  ;
  assign n21274 = n21272 & n21273 ;
  assign n21275 = ~n2165 & ~n6761 ;
  assign n21276 = n6716 & ~n6717 ;
  assign n21277 = ~\pi0287  & ~n21276 ;
  assign n21278 = ~\pi0120  & n1689 ;
  assign n21279 = n21277 & n21278 ;
  assign n21280 = n1281 & n21279 ;
  assign n21281 = n1260 & n21280 ;
  assign n21282 = \pi0120  & n1689 ;
  assign n21283 = n1281 & n21282 ;
  assign n21284 = n1260 & n21283 ;
  assign n21285 = ~n21281 & ~n21284 ;
  assign n21286 = ~n6706 & ~n21285 ;
  assign n21287 = \pi1092  & \pi1093  ;
  assign n21288 = n1281 & n21287 ;
  assign n21289 = n1260 & n21288 ;
  assign n21290 = \pi0120  & ~n21289 ;
  assign n21291 = ~\pi1091  & ~n21290 ;
  assign n21292 = ~\pi0287  & ~n6716 ;
  assign n21293 = ~\pi0287  & \pi0835  ;
  assign n21294 = ~n11879 & n21293 ;
  assign n21295 = ~n21292 & ~n21294 ;
  assign n21296 = \pi1092  & ~n21295 ;
  assign n21297 = n1281 & n21296 ;
  assign n21298 = n1260 & n21297 ;
  assign n21299 = ~n13053 & ~n21298 ;
  assign n21300 = n1281 & n21277 ;
  assign n21301 = n1260 & n21300 ;
  assign n21302 = ~\pi0824  & ~n21301 ;
  assign n21303 = \pi1093  & ~n21302 ;
  assign n21304 = ~n21299 & n21303 ;
  assign n21305 = ~\pi0120  & ~n21304 ;
  assign n21306 = n21291 & ~n21305 ;
  assign n21307 = n6706 & n21306 ;
  assign n21308 = ~\pi0824  & ~\pi0829  ;
  assign n21309 = ~n21301 & n21308 ;
  assign n21310 = ~\pi0829  & ~n13053 ;
  assign n21311 = ~n21298 & n21310 ;
  assign n21312 = ~n21309 & ~n21311 ;
  assign n21313 = ~\pi0829  & \pi1093  ;
  assign n21314 = ~n1686 & n21313 ;
  assign n21315 = \pi1093  & ~n1686 ;
  assign n21316 = n21298 & n21315 ;
  assign n21317 = ~n21314 & ~n21316 ;
  assign n21318 = \pi1091  & ~n21317 ;
  assign n21319 = n21312 & n21318 ;
  assign n21320 = n1689 & n21277 ;
  assign n21321 = n1281 & n21320 ;
  assign n21322 = n1260 & n21321 ;
  assign n21323 = n16968 & n21322 ;
  assign n21324 = ~\pi0120  & ~n21323 ;
  assign n21325 = ~n21319 & n21324 ;
  assign n21326 = n6706 & ~n21290 ;
  assign n21327 = ~n21325 & n21326 ;
  assign n21328 = ~n21307 & ~n21327 ;
  assign n21329 = ~n21286 & n21328 ;
  assign n21330 = n6713 & ~n21329 ;
  assign n21331 = ~n6713 & n21306 ;
  assign n21332 = ~n6713 & ~n21290 ;
  assign n21333 = ~n21325 & n21332 ;
  assign n21334 = ~n21331 & ~n21333 ;
  assign n21335 = ~n21330 & n21334 ;
  assign n21336 = ~\pi0603  & ~n21286 ;
  assign n21337 = n21328 & n21336 ;
  assign n21338 = \pi0603  & ~n21286 ;
  assign n21339 = ~n21327 & n21338 ;
  assign n21340 = ~n20784 & ~n21339 ;
  assign n21341 = ~n21337 & n21340 ;
  assign n21342 = n20783 & ~n21290 ;
  assign n21343 = ~n21325 & n21342 ;
  assign n21344 = ~\pi0621  & ~n21290 ;
  assign n21345 = ~n21325 & n21344 ;
  assign n21346 = ~n21306 & ~n21345 ;
  assign n21347 = ~\pi0603  & ~n21346 ;
  assign n21348 = ~n21343 & ~n21347 ;
  assign n21349 = ~n21341 & n21348 ;
  assign n21350 = ~n21335 & ~n21349 ;
  assign n21351 = n21275 & n21350 ;
  assign n21352 = n6706 & n21285 ;
  assign n21353 = ~n6706 & ~n21291 ;
  assign n21354 = n17064 & ~n21304 ;
  assign n21355 = ~n21353 & ~n21354 ;
  assign n21356 = ~n21352 & n21355 ;
  assign n21357 = ~n21290 & ~n21352 ;
  assign n21358 = ~n21325 & n21357 ;
  assign n21359 = ~n21356 & ~n21358 ;
  assign n21360 = n20783 & ~n21285 ;
  assign n21361 = \pi0603  & n6706 ;
  assign n21362 = ~n21360 & n21361 ;
  assign n21363 = \pi0603  & ~n6706 ;
  assign n21364 = ~n21343 & n21363 ;
  assign n21365 = ~n21362 & ~n21364 ;
  assign n21366 = ~n21359 & n21365 ;
  assign n21367 = n6709 & ~n21366 ;
  assign n21368 = ~n2165 & n6761 ;
  assign n21369 = ~\pi0614  & ~\pi0642  ;
  assign n21370 = ~\pi0616  & n21369 ;
  assign n21371 = ~\pi0603  & n21285 ;
  assign n21372 = n21370 & ~n21371 ;
  assign n21373 = ~n21362 & n21372 ;
  assign n21374 = ~n21364 & n21373 ;
  assign n21375 = ~n20784 & ~n21370 ;
  assign n21376 = ~n21285 & n21375 ;
  assign n21377 = ~n6709 & ~n21376 ;
  assign n21378 = ~n21374 & n21377 ;
  assign n21379 = n21368 & ~n21378 ;
  assign n21380 = ~n21367 & n21379 ;
  assign n21381 = n6720 & n16927 ;
  assign n21382 = n6719 & n21381 ;
  assign n21383 = n1689 & ~n21382 ;
  assign n21384 = n1281 & n21383 ;
  assign n21385 = n1260 & n21384 ;
  assign n21386 = \pi0120  & n20783 ;
  assign n21387 = n21385 & n21386 ;
  assign n21388 = ~\pi0120  & n20783 ;
  assign n21389 = n21322 & n21388 ;
  assign n21390 = ~n21387 & ~n21389 ;
  assign n21391 = n21363 & n21390 ;
  assign n21392 = ~n21362 & ~n21391 ;
  assign n21393 = ~\pi0120  & ~n21322 ;
  assign n21394 = \pi0120  & \pi0824  ;
  assign n21395 = n6720 & n21394 ;
  assign n21396 = n6719 & n21395 ;
  assign n21397 = ~\pi1091  & ~n21396 ;
  assign n21398 = ~n21290 & n21397 ;
  assign n21399 = ~n21393 & n21398 ;
  assign n21400 = n16869 & n21385 ;
  assign n21401 = ~\pi0120  & \pi1091  ;
  assign n21402 = n21322 & n21401 ;
  assign n21403 = ~n21400 & ~n21402 ;
  assign n21404 = ~n6706 & n21403 ;
  assign n21405 = ~n21399 & n21404 ;
  assign n21406 = n6709 & ~n21352 ;
  assign n21407 = ~n21405 & n21406 ;
  assign n21408 = n21392 & n21407 ;
  assign n21409 = ~n6709 & n21370 ;
  assign n21410 = ~n21371 & n21409 ;
  assign n21411 = n21392 & n21410 ;
  assign n21412 = ~n6709 & n21375 ;
  assign n21413 = ~n21285 & n21412 ;
  assign n21414 = n6761 & ~n21413 ;
  assign n21415 = ~n21411 & n21414 ;
  assign n21416 = ~n21408 & n21415 ;
  assign n21417 = n1689 & ~n20784 ;
  assign n21418 = ~n6706 & n21417 ;
  assign n21419 = ~n21285 & n21418 ;
  assign n21420 = n6712 & n21403 ;
  assign n21421 = n21419 & ~n21420 ;
  assign n21422 = ~n21403 & n21417 ;
  assign n21423 = ~n21393 & n21417 ;
  assign n21424 = n21398 & n21423 ;
  assign n21425 = ~n21422 & ~n21424 ;
  assign n21426 = n6706 & ~n21420 ;
  assign n21427 = ~n21425 & n21426 ;
  assign n21428 = ~n21421 & ~n21427 ;
  assign n21429 = ~n6709 & ~n6761 ;
  assign n21430 = n21428 & n21429 ;
  assign n21431 = n6709 & ~n6761 ;
  assign n21432 = n21425 & n21431 ;
  assign n21433 = \pi0223  & ~n21432 ;
  assign n21434 = ~n21430 & n21433 ;
  assign n21435 = ~n21416 & n21434 ;
  assign n21436 = n2165 & ~n20784 ;
  assign n21437 = ~n21285 & n21436 ;
  assign n21438 = ~n21435 & ~n21437 ;
  assign n21439 = ~n21380 & n21438 ;
  assign n21440 = ~n21351 & n21439 ;
  assign n21441 = \pi0223  & ~n21435 ;
  assign n21442 = n6205 & ~n21441 ;
  assign n21443 = ~n21440 & n21442 ;
  assign n21444 = ~n2352 & ~n6732 ;
  assign n21445 = n21350 & n21444 ;
  assign n21446 = ~n2352 & n6732 ;
  assign n21447 = ~n21378 & n21446 ;
  assign n21448 = ~n21367 & n21447 ;
  assign n21449 = n6732 & ~n21413 ;
  assign n21450 = ~n21411 & n21449 ;
  assign n21451 = ~n21408 & n21450 ;
  assign n21452 = ~n6709 & ~n6732 ;
  assign n21453 = n21428 & n21452 ;
  assign n21454 = n6709 & ~n6732 ;
  assign n21455 = n21425 & n21454 ;
  assign n21456 = \pi0215  & ~n21455 ;
  assign n21457 = ~n21453 & n21456 ;
  assign n21458 = ~n21451 & n21457 ;
  assign n21459 = n2352 & ~n20784 ;
  assign n21460 = ~n21285 & n21459 ;
  assign n21461 = ~n21458 & ~n21460 ;
  assign n21462 = ~n21448 & n21461 ;
  assign n21463 = ~n21445 & n21462 ;
  assign n21464 = \pi0215  & ~n21458 ;
  assign n21465 = n2297 & ~n21464 ;
  assign n21466 = ~n21463 & n21465 ;
  assign n21467 = ~n21443 & ~n21466 ;
  assign n21468 = ~\pi0761  & ~n21467 ;
  assign n21469 = ~\pi0140  & ~n21468 ;
  assign n21470 = ~n21274 & n21469 ;
  assign n21471 = ~\pi0039  & \pi0299  ;
  assign n21472 = n21237 & n21262 ;
  assign n21473 = n21204 & ~n21254 ;
  assign n21474 = \pi0603  & ~n21473 ;
  assign n21475 = ~n21472 & n21474 ;
  assign n21476 = n21471 & ~n21475 ;
  assign n21477 = \pi0198  & \pi0603  ;
  assign n21478 = ~n21263 & n21477 ;
  assign n21479 = ~\pi0039  & ~\pi0299  ;
  assign n21480 = ~\pi0198  & \pi0603  ;
  assign n21481 = ~n21255 & n21480 ;
  assign n21482 = n21479 & ~n21481 ;
  assign n21483 = ~n21478 & n21482 ;
  assign n21484 = ~n21476 & ~n21483 ;
  assign n21485 = \pi0140  & ~\pi0761  ;
  assign n21486 = n20784 & ~n21359 ;
  assign n21487 = n6709 & ~n21486 ;
  assign n21488 = n20784 & n21370 ;
  assign n21489 = ~n21359 & n21488 ;
  assign n21490 = n20784 & ~n21370 ;
  assign n21491 = ~n21285 & n21490 ;
  assign n21492 = ~n6709 & ~n21491 ;
  assign n21493 = ~n21489 & n21492 ;
  assign n21494 = ~n21487 & ~n21493 ;
  assign n21495 = n21446 & n21494 ;
  assign n21496 = n20784 & ~n21334 ;
  assign n21497 = n6713 & n20784 ;
  assign n21498 = ~n21329 & n21497 ;
  assign n21499 = ~n21496 & ~n21498 ;
  assign n21500 = n21444 & ~n21499 ;
  assign n21501 = ~n21495 & ~n21500 ;
  assign n21502 = ~\pi0120  & n2352 ;
  assign n21503 = n21277 & n21502 ;
  assign n21504 = n1281 & n21503 ;
  assign n21505 = n1260 & n21504 ;
  assign n21506 = \pi0120  & n2352 ;
  assign n21507 = n1281 & n21506 ;
  assign n21508 = n1260 & n21507 ;
  assign n21509 = ~n21505 & ~n21508 ;
  assign n21510 = n1689 & n20784 ;
  assign n21511 = ~n21509 & n21510 ;
  assign n21512 = ~\pi0215  & ~n21511 ;
  assign n21513 = n21501 & n21512 ;
  assign n21514 = ~n6706 & n20784 ;
  assign n21515 = ~n21285 & n21514 ;
  assign n21516 = n20784 & ~n21285 ;
  assign n21517 = n6706 & ~n21403 ;
  assign n21518 = n6706 & ~n21393 ;
  assign n21519 = n21398 & n21518 ;
  assign n21520 = ~n21517 & ~n21519 ;
  assign n21521 = n21516 & ~n21520 ;
  assign n21522 = ~n21515 & ~n21521 ;
  assign n21523 = ~n6706 & n21370 ;
  assign n21524 = n21403 & n21523 ;
  assign n21525 = ~n21399 & n21524 ;
  assign n21526 = ~n6709 & ~n21525 ;
  assign n21527 = ~n21522 & n21526 ;
  assign n21528 = ~n21405 & n21516 ;
  assign n21529 = \pi0215  & ~n21528 ;
  assign n21530 = ~n21527 & n21529 ;
  assign n21531 = ~n6732 & ~n21286 ;
  assign n21532 = \pi0215  & n21531 ;
  assign n21533 = n21520 & n21532 ;
  assign n21534 = \pi0299  & ~n21533 ;
  assign n21535 = ~n21530 & n21534 ;
  assign n21536 = ~n21513 & n21535 ;
  assign n21537 = \pi0223  & ~n21528 ;
  assign n21538 = ~n21527 & n21537 ;
  assign n21539 = ~n6761 & ~n21286 ;
  assign n21540 = \pi0223  & n21539 ;
  assign n21541 = n21520 & n21540 ;
  assign n21542 = ~\pi0299  & ~n21541 ;
  assign n21543 = ~n21538 & n21542 ;
  assign n21544 = \pi0039  & ~n21543 ;
  assign n21545 = ~n2165 & n20784 ;
  assign n21546 = ~n21334 & n21545 ;
  assign n21547 = n6713 & n21545 ;
  assign n21548 = ~n21329 & n21547 ;
  assign n21549 = ~n21546 & ~n21548 ;
  assign n21550 = ~n21368 & n21549 ;
  assign n21551 = n6761 & ~n21494 ;
  assign n21552 = ~n21550 & ~n21551 ;
  assign n21553 = ~\pi0120  & n2165 ;
  assign n21554 = n21277 & n21553 ;
  assign n21555 = n1281 & n21554 ;
  assign n21556 = n1260 & n21555 ;
  assign n21557 = \pi0120  & n2165 ;
  assign n21558 = n1281 & n21557 ;
  assign n21559 = n1260 & n21558 ;
  assign n21560 = ~n21556 & ~n21559 ;
  assign n21561 = n21510 & ~n21560 ;
  assign n21562 = ~\pi0223  & ~n21561 ;
  assign n21563 = \pi0039  & n21562 ;
  assign n21564 = ~n21552 & n21563 ;
  assign n21565 = ~n21544 & ~n21564 ;
  assign n21566 = ~n21536 & ~n21565 ;
  assign n21567 = n21485 & ~n21566 ;
  assign n21568 = n21484 & n21567 ;
  assign n21569 = ~n21470 & ~n21568 ;
  assign n21570 = \pi0616  & n21285 ;
  assign n21571 = \pi0616  & ~n21570 ;
  assign n21572 = \pi0603  & ~\pi0642  ;
  assign n21573 = ~n21359 & n21572 ;
  assign n21574 = ~n21285 & ~n21572 ;
  assign n21575 = ~\pi0614  & ~n21574 ;
  assign n21576 = ~n21573 & n21575 ;
  assign n21577 = \pi0614  & n21285 ;
  assign n21578 = ~n21570 & ~n21577 ;
  assign n21579 = ~n21576 & n21578 ;
  assign n21580 = ~n21571 & ~n21579 ;
  assign n21581 = \pi0681  & n21580 ;
  assign n21582 = ~\pi0680  & n21285 ;
  assign n21583 = \pi0614  & ~\pi0662  ;
  assign n21584 = n6708 & n21583 ;
  assign n21585 = ~n21582 & n21584 ;
  assign n21586 = ~\pi0662  & n6708 ;
  assign n21587 = \pi0614  & ~n21586 ;
  assign n21588 = ~n21285 & n21587 ;
  assign n21589 = ~\pi0681  & ~n21588 ;
  assign n21590 = ~n21585 & n21589 ;
  assign n21591 = \pi0680  & n21589 ;
  assign n21592 = n21359 & n21591 ;
  assign n21593 = ~n21590 & ~n21592 ;
  assign n21594 = n6761 & n21593 ;
  assign n21595 = ~n21573 & ~n21574 ;
  assign n21596 = ~\pi0614  & n6709 ;
  assign n21597 = ~n21359 & n21596 ;
  assign n21598 = ~\pi0616  & ~n21597 ;
  assign n21599 = n21595 & n21598 ;
  assign n21600 = ~\pi0614  & ~n6709 ;
  assign n21601 = ~n21570 & n21600 ;
  assign n21602 = ~n21597 & ~n21601 ;
  assign n21603 = n6761 & ~n21602 ;
  assign n21604 = ~n21599 & n21603 ;
  assign n21605 = ~n21594 & ~n21604 ;
  assign n21606 = ~n21581 & ~n21605 ;
  assign n21607 = n2165 & ~n21285 ;
  assign n21608 = ~\pi0223  & ~n21607 ;
  assign n21609 = ~n6761 & ~n21334 ;
  assign n21610 = n6713 & ~n6761 ;
  assign n21611 = ~n21329 & n21610 ;
  assign n21612 = ~n21609 & ~n21611 ;
  assign n21613 = n21608 & n21612 ;
  assign n21614 = ~n21606 & n21613 ;
  assign n21615 = ~n21286 & n21520 ;
  assign n21616 = \pi0681  & n21615 ;
  assign n21617 = ~n6706 & n6710 ;
  assign n21618 = n21403 & n21617 ;
  assign n21619 = ~n21399 & n21618 ;
  assign n21620 = ~n6710 & n21285 ;
  assign n21621 = n6706 & n6710 ;
  assign n21622 = n21285 & n21621 ;
  assign n21623 = ~n21620 & ~n21622 ;
  assign n21624 = ~n21619 & n21623 ;
  assign n21625 = \pi0681  & n6711 ;
  assign n21626 = ~n21624 & n21625 ;
  assign n21627 = ~n21616 & ~n21626 ;
  assign n21628 = ~n6761 & ~n21627 ;
  assign n21629 = ~\pi0661  & ~n21520 ;
  assign n21630 = ~n21577 & n21623 ;
  assign n21631 = ~n21619 & n21630 ;
  assign n21632 = \pi0614  & ~n21285 ;
  assign n21633 = ~\pi0616  & ~n6707 ;
  assign n21634 = ~n21632 & n21633 ;
  assign n21635 = ~n21631 & n21634 ;
  assign n21636 = \pi0616  & ~n6707 ;
  assign n21637 = n21285 & n21636 ;
  assign n21638 = n6707 & n21403 ;
  assign n21639 = ~n21399 & n21638 ;
  assign n21640 = ~\pi0661  & ~n6706 ;
  assign n21641 = ~n21639 & n21640 ;
  assign n21642 = ~n21637 & n21641 ;
  assign n21643 = ~n21635 & n21642 ;
  assign n21644 = ~n21629 & ~n21643 ;
  assign n21645 = n6711 & ~n21624 ;
  assign n21646 = \pi0661  & ~n21615 ;
  assign n21647 = ~n21645 & n21646 ;
  assign n21648 = ~\pi0681  & ~n6761 ;
  assign n21649 = ~n21647 & n21648 ;
  assign n21650 = n21644 & n21649 ;
  assign n21651 = ~n21628 & ~n21650 ;
  assign n21652 = \pi0223  & ~n21651 ;
  assign n21653 = \pi0616  & \pi0681  ;
  assign n21654 = n21285 & n21653 ;
  assign n21655 = ~\pi0616  & \pi0681  ;
  assign n21656 = ~n21632 & n21655 ;
  assign n21657 = ~n21631 & n21656 ;
  assign n21658 = ~n21654 & ~n21657 ;
  assign n21659 = ~n21631 & ~n21632 ;
  assign n21660 = ~\pi0616  & ~n21586 ;
  assign n21661 = ~n21659 & n21660 ;
  assign n21662 = \pi0616  & ~\pi0662  ;
  assign n21663 = n6708 & n21662 ;
  assign n21664 = ~n21582 & n21663 ;
  assign n21665 = ~\pi0680  & n21664 ;
  assign n21666 = ~n21352 & n21664 ;
  assign n21667 = ~n21405 & n21666 ;
  assign n21668 = ~n21665 & ~n21667 ;
  assign n21669 = ~n21661 & n21668 ;
  assign n21670 = ~\pi0616  & ~\pi0680  ;
  assign n21671 = ~n21632 & n21670 ;
  assign n21672 = ~n21631 & n21671 ;
  assign n21673 = ~\pi0616  & ~\pi0662  ;
  assign n21674 = n6708 & n21673 ;
  assign n21675 = ~\pi0680  & n21674 ;
  assign n21676 = ~n21352 & n21674 ;
  assign n21677 = ~n21405 & n21676 ;
  assign n21678 = ~n21675 & ~n21677 ;
  assign n21679 = ~n21672 & ~n21678 ;
  assign n21680 = \pi0616  & ~n21586 ;
  assign n21681 = ~n21285 & n21680 ;
  assign n21682 = ~\pi0681  & ~n21681 ;
  assign n21683 = ~n21679 & n21682 ;
  assign n21684 = n21669 & n21683 ;
  assign n21685 = n21658 & ~n21684 ;
  assign n21686 = \pi0223  & n6761 ;
  assign n21687 = ~n21685 & n21686 ;
  assign n21688 = ~n21652 & ~n21687 ;
  assign n21689 = ~\pi0223  & n2165 ;
  assign n21690 = n21285 & n21689 ;
  assign n21691 = n21688 & ~n21690 ;
  assign n21692 = ~n21614 & n21691 ;
  assign n21693 = ~\pi0299  & ~n21692 ;
  assign n21694 = n6728 & n6729 ;
  assign n21695 = n21334 & ~n21694 ;
  assign n21696 = ~n21330 & n21695 ;
  assign n21697 = ~n2352 & n6730 ;
  assign n21698 = ~n21696 & n21697 ;
  assign n21699 = ~n2352 & ~n6730 ;
  assign n21700 = ~n21334 & n21699 ;
  assign n21701 = n6713 & n21699 ;
  assign n21702 = ~n21329 & n21701 ;
  assign n21703 = ~n21700 & ~n21702 ;
  assign n21704 = n2352 & ~n21285 ;
  assign n21705 = ~\pi0215  & ~n21704 ;
  assign n21706 = \pi0299  & n21705 ;
  assign n21707 = n21703 & n21706 ;
  assign n21708 = ~n21698 & n21707 ;
  assign n21709 = ~n21599 & ~n21602 ;
  assign n21710 = ~n21593 & ~n21709 ;
  assign n21711 = ~n21581 & ~n21710 ;
  assign n21712 = n21694 & n21707 ;
  assign n21713 = ~n21711 & n21712 ;
  assign n21714 = ~n21708 & ~n21713 ;
  assign n21715 = n6730 & ~n21694 ;
  assign n21716 = n6730 & n21658 ;
  assign n21717 = ~n21684 & n21716 ;
  assign n21718 = ~n21715 & ~n21717 ;
  assign n21719 = ~\pi0681  & ~n21694 ;
  assign n21720 = ~n21647 & n21719 ;
  assign n21721 = n21644 & n21720 ;
  assign n21722 = ~n21627 & ~n21694 ;
  assign n21723 = ~n21721 & ~n21722 ;
  assign n21724 = ~n21718 & n21723 ;
  assign n21725 = ~\pi0681  & ~n21647 ;
  assign n21726 = n21644 & n21725 ;
  assign n21727 = ~n6730 & n21627 ;
  assign n21728 = ~n21726 & n21727 ;
  assign n21729 = \pi0215  & ~n21728 ;
  assign n21730 = \pi0299  & n21729 ;
  assign n21731 = ~n21724 & n21730 ;
  assign n21732 = \pi0039  & ~n21731 ;
  assign n21733 = n21714 & n21732 ;
  assign n21734 = ~n21693 & n21733 ;
  assign n21735 = ~n21205 & n21471 ;
  assign n21736 = ~n21238 & n21735 ;
  assign n21737 = \pi0198  & n21236 ;
  assign n21738 = n21232 & n21737 ;
  assign n21739 = ~\pi0198  & n21203 ;
  assign n21740 = ~n21199 & n21739 ;
  assign n21741 = n21479 & ~n21740 ;
  assign n21742 = ~n21738 & n21741 ;
  assign n21743 = ~n21736 & ~n21742 ;
  assign n21744 = ~n21734 & n21743 ;
  assign n21745 = \pi0761  & ~n21744 ;
  assign n21746 = ~n21569 & ~n21745 ;
  assign n21747 = ~\pi0038  & n21746 ;
  assign n21748 = \pi0038  & \pi0603  ;
  assign n21749 = ~n20783 & n21748 ;
  assign n21750 = n20785 & n21749 ;
  assign n21751 = n1354 & n21750 ;
  assign n21752 = n8413 & n21751 ;
  assign n21753 = n1358 & n21752 ;
  assign n21754 = n1689 & n6784 ;
  assign n21755 = n1266 & n21754 ;
  assign n21756 = n1354 & n21755 ;
  assign n21757 = n1358 & n21756 ;
  assign n21758 = \pi0038  & ~\pi0140  ;
  assign n21759 = ~n21757 & n21758 ;
  assign n21760 = ~n21753 & ~n21759 ;
  assign n21761 = n6861 & n21760 ;
  assign n21762 = ~n21747 & n21761 ;
  assign n21763 = \pi0140  & ~n6861 ;
  assign n21764 = ~\pi0038  & n6861 ;
  assign n21765 = n1689 & n4520 ;
  assign n21766 = n6861 & n21765 ;
  assign n21767 = n1638 & n21766 ;
  assign n21768 = ~n21764 & ~n21767 ;
  assign n21769 = ~\pi0140  & n21768 ;
  assign n21770 = ~\pi0038  & n21743 ;
  assign n21771 = ~\pi0140  & n21770 ;
  assign n21772 = ~n21734 & n21771 ;
  assign n21773 = ~n21769 & ~n21772 ;
  assign n21774 = \pi0609  & \pi1155  ;
  assign n21775 = \pi0785  & ~n20999 ;
  assign n21776 = ~n21774 & n21775 ;
  assign n21777 = ~n20985 & ~n21776 ;
  assign n21778 = n21773 & ~n21777 ;
  assign n21779 = ~n21763 & ~n21778 ;
  assign n21780 = ~n21762 & n21779 ;
  assign n21781 = ~n21773 & ~n21777 ;
  assign n21782 = ~\pi0781  & ~n21781 ;
  assign n21783 = ~n21780 & n21782 ;
  assign n21784 = ~\pi0789  & n21783 ;
  assign n21785 = ~\pi0140  & ~\pi0618  ;
  assign n21786 = n21768 & n21785 ;
  assign n21787 = n21770 & n21785 ;
  assign n21788 = ~n21734 & n21787 ;
  assign n21789 = ~n21786 & ~n21788 ;
  assign n21790 = \pi1154  & n21789 ;
  assign n21791 = ~\pi0618  & n21790 ;
  assign n21792 = ~n21781 & n21790 ;
  assign n21793 = ~n21780 & n21792 ;
  assign n21794 = ~n21791 & ~n21793 ;
  assign n21795 = ~\pi0140  & \pi0618  ;
  assign n21796 = n21768 & n21795 ;
  assign n21797 = n21770 & n21795 ;
  assign n21798 = ~n21734 & n21797 ;
  assign n21799 = ~n21796 & ~n21798 ;
  assign n21800 = ~\pi1154  & n21799 ;
  assign n21801 = \pi0618  & n21800 ;
  assign n21802 = ~n21781 & n21800 ;
  assign n21803 = ~n21780 & n21802 ;
  assign n21804 = ~n21801 & ~n21803 ;
  assign n21805 = n21794 & n21804 ;
  assign n21806 = \pi0781  & ~\pi0789  ;
  assign n21807 = ~n21805 & n21806 ;
  assign n21808 = ~n21784 & ~n21807 ;
  assign n21809 = ~\pi0788  & ~n21808 ;
  assign n21810 = ~\pi0619  & ~n21783 ;
  assign n21811 = n20823 & n21768 ;
  assign n21812 = n20823 & n21770 ;
  assign n21813 = ~n21734 & n21812 ;
  assign n21814 = ~n21811 & ~n21813 ;
  assign n21815 = ~\pi1159  & n21814 ;
  assign n21816 = ~n21810 & n21815 ;
  assign n21817 = \pi0781  & n21815 ;
  assign n21818 = ~n21805 & n21817 ;
  assign n21819 = ~n21816 & ~n21818 ;
  assign n21820 = \pi0619  & ~n21783 ;
  assign n21821 = ~\pi0140  & ~\pi0619  ;
  assign n21822 = n21768 & n21821 ;
  assign n21823 = n21770 & n21821 ;
  assign n21824 = ~n21734 & n21823 ;
  assign n21825 = ~n21822 & ~n21824 ;
  assign n21826 = \pi1159  & n21825 ;
  assign n21827 = ~n21820 & n21826 ;
  assign n21828 = \pi0781  & n21826 ;
  assign n21829 = ~n21805 & n21828 ;
  assign n21830 = ~n21827 & ~n21829 ;
  assign n21831 = n21819 & n21830 ;
  assign n21832 = ~\pi0788  & \pi0789  ;
  assign n21833 = ~n21831 & n21832 ;
  assign n21834 = ~n21809 & ~n21833 ;
  assign n21835 = ~\pi0628  & n21834 ;
  assign n21836 = \pi1156  & ~n21835 ;
  assign n21837 = ~\pi0626  & n21808 ;
  assign n21838 = ~\pi0140  & \pi0626  ;
  assign n21839 = n21768 & n21838 ;
  assign n21840 = n21770 & n21838 ;
  assign n21841 = ~n21734 & n21840 ;
  assign n21842 = ~n21839 & ~n21841 ;
  assign n21843 = ~\pi1158  & n21842 ;
  assign n21844 = ~n21837 & n21843 ;
  assign n21845 = \pi0789  & n21843 ;
  assign n21846 = ~n21831 & n21845 ;
  assign n21847 = ~n21844 & ~n21846 ;
  assign n21848 = \pi0626  & n21808 ;
  assign n21849 = ~\pi0140  & ~\pi0626  ;
  assign n21850 = n21768 & n21849 ;
  assign n21851 = n21770 & n21849 ;
  assign n21852 = ~n21734 & n21851 ;
  assign n21853 = ~n21850 & ~n21852 ;
  assign n21854 = \pi1158  & n21853 ;
  assign n21855 = ~n21848 & n21854 ;
  assign n21856 = \pi0789  & n21854 ;
  assign n21857 = ~n21831 & n21856 ;
  assign n21858 = ~n21855 & ~n21857 ;
  assign n21859 = n21847 & n21858 ;
  assign n21860 = \pi0788  & \pi1156  ;
  assign n21861 = ~n21859 & n21860 ;
  assign n21862 = ~n21836 & ~n21861 ;
  assign n21863 = ~\pi0140  & \pi0628  ;
  assign n21864 = n21768 & n21863 ;
  assign n21865 = n21770 & n21863 ;
  assign n21866 = ~n21734 & n21865 ;
  assign n21867 = ~n21864 & ~n21866 ;
  assign n21868 = ~\pi1156  & n21867 ;
  assign n21869 = \pi0629  & ~n21868 ;
  assign n21870 = ~\pi0140  & ~\pi0625  ;
  assign n21871 = n21768 & n21870 ;
  assign n21872 = n21770 & n21870 ;
  assign n21873 = ~n21734 & n21872 ;
  assign n21874 = ~n21871 & ~n21873 ;
  assign n21875 = \pi1153  & n21874 ;
  assign n21876 = n20854 & ~n21285 ;
  assign n21877 = \pi0680  & n6706 ;
  assign n21878 = ~n21876 & n21877 ;
  assign n21879 = n21586 & n21878 ;
  assign n21880 = n20854 & ~n21290 ;
  assign n21881 = ~n21325 & n21880 ;
  assign n21882 = \pi0680  & ~n6706 ;
  assign n21883 = n21586 & n21882 ;
  assign n21884 = ~n21881 & n21883 ;
  assign n21885 = ~n21879 & ~n21884 ;
  assign n21886 = ~n6706 & ~n21881 ;
  assign n21887 = n6706 & ~n21876 ;
  assign n21888 = n6712 & ~n21887 ;
  assign n21889 = ~n21886 & n21888 ;
  assign n21890 = ~n6712 & n20854 ;
  assign n21891 = ~n21285 & n21890 ;
  assign n21892 = \pi0680  & ~n21891 ;
  assign n21893 = ~n21586 & n21892 ;
  assign n21894 = ~n21889 & n21893 ;
  assign n21895 = n21885 & ~n21894 ;
  assign n21896 = n2165 & ~n20855 ;
  assign n21897 = ~n21285 & n21896 ;
  assign n21898 = n6761 & ~n21897 ;
  assign n21899 = ~n21895 & n21898 ;
  assign n21900 = ~\pi0680  & n21898 ;
  assign n21901 = n21580 & n21900 ;
  assign n21902 = ~n21899 & ~n21901 ;
  assign n21903 = ~n21290 & ~n21325 ;
  assign n21904 = n6712 & ~n21306 ;
  assign n21905 = ~n21903 & n21904 ;
  assign n21906 = ~\pi0680  & ~n6761 ;
  assign n21907 = n21905 & n21906 ;
  assign n21908 = ~n6712 & ~n21286 ;
  assign n21909 = n21906 & n21908 ;
  assign n21910 = n21328 & n21909 ;
  assign n21911 = ~n21907 & ~n21910 ;
  assign n21912 = ~n6735 & n20854 ;
  assign n21913 = ~n21290 & n21912 ;
  assign n21914 = ~n21325 & n21913 ;
  assign n21915 = ~n6706 & n20854 ;
  assign n21916 = ~n6712 & n21915 ;
  assign n21917 = ~n21285 & n21916 ;
  assign n21918 = ~n21914 & ~n21917 ;
  assign n21919 = ~n21586 & ~n21918 ;
  assign n21920 = n20854 & n21586 ;
  assign n21921 = ~n21290 & n21920 ;
  assign n21922 = ~n21325 & n21921 ;
  assign n21923 = \pi0680  & ~n21922 ;
  assign n21924 = ~n6761 & n21923 ;
  assign n21925 = ~n21919 & n21924 ;
  assign n21926 = ~n2165 & ~n21925 ;
  assign n21927 = n21911 & n21926 ;
  assign n21928 = ~n21897 & ~n21927 ;
  assign n21929 = n3058 & ~n21928 ;
  assign n21930 = n21902 & n21929 ;
  assign n21931 = n1689 & ~n20855 ;
  assign n21932 = ~n21509 & n21931 ;
  assign n21933 = n6732 & ~n21932 ;
  assign n21934 = ~n21895 & n21933 ;
  assign n21935 = ~\pi0680  & n21933 ;
  assign n21936 = n21580 & n21935 ;
  assign n21937 = ~n21934 & ~n21936 ;
  assign n21938 = ~\pi0680  & ~n6732 ;
  assign n21939 = n21905 & n21938 ;
  assign n21940 = n21908 & n21938 ;
  assign n21941 = n21328 & n21940 ;
  assign n21942 = ~n21939 & ~n21941 ;
  assign n21943 = ~n6732 & n21923 ;
  assign n21944 = ~n21919 & n21943 ;
  assign n21945 = ~n2352 & ~n21944 ;
  assign n21946 = n21942 & n21945 ;
  assign n21947 = ~n21932 & ~n21946 ;
  assign n21948 = ~\pi0215  & \pi0299  ;
  assign n21949 = ~n21947 & n21948 ;
  assign n21950 = n21937 & n21949 ;
  assign n21951 = ~\pi0680  & n21615 ;
  assign n21952 = ~\pi0680  & n6711 ;
  assign n21953 = ~n21624 & n21952 ;
  assign n21954 = ~n21951 & ~n21953 ;
  assign n21955 = \pi0120  & n20854 ;
  assign n21956 = n21385 & n21955 ;
  assign n21957 = ~\pi0120  & n20854 ;
  assign n21958 = n21322 & n21957 ;
  assign n21959 = ~n21956 & ~n21958 ;
  assign n21960 = \pi0680  & n21959 ;
  assign n21961 = ~n21917 & n21960 ;
  assign n21962 = ~n6706 & n21959 ;
  assign n21963 = ~n21887 & ~n21962 ;
  assign n21964 = ~n6709 & ~n21892 ;
  assign n21965 = ~n21963 & ~n21964 ;
  assign n21966 = \pi0215  & ~n21965 ;
  assign n21967 = ~n21961 & n21966 ;
  assign n21968 = n21954 & n21967 ;
  assign n21969 = ~n6734 & ~n21968 ;
  assign n21970 = n21892 & ~n21963 ;
  assign n21971 = \pi0616  & ~\pi0680  ;
  assign n21972 = n21285 & n21971 ;
  assign n21973 = ~n6706 & n6709 ;
  assign n21974 = n21959 & n21973 ;
  assign n21975 = n6706 & n6709 ;
  assign n21976 = ~n21876 & n21975 ;
  assign n21977 = ~n21974 & ~n21976 ;
  assign n21978 = ~n21972 & n21977 ;
  assign n21979 = ~n21970 & n21978 ;
  assign n21980 = ~n21672 & n21979 ;
  assign n21981 = n6732 & ~n21980 ;
  assign n21982 = \pi0299  & ~n21981 ;
  assign n21983 = ~n21969 & n21982 ;
  assign n21984 = \pi0223  & ~n21965 ;
  assign n21985 = ~n21961 & n21984 ;
  assign n21986 = n21954 & n21985 ;
  assign n21987 = ~n21686 & ~n21986 ;
  assign n21988 = n6761 & ~n21980 ;
  assign n21989 = ~\pi0299  & ~n21988 ;
  assign n21990 = ~n21987 & n21989 ;
  assign n21991 = ~n21983 & ~n21990 ;
  assign n21992 = ~n21950 & n21991 ;
  assign n21993 = ~n21930 & n21992 ;
  assign n21994 = \pi0039  & ~n21993 ;
  assign n21995 = \pi0665  & ~n21198 ;
  assign n21996 = ~n21194 & n21995 ;
  assign n21997 = ~\pi0210  & \pi0680  ;
  assign n21998 = ~n21996 & n21997 ;
  assign n21999 = n1686 & n21995 ;
  assign n22000 = \pi1093  & n21995 ;
  assign n22001 = ~n21229 & n22000 ;
  assign n22002 = ~n21999 & ~n22001 ;
  assign n22003 = \pi0210  & \pi0680  ;
  assign n22004 = n22002 & n22003 ;
  assign n22005 = ~n21998 & ~n22004 ;
  assign n22006 = n21239 & n22005 ;
  assign n22007 = \pi0299  & ~n22006 ;
  assign n22008 = ~\pi0198  & \pi0680  ;
  assign n22009 = ~n21996 & n22008 ;
  assign n22010 = ~n21740 & ~n22009 ;
  assign n22011 = ~n21738 & n22010 ;
  assign n22012 = \pi0198  & \pi0680  ;
  assign n22013 = n22002 & n22012 ;
  assign n22014 = ~\pi0039  & ~n22013 ;
  assign n22015 = n22011 & n22014 ;
  assign n22016 = ~n21471 & ~n22015 ;
  assign n22017 = ~n22007 & ~n22016 ;
  assign n22018 = ~\pi0140  & ~n22017 ;
  assign n22019 = ~n21994 & n22018 ;
  assign n22020 = ~\pi0038  & ~\pi0140  ;
  assign n22021 = ~\pi0665  & ~n21290 ;
  assign n22022 = ~n21325 & n22021 ;
  assign n22023 = ~n20854 & ~n21285 ;
  assign n22024 = ~n21306 & ~n22023 ;
  assign n22025 = ~n22022 & n22024 ;
  assign n22026 = ~n21359 & ~n22025 ;
  assign n22027 = n21586 & ~n22026 ;
  assign n22028 = \pi0680  & ~n22027 ;
  assign n22029 = ~n6712 & ~n20854 ;
  assign n22030 = ~n21285 & n22029 ;
  assign n22031 = ~n21586 & ~n22030 ;
  assign n22032 = ~n2352 & ~n22031 ;
  assign n22033 = n6712 & ~n21359 ;
  assign n22034 = ~n2352 & ~n22025 ;
  assign n22035 = n22033 & n22034 ;
  assign n22036 = ~n22032 & ~n22035 ;
  assign n22037 = n22028 & ~n22036 ;
  assign n22038 = ~n21444 & ~n22037 ;
  assign n22039 = n21328 & n21908 ;
  assign n22040 = n20855 & ~n21586 ;
  assign n22041 = ~n21905 & n22040 ;
  assign n22042 = ~n22039 & n22041 ;
  assign n22043 = ~n6732 & ~n21306 ;
  assign n22044 = ~n22022 & n22043 ;
  assign n22045 = ~n21452 & ~n22044 ;
  assign n22046 = ~n22042 & ~n22045 ;
  assign n22047 = ~\pi0215  & ~n22046 ;
  assign n22048 = ~n22038 & n22047 ;
  assign n22049 = n2352 & n20855 ;
  assign n22050 = ~\pi0215  & n22049 ;
  assign n22051 = ~n21285 & n22050 ;
  assign n22052 = \pi0680  & n22023 ;
  assign n22053 = n21405 & ~n22030 ;
  assign n22054 = n22052 & ~n22053 ;
  assign n22055 = n21520 & n21531 ;
  assign n22056 = \pi0215  & ~n21586 ;
  assign n22057 = \pi0215  & n22023 ;
  assign n22058 = ~n21405 & n22057 ;
  assign n22059 = ~n22056 & ~n22058 ;
  assign n22060 = ~n22055 & ~n22059 ;
  assign n22061 = n22054 & n22060 ;
  assign n22062 = ~n22051 & ~n22061 ;
  assign n22063 = ~n22048 & n22062 ;
  assign n22064 = n2297 & ~n22063 ;
  assign n22065 = ~n22025 & n22033 ;
  assign n22066 = n22031 & ~n22065 ;
  assign n22067 = n22028 & ~n22066 ;
  assign n22068 = n6761 & ~n22067 ;
  assign n22069 = ~n6761 & ~n21306 ;
  assign n22070 = ~n22022 & n22069 ;
  assign n22071 = ~n21429 & ~n22070 ;
  assign n22072 = ~n22042 & ~n22071 ;
  assign n22073 = ~\pi0223  & ~n22072 ;
  assign n22074 = ~n2165 & n22073 ;
  assign n22075 = ~n22068 & n22074 ;
  assign n22076 = n2165 & n20855 ;
  assign n22077 = ~\pi0223  & n22076 ;
  assign n22078 = ~n21285 & n22077 ;
  assign n22079 = n21520 & n21539 ;
  assign n22080 = \pi0223  & ~n21586 ;
  assign n22081 = \pi0223  & n22023 ;
  assign n22082 = ~n21405 & n22081 ;
  assign n22083 = ~n22080 & ~n22082 ;
  assign n22084 = ~n22079 & ~n22083 ;
  assign n22085 = n22054 & n22084 ;
  assign n22086 = ~n22078 & ~n22085 ;
  assign n22087 = ~n22075 & n22086 ;
  assign n22088 = n6205 & ~n22087 ;
  assign n22089 = ~n22064 & ~n22088 ;
  assign n22090 = ~\pi0665  & ~n21198 ;
  assign n22091 = n1686 & n22090 ;
  assign n22092 = \pi1093  & n22090 ;
  assign n22093 = ~n21229 & n22092 ;
  assign n22094 = ~n22091 & ~n22093 ;
  assign n22095 = n21237 & n22094 ;
  assign n22096 = ~n21194 & n22090 ;
  assign n22097 = n21204 & ~n22096 ;
  assign n22098 = \pi0680  & ~n22097 ;
  assign n22099 = ~n22095 & n22098 ;
  assign n22100 = \pi0299  & ~n22099 ;
  assign n22101 = n21737 & n22094 ;
  assign n22102 = n21739 & ~n22096 ;
  assign n22103 = \pi0680  & ~n22102 ;
  assign n22104 = ~\pi0039  & n22103 ;
  assign n22105 = ~n22101 & n22104 ;
  assign n22106 = ~n21471 & ~n22105 ;
  assign n22107 = ~n22100 & ~n22106 ;
  assign n22108 = ~\pi0038  & ~n22107 ;
  assign n22109 = n22089 & n22108 ;
  assign n22110 = ~n22020 & ~n22109 ;
  assign n22111 = ~n22019 & ~n22110 ;
  assign n22112 = ~\pi0140  & ~n21757 ;
  assign n22113 = n1689 & n20855 ;
  assign n22114 = n8413 & n22113 ;
  assign n22115 = n1354 & n22114 ;
  assign n22116 = n1358 & n22115 ;
  assign n22117 = \pi0038  & ~n22116 ;
  assign n22118 = ~n22112 & n22117 ;
  assign n22119 = ~\pi0738  & ~n21763 ;
  assign n22120 = ~n22118 & n22119 ;
  assign n22121 = ~n22111 & n22120 ;
  assign n22122 = \pi0625  & n22121 ;
  assign n22123 = n1638 & n21765 ;
  assign n22124 = \pi0038  & ~n22123 ;
  assign n22125 = ~\pi0140  & \pi0738  ;
  assign n22126 = n22124 & n22125 ;
  assign n22127 = n21770 & n22125 ;
  assign n22128 = ~n21734 & n22127 ;
  assign n22129 = ~n22126 & ~n22128 ;
  assign n22130 = n6861 & n22129 ;
  assign n22131 = \pi0625  & ~n21763 ;
  assign n22132 = ~n22130 & n22131 ;
  assign n22133 = ~n22122 & ~n22132 ;
  assign n22134 = n21875 & n22133 ;
  assign n22135 = ~\pi0140  & \pi0625  ;
  assign n22136 = n21768 & n22135 ;
  assign n22137 = n21770 & n22135 ;
  assign n22138 = ~n21734 & n22137 ;
  assign n22139 = ~n22136 & ~n22138 ;
  assign n22140 = ~\pi1153  & n22139 ;
  assign n22141 = ~\pi0625  & n22121 ;
  assign n22142 = ~\pi0625  & ~n21763 ;
  assign n22143 = ~n22130 & n22142 ;
  assign n22144 = ~n22141 & ~n22143 ;
  assign n22145 = n22140 & n22144 ;
  assign n22146 = ~n22134 & ~n22145 ;
  assign n22147 = \pi0785  & ~n20866 ;
  assign n22148 = \pi0778  & ~n22147 ;
  assign n22149 = ~n22146 & n22148 ;
  assign n22150 = ~n21763 & ~n22130 ;
  assign n22151 = ~\pi0778  & ~n22147 ;
  assign n22152 = ~n22121 & n22151 ;
  assign n22153 = ~n22150 & n22152 ;
  assign n22154 = n21773 & n22147 ;
  assign n22155 = \pi0781  & n20871 ;
  assign n22156 = ~n22154 & ~n22155 ;
  assign n22157 = ~n22153 & n22156 ;
  assign n22158 = ~n22149 & n22157 ;
  assign n22159 = ~n21773 & n22155 ;
  assign n22160 = \pi0789  & ~n20876 ;
  assign n22161 = \pi0788  & ~n20883 ;
  assign n22162 = ~n22160 & ~n22161 ;
  assign n22163 = ~n22159 & n22162 ;
  assign n22164 = ~n22158 & n22163 ;
  assign n22165 = n21773 & ~n22162 ;
  assign n22166 = ~\pi0628  & \pi0629  ;
  assign n22167 = ~n22165 & n22166 ;
  assign n22168 = ~n22164 & n22167 ;
  assign n22169 = ~n21869 & ~n22168 ;
  assign n22170 = n21862 & ~n22169 ;
  assign n22171 = \pi0738  & n21753 ;
  assign n22172 = \pi0738  & n21758 ;
  assign n22173 = ~n21757 & n22172 ;
  assign n22174 = ~n22171 & ~n22173 ;
  assign n22175 = ~\pi0038  & \pi0738  ;
  assign n22176 = n21746 & n22175 ;
  assign n22177 = n22174 & ~n22176 ;
  assign n22178 = ~n21763 & ~n22177 ;
  assign n22179 = ~\pi0140  & \pi0299  ;
  assign n22180 = \pi0680  & ~n21586 ;
  assign n22181 = n6709 & n21959 ;
  assign n22182 = ~n22180 & ~n22181 ;
  assign n22183 = ~n21399 & n21403 ;
  assign n22184 = n21516 & ~n22180 ;
  assign n22185 = ~n22183 & n22184 ;
  assign n22186 = ~n22182 & ~n22185 ;
  assign n22187 = ~n21285 & n21915 ;
  assign n22188 = n21959 & ~n22187 ;
  assign n22189 = ~n21370 & n22188 ;
  assign n22190 = ~n21515 & n22189 ;
  assign n22191 = ~n21521 & n22190 ;
  assign n22192 = n21516 & ~n22183 ;
  assign n22193 = ~\pi0603  & ~n6706 ;
  assign n22194 = n20854 & n22193 ;
  assign n22195 = ~n21285 & n22194 ;
  assign n22196 = n21959 & ~n22195 ;
  assign n22197 = n21370 & n22196 ;
  assign n22198 = ~n22181 & ~n22197 ;
  assign n22199 = ~n22192 & ~n22198 ;
  assign n22200 = ~n22191 & ~n22199 ;
  assign n22201 = n22186 & ~n22200 ;
  assign n22202 = ~n6732 & n21954 ;
  assign n22203 = ~n22201 & n22202 ;
  assign n22204 = ~n21672 & ~n21972 ;
  assign n22205 = ~n21528 & ~n21977 ;
  assign n22206 = n6732 & ~n22205 ;
  assign n22207 = n22204 & n22206 ;
  assign n22208 = \pi0215  & ~n22207 ;
  assign n22209 = ~\pi0642  & ~n6706 ;
  assign n22210 = n21959 & n22209 ;
  assign n22211 = ~\pi0642  & n6706 ;
  assign n22212 = ~n21876 & n22211 ;
  assign n22213 = ~n22210 & ~n22212 ;
  assign n22214 = ~n21528 & ~n22213 ;
  assign n22215 = ~\pi0614  & n22196 ;
  assign n22216 = ~n22192 & n22215 ;
  assign n22217 = n22214 & n22216 ;
  assign n22218 = ~n20784 & ~n20854 ;
  assign n22219 = ~n21285 & ~n22218 ;
  assign n22220 = ~\pi0614  & \pi0642  ;
  assign n22221 = ~n22219 & n22220 ;
  assign n22222 = ~n6711 & ~n22219 ;
  assign n22223 = ~n22221 & ~n22222 ;
  assign n22224 = ~n22217 & n22223 ;
  assign n22225 = \pi0616  & ~n22218 ;
  assign n22226 = ~n21285 & n22225 ;
  assign n22227 = n22180 & ~n22226 ;
  assign n22228 = \pi0215  & n22227 ;
  assign n22229 = ~n22224 & n22228 ;
  assign n22230 = ~n22208 & ~n22229 ;
  assign n22231 = ~n22203 & ~n22230 ;
  assign n22232 = ~n20784 & n20855 ;
  assign n22233 = n2352 & ~n22232 ;
  assign n22234 = ~n21285 & n22233 ;
  assign n22235 = ~\pi0215  & ~n22234 ;
  assign n22236 = ~n22231 & ~n22235 ;
  assign n22237 = ~n21881 & n22193 ;
  assign n22238 = ~\pi0603  & n6706 ;
  assign n22239 = ~n21876 & n22238 ;
  assign n22240 = ~\pi0603  & ~n22239 ;
  assign n22241 = \pi0603  & ~\pi0665  ;
  assign n22242 = n20783 & n22241 ;
  assign n22243 = ~n22239 & ~n22242 ;
  assign n22244 = ~n21359 & n22243 ;
  assign n22245 = ~n22240 & ~n22244 ;
  assign n22246 = ~n22237 & ~n22245 ;
  assign n22247 = n6709 & ~n22246 ;
  assign n22248 = n6732 & n22247 ;
  assign n22249 = ~\pi0680  & n6732 ;
  assign n22250 = n21580 & n22249 ;
  assign n22251 = ~n22248 & ~n22250 ;
  assign n22252 = ~\pi0642  & ~n22218 ;
  assign n22253 = ~n22219 & ~n22252 ;
  assign n22254 = ~n21371 & ~n22253 ;
  assign n22255 = ~n21359 & n22254 ;
  assign n22256 = ~\pi0603  & ~n21371 ;
  assign n22257 = ~n22253 & n22256 ;
  assign n22258 = ~n22255 & ~n22257 ;
  assign n22259 = \pi0642  & ~n22218 ;
  assign n22260 = ~n21285 & n22259 ;
  assign n22261 = n6711 & ~n22260 ;
  assign n22262 = n22258 & n22261 ;
  assign n22263 = \pi0616  & ~n22219 ;
  assign n22264 = \pi0614  & ~\pi0616  ;
  assign n22265 = ~n22219 & n22264 ;
  assign n22266 = ~n22263 & ~n22265 ;
  assign n22267 = ~n22262 & n22266 ;
  assign n22268 = n6732 & n22180 ;
  assign n22269 = ~n22267 & n22268 ;
  assign n22270 = n22251 & ~n22269 ;
  assign n22271 = ~\pi0680  & n21905 ;
  assign n22272 = ~\pi0680  & n21908 ;
  assign n22273 = n21328 & n22272 ;
  assign n22274 = ~n22271 & ~n22273 ;
  assign n22275 = \pi0603  & ~\pi0621  ;
  assign n22276 = n20854 & ~n22275 ;
  assign n22277 = ~n21290 & n22276 ;
  assign n22278 = ~n21325 & n22277 ;
  assign n22279 = n6709 & ~n22278 ;
  assign n22280 = \pi0603  & ~n21346 ;
  assign n22281 = n22279 & ~n22280 ;
  assign n22282 = n22274 & ~n22281 ;
  assign n22283 = ~n21905 & ~n22218 ;
  assign n22284 = ~n22039 & n22283 ;
  assign n22285 = n22180 & ~n22284 ;
  assign n22286 = ~n2352 & ~n22285 ;
  assign n22287 = n22282 & n22286 ;
  assign n22288 = ~n21446 & ~n22287 ;
  assign n22289 = ~n22231 & ~n22288 ;
  assign n22290 = n22270 & n22289 ;
  assign n22291 = ~n22236 & ~n22290 ;
  assign n22292 = n22179 & ~n22291 ;
  assign n22293 = ~n21306 & ~n22022 ;
  assign n22294 = n6709 & ~n22293 ;
  assign n22295 = ~\pi0665  & n20783 ;
  assign n22296 = ~n21290 & n22295 ;
  assign n22297 = ~n21325 & n22296 ;
  assign n22298 = \pi0603  & ~n22297 ;
  assign n22299 = n21586 & ~n22298 ;
  assign n22300 = n22294 & n22299 ;
  assign n22301 = ~\pi0603  & n22025 ;
  assign n22302 = ~n21337 & ~n22301 ;
  assign n22303 = n21369 & ~n22298 ;
  assign n22304 = n22302 & n22303 ;
  assign n22305 = ~n21369 & ~n22025 ;
  assign n22306 = n21341 & n22305 ;
  assign n22307 = ~\pi0616  & ~n22306 ;
  assign n22308 = ~n22304 & n22307 ;
  assign n22309 = n22294 & ~n22298 ;
  assign n22310 = ~n22180 & ~n22309 ;
  assign n22311 = n21341 & ~n22025 ;
  assign n22312 = \pi0616  & ~n22311 ;
  assign n22313 = ~n22310 & ~n22312 ;
  assign n22314 = ~n22308 & n22313 ;
  assign n22315 = ~n22300 & ~n22314 ;
  assign n22316 = ~\pi0223  & ~n2165 ;
  assign n22317 = ~n20784 & ~n20855 ;
  assign n22318 = ~\pi0223  & ~n22317 ;
  assign n22319 = ~n21285 & n22318 ;
  assign n22320 = ~n22316 & ~n22319 ;
  assign n22321 = ~n6761 & ~n21561 ;
  assign n22322 = ~n22320 & n22321 ;
  assign n22323 = ~n22315 & n22322 ;
  assign n22324 = n6709 & ~n21359 ;
  assign n22325 = ~n22246 & n22324 ;
  assign n22326 = ~\pi0616  & n22180 ;
  assign n22327 = n22180 & n22218 ;
  assign n22328 = ~n21285 & n22327 ;
  assign n22329 = ~n22326 & ~n22328 ;
  assign n22330 = \pi0603  & \pi0665  ;
  assign n22331 = ~n20854 & ~n22330 ;
  assign n22332 = ~n21285 & n22331 ;
  assign n22333 = ~n22241 & ~n22332 ;
  assign n22334 = ~n21362 & n21369 ;
  assign n22335 = ~n22333 & n22334 ;
  assign n22336 = ~n21364 & n22335 ;
  assign n22337 = ~n20854 & ~n21369 ;
  assign n22338 = ~n20784 & n22337 ;
  assign n22339 = ~n21285 & n22338 ;
  assign n22340 = ~\pi0616  & ~n22339 ;
  assign n22341 = ~n22336 & n22340 ;
  assign n22342 = ~n22329 & ~n22341 ;
  assign n22343 = ~n2165 & ~n22342 ;
  assign n22344 = ~n22325 & n22343 ;
  assign n22345 = ~n21275 & ~n22344 ;
  assign n22346 = ~n21561 & ~n22320 ;
  assign n22347 = n22345 & n22346 ;
  assign n22348 = ~n20854 & n21370 ;
  assign n22349 = ~n21371 & n22348 ;
  assign n22350 = n21392 & n22349 ;
  assign n22351 = ~n20854 & n21375 ;
  assign n22352 = ~n21285 & n22351 ;
  assign n22353 = ~\pi0616  & ~n22352 ;
  assign n22354 = ~n22350 & n22353 ;
  assign n22355 = ~n22329 & ~n22354 ;
  assign n22356 = n21392 & ~n22333 ;
  assign n22357 = n21407 & n22356 ;
  assign n22358 = n6761 & ~n22357 ;
  assign n22359 = ~n22355 & n22358 ;
  assign n22360 = n21419 & ~n22333 ;
  assign n22361 = n6706 & ~n22333 ;
  assign n22362 = ~n21425 & n22361 ;
  assign n22363 = ~n22360 & ~n22362 ;
  assign n22364 = ~n21403 & n22232 ;
  assign n22365 = ~n21393 & n22232 ;
  assign n22366 = n21398 & n22365 ;
  assign n22367 = ~n22364 & ~n22366 ;
  assign n22368 = ~n22180 & n22367 ;
  assign n22369 = n21370 & ~n21392 ;
  assign n22370 = ~n22368 & ~n22369 ;
  assign n22371 = ~n22363 & n22370 ;
  assign n22372 = n21586 & ~n22367 ;
  assign n22373 = ~n6761 & ~n22372 ;
  assign n22374 = ~n22371 & n22373 ;
  assign n22375 = \pi0223  & ~n22374 ;
  assign n22376 = ~n22359 & n22375 ;
  assign n22377 = ~\pi0299  & ~n22376 ;
  assign n22378 = ~n22347 & n22377 ;
  assign n22379 = ~n22323 & n22378 ;
  assign n22380 = \pi0140  & n22379 ;
  assign n22381 = \pi0761  & ~n22380 ;
  assign n22382 = ~\pi0140  & ~\pi0299  ;
  assign n22383 = ~n22224 & n22227 ;
  assign n22384 = n6761 & ~n22205 ;
  assign n22385 = n22204 & n22384 ;
  assign n22386 = ~n22383 & n22385 ;
  assign n22387 = ~n6761 & n21954 ;
  assign n22388 = ~n22201 & n22387 ;
  assign n22389 = \pi0223  & ~n22388 ;
  assign n22390 = ~n22386 & n22389 ;
  assign n22391 = n2165 & ~n22232 ;
  assign n22392 = ~n21285 & n22391 ;
  assign n22393 = ~\pi0223  & ~n22392 ;
  assign n22394 = ~n22390 & ~n22393 ;
  assign n22395 = n6761 & n22247 ;
  assign n22396 = ~\pi0680  & n6761 ;
  assign n22397 = n21580 & n22396 ;
  assign n22398 = ~n22395 & ~n22397 ;
  assign n22399 = n6761 & n22180 ;
  assign n22400 = ~n22267 & n22399 ;
  assign n22401 = n22398 & ~n22400 ;
  assign n22402 = ~n2165 & ~n22285 ;
  assign n22403 = n22282 & n22402 ;
  assign n22404 = ~n21368 & ~n22403 ;
  assign n22405 = ~n22390 & ~n22404 ;
  assign n22406 = n22401 & n22405 ;
  assign n22407 = ~n22394 & ~n22406 ;
  assign n22408 = n22382 & ~n22407 ;
  assign n22409 = \pi0140  & \pi0299  ;
  assign n22410 = n6732 & ~n22342 ;
  assign n22411 = ~n22325 & n22410 ;
  assign n22412 = ~n2352 & ~n22411 ;
  assign n22413 = ~n20784 & n22049 ;
  assign n22414 = ~n21285 & n22413 ;
  assign n22415 = ~\pi0215  & ~n22414 ;
  assign n22416 = ~n22412 & n22415 ;
  assign n22417 = ~\pi0215  & ~n6732 ;
  assign n22418 = ~n22414 & n22417 ;
  assign n22419 = ~n22300 & n22418 ;
  assign n22420 = ~n22314 & n22419 ;
  assign n22421 = ~n22416 & ~n22420 ;
  assign n22422 = n6732 & n22357 ;
  assign n22423 = n6732 & ~n22329 ;
  assign n22424 = ~n22354 & n22423 ;
  assign n22425 = ~n22422 & ~n22424 ;
  assign n22426 = \pi0215  & n6732 ;
  assign n22427 = \pi0215  & ~n22372 ;
  assign n22428 = ~n22371 & n22427 ;
  assign n22429 = ~n22426 & ~n22428 ;
  assign n22430 = n22425 & ~n22429 ;
  assign n22431 = n22421 & ~n22430 ;
  assign n22432 = n22409 & ~n22431 ;
  assign n22433 = ~n22408 & ~n22432 ;
  assign n22434 = n22381 & n22433 ;
  assign n22435 = ~n22292 & n22434 ;
  assign n22436 = ~n21370 & ~n22276 ;
  assign n22437 = ~n21285 & n22436 ;
  assign n22438 = n22180 & ~n22437 ;
  assign n22439 = n21370 & n21528 ;
  assign n22440 = n21370 & n22023 ;
  assign n22441 = ~n22053 & n22440 ;
  assign n22442 = ~n22439 & ~n22441 ;
  assign n22443 = n22438 & n22442 ;
  assign n22444 = ~n21405 & n22052 ;
  assign n22445 = ~n22180 & ~n22444 ;
  assign n22446 = ~n21528 & n22445 ;
  assign n22447 = ~n21527 & n22446 ;
  assign n22448 = ~n22443 & ~n22447 ;
  assign n22449 = ~\pi0299  & n6761 ;
  assign n22450 = ~n22448 & n22449 ;
  assign n22451 = n22320 & n22450 ;
  assign n22452 = n22023 & ~n22053 ;
  assign n22453 = ~n6706 & ~n20854 ;
  assign n22454 = ~n21285 & n22453 ;
  assign n22455 = ~n21520 & n22023 ;
  assign n22456 = ~n22454 & ~n22455 ;
  assign n22457 = n22452 & ~n22456 ;
  assign n22458 = ~n22445 & n22457 ;
  assign n22459 = ~n6761 & ~n21516 ;
  assign n22460 = ~n6761 & n21403 ;
  assign n22461 = ~n21399 & n22460 ;
  assign n22462 = ~n22459 & ~n22461 ;
  assign n22463 = ~n21527 & ~n22462 ;
  assign n22464 = ~n22458 & n22463 ;
  assign n22465 = \pi0223  & ~n22464 ;
  assign n22466 = ~\pi0299  & n22320 ;
  assign n22467 = ~n22465 & n22466 ;
  assign n22468 = ~n22451 & ~n22467 ;
  assign n22469 = \pi0140  & ~n22468 ;
  assign n22470 = ~\pi0299  & ~n22465 ;
  assign n22471 = ~n22450 & ~n22470 ;
  assign n22472 = ~\pi0680  & ~n21491 ;
  assign n22473 = ~n21489 & n22472 ;
  assign n22474 = n6761 & ~n22473 ;
  assign n22475 = ~n21362 & n21370 ;
  assign n22476 = ~n22333 & n22475 ;
  assign n22477 = ~n21364 & n22476 ;
  assign n22478 = ~n21489 & ~n22477 ;
  assign n22479 = n22438 & n22478 ;
  assign n22480 = n6709 & n21359 ;
  assign n22481 = n6709 & ~n20784 ;
  assign n22482 = n22025 & n22481 ;
  assign n22483 = ~n22480 & ~n22482 ;
  assign n22484 = ~n22479 & n22483 ;
  assign n22485 = n22474 & n22484 ;
  assign n22486 = ~n2165 & ~n22485 ;
  assign n22487 = ~n22471 & n22486 ;
  assign n22488 = n21375 & ~n22023 ;
  assign n22489 = ~n21306 & n22488 ;
  assign n22490 = ~n22022 & n22489 ;
  assign n22491 = ~n21286 & ~n21370 ;
  assign n22492 = n21328 & n22491 ;
  assign n22493 = ~n22490 & ~n22492 ;
  assign n22494 = n22180 & ~n22493 ;
  assign n22495 = \pi0603  & n21370 ;
  assign n22496 = ~n22297 & n22495 ;
  assign n22497 = ~\pi0603  & n22180 ;
  assign n22498 = ~n21306 & n22180 ;
  assign n22499 = ~n21345 & n22498 ;
  assign n22500 = ~n22497 & ~n22499 ;
  assign n22501 = n22496 & ~n22500 ;
  assign n22502 = n21370 & ~n22500 ;
  assign n22503 = ~n22302 & n22502 ;
  assign n22504 = ~n22501 & ~n22503 ;
  assign n22505 = ~n22494 & n22504 ;
  assign n22506 = ~n22180 & ~n22294 ;
  assign n22507 = n21499 & n22506 ;
  assign n22508 = ~n6761 & ~n22507 ;
  assign n22509 = n22505 & n22508 ;
  assign n22510 = \pi0140  & ~n22509 ;
  assign n22511 = n22487 & n22510 ;
  assign n22512 = ~n22469 & ~n22511 ;
  assign n22513 = n2352 & ~n22317 ;
  assign n22514 = ~n21285 & n22513 ;
  assign n22515 = ~\pi0215  & ~n22514 ;
  assign n22516 = n2352 & n22515 ;
  assign n22517 = ~n6732 & ~n22507 ;
  assign n22518 = n22505 & n22517 ;
  assign n22519 = n6732 & ~n22473 ;
  assign n22520 = n22484 & n22519 ;
  assign n22521 = n22515 & ~n22520 ;
  assign n22522 = ~n22518 & n22521 ;
  assign n22523 = ~n22516 & ~n22522 ;
  assign n22524 = ~n21527 & ~n22192 ;
  assign n22525 = ~n22458 & n22524 ;
  assign n22526 = \pi0215  & ~n6732 ;
  assign n22527 = n22525 & n22526 ;
  assign n22528 = n22426 & ~n22448 ;
  assign n22529 = ~n22527 & ~n22528 ;
  assign n22530 = n22523 & n22529 ;
  assign n22531 = n22409 & ~n22530 ;
  assign n22532 = ~\pi0120  & ~n21301 ;
  assign n22533 = n1689 & n22317 ;
  assign n22534 = n1259 & n22533 ;
  assign n22535 = n1249 & n22534 ;
  assign n22536 = n1281 & n22535 ;
  assign n22537 = n2165 & n22536 ;
  assign n22538 = ~n22532 & n22537 ;
  assign n22539 = ~\pi0223  & ~n22538 ;
  assign n22540 = ~\pi0680  & n21428 ;
  assign n22541 = n21372 & ~n22188 ;
  assign n22542 = n21392 & n22541 ;
  assign n22543 = n21376 & ~n22188 ;
  assign n22544 = n22180 & ~n22543 ;
  assign n22545 = ~n22542 & n22544 ;
  assign n22546 = n6709 & n22275 ;
  assign n22547 = \pi0680  & n6709 ;
  assign n22548 = n21959 & n22547 ;
  assign n22549 = ~n22546 & ~n22548 ;
  assign n22550 = ~n6761 & n22549 ;
  assign n22551 = ~n22545 & n22550 ;
  assign n22552 = ~n22540 & n22551 ;
  assign n22553 = n6761 & ~n20855 ;
  assign n22554 = n21413 & n22553 ;
  assign n22555 = n21410 & n22553 ;
  assign n22556 = n21392 & n22555 ;
  assign n22557 = ~n22554 & ~n22556 ;
  assign n22558 = n6709 & ~n22275 ;
  assign n22559 = ~n6706 & n22558 ;
  assign n22560 = n20854 & n22558 ;
  assign n22561 = ~n21285 & n22560 ;
  assign n22562 = ~n22559 & ~n22561 ;
  assign n22563 = ~n21962 & ~n22562 ;
  assign n22564 = n6761 & n22563 ;
  assign n22565 = \pi0223  & ~n22564 ;
  assign n22566 = n22557 & n22565 ;
  assign n22567 = ~n22552 & n22566 ;
  assign n22568 = ~n22539 & ~n22567 ;
  assign n22569 = ~\pi0680  & ~n21376 ;
  assign n22570 = ~n21374 & n22569 ;
  assign n22571 = ~n6706 & n22276 ;
  assign n22572 = n20854 & n22276 ;
  assign n22573 = ~n21285 & n22572 ;
  assign n22574 = ~n22571 & ~n22573 ;
  assign n22575 = n6709 & n22574 ;
  assign n22576 = ~n21881 & n21973 ;
  assign n22577 = ~n22575 & ~n22576 ;
  assign n22578 = ~n22570 & n22577 ;
  assign n22579 = n20854 & n21372 ;
  assign n22580 = ~n21362 & n22579 ;
  assign n22581 = ~n21364 & n22580 ;
  assign n22582 = ~n21370 & n22276 ;
  assign n22583 = ~n21285 & n22582 ;
  assign n22584 = n22180 & ~n22583 ;
  assign n22585 = ~n22581 & n22584 ;
  assign n22586 = n6761 & ~n22585 ;
  assign n22587 = n22578 & n22586 ;
  assign n22588 = ~n20784 & ~n21905 ;
  assign n22589 = ~n22039 & n22588 ;
  assign n22590 = ~\pi0680  & ~n22589 ;
  assign n22591 = n22180 & ~n22276 ;
  assign n22592 = ~n21917 & n22180 ;
  assign n22593 = ~n21914 & n22592 ;
  assign n22594 = ~n22591 & ~n22593 ;
  assign n22595 = ~n6761 & ~n22279 ;
  assign n22596 = n22594 & n22595 ;
  assign n22597 = ~n22590 & n22596 ;
  assign n22598 = ~n22587 & ~n22597 ;
  assign n22599 = ~n2165 & ~n22567 ;
  assign n22600 = ~n22598 & n22599 ;
  assign n22601 = ~n22568 & ~n22600 ;
  assign n22602 = n22382 & ~n22601 ;
  assign n22603 = n1281 & n2352 ;
  assign n22604 = n22535 & n22603 ;
  assign n22605 = ~\pi0215  & ~n22604 ;
  assign n22606 = ~\pi0120  & ~\pi0215  ;
  assign n22607 = ~n21301 & n22606 ;
  assign n22608 = ~n22605 & ~n22607 ;
  assign n22609 = ~n6732 & n22549 ;
  assign n22610 = ~n22545 & n22609 ;
  assign n22611 = ~n22540 & n22610 ;
  assign n22612 = n6732 & ~n20855 ;
  assign n22613 = n21413 & n22612 ;
  assign n22614 = n21410 & n22612 ;
  assign n22615 = n21392 & n22614 ;
  assign n22616 = ~n22613 & ~n22615 ;
  assign n22617 = n6732 & n22563 ;
  assign n22618 = \pi0215  & ~n22617 ;
  assign n22619 = n22616 & n22618 ;
  assign n22620 = ~n22611 & n22619 ;
  assign n22621 = n22608 & ~n22620 ;
  assign n22622 = n6732 & ~n22585 ;
  assign n22623 = n22578 & n22622 ;
  assign n22624 = ~n6732 & ~n22279 ;
  assign n22625 = n22594 & n22624 ;
  assign n22626 = ~n22590 & n22625 ;
  assign n22627 = ~n22623 & ~n22626 ;
  assign n22628 = ~n2352 & ~n22620 ;
  assign n22629 = ~n22627 & n22628 ;
  assign n22630 = ~n22621 & ~n22629 ;
  assign n22631 = n22179 & ~n22630 ;
  assign n22632 = ~\pi0761  & ~n22631 ;
  assign n22633 = ~n22602 & n22632 ;
  assign n22634 = ~n22531 & n22633 ;
  assign n22635 = n22512 & n22634 ;
  assign n22636 = ~\pi0038  & ~n22635 ;
  assign n22637 = ~n22435 & n22636 ;
  assign n22638 = ~n1288 & ~n22637 ;
  assign n22639 = ~\pi0299  & \pi0680  ;
  assign n22640 = n21481 & n22639 ;
  assign n22641 = n21477 & n22639 ;
  assign n22642 = ~n21263 & n22641 ;
  assign n22643 = ~n22640 & ~n22642 ;
  assign n22644 = \pi0299  & \pi0680  ;
  assign n22645 = n21474 & n22644 ;
  assign n22646 = ~n21472 & n22645 ;
  assign n22647 = \pi0299  & ~n22646 ;
  assign n22648 = ~n22006 & n22647 ;
  assign n22649 = n22011 & ~n22013 ;
  assign n22650 = ~\pi0299  & ~n22646 ;
  assign n22651 = ~n22649 & n22650 ;
  assign n22652 = ~n22648 & ~n22651 ;
  assign n22653 = n22643 & ~n22652 ;
  assign n22654 = ~\pi0140  & ~n22653 ;
  assign n22655 = ~\pi0210  & ~\pi0603  ;
  assign n22656 = n21203 & n22655 ;
  assign n22657 = ~n22096 & n22656 ;
  assign n22658 = \pi0210  & ~\pi0603  ;
  assign n22659 = n21236 & n22658 ;
  assign n22660 = n22094 & n22659 ;
  assign n22661 = ~n22657 & ~n22660 ;
  assign n22662 = \pi0680  & ~n22330 ;
  assign n22663 = ~n21243 & n22662 ;
  assign n22664 = ~n21249 & n22663 ;
  assign n22665 = n22661 & n22664 ;
  assign n22666 = n22409 & ~n22665 ;
  assign n22667 = \pi0603  & n21266 ;
  assign n22668 = n21247 & n21477 ;
  assign n22669 = ~n22667 & ~n22668 ;
  assign n22670 = n21236 & n21258 ;
  assign n22671 = n22094 & n22670 ;
  assign n22672 = n21203 & n21256 ;
  assign n22673 = ~n22096 & n22672 ;
  assign n22674 = n22662 & ~n22673 ;
  assign n22675 = ~n22671 & n22674 ;
  assign n22676 = n22669 & n22675 ;
  assign n22677 = n18434 & ~n22676 ;
  assign n22678 = ~n22666 & ~n22677 ;
  assign n22679 = \pi0761  & n22678 ;
  assign n22680 = ~n22654 & n22679 ;
  assign n22681 = ~\pi0299  & ~n22649 ;
  assign n22682 = ~n22007 & ~n22681 ;
  assign n22683 = n21272 & n22682 ;
  assign n22684 = ~\pi0140  & ~\pi0761  ;
  assign n22685 = ~n22683 & n22684 ;
  assign n22686 = ~n22101 & n22103 ;
  assign n22687 = ~\pi0299  & ~n22686 ;
  assign n22688 = ~n22100 & ~n22687 ;
  assign n22689 = ~\pi0299  & ~n21481 ;
  assign n22690 = ~n21478 & n22689 ;
  assign n22691 = \pi0299  & ~n21475 ;
  assign n22692 = ~n22690 & ~n22691 ;
  assign n22693 = ~n22688 & ~n22692 ;
  assign n22694 = n21485 & ~n22693 ;
  assign n22695 = ~n22685 & ~n22694 ;
  assign n22696 = ~n22680 & n22695 ;
  assign n22697 = ~\pi0039  & ~n22696 ;
  assign n22698 = n1287 & n1289 ;
  assign n22699 = ~n22697 & n22698 ;
  assign n22700 = ~n22638 & n22699 ;
  assign n22701 = \pi0738  & n6861 ;
  assign n22702 = \pi0038  & ~n22112 ;
  assign n22703 = \pi0603  & \pi0761  ;
  assign n22704 = ~n20783 & n22703 ;
  assign n22705 = n8413 & ~n22317 ;
  assign n22706 = n1354 & n1689 ;
  assign n22707 = n22705 & n22706 ;
  assign n22708 = n1358 & n22707 ;
  assign n22709 = ~n22704 & n22708 ;
  assign n22710 = n6861 & ~n22709 ;
  assign n22711 = n22702 & n22710 ;
  assign n22712 = ~n22701 & ~n22711 ;
  assign n22713 = ~n21763 & n22712 ;
  assign n22714 = ~n22700 & n22713 ;
  assign n22715 = ~n22178 & ~n22714 ;
  assign n22716 = ~\pi0778  & n22715 ;
  assign n22717 = \pi0609  & ~n22716 ;
  assign n22718 = ~\pi0778  & ~n22121 ;
  assign n22719 = ~n22150 & n22718 ;
  assign n22720 = ~\pi0609  & ~n22719 ;
  assign n22721 = \pi1155  & ~n22720 ;
  assign n22722 = \pi0778  & \pi1155  ;
  assign n22723 = ~n22146 & n22722 ;
  assign n22724 = ~n22721 & ~n22723 ;
  assign n22725 = ~n22717 & ~n22724 ;
  assign n22726 = \pi0625  & n1289 ;
  assign n22727 = n1287 & n22726 ;
  assign n22728 = ~n22135 & ~n22727 ;
  assign n22729 = ~n22177 & ~n22728 ;
  assign n22730 = n22712 & ~n22728 ;
  assign n22731 = ~n22700 & n22730 ;
  assign n22732 = ~n22729 & ~n22731 ;
  assign n22733 = ~\pi0625  & n1289 ;
  assign n22734 = n1287 & n22733 ;
  assign n22735 = ~n21870 & ~n22734 ;
  assign n22736 = ~n21762 & ~n22735 ;
  assign n22737 = \pi1153  & ~n22736 ;
  assign n22738 = n22732 & n22737 ;
  assign n22739 = \pi0608  & ~n22140 ;
  assign n22740 = \pi0608  & ~\pi0625  ;
  assign n22741 = n22121 & n22740 ;
  assign n22742 = ~n21763 & n22740 ;
  assign n22743 = ~n22130 & n22742 ;
  assign n22744 = ~n22741 & ~n22743 ;
  assign n22745 = ~n22739 & n22744 ;
  assign n22746 = ~n22738 & ~n22745 ;
  assign n22747 = ~n22177 & ~n22735 ;
  assign n22748 = n22712 & ~n22735 ;
  assign n22749 = ~n22700 & n22748 ;
  assign n22750 = ~n22747 & ~n22749 ;
  assign n22751 = ~n21762 & ~n22728 ;
  assign n22752 = ~\pi1153  & ~n22751 ;
  assign n22753 = n22750 & n22752 ;
  assign n22754 = ~\pi0608  & ~n21875 ;
  assign n22755 = ~\pi0608  & \pi0625  ;
  assign n22756 = n22121 & n22755 ;
  assign n22757 = ~n21763 & n22755 ;
  assign n22758 = ~n22130 & n22757 ;
  assign n22759 = ~n22756 & ~n22758 ;
  assign n22760 = ~n22754 & n22759 ;
  assign n22761 = ~n22753 & ~n22760 ;
  assign n22762 = ~n22746 & ~n22761 ;
  assign n22763 = \pi0778  & ~n22724 ;
  assign n22764 = n22762 & n22763 ;
  assign n22765 = ~n22725 & ~n22764 ;
  assign n22766 = \pi0660  & \pi1155  ;
  assign n22767 = ~\pi0609  & ~n20985 ;
  assign n22768 = n21773 & ~n22767 ;
  assign n22769 = \pi0660  & ~n22768 ;
  assign n22770 = ~n22767 & n22769 ;
  assign n22771 = ~n21763 & n22769 ;
  assign n22772 = ~n21762 & n22771 ;
  assign n22773 = ~n22770 & ~n22772 ;
  assign n22774 = ~n22766 & n22773 ;
  assign n22775 = n22765 & ~n22774 ;
  assign n22776 = ~\pi0618  & \pi0785  ;
  assign n22777 = n22775 & n22776 ;
  assign n22778 = ~\pi0609  & ~n22716 ;
  assign n22779 = \pi0778  & ~n22146 ;
  assign n22780 = \pi0609  & ~n22719 ;
  assign n22781 = ~n22779 & n22780 ;
  assign n22782 = ~n22778 & ~n22781 ;
  assign n22783 = \pi0778  & ~n22781 ;
  assign n22784 = n22762 & n22783 ;
  assign n22785 = ~n22782 & ~n22784 ;
  assign n22786 = ~\pi1155  & ~n22785 ;
  assign n22787 = ~\pi0660  & ~\pi1155  ;
  assign n22788 = \pi0609  & ~n20985 ;
  assign n22789 = n21773 & ~n22788 ;
  assign n22790 = ~\pi0660  & ~n22789 ;
  assign n22791 = ~n22788 & n22790 ;
  assign n22792 = ~n21763 & n22790 ;
  assign n22793 = ~n21762 & n22792 ;
  assign n22794 = ~n22791 & ~n22793 ;
  assign n22795 = ~n22787 & n22794 ;
  assign n22796 = n22776 & ~n22795 ;
  assign n22797 = ~n22786 & n22796 ;
  assign n22798 = ~n22777 & ~n22797 ;
  assign n22799 = \pi0778  & n22762 ;
  assign n22800 = ~\pi0785  & ~n22716 ;
  assign n22801 = ~\pi0618  & n22800 ;
  assign n22802 = ~n22799 & n22801 ;
  assign n22803 = \pi0618  & ~n22154 ;
  assign n22804 = ~n22153 & n22803 ;
  assign n22805 = ~n22149 & n22804 ;
  assign n22806 = ~\pi1154  & ~n22805 ;
  assign n22807 = ~n22802 & n22806 ;
  assign n22808 = n22798 & n22807 ;
  assign n22809 = ~\pi0627  & ~n21790 ;
  assign n22810 = \pi0618  & ~\pi0627  ;
  assign n22811 = ~n22809 & ~n22810 ;
  assign n22812 = ~n21781 & ~n22809 ;
  assign n22813 = ~n21780 & n22812 ;
  assign n22814 = ~n22811 & ~n22813 ;
  assign n22815 = ~n22808 & n22814 ;
  assign n22816 = \pi0618  & \pi0785  ;
  assign n22817 = n22775 & n22816 ;
  assign n22818 = ~n22795 & n22816 ;
  assign n22819 = ~n22786 & n22818 ;
  assign n22820 = ~n22817 & ~n22819 ;
  assign n22821 = \pi0618  & n22800 ;
  assign n22822 = ~n22799 & n22821 ;
  assign n22823 = ~\pi0618  & ~n22154 ;
  assign n22824 = ~n22153 & n22823 ;
  assign n22825 = ~n22149 & n22824 ;
  assign n22826 = \pi1154  & ~n22825 ;
  assign n22827 = ~n22822 & n22826 ;
  assign n22828 = n22820 & n22827 ;
  assign n22829 = \pi0627  & ~n21800 ;
  assign n22830 = ~\pi0618  & \pi0627  ;
  assign n22831 = ~n22829 & ~n22830 ;
  assign n22832 = ~n21781 & ~n22829 ;
  assign n22833 = ~n21780 & n22832 ;
  assign n22834 = ~n22831 & ~n22833 ;
  assign n22835 = ~n22828 & n22834 ;
  assign n22836 = ~n22815 & ~n22835 ;
  assign n22837 = n21806 & ~n22836 ;
  assign n22838 = ~\pi0781  & n22800 ;
  assign n22839 = ~n22799 & n22838 ;
  assign n22840 = ~\pi0781  & \pi0785  ;
  assign n22841 = n22775 & n22840 ;
  assign n22842 = ~n22795 & n22840 ;
  assign n22843 = ~n22786 & n22842 ;
  assign n22844 = ~n22841 & ~n22843 ;
  assign n22845 = ~n22839 & n22844 ;
  assign n22846 = ~\pi0789  & ~n22845 ;
  assign n22847 = \pi0626  & ~n22846 ;
  assign n22848 = ~n22837 & n22847 ;
  assign n22849 = ~n22155 & ~n22160 ;
  assign n22850 = n21773 & ~n22849 ;
  assign n22851 = ~\pi0626  & n22850 ;
  assign n22852 = ~n22153 & ~n22154 ;
  assign n22853 = ~n22149 & n22852 ;
  assign n22854 = ~\pi0626  & n22849 ;
  assign n22855 = ~n22853 & n22854 ;
  assign n22856 = ~n22851 & ~n22855 ;
  assign n22857 = \pi0641  & n22856 ;
  assign n22858 = ~n22848 & n22857 ;
  assign n22859 = \pi0619  & \pi0781  ;
  assign n22860 = ~n22836 & n22859 ;
  assign n22861 = \pi0619  & ~n22845 ;
  assign n22862 = \pi1159  & ~n22159 ;
  assign n22863 = ~n22158 & n22862 ;
  assign n22864 = ~n20830 & ~n22863 ;
  assign n22865 = ~n22861 & ~n22864 ;
  assign n22866 = ~n22860 & n22865 ;
  assign n22867 = \pi0648  & n21819 ;
  assign n22868 = ~n22866 & n22867 ;
  assign n22869 = ~\pi0619  & \pi0781  ;
  assign n22870 = ~n22836 & n22869 ;
  assign n22871 = ~\pi0619  & ~n22845 ;
  assign n22872 = ~\pi0619  & ~\pi1159  ;
  assign n22873 = ~\pi1159  & ~n22159 ;
  assign n22874 = ~n22158 & n22873 ;
  assign n22875 = ~n22872 & ~n22874 ;
  assign n22876 = ~n22871 & ~n22875 ;
  assign n22877 = ~n22870 & n22876 ;
  assign n22878 = ~\pi0648  & n21830 ;
  assign n22879 = ~n22877 & n22878 ;
  assign n22880 = ~n22868 & ~n22879 ;
  assign n22881 = \pi0789  & n22857 ;
  assign n22882 = ~n22880 & n22881 ;
  assign n22883 = ~n22858 & ~n22882 ;
  assign n22884 = \pi0641  & \pi1158  ;
  assign n22885 = n21858 & ~n22884 ;
  assign n22886 = n22883 & ~n22885 ;
  assign n22887 = \pi0788  & n22886 ;
  assign n22888 = ~\pi0626  & ~n22846 ;
  assign n22889 = ~n22837 & n22888 ;
  assign n22890 = \pi0626  & n22850 ;
  assign n22891 = \pi0626  & n22849 ;
  assign n22892 = ~n22853 & n22891 ;
  assign n22893 = ~n22890 & ~n22892 ;
  assign n22894 = ~n22889 & n22893 ;
  assign n22895 = \pi0789  & n22893 ;
  assign n22896 = ~n22880 & n22895 ;
  assign n22897 = ~n22894 & ~n22896 ;
  assign n22898 = ~\pi0641  & ~n22897 ;
  assign n22899 = ~\pi0641  & ~\pi1158  ;
  assign n22900 = n21847 & ~n22899 ;
  assign n22901 = \pi0788  & ~n22900 ;
  assign n22902 = ~n22898 & n22901 ;
  assign n22903 = ~n22887 & ~n22902 ;
  assign n22904 = ~\pi0788  & ~n22846 ;
  assign n22905 = ~n22837 & n22904 ;
  assign n22906 = \pi0628  & ~n22905 ;
  assign n22907 = \pi0628  & \pi0789  ;
  assign n22908 = ~n22880 & n22907 ;
  assign n22909 = ~n22906 & ~n22908 ;
  assign n22910 = ~n22169 & ~n22909 ;
  assign n22911 = n22903 & n22910 ;
  assign n22912 = ~n22170 & ~n22911 ;
  assign n22913 = ~\pi0647  & \pi0792  ;
  assign n22914 = ~n22912 & n22913 ;
  assign n22915 = ~\pi0628  & ~n22905 ;
  assign n22916 = ~\pi0628  & \pi0789  ;
  assign n22917 = ~n22880 & n22916 ;
  assign n22918 = ~n22915 & ~n22917 ;
  assign n22919 = n22903 & ~n22918 ;
  assign n22920 = \pi0788  & ~n21859 ;
  assign n22921 = \pi0628  & n21834 ;
  assign n22922 = ~n22920 & n22921 ;
  assign n22923 = ~\pi1156  & ~n22922 ;
  assign n22924 = ~n22919 & n22923 ;
  assign n22925 = ~\pi0140  & ~\pi0628  ;
  assign n22926 = n21768 & n22925 ;
  assign n22927 = n21770 & n22925 ;
  assign n22928 = ~n21734 & n22927 ;
  assign n22929 = ~n22926 & ~n22928 ;
  assign n22930 = \pi1156  & n22929 ;
  assign n22931 = ~\pi0629  & ~n22930 ;
  assign n22932 = \pi0628  & ~\pi0629  ;
  assign n22933 = ~n22165 & n22932 ;
  assign n22934 = ~n22164 & n22933 ;
  assign n22935 = ~n22931 & ~n22934 ;
  assign n22936 = n22913 & ~n22935 ;
  assign n22937 = ~n22924 & n22936 ;
  assign n22938 = ~n22914 & ~n22937 ;
  assign n22939 = ~\pi0792  & ~n22905 ;
  assign n22940 = \pi0789  & ~\pi0792  ;
  assign n22941 = ~n22880 & n22940 ;
  assign n22942 = ~n22939 & ~n22941 ;
  assign n22943 = ~\pi0647  & ~n22942 ;
  assign n22944 = n22903 & n22943 ;
  assign n22945 = ~\pi0647  & ~\pi1157  ;
  assign n22946 = ~n20846 & n21834 ;
  assign n22947 = n20846 & ~n21773 ;
  assign n22948 = ~\pi1157  & ~n22947 ;
  assign n22949 = ~n22946 & n22948 ;
  assign n22950 = \pi0788  & n22948 ;
  assign n22951 = ~n21859 & n22950 ;
  assign n22952 = ~n22949 & ~n22951 ;
  assign n22953 = ~n22945 & n22952 ;
  assign n22954 = ~n22944 & ~n22953 ;
  assign n22955 = n22938 & n22954 ;
  assign n22956 = \pi0647  & \pi0792  ;
  assign n22957 = \pi0647  & ~n22165 ;
  assign n22958 = ~n22164 & n22957 ;
  assign n22959 = ~n22956 & ~n22958 ;
  assign n22960 = ~\pi0140  & ~\pi0647  ;
  assign n22961 = n21768 & n22960 ;
  assign n22962 = n21770 & n22960 ;
  assign n22963 = ~n21734 & n22962 ;
  assign n22964 = ~n22961 & ~n22963 ;
  assign n22965 = \pi1157  & n22964 ;
  assign n22966 = n22959 & n22965 ;
  assign n22967 = \pi0628  & ~n22165 ;
  assign n22968 = ~n22164 & n22967 ;
  assign n22969 = n22930 & ~n22968 ;
  assign n22970 = ~\pi0628  & ~n22165 ;
  assign n22971 = ~n22164 & n22970 ;
  assign n22972 = n21868 & ~n22971 ;
  assign n22973 = ~n22969 & ~n22972 ;
  assign n22974 = \pi0792  & n22965 ;
  assign n22975 = ~n22973 & n22974 ;
  assign n22976 = ~n22966 & ~n22975 ;
  assign n22977 = ~\pi0630  & n22976 ;
  assign n22978 = ~n22955 & n22977 ;
  assign n22979 = ~n22912 & n22956 ;
  assign n22980 = ~n22935 & n22956 ;
  assign n22981 = ~n22924 & n22980 ;
  assign n22982 = ~n22979 & ~n22981 ;
  assign n22983 = \pi0647  & ~n22942 ;
  assign n22984 = n22903 & n22983 ;
  assign n22985 = \pi1157  & ~n22947 ;
  assign n22986 = ~n22946 & n22985 ;
  assign n22987 = \pi0788  & n22985 ;
  assign n22988 = ~n21859 & n22987 ;
  assign n22989 = ~n22986 & ~n22988 ;
  assign n22990 = ~n20925 & n22989 ;
  assign n22991 = ~n22984 & ~n22990 ;
  assign n22992 = n22982 & n22991 ;
  assign n22993 = ~\pi0647  & ~n22165 ;
  assign n22994 = ~n22164 & n22993 ;
  assign n22995 = ~n22913 & ~n22994 ;
  assign n22996 = n20898 & n21768 ;
  assign n22997 = n20898 & n21770 ;
  assign n22998 = ~n21734 & n22997 ;
  assign n22999 = ~n22996 & ~n22998 ;
  assign n23000 = ~\pi1157  & n22999 ;
  assign n23001 = n22995 & n23000 ;
  assign n23002 = \pi0792  & n23000 ;
  assign n23003 = ~n22973 & n23002 ;
  assign n23004 = ~n23001 & ~n23003 ;
  assign n23005 = \pi0630  & n23004 ;
  assign n23006 = ~n22992 & n23005 ;
  assign n23007 = ~n22978 & ~n23006 ;
  assign n23008 = \pi0787  & ~n23007 ;
  assign n23009 = ~\pi0787  & ~n22942 ;
  assign n23010 = n22903 & n23009 ;
  assign n23011 = ~\pi0787  & \pi0792  ;
  assign n23012 = ~n22912 & n23011 ;
  assign n23013 = ~n22935 & n23011 ;
  assign n23014 = ~n22924 & n23013 ;
  assign n23015 = ~n23012 & ~n23014 ;
  assign n23016 = ~n23010 & n23015 ;
  assign n23017 = ~\pi0790  & n23016 ;
  assign n23018 = ~n23008 & n23017 ;
  assign n23019 = n9948 & ~n23018 ;
  assign n23020 = ~n21133 & ~n23019 ;
  assign n23021 = ~\pi0644  & \pi0787  ;
  assign n23022 = ~n23007 & n23021 ;
  assign n23023 = ~\pi0644  & ~n23016 ;
  assign n23024 = n22976 & n23004 ;
  assign n23025 = \pi0787  & ~n23024 ;
  assign n23026 = ~n22164 & ~n22165 ;
  assign n23027 = ~\pi0792  & ~n23026 ;
  assign n23028 = ~\pi0787  & n23027 ;
  assign n23029 = ~n22973 & n23011 ;
  assign n23030 = ~n23028 & ~n23029 ;
  assign n23031 = \pi0644  & n23030 ;
  assign n23032 = ~n23025 & n23031 ;
  assign n23033 = ~\pi0715  & ~n23032 ;
  assign n23034 = ~n23023 & n23033 ;
  assign n23035 = ~n23022 & n23034 ;
  assign n23036 = ~n21088 & ~n22947 ;
  assign n23037 = ~n22946 & n23036 ;
  assign n23038 = \pi0788  & n23036 ;
  assign n23039 = ~n21859 & n23038 ;
  assign n23040 = ~n23037 & ~n23039 ;
  assign n23041 = n21088 & n21773 ;
  assign n23042 = ~\pi0644  & ~n23041 ;
  assign n23043 = n23040 & n23042 ;
  assign n23044 = n21096 & n21768 ;
  assign n23045 = n21096 & n21770 ;
  assign n23046 = ~n21734 & n23045 ;
  assign n23047 = ~n23044 & ~n23046 ;
  assign n23048 = \pi0715  & n23047 ;
  assign n23049 = ~n23043 & n23048 ;
  assign n23050 = ~\pi1160  & ~n23049 ;
  assign n23051 = ~n23035 & n23050 ;
  assign n23052 = n21113 & n21768 ;
  assign n23053 = n21113 & n21770 ;
  assign n23054 = ~n21734 & n23053 ;
  assign n23055 = ~n23052 & ~n23054 ;
  assign n23056 = ~\pi0715  & n23055 ;
  assign n23057 = \pi1160  & ~n23056 ;
  assign n23058 = \pi0644  & ~n23041 ;
  assign n23059 = \pi1160  & n23058 ;
  assign n23060 = n23040 & n23059 ;
  assign n23061 = ~n23057 & ~n23060 ;
  assign n23062 = \pi0790  & n23061 ;
  assign n23063 = ~\pi0644  & n23030 ;
  assign n23064 = \pi0790  & ~n23063 ;
  assign n23065 = \pi0787  & \pi0790  ;
  assign n23066 = ~n23024 & n23065 ;
  assign n23067 = ~n23064 & ~n23066 ;
  assign n23068 = \pi0715  & ~n23067 ;
  assign n23069 = ~\pi0644  & n23068 ;
  assign n23070 = ~n23010 & n23068 ;
  assign n23071 = n23015 & n23070 ;
  assign n23072 = ~n23069 & ~n23071 ;
  assign n23073 = ~n23062 & n23072 ;
  assign n23074 = \pi0644  & \pi0787  ;
  assign n23075 = ~n23062 & n23074 ;
  assign n23076 = ~n23007 & n23075 ;
  assign n23077 = ~n23073 & ~n23076 ;
  assign n23078 = ~n21133 & n23077 ;
  assign n23079 = ~n23051 & n23078 ;
  assign n23080 = ~n23020 & ~n23079 ;
  assign n23081 = ~n21129 & n23080 ;
  assign n23082 = ~\pi0141  & \pi0788  ;
  assign n23083 = ~n1689 & n23082 ;
  assign n23084 = ~n20778 & n23083 ;
  assign n23085 = ~\pi0141  & ~n1689 ;
  assign n23086 = \pi0749  & n1689 ;
  assign n23087 = n20784 & n23086 ;
  assign n23088 = ~n23085 & ~n23087 ;
  assign n23089 = n20794 & ~n23088 ;
  assign n23090 = n20796 & ~n23089 ;
  assign n23091 = n20799 & ~n23088 ;
  assign n23092 = n20801 & ~n23091 ;
  assign n23093 = ~n23090 & ~n23092 ;
  assign n23094 = ~\pi0785  & ~n23085 ;
  assign n23095 = ~n23087 & n23094 ;
  assign n23096 = ~n20804 & ~n23095 ;
  assign n23097 = ~n20812 & n23096 ;
  assign n23098 = ~\pi0789  & n23097 ;
  assign n23099 = n23093 & n23098 ;
  assign n23100 = n20816 & n23099 ;
  assign n23101 = n23093 & n23097 ;
  assign n23102 = ~\pi0789  & ~n23101 ;
  assign n23103 = n20820 & n23096 ;
  assign n23104 = n23093 & n23103 ;
  assign n23105 = ~\pi0141  & \pi0619  ;
  assign n23106 = ~n1689 & n23105 ;
  assign n23107 = ~\pi1159  & ~n23106 ;
  assign n23108 = ~n23104 & n23107 ;
  assign n23109 = ~n23102 & ~n23108 ;
  assign n23110 = n20828 & ~n23085 ;
  assign n23111 = ~n20830 & ~n23110 ;
  assign n23112 = n23097 & ~n23110 ;
  assign n23113 = n23093 & n23112 ;
  assign n23114 = ~n23111 & ~n23113 ;
  assign n23115 = n20816 & ~n23114 ;
  assign n23116 = n23109 & n23115 ;
  assign n23117 = ~n23100 & ~n23116 ;
  assign n23118 = ~n23084 & n23117 ;
  assign n23119 = ~\pi0788  & n23099 ;
  assign n23120 = ~\pi0788  & ~n23114 ;
  assign n23121 = n23109 & n23120 ;
  assign n23122 = ~n23119 & ~n23121 ;
  assign n23123 = ~n20846 & n23122 ;
  assign n23124 = n23118 & n23123 ;
  assign n23125 = n20850 & ~n23085 ;
  assign n23126 = ~n20852 & ~n23125 ;
  assign n23127 = \pi0706  & n1689 ;
  assign n23128 = n20855 & n23127 ;
  assign n23129 = ~n20861 & n23128 ;
  assign n23130 = ~n23085 & ~n23129 ;
  assign n23131 = n20879 & ~n23130 ;
  assign n23132 = n20891 & ~n23125 ;
  assign n23133 = n23131 & n23132 ;
  assign n23134 = ~n23126 & ~n23133 ;
  assign n23135 = n20895 & n23131 ;
  assign n23136 = ~\pi0141  & \pi0647  ;
  assign n23137 = ~n1689 & n23136 ;
  assign n23138 = n20897 & ~n23137 ;
  assign n23139 = ~n23135 & n23138 ;
  assign n23140 = ~n23134 & ~n23139 ;
  assign n23141 = n20846 & ~n23085 ;
  assign n23142 = n23140 & ~n23141 ;
  assign n23143 = ~n23124 & n23142 ;
  assign n23144 = n20910 & n23140 ;
  assign n23145 = \pi0787  & ~n23144 ;
  assign n23146 = ~n23143 & n23145 ;
  assign n23147 = ~\pi0644  & ~n23146 ;
  assign n23148 = n20915 & n23131 ;
  assign n23149 = \pi0644  & n23148 ;
  assign n23150 = n20891 & n23131 ;
  assign n23151 = ~\pi0787  & ~n23150 ;
  assign n23152 = ~\pi1157  & ~n23137 ;
  assign n23153 = ~n23135 & n23152 ;
  assign n23154 = ~n23151 & ~n23153 ;
  assign n23155 = n20923 & ~n23085 ;
  assign n23156 = ~n20925 & ~n23155 ;
  assign n23157 = n20891 & ~n23155 ;
  assign n23158 = n23131 & n23157 ;
  assign n23159 = ~n23156 & ~n23158 ;
  assign n23160 = \pi0644  & ~n23159 ;
  assign n23161 = n23154 & n23160 ;
  assign n23162 = ~n23149 & ~n23161 ;
  assign n23163 = ~\pi0715  & n23162 ;
  assign n23164 = ~n23147 & n23163 ;
  assign n23165 = n20947 & n23099 ;
  assign n23166 = n20947 & ~n23114 ;
  assign n23167 = n23109 & n23166 ;
  assign n23168 = ~n23165 & ~n23167 ;
  assign n23169 = ~n20878 & n20951 ;
  assign n23170 = n20873 & n23169 ;
  assign n23171 = ~n23130 & n23170 ;
  assign n23172 = ~n20778 & n23085 ;
  assign n23173 = ~n20883 & n23172 ;
  assign n23174 = ~n23171 & ~n23173 ;
  assign n23175 = n23168 & n23174 ;
  assign n23176 = \pi0788  & ~n23175 ;
  assign n23177 = ~\pi0789  & ~n21038 ;
  assign n23178 = n20874 & ~n23106 ;
  assign n23179 = ~n23104 & n23178 ;
  assign n23180 = n21050 & ~n23085 ;
  assign n23181 = ~n23129 & n23180 ;
  assign n23182 = ~n21051 & ~n23181 ;
  assign n23183 = ~n23179 & n23182 ;
  assign n23184 = n21039 & ~n23085 ;
  assign n23185 = ~n21041 & ~n23184 ;
  assign n23186 = n23097 & ~n23184 ;
  assign n23187 = n23093 & n23186 ;
  assign n23188 = ~n23185 & ~n23187 ;
  assign n23189 = ~n21038 & ~n23188 ;
  assign n23190 = n23183 & n23189 ;
  assign n23191 = ~n23177 & ~n23190 ;
  assign n23192 = ~\pi0628  & n23191 ;
  assign n23193 = n20964 & n23096 ;
  assign n23194 = n23093 & n23193 ;
  assign n23195 = \pi0627  & ~n23085 ;
  assign n23196 = ~n23129 & n23195 ;
  assign n23197 = ~n20968 & ~n23196 ;
  assign n23198 = ~n23194 & ~n23197 ;
  assign n23199 = n20974 & n23096 ;
  assign n23200 = n23093 & n23199 ;
  assign n23201 = ~\pi0627  & ~n23085 ;
  assign n23202 = ~n23129 & n23201 ;
  assign n23203 = ~n20978 & ~n23202 ;
  assign n23204 = ~n23200 & ~n23203 ;
  assign n23205 = ~n23198 & ~n23204 ;
  assign n23206 = \pi0781  & n23205 ;
  assign n23207 = ~n21034 & ~n23206 ;
  assign n23208 = \pi0680  & \pi0706  ;
  assign n23209 = ~n20854 & n23208 ;
  assign n23210 = ~n20861 & n23209 ;
  assign n23211 = ~n20986 & n23210 ;
  assign n23212 = \pi0603  & \pi0749  ;
  assign n23213 = ~n20783 & n23212 ;
  assign n23214 = ~n20985 & n23213 ;
  assign n23215 = ~n23085 & ~n23214 ;
  assign n23216 = ~n23211 & n23215 ;
  assign n23217 = \pi0141  & ~n1689 ;
  assign n23218 = ~\pi0609  & ~n23217 ;
  assign n23219 = ~n23216 & n23218 ;
  assign n23220 = ~\pi1155  & ~n23085 ;
  assign n23221 = ~n23129 & n23220 ;
  assign n23222 = ~n20999 & ~n23221 ;
  assign n23223 = ~n23219 & ~n23222 ;
  assign n23224 = \pi1155  & ~n23091 ;
  assign n23225 = ~\pi0660  & ~n23224 ;
  assign n23226 = ~n23223 & n23225 ;
  assign n23227 = ~n21007 & ~n23090 ;
  assign n23228 = \pi0609  & ~n23217 ;
  assign n23229 = ~n23216 & n23228 ;
  assign n23230 = ~\pi0609  & ~n23130 ;
  assign n23231 = n20801 & ~n23230 ;
  assign n23232 = ~n23229 & n23231 ;
  assign n23233 = n23227 & ~n23232 ;
  assign n23234 = ~n23226 & ~n23233 ;
  assign n23235 = ~n23216 & ~n23217 ;
  assign n23236 = ~\pi0785  & ~n23235 ;
  assign n23237 = n21022 & ~n23236 ;
  assign n23238 = ~n23234 & n23237 ;
  assign n23239 = ~\pi0628  & ~n23238 ;
  assign n23240 = n23207 & n23239 ;
  assign n23241 = ~n23192 & ~n23240 ;
  assign n23242 = ~n23176 & ~n23241 ;
  assign n23243 = \pi0628  & n23122 ;
  assign n23244 = n23118 & n23243 ;
  assign n23245 = ~\pi1156  & ~n23244 ;
  assign n23246 = ~n23242 & n23245 ;
  assign n23247 = n21077 & n23131 ;
  assign n23248 = ~\pi0629  & ~n23247 ;
  assign n23249 = ~n23246 & n23248 ;
  assign n23250 = n20939 & n23131 ;
  assign n23251 = ~n20935 & ~n23250 ;
  assign n23252 = ~\pi0628  & n23122 ;
  assign n23253 = n23118 & n23252 ;
  assign n23254 = n20944 & ~n23253 ;
  assign n23255 = n23251 & ~n23254 ;
  assign n23256 = n23207 & ~n23238 ;
  assign n23257 = ~n23191 & ~n23256 ;
  assign n23258 = ~n23176 & ~n23257 ;
  assign n23259 = \pi0628  & n23251 ;
  assign n23260 = n23258 & n23259 ;
  assign n23261 = ~n23255 & ~n23260 ;
  assign n23262 = ~n23249 & n23261 ;
  assign n23263 = \pi0788  & ~\pi0792  ;
  assign n23264 = ~n23175 & n23263 ;
  assign n23265 = ~\pi0792  & ~n23191 ;
  assign n23266 = ~n23256 & n23265 ;
  assign n23267 = ~n21067 & ~n23266 ;
  assign n23268 = ~n23264 & n23267 ;
  assign n23269 = n23163 & n23268 ;
  assign n23270 = ~n23262 & n23269 ;
  assign n23271 = ~n23164 & ~n23270 ;
  assign n23272 = ~n21088 & ~n23084 ;
  assign n23273 = n23117 & n23272 ;
  assign n23274 = n23123 & n23273 ;
  assign n23275 = ~n21092 & ~n23085 ;
  assign n23276 = ~\pi0644  & ~n23275 ;
  assign n23277 = ~n23274 & n23276 ;
  assign n23278 = ~\pi0141  & \pi0644  ;
  assign n23279 = ~n1689 & n23278 ;
  assign n23280 = \pi0715  & ~n23279 ;
  assign n23281 = ~n23277 & n23280 ;
  assign n23282 = ~\pi1160  & ~n23281 ;
  assign n23283 = n23271 & n23282 ;
  assign n23284 = \pi0790  & n23283 ;
  assign n23285 = \pi0644  & ~n23146 ;
  assign n23286 = ~\pi0644  & n23148 ;
  assign n23287 = ~\pi0644  & ~n23159 ;
  assign n23288 = n23154 & n23287 ;
  assign n23289 = ~n23286 & ~n23288 ;
  assign n23290 = ~n23285 & n23289 ;
  assign n23291 = n23268 & n23289 ;
  assign n23292 = ~n23262 & n23291 ;
  assign n23293 = ~n23290 & ~n23292 ;
  assign n23294 = \pi0715  & ~n23293 ;
  assign n23295 = ~\pi0141  & ~\pi0644  ;
  assign n23296 = ~n1689 & n23295 ;
  assign n23297 = ~\pi0715  & ~n23296 ;
  assign n23298 = \pi1160  & ~n23297 ;
  assign n23299 = \pi0644  & ~n23275 ;
  assign n23300 = \pi1160  & n23299 ;
  assign n23301 = ~n23274 & n23300 ;
  assign n23302 = ~n23298 & ~n23301 ;
  assign n23303 = \pi0790  & ~n23302 ;
  assign n23304 = ~n23294 & n23303 ;
  assign n23305 = ~n23284 & ~n23304 ;
  assign n23306 = ~\pi0790  & ~n23146 ;
  assign n23307 = \pi0832  & ~n23306 ;
  assign n23308 = \pi0832  & n23268 ;
  assign n23309 = ~n23262 & n23308 ;
  assign n23310 = ~n23307 & ~n23309 ;
  assign n23311 = n23305 & ~n23310 ;
  assign n23312 = \pi0644  & ~\pi0715  ;
  assign n23313 = ~\pi0644  & \pi0715  ;
  assign n23314 = ~n23312 & ~n23313 ;
  assign n23315 = \pi0715  & \pi1160  ;
  assign n23316 = ~\pi0715  & ~\pi1160  ;
  assign n23317 = ~n23315 & ~n23316 ;
  assign n23318 = n23314 & ~n23317 ;
  assign n23319 = n9948 & n23318 ;
  assign n23320 = ~\pi0141  & \pi0628  ;
  assign n23321 = n21768 & n23320 ;
  assign n23322 = n21770 & n23320 ;
  assign n23323 = ~n21734 & n23322 ;
  assign n23324 = ~n23321 & ~n23323 ;
  assign n23325 = n20887 & n23324 ;
  assign n23326 = \pi0141  & ~n6861 ;
  assign n23327 = ~\pi0141  & ~\pi0706  ;
  assign n23328 = n22124 & n23327 ;
  assign n23329 = n21770 & n23327 ;
  assign n23330 = ~n21734 & n23329 ;
  assign n23331 = ~n23328 & ~n23330 ;
  assign n23332 = n6861 & n23331 ;
  assign n23333 = ~n23326 & ~n23332 ;
  assign n23334 = ~\pi0039  & ~\pi0141  ;
  assign n23335 = ~\pi0141  & ~n21930 ;
  assign n23336 = n21992 & n23335 ;
  assign n23337 = ~n23334 & ~n23336 ;
  assign n23338 = ~n22017 & ~n23337 ;
  assign n23339 = ~\pi0038  & ~\pi0141  ;
  assign n23340 = ~n22109 & ~n23339 ;
  assign n23341 = ~n23338 & ~n23340 ;
  assign n23342 = ~\pi0141  & ~n21757 ;
  assign n23343 = n22117 & ~n23342 ;
  assign n23344 = \pi0706  & ~n23326 ;
  assign n23345 = ~n23343 & n23344 ;
  assign n23346 = ~n23341 & n23345 ;
  assign n23347 = n22151 & ~n23346 ;
  assign n23348 = ~n23333 & n23347 ;
  assign n23349 = n22849 & n23348 ;
  assign n23350 = \pi0625  & n23346 ;
  assign n23351 = \pi0625  & ~n23326 ;
  assign n23352 = ~n23332 & n23351 ;
  assign n23353 = ~n23350 & ~n23352 ;
  assign n23354 = ~\pi0141  & ~\pi0625  ;
  assign n23355 = n21768 & n23354 ;
  assign n23356 = n21770 & n23354 ;
  assign n23357 = ~n21734 & n23356 ;
  assign n23358 = ~n23355 & ~n23357 ;
  assign n23359 = \pi1153  & n23358 ;
  assign n23360 = n23353 & n23359 ;
  assign n23361 = ~\pi0625  & n23346 ;
  assign n23362 = ~\pi0625  & ~n23326 ;
  assign n23363 = ~n23332 & n23362 ;
  assign n23364 = ~n23361 & ~n23363 ;
  assign n23365 = ~\pi0141  & \pi0625  ;
  assign n23366 = n21768 & n23365 ;
  assign n23367 = n21770 & n23365 ;
  assign n23368 = ~n21734 & n23367 ;
  assign n23369 = ~n23366 & ~n23368 ;
  assign n23370 = ~\pi1153  & n23369 ;
  assign n23371 = n23364 & n23370 ;
  assign n23372 = ~n23360 & ~n23371 ;
  assign n23373 = n22148 & n22849 ;
  assign n23374 = ~n23372 & n23373 ;
  assign n23375 = ~n23349 & ~n23374 ;
  assign n23376 = ~\pi0141  & n21768 ;
  assign n23377 = ~\pi0141  & n21770 ;
  assign n23378 = ~n21734 & n23377 ;
  assign n23379 = ~n23376 & ~n23378 ;
  assign n23380 = ~n22147 & ~n22155 ;
  assign n23381 = ~n22160 & ~n23380 ;
  assign n23382 = n23379 & n23381 ;
  assign n23383 = n22160 & n23379 ;
  assign n23384 = ~n22161 & ~n23383 ;
  assign n23385 = ~n23382 & n23384 ;
  assign n23386 = n23375 & n23385 ;
  assign n23387 = n22161 & ~n23379 ;
  assign n23388 = ~\pi1156  & n23324 ;
  assign n23389 = ~n23387 & n23388 ;
  assign n23390 = ~n23386 & n23389 ;
  assign n23391 = ~n23325 & ~n23390 ;
  assign n23392 = ~\pi0141  & ~\pi0628  ;
  assign n23393 = n21768 & n23392 ;
  assign n23394 = n21770 & n23392 ;
  assign n23395 = ~n21734 & n23394 ;
  assign n23396 = ~n23393 & ~n23395 ;
  assign n23397 = n20886 & n23396 ;
  assign n23398 = \pi1156  & n23396 ;
  assign n23399 = ~n23387 & n23398 ;
  assign n23400 = ~n23386 & n23399 ;
  assign n23401 = ~n23397 & ~n23400 ;
  assign n23402 = n23391 & n23401 ;
  assign n23403 = n22956 & ~n23402 ;
  assign n23404 = ~\pi0792  & ~n23387 ;
  assign n23405 = \pi0647  & n23404 ;
  assign n23406 = ~n23386 & n23405 ;
  assign n23407 = ~\pi0647  & n23379 ;
  assign n23408 = \pi1157  & ~n23407 ;
  assign n23409 = ~n23406 & n23408 ;
  assign n23410 = ~n23403 & n23409 ;
  assign n23411 = \pi0787  & ~n23410 ;
  assign n23412 = ~\pi0715  & \pi1160  ;
  assign n23413 = \pi0715  & ~\pi1160  ;
  assign n23414 = ~n23412 & ~n23413 ;
  assign n23415 = ~n21088 & ~n23314 ;
  assign n23416 = ~n23414 & ~n23415 ;
  assign n23417 = ~n23379 & n23416 ;
  assign n23418 = ~n23314 & ~n23414 ;
  assign n23419 = ~n21088 & n23418 ;
  assign n23420 = \pi0790  & ~n23419 ;
  assign n23421 = ~n23417 & n23420 ;
  assign n23422 = ~n20811 & ~n23379 ;
  assign n23423 = \pi0789  & ~n21032 ;
  assign n23424 = \pi0781  & ~n23423 ;
  assign n23425 = n23422 & n23424 ;
  assign n23426 = n21777 & n23326 ;
  assign n23427 = ~\pi0749  & ~n21731 ;
  assign n23428 = n21714 & n23427 ;
  assign n23429 = ~n21693 & n23428 ;
  assign n23430 = ~n21552 & n21562 ;
  assign n23431 = n21543 & ~n23430 ;
  assign n23432 = \pi0141  & ~n21536 ;
  assign n23433 = ~n23431 & n23432 ;
  assign n23434 = ~\pi0038  & ~n23433 ;
  assign n23435 = ~n23429 & n23434 ;
  assign n23436 = ~n1288 & ~n23435 ;
  assign n23437 = n1354 & n23087 ;
  assign n23438 = n8413 & n23437 ;
  assign n23439 = n1358 & n23438 ;
  assign n23440 = \pi0038  & n23439 ;
  assign n23441 = \pi0038  & ~\pi0141  ;
  assign n23442 = ~n21757 & n23441 ;
  assign n23443 = ~n23440 & ~n23442 ;
  assign n23444 = n23436 & n23443 ;
  assign n23445 = ~\pi0141  & ~n21467 ;
  assign n23446 = n21272 & n23334 ;
  assign n23447 = ~n23445 & ~n23446 ;
  assign n23448 = \pi0141  & ~n21484 ;
  assign n23449 = \pi0749  & ~n23448 ;
  assign n23450 = n23447 & n23449 ;
  assign n23451 = ~\pi0141  & ~\pi0749  ;
  assign n23452 = n21743 & n23451 ;
  assign n23453 = n23443 & ~n23452 ;
  assign n23454 = ~n23450 & n23453 ;
  assign n23455 = ~n23444 & ~n23454 ;
  assign n23456 = n6861 & n21777 ;
  assign n23457 = ~n23455 & n23456 ;
  assign n23458 = ~n23426 & ~n23457 ;
  assign n23459 = ~n21777 & n23379 ;
  assign n23460 = n20811 & ~n23459 ;
  assign n23461 = n23424 & n23460 ;
  assign n23462 = n23458 & n23461 ;
  assign n23463 = ~n23425 & ~n23462 ;
  assign n23464 = ~\pi0781  & ~n23459 ;
  assign n23465 = ~n23423 & n23464 ;
  assign n23466 = n23458 & n23465 ;
  assign n23467 = ~n23379 & n23423 ;
  assign n23468 = ~\pi0788  & ~n23467 ;
  assign n23469 = ~n23466 & n23468 ;
  assign n23470 = n23463 & n23469 ;
  assign n23471 = ~n20846 & ~n23470 ;
  assign n23472 = \pi0790  & n23379 ;
  assign n23473 = \pi0790  & ~n20846 ;
  assign n23474 = ~n23416 & n23473 ;
  assign n23475 = ~n23472 & ~n23474 ;
  assign n23476 = ~n23471 & ~n23475 ;
  assign n23477 = ~\pi0141  & \pi0626  ;
  assign n23478 = n21768 & n23477 ;
  assign n23479 = n21770 & n23477 ;
  assign n23480 = ~n21734 & n23479 ;
  assign n23481 = ~n23478 & ~n23480 ;
  assign n23482 = n20777 & n23481 ;
  assign n23483 = ~\pi1158  & n23481 ;
  assign n23484 = ~n23467 & n23483 ;
  assign n23485 = ~n23466 & n23484 ;
  assign n23486 = n23463 & n23485 ;
  assign n23487 = ~n23482 & ~n23486 ;
  assign n23488 = ~\pi0141  & ~\pi0626  ;
  assign n23489 = n21768 & n23488 ;
  assign n23490 = n21770 & n23488 ;
  assign n23491 = ~n21734 & n23490 ;
  assign n23492 = ~n23489 & ~n23491 ;
  assign n23493 = n20776 & n23492 ;
  assign n23494 = \pi1158  & n23492 ;
  assign n23495 = ~n23467 & n23494 ;
  assign n23496 = ~n23466 & n23495 ;
  assign n23497 = n23463 & n23496 ;
  assign n23498 = ~n23493 & ~n23497 ;
  assign n23499 = n23487 & n23498 ;
  assign n23500 = \pi0788  & ~n23475 ;
  assign n23501 = ~n23499 & n23500 ;
  assign n23502 = ~n23476 & ~n23501 ;
  assign n23503 = ~n23421 & n23502 ;
  assign n23504 = n22913 & ~n23402 ;
  assign n23505 = ~\pi0647  & n23404 ;
  assign n23506 = ~n23386 & n23505 ;
  assign n23507 = \pi0647  & n23379 ;
  assign n23508 = ~\pi1157  & ~n23507 ;
  assign n23509 = ~n23506 & n23508 ;
  assign n23510 = ~n23504 & n23509 ;
  assign n23511 = ~n23503 & ~n23510 ;
  assign n23512 = n23411 & n23511 ;
  assign n23513 = n23011 & ~n23402 ;
  assign n23514 = ~\pi0787  & n23404 ;
  assign n23515 = ~n23386 & n23514 ;
  assign n23516 = ~\pi0644  & ~n23315 ;
  assign n23517 = \pi0644  & ~n23316 ;
  assign n23518 = ~n23516 & ~n23517 ;
  assign n23519 = ~n23515 & n23518 ;
  assign n23520 = ~n23513 & n23519 ;
  assign n23521 = ~n23503 & ~n23520 ;
  assign n23522 = n9948 & ~n23521 ;
  assign n23523 = ~n23512 & n23522 ;
  assign n23524 = ~n23319 & ~n23523 ;
  assign n23525 = ~n23406 & ~n23407 ;
  assign n23526 = ~n23403 & n23525 ;
  assign n23527 = n20849 & ~n23526 ;
  assign n23528 = n20846 & ~n23379 ;
  assign n23529 = ~n20910 & ~n23528 ;
  assign n23530 = ~n23471 & n23529 ;
  assign n23531 = \pi0788  & n23529 ;
  assign n23532 = ~n23499 & n23531 ;
  assign n23533 = ~n23530 & ~n23532 ;
  assign n23534 = ~n20897 & n23533 ;
  assign n23535 = ~n23506 & ~n23507 ;
  assign n23536 = n23533 & n23535 ;
  assign n23537 = ~n23504 & n23536 ;
  assign n23538 = ~n23534 & ~n23537 ;
  assign n23539 = ~n23527 & ~n23538 ;
  assign n23540 = n21067 & n23539 ;
  assign n23541 = \pi0790  & ~n23521 ;
  assign n23542 = ~n23512 & n23541 ;
  assign n23543 = ~n23540 & ~n23542 ;
  assign n23544 = ~n23524 & ~n23543 ;
  assign n23545 = ~n22683 & n23334 ;
  assign n23546 = n2297 & n22630 ;
  assign n23547 = n6205 & n22601 ;
  assign n23548 = ~n23546 & ~n23547 ;
  assign n23549 = ~\pi0141  & ~n23548 ;
  assign n23550 = \pi0749  & ~n23549 ;
  assign n23551 = ~n23545 & n23550 ;
  assign n23552 = \pi0039  & ~n22468 ;
  assign n23553 = \pi0039  & ~n22509 ;
  assign n23554 = n22487 & n23553 ;
  assign n23555 = ~n23552 & ~n23554 ;
  assign n23556 = n2297 & ~n22530 ;
  assign n23557 = n23555 & ~n23556 ;
  assign n23558 = ~\pi0039  & n22693 ;
  assign n23559 = \pi0141  & ~n23558 ;
  assign n23560 = n23557 & n23559 ;
  assign n23561 = ~\pi0038  & ~n23560 ;
  assign n23562 = n23551 & n23561 ;
  assign n23563 = n6205 & n22407 ;
  assign n23564 = n2297 & n22291 ;
  assign n23565 = ~n23563 & ~n23564 ;
  assign n23566 = ~\pi0039  & n22643 ;
  assign n23567 = ~n22652 & n23566 ;
  assign n23568 = n23565 & ~n23567 ;
  assign n23569 = ~\pi0141  & ~n23568 ;
  assign n23570 = \pi0039  & n22379 ;
  assign n23571 = n2297 & ~n22431 ;
  assign n23572 = ~n23570 & ~n23571 ;
  assign n23573 = n21471 & ~n22665 ;
  assign n23574 = n21479 & ~n22676 ;
  assign n23575 = ~n23573 & ~n23574 ;
  assign n23576 = \pi0141  & n23575 ;
  assign n23577 = n23572 & n23576 ;
  assign n23578 = ~\pi0038  & ~\pi0749  ;
  assign n23579 = ~n23577 & n23578 ;
  assign n23580 = ~n23569 & n23579 ;
  assign n23581 = ~n23562 & ~n23580 ;
  assign n23582 = ~n23342 & ~n23439 ;
  assign n23583 = n20855 & n21417 ;
  assign n23584 = n8413 & n23583 ;
  assign n23585 = n1354 & n23584 ;
  assign n23586 = n1358 & n23585 ;
  assign n23587 = \pi0038  & ~n23586 ;
  assign n23588 = n23582 & n23587 ;
  assign n23589 = \pi0706  & ~n23588 ;
  assign n23590 = n23581 & n23589 ;
  assign n23591 = ~\pi0706  & n23455 ;
  assign n23592 = n22698 & ~n23591 ;
  assign n23593 = ~n23590 & n23592 ;
  assign n23594 = ~n22734 & ~n23354 ;
  assign n23595 = ~n23593 & ~n23594 ;
  assign n23596 = ~n22727 & ~n23365 ;
  assign n23597 = ~\pi1153  & n23596 ;
  assign n23598 = ~\pi1153  & n6861 ;
  assign n23599 = ~n23455 & n23598 ;
  assign n23600 = ~n23597 & ~n23599 ;
  assign n23601 = ~n23595 & ~n23600 ;
  assign n23602 = ~\pi0608  & ~n23360 ;
  assign n23603 = ~n23601 & n23602 ;
  assign n23604 = ~n23593 & ~n23596 ;
  assign n23605 = \pi1153  & n23594 ;
  assign n23606 = \pi1153  & n6861 ;
  assign n23607 = ~n23455 & n23606 ;
  assign n23608 = ~n23605 & ~n23607 ;
  assign n23609 = ~n23604 & ~n23608 ;
  assign n23610 = \pi0608  & ~n23371 ;
  assign n23611 = ~n23609 & n23610 ;
  assign n23612 = ~n23603 & ~n23611 ;
  assign n23613 = ~\pi0609  & \pi0778  ;
  assign n23614 = ~n23612 & n23613 ;
  assign n23615 = \pi0778  & ~n23372 ;
  assign n23616 = ~\pi0778  & ~n23346 ;
  assign n23617 = ~n23333 & n23616 ;
  assign n23618 = \pi0609  & ~n23617 ;
  assign n23619 = ~n23615 & n23618 ;
  assign n23620 = ~\pi0141  & ~\pi0778  ;
  assign n23621 = ~\pi0778  & n1289 ;
  assign n23622 = n1287 & n23621 ;
  assign n23623 = ~n23620 & ~n23622 ;
  assign n23624 = ~\pi0609  & ~n23623 ;
  assign n23625 = ~n23593 & n23624 ;
  assign n23626 = ~\pi1155  & ~n23625 ;
  assign n23627 = ~n23619 & n23626 ;
  assign n23628 = ~n23614 & n23627 ;
  assign n23629 = n22788 & n23326 ;
  assign n23630 = n6861 & n22788 ;
  assign n23631 = ~n23455 & n23630 ;
  assign n23632 = ~n23629 & ~n23631 ;
  assign n23633 = ~n22788 & n23379 ;
  assign n23634 = ~\pi0660  & ~n23633 ;
  assign n23635 = n23632 & n23634 ;
  assign n23636 = ~n22787 & ~n23635 ;
  assign n23637 = ~n23628 & ~n23636 ;
  assign n23638 = \pi0609  & \pi0778  ;
  assign n23639 = ~n23612 & n23638 ;
  assign n23640 = \pi0609  & ~n23623 ;
  assign n23641 = ~n23593 & n23640 ;
  assign n23642 = ~\pi0609  & ~n23617 ;
  assign n23643 = \pi1155  & ~n23642 ;
  assign n23644 = n22722 & ~n23372 ;
  assign n23645 = ~n23643 & ~n23644 ;
  assign n23646 = ~n23641 & ~n23645 ;
  assign n23647 = ~n23639 & n23646 ;
  assign n23648 = n22767 & n23326 ;
  assign n23649 = n6861 & n22767 ;
  assign n23650 = ~n23455 & n23649 ;
  assign n23651 = ~n23648 & ~n23650 ;
  assign n23652 = ~n22767 & n23379 ;
  assign n23653 = \pi0660  & ~n23652 ;
  assign n23654 = n23651 & n23653 ;
  assign n23655 = ~n22766 & ~n23654 ;
  assign n23656 = ~n23647 & ~n23655 ;
  assign n23657 = ~n23637 & ~n23656 ;
  assign n23658 = n22148 & ~n23372 ;
  assign n23659 = ~n23348 & ~n23658 ;
  assign n23660 = n23458 & n23460 ;
  assign n23661 = n20871 & ~n23422 ;
  assign n23662 = ~n23660 & n23661 ;
  assign n23663 = n22147 & n23379 ;
  assign n23664 = ~n23662 & ~n23663 ;
  assign n23665 = n23659 & n23664 ;
  assign n23666 = ~n21016 & ~n21019 ;
  assign n23667 = ~n20811 & n23666 ;
  assign n23668 = ~n23662 & ~n23667 ;
  assign n23669 = \pi0781  & ~n23668 ;
  assign n23670 = ~n23665 & n23669 ;
  assign n23671 = \pi0785  & ~n23670 ;
  assign n23672 = ~n23657 & n23671 ;
  assign n23673 = \pi0778  & ~\pi0785  ;
  assign n23674 = ~n23612 & n23673 ;
  assign n23675 = ~\pi0785  & ~n23623 ;
  assign n23676 = ~n23593 & n23675 ;
  assign n23677 = n21022 & ~n23676 ;
  assign n23678 = ~n23674 & n23677 ;
  assign n23679 = ~n23670 & ~n23678 ;
  assign n23680 = ~\pi0788  & ~n21034 ;
  assign n23681 = ~n23679 & n23680 ;
  assign n23682 = ~n23672 & n23681 ;
  assign n23683 = \pi0781  & n21032 ;
  assign n23684 = n23422 & n23683 ;
  assign n23685 = n23460 & n23683 ;
  assign n23686 = n23458 & n23685 ;
  assign n23687 = ~n23684 & ~n23686 ;
  assign n23688 = n21032 & n23464 ;
  assign n23689 = n23458 & n23688 ;
  assign n23690 = ~n21032 & ~n23379 ;
  assign n23691 = ~n20876 & ~n23690 ;
  assign n23692 = ~n23689 & n23691 ;
  assign n23693 = n23687 & n23692 ;
  assign n23694 = \pi0789  & n23693 ;
  assign n23695 = n23379 & ~n23380 ;
  assign n23696 = ~n22155 & n23348 ;
  assign n23697 = n22148 & ~n22155 ;
  assign n23698 = ~n23372 & n23697 ;
  assign n23699 = ~n23696 & ~n23698 ;
  assign n23700 = ~n23695 & n23699 ;
  assign n23701 = \pi0789  & n21050 ;
  assign n23702 = ~n23700 & n23701 ;
  assign n23703 = ~n23694 & ~n23702 ;
  assign n23704 = ~\pi0788  & ~n23703 ;
  assign n23705 = ~\pi0628  & ~n23704 ;
  assign n23706 = ~n23682 & n23705 ;
  assign n23707 = \pi0628  & ~n23470 ;
  assign n23708 = ~\pi1156  & ~n23707 ;
  assign n23709 = \pi0788  & ~\pi1156  ;
  assign n23710 = ~n23499 & n23709 ;
  assign n23711 = ~n23708 & ~n23710 ;
  assign n23712 = ~n23706 & ~n23711 ;
  assign n23713 = ~n22899 & ~n23482 ;
  assign n23714 = ~n23486 & n23713 ;
  assign n23715 = ~\pi0626  & ~n21034 ;
  assign n23716 = ~n23679 & n23715 ;
  assign n23717 = ~n23672 & n23716 ;
  assign n23718 = ~\pi0626  & ~n23703 ;
  assign n23719 = ~\pi0626  & ~\pi0641  ;
  assign n23720 = ~\pi0641  & ~n23383 ;
  assign n23721 = ~n23382 & n23720 ;
  assign n23722 = n23375 & n23721 ;
  assign n23723 = ~n23719 & ~n23722 ;
  assign n23724 = ~n23718 & ~n23723 ;
  assign n23725 = ~n23717 & n23724 ;
  assign n23726 = ~n23714 & ~n23725 ;
  assign n23727 = ~n22884 & ~n23493 ;
  assign n23728 = ~n23497 & n23727 ;
  assign n23729 = \pi0626  & ~n21034 ;
  assign n23730 = ~n23679 & n23729 ;
  assign n23731 = ~n23672 & n23730 ;
  assign n23732 = \pi0626  & ~n23703 ;
  assign n23733 = \pi0626  & \pi0641  ;
  assign n23734 = \pi0641  & ~n23383 ;
  assign n23735 = ~n23382 & n23734 ;
  assign n23736 = n23375 & n23735 ;
  assign n23737 = ~n23733 & ~n23736 ;
  assign n23738 = ~n23732 & ~n23737 ;
  assign n23739 = ~n23731 & n23738 ;
  assign n23740 = ~n23728 & ~n23739 ;
  assign n23741 = ~n23726 & ~n23740 ;
  assign n23742 = \pi0788  & ~n23711 ;
  assign n23743 = ~n23741 & n23742 ;
  assign n23744 = ~n23712 & ~n23743 ;
  assign n23745 = ~\pi0629  & n23401 ;
  assign n23746 = n23744 & n23745 ;
  assign n23747 = \pi0629  & ~n23325 ;
  assign n23748 = ~n23390 & n23747 ;
  assign n23749 = \pi0792  & ~n23748 ;
  assign n23750 = \pi0628  & ~n23704 ;
  assign n23751 = ~n23682 & n23750 ;
  assign n23752 = ~\pi0628  & ~n23470 ;
  assign n23753 = \pi1156  & ~n23752 ;
  assign n23754 = n21860 & ~n23499 ;
  assign n23755 = ~n23753 & ~n23754 ;
  assign n23756 = \pi0792  & ~n23755 ;
  assign n23757 = ~n23751 & n23756 ;
  assign n23758 = \pi0788  & n23756 ;
  assign n23759 = ~n23741 & n23758 ;
  assign n23760 = ~n23757 & ~n23759 ;
  assign n23761 = ~n23749 & n23760 ;
  assign n23762 = ~n23746 & ~n23761 ;
  assign n23763 = ~n23682 & ~n23704 ;
  assign n23764 = ~\pi0792  & ~n23763 ;
  assign n23765 = n23263 & ~n23741 ;
  assign n23766 = ~n23764 & ~n23765 ;
  assign n23767 = \pi0787  & ~n23539 ;
  assign n23768 = n23766 & ~n23767 ;
  assign n23769 = ~n23524 & n23768 ;
  assign n23770 = ~n23762 & n23769 ;
  assign n23771 = ~n23544 & ~n23770 ;
  assign n23772 = \pi0141  & ~\pi0832  ;
  assign n23773 = ~n21132 & ~n23772 ;
  assign n23774 = n23771 & ~n23773 ;
  assign n23775 = ~n23311 & ~n23774 ;
  assign n23776 = \pi0735  & n1689 ;
  assign n23777 = ~\pi0625  & \pi0680  ;
  assign n23778 = ~n20854 & n23777 ;
  assign n23779 = n23776 & n23778 ;
  assign n23780 = \pi0142  & ~n1689 ;
  assign n23781 = \pi0608  & ~\pi1153  ;
  assign n23782 = ~n23780 & n23781 ;
  assign n23783 = ~n23779 & n23782 ;
  assign n23784 = n20855 & n23776 ;
  assign n23785 = ~\pi0608  & ~n23784 ;
  assign n23786 = \pi0625  & ~n23785 ;
  assign n23787 = \pi1153  & ~n23780 ;
  assign n23788 = \pi0608  & \pi0743  ;
  assign n23789 = n1689 & n23788 ;
  assign n23790 = n20784 & n23789 ;
  assign n23791 = n23787 & ~n23790 ;
  assign n23792 = ~n23786 & n23791 ;
  assign n23793 = ~n23783 & ~n23792 ;
  assign n23794 = ~n20986 & n23784 ;
  assign n23795 = \pi0743  & n1689 ;
  assign n23796 = n20784 & n23795 ;
  assign n23797 = ~n23780 & ~n23796 ;
  assign n23798 = ~n23794 & n23797 ;
  assign n23799 = ~\pi0608  & n20858 ;
  assign n23800 = ~n20784 & n23799 ;
  assign n23801 = n23784 & n23800 ;
  assign n23802 = ~n23798 & ~n23801 ;
  assign n23803 = n23793 & n23802 ;
  assign n23804 = \pi0609  & ~\pi0660  ;
  assign n23805 = ~\pi0609  & \pi0660  ;
  assign n23806 = ~n23804 & ~n23805 ;
  assign n23807 = n20866 & n23806 ;
  assign n23808 = \pi0785  & ~n23807 ;
  assign n23809 = ~\pi0778  & ~n23798 ;
  assign n23810 = ~n23808 & ~n23809 ;
  assign n23811 = ~n23803 & n23810 ;
  assign n23812 = ~n20861 & n23784 ;
  assign n23813 = ~\pi0609  & ~n23812 ;
  assign n23814 = \pi0660  & ~n23813 ;
  assign n23815 = n22788 & n23796 ;
  assign n23816 = \pi1155  & ~n23815 ;
  assign n23817 = ~n23814 & n23816 ;
  assign n23818 = ~n20985 & n23796 ;
  assign n23819 = \pi0660  & ~n23818 ;
  assign n23820 = ~\pi0609  & ~n23819 ;
  assign n23821 = ~\pi0660  & n23812 ;
  assign n23822 = ~\pi1155  & ~n23821 ;
  assign n23823 = ~n23820 & n23822 ;
  assign n23824 = ~n23817 & ~n23823 ;
  assign n23825 = \pi0785  & ~n23780 ;
  assign n23826 = ~n23824 & n23825 ;
  assign n23827 = ~n23811 & ~n23826 ;
  assign n23828 = n21022 & n23827 ;
  assign n23829 = ~n20883 & n23780 ;
  assign n23830 = \pi0781  & ~n20811 ;
  assign n23831 = ~n23423 & ~n23830 ;
  assign n23832 = n21777 & n23831 ;
  assign n23833 = n20947 & n23796 ;
  assign n23834 = n23832 & n23833 ;
  assign n23835 = ~n23829 & ~n23834 ;
  assign n23836 = n20951 & n23780 ;
  assign n23837 = n23380 & n23812 ;
  assign n23838 = n20951 & ~n22160 ;
  assign n23839 = n23837 & n23838 ;
  assign n23840 = ~n23836 & ~n23839 ;
  assign n23841 = n23835 & n23840 ;
  assign n23842 = \pi0788  & ~n23841 ;
  assign n23843 = n20811 & n23666 ;
  assign n23844 = n23796 & n23843 ;
  assign n23845 = n21777 & n23844 ;
  assign n23846 = ~n22147 & n23667 ;
  assign n23847 = n23812 & n23846 ;
  assign n23848 = ~\pi1154  & n21016 ;
  assign n23849 = \pi1154  & n21019 ;
  assign n23850 = n23780 & ~n23849 ;
  assign n23851 = ~n23848 & n23850 ;
  assign n23852 = ~n23847 & ~n23851 ;
  assign n23853 = ~n23845 & n23852 ;
  assign n23854 = \pi0781  & ~n23853 ;
  assign n23855 = n20845 & n20888 ;
  assign n23856 = \pi0792  & ~n23855 ;
  assign n23857 = ~n21034 & ~n23856 ;
  assign n23858 = ~n23854 & n23857 ;
  assign n23859 = ~n23842 & n23858 ;
  assign n23860 = ~n23828 & n23859 ;
  assign n23861 = ~n23842 & ~n23856 ;
  assign n23862 = ~\pi0619  & ~n23837 ;
  assign n23863 = \pi0648  & ~n23862 ;
  assign n23864 = n23796 & ~n23830 ;
  assign n23865 = n21777 & n23864 ;
  assign n23866 = \pi0619  & n23865 ;
  assign n23867 = \pi1159  & ~n23866 ;
  assign n23868 = ~n23863 & n23867 ;
  assign n23869 = \pi0648  & ~n23865 ;
  assign n23870 = ~\pi0619  & ~n23869 ;
  assign n23871 = ~\pi0648  & n23837 ;
  assign n23872 = ~\pi1159  & ~n23871 ;
  assign n23873 = ~n23870 & n23872 ;
  assign n23874 = ~n23868 & ~n23873 ;
  assign n23875 = \pi0789  & ~n23780 ;
  assign n23876 = ~n23874 & n23875 ;
  assign n23877 = ~n21038 & ~n23876 ;
  assign n23878 = n23861 & ~n23877 ;
  assign n23879 = ~n23860 & ~n23878 ;
  assign n23880 = \pi0788  & ~n20778 ;
  assign n23881 = n23796 & ~n23880 ;
  assign n23882 = n23832 & n23881 ;
  assign n23883 = n20887 & ~n23882 ;
  assign n23884 = ~n23780 & ~n23812 ;
  assign n23885 = n22162 & n23380 ;
  assign n23886 = ~n23884 & n23885 ;
  assign n23887 = ~\pi0628  & n23886 ;
  assign n23888 = n20844 & ~n23887 ;
  assign n23889 = ~n23883 & ~n23888 ;
  assign n23890 = ~\pi0628  & ~n23882 ;
  assign n23891 = \pi0629  & ~n23890 ;
  assign n23892 = \pi0628  & n23886 ;
  assign n23893 = \pi1156  & ~n23892 ;
  assign n23894 = ~n23891 & n23893 ;
  assign n23895 = n23889 & ~n23894 ;
  assign n23896 = \pi0792  & ~n23780 ;
  assign n23897 = ~n23895 & n23896 ;
  assign n23898 = ~\pi0647  & ~n23897 ;
  assign n23899 = n23879 & n23898 ;
  assign n23900 = ~n20846 & n23796 ;
  assign n23901 = ~n23880 & n23900 ;
  assign n23902 = n23832 & n23901 ;
  assign n23903 = ~\pi1157  & ~n23780 ;
  assign n23904 = ~n23902 & n23903 ;
  assign n23905 = ~n22945 & ~n23904 ;
  assign n23906 = ~n23899 & ~n23905 ;
  assign n23907 = \pi0792  & ~n20888 ;
  assign n23908 = \pi0647  & ~n23907 ;
  assign n23909 = n23886 & n23908 ;
  assign n23910 = \pi1157  & ~n23780 ;
  assign n23911 = ~n23909 & n23910 ;
  assign n23912 = ~\pi0630  & ~n23911 ;
  assign n23913 = ~n23906 & n23912 ;
  assign n23914 = \pi0647  & ~n23897 ;
  assign n23915 = n23879 & n23914 ;
  assign n23916 = ~n23902 & n23910 ;
  assign n23917 = ~n20925 & ~n23916 ;
  assign n23918 = ~n23915 & ~n23917 ;
  assign n23919 = \pi0630  & ~n23903 ;
  assign n23920 = ~\pi0647  & ~n23907 ;
  assign n23921 = \pi0630  & n23920 ;
  assign n23922 = n23886 & n23921 ;
  assign n23923 = ~n23919 & ~n23922 ;
  assign n23924 = ~n23918 & ~n23923 ;
  assign n23925 = ~n23913 & ~n23924 ;
  assign n23926 = \pi0787  & ~\pi0790  ;
  assign n23927 = ~n23925 & n23926 ;
  assign n23928 = ~\pi0787  & ~n23897 ;
  assign n23929 = ~\pi0790  & n23928 ;
  assign n23930 = n23879 & n23929 ;
  assign n23931 = \pi0832  & ~n23930 ;
  assign n23932 = ~n23927 & n23931 ;
  assign n23933 = \pi0057  & \pi0142  ;
  assign n23934 = ~\pi0832  & ~n23933 ;
  assign n23935 = ~n23932 & ~n23934 ;
  assign n23936 = n23074 & ~n23925 ;
  assign n23937 = \pi0644  & n23928 ;
  assign n23938 = n23879 & n23937 ;
  assign n23939 = \pi0644  & \pi0715  ;
  assign n23940 = \pi0715  & ~n23780 ;
  assign n23941 = ~n23939 & ~n23940 ;
  assign n23942 = \pi0787  & ~n21065 ;
  assign n23943 = ~n23907 & ~n23942 ;
  assign n23944 = ~n23939 & n23943 ;
  assign n23945 = n23886 & n23944 ;
  assign n23946 = ~n23941 & ~n23945 ;
  assign n23947 = ~n23938 & n23946 ;
  assign n23948 = ~n23936 & n23947 ;
  assign n23949 = \pi0644  & ~n21088 ;
  assign n23950 = n23902 & n23949 ;
  assign n23951 = ~\pi0715  & ~n23780 ;
  assign n23952 = ~n23950 & n23951 ;
  assign n23953 = \pi1160  & ~n23952 ;
  assign n23954 = ~n23948 & n23953 ;
  assign n23955 = n23021 & ~n23925 ;
  assign n23956 = ~\pi0644  & n23928 ;
  assign n23957 = n23879 & n23956 ;
  assign n23958 = ~\pi0644  & ~\pi0715  ;
  assign n23959 = ~n23951 & ~n23958 ;
  assign n23960 = n23943 & ~n23958 ;
  assign n23961 = n23886 & n23960 ;
  assign n23962 = ~n23959 & ~n23961 ;
  assign n23963 = ~n23957 & n23962 ;
  assign n23964 = ~n23955 & n23963 ;
  assign n23965 = ~\pi1160  & ~n23940 ;
  assign n23966 = ~\pi0644  & ~n21088 ;
  assign n23967 = ~\pi1160  & n23966 ;
  assign n23968 = n23902 & n23967 ;
  assign n23969 = ~n23965 & ~n23968 ;
  assign n23970 = ~n23964 & ~n23969 ;
  assign n23971 = ~n23954 & ~n23970 ;
  assign n23972 = \pi0790  & ~n23934 ;
  assign n23973 = ~n23971 & n23972 ;
  assign n23974 = ~n23935 & ~n23973 ;
  assign n23975 = ~\pi0142  & n6732 ;
  assign n23976 = n6732 & n21658 ;
  assign n23977 = ~n21684 & n23976 ;
  assign n23978 = ~n23975 & ~n23977 ;
  assign n23979 = \pi0039  & \pi0215  ;
  assign n23980 = \pi0299  & n23979 ;
  assign n23981 = n23978 & n23980 ;
  assign n23982 = ~\pi0142  & ~n6732 ;
  assign n23983 = ~n6732 & n21627 ;
  assign n23984 = ~n21726 & n23983 ;
  assign n23985 = ~n23982 & ~n23984 ;
  assign n23986 = n15410 & n23985 ;
  assign n23987 = n23981 & n23986 ;
  assign n23988 = \pi0142  & n15410 ;
  assign n23989 = n21743 & n23988 ;
  assign n23990 = ~n23987 & ~n23989 ;
  assign n23991 = \pi0039  & ~n21693 ;
  assign n23992 = n6730 & n21694 ;
  assign n23993 = ~n21711 & n23992 ;
  assign n23994 = ~n6732 & n21334 ;
  assign n23995 = ~n21330 & n23994 ;
  assign n23996 = ~n2352 & ~n23995 ;
  assign n23997 = ~n23993 & n23996 ;
  assign n23998 = ~n21704 & n21948 ;
  assign n23999 = ~n23997 & n23998 ;
  assign n24000 = ~n23987 & ~n23999 ;
  assign n24001 = n23991 & n24000 ;
  assign n24002 = ~n23990 & ~n24001 ;
  assign n24003 = \pi0142  & n21768 ;
  assign n24004 = ~n20811 & ~n24003 ;
  assign n24005 = ~n24002 & n24004 ;
  assign n24006 = \pi0142  & ~n21205 ;
  assign n24007 = ~n21238 & n24006 ;
  assign n24008 = n21250 & n24007 ;
  assign n24009 = ~\pi0142  & ~n21475 ;
  assign n24010 = \pi0142  & n21205 ;
  assign n24011 = \pi0142  & n21237 ;
  assign n24012 = n21232 & n24011 ;
  assign n24013 = ~n24010 & ~n24012 ;
  assign n24014 = ~\pi0743  & n24013 ;
  assign n24015 = ~n24009 & ~n24014 ;
  assign n24016 = ~n24008 & n24015 ;
  assign n24017 = \pi0299  & ~n24016 ;
  assign n24018 = ~\pi0142  & ~n21481 ;
  assign n24019 = ~n21478 & n24018 ;
  assign n24020 = \pi0743  & ~n24019 ;
  assign n24021 = \pi0142  & ~\pi0743  ;
  assign n24022 = n21740 & n24021 ;
  assign n24023 = n21737 & n24021 ;
  assign n24024 = n21232 & n24023 ;
  assign n24025 = ~n24022 & ~n24024 ;
  assign n24026 = ~\pi0299  & n24025 ;
  assign n24027 = ~n24020 & n24026 ;
  assign n24028 = \pi0198  & n21247 ;
  assign n24029 = ~n21266 & ~n24028 ;
  assign n24030 = n21265 & ~n24029 ;
  assign n24031 = \pi0142  & n24026 ;
  assign n24032 = ~n24030 & n24031 ;
  assign n24033 = ~n24027 & ~n24032 ;
  assign n24034 = ~n24017 & n24033 ;
  assign n24035 = ~\pi0039  & n24034 ;
  assign n24036 = \pi0142  & ~n6861 ;
  assign n24037 = ~\pi0142  & ~n21494 ;
  assign n24038 = \pi0743  & ~n24037 ;
  assign n24039 = \pi0142  & ~n21378 ;
  assign n24040 = ~n21367 & n24039 ;
  assign n24041 = n6761 & ~n24040 ;
  assign n24042 = n24038 & n24041 ;
  assign n24043 = ~\pi0743  & n6761 ;
  assign n24044 = \pi0142  & n24043 ;
  assign n24045 = ~n21711 & n24044 ;
  assign n24046 = ~n24042 & ~n24045 ;
  assign n24047 = \pi0142  & ~n21350 ;
  assign n24048 = \pi0743  & n21499 ;
  assign n24049 = ~n24047 & n24048 ;
  assign n24050 = \pi0142  & n21334 ;
  assign n24051 = ~n21330 & n24050 ;
  assign n24052 = ~\pi0743  & ~n24051 ;
  assign n24053 = ~n6761 & ~n24052 ;
  assign n24054 = ~n24049 & n24053 ;
  assign n24055 = \pi0743  & ~n21516 ;
  assign n24056 = \pi0743  & n21403 ;
  assign n24057 = ~n21399 & n24056 ;
  assign n24058 = ~n24055 & ~n24057 ;
  assign n24059 = ~n21527 & ~n24058 ;
  assign n24060 = \pi0142  & ~n6709 ;
  assign n24061 = n21428 & n24060 ;
  assign n24062 = \pi0142  & n6709 ;
  assign n24063 = n21425 & n24062 ;
  assign n24064 = ~n6761 & ~n24063 ;
  assign n24065 = ~n24061 & n24064 ;
  assign n24066 = n24059 & n24065 ;
  assign n24067 = ~\pi0743  & ~n6761 ;
  assign n24068 = ~\pi0142  & n24067 ;
  assign n24069 = n21627 & n24067 ;
  assign n24070 = ~n21726 & n24069 ;
  assign n24071 = ~n24068 & ~n24070 ;
  assign n24072 = ~n24066 & n24071 ;
  assign n24073 = \pi0743  & n21528 ;
  assign n24074 = \pi0743  & n21526 ;
  assign n24075 = ~n21522 & n24074 ;
  assign n24076 = ~n24073 & ~n24075 ;
  assign n24077 = \pi0142  & \pi0743  ;
  assign n24078 = ~n21413 & n24077 ;
  assign n24079 = ~n21411 & n24078 ;
  assign n24080 = ~n21408 & n24079 ;
  assign n24081 = n6761 & ~n24080 ;
  assign n24082 = n24076 & n24081 ;
  assign n24083 = \pi0223  & ~n24082 ;
  assign n24084 = \pi0223  & n24021 ;
  assign n24085 = ~n21685 & n24084 ;
  assign n24086 = ~n24083 & ~n24085 ;
  assign n24087 = n24072 & ~n24086 ;
  assign n24088 = ~n2165 & ~n24087 ;
  assign n24089 = ~n24054 & n24088 ;
  assign n24090 = n24046 & n24089 ;
  assign n24091 = \pi0603  & \pi0743  ;
  assign n24092 = ~n20783 & n24091 ;
  assign n24093 = n2165 & ~n24092 ;
  assign n24094 = ~n21285 & n24093 ;
  assign n24095 = ~\pi0142  & n2165 ;
  assign n24096 = n21285 & n24095 ;
  assign n24097 = ~n24094 & ~n24096 ;
  assign n24098 = ~\pi0223  & n24097 ;
  assign n24099 = ~n24087 & ~n24098 ;
  assign n24100 = n6205 & ~n24099 ;
  assign n24101 = ~n24090 & n24100 ;
  assign n24102 = ~n24036 & ~n24101 ;
  assign n24103 = ~n6732 & ~n24052 ;
  assign n24104 = ~n24049 & n24103 ;
  assign n24105 = ~n21685 & n24021 ;
  assign n24106 = n6732 & ~n24080 ;
  assign n24107 = n24076 & n24106 ;
  assign n24108 = ~n24105 & n24107 ;
  assign n24109 = ~\pi0743  & ~n6732 ;
  assign n24110 = ~\pi0142  & n24109 ;
  assign n24111 = n21627 & n24109 ;
  assign n24112 = ~n21726 & n24111 ;
  assign n24113 = ~n24110 & ~n24112 ;
  assign n24114 = ~n6732 & ~n24063 ;
  assign n24115 = ~n24061 & n24114 ;
  assign n24116 = n24059 & n24115 ;
  assign n24117 = \pi0215  & ~n24116 ;
  assign n24118 = n24113 & n24117 ;
  assign n24119 = ~n24108 & n24118 ;
  assign n24120 = ~n2352 & ~n24119 ;
  assign n24121 = ~n24104 & n24120 ;
  assign n24122 = ~\pi0743  & n6732 ;
  assign n24123 = \pi0142  & n24122 ;
  assign n24124 = ~n21711 & n24123 ;
  assign n24125 = n6732 & ~n24040 ;
  assign n24126 = n24038 & n24125 ;
  assign n24127 = ~n24124 & ~n24126 ;
  assign n24128 = n24121 & n24127 ;
  assign n24129 = n2352 & ~n24092 ;
  assign n24130 = ~n21285 & n24129 ;
  assign n24131 = ~\pi0142  & n2352 ;
  assign n24132 = n21285 & n24131 ;
  assign n24133 = ~n24130 & ~n24132 ;
  assign n24134 = ~\pi0215  & n24133 ;
  assign n24135 = ~n24119 & ~n24134 ;
  assign n24136 = n2297 & ~n24135 ;
  assign n24137 = ~n24128 & n24136 ;
  assign n24138 = ~\pi0038  & ~n24137 ;
  assign n24139 = n24102 & n24138 ;
  assign n24140 = ~n24035 & n24139 ;
  assign n24141 = ~\pi0039  & \pi0142  ;
  assign n24142 = ~n21289 & n24141 ;
  assign n24143 = n1259 & n23796 ;
  assign n24144 = n1249 & n24143 ;
  assign n24145 = ~\pi0039  & n1281 ;
  assign n24146 = n24144 & n24145 ;
  assign n24147 = \pi0039  & \pi0142  ;
  assign n24148 = \pi0038  & ~n24147 ;
  assign n24149 = ~n24146 & n24148 ;
  assign n24150 = ~n24142 & n24149 ;
  assign n24151 = n6861 & ~n24150 ;
  assign n24152 = ~n24036 & ~n24151 ;
  assign n24153 = n21777 & ~n24152 ;
  assign n24154 = ~n24140 & n24153 ;
  assign n24155 = n20811 & n21777 ;
  assign n24156 = n20811 & ~n24003 ;
  assign n24157 = ~n24002 & n24156 ;
  assign n24158 = ~n24155 & ~n24157 ;
  assign n24159 = ~n24154 & ~n24158 ;
  assign n24160 = ~n24005 & ~n24159 ;
  assign n24161 = n23424 & ~n24160 ;
  assign n24162 = ~\pi0781  & n21777 ;
  assign n24163 = ~\pi0781  & ~n24003 ;
  assign n24164 = ~n24002 & n24163 ;
  assign n24165 = ~n24162 & ~n24164 ;
  assign n24166 = ~n24154 & ~n24165 ;
  assign n24167 = ~n23423 & n24166 ;
  assign n24168 = n23423 & ~n24003 ;
  assign n24169 = ~n24002 & n24168 ;
  assign n24170 = ~\pi0626  & ~n24003 ;
  assign n24171 = ~n24002 & n24170 ;
  assign n24172 = \pi1158  & ~n24171 ;
  assign n24173 = ~n24169 & n24172 ;
  assign n24174 = ~n24167 & n24173 ;
  assign n24175 = ~n24161 & n24174 ;
  assign n24176 = n20776 & ~n24171 ;
  assign n24177 = ~n22884 & ~n24176 ;
  assign n24178 = ~n24175 & n24177 ;
  assign n24179 = n22155 & ~n24005 ;
  assign n24180 = ~n24159 & n24179 ;
  assign n24181 = n1281 & n23784 ;
  assign n24182 = ~\pi0039  & n1259 ;
  assign n24183 = n1249 & n24182 ;
  assign n24184 = n24181 & n24183 ;
  assign n24185 = n24148 & ~n24184 ;
  assign n24186 = ~n24142 & n24185 ;
  assign n24187 = ~n21961 & ~n21965 ;
  assign n24188 = n21954 & n24187 ;
  assign n24189 = \pi0142  & ~n24188 ;
  assign n24190 = ~\pi0142  & n22023 ;
  assign n24191 = ~n22053 & n24190 ;
  assign n24192 = ~n22445 & n24191 ;
  assign n24193 = ~n22456 & n24192 ;
  assign n24194 = \pi0735  & ~n6761 ;
  assign n24195 = ~n24193 & n24194 ;
  assign n24196 = ~n24189 & n24195 ;
  assign n24197 = ~\pi0735  & ~n6761 ;
  assign n24198 = ~\pi0142  & n24197 ;
  assign n24199 = n21627 & n24197 ;
  assign n24200 = ~n21726 & n24199 ;
  assign n24201 = ~n24198 & ~n24200 ;
  assign n24202 = ~n24196 & n24201 ;
  assign n24203 = ~\pi0142  & ~\pi0735  ;
  assign n24204 = ~\pi0735  & n21658 ;
  assign n24205 = ~n21684 & n24204 ;
  assign n24206 = ~n24203 & ~n24205 ;
  assign n24207 = \pi0142  & ~n21980 ;
  assign n24208 = \pi0735  & ~n24192 ;
  assign n24209 = ~n24207 & n24208 ;
  assign n24210 = \pi0223  & ~n24209 ;
  assign n24211 = n24206 & n24210 ;
  assign n24212 = ~n6764 & ~n24211 ;
  assign n24213 = n24202 & ~n24212 ;
  assign n24214 = ~\pi0299  & ~n24213 ;
  assign n24215 = \pi0142  & n21285 ;
  assign n24216 = ~\pi0120  & n21277 ;
  assign n24217 = n1281 & n24216 ;
  assign n24218 = n1260 & n24217 ;
  assign n24219 = n23784 & n24218 ;
  assign n24220 = \pi0120  & n23784 ;
  assign n24221 = n1281 & n24220 ;
  assign n24222 = n1260 & n24221 ;
  assign n24223 = n2165 & ~n24222 ;
  assign n24224 = ~n24219 & n24223 ;
  assign n24225 = ~n24215 & n24224 ;
  assign n24226 = ~\pi0223  & ~n24225 ;
  assign n24227 = ~n21919 & n21923 ;
  assign n24228 = n22274 & ~n24227 ;
  assign n24229 = \pi0142  & n24228 ;
  assign n24230 = ~\pi0142  & ~n6709 ;
  assign n24231 = ~\pi0142  & ~n21306 ;
  assign n24232 = ~n22022 & n24231 ;
  assign n24233 = ~n24230 & ~n24232 ;
  assign n24234 = ~n22042 & ~n24233 ;
  assign n24235 = \pi0735  & ~n24234 ;
  assign n24236 = ~n24229 & n24235 ;
  assign n24237 = \pi0142  & ~\pi0735  ;
  assign n24238 = n21334 & n24237 ;
  assign n24239 = ~n21330 & n24238 ;
  assign n24240 = ~n2165 & ~n24239 ;
  assign n24241 = ~n24236 & n24240 ;
  assign n24242 = ~n21368 & ~n24241 ;
  assign n24243 = n24226 & n24242 ;
  assign n24244 = \pi0735  & n6761 ;
  assign n24245 = \pi0142  & n6761 ;
  assign n24246 = ~n21711 & n24245 ;
  assign n24247 = ~n24244 & ~n24246 ;
  assign n24248 = ~\pi0142  & \pi0735  ;
  assign n24249 = ~n22067 & n24248 ;
  assign n24250 = ~\pi0680  & n21580 ;
  assign n24251 = \pi0142  & \pi0735  ;
  assign n24252 = n21895 & n24251 ;
  assign n24253 = ~n24250 & n24252 ;
  assign n24254 = ~n24249 & ~n24253 ;
  assign n24255 = n24226 & n24254 ;
  assign n24256 = ~n24247 & n24255 ;
  assign n24257 = ~n24243 & ~n24256 ;
  assign n24258 = n24214 & n24257 ;
  assign n24259 = \pi0735  & n6732 ;
  assign n24260 = \pi0142  & n6732 ;
  assign n24261 = ~n21711 & n24260 ;
  assign n24262 = ~n24259 & ~n24261 ;
  assign n24263 = n24254 & ~n24262 ;
  assign n24264 = \pi0735  & ~n6732 ;
  assign n24265 = ~n24193 & n24264 ;
  assign n24266 = ~n24189 & n24265 ;
  assign n24267 = ~\pi0735  & ~n6732 ;
  assign n24268 = ~\pi0142  & n24267 ;
  assign n24269 = n21627 & n24267 ;
  assign n24270 = ~n21726 & n24269 ;
  assign n24271 = ~n24268 & ~n24270 ;
  assign n24272 = ~n24266 & n24271 ;
  assign n24273 = \pi0215  & ~n24209 ;
  assign n24274 = n24206 & n24273 ;
  assign n24275 = ~n22526 & ~n24274 ;
  assign n24276 = n24272 & ~n24275 ;
  assign n24277 = \pi0299  & ~n24276 ;
  assign n24278 = ~n2352 & ~n24239 ;
  assign n24279 = ~n24236 & n24278 ;
  assign n24280 = ~n21446 & ~n24279 ;
  assign n24281 = n24277 & ~n24280 ;
  assign n24282 = ~n24263 & n24281 ;
  assign n24283 = n2352 & ~n24222 ;
  assign n24284 = ~n24219 & n24283 ;
  assign n24285 = ~n24215 & n24284 ;
  assign n24286 = ~\pi0215  & ~n24285 ;
  assign n24287 = \pi0299  & ~n24286 ;
  assign n24288 = ~n24276 & n24287 ;
  assign n24289 = \pi0039  & ~n24288 ;
  assign n24290 = n6861 & n24289 ;
  assign n24291 = ~n24282 & n24290 ;
  assign n24292 = ~n24258 & n24291 ;
  assign n24293 = ~n24186 & n24292 ;
  assign n24294 = \pi0142  & \pi0299  ;
  assign n24295 = ~n22006 & n24294 ;
  assign n24296 = \pi0735  & ~n24295 ;
  assign n24297 = n11698 & ~n22649 ;
  assign n24298 = ~\pi0142  & ~\pi0299  ;
  assign n24299 = n22103 & n24298 ;
  assign n24300 = ~n22101 & n24299 ;
  assign n24301 = ~\pi0142  & \pi0299  ;
  assign n24302 = n22098 & n24301 ;
  assign n24303 = ~n22095 & n24302 ;
  assign n24304 = ~\pi0038  & ~n24303 ;
  assign n24305 = ~n24300 & n24304 ;
  assign n24306 = ~n24297 & n24305 ;
  assign n24307 = n24296 & n24306 ;
  assign n24308 = n21205 & n24294 ;
  assign n24309 = n21237 & n24294 ;
  assign n24310 = n21232 & n24309 ;
  assign n24311 = ~n24308 & ~n24310 ;
  assign n24312 = ~\pi0735  & n24311 ;
  assign n24313 = n11698 & n21740 ;
  assign n24314 = n11698 & n21737 ;
  assign n24315 = n21232 & n24314 ;
  assign n24316 = ~n24313 & ~n24315 ;
  assign n24317 = ~\pi0038  & n24316 ;
  assign n24318 = n24312 & n24317 ;
  assign n24319 = ~n9627 & ~n24318 ;
  assign n24320 = n6861 & ~n24186 ;
  assign n24321 = n24319 & n24320 ;
  assign n24322 = ~n24307 & n24321 ;
  assign n24323 = ~\pi0142  & ~\pi0625  ;
  assign n24324 = ~n22734 & ~n24323 ;
  assign n24325 = ~n24322 & ~n24324 ;
  assign n24326 = ~n24293 & n24325 ;
  assign n24327 = \pi0625  & ~n24003 ;
  assign n24328 = ~n24002 & n24327 ;
  assign n24329 = ~\pi1153  & ~n24328 ;
  assign n24330 = ~n24326 & n24329 ;
  assign n24331 = ~\pi0142  & \pi0625  ;
  assign n24332 = ~n22727 & ~n24331 ;
  assign n24333 = ~n24322 & ~n24332 ;
  assign n24334 = ~n24293 & n24333 ;
  assign n24335 = ~\pi0625  & ~n24003 ;
  assign n24336 = ~n24002 & n24335 ;
  assign n24337 = \pi1153  & ~n24336 ;
  assign n24338 = ~n24334 & n24337 ;
  assign n24339 = ~n24330 & ~n24338 ;
  assign n24340 = \pi0778  & ~n24339 ;
  assign n24341 = ~n24036 & ~n24322 ;
  assign n24342 = ~n24293 & n24341 ;
  assign n24343 = ~\pi0778  & ~n24342 ;
  assign n24344 = ~n22147 & ~n24343 ;
  assign n24345 = ~n24340 & n24344 ;
  assign n24346 = n22147 & ~n24003 ;
  assign n24347 = ~n24002 & n24346 ;
  assign n24348 = \pi0781  & n23667 ;
  assign n24349 = ~n24347 & n24348 ;
  assign n24350 = ~n24345 & n24349 ;
  assign n24351 = ~n24180 & ~n24350 ;
  assign n24352 = n6861 & ~n24148 ;
  assign n24353 = \pi0142  & ~n21289 ;
  assign n24354 = n1281 & n24144 ;
  assign n24355 = ~n20784 & n23784 ;
  assign n24356 = n1259 & n24355 ;
  assign n24357 = n1249 & n24356 ;
  assign n24358 = n1281 & n24357 ;
  assign n24359 = ~n24354 & ~n24358 ;
  assign n24360 = ~n24353 & n24359 ;
  assign n24361 = ~\pi0039  & n6861 ;
  assign n24362 = ~n24360 & n24361 ;
  assign n24363 = ~n24352 & ~n24362 ;
  assign n24364 = ~n24332 & n24363 ;
  assign n24365 = \pi0142  & ~n22279 ;
  assign n24366 = n22594 & n24365 ;
  assign n24367 = \pi0743  & ~n24366 ;
  assign n24368 = ~\pi0680  & \pi0743  ;
  assign n24369 = ~n22589 & n24368 ;
  assign n24370 = ~n24367 & ~n24369 ;
  assign n24371 = \pi0142  & ~n24370 ;
  assign n24372 = ~n22507 & ~n24370 ;
  assign n24373 = n22505 & n24372 ;
  assign n24374 = ~n24371 & ~n24373 ;
  assign n24375 = \pi0735  & ~n24374 ;
  assign n24376 = ~\pi0142  & ~n22300 ;
  assign n24377 = ~n22314 & n24376 ;
  assign n24378 = \pi0142  & ~n22285 ;
  assign n24379 = n22282 & n24378 ;
  assign n24380 = ~\pi0743  & ~n24379 ;
  assign n24381 = \pi0735  & n24380 ;
  assign n24382 = ~n24377 & n24381 ;
  assign n24383 = ~n24375 & ~n24382 ;
  assign n24384 = ~\pi0735  & ~n24052 ;
  assign n24385 = ~n24049 & n24384 ;
  assign n24386 = ~n2352 & ~n24385 ;
  assign n24387 = n24383 & n24386 ;
  assign n24388 = ~\pi0215  & ~n2352 ;
  assign n24389 = n1689 & n22232 ;
  assign n24390 = n1281 & n24389 ;
  assign n24391 = n1260 & n24390 ;
  assign n24392 = ~n24354 & ~n24391 ;
  assign n24393 = ~n24353 & n24392 ;
  assign n24394 = ~n22532 & ~n24393 ;
  assign n24395 = \pi0735  & ~n24215 ;
  assign n24396 = ~n24394 & n24395 ;
  assign n24397 = ~\pi0735  & ~n24092 ;
  assign n24398 = ~n21285 & n24397 ;
  assign n24399 = n21285 & n24203 ;
  assign n24400 = ~n24398 & ~n24399 ;
  assign n24401 = ~\pi0215  & n24400 ;
  assign n24402 = ~n24396 & n24401 ;
  assign n24403 = ~n24388 & ~n24402 ;
  assign n24404 = ~n21446 & ~n24403 ;
  assign n24405 = ~n24387 & n24404 ;
  assign n24406 = ~n22247 & ~n24250 ;
  assign n24407 = n22180 & ~n22267 ;
  assign n24408 = \pi0142  & ~n24407 ;
  assign n24409 = n24406 & n24408 ;
  assign n24410 = ~\pi0142  & ~n22342 ;
  assign n24411 = ~n22325 & n24410 ;
  assign n24412 = \pi0735  & ~\pi0743  ;
  assign n24413 = ~n24411 & n24412 ;
  assign n24414 = ~n24409 & n24413 ;
  assign n24415 = ~\pi0735  & ~\pi0743  ;
  assign n24416 = \pi0142  & n24415 ;
  assign n24417 = ~n21711 & n24416 ;
  assign n24418 = ~n22473 & n22483 ;
  assign n24419 = ~n22479 & n24418 ;
  assign n24420 = ~\pi0142  & ~n24419 ;
  assign n24421 = \pi0142  & ~n22585 ;
  assign n24422 = n22578 & n24421 ;
  assign n24423 = \pi0735  & \pi0743  ;
  assign n24424 = ~n24422 & n24423 ;
  assign n24425 = ~n24420 & n24424 ;
  assign n24426 = ~\pi0735  & ~n24040 ;
  assign n24427 = n24038 & n24426 ;
  assign n24428 = ~n24425 & ~n24427 ;
  assign n24429 = ~n24417 & n24428 ;
  assign n24430 = ~n24414 & n24429 ;
  assign n24431 = n6732 & ~n24403 ;
  assign n24432 = ~n24430 & n24431 ;
  assign n24433 = ~\pi0142  & ~\pi0743  ;
  assign n24434 = ~\pi0743  & n21627 ;
  assign n24435 = ~n21726 & n24434 ;
  assign n24436 = ~n24433 & ~n24435 ;
  assign n24437 = ~n24061 & ~n24063 ;
  assign n24438 = n24059 & n24437 ;
  assign n24439 = ~\pi0735  & ~n24438 ;
  assign n24440 = n24436 & n24439 ;
  assign n24441 = ~\pi0142  & ~n21516 ;
  assign n24442 = ~\pi0142  & n21403 ;
  assign n24443 = ~n21399 & n24442 ;
  assign n24444 = ~n24441 & ~n24443 ;
  assign n24445 = ~n21527 & ~n24444 ;
  assign n24446 = ~n22458 & n24445 ;
  assign n24447 = \pi0142  & n22549 ;
  assign n24448 = ~n22545 & n24447 ;
  assign n24449 = ~n22540 & n24448 ;
  assign n24450 = \pi0743  & ~n24449 ;
  assign n24451 = ~n24446 & n24450 ;
  assign n24452 = \pi0142  & n21954 ;
  assign n24453 = ~n22201 & n24452 ;
  assign n24454 = ~\pi0142  & ~n22372 ;
  assign n24455 = ~n22371 & n24454 ;
  assign n24456 = ~\pi0743  & ~n24455 ;
  assign n24457 = ~n24453 & n24456 ;
  assign n24458 = ~n24451 & ~n24457 ;
  assign n24459 = \pi0735  & ~n24458 ;
  assign n24460 = ~n6732 & ~n24459 ;
  assign n24461 = ~n24440 & n24460 ;
  assign n24462 = ~\pi0142  & ~n22448 ;
  assign n24463 = \pi0142  & ~n20855 ;
  assign n24464 = n21413 & n24463 ;
  assign n24465 = n21410 & n24463 ;
  assign n24466 = n21392 & n24465 ;
  assign n24467 = ~n24464 & ~n24466 ;
  assign n24468 = \pi0142  & n22563 ;
  assign n24469 = \pi0743  & ~n24468 ;
  assign n24470 = n24467 & n24469 ;
  assign n24471 = \pi0735  & n24470 ;
  assign n24472 = ~n24462 & n24471 ;
  assign n24473 = ~\pi0142  & ~n22357 ;
  assign n24474 = ~n22355 & n24473 ;
  assign n24475 = ~\pi0743  & ~n24474 ;
  assign n24476 = \pi0142  & ~n22205 ;
  assign n24477 = n22204 & n24476 ;
  assign n24478 = \pi0735  & ~n24477 ;
  assign n24479 = \pi0735  & n22227 ;
  assign n24480 = ~n22224 & n24479 ;
  assign n24481 = ~n24478 & ~n24480 ;
  assign n24482 = n24475 & ~n24481 ;
  assign n24483 = ~n24472 & ~n24482 ;
  assign n24484 = n24076 & ~n24080 ;
  assign n24485 = ~\pi0735  & ~n24484 ;
  assign n24486 = ~\pi0735  & n24021 ;
  assign n24487 = ~n21685 & n24486 ;
  assign n24488 = ~n24485 & ~n24487 ;
  assign n24489 = n24483 & n24488 ;
  assign n24490 = n6732 & n24489 ;
  assign n24491 = \pi0215  & ~n24490 ;
  assign n24492 = ~n24461 & n24491 ;
  assign n24493 = ~n24432 & ~n24492 ;
  assign n24494 = ~n24405 & n24493 ;
  assign n24495 = \pi0299  & ~n24494 ;
  assign n24496 = ~n2165 & ~n24385 ;
  assign n24497 = n24383 & n24496 ;
  assign n24498 = ~\pi0223  & n24400 ;
  assign n24499 = ~n24396 & n24498 ;
  assign n24500 = ~n22316 & ~n24499 ;
  assign n24501 = ~n21368 & ~n24500 ;
  assign n24502 = ~n24497 & n24501 ;
  assign n24503 = n6761 & ~n24500 ;
  assign n24504 = ~n24430 & n24503 ;
  assign n24505 = ~n24440 & ~n24459 ;
  assign n24506 = n6764 & ~n24505 ;
  assign n24507 = n21686 & ~n24489 ;
  assign n24508 = ~n24506 & ~n24507 ;
  assign n24509 = \pi0039  & n24508 ;
  assign n24510 = ~n24504 & n24509 ;
  assign n24511 = ~n24502 & n24510 ;
  assign n24512 = ~n2297 & ~n24511 ;
  assign n24513 = ~n24495 & ~n24512 ;
  assign n24514 = \pi0142  & n22649 ;
  assign n24515 = ~n24030 & n24514 ;
  assign n24516 = ~n22686 & n24019 ;
  assign n24517 = ~\pi0299  & ~n24516 ;
  assign n24518 = ~n24515 & n24517 ;
  assign n24519 = ~n22099 & n24009 ;
  assign n24520 = n22005 & n24008 ;
  assign n24521 = \pi0299  & ~n24520 ;
  assign n24522 = ~n24519 & n24521 ;
  assign n24523 = ~n24518 & ~n24522 ;
  assign n24524 = \pi0743  & n24523 ;
  assign n24525 = \pi0142  & ~n21475 ;
  assign n24526 = ~n22006 & n24525 ;
  assign n24527 = ~\pi0142  & ~n22657 ;
  assign n24528 = ~n22660 & n24527 ;
  assign n24529 = n22664 & n24528 ;
  assign n24530 = \pi0299  & ~n24529 ;
  assign n24531 = ~n24526 & n24530 ;
  assign n24532 = ~\pi0743  & n24531 ;
  assign n24533 = \pi0142  & ~n21481 ;
  assign n24534 = ~n21478 & n24533 ;
  assign n24535 = ~n22649 & n24534 ;
  assign n24536 = ~\pi0299  & ~n24535 ;
  assign n24537 = ~\pi0142  & n22676 ;
  assign n24538 = ~\pi0743  & ~n24537 ;
  assign n24539 = n24536 & n24538 ;
  assign n24540 = ~n24532 & ~n24539 ;
  assign n24541 = \pi0735  & n24540 ;
  assign n24542 = ~n24524 & n24541 ;
  assign n24543 = ~\pi0735  & n24034 ;
  assign n24544 = ~\pi0039  & ~n24543 ;
  assign n24545 = ~n24542 & n24544 ;
  assign n24546 = ~n24513 & ~n24545 ;
  assign n24547 = ~\pi0038  & ~n24332 ;
  assign n24548 = ~n24546 & n24547 ;
  assign n24549 = ~n24364 & ~n24548 ;
  assign n24550 = \pi0625  & \pi1153  ;
  assign n24551 = \pi1153  & ~n24152 ;
  assign n24552 = ~n24140 & n24551 ;
  assign n24553 = ~n24550 & ~n24552 ;
  assign n24554 = n24549 & ~n24553 ;
  assign n24555 = \pi0608  & ~n24330 ;
  assign n24556 = ~n24554 & n24555 ;
  assign n24557 = ~n24324 & n24363 ;
  assign n24558 = ~\pi0038  & ~n24324 ;
  assign n24559 = ~n24546 & n24558 ;
  assign n24560 = ~n24557 & ~n24559 ;
  assign n24561 = ~\pi0625  & ~\pi1153  ;
  assign n24562 = ~\pi1153  & ~n24152 ;
  assign n24563 = ~n24140 & n24562 ;
  assign n24564 = ~n24561 & ~n24563 ;
  assign n24565 = n24560 & ~n24564 ;
  assign n24566 = ~\pi0608  & ~n24338 ;
  assign n24567 = ~n24565 & n24566 ;
  assign n24568 = ~n24556 & ~n24567 ;
  assign n24569 = n23673 & ~n24568 ;
  assign n24570 = ~\pi0142  & ~\pi0778  ;
  assign n24571 = ~n23622 & ~n24570 ;
  assign n24572 = n24363 & ~n24571 ;
  assign n24573 = ~\pi0038  & ~n24571 ;
  assign n24574 = ~n24546 & n24573 ;
  assign n24575 = ~n24572 & ~n24574 ;
  assign n24576 = ~\pi0785  & ~n24575 ;
  assign n24577 = n21022 & ~n24576 ;
  assign n24578 = ~n24569 & n24577 ;
  assign n24579 = n24351 & ~n24578 ;
  assign n24580 = n23613 & ~n24568 ;
  assign n24581 = ~\pi0609  & ~n24575 ;
  assign n24582 = \pi0609  & ~n24343 ;
  assign n24583 = ~\pi1155  & ~n24582 ;
  assign n24584 = \pi0778  & ~\pi1155  ;
  assign n24585 = ~n24339 & n24584 ;
  assign n24586 = ~n24583 & ~n24585 ;
  assign n24587 = ~n24581 & ~n24586 ;
  assign n24588 = ~n24580 & n24587 ;
  assign n24589 = n22788 & ~n24152 ;
  assign n24590 = ~n24140 & n24589 ;
  assign n24591 = ~\pi0660  & n22788 ;
  assign n24592 = ~\pi0660  & ~n24003 ;
  assign n24593 = ~n24002 & n24592 ;
  assign n24594 = ~n24591 & ~n24593 ;
  assign n24595 = ~n24590 & ~n24594 ;
  assign n24596 = ~n22787 & ~n24595 ;
  assign n24597 = ~n24588 & ~n24596 ;
  assign n24598 = n23638 & ~n24568 ;
  assign n24599 = \pi0609  & ~n24575 ;
  assign n24600 = ~\pi0609  & ~n24343 ;
  assign n24601 = \pi1155  & ~n24600 ;
  assign n24602 = n22722 & ~n24339 ;
  assign n24603 = ~n24601 & ~n24602 ;
  assign n24604 = ~n24599 & ~n24603 ;
  assign n24605 = ~n24598 & n24604 ;
  assign n24606 = n22767 & ~n24152 ;
  assign n24607 = ~n24140 & n24606 ;
  assign n24608 = \pi0660  & n22767 ;
  assign n24609 = \pi0660  & ~n24003 ;
  assign n24610 = ~n24002 & n24609 ;
  assign n24611 = ~n24608 & ~n24610 ;
  assign n24612 = ~n24607 & ~n24611 ;
  assign n24613 = ~n22766 & ~n24612 ;
  assign n24614 = ~n24605 & ~n24613 ;
  assign n24615 = ~n24597 & ~n24614 ;
  assign n24616 = \pi0785  & n24351 ;
  assign n24617 = ~n24615 & n24616 ;
  assign n24618 = ~n24579 & ~n24617 ;
  assign n24619 = n23729 & n24618 ;
  assign n24620 = n23380 & ~n24343 ;
  assign n24621 = ~n23380 & ~n24003 ;
  assign n24622 = ~n24002 & n24621 ;
  assign n24623 = ~n24620 & ~n24622 ;
  assign n24624 = \pi0778  & ~n24622 ;
  assign n24625 = ~n24339 & n24624 ;
  assign n24626 = ~n24623 & ~n24625 ;
  assign n24627 = n23701 & ~n24626 ;
  assign n24628 = n23683 & ~n24160 ;
  assign n24629 = n21032 & n24166 ;
  assign n24630 = ~n21032 & ~n24003 ;
  assign n24631 = ~n24002 & n24630 ;
  assign n24632 = n22160 & ~n24631 ;
  assign n24633 = ~n24629 & n24632 ;
  assign n24634 = ~n24628 & n24633 ;
  assign n24635 = ~n24627 & ~n24634 ;
  assign n24636 = \pi0626  & ~n24635 ;
  assign n24637 = ~n22160 & ~n24622 ;
  assign n24638 = ~n24620 & n24637 ;
  assign n24639 = \pi0778  & n24637 ;
  assign n24640 = ~n24339 & n24639 ;
  assign n24641 = ~n24638 & ~n24640 ;
  assign n24642 = \pi0641  & ~n22160 ;
  assign n24643 = \pi0641  & ~n24003 ;
  assign n24644 = ~n24002 & n24643 ;
  assign n24645 = ~n24642 & ~n24644 ;
  assign n24646 = n24641 & ~n24645 ;
  assign n24647 = ~n23733 & ~n24646 ;
  assign n24648 = ~n24636 & ~n24647 ;
  assign n24649 = ~n24619 & n24648 ;
  assign n24650 = ~n24178 & ~n24649 ;
  assign n24651 = \pi0626  & ~n24003 ;
  assign n24652 = ~n24002 & n24651 ;
  assign n24653 = ~\pi1158  & ~n24652 ;
  assign n24654 = ~n24169 & n24653 ;
  assign n24655 = ~n24167 & n24654 ;
  assign n24656 = ~n24161 & n24655 ;
  assign n24657 = n20777 & ~n24652 ;
  assign n24658 = \pi0788  & ~n22899 ;
  assign n24659 = ~n24657 & n24658 ;
  assign n24660 = ~n24656 & n24659 ;
  assign n24661 = n23715 & n24618 ;
  assign n24662 = ~\pi0626  & ~n24635 ;
  assign n24663 = \pi0788  & n23719 ;
  assign n24664 = ~\pi0641  & ~n22160 ;
  assign n24665 = ~\pi0641  & ~n24003 ;
  assign n24666 = ~n24002 & n24665 ;
  assign n24667 = ~n24664 & ~n24666 ;
  assign n24668 = \pi0788  & ~n24667 ;
  assign n24669 = n24641 & n24668 ;
  assign n24670 = ~n24663 & ~n24669 ;
  assign n24671 = ~n24662 & ~n24670 ;
  assign n24672 = ~n24661 & n24671 ;
  assign n24673 = ~n24660 & ~n24672 ;
  assign n24674 = ~n24650 & ~n24673 ;
  assign n24675 = ~\pi0788  & ~n24634 ;
  assign n24676 = ~n24627 & n24675 ;
  assign n24677 = ~n23856 & ~n24676 ;
  assign n24678 = n23857 & n24618 ;
  assign n24679 = ~n24677 & ~n24678 ;
  assign n24680 = ~n21067 & ~n24679 ;
  assign n24681 = ~n24674 & n24680 ;
  assign n24682 = ~n24656 & ~n24657 ;
  assign n24683 = ~n24175 & ~n24176 ;
  assign n24684 = n24682 & n24683 ;
  assign n24685 = n21860 & n22166 ;
  assign n24686 = n22932 & n23709 ;
  assign n24687 = ~n24685 & ~n24686 ;
  assign n24688 = ~n24684 & ~n24687 ;
  assign n24689 = ~\pi1156  & ~n22932 ;
  assign n24690 = \pi1156  & ~n22166 ;
  assign n24691 = ~n24689 & ~n24690 ;
  assign n24692 = ~\pi0788  & ~n24169 ;
  assign n24693 = ~n24167 & n24692 ;
  assign n24694 = ~n24161 & n24693 ;
  assign n24695 = n24691 & n24694 ;
  assign n24696 = ~n24688 & ~n24695 ;
  assign n24697 = ~\pi0628  & ~n24003 ;
  assign n24698 = ~n24002 & n24697 ;
  assign n24699 = n20886 & ~n24698 ;
  assign n24700 = n22161 & ~n24003 ;
  assign n24701 = ~n24002 & n24700 ;
  assign n24702 = \pi1156  & ~n24698 ;
  assign n24703 = ~n24701 & n24702 ;
  assign n24704 = ~n24699 & ~n24703 ;
  assign n24705 = ~n22161 & ~n24003 ;
  assign n24706 = ~n24002 & n24705 ;
  assign n24707 = ~n22162 & ~n24706 ;
  assign n24708 = ~n24699 & ~n24707 ;
  assign n24709 = n24641 & n24708 ;
  assign n24710 = ~n24704 & ~n24709 ;
  assign n24711 = ~\pi0629  & n24710 ;
  assign n24712 = \pi0628  & ~n24003 ;
  assign n24713 = ~n24002 & n24712 ;
  assign n24714 = n20887 & ~n24713 ;
  assign n24715 = ~\pi1156  & ~n24713 ;
  assign n24716 = ~n24701 & n24715 ;
  assign n24717 = ~n24714 & ~n24716 ;
  assign n24718 = ~n24707 & ~n24714 ;
  assign n24719 = n24641 & n24718 ;
  assign n24720 = ~n24717 & ~n24719 ;
  assign n24721 = \pi0629  & n24720 ;
  assign n24722 = ~n24711 & ~n24721 ;
  assign n24723 = n24696 & n24722 ;
  assign n24724 = \pi0792  & ~n21067 ;
  assign n24725 = ~n24723 & n24724 ;
  assign n24726 = n24641 & ~n24707 ;
  assign n24727 = ~\pi0792  & ~n24701 ;
  assign n24728 = ~n24726 & n24727 ;
  assign n24729 = ~\pi0647  & n24728 ;
  assign n24730 = ~n24710 & ~n24720 ;
  assign n24731 = n22913 & ~n24730 ;
  assign n24732 = ~n24729 & ~n24731 ;
  assign n24733 = ~n24002 & ~n24003 ;
  assign n24734 = \pi0647  & ~n24733 ;
  assign n24735 = n24732 & ~n24734 ;
  assign n24736 = n20897 & ~n24735 ;
  assign n24737 = \pi0788  & ~n20846 ;
  assign n24738 = ~n24684 & n24737 ;
  assign n24739 = ~\pi0788  & ~n20846 ;
  assign n24740 = ~n24169 & n24739 ;
  assign n24741 = ~n24167 & n24740 ;
  assign n24742 = ~n24161 & n24741 ;
  assign n24743 = n20846 & ~n24733 ;
  assign n24744 = ~n24742 & ~n24743 ;
  assign n24745 = ~n24738 & n24744 ;
  assign n24746 = ~n20910 & ~n24745 ;
  assign n24747 = \pi0647  & ~n24727 ;
  assign n24748 = \pi0647  & ~n24707 ;
  assign n24749 = n24641 & n24748 ;
  assign n24750 = ~n24747 & ~n24749 ;
  assign n24751 = ~\pi0647  & ~n24003 ;
  assign n24752 = ~n24002 & n24751 ;
  assign n24753 = n20849 & ~n24752 ;
  assign n24754 = n24750 & n24753 ;
  assign n24755 = \pi0792  & n24753 ;
  assign n24756 = ~n24730 & n24755 ;
  assign n24757 = ~n24754 & ~n24756 ;
  assign n24758 = ~n24746 & n24757 ;
  assign n24759 = ~n24736 & n24758 ;
  assign n24760 = \pi0787  & ~n24759 ;
  assign n24761 = \pi0790  & ~n23318 ;
  assign n24762 = n6848 & ~n24761 ;
  assign n24763 = ~n24760 & n24762 ;
  assign n24764 = ~n24725 & n24763 ;
  assign n24765 = ~n24681 & n24764 ;
  assign n24766 = ~n21088 & n23413 ;
  assign n24767 = ~n20846 & n24766 ;
  assign n24768 = ~n24003 & n24766 ;
  assign n24769 = ~n24002 & n24768 ;
  assign n24770 = ~n24767 & ~n24769 ;
  assign n24771 = ~n24742 & ~n24770 ;
  assign n24772 = ~n24738 & n24771 ;
  assign n24773 = n23412 & ~n24003 ;
  assign n24774 = ~n24002 & n24773 ;
  assign n24775 = ~n24772 & ~n24774 ;
  assign n24776 = ~\pi0644  & ~n24775 ;
  assign n24777 = n21088 & ~n23414 ;
  assign n24778 = ~n24003 & n24777 ;
  assign n24779 = ~n24002 & n24778 ;
  assign n24780 = ~\pi0644  & ~n24779 ;
  assign n24781 = ~n21088 & n23412 ;
  assign n24782 = ~n20846 & n24781 ;
  assign n24783 = ~n24003 & n24781 ;
  assign n24784 = ~n24002 & n24783 ;
  assign n24785 = ~n24782 & ~n24784 ;
  assign n24786 = ~n24742 & ~n24785 ;
  assign n24787 = ~n24738 & n24786 ;
  assign n24788 = n23413 & ~n24003 ;
  assign n24789 = ~n24002 & n24788 ;
  assign n24790 = ~n24779 & ~n24789 ;
  assign n24791 = ~n24787 & n24790 ;
  assign n24792 = ~n24780 & ~n24791 ;
  assign n24793 = ~n24776 & ~n24792 ;
  assign n24794 = \pi0790  & ~n24793 ;
  assign n24795 = \pi0787  & ~\pi1157  ;
  assign n24796 = ~n24735 & n24795 ;
  assign n24797 = \pi1157  & ~n24752 ;
  assign n24798 = \pi0787  & n24750 ;
  assign n24799 = \pi0787  & \pi0792  ;
  assign n24800 = ~n24730 & n24799 ;
  assign n24801 = ~n24798 & ~n24800 ;
  assign n24802 = n24797 & ~n24801 ;
  assign n24803 = ~\pi0787  & n24728 ;
  assign n24804 = n23011 & ~n24730 ;
  assign n24805 = ~n24803 & ~n24804 ;
  assign n24806 = \pi0790  & ~n23517 ;
  assign n24807 = ~n23516 & n24806 ;
  assign n24808 = n24805 & n24807 ;
  assign n24809 = ~n24802 & n24808 ;
  assign n24810 = ~n24796 & n24809 ;
  assign n24811 = ~n24794 & ~n24810 ;
  assign n24812 = n6848 & ~n24811 ;
  assign n24813 = ~\pi0142  & ~n6848 ;
  assign n24814 = ~\pi0057  & ~n24813 ;
  assign n24815 = ~n23932 & n24814 ;
  assign n24816 = \pi0790  & n24814 ;
  assign n24817 = ~n23971 & n24816 ;
  assign n24818 = ~n24815 & ~n24817 ;
  assign n24819 = ~n24812 & ~n24818 ;
  assign n24820 = ~n24765 & n24819 ;
  assign n24821 = n23974 & ~n24820 ;
  assign n24822 = \pi0143  & ~\pi0832  ;
  assign n24823 = ~n21132 & ~n24822 ;
  assign n24824 = \pi0687  & n1689 ;
  assign n24825 = n20855 & n24824 ;
  assign n24826 = ~n20861 & n24825 ;
  assign n24827 = ~\pi0143  & ~n1689 ;
  assign n24828 = ~n24826 & ~n24827 ;
  assign n24829 = n20879 & ~n24828 ;
  assign n24830 = \pi0647  & n20891 ;
  assign n24831 = n24829 & n24830 ;
  assign n24832 = ~\pi0143  & ~\pi0647  ;
  assign n24833 = ~n1689 & n24832 ;
  assign n24834 = \pi1157  & ~n24833 ;
  assign n24835 = ~n24831 & n24834 ;
  assign n24836 = n20895 & n24829 ;
  assign n24837 = ~\pi0143  & \pi0647  ;
  assign n24838 = ~n1689 & n24837 ;
  assign n24839 = ~\pi1157  & ~n24838 ;
  assign n24840 = ~n24836 & n24839 ;
  assign n24841 = ~n24835 & ~n24840 ;
  assign n24842 = \pi0787  & ~n24841 ;
  assign n24843 = \pi0787  & \pi1160  ;
  assign n24844 = \pi1160  & n20891 ;
  assign n24845 = n24829 & n24844 ;
  assign n24846 = ~n24843 & ~n24845 ;
  assign n24847 = n23313 & ~n24846 ;
  assign n24848 = ~n24842 & n24847 ;
  assign n24849 = ~n21032 & ~n24827 ;
  assign n24850 = \pi0789  & n24849 ;
  assign n24851 = ~\pi0788  & ~n24850 ;
  assign n24852 = n23423 & n24851 ;
  assign n24853 = ~\pi0774  & n1689 ;
  assign n24854 = n20784 & n24853 ;
  assign n24855 = ~n24827 & ~n24854 ;
  assign n24856 = n20794 & ~n24855 ;
  assign n24857 = n20796 & ~n24856 ;
  assign n24858 = n20799 & ~n24855 ;
  assign n24859 = n20801 & ~n24858 ;
  assign n24860 = ~n24857 & ~n24859 ;
  assign n24861 = ~\pi0785  & ~n24827 ;
  assign n24862 = ~n24854 & n24861 ;
  assign n24863 = ~n20804 & ~n24862 ;
  assign n24864 = ~n20812 & n24863 ;
  assign n24865 = n24851 & n24864 ;
  assign n24866 = n24860 & n24865 ;
  assign n24867 = ~n24852 & ~n24866 ;
  assign n24868 = ~n20846 & ~n24867 ;
  assign n24869 = ~n20778 & n24827 ;
  assign n24870 = n24737 & n24869 ;
  assign n24871 = n23423 & ~n24850 ;
  assign n24872 = ~n24850 & n24864 ;
  assign n24873 = n24860 & n24872 ;
  assign n24874 = ~n24871 & ~n24873 ;
  assign n24875 = n20778 & n24737 ;
  assign n24876 = ~n24874 & n24875 ;
  assign n24877 = ~n24870 & ~n24876 ;
  assign n24878 = ~n24868 & n24877 ;
  assign n24879 = ~\pi1160  & n23313 ;
  assign n24880 = ~n21088 & n24879 ;
  assign n24881 = ~n24878 & n24880 ;
  assign n24882 = ~n24848 & ~n24881 ;
  assign n24883 = \pi1160  & n23312 ;
  assign n24884 = ~n21088 & n24883 ;
  assign n24885 = ~n24878 & n24884 ;
  assign n24886 = ~n20846 & n23415 ;
  assign n24887 = ~n23414 & n24827 ;
  assign n24888 = ~n24886 & n24887 ;
  assign n24889 = n20891 & n24829 ;
  assign n24890 = ~\pi0787  & ~n24889 ;
  assign n24891 = ~\pi1160  & n23312 ;
  assign n24892 = ~n24890 & n24891 ;
  assign n24893 = ~n24842 & n24892 ;
  assign n24894 = ~n24888 & ~n24893 ;
  assign n24895 = ~n24885 & n24894 ;
  assign n24896 = n24882 & n24895 ;
  assign n24897 = \pi0790  & ~n24896 ;
  assign n24898 = n24823 & n24897 ;
  assign n24899 = \pi0788  & n24869 ;
  assign n24900 = n20816 & ~n24874 ;
  assign n24901 = ~n24899 & ~n24900 ;
  assign n24902 = n24691 & n24867 ;
  assign n24903 = n24901 & n24902 ;
  assign n24904 = ~n20885 & ~n21075 ;
  assign n24905 = n24829 & n24904 ;
  assign n24906 = n20843 & ~n24905 ;
  assign n24907 = ~n20878 & ~n20936 ;
  assign n24908 = n20873 & n24907 ;
  assign n24909 = ~n24828 & n24908 ;
  assign n24910 = ~n20885 & n24909 ;
  assign n24911 = n20844 & ~n24910 ;
  assign n24912 = ~n24906 & ~n24911 ;
  assign n24913 = ~n24903 & n24912 ;
  assign n24914 = \pi0792  & ~n24913 ;
  assign n24915 = n20855 & ~n20861 ;
  assign n24916 = \pi0687  & ~n20784 ;
  assign n24917 = \pi0687  & ~n20790 ;
  assign n24918 = n20789 & n24917 ;
  assign n24919 = ~n24916 & ~n24918 ;
  assign n24920 = n24915 & ~n24919 ;
  assign n24921 = \pi0603  & ~\pi0774  ;
  assign n24922 = ~n20783 & n24921 ;
  assign n24923 = ~n20985 & n24922 ;
  assign n24924 = ~n24827 & ~n24923 ;
  assign n24925 = ~n24920 & n24924 ;
  assign n24926 = \pi0143  & ~n1689 ;
  assign n24927 = ~\pi0609  & ~n24926 ;
  assign n24928 = ~n24925 & n24927 ;
  assign n24929 = ~\pi1155  & ~n24827 ;
  assign n24930 = ~n24826 & n24929 ;
  assign n24931 = ~n20999 & ~n24930 ;
  assign n24932 = ~n24928 & ~n24931 ;
  assign n24933 = \pi1155  & ~n24858 ;
  assign n24934 = ~\pi0660  & ~n24933 ;
  assign n24935 = ~n24932 & n24934 ;
  assign n24936 = ~n21007 & ~n24857 ;
  assign n24937 = \pi0609  & ~n24926 ;
  assign n24938 = ~n24925 & n24937 ;
  assign n24939 = ~\pi0609  & ~n24828 ;
  assign n24940 = n20801 & ~n24939 ;
  assign n24941 = ~n24938 & n24940 ;
  assign n24942 = n24936 & ~n24941 ;
  assign n24943 = ~n24935 & ~n24942 ;
  assign n24944 = ~n24925 & ~n24926 ;
  assign n24945 = ~\pi0785  & ~n24944 ;
  assign n24946 = n21022 & ~n24945 ;
  assign n24947 = ~n24943 & n24946 ;
  assign n24948 = n20964 & n24863 ;
  assign n24949 = n24860 & n24948 ;
  assign n24950 = \pi0627  & ~n24827 ;
  assign n24951 = ~n24826 & n24950 ;
  assign n24952 = ~n20968 & ~n24951 ;
  assign n24953 = ~n24949 & ~n24952 ;
  assign n24954 = ~\pi0627  & ~n24827 ;
  assign n24955 = ~n24826 & n24954 ;
  assign n24956 = ~n20978 & ~n24955 ;
  assign n24957 = \pi0781  & n24956 ;
  assign n24958 = n20974 & n24863 ;
  assign n24959 = \pi0781  & n24958 ;
  assign n24960 = n24860 & n24959 ;
  assign n24961 = ~n24957 & ~n24960 ;
  assign n24962 = ~n24953 & ~n24961 ;
  assign n24963 = ~n21034 & ~n24962 ;
  assign n24964 = ~n24947 & n24963 ;
  assign n24965 = n21050 & ~n24827 ;
  assign n24966 = ~n24826 & n24965 ;
  assign n24967 = ~n21051 & ~n24966 ;
  assign n24968 = ~n20876 & n24849 ;
  assign n24969 = ~n20876 & n21032 ;
  assign n24970 = ~n24968 & ~n24969 ;
  assign n24971 = n24864 & ~n24968 ;
  assign n24972 = n24860 & n24971 ;
  assign n24973 = ~n24970 & ~n24972 ;
  assign n24974 = n24967 & ~n24973 ;
  assign n24975 = \pi0789  & ~n24974 ;
  assign n24976 = ~n21038 & ~n24975 ;
  assign n24977 = ~n24964 & n24976 ;
  assign n24978 = n20778 & ~n24874 ;
  assign n24979 = n23170 & ~n24828 ;
  assign n24980 = ~n24869 & ~n24979 ;
  assign n24981 = ~n24978 & n24980 ;
  assign n24982 = n20883 & ~n24979 ;
  assign n24983 = \pi0788  & ~n24982 ;
  assign n24984 = ~n24981 & n24983 ;
  assign n24985 = ~n23856 & ~n24984 ;
  assign n24986 = ~n24977 & n24985 ;
  assign n24987 = ~n24914 & ~n24986 ;
  assign n24988 = \pi0832  & ~n21067 ;
  assign n24989 = ~n24987 & n24988 ;
  assign n24990 = ~\pi0143  & \pi0792  ;
  assign n24991 = ~n1689 & n24990 ;
  assign n24992 = ~n20845 & n24991 ;
  assign n24993 = n20908 & n24795 ;
  assign n24994 = \pi0787  & \pi1157  ;
  assign n24995 = n20906 & n24994 ;
  assign n24996 = ~n24993 & ~n24995 ;
  assign n24997 = ~n24992 & ~n24996 ;
  assign n24998 = ~n24868 & n24997 ;
  assign n24999 = n24877 & n24998 ;
  assign n25000 = \pi0630  & n24839 ;
  assign n25001 = ~n24836 & n25000 ;
  assign n25002 = n20849 & ~n24833 ;
  assign n25003 = ~n24831 & n25002 ;
  assign n25004 = ~n25001 & ~n25003 ;
  assign n25005 = \pi0787  & ~n25004 ;
  assign n25006 = ~n24761 & ~n25005 ;
  assign n25007 = ~n24999 & n25006 ;
  assign n25008 = \pi0832  & ~n25007 ;
  assign n25009 = n24823 & ~n25008 ;
  assign n25010 = ~n24989 & n25009 ;
  assign n25011 = ~n24898 & ~n25010 ;
  assign n25012 = ~\pi0143  & n21770 ;
  assign n25013 = ~n21734 & n25012 ;
  assign n25014 = ~\pi0143  & n21768 ;
  assign n25015 = ~n25013 & ~n25014 ;
  assign n25016 = ~n21777 & n25015 ;
  assign n25017 = ~\pi0781  & n25016 ;
  assign n25018 = \pi0143  & ~n6861 ;
  assign n25019 = ~\pi0143  & n22124 ;
  assign n25020 = ~n25013 & ~n25019 ;
  assign n25021 = \pi0774  & n25020 ;
  assign n25022 = n6861 & n25021 ;
  assign n25023 = n21484 & ~n21566 ;
  assign n25024 = ~\pi0038  & n25023 ;
  assign n25025 = \pi0143  & ~n25024 ;
  assign n25026 = ~\pi0039  & n21272 ;
  assign n25027 = ~\pi0038  & n21467 ;
  assign n25028 = ~n25026 & n25027 ;
  assign n25029 = ~\pi0143  & ~\pi0774  ;
  assign n25030 = n8413 & n21417 ;
  assign n25031 = n1354 & n25030 ;
  assign n25032 = n1358 & n25031 ;
  assign n25033 = \pi0038  & ~n25032 ;
  assign n25034 = n25029 & ~n25033 ;
  assign n25035 = ~n25028 & n25034 ;
  assign n25036 = ~n25025 & ~n25035 ;
  assign n25037 = \pi0038  & n1689 ;
  assign n25038 = n4520 & n25037 ;
  assign n25039 = n1638 & n25038 ;
  assign n25040 = n20784 & n25039 ;
  assign n25041 = n6861 & ~n25040 ;
  assign n25042 = ~n25036 & n25041 ;
  assign n25043 = ~n25022 & ~n25042 ;
  assign n25044 = ~n25018 & n25043 ;
  assign n25045 = n24162 & ~n25044 ;
  assign n25046 = ~n25017 & ~n25045 ;
  assign n25047 = ~\pi0789  & ~n25046 ;
  assign n25048 = \pi0618  & ~n25016 ;
  assign n25049 = ~n21777 & n25048 ;
  assign n25050 = ~n25018 & n25048 ;
  assign n25051 = n25043 & n25050 ;
  assign n25052 = ~n25049 & ~n25051 ;
  assign n25053 = ~\pi0143  & ~\pi0618  ;
  assign n25054 = n21768 & n25053 ;
  assign n25055 = n21770 & n25053 ;
  assign n25056 = ~n21734 & n25055 ;
  assign n25057 = ~n25054 & ~n25056 ;
  assign n25058 = \pi1154  & n25057 ;
  assign n25059 = n25052 & n25058 ;
  assign n25060 = ~\pi0618  & ~n25016 ;
  assign n25061 = ~n21777 & n25060 ;
  assign n25062 = ~n25018 & n25060 ;
  assign n25063 = n25043 & n25062 ;
  assign n25064 = ~n25061 & ~n25063 ;
  assign n25065 = ~\pi0143  & \pi0618  ;
  assign n25066 = n21768 & n25065 ;
  assign n25067 = n21770 & n25065 ;
  assign n25068 = ~n21734 & n25067 ;
  assign n25069 = ~n25066 & ~n25068 ;
  assign n25070 = ~\pi1154  & n25069 ;
  assign n25071 = n25064 & n25070 ;
  assign n25072 = ~n25059 & ~n25071 ;
  assign n25073 = n21806 & ~n25072 ;
  assign n25074 = ~n25047 & ~n25073 ;
  assign n25075 = ~\pi0788  & ~n25074 ;
  assign n25076 = ~\pi0619  & n25046 ;
  assign n25077 = ~\pi0143  & \pi0619  ;
  assign n25078 = n21768 & n25077 ;
  assign n25079 = n21770 & n25077 ;
  assign n25080 = ~n21734 & n25079 ;
  assign n25081 = ~n25078 & ~n25080 ;
  assign n25082 = ~\pi1159  & n25081 ;
  assign n25083 = ~n25076 & n25082 ;
  assign n25084 = \pi0781  & n25082 ;
  assign n25085 = ~n25072 & n25084 ;
  assign n25086 = ~n25083 & ~n25085 ;
  assign n25087 = \pi0619  & n25046 ;
  assign n25088 = ~\pi0143  & ~\pi0619  ;
  assign n25089 = n21768 & n25088 ;
  assign n25090 = n21770 & n25088 ;
  assign n25091 = ~n21734 & n25090 ;
  assign n25092 = ~n25089 & ~n25091 ;
  assign n25093 = \pi1159  & n25092 ;
  assign n25094 = ~n25087 & n25093 ;
  assign n25095 = \pi0781  & n25093 ;
  assign n25096 = ~n25072 & n25095 ;
  assign n25097 = ~n25094 & ~n25096 ;
  assign n25098 = n25086 & n25097 ;
  assign n25099 = n21832 & ~n25098 ;
  assign n25100 = ~n25075 & ~n25099 ;
  assign n25101 = ~\pi0628  & n25100 ;
  assign n25102 = \pi1156  & ~n25101 ;
  assign n25103 = ~\pi0626  & n25074 ;
  assign n25104 = ~\pi0143  & \pi0626  ;
  assign n25105 = n21768 & n25104 ;
  assign n25106 = n21770 & n25104 ;
  assign n25107 = ~n21734 & n25106 ;
  assign n25108 = ~n25105 & ~n25107 ;
  assign n25109 = ~\pi1158  & n25108 ;
  assign n25110 = ~n25103 & n25109 ;
  assign n25111 = \pi0789  & n25109 ;
  assign n25112 = ~n25098 & n25111 ;
  assign n25113 = ~n25110 & ~n25112 ;
  assign n25114 = \pi0626  & n25074 ;
  assign n25115 = ~\pi0143  & ~\pi0626  ;
  assign n25116 = n21768 & n25115 ;
  assign n25117 = n21770 & n25115 ;
  assign n25118 = ~n21734 & n25117 ;
  assign n25119 = ~n25116 & ~n25118 ;
  assign n25120 = \pi1158  & n25119 ;
  assign n25121 = ~n25114 & n25120 ;
  assign n25122 = \pi0789  & n25120 ;
  assign n25123 = ~n25098 & n25122 ;
  assign n25124 = ~n25121 & ~n25123 ;
  assign n25125 = n25113 & n25124 ;
  assign n25126 = n21860 & ~n25125 ;
  assign n25127 = ~n25102 & ~n25126 ;
  assign n25128 = ~\pi0143  & \pi0628  ;
  assign n25129 = n21768 & n25128 ;
  assign n25130 = n21770 & n25128 ;
  assign n25131 = ~n21734 & n25130 ;
  assign n25132 = ~n25129 & ~n25131 ;
  assign n25133 = ~\pi1156  & n25132 ;
  assign n25134 = \pi0629  & ~n25133 ;
  assign n25135 = ~\pi0143  & ~\pi0625  ;
  assign n25136 = ~n22734 & ~n25135 ;
  assign n25137 = ~\pi0143  & \pi0625  ;
  assign n25138 = n21768 & n25137 ;
  assign n25139 = n21770 & n25137 ;
  assign n25140 = ~n21734 & n25139 ;
  assign n25141 = ~n25138 & ~n25140 ;
  assign n25142 = ~\pi1153  & n25141 ;
  assign n25143 = n25136 & n25142 ;
  assign n25144 = ~\pi0143  & ~n22017 ;
  assign n25145 = ~n21994 & n25144 ;
  assign n25146 = ~\pi0038  & ~\pi0143  ;
  assign n25147 = ~n22109 & ~n25146 ;
  assign n25148 = ~n25145 & ~n25147 ;
  assign n25149 = ~\pi0143  & ~n21757 ;
  assign n25150 = n22117 & ~n25149 ;
  assign n25151 = \pi0687  & ~n25150 ;
  assign n25152 = ~n25148 & n25151 ;
  assign n25153 = ~\pi0687  & ~n25020 ;
  assign n25154 = ~n25152 & ~n25153 ;
  assign n25155 = n6861 & n25142 ;
  assign n25156 = n25154 & n25155 ;
  assign n25157 = ~n25143 & ~n25156 ;
  assign n25158 = ~n22727 & ~n25137 ;
  assign n25159 = n21768 & n25135 ;
  assign n25160 = n21770 & n25135 ;
  assign n25161 = ~n21734 & n25160 ;
  assign n25162 = ~n25159 & ~n25161 ;
  assign n25163 = \pi1153  & n25162 ;
  assign n25164 = n25158 & n25163 ;
  assign n25165 = n6861 & n25163 ;
  assign n25166 = n25154 & n25165 ;
  assign n25167 = ~n25164 & ~n25166 ;
  assign n25168 = n25157 & n25167 ;
  assign n25169 = n22148 & ~n25168 ;
  assign n25170 = ~\pi0778  & n25018 ;
  assign n25171 = ~\pi0778  & n6861 ;
  assign n25172 = n25154 & n25171 ;
  assign n25173 = ~n25170 & ~n25172 ;
  assign n25174 = ~n22147 & ~n25173 ;
  assign n25175 = n22147 & n25015 ;
  assign n25176 = ~n22155 & ~n25175 ;
  assign n25177 = ~n25174 & n25176 ;
  assign n25178 = ~n25169 & n25177 ;
  assign n25179 = n22155 & ~n25015 ;
  assign n25180 = n22162 & ~n25179 ;
  assign n25181 = ~n25178 & n25180 ;
  assign n25182 = ~n22162 & n25015 ;
  assign n25183 = n22166 & ~n25182 ;
  assign n25184 = ~n25181 & n25183 ;
  assign n25185 = ~n25134 & ~n25184 ;
  assign n25186 = n25127 & ~n25185 ;
  assign n25187 = n1281 & n12800 ;
  assign n25188 = n22535 & n25187 ;
  assign n25189 = ~\pi0039  & ~n25188 ;
  assign n25190 = ~n22683 & n25189 ;
  assign n25191 = \pi0038  & ~n25188 ;
  assign n25192 = n23548 & ~n25191 ;
  assign n25193 = ~n25190 & n25192 ;
  assign n25194 = ~\pi0143  & ~n25193 ;
  assign n25195 = \pi0038  & ~n22708 ;
  assign n25196 = \pi0143  & ~n25195 ;
  assign n25197 = \pi0038  & n25196 ;
  assign n25198 = ~n23558 & n25196 ;
  assign n25199 = n23557 & n25198 ;
  assign n25200 = ~n25197 & ~n25199 ;
  assign n25201 = ~n25194 & n25200 ;
  assign n25202 = ~\pi0774  & n25201 ;
  assign n25203 = ~\pi0038  & ~n23567 ;
  assign n25204 = n23565 & n25203 ;
  assign n25205 = n21754 & ~n22232 ;
  assign n25206 = n1266 & n25205 ;
  assign n25207 = \pi0038  & n1354 ;
  assign n25208 = n25206 & n25207 ;
  assign n25209 = n1358 & n25208 ;
  assign n25210 = ~\pi0143  & ~n25209 ;
  assign n25211 = ~n25204 & n25210 ;
  assign n25212 = ~\pi0038  & \pi0143  ;
  assign n25213 = n23575 & n25212 ;
  assign n25214 = n23572 & n25213 ;
  assign n25215 = n12800 & n24389 ;
  assign n25216 = n1281 & n25215 ;
  assign n25217 = n1260 & n25216 ;
  assign n25218 = \pi0774  & ~n25217 ;
  assign n25219 = ~n25214 & n25218 ;
  assign n25220 = ~n25211 & n25219 ;
  assign n25221 = \pi0687  & ~n25220 ;
  assign n25222 = ~n25202 & n25221 ;
  assign n25223 = ~\pi0687  & n25040 ;
  assign n25224 = ~\pi0687  & ~n25025 ;
  assign n25225 = ~n25035 & n25224 ;
  assign n25226 = ~n25223 & ~n25225 ;
  assign n25227 = ~n25021 & ~n25226 ;
  assign n25228 = n6861 & ~n25227 ;
  assign n25229 = ~n25222 & n25228 ;
  assign n25230 = \pi0609  & ~n25018 ;
  assign n25231 = ~n25229 & n25230 ;
  assign n25232 = ~n23638 & ~n25231 ;
  assign n25233 = ~\pi0609  & n25173 ;
  assign n25234 = \pi1155  & ~n25233 ;
  assign n25235 = n22722 & ~n25168 ;
  assign n25236 = ~n25234 & ~n25235 ;
  assign n25237 = n25232 & ~n25236 ;
  assign n25238 = ~n25158 & ~n25229 ;
  assign n25239 = n25043 & ~n25136 ;
  assign n25240 = \pi1153  & ~n25239 ;
  assign n25241 = ~n25238 & n25240 ;
  assign n25242 = \pi0608  & n25157 ;
  assign n25243 = ~n25241 & n25242 ;
  assign n25244 = ~n25136 & ~n25229 ;
  assign n25245 = n25043 & ~n25158 ;
  assign n25246 = ~\pi1153  & ~n25245 ;
  assign n25247 = ~n25244 & n25246 ;
  assign n25248 = ~\pi0608  & n25167 ;
  assign n25249 = ~n25247 & n25248 ;
  assign n25250 = ~n25243 & ~n25249 ;
  assign n25251 = \pi0778  & ~n25236 ;
  assign n25252 = n25250 & n25251 ;
  assign n25253 = ~n25237 & ~n25252 ;
  assign n25254 = ~n22767 & n25015 ;
  assign n25255 = \pi0660  & ~n25254 ;
  assign n25256 = ~n22767 & n25255 ;
  assign n25257 = ~n25018 & n25255 ;
  assign n25258 = n25043 & n25257 ;
  assign n25259 = ~n25256 & ~n25258 ;
  assign n25260 = ~n22766 & n25259 ;
  assign n25261 = n25253 & ~n25260 ;
  assign n25262 = n22776 & n25261 ;
  assign n25263 = ~\pi0609  & ~n25018 ;
  assign n25264 = ~n25229 & n25263 ;
  assign n25265 = ~n23613 & ~n25264 ;
  assign n25266 = \pi0778  & ~n25168 ;
  assign n25267 = \pi0609  & n25173 ;
  assign n25268 = ~n25266 & n25267 ;
  assign n25269 = n25265 & ~n25268 ;
  assign n25270 = \pi0778  & ~n25268 ;
  assign n25271 = n25250 & n25270 ;
  assign n25272 = ~n25269 & ~n25271 ;
  assign n25273 = ~\pi1155  & ~n25272 ;
  assign n25274 = ~n22788 & n25015 ;
  assign n25275 = ~\pi0660  & ~n25274 ;
  assign n25276 = ~n22788 & n25275 ;
  assign n25277 = ~n25018 & n25275 ;
  assign n25278 = n25043 & n25277 ;
  assign n25279 = ~n25276 & ~n25278 ;
  assign n25280 = ~n22787 & n25279 ;
  assign n25281 = n22776 & ~n25280 ;
  assign n25282 = ~n25273 & n25281 ;
  assign n25283 = ~n25262 & ~n25282 ;
  assign n25284 = \pi0778  & n25250 ;
  assign n25285 = ~\pi0785  & ~n25018 ;
  assign n25286 = ~n25229 & n25285 ;
  assign n25287 = ~n23673 & ~n25286 ;
  assign n25288 = ~\pi0618  & ~n25287 ;
  assign n25289 = ~n25284 & n25288 ;
  assign n25290 = \pi0618  & ~n25175 ;
  assign n25291 = ~n25174 & n25290 ;
  assign n25292 = ~n25169 & n25291 ;
  assign n25293 = ~\pi1154  & ~n25292 ;
  assign n25294 = ~n25289 & n25293 ;
  assign n25295 = n25283 & n25294 ;
  assign n25296 = ~\pi0627  & ~n25059 ;
  assign n25297 = ~n25295 & n25296 ;
  assign n25298 = n22816 & n25261 ;
  assign n25299 = n22816 & ~n25280 ;
  assign n25300 = ~n25273 & n25299 ;
  assign n25301 = ~n25298 & ~n25300 ;
  assign n25302 = \pi0618  & ~n25287 ;
  assign n25303 = ~n25284 & n25302 ;
  assign n25304 = ~\pi0618  & ~n25175 ;
  assign n25305 = ~n25174 & n25304 ;
  assign n25306 = ~n25169 & n25305 ;
  assign n25307 = \pi1154  & ~n25306 ;
  assign n25308 = ~n25303 & n25307 ;
  assign n25309 = n25301 & n25308 ;
  assign n25310 = \pi0627  & ~n25071 ;
  assign n25311 = ~n25309 & n25310 ;
  assign n25312 = ~n25297 & ~n25311 ;
  assign n25313 = n21806 & ~n25312 ;
  assign n25314 = ~\pi0781  & ~n25287 ;
  assign n25315 = ~n25284 & n25314 ;
  assign n25316 = n22840 & n25261 ;
  assign n25317 = n22840 & ~n25280 ;
  assign n25318 = ~n25273 & n25317 ;
  assign n25319 = ~n25316 & ~n25318 ;
  assign n25320 = ~n25315 & n25319 ;
  assign n25321 = ~\pi0789  & ~n25320 ;
  assign n25322 = \pi0626  & ~n25321 ;
  assign n25323 = ~n25313 & n25322 ;
  assign n25324 = ~n22849 & n25015 ;
  assign n25325 = ~\pi0626  & n25324 ;
  assign n25326 = ~n25174 & ~n25175 ;
  assign n25327 = ~n25169 & n25326 ;
  assign n25328 = n22854 & ~n25327 ;
  assign n25329 = ~n25325 & ~n25328 ;
  assign n25330 = \pi0641  & n25329 ;
  assign n25331 = ~n25323 & n25330 ;
  assign n25332 = n22859 & ~n25312 ;
  assign n25333 = \pi0619  & ~n25320 ;
  assign n25334 = \pi1159  & ~n25179 ;
  assign n25335 = ~n25178 & n25334 ;
  assign n25336 = ~n20830 & ~n25335 ;
  assign n25337 = ~n25333 & ~n25336 ;
  assign n25338 = ~n25332 & n25337 ;
  assign n25339 = \pi0648  & n25086 ;
  assign n25340 = ~n25338 & n25339 ;
  assign n25341 = n22869 & ~n25312 ;
  assign n25342 = ~\pi0619  & ~n25320 ;
  assign n25343 = ~\pi1159  & ~n25179 ;
  assign n25344 = ~n25178 & n25343 ;
  assign n25345 = ~n22872 & ~n25344 ;
  assign n25346 = ~n25342 & ~n25345 ;
  assign n25347 = ~n25341 & n25346 ;
  assign n25348 = ~\pi0648  & n25097 ;
  assign n25349 = ~n25347 & n25348 ;
  assign n25350 = ~n25340 & ~n25349 ;
  assign n25351 = \pi0789  & n25330 ;
  assign n25352 = ~n25350 & n25351 ;
  assign n25353 = ~n25331 & ~n25352 ;
  assign n25354 = ~n22884 & n25124 ;
  assign n25355 = n25353 & ~n25354 ;
  assign n25356 = \pi0788  & n25355 ;
  assign n25357 = ~\pi0626  & ~n25321 ;
  assign n25358 = ~n25313 & n25357 ;
  assign n25359 = \pi0626  & n25324 ;
  assign n25360 = n22891 & ~n25327 ;
  assign n25361 = ~n25359 & ~n25360 ;
  assign n25362 = ~n25358 & n25361 ;
  assign n25363 = \pi0789  & n25361 ;
  assign n25364 = ~n25350 & n25363 ;
  assign n25365 = ~n25362 & ~n25364 ;
  assign n25366 = ~\pi0641  & ~n25365 ;
  assign n25367 = ~n22899 & n25113 ;
  assign n25368 = \pi0788  & ~n25367 ;
  assign n25369 = ~n25366 & n25368 ;
  assign n25370 = ~n25356 & ~n25369 ;
  assign n25371 = ~\pi0788  & ~n25321 ;
  assign n25372 = ~n25313 & n25371 ;
  assign n25373 = \pi0628  & ~n25372 ;
  assign n25374 = n22907 & ~n25350 ;
  assign n25375 = ~n25373 & ~n25374 ;
  assign n25376 = ~n25185 & ~n25375 ;
  assign n25377 = n25370 & n25376 ;
  assign n25378 = ~n25186 & ~n25377 ;
  assign n25379 = n22913 & ~n25378 ;
  assign n25380 = ~\pi0628  & ~n25372 ;
  assign n25381 = n22916 & ~n25350 ;
  assign n25382 = ~n25380 & ~n25381 ;
  assign n25383 = n25370 & ~n25382 ;
  assign n25384 = \pi0788  & ~n25125 ;
  assign n25385 = \pi0628  & n25100 ;
  assign n25386 = ~n25384 & n25385 ;
  assign n25387 = ~\pi1156  & ~n25386 ;
  assign n25388 = ~n25383 & n25387 ;
  assign n25389 = ~\pi0143  & ~\pi0628  ;
  assign n25390 = n21768 & n25389 ;
  assign n25391 = n21770 & n25389 ;
  assign n25392 = ~n21734 & n25391 ;
  assign n25393 = ~n25390 & ~n25392 ;
  assign n25394 = \pi1156  & n25393 ;
  assign n25395 = \pi0628  & ~n25182 ;
  assign n25396 = ~n25181 & n25395 ;
  assign n25397 = n25394 & ~n25396 ;
  assign n25398 = ~\pi0629  & ~n25397 ;
  assign n25399 = n22913 & n25398 ;
  assign n25400 = ~n25388 & n25399 ;
  assign n25401 = ~n25379 & ~n25400 ;
  assign n25402 = ~\pi0792  & ~n25372 ;
  assign n25403 = n22940 & ~n25350 ;
  assign n25404 = ~n25402 & ~n25403 ;
  assign n25405 = ~\pi0647  & ~n25404 ;
  assign n25406 = n25370 & n25405 ;
  assign n25407 = ~n20846 & n25100 ;
  assign n25408 = n20846 & ~n25015 ;
  assign n25409 = ~\pi1157  & ~n25408 ;
  assign n25410 = ~n25407 & n25409 ;
  assign n25411 = \pi0788  & n25409 ;
  assign n25412 = ~n25125 & n25411 ;
  assign n25413 = ~n25410 & ~n25412 ;
  assign n25414 = ~n22945 & n25413 ;
  assign n25415 = ~n25406 & ~n25414 ;
  assign n25416 = n25401 & n25415 ;
  assign n25417 = \pi0647  & ~n25182 ;
  assign n25418 = ~n25181 & n25417 ;
  assign n25419 = ~n22956 & ~n25418 ;
  assign n25420 = n21768 & n24832 ;
  assign n25421 = n21770 & n24832 ;
  assign n25422 = ~n21734 & n25421 ;
  assign n25423 = ~n25420 & ~n25422 ;
  assign n25424 = \pi1157  & n25423 ;
  assign n25425 = n25419 & n25424 ;
  assign n25426 = ~\pi0628  & ~n25182 ;
  assign n25427 = ~n25181 & n25426 ;
  assign n25428 = n25133 & ~n25427 ;
  assign n25429 = ~n25397 & ~n25428 ;
  assign n25430 = \pi0792  & n25424 ;
  assign n25431 = ~n25429 & n25430 ;
  assign n25432 = ~n25425 & ~n25431 ;
  assign n25433 = ~\pi0630  & n25432 ;
  assign n25434 = ~n25416 & n25433 ;
  assign n25435 = n22956 & ~n25378 ;
  assign n25436 = n22956 & n25398 ;
  assign n25437 = ~n25388 & n25436 ;
  assign n25438 = ~n25435 & ~n25437 ;
  assign n25439 = \pi0647  & ~n25404 ;
  assign n25440 = n25370 & n25439 ;
  assign n25441 = \pi1157  & ~n25408 ;
  assign n25442 = ~n25407 & n25441 ;
  assign n25443 = \pi0788  & n25441 ;
  assign n25444 = ~n25125 & n25443 ;
  assign n25445 = ~n25442 & ~n25444 ;
  assign n25446 = ~n20925 & n25445 ;
  assign n25447 = ~n25440 & ~n25446 ;
  assign n25448 = n25438 & n25447 ;
  assign n25449 = ~\pi0647  & ~n25182 ;
  assign n25450 = ~n25181 & n25449 ;
  assign n25451 = ~n22913 & ~n25450 ;
  assign n25452 = n21768 & n24837 ;
  assign n25453 = n21770 & n24837 ;
  assign n25454 = ~n21734 & n25453 ;
  assign n25455 = ~n25452 & ~n25454 ;
  assign n25456 = ~\pi1157  & n25455 ;
  assign n25457 = n25451 & n25456 ;
  assign n25458 = \pi0792  & n25456 ;
  assign n25459 = ~n25429 & n25458 ;
  assign n25460 = ~n25457 & ~n25459 ;
  assign n25461 = \pi0630  & n25460 ;
  assign n25462 = ~n25448 & n25461 ;
  assign n25463 = ~n25434 & ~n25462 ;
  assign n25464 = \pi0787  & ~n25463 ;
  assign n25465 = ~\pi0787  & ~n25404 ;
  assign n25466 = n25370 & n25465 ;
  assign n25467 = n23011 & ~n25378 ;
  assign n25468 = n23011 & n25398 ;
  assign n25469 = ~n25388 & n25468 ;
  assign n25470 = ~n25467 & ~n25469 ;
  assign n25471 = ~n25466 & n25470 ;
  assign n25472 = ~\pi0790  & n25471 ;
  assign n25473 = ~n25464 & n25472 ;
  assign n25474 = ~n24989 & ~n25008 ;
  assign n25475 = ~n24897 & ~n25474 ;
  assign n25476 = n9948 & ~n25475 ;
  assign n25477 = ~n25473 & n25476 ;
  assign n25478 = n25011 & ~n25477 ;
  assign n25479 = n23021 & ~n25463 ;
  assign n25480 = ~\pi0644  & ~n25471 ;
  assign n25481 = n25432 & n25460 ;
  assign n25482 = \pi0787  & ~n25481 ;
  assign n25483 = ~n25181 & ~n25182 ;
  assign n25484 = ~\pi0792  & ~n25483 ;
  assign n25485 = ~\pi0787  & n25484 ;
  assign n25486 = n23011 & ~n25429 ;
  assign n25487 = ~n25485 & ~n25486 ;
  assign n25488 = \pi0644  & n25487 ;
  assign n25489 = ~n25482 & n25488 ;
  assign n25490 = ~\pi0715  & ~n25489 ;
  assign n25491 = ~n25480 & n25490 ;
  assign n25492 = ~n25479 & n25491 ;
  assign n25493 = ~n21088 & ~n25408 ;
  assign n25494 = ~n25407 & n25493 ;
  assign n25495 = \pi0788  & n25493 ;
  assign n25496 = ~n25125 & n25495 ;
  assign n25497 = ~n25494 & ~n25496 ;
  assign n25498 = n21088 & n25015 ;
  assign n25499 = ~\pi0644  & ~n25498 ;
  assign n25500 = n25497 & n25499 ;
  assign n25501 = ~\pi0143  & \pi0644  ;
  assign n25502 = n21768 & n25501 ;
  assign n25503 = n21770 & n25501 ;
  assign n25504 = ~n21734 & n25503 ;
  assign n25505 = ~n25502 & ~n25504 ;
  assign n25506 = \pi0715  & n25505 ;
  assign n25507 = ~n25500 & n25506 ;
  assign n25508 = ~\pi1160  & ~n25507 ;
  assign n25509 = ~n25492 & n25508 ;
  assign n25510 = ~\pi0143  & ~\pi0644  ;
  assign n25511 = n21768 & n25510 ;
  assign n25512 = n21770 & n25510 ;
  assign n25513 = ~n21734 & n25512 ;
  assign n25514 = ~n25511 & ~n25513 ;
  assign n25515 = ~\pi0715  & n25514 ;
  assign n25516 = \pi1160  & ~n25515 ;
  assign n25517 = \pi0644  & ~n25498 ;
  assign n25518 = \pi1160  & n25517 ;
  assign n25519 = n25497 & n25518 ;
  assign n25520 = ~n25516 & ~n25519 ;
  assign n25521 = \pi0790  & n25520 ;
  assign n25522 = ~\pi0644  & n25487 ;
  assign n25523 = \pi0790  & ~n25522 ;
  assign n25524 = n23065 & ~n25481 ;
  assign n25525 = ~n25523 & ~n25524 ;
  assign n25526 = \pi0715  & ~n25525 ;
  assign n25527 = ~\pi0644  & n25526 ;
  assign n25528 = ~n25466 & n25526 ;
  assign n25529 = n25470 & n25528 ;
  assign n25530 = ~n25527 & ~n25529 ;
  assign n25531 = ~n25521 & n25530 ;
  assign n25532 = n23074 & ~n25521 ;
  assign n25533 = ~n25463 & n25532 ;
  assign n25534 = ~n25531 & ~n25533 ;
  assign n25535 = n25011 & n25534 ;
  assign n25536 = ~n25509 & n25535 ;
  assign n25537 = ~n25478 & ~n25536 ;
  assign n25538 = \pi0057  & \pi0144  ;
  assign n25539 = ~\pi0832  & ~n25538 ;
  assign n25540 = ~\pi0144  & ~n6861 ;
  assign n25541 = n21714 & ~n21731 ;
  assign n25542 = ~n21693 & n25541 ;
  assign n25543 = ~\pi0758  & ~n25542 ;
  assign n25544 = \pi0758  & n21272 ;
  assign n25545 = \pi0299  & ~\pi0758  ;
  assign n25546 = ~n21205 & n25545 ;
  assign n25547 = ~n21238 & n25546 ;
  assign n25548 = ~\pi0299  & ~\pi0758  ;
  assign n25549 = ~n21740 & n25548 ;
  assign n25550 = ~n21738 & n25549 ;
  assign n25551 = ~\pi0039  & ~n25550 ;
  assign n25552 = ~n25547 & n25551 ;
  assign n25553 = ~n25544 & n25552 ;
  assign n25554 = ~n21440 & ~n21441 ;
  assign n25555 = ~\pi0299  & \pi0758  ;
  assign n25556 = ~n25554 & n25555 ;
  assign n25557 = ~n21463 & ~n21464 ;
  assign n25558 = \pi0299  & \pi0758  ;
  assign n25559 = ~n25557 & n25558 ;
  assign n25560 = ~n25556 & ~n25559 ;
  assign n25561 = ~n25553 & n25560 ;
  assign n25562 = ~n25543 & n25561 ;
  assign n25563 = ~\pi0039  & ~n25552 ;
  assign n25564 = ~\pi0039  & \pi0758  ;
  assign n25565 = n21272 & n25564 ;
  assign n25566 = ~n25563 & ~n25565 ;
  assign n25567 = ~\pi0038  & \pi0144  ;
  assign n25568 = n25566 & n25567 ;
  assign n25569 = ~n25562 & n25568 ;
  assign n25570 = ~\pi0144  & \pi0758  ;
  assign n25571 = ~\pi0038  & n25570 ;
  assign n25572 = n25023 & n25571 ;
  assign n25573 = ~\pi0144  & ~n21757 ;
  assign n25574 = \pi0603  & \pi0758  ;
  assign n25575 = ~n20783 & n25574 ;
  assign n25576 = n1689 & ~n25575 ;
  assign n25577 = n8413 & n25576 ;
  assign n25578 = n1354 & n25577 ;
  assign n25579 = n1358 & n25578 ;
  assign n25580 = \pi0038  & ~n25579 ;
  assign n25581 = ~n25573 & n25580 ;
  assign n25582 = \pi0144  & ~n6861 ;
  assign n25583 = ~n25581 & ~n25582 ;
  assign n25584 = ~n25572 & n25583 ;
  assign n25585 = ~n25569 & n25584 ;
  assign n25586 = ~n25540 & ~n25585 ;
  assign n25587 = ~n20999 & ~n21774 ;
  assign n25588 = \pi0785  & n25587 ;
  assign n25589 = ~n20985 & ~n25588 ;
  assign n25590 = ~n25586 & n25589 ;
  assign n25591 = \pi0144  & n21768 ;
  assign n25592 = \pi0144  & n21770 ;
  assign n25593 = ~n21734 & n25592 ;
  assign n25594 = ~n25591 & ~n25593 ;
  assign n25595 = n20985 & ~n25588 ;
  assign n25596 = n25594 & n25595 ;
  assign n25597 = n21776 & n25594 ;
  assign n25598 = ~\pi0781  & ~n25597 ;
  assign n25599 = ~n25596 & n25598 ;
  assign n25600 = ~n25590 & n25599 ;
  assign n25601 = ~\pi0789  & n25600 ;
  assign n25602 = n20809 & ~n25594 ;
  assign n25603 = \pi1154  & ~n25594 ;
  assign n25604 = \pi0618  & \pi1154  ;
  assign n25605 = ~n21776 & n25604 ;
  assign n25606 = ~n25603 & ~n25605 ;
  assign n25607 = ~n25596 & ~n25606 ;
  assign n25608 = ~n25590 & n25607 ;
  assign n25609 = ~n25602 & ~n25608 ;
  assign n25610 = n20810 & ~n25594 ;
  assign n25611 = ~\pi1154  & ~n25594 ;
  assign n25612 = ~\pi0618  & ~\pi1154  ;
  assign n25613 = ~n21776 & n25612 ;
  assign n25614 = ~n25611 & ~n25613 ;
  assign n25615 = ~n25596 & ~n25614 ;
  assign n25616 = ~n25590 & n25615 ;
  assign n25617 = ~n25610 & ~n25616 ;
  assign n25618 = n25609 & n25617 ;
  assign n25619 = n21806 & ~n25618 ;
  assign n25620 = ~n25601 & ~n25619 ;
  assign n25621 = ~\pi0788  & ~n25620 ;
  assign n25622 = ~\pi0619  & ~n25600 ;
  assign n25623 = \pi0619  & n25594 ;
  assign n25624 = ~\pi1159  & ~n25623 ;
  assign n25625 = ~n25622 & n25624 ;
  assign n25626 = \pi0781  & n25624 ;
  assign n25627 = ~n25618 & n25626 ;
  assign n25628 = ~n25625 & ~n25627 ;
  assign n25629 = \pi0619  & ~n25600 ;
  assign n25630 = ~\pi0619  & n25594 ;
  assign n25631 = \pi1159  & ~n25630 ;
  assign n25632 = ~n25629 & n25631 ;
  assign n25633 = \pi0781  & n25631 ;
  assign n25634 = ~n25618 & n25633 ;
  assign n25635 = ~n25632 & ~n25634 ;
  assign n25636 = n25628 & n25635 ;
  assign n25637 = n21832 & ~n25636 ;
  assign n25638 = ~n25621 & ~n25637 ;
  assign n25639 = ~\pi0628  & n25638 ;
  assign n25640 = \pi1156  & ~n25639 ;
  assign n25641 = ~\pi0626  & n25620 ;
  assign n25642 = \pi0626  & n25594 ;
  assign n25643 = ~\pi1158  & ~n25642 ;
  assign n25644 = ~n25641 & n25643 ;
  assign n25645 = \pi0789  & n25643 ;
  assign n25646 = ~n25636 & n25645 ;
  assign n25647 = ~n25644 & ~n25646 ;
  assign n25648 = \pi0626  & n25620 ;
  assign n25649 = ~\pi0626  & n25594 ;
  assign n25650 = \pi1158  & ~n25649 ;
  assign n25651 = ~n25648 & n25650 ;
  assign n25652 = \pi0789  & n25650 ;
  assign n25653 = ~n25636 & n25652 ;
  assign n25654 = ~n25651 & ~n25653 ;
  assign n25655 = n25647 & n25654 ;
  assign n25656 = n21860 & ~n25655 ;
  assign n25657 = ~n25640 & ~n25656 ;
  assign n25658 = \pi0629  & \pi1156  ;
  assign n25659 = \pi0628  & \pi0629  ;
  assign n25660 = n25594 & n25659 ;
  assign n25661 = ~n25658 & ~n25660 ;
  assign n25662 = ~n22166 & n25661 ;
  assign n25663 = ~\pi0074  & \pi0736  ;
  assign n25664 = ~\pi0100  & n25663 ;
  assign n25665 = n1287 & n25664 ;
  assign n25666 = n8413 & n21931 ;
  assign n25667 = n1354 & n25666 ;
  assign n25668 = n1358 & n25667 ;
  assign n25669 = \pi0038  & ~n25668 ;
  assign n25670 = ~n25573 & n25669 ;
  assign n25671 = \pi0144  & n22017 ;
  assign n25672 = \pi0039  & \pi0144  ;
  assign n25673 = ~n21993 & n25672 ;
  assign n25674 = ~n25671 & ~n25673 ;
  assign n25675 = ~\pi0144  & ~n22107 ;
  assign n25676 = n22089 & n25675 ;
  assign n25677 = ~\pi0038  & ~n25676 ;
  assign n25678 = n25674 & n25677 ;
  assign n25679 = ~n25670 & ~n25678 ;
  assign n25680 = n25665 & ~n25679 ;
  assign n25681 = \pi0144  & ~n25665 ;
  assign n25682 = n21768 & n25681 ;
  assign n25683 = n21770 & n25681 ;
  assign n25684 = ~n21734 & n25683 ;
  assign n25685 = ~n25682 & ~n25684 ;
  assign n25686 = \pi0625  & n25685 ;
  assign n25687 = ~n25680 & n25686 ;
  assign n25688 = \pi0144  & \pi1153  ;
  assign n25689 = n21768 & n25688 ;
  assign n25690 = n21770 & n25688 ;
  assign n25691 = ~n21734 & n25690 ;
  assign n25692 = ~n25689 & ~n25691 ;
  assign n25693 = ~n24550 & n25692 ;
  assign n25694 = ~n25687 & ~n25693 ;
  assign n25695 = ~\pi0625  & n25685 ;
  assign n25696 = ~n25680 & n25695 ;
  assign n25697 = \pi0144  & ~\pi1153  ;
  assign n25698 = n21768 & n25697 ;
  assign n25699 = n21770 & n25697 ;
  assign n25700 = ~n21734 & n25699 ;
  assign n25701 = ~n25698 & ~n25700 ;
  assign n25702 = ~n24561 & n25701 ;
  assign n25703 = ~n25696 & ~n25702 ;
  assign n25704 = ~n25694 & ~n25703 ;
  assign n25705 = \pi0778  & ~n25704 ;
  assign n25706 = ~\pi0778  & ~n25685 ;
  assign n25707 = ~\pi0778  & n25665 ;
  assign n25708 = ~n25679 & n25707 ;
  assign n25709 = ~n25706 & ~n25708 ;
  assign n25710 = ~n22147 & n25709 ;
  assign n25711 = ~n25705 & n25710 ;
  assign n25712 = n22147 & n25594 ;
  assign n25713 = ~n22155 & ~n25712 ;
  assign n25714 = ~n25711 & n25713 ;
  assign n25715 = n22155 & ~n25594 ;
  assign n25716 = n22162 & ~n25715 ;
  assign n25717 = ~n25714 & n25716 ;
  assign n25718 = ~n22162 & n25594 ;
  assign n25719 = n25661 & ~n25718 ;
  assign n25720 = ~n25717 & n25719 ;
  assign n25721 = ~n25662 & ~n25720 ;
  assign n25722 = n25657 & n25721 ;
  assign n25723 = ~\pi0736  & ~n25581 ;
  assign n25724 = ~n25572 & n25723 ;
  assign n25725 = ~n25569 & n25724 ;
  assign n25726 = ~\pi0144  & ~\pi0778  ;
  assign n25727 = ~n23622 & ~n25726 ;
  assign n25728 = n25725 & ~n25727 ;
  assign n25729 = ~\pi0144  & ~n22468 ;
  assign n25730 = ~\pi0144  & ~n22509 ;
  assign n25731 = n22487 & n25730 ;
  assign n25732 = ~n25729 & ~n25731 ;
  assign n25733 = ~\pi0144  & \pi0299  ;
  assign n25734 = ~n22530 & n25733 ;
  assign n25735 = \pi0144  & ~\pi0299  ;
  assign n25736 = ~n22601 & n25735 ;
  assign n25737 = \pi0144  & \pi0299  ;
  assign n25738 = ~n22630 & n25737 ;
  assign n25739 = \pi0758  & ~n25738 ;
  assign n25740 = ~n25736 & n25739 ;
  assign n25741 = ~n25734 & n25740 ;
  assign n25742 = n25732 & n25741 ;
  assign n25743 = \pi0039  & ~n25742 ;
  assign n25744 = ~n22407 & n25735 ;
  assign n25745 = ~n22291 & n25737 ;
  assign n25746 = ~n25744 & ~n25745 ;
  assign n25747 = ~n22431 & n25733 ;
  assign n25748 = ~\pi0144  & n22379 ;
  assign n25749 = ~\pi0758  & ~n25748 ;
  assign n25750 = ~n25747 & n25749 ;
  assign n25751 = n25746 & n25750 ;
  assign n25752 = n25743 & ~n25751 ;
  assign n25753 = ~\pi0038  & ~n25752 ;
  assign n25754 = n22693 & n25570 ;
  assign n25755 = \pi0144  & \pi0758  ;
  assign n25756 = n22683 & n25755 ;
  assign n25757 = ~n25754 & ~n25756 ;
  assign n25758 = \pi0144  & n22643 ;
  assign n25759 = ~n22652 & n25758 ;
  assign n25760 = n11250 & n22676 ;
  assign n25761 = ~n22657 & n25733 ;
  assign n25762 = ~n22660 & n25761 ;
  assign n25763 = n22664 & n25762 ;
  assign n25764 = ~\pi0758  & ~n25763 ;
  assign n25765 = ~n25760 & n25764 ;
  assign n25766 = ~n25759 & n25765 ;
  assign n25767 = n25757 & ~n25766 ;
  assign n25768 = ~\pi0039  & ~n25767 ;
  assign n25769 = n6861 & ~n25768 ;
  assign n25770 = n25753 & n25769 ;
  assign n25771 = \pi0736  & ~n25217 ;
  assign n25772 = ~n25581 & n25771 ;
  assign n25773 = n6861 & ~n25772 ;
  assign n25774 = ~n25727 & ~n25773 ;
  assign n25775 = ~n25770 & n25774 ;
  assign n25776 = ~n25728 & ~n25775 ;
  assign n25777 = ~\pi0785  & ~n25776 ;
  assign n25778 = \pi0618  & n25777 ;
  assign n25779 = ~\pi0144  & ~\pi0625  ;
  assign n25780 = ~n22734 & ~n25779 ;
  assign n25781 = n25725 & ~n25780 ;
  assign n25782 = ~n25773 & ~n25780 ;
  assign n25783 = ~n25770 & n25782 ;
  assign n25784 = ~n25781 & ~n25783 ;
  assign n25785 = \pi0625  & ~n25586 ;
  assign n25786 = ~\pi1153  & ~n25785 ;
  assign n25787 = n25784 & n25786 ;
  assign n25788 = ~\pi0608  & ~n25694 ;
  assign n25789 = ~n25787 & n25788 ;
  assign n25790 = ~\pi0144  & \pi0625  ;
  assign n25791 = ~n22727 & ~n25790 ;
  assign n25792 = n25725 & ~n25791 ;
  assign n25793 = ~n25773 & ~n25791 ;
  assign n25794 = ~n25770 & n25793 ;
  assign n25795 = ~n25792 & ~n25794 ;
  assign n25796 = \pi1153  & ~n25540 ;
  assign n25797 = ~n25585 & n25796 ;
  assign n25798 = ~n24550 & ~n25797 ;
  assign n25799 = n25795 & ~n25798 ;
  assign n25800 = \pi0608  & ~n25703 ;
  assign n25801 = ~n25799 & n25800 ;
  assign n25802 = ~n25789 & ~n25801 ;
  assign n25803 = \pi0618  & n23673 ;
  assign n25804 = ~n25802 & n25803 ;
  assign n25805 = ~n25778 & ~n25804 ;
  assign n25806 = \pi1154  & ~n25712 ;
  assign n25807 = ~n25711 & n25806 ;
  assign n25808 = ~n25604 & ~n25807 ;
  assign n25809 = n25805 & ~n25808 ;
  assign n25810 = \pi0627  & ~n25610 ;
  assign n25811 = ~n25616 & n25810 ;
  assign n25812 = ~n25809 & n25811 ;
  assign n25813 = n23613 & ~n25802 ;
  assign n25814 = \pi0609  & n25709 ;
  assign n25815 = ~n25705 & n25814 ;
  assign n25816 = ~\pi0609  & ~n25776 ;
  assign n25817 = ~\pi1155  & ~n25816 ;
  assign n25818 = ~n25815 & n25817 ;
  assign n25819 = ~n25813 & n25818 ;
  assign n25820 = \pi0609  & n20985 ;
  assign n25821 = n25594 & n25820 ;
  assign n25822 = ~\pi0609  & n25594 ;
  assign n25823 = \pi1155  & ~n25822 ;
  assign n25824 = ~n22788 & n25823 ;
  assign n25825 = ~n25540 & n25823 ;
  assign n25826 = ~n25585 & n25825 ;
  assign n25827 = ~n25824 & ~n25826 ;
  assign n25828 = ~n25821 & ~n25827 ;
  assign n25829 = ~\pi0660  & ~n25828 ;
  assign n25830 = ~n25819 & n25829 ;
  assign n25831 = n23638 & ~n25802 ;
  assign n25832 = \pi0609  & ~n25776 ;
  assign n25833 = ~\pi0609  & n25709 ;
  assign n25834 = \pi1155  & ~n25833 ;
  assign n25835 = n22722 & ~n25704 ;
  assign n25836 = ~n25834 & ~n25835 ;
  assign n25837 = ~n25832 & ~n25836 ;
  assign n25838 = ~n25831 & n25837 ;
  assign n25839 = ~\pi0609  & n20985 ;
  assign n25840 = n25594 & n25839 ;
  assign n25841 = \pi0609  & n25594 ;
  assign n25842 = ~\pi1155  & ~n25841 ;
  assign n25843 = ~n22767 & n25842 ;
  assign n25844 = ~n25540 & n25842 ;
  assign n25845 = ~n25585 & n25844 ;
  assign n25846 = ~n25843 & ~n25845 ;
  assign n25847 = ~n25840 & ~n25846 ;
  assign n25848 = \pi0660  & ~n25847 ;
  assign n25849 = ~n25838 & n25848 ;
  assign n25850 = ~n25830 & ~n25849 ;
  assign n25851 = n22816 & n25811 ;
  assign n25852 = ~n25850 & n25851 ;
  assign n25853 = ~n25812 & ~n25852 ;
  assign n25854 = n21806 & ~n25853 ;
  assign n25855 = n22776 & ~n25850 ;
  assign n25856 = ~\pi0618  & n25777 ;
  assign n25857 = ~\pi0618  & n23673 ;
  assign n25858 = ~n25802 & n25857 ;
  assign n25859 = ~n25856 & ~n25858 ;
  assign n25860 = ~\pi1154  & ~n25712 ;
  assign n25861 = ~n25711 & n25860 ;
  assign n25862 = ~n25612 & ~n25861 ;
  assign n25863 = n25859 & ~n25862 ;
  assign n25864 = ~n25855 & n25863 ;
  assign n25865 = ~\pi0627  & ~n25602 ;
  assign n25866 = ~n25608 & n25865 ;
  assign n25867 = n21806 & n25866 ;
  assign n25868 = ~n25864 & n25867 ;
  assign n25869 = ~n25854 & ~n25868 ;
  assign n25870 = ~\pi0781  & n25777 ;
  assign n25871 = ~\pi0781  & n23673 ;
  assign n25872 = ~n25802 & n25871 ;
  assign n25873 = ~n25870 & ~n25872 ;
  assign n25874 = ~\pi0789  & ~n25873 ;
  assign n25875 = ~\pi0789  & n22840 ;
  assign n25876 = ~n25850 & n25875 ;
  assign n25877 = ~n25874 & ~n25876 ;
  assign n25878 = \pi0626  & n25877 ;
  assign n25879 = n25869 & n25878 ;
  assign n25880 = ~n25711 & ~n25712 ;
  assign n25881 = n22849 & ~n25880 ;
  assign n25882 = ~n22849 & n25594 ;
  assign n25883 = ~\pi0626  & ~n25882 ;
  assign n25884 = ~n25881 & n25883 ;
  assign n25885 = \pi0641  & ~n25884 ;
  assign n25886 = ~n25879 & n25885 ;
  assign n25887 = n22859 & ~n25853 ;
  assign n25888 = n22859 & n25866 ;
  assign n25889 = ~n25864 & n25888 ;
  assign n25890 = ~n25887 & ~n25889 ;
  assign n25891 = \pi0619  & ~n25873 ;
  assign n25892 = \pi0619  & n22840 ;
  assign n25893 = ~n25850 & n25892 ;
  assign n25894 = ~n25891 & ~n25893 ;
  assign n25895 = ~\pi0619  & ~n25715 ;
  assign n25896 = ~n25714 & n25895 ;
  assign n25897 = \pi1159  & ~n25896 ;
  assign n25898 = n25894 & n25897 ;
  assign n25899 = n25890 & n25898 ;
  assign n25900 = \pi0648  & n25628 ;
  assign n25901 = ~n25899 & n25900 ;
  assign n25902 = n22869 & ~n25853 ;
  assign n25903 = n22869 & n25866 ;
  assign n25904 = ~n25864 & n25903 ;
  assign n25905 = ~n25902 & ~n25904 ;
  assign n25906 = ~\pi0619  & ~n25873 ;
  assign n25907 = ~\pi0619  & n22840 ;
  assign n25908 = ~n25850 & n25907 ;
  assign n25909 = ~n25906 & ~n25908 ;
  assign n25910 = \pi0619  & ~n25715 ;
  assign n25911 = ~n25714 & n25910 ;
  assign n25912 = ~\pi1159  & ~n25911 ;
  assign n25913 = n25909 & n25912 ;
  assign n25914 = n25905 & n25913 ;
  assign n25915 = ~\pi0648  & n25635 ;
  assign n25916 = ~n25914 & n25915 ;
  assign n25917 = ~n25901 & ~n25916 ;
  assign n25918 = \pi0789  & n25885 ;
  assign n25919 = ~n25917 & n25918 ;
  assign n25920 = ~n25886 & ~n25919 ;
  assign n25921 = ~n22884 & n25654 ;
  assign n25922 = n25920 & ~n25921 ;
  assign n25923 = \pi0788  & n25922 ;
  assign n25924 = ~\pi0626  & n25877 ;
  assign n25925 = n25869 & n25924 ;
  assign n25926 = \pi0626  & ~n25882 ;
  assign n25927 = ~n25881 & n25926 ;
  assign n25928 = ~n25925 & ~n25927 ;
  assign n25929 = \pi0789  & ~n25927 ;
  assign n25930 = ~n25917 & n25929 ;
  assign n25931 = ~n25928 & ~n25930 ;
  assign n25932 = ~\pi0641  & ~n25931 ;
  assign n25933 = ~n22899 & n25647 ;
  assign n25934 = \pi0788  & ~n25933 ;
  assign n25935 = ~n25932 & n25934 ;
  assign n25936 = ~n25923 & ~n25935 ;
  assign n25937 = ~\pi0788  & n25877 ;
  assign n25938 = n25869 & n25937 ;
  assign n25939 = \pi0628  & ~n25938 ;
  assign n25940 = n22907 & ~n25917 ;
  assign n25941 = ~n25939 & ~n25940 ;
  assign n25942 = n25721 & ~n25941 ;
  assign n25943 = n25936 & n25942 ;
  assign n25944 = ~n25722 & ~n25943 ;
  assign n25945 = n23011 & ~n25944 ;
  assign n25946 = ~\pi0628  & ~n25938 ;
  assign n25947 = n22916 & ~n25917 ;
  assign n25948 = ~n25946 & ~n25947 ;
  assign n25949 = n25936 & ~n25948 ;
  assign n25950 = \pi0788  & ~n25655 ;
  assign n25951 = \pi0628  & n25638 ;
  assign n25952 = ~n25950 & n25951 ;
  assign n25953 = ~\pi1156  & ~n25952 ;
  assign n25954 = ~n25949 & n25953 ;
  assign n25955 = ~\pi0629  & ~\pi1156  ;
  assign n25956 = ~\pi0628  & ~\pi0629  ;
  assign n25957 = n25594 & n25956 ;
  assign n25958 = ~n25955 & ~n25957 ;
  assign n25959 = ~n22932 & n25958 ;
  assign n25960 = ~n25718 & n25958 ;
  assign n25961 = ~n25717 & n25960 ;
  assign n25962 = ~n25959 & ~n25961 ;
  assign n25963 = n23011 & n25962 ;
  assign n25964 = ~n25954 & n25963 ;
  assign n25965 = ~n25945 & ~n25964 ;
  assign n25966 = ~\pi0792  & ~n25938 ;
  assign n25967 = n22940 & ~n25917 ;
  assign n25968 = ~n25966 & ~n25967 ;
  assign n25969 = ~\pi0787  & ~n25968 ;
  assign n25970 = n25936 & n25969 ;
  assign n25971 = ~\pi0790  & ~n25970 ;
  assign n25972 = n25965 & n25971 ;
  assign n25973 = n25539 & ~n25972 ;
  assign n25974 = n22913 & ~n25944 ;
  assign n25975 = n22913 & n25962 ;
  assign n25976 = ~n25954 & n25975 ;
  assign n25977 = ~n25974 & ~n25976 ;
  assign n25978 = ~\pi0647  & ~n25968 ;
  assign n25979 = n25936 & n25978 ;
  assign n25980 = ~n20846 & ~n25638 ;
  assign n25981 = n24737 & ~n25655 ;
  assign n25982 = ~n25980 & ~n25981 ;
  assign n25983 = n20846 & ~n25594 ;
  assign n25984 = \pi0647  & ~n25983 ;
  assign n25985 = n25982 & n25984 ;
  assign n25986 = ~\pi1157  & ~n25985 ;
  assign n25987 = ~n25979 & n25986 ;
  assign n25988 = n25977 & n25987 ;
  assign n25989 = ~\pi0792  & ~n25718 ;
  assign n25990 = ~n25717 & n25989 ;
  assign n25991 = \pi0647  & ~n25990 ;
  assign n25992 = \pi0144  & \pi1157  ;
  assign n25993 = n21768 & n25992 ;
  assign n25994 = n21770 & n25992 ;
  assign n25995 = ~n21734 & n25994 ;
  assign n25996 = ~n25993 & ~n25995 ;
  assign n25997 = ~n20925 & n25996 ;
  assign n25998 = ~n25991 & ~n25997 ;
  assign n25999 = ~\pi0628  & n25594 ;
  assign n26000 = \pi1156  & ~n25999 ;
  assign n26001 = ~\pi0628  & n26000 ;
  assign n26002 = ~n25718 & n26000 ;
  assign n26003 = ~n25717 & n26002 ;
  assign n26004 = ~n26001 & ~n26003 ;
  assign n26005 = \pi0628  & n25594 ;
  assign n26006 = ~\pi1156  & ~n26005 ;
  assign n26007 = \pi0628  & n26006 ;
  assign n26008 = ~n25718 & n26006 ;
  assign n26009 = ~n25717 & n26008 ;
  assign n26010 = ~n26007 & ~n26009 ;
  assign n26011 = n26004 & n26010 ;
  assign n26012 = \pi0792  & ~n25997 ;
  assign n26013 = ~n26011 & n26012 ;
  assign n26014 = ~n25998 & ~n26013 ;
  assign n26015 = ~\pi0630  & n26014 ;
  assign n26016 = ~n25988 & n26015 ;
  assign n26017 = n22956 & ~n25944 ;
  assign n26018 = n22956 & n25962 ;
  assign n26019 = ~n25954 & n26018 ;
  assign n26020 = ~n26017 & ~n26019 ;
  assign n26021 = \pi0647  & ~n25968 ;
  assign n26022 = n25936 & n26021 ;
  assign n26023 = ~\pi0647  & ~n25983 ;
  assign n26024 = n25982 & n26023 ;
  assign n26025 = \pi1157  & ~n26024 ;
  assign n26026 = ~n26022 & n26025 ;
  assign n26027 = n26020 & n26026 ;
  assign n26028 = ~\pi0647  & ~n25990 ;
  assign n26029 = \pi0144  & ~\pi1157  ;
  assign n26030 = n21768 & n26029 ;
  assign n26031 = n21770 & n26029 ;
  assign n26032 = ~n21734 & n26031 ;
  assign n26033 = ~n26030 & ~n26032 ;
  assign n26034 = ~n22945 & n26033 ;
  assign n26035 = ~n26028 & ~n26034 ;
  assign n26036 = \pi0792  & ~n26034 ;
  assign n26037 = ~n26011 & n26036 ;
  assign n26038 = ~n26035 & ~n26037 ;
  assign n26039 = \pi0630  & n26038 ;
  assign n26040 = ~n26027 & n26039 ;
  assign n26041 = ~n26016 & ~n26040 ;
  assign n26042 = \pi0787  & n25539 ;
  assign n26043 = ~n26041 & n26042 ;
  assign n26044 = ~n25973 & ~n26043 ;
  assign n26045 = n6848 & ~n26044 ;
  assign n26046 = ~\pi0144  & ~\pi0832  ;
  assign n26047 = ~n6848 & n26046 ;
  assign n26048 = \pi0057  & ~\pi0144  ;
  assign n26049 = ~\pi0832  & n26048 ;
  assign n26050 = ~n26047 & ~n26049 ;
  assign n26051 = \pi0144  & ~n1689 ;
  assign n26052 = \pi0736  & n1689 ;
  assign n26053 = n20855 & n26052 ;
  assign n26054 = ~n26051 & ~n26053 ;
  assign n26055 = ~\pi0778  & ~n26054 ;
  assign n26056 = n23885 & n26055 ;
  assign n26057 = \pi0625  & \pi0736  ;
  assign n26058 = n1689 & n26057 ;
  assign n26059 = n20855 & n26058 ;
  assign n26060 = ~n26051 & ~n26059 ;
  assign n26061 = \pi1153  & ~n26060 ;
  assign n26062 = ~\pi1153  & ~n26059 ;
  assign n26063 = ~n26054 & n26062 ;
  assign n26064 = ~n26061 & ~n26063 ;
  assign n26065 = \pi0778  & n23885 ;
  assign n26066 = ~n26064 & n26065 ;
  assign n26067 = ~n26056 & ~n26066 ;
  assign n26068 = n23518 & ~n23942 ;
  assign n26069 = ~n23907 & n26068 ;
  assign n26070 = ~n26067 & n26069 ;
  assign n26071 = \pi0758  & n1689 ;
  assign n26072 = n20784 & n26071 ;
  assign n26073 = ~n20846 & n26072 ;
  assign n26074 = ~n23880 & n26073 ;
  assign n26075 = n23832 & n26074 ;
  assign n26076 = ~\pi0644  & ~n23316 ;
  assign n26077 = ~\pi1160  & n26076 ;
  assign n26078 = ~n21088 & n26077 ;
  assign n26079 = n26075 & n26078 ;
  assign n26080 = \pi0644  & ~n23315 ;
  assign n26081 = \pi1160  & n26080 ;
  assign n26082 = ~n21088 & n26081 ;
  assign n26083 = n26075 & n26082 ;
  assign n26084 = n26051 & n26080 ;
  assign n26085 = n26051 & n26076 ;
  assign n26086 = ~n26084 & ~n26085 ;
  assign n26087 = ~n26083 & n26086 ;
  assign n26088 = ~n26079 & n26087 ;
  assign n26089 = ~n26070 & n26088 ;
  assign n26090 = \pi0790  & ~n26089 ;
  assign n26091 = \pi0832  & ~n26090 ;
  assign n26092 = ~\pi0630  & ~n23880 ;
  assign n26093 = n26073 & n26092 ;
  assign n26094 = n23832 & n26093 ;
  assign n26095 = n21064 & ~n26094 ;
  assign n26096 = n20897 & n23907 ;
  assign n26097 = n20897 & ~n26056 ;
  assign n26098 = ~n26066 & n26097 ;
  assign n26099 = ~n26096 & ~n26098 ;
  assign n26100 = ~n26095 & n26099 ;
  assign n26101 = \pi0787  & ~n26051 ;
  assign n26102 = ~n26100 & n26101 ;
  assign n26103 = ~\pi0630  & n23907 ;
  assign n26104 = ~\pi0630  & ~n26056 ;
  assign n26105 = ~n26066 & n26104 ;
  assign n26106 = ~n26103 & ~n26105 ;
  assign n26107 = \pi0647  & n26106 ;
  assign n26108 = \pi0630  & ~n23880 ;
  assign n26109 = n26073 & n26108 ;
  assign n26110 = n23832 & n26109 ;
  assign n26111 = \pi1157  & ~n26110 ;
  assign n26112 = n26101 & n26111 ;
  assign n26113 = ~n26107 & n26112 ;
  assign n26114 = ~n26102 & ~n26113 ;
  assign n26115 = ~n24761 & n26114 ;
  assign n26116 = n26091 & ~n26115 ;
  assign n26117 = n22787 & n23638 ;
  assign n26118 = n22766 & n23613 ;
  assign n26119 = ~n26117 & ~n26118 ;
  assign n26120 = ~n26064 & ~n26119 ;
  assign n26121 = ~\pi0609  & \pi1155  ;
  assign n26122 = \pi0660  & n26121 ;
  assign n26123 = ~\pi1155  & n23804 ;
  assign n26124 = ~n26122 & ~n26123 ;
  assign n26125 = ~\pi0778  & ~n26124 ;
  assign n26126 = ~n26054 & n26125 ;
  assign n26127 = ~n20866 & n26051 ;
  assign n26128 = ~n20985 & ~n23806 ;
  assign n26129 = ~n20866 & n26072 ;
  assign n26130 = n26128 & n26129 ;
  assign n26131 = ~n26127 & ~n26130 ;
  assign n26132 = ~n26126 & n26131 ;
  assign n26133 = ~n26120 & n26132 ;
  assign n26134 = \pi0785  & ~n26133 ;
  assign n26135 = n21022 & n23808 ;
  assign n26136 = n20784 & ~n26051 ;
  assign n26137 = ~n20985 & n26136 ;
  assign n26138 = ~n26054 & ~n26137 ;
  assign n26139 = n21022 & ~n26072 ;
  assign n26140 = ~n26138 & n26139 ;
  assign n26141 = ~n26135 & ~n26140 ;
  assign n26142 = ~n21034 & ~n26141 ;
  assign n26143 = \pi0608  & n26059 ;
  assign n26144 = \pi0608  & ~n26051 ;
  assign n26145 = ~n26053 & n26144 ;
  assign n26146 = ~n26143 & ~n26145 ;
  assign n26147 = \pi0625  & ~n20784 ;
  assign n26148 = n26053 & n26147 ;
  assign n26149 = ~\pi1153  & ~n26148 ;
  assign n26150 = n26146 & n26149 ;
  assign n26151 = ~\pi0625  & ~n26072 ;
  assign n26152 = n20788 & ~n26151 ;
  assign n26153 = \pi0778  & ~n26152 ;
  assign n26154 = ~n26150 & n26153 ;
  assign n26155 = n21022 & ~n26061 ;
  assign n26156 = ~n21034 & n26155 ;
  assign n26157 = n26154 & n26156 ;
  assign n26158 = ~n26142 & ~n26157 ;
  assign n26159 = ~n26134 & ~n26158 ;
  assign n26160 = n23666 & n26072 ;
  assign n26161 = n21777 & n26160 ;
  assign n26162 = \pi0781  & ~n26051 ;
  assign n26163 = n20871 & n26162 ;
  assign n26164 = ~n26161 & n26163 ;
  assign n26165 = n22148 & ~n26064 ;
  assign n26166 = n22151 & ~n26054 ;
  assign n26167 = n23667 & n26162 ;
  assign n26168 = ~n26166 & n26167 ;
  assign n26169 = ~n26165 & n26168 ;
  assign n26170 = ~n26164 & ~n26169 ;
  assign n26171 = ~n21034 & ~n26170 ;
  assign n26172 = n21050 & n23380 ;
  assign n26173 = n26055 & n26172 ;
  assign n26174 = \pi0778  & n26172 ;
  assign n26175 = ~n26064 & n26174 ;
  assign n26176 = n21032 & ~n23830 ;
  assign n26177 = n21777 & n26176 ;
  assign n26178 = n26072 & n26177 ;
  assign n26179 = n21034 & ~n26051 ;
  assign n26180 = ~n26178 & n26179 ;
  assign n26181 = ~n26175 & n26180 ;
  assign n26182 = ~n26173 & n26181 ;
  assign n26183 = ~n21038 & ~n26182 ;
  assign n26184 = ~n26171 & n26183 ;
  assign n26185 = ~n26159 & n26184 ;
  assign n26186 = ~n22160 & n23380 ;
  assign n26187 = \pi0778  & n26186 ;
  assign n26188 = ~n26064 & n26187 ;
  assign n26189 = n26055 & n26186 ;
  assign n26190 = ~n26051 & ~n26189 ;
  assign n26191 = ~n26188 & n26190 ;
  assign n26192 = n20777 & ~n26191 ;
  assign n26193 = ~\pi0641  & ~n26051 ;
  assign n26194 = ~n22899 & ~n26193 ;
  assign n26195 = \pi0603  & \pi0626  ;
  assign n26196 = ~n20783 & n26195 ;
  assign n26197 = n26071 & n26196 ;
  assign n26198 = ~n22899 & n26197 ;
  assign n26199 = n23832 & n26198 ;
  assign n26200 = ~n26194 & ~n26199 ;
  assign n26201 = ~n26192 & n26200 ;
  assign n26202 = \pi0641  & ~n26051 ;
  assign n26203 = ~n22884 & ~n26202 ;
  assign n26204 = \pi0603  & ~\pi0626  ;
  assign n26205 = ~n20783 & n26204 ;
  assign n26206 = n26071 & n26205 ;
  assign n26207 = ~n22884 & n26206 ;
  assign n26208 = n23832 & n26207 ;
  assign n26209 = ~n26203 & ~n26208 ;
  assign n26210 = \pi0788  & ~n26209 ;
  assign n26211 = \pi0788  & n20776 ;
  assign n26212 = ~n26191 & n26211 ;
  assign n26213 = ~n26210 & ~n26212 ;
  assign n26214 = ~n26201 & ~n26213 ;
  assign n26215 = ~n23856 & ~n26214 ;
  assign n26216 = ~n26185 & n26215 ;
  assign n26217 = ~\pi0628  & ~n26067 ;
  assign n26218 = \pi0792  & ~\pi1156  ;
  assign n26219 = ~n26051 & n26218 ;
  assign n26220 = \pi0629  & n26219 ;
  assign n26221 = ~n23880 & n26072 ;
  assign n26222 = n23832 & n26221 ;
  assign n26223 = \pi0628  & n26219 ;
  assign n26224 = ~n26222 & n26223 ;
  assign n26225 = ~n26220 & ~n26224 ;
  assign n26226 = ~n26217 & ~n26225 ;
  assign n26227 = \pi0628  & ~n26067 ;
  assign n26228 = \pi0792  & ~n26051 ;
  assign n26229 = n20886 & ~n26222 ;
  assign n26230 = ~n20843 & ~n26229 ;
  assign n26231 = n26228 & ~n26230 ;
  assign n26232 = ~n26227 & n26231 ;
  assign n26233 = ~n26226 & ~n26232 ;
  assign n26234 = ~n26216 & n26233 ;
  assign n26235 = ~n21067 & n26091 ;
  assign n26236 = ~n26234 & n26235 ;
  assign n26237 = ~n26116 & ~n26236 ;
  assign n26238 = n26050 & n26237 ;
  assign n26239 = ~n26045 & n26238 ;
  assign n26240 = n23021 & ~n26041 ;
  assign n26241 = n25965 & ~n25970 ;
  assign n26242 = ~\pi0644  & ~n26241 ;
  assign n26243 = n26014 & n26038 ;
  assign n26244 = \pi0787  & ~n26243 ;
  assign n26245 = ~\pi0787  & n25990 ;
  assign n26246 = n23011 & ~n26011 ;
  assign n26247 = ~n26245 & ~n26246 ;
  assign n26248 = \pi0644  & n26247 ;
  assign n26249 = ~n26244 & n26248 ;
  assign n26250 = ~\pi0715  & ~n26249 ;
  assign n26251 = ~n26242 & n26250 ;
  assign n26252 = ~n26240 & n26251 ;
  assign n26253 = \pi0144  & \pi0715  ;
  assign n26254 = n21768 & n26253 ;
  assign n26255 = n21770 & n26253 ;
  assign n26256 = ~n21734 & n26255 ;
  assign n26257 = ~n26254 & ~n26256 ;
  assign n26258 = ~n23313 & n26257 ;
  assign n26259 = n21088 & n25594 ;
  assign n26260 = ~n26258 & ~n26259 ;
  assign n26261 = \pi0644  & ~n26257 ;
  assign n26262 = ~\pi1160  & ~n26261 ;
  assign n26263 = ~n26260 & n26262 ;
  assign n26264 = ~n21088 & ~n25983 ;
  assign n26265 = n26262 & n26264 ;
  assign n26266 = n25982 & n26265 ;
  assign n26267 = ~n26263 & ~n26266 ;
  assign n26268 = ~n26252 & ~n26267 ;
  assign n26269 = \pi0144  & ~\pi0715  ;
  assign n26270 = n21768 & n26269 ;
  assign n26271 = n21770 & n26269 ;
  assign n26272 = ~n21734 & n26271 ;
  assign n26273 = ~n26270 & ~n26272 ;
  assign n26274 = ~n23312 & n26273 ;
  assign n26275 = ~n26259 & ~n26274 ;
  assign n26276 = ~\pi0644  & ~n26273 ;
  assign n26277 = \pi1160  & ~n26276 ;
  assign n26278 = ~n26275 & n26277 ;
  assign n26279 = n26264 & n26277 ;
  assign n26280 = n25982 & n26279 ;
  assign n26281 = ~n26278 & ~n26280 ;
  assign n26282 = \pi0790  & n26281 ;
  assign n26283 = ~\pi0644  & n26247 ;
  assign n26284 = \pi0790  & ~n26283 ;
  assign n26285 = n23065 & ~n26243 ;
  assign n26286 = ~n26284 & ~n26285 ;
  assign n26287 = \pi0715  & ~n26286 ;
  assign n26288 = ~\pi0644  & n26287 ;
  assign n26289 = ~n25970 & n26287 ;
  assign n26290 = n25965 & n26289 ;
  assign n26291 = ~n26288 & ~n26290 ;
  assign n26292 = ~n26282 & n26291 ;
  assign n26293 = n23074 & ~n26282 ;
  assign n26294 = ~n26041 & n26293 ;
  assign n26295 = ~n26292 & ~n26294 ;
  assign n26296 = n26238 & n26295 ;
  assign n26297 = ~n26268 & n26296 ;
  assign n26298 = ~n26239 & ~n26297 ;
  assign n26299 = \pi0145  & ~\pi0832  ;
  assign n26300 = ~n21132 & ~n26299 ;
  assign n26301 = ~\pi0698  & n1689 ;
  assign n26302 = n20855 & n26301 ;
  assign n26303 = ~\pi0145  & ~n1689 ;
  assign n26304 = ~\pi0778  & ~n26303 ;
  assign n26305 = ~n26302 & n26304 ;
  assign n26306 = ~\pi0778  & ~n26305 ;
  assign n26307 = ~\pi0625  & ~\pi0698  ;
  assign n26308 = n1689 & n26307 ;
  assign n26309 = n20855 & n26308 ;
  assign n26310 = \pi1153  & n26309 ;
  assign n26311 = \pi1153  & ~n26303 ;
  assign n26312 = ~n26302 & n26311 ;
  assign n26313 = ~n26310 & ~n26312 ;
  assign n26314 = ~\pi1153  & ~n26303 ;
  assign n26315 = ~n26309 & n26314 ;
  assign n26316 = ~n26305 & ~n26315 ;
  assign n26317 = n26313 & n26316 ;
  assign n26318 = ~n26306 & ~n26317 ;
  assign n26319 = n20879 & n20895 ;
  assign n26320 = ~n26318 & n26319 ;
  assign n26321 = ~\pi0145  & \pi0647  ;
  assign n26322 = ~n1689 & n26321 ;
  assign n26323 = ~\pi1157  & ~n26322 ;
  assign n26324 = ~n26320 & n26323 ;
  assign n26325 = n20879 & n24830 ;
  assign n26326 = ~n26318 & n26325 ;
  assign n26327 = ~\pi0145  & ~\pi0647  ;
  assign n26328 = ~n1689 & n26327 ;
  assign n26329 = \pi1157  & ~n26328 ;
  assign n26330 = ~n26326 & n26329 ;
  assign n26331 = ~n26324 & ~n26330 ;
  assign n26332 = \pi0787  & ~n26331 ;
  assign n26333 = n20879 & n20891 ;
  assign n26334 = ~n26318 & n26333 ;
  assign n26335 = ~\pi0787  & ~n26334 ;
  assign n26336 = ~\pi1160  & ~n26335 ;
  assign n26337 = n23312 & n26336 ;
  assign n26338 = ~n26332 & n26337 ;
  assign n26339 = ~n21032 & ~n26303 ;
  assign n26340 = \pi0789  & n26339 ;
  assign n26341 = ~\pi0788  & ~n26340 ;
  assign n26342 = n23423 & n26341 ;
  assign n26343 = ~\pi0767  & n1689 ;
  assign n26344 = n20784 & n26343 ;
  assign n26345 = ~n26303 & ~n26344 ;
  assign n26346 = n20794 & ~n26345 ;
  assign n26347 = n20796 & ~n26346 ;
  assign n26348 = n20799 & ~n26345 ;
  assign n26349 = n20801 & ~n26348 ;
  assign n26350 = ~n26347 & ~n26349 ;
  assign n26351 = ~\pi0785  & ~n26303 ;
  assign n26352 = ~n26344 & n26351 ;
  assign n26353 = ~n20804 & ~n26352 ;
  assign n26354 = ~n20812 & n26353 ;
  assign n26355 = n26341 & n26354 ;
  assign n26356 = n26350 & n26355 ;
  assign n26357 = ~n26342 & ~n26356 ;
  assign n26358 = ~n20846 & ~n26357 ;
  assign n26359 = ~n20778 & n26303 ;
  assign n26360 = n24737 & n26359 ;
  assign n26361 = n23423 & ~n26340 ;
  assign n26362 = ~n26340 & n26354 ;
  assign n26363 = n26350 & n26362 ;
  assign n26364 = ~n26361 & ~n26363 ;
  assign n26365 = n24875 & ~n26364 ;
  assign n26366 = ~n26360 & ~n26365 ;
  assign n26367 = ~n26358 & n26366 ;
  assign n26368 = n24884 & ~n26367 ;
  assign n26369 = ~n26338 & ~n26368 ;
  assign n26370 = n24880 & ~n26367 ;
  assign n26371 = ~n23414 & n26303 ;
  assign n26372 = ~n24886 & n26371 ;
  assign n26373 = \pi1160  & n23313 ;
  assign n26374 = ~n26335 & n26373 ;
  assign n26375 = ~n26332 & n26374 ;
  assign n26376 = ~n26372 & ~n26375 ;
  assign n26377 = ~n26370 & n26376 ;
  assign n26378 = n26369 & n26377 ;
  assign n26379 = \pi0790  & ~n26378 ;
  assign n26380 = n26300 & n26379 ;
  assign n26381 = ~n21067 & n23856 ;
  assign n26382 = n20967 & ~n26318 ;
  assign n26383 = n20964 & n26353 ;
  assign n26384 = n26350 & n26383 ;
  assign n26385 = \pi0627  & ~n26384 ;
  assign n26386 = ~n26382 & n26385 ;
  assign n26387 = n20974 & n26353 ;
  assign n26388 = n26350 & n26387 ;
  assign n26389 = ~\pi0627  & ~n26306 ;
  assign n26390 = ~n26317 & n26389 ;
  assign n26391 = ~n20978 & ~n26390 ;
  assign n26392 = ~n26388 & ~n26391 ;
  assign n26393 = \pi0781  & ~n26392 ;
  assign n26394 = ~n26386 & n26393 ;
  assign n26395 = ~n21034 & ~n26394 ;
  assign n26396 = ~n20876 & n26339 ;
  assign n26397 = ~n24969 & ~n26396 ;
  assign n26398 = n26354 & ~n26396 ;
  assign n26399 = n26350 & n26398 ;
  assign n26400 = ~n26397 & ~n26399 ;
  assign n26401 = n21050 & ~n26306 ;
  assign n26402 = ~n26317 & n26401 ;
  assign n26403 = ~n21051 & ~n26402 ;
  assign n26404 = ~n21038 & n26403 ;
  assign n26405 = ~n26400 & n26404 ;
  assign n26406 = ~n23177 & ~n26405 ;
  assign n26407 = ~n26395 & ~n26406 ;
  assign n26408 = ~n26302 & ~n26303 ;
  assign n26409 = n26147 & ~n26408 ;
  assign n26410 = ~\pi0698  & ~n20784 ;
  assign n26411 = n22113 & n26410 ;
  assign n26412 = n26345 & ~n26411 ;
  assign n26413 = ~n26409 & ~n26412 ;
  assign n26414 = n26314 & ~n26413 ;
  assign n26415 = ~\pi0608  & \pi0778  ;
  assign n26416 = n26313 & n26415 ;
  assign n26417 = ~n26414 & n26416 ;
  assign n26418 = \pi0608  & ~n26315 ;
  assign n26419 = n26311 & ~n26344 ;
  assign n26420 = \pi0778  & ~n26419 ;
  assign n26421 = \pi0778  & n26147 ;
  assign n26422 = ~n26408 & n26421 ;
  assign n26423 = ~n26420 & ~n26422 ;
  assign n26424 = n26418 & ~n26423 ;
  assign n26425 = ~\pi0778  & ~n26412 ;
  assign n26426 = ~\pi0785  & ~n26425 ;
  assign n26427 = ~n26424 & n26426 ;
  assign n26428 = ~n26417 & n26427 ;
  assign n26429 = n21022 & ~n26428 ;
  assign n26430 = ~n26406 & n26429 ;
  assign n26431 = ~\pi1155  & ~n26306 ;
  assign n26432 = ~n26317 & n26431 ;
  assign n26433 = ~n20999 & ~n26432 ;
  assign n26434 = \pi1155  & ~n26348 ;
  assign n26435 = ~\pi0660  & ~n26434 ;
  assign n26436 = n26433 & n26435 ;
  assign n26437 = ~n26424 & ~n26425 ;
  assign n26438 = ~n26417 & n26437 ;
  assign n26439 = ~\pi0609  & ~\pi0660  ;
  assign n26440 = ~n26434 & n26439 ;
  assign n26441 = ~n26438 & n26440 ;
  assign n26442 = ~n26436 & ~n26441 ;
  assign n26443 = ~\pi1155  & ~n26346 ;
  assign n26444 = \pi0609  & \pi0660  ;
  assign n26445 = ~n26443 & n26444 ;
  assign n26446 = ~n26438 & n26445 ;
  assign n26447 = \pi0660  & ~n26443 ;
  assign n26448 = \pi1155  & ~n26306 ;
  assign n26449 = ~n26317 & n26448 ;
  assign n26450 = ~n21774 & ~n26449 ;
  assign n26451 = n26447 & n26450 ;
  assign n26452 = \pi0785  & ~n26451 ;
  assign n26453 = ~n26446 & n26452 ;
  assign n26454 = n26442 & n26453 ;
  assign n26455 = n26430 & ~n26454 ;
  assign n26456 = ~n26407 & ~n26455 ;
  assign n26457 = n20778 & ~n26364 ;
  assign n26458 = n20879 & n20951 ;
  assign n26459 = ~n26318 & n26458 ;
  assign n26460 = ~n26359 & ~n26459 ;
  assign n26461 = ~n26457 & n26460 ;
  assign n26462 = n20883 & ~n26459 ;
  assign n26463 = \pi0788  & ~n26462 ;
  assign n26464 = ~n26461 & n26463 ;
  assign n26465 = ~n21067 & ~n26464 ;
  assign n26466 = n26456 & n26465 ;
  assign n26467 = ~n26381 & ~n26466 ;
  assign n26468 = \pi0788  & n20886 ;
  assign n26469 = n26359 & n26468 ;
  assign n26470 = n20778 & n26468 ;
  assign n26471 = ~n26364 & n26470 ;
  assign n26472 = ~n26469 & ~n26471 ;
  assign n26473 = n20886 & ~n26357 ;
  assign n26474 = n20879 & n20938 ;
  assign n26475 = ~n26318 & n26474 ;
  assign n26476 = \pi0629  & ~n26475 ;
  assign n26477 = ~n26473 & n26476 ;
  assign n26478 = n26472 & n26477 ;
  assign n26479 = \pi0788  & n20887 ;
  assign n26480 = n26359 & n26479 ;
  assign n26481 = n20778 & n26479 ;
  assign n26482 = ~n26364 & n26481 ;
  assign n26483 = ~n26480 & ~n26482 ;
  assign n26484 = n20887 & ~n26357 ;
  assign n26485 = n20879 & n21077 ;
  assign n26486 = ~n26318 & n26485 ;
  assign n26487 = ~\pi0629  & ~n26486 ;
  assign n26488 = ~n26484 & n26487 ;
  assign n26489 = n26483 & n26488 ;
  assign n26490 = \pi0792  & ~n26489 ;
  assign n26491 = ~n26478 & n26490 ;
  assign n26492 = \pi0832  & ~n26491 ;
  assign n26493 = ~n26467 & n26492 ;
  assign n26494 = ~\pi0145  & \pi0792  ;
  assign n26495 = ~n1689 & n26494 ;
  assign n26496 = ~n20845 & n26495 ;
  assign n26497 = ~n24996 & ~n26496 ;
  assign n26498 = ~n26358 & n26497 ;
  assign n26499 = n26366 & n26498 ;
  assign n26500 = \pi0630  & n26323 ;
  assign n26501 = ~n26320 & n26500 ;
  assign n26502 = n20849 & ~n26328 ;
  assign n26503 = ~n26326 & n26502 ;
  assign n26504 = ~n26501 & ~n26503 ;
  assign n26505 = \pi0787  & ~n26504 ;
  assign n26506 = ~n24761 & ~n26505 ;
  assign n26507 = ~n26499 & n26506 ;
  assign n26508 = \pi0832  & ~n26507 ;
  assign n26509 = n26300 & ~n26508 ;
  assign n26510 = ~n26493 & n26509 ;
  assign n26511 = ~n26380 & ~n26510 ;
  assign n26512 = \pi0038  & n26344 ;
  assign n26513 = n8413 & n26512 ;
  assign n26514 = n1354 & n26513 ;
  assign n26515 = n1358 & n26514 ;
  assign n26516 = \pi0038  & ~\pi0145  ;
  assign n26517 = ~n21757 & n26516 ;
  assign n26518 = ~n26515 & ~n26517 ;
  assign n26519 = \pi0038  & n26518 ;
  assign n26520 = ~\pi0145  & ~n21467 ;
  assign n26521 = ~\pi0039  & ~\pi0145  ;
  assign n26522 = n21272 & n26521 ;
  assign n26523 = ~n26520 & ~n26522 ;
  assign n26524 = ~\pi0145  & ~\pi0767  ;
  assign n26525 = ~\pi0767  & n25023 ;
  assign n26526 = ~n26524 & ~n26525 ;
  assign n26527 = n26523 & ~n26526 ;
  assign n26528 = ~\pi0145  & \pi0767  ;
  assign n26529 = n21743 & n26528 ;
  assign n26530 = ~n21734 & n26529 ;
  assign n26531 = n26518 & ~n26530 ;
  assign n26532 = ~n26527 & n26531 ;
  assign n26533 = ~n26519 & ~n26532 ;
  assign n26534 = \pi0698  & n26533 ;
  assign n26535 = ~\pi0145  & ~\pi0778  ;
  assign n26536 = ~n23622 & ~n26535 ;
  assign n26537 = n26534 & ~n26536 ;
  assign n26538 = n23557 & ~n23558 ;
  assign n26539 = \pi0145  & ~n26538 ;
  assign n26540 = ~\pi0039  & ~n22683 ;
  assign n26541 = ~\pi0145  & n23548 ;
  assign n26542 = ~n26540 & n26541 ;
  assign n26543 = ~\pi0767  & ~n26542 ;
  assign n26544 = ~n26539 & n26543 ;
  assign n26545 = ~\pi0038  & ~n26544 ;
  assign n26546 = ~\pi0145  & ~n23567 ;
  assign n26547 = n23565 & n26546 ;
  assign n26548 = \pi0767  & n23575 ;
  assign n26549 = n23572 & n26548 ;
  assign n26550 = ~n26528 & ~n26549 ;
  assign n26551 = ~n26547 & ~n26550 ;
  assign n26552 = n6861 & ~n26551 ;
  assign n26553 = n26545 & n26552 ;
  assign n26554 = n1354 & n8413 ;
  assign n26555 = \pi0145  & \pi0603  ;
  assign n26556 = ~n20783 & n26555 ;
  assign n26557 = n26343 & n26556 ;
  assign n26558 = \pi0145  & ~n20784 ;
  assign n26559 = n22113 & n26558 ;
  assign n26560 = ~n26557 & ~n26559 ;
  assign n26561 = n26554 & ~n26560 ;
  assign n26562 = n1358 & n26561 ;
  assign n26563 = \pi0038  & ~n26562 ;
  assign n26564 = ~\pi0698  & ~n26563 ;
  assign n26565 = n1354 & n25206 ;
  assign n26566 = n1358 & n26565 ;
  assign n26567 = ~\pi0145  & ~\pi0698  ;
  assign n26568 = ~n26566 & n26567 ;
  assign n26569 = ~\pi0767  & n26567 ;
  assign n26570 = ~n22536 & n26569 ;
  assign n26571 = ~n26568 & ~n26570 ;
  assign n26572 = ~n26564 & n26571 ;
  assign n26573 = n6861 & n26572 ;
  assign n26574 = ~n26536 & ~n26573 ;
  assign n26575 = ~n26553 & n26574 ;
  assign n26576 = ~n26537 & ~n26575 ;
  assign n26577 = \pi0609  & ~n26576 ;
  assign n26578 = ~\pi0145  & ~\pi0625  ;
  assign n26579 = ~n22734 & ~n26578 ;
  assign n26580 = n26534 & ~n26579 ;
  assign n26581 = ~n26573 & ~n26579 ;
  assign n26582 = ~n26553 & n26581 ;
  assign n26583 = ~n26580 & ~n26582 ;
  assign n26584 = n6861 & ~n26533 ;
  assign n26585 = ~\pi0145  & \pi0625  ;
  assign n26586 = ~n22727 & ~n26585 ;
  assign n26587 = ~n26584 & ~n26586 ;
  assign n26588 = ~\pi1153  & ~n26587 ;
  assign n26589 = n26583 & n26588 ;
  assign n26590 = ~\pi0074  & ~\pi0698  ;
  assign n26591 = ~\pi0100  & n26590 ;
  assign n26592 = n1287 & n26591 ;
  assign n26593 = ~\pi0145  & ~n26592 ;
  assign n26594 = n21768 & n26593 ;
  assign n26595 = n21770 & n26593 ;
  assign n26596 = ~n21734 & n26595 ;
  assign n26597 = ~n26594 & ~n26596 ;
  assign n26598 = \pi0625  & ~n26597 ;
  assign n26599 = ~\pi0145  & ~n22017 ;
  assign n26600 = ~n21994 & n26599 ;
  assign n26601 = ~\pi0038  & ~\pi0145  ;
  assign n26602 = n6861 & ~n26601 ;
  assign n26603 = ~n22109 & n26602 ;
  assign n26604 = ~n26600 & ~n26603 ;
  assign n26605 = ~\pi0145  & ~n21757 ;
  assign n26606 = n22117 & ~n26605 ;
  assign n26607 = ~\pi0698  & ~n26606 ;
  assign n26608 = \pi0625  & n26607 ;
  assign n26609 = ~n26604 & n26608 ;
  assign n26610 = ~n26598 & ~n26609 ;
  assign n26611 = n21768 & n26578 ;
  assign n26612 = n21770 & n26578 ;
  assign n26613 = ~n21734 & n26612 ;
  assign n26614 = ~n26611 & ~n26613 ;
  assign n26615 = \pi1153  & n26614 ;
  assign n26616 = n26610 & n26615 ;
  assign n26617 = ~\pi0608  & ~n26616 ;
  assign n26618 = ~n26589 & n26617 ;
  assign n26619 = n26534 & ~n26586 ;
  assign n26620 = ~n26573 & ~n26586 ;
  assign n26621 = ~n26553 & n26620 ;
  assign n26622 = ~n26619 & ~n26621 ;
  assign n26623 = \pi1153  & n26579 ;
  assign n26624 = n23606 & ~n26533 ;
  assign n26625 = ~n26623 & ~n26624 ;
  assign n26626 = n26622 & ~n26625 ;
  assign n26627 = ~\pi0625  & ~n26597 ;
  assign n26628 = ~\pi0625  & n26607 ;
  assign n26629 = ~n26604 & n26628 ;
  assign n26630 = ~n26627 & ~n26629 ;
  assign n26631 = n21768 & n26585 ;
  assign n26632 = n21770 & n26585 ;
  assign n26633 = ~n21734 & n26632 ;
  assign n26634 = ~n26631 & ~n26633 ;
  assign n26635 = ~\pi1153  & n26634 ;
  assign n26636 = n26630 & n26635 ;
  assign n26637 = \pi0608  & ~n26636 ;
  assign n26638 = ~n26626 & n26637 ;
  assign n26639 = ~n26618 & ~n26638 ;
  assign n26640 = n23638 & ~n26639 ;
  assign n26641 = ~n26577 & ~n26640 ;
  assign n26642 = \pi0145  & ~n6861 ;
  assign n26643 = ~n20985 & n26642 ;
  assign n26644 = n21774 & n26643 ;
  assign n26645 = n6861 & ~n20985 ;
  assign n26646 = n21774 & n26645 ;
  assign n26647 = ~n26533 & n26646 ;
  assign n26648 = ~n26644 & ~n26647 ;
  assign n26649 = ~\pi0145  & n21768 ;
  assign n26650 = ~\pi0145  & n21770 ;
  assign n26651 = ~n21734 & n26650 ;
  assign n26652 = ~n26649 & ~n26651 ;
  assign n26653 = \pi1155  & ~n22788 ;
  assign n26654 = n26652 & n26653 ;
  assign n26655 = ~\pi0660  & ~n26654 ;
  assign n26656 = n26648 & n26655 ;
  assign n26657 = ~n26604 & n26607 ;
  assign n26658 = ~\pi0778  & n26597 ;
  assign n26659 = ~n26657 & n26658 ;
  assign n26660 = ~\pi0609  & ~n26659 ;
  assign n26661 = \pi1155  & ~n26660 ;
  assign n26662 = ~n26616 & ~n26636 ;
  assign n26663 = n22722 & ~n26662 ;
  assign n26664 = ~n26661 & ~n26663 ;
  assign n26665 = ~n26656 & ~n26664 ;
  assign n26666 = n26641 & n26665 ;
  assign n26667 = \pi0778  & ~n26639 ;
  assign n26668 = \pi0778  & ~n26662 ;
  assign n26669 = \pi0609  & ~n26659 ;
  assign n26670 = ~n26668 & n26669 ;
  assign n26671 = ~\pi1155  & n26643 ;
  assign n26672 = ~\pi1155  & n26645 ;
  assign n26673 = ~n26533 & n26672 ;
  assign n26674 = ~n26671 & ~n26673 ;
  assign n26675 = ~\pi0609  & ~n26674 ;
  assign n26676 = ~\pi1155  & ~n22767 ;
  assign n26677 = n26652 & n26676 ;
  assign n26678 = ~n22787 & ~n26677 ;
  assign n26679 = ~n26675 & n26678 ;
  assign n26680 = ~n26670 & ~n26679 ;
  assign n26681 = \pi0785  & ~n26680 ;
  assign n26682 = n26576 & ~n26681 ;
  assign n26683 = ~n26667 & n26682 ;
  assign n26684 = n20999 & n26643 ;
  assign n26685 = n20999 & n26645 ;
  assign n26686 = ~n26533 & n26685 ;
  assign n26687 = ~n26684 & ~n26686 ;
  assign n26688 = \pi0660  & ~n26677 ;
  assign n26689 = n26687 & n26688 ;
  assign n26690 = ~n26656 & ~n26689 ;
  assign n26691 = \pi0609  & ~n26678 ;
  assign n26692 = n26659 & n26691 ;
  assign n26693 = \pi0778  & n26691 ;
  assign n26694 = ~n26662 & n26693 ;
  assign n26695 = ~n26692 & ~n26694 ;
  assign n26696 = ~n26690 & n26695 ;
  assign n26697 = ~n26683 & n26696 ;
  assign n26698 = ~n26666 & n26697 ;
  assign n26699 = ~\pi0785  & ~n26683 ;
  assign n26700 = n21022 & ~n21034 ;
  assign n26701 = ~n26699 & n26700 ;
  assign n26702 = ~n26698 & n26701 ;
  assign n26703 = ~\pi0145  & ~n20778 ;
  assign n26704 = n21768 & n26703 ;
  assign n26705 = n21770 & n26703 ;
  assign n26706 = ~n21734 & n26705 ;
  assign n26707 = ~n26704 & ~n26706 ;
  assign n26708 = \pi0788  & ~n26707 ;
  assign n26709 = n23456 & ~n26533 ;
  assign n26710 = ~n21777 & n26652 ;
  assign n26711 = ~\pi0781  & ~n26710 ;
  assign n26712 = n21777 & n26642 ;
  assign n26713 = ~n23423 & ~n26712 ;
  assign n26714 = n26711 & n26713 ;
  assign n26715 = ~n26709 & n26714 ;
  assign n26716 = n23423 & ~n26652 ;
  assign n26717 = ~n26715 & ~n26716 ;
  assign n26718 = n20816 & ~n26717 ;
  assign n26719 = ~\pi0145  & ~n20811 ;
  assign n26720 = n21768 & n26719 ;
  assign n26721 = n21770 & n26719 ;
  assign n26722 = ~n21734 & n26721 ;
  assign n26723 = ~n26720 & ~n26722 ;
  assign n26724 = n20811 & ~n26710 ;
  assign n26725 = ~n26712 & n26724 ;
  assign n26726 = ~n26709 & n26725 ;
  assign n26727 = n26723 & ~n26726 ;
  assign n26728 = n20816 & n23424 ;
  assign n26729 = ~n26727 & n26728 ;
  assign n26730 = ~n26718 & ~n26729 ;
  assign n26731 = ~n26708 & n26730 ;
  assign n26732 = ~\pi0788  & ~n26717 ;
  assign n26733 = ~\pi0788  & n23424 ;
  assign n26734 = ~n26727 & n26733 ;
  assign n26735 = ~n26732 & ~n26734 ;
  assign n26736 = n24691 & n26735 ;
  assign n26737 = n26731 & n26736 ;
  assign n26738 = n26065 & ~n26662 ;
  assign n26739 = ~\pi0778  & n23885 ;
  assign n26740 = n26597 & n26739 ;
  assign n26741 = ~n26657 & n26740 ;
  assign n26742 = ~n23885 & n26652 ;
  assign n26743 = ~\pi0628  & ~n26742 ;
  assign n26744 = ~n26741 & n26743 ;
  assign n26745 = ~n26738 & n26744 ;
  assign n26746 = ~\pi0145  & \pi0628  ;
  assign n26747 = n21768 & n26746 ;
  assign n26748 = n21770 & n26746 ;
  assign n26749 = ~n21734 & n26748 ;
  assign n26750 = ~n26747 & ~n26749 ;
  assign n26751 = n20844 & n26750 ;
  assign n26752 = ~n26745 & n26751 ;
  assign n26753 = \pi0628  & ~n26742 ;
  assign n26754 = ~n26741 & n26753 ;
  assign n26755 = ~n26738 & n26754 ;
  assign n26756 = ~\pi0145  & ~\pi0628  ;
  assign n26757 = n21768 & n26756 ;
  assign n26758 = n21770 & n26756 ;
  assign n26759 = ~n21734 & n26758 ;
  assign n26760 = ~n26757 & ~n26759 ;
  assign n26761 = n20843 & n26760 ;
  assign n26762 = ~n26755 & n26761 ;
  assign n26763 = ~n26752 & ~n26762 ;
  assign n26764 = ~n26737 & n26763 ;
  assign n26765 = \pi0792  & ~n26764 ;
  assign n26766 = n23380 & ~n26659 ;
  assign n26767 = n21768 & ~n23380 ;
  assign n26768 = n21770 & ~n23380 ;
  assign n26769 = ~n21734 & n26768 ;
  assign n26770 = ~n26767 & ~n26769 ;
  assign n26771 = ~\pi0145  & ~n26770 ;
  assign n26772 = n21050 & ~n26771 ;
  assign n26773 = ~n26766 & n26772 ;
  assign n26774 = \pi0778  & n26772 ;
  assign n26775 = ~n26662 & n26774 ;
  assign n26776 = ~n26773 & ~n26775 ;
  assign n26777 = \pi0789  & ~n26776 ;
  assign n26778 = n23683 & ~n26727 ;
  assign n26779 = n21032 & ~n26712 ;
  assign n26780 = n26711 & n26779 ;
  assign n26781 = ~n26709 & n26780 ;
  assign n26782 = ~n21032 & ~n26652 ;
  assign n26783 = ~n20876 & ~n26782 ;
  assign n26784 = ~n26781 & n26783 ;
  assign n26785 = \pi0789  & n26784 ;
  assign n26786 = ~n26778 & n26785 ;
  assign n26787 = ~n26777 & ~n26786 ;
  assign n26788 = n22155 & n26723 ;
  assign n26789 = ~n26726 & n26788 ;
  assign n26790 = ~n22147 & ~n26659 ;
  assign n26791 = n22147 & ~n26652 ;
  assign n26792 = n24348 & ~n26791 ;
  assign n26793 = ~n26790 & n26792 ;
  assign n26794 = \pi0778  & n26792 ;
  assign n26795 = ~n26662 & n26794 ;
  assign n26796 = ~n26793 & ~n26795 ;
  assign n26797 = ~n26789 & n26796 ;
  assign n26798 = ~n21034 & ~n26797 ;
  assign n26799 = ~n21038 & ~n26798 ;
  assign n26800 = n26787 & n26799 ;
  assign n26801 = ~n26765 & n26800 ;
  assign n26802 = ~n26702 & n26801 ;
  assign n26803 = ~\pi0788  & ~n23856 ;
  assign n26804 = ~n20883 & ~n26707 ;
  assign n26805 = n20947 & ~n26717 ;
  assign n26806 = n20947 & n23424 ;
  assign n26807 = ~n26727 & n26806 ;
  assign n26808 = ~n26805 & ~n26807 ;
  assign n26809 = ~n26804 & n26808 ;
  assign n26810 = ~n22160 & ~n26771 ;
  assign n26811 = ~n26766 & n26810 ;
  assign n26812 = \pi0778  & n26810 ;
  assign n26813 = ~n26662 & n26812 ;
  assign n26814 = ~n26811 & ~n26813 ;
  assign n26815 = n20951 & ~n26652 ;
  assign n26816 = ~n23838 & ~n26815 ;
  assign n26817 = n26814 & ~n26816 ;
  assign n26818 = ~n23856 & ~n26817 ;
  assign n26819 = n26809 & n26818 ;
  assign n26820 = ~n26803 & ~n26819 ;
  assign n26821 = ~n26765 & n26820 ;
  assign n26822 = ~n21067 & ~n26821 ;
  assign n26823 = ~n26802 & n26822 ;
  assign n26824 = \pi0644  & \pi1160  ;
  assign n26825 = ~\pi0145  & ~\pi0644  ;
  assign n26826 = n21768 & n26825 ;
  assign n26827 = n21770 & n26825 ;
  assign n26828 = ~n21734 & n26827 ;
  assign n26829 = ~n26826 & ~n26828 ;
  assign n26830 = ~\pi0715  & n26829 ;
  assign n26831 = n26824 & ~n26830 ;
  assign n26832 = n21092 & n26735 ;
  assign n26833 = n26731 & n26832 ;
  assign n26834 = ~n21092 & n26652 ;
  assign n26835 = n26824 & ~n26834 ;
  assign n26836 = ~n26833 & n26835 ;
  assign n26837 = ~n26831 & ~n26836 ;
  assign n26838 = \pi0790  & n26837 ;
  assign n26839 = ~n26741 & ~n26742 ;
  assign n26840 = ~n26738 & n26839 ;
  assign n26841 = ~\pi0792  & ~n26840 ;
  assign n26842 = ~\pi0647  & ~n26841 ;
  assign n26843 = n21768 & n26321 ;
  assign n26844 = n21770 & n26321 ;
  assign n26845 = ~n21734 & n26844 ;
  assign n26846 = ~n26843 & ~n26845 ;
  assign n26847 = n20897 & n26846 ;
  assign n26848 = ~n26842 & n26847 ;
  assign n26849 = \pi1156  & n26760 ;
  assign n26850 = ~n26755 & n26849 ;
  assign n26851 = ~\pi1156  & n26750 ;
  assign n26852 = ~n26745 & n26851 ;
  assign n26853 = ~n26850 & ~n26852 ;
  assign n26854 = \pi0792  & n26847 ;
  assign n26855 = ~n26853 & n26854 ;
  assign n26856 = ~n26848 & ~n26855 ;
  assign n26857 = n20846 & ~n26652 ;
  assign n26858 = ~n20910 & ~n26857 ;
  assign n26859 = n20846 & n26858 ;
  assign n26860 = n26735 & n26858 ;
  assign n26861 = n26731 & n26860 ;
  assign n26862 = ~n26859 & ~n26861 ;
  assign n26863 = \pi0647  & ~n26841 ;
  assign n26864 = n21768 & n26327 ;
  assign n26865 = n21770 & n26327 ;
  assign n26866 = ~n21734 & n26865 ;
  assign n26867 = ~n26864 & ~n26866 ;
  assign n26868 = n20849 & n26867 ;
  assign n26869 = ~n26863 & n26868 ;
  assign n26870 = \pi0792  & n26868 ;
  assign n26871 = ~n26853 & n26870 ;
  assign n26872 = ~n26869 & ~n26871 ;
  assign n26873 = n26862 & n26872 ;
  assign n26874 = n26856 & n26873 ;
  assign n26875 = \pi0787  & ~n26874 ;
  assign n26876 = ~n26838 & ~n26875 ;
  assign n26877 = ~n26823 & n26876 ;
  assign n26878 = n9948 & n26379 ;
  assign n26879 = n9948 & ~n26508 ;
  assign n26880 = ~n26493 & n26879 ;
  assign n26881 = ~n26878 & ~n26880 ;
  assign n26882 = n26877 & ~n26881 ;
  assign n26883 = ~\pi0787  & n26841 ;
  assign n26884 = n23011 & ~n26853 ;
  assign n26885 = ~n26883 & ~n26884 ;
  assign n26886 = \pi0644  & ~n26885 ;
  assign n26887 = \pi1157  & n26867 ;
  assign n26888 = ~n26863 & n26887 ;
  assign n26889 = \pi0792  & n26887 ;
  assign n26890 = ~n26853 & n26889 ;
  assign n26891 = ~n26888 & ~n26890 ;
  assign n26892 = ~\pi1157  & n26846 ;
  assign n26893 = ~n26842 & n26892 ;
  assign n26894 = \pi0792  & n26892 ;
  assign n26895 = ~n26853 & n26894 ;
  assign n26896 = ~n26893 & ~n26895 ;
  assign n26897 = n26891 & n26896 ;
  assign n26898 = n23074 & ~n26897 ;
  assign n26899 = ~n26886 & ~n26898 ;
  assign n26900 = \pi0644  & n26899 ;
  assign n26901 = ~n26875 & n26899 ;
  assign n26902 = ~n26823 & n26901 ;
  assign n26903 = ~n26900 & ~n26902 ;
  assign n26904 = n23316 & ~n26903 ;
  assign n26905 = ~\pi0145  & \pi0715  ;
  assign n26906 = n21768 & n26905 ;
  assign n26907 = n21770 & n26905 ;
  assign n26908 = ~n21734 & n26907 ;
  assign n26909 = ~n26906 & ~n26908 ;
  assign n26910 = ~n23313 & n26909 ;
  assign n26911 = \pi0644  & ~\pi1160  ;
  assign n26912 = ~\pi1160  & ~n26834 ;
  assign n26913 = ~n26833 & n26912 ;
  assign n26914 = ~n26911 & ~n26913 ;
  assign n26915 = ~n26910 & ~n26914 ;
  assign n26916 = ~\pi0644  & n26885 ;
  assign n26917 = \pi0715  & ~n26916 ;
  assign n26918 = \pi0715  & \pi0787  ;
  assign n26919 = ~n26897 & n26918 ;
  assign n26920 = ~n26917 & ~n26919 ;
  assign n26921 = \pi1160  & ~n26830 ;
  assign n26922 = ~n26836 & ~n26921 ;
  assign n26923 = n26920 & ~n26922 ;
  assign n26924 = ~n26915 & ~n26923 ;
  assign n26925 = ~n26904 & n26924 ;
  assign n26926 = \pi0790  & ~n26881 ;
  assign n26927 = ~n26925 & n26926 ;
  assign n26928 = ~n26882 & ~n26927 ;
  assign n26929 = n26511 & n26928 ;
  assign n26930 = \pi0907  & ~\pi0947  ;
  assign n26931 = \pi0735  & n26930 ;
  assign n26932 = \pi0743  & \pi0947  ;
  assign n26933 = n1689 & ~n26932 ;
  assign n26934 = ~n26931 & n26933 ;
  assign n26935 = ~\pi0146  & ~n1689 ;
  assign n26936 = \pi0832  & ~n26935 ;
  assign n26937 = ~n26934 & n26936 ;
  assign n26938 = ~\pi0146  & ~n21757 ;
  assign n26939 = n1354 & n1356 ;
  assign n26940 = n8413 & n26934 ;
  assign n26941 = n26939 & n26940 ;
  assign n26942 = n10323 & n26941 ;
  assign n26943 = \pi0038  & ~n26942 ;
  assign n26944 = ~n26938 & n26943 ;
  assign n26945 = n11834 & ~n26944 ;
  assign n26946 = ~\pi0146  & n21740 ;
  assign n26947 = ~\pi0146  & n21737 ;
  assign n26948 = n21232 & n26947 ;
  assign n26949 = ~n26946 & ~n26948 ;
  assign n26950 = ~\pi0299  & n26949 ;
  assign n26951 = ~n26931 & ~n26932 ;
  assign n26952 = ~n21740 & n26951 ;
  assign n26953 = ~n21738 & n26952 ;
  assign n26954 = n26950 & ~n26953 ;
  assign n26955 = ~n21205 & n26951 ;
  assign n26956 = ~n21238 & n26955 ;
  assign n26957 = \pi0299  & ~n21205 ;
  assign n26958 = ~n11696 & ~n26957 ;
  assign n26959 = ~n11696 & n21237 ;
  assign n26960 = n21232 & n26959 ;
  assign n26961 = ~n26958 & ~n26960 ;
  assign n26962 = ~n26956 & n26961 ;
  assign n26963 = ~\pi0039  & ~n26962 ;
  assign n26964 = ~n26954 & n26963 ;
  assign n26965 = ~\pi0038  & ~n26964 ;
  assign n26966 = n26945 & ~n26965 ;
  assign n26967 = n21711 & ~n26951 ;
  assign n26968 = \pi0146  & ~n21593 ;
  assign n26969 = ~n21709 & n26968 ;
  assign n26970 = n6761 & ~n26969 ;
  assign n26971 = n2165 & ~n26951 ;
  assign n26972 = ~n21285 & n26971 ;
  assign n26973 = \pi0146  & n2165 ;
  assign n26974 = n21285 & n26973 ;
  assign n26975 = ~\pi0223  & ~n26974 ;
  assign n26976 = ~n26972 & n26975 ;
  assign n26977 = \pi0146  & \pi0681  ;
  assign n26978 = n21580 & n26977 ;
  assign n26979 = n26976 & ~n26978 ;
  assign n26980 = n26970 & n26979 ;
  assign n26981 = ~n26967 & n26980 ;
  assign n26982 = ~\pi0146  & ~n6761 ;
  assign n26983 = n21334 & n26982 ;
  assign n26984 = ~n21330 & n26983 ;
  assign n26985 = ~n6761 & n26951 ;
  assign n26986 = ~n21334 & n26985 ;
  assign n26987 = n6713 & n26985 ;
  assign n26988 = ~n21329 & n26987 ;
  assign n26989 = ~n26986 & ~n26988 ;
  assign n26990 = ~n2165 & n26989 ;
  assign n26991 = ~n26984 & n26990 ;
  assign n26992 = n26976 & ~n26991 ;
  assign n26993 = n21627 & ~n26951 ;
  assign n26994 = ~n21726 & n26993 ;
  assign n26995 = ~n6761 & n26994 ;
  assign n26996 = n21627 & ~n21726 ;
  assign n26997 = \pi0146  & ~n6761 ;
  assign n26998 = ~n26996 & n26997 ;
  assign n26999 = ~n26995 & ~n26998 ;
  assign n27000 = ~n21654 & n26951 ;
  assign n27001 = ~n21657 & n27000 ;
  assign n27002 = ~n21684 & n27001 ;
  assign n27003 = \pi0223  & n27002 ;
  assign n27004 = n6761 & ~n21654 ;
  assign n27005 = ~n21657 & n27004 ;
  assign n27006 = ~n21684 & n27005 ;
  assign n27007 = \pi0146  & n6761 ;
  assign n27008 = \pi0223  & ~n27007 ;
  assign n27009 = ~n27006 & n27008 ;
  assign n27010 = ~n27003 & ~n27009 ;
  assign n27011 = n26999 & ~n27010 ;
  assign n27012 = ~n26992 & ~n27011 ;
  assign n27013 = ~n26981 & n27012 ;
  assign n27014 = ~\pi0299  & ~n27013 ;
  assign n27015 = \pi0146  & n6730 ;
  assign n27016 = n21694 & n27015 ;
  assign n27017 = ~n21711 & n27016 ;
  assign n27018 = \pi0146  & ~n6732 ;
  assign n27019 = n21334 & n27018 ;
  assign n27020 = ~n21330 & n27019 ;
  assign n27021 = ~n21334 & ~n26951 ;
  assign n27022 = n6713 & ~n26951 ;
  assign n27023 = ~n21329 & n27022 ;
  assign n27024 = ~n27021 & ~n27023 ;
  assign n27025 = ~n2352 & n27024 ;
  assign n27026 = ~n27020 & n27025 ;
  assign n27027 = ~n27017 & n27026 ;
  assign n27028 = n2352 & ~n26932 ;
  assign n27029 = ~n26931 & n27028 ;
  assign n27030 = ~\pi0215  & ~n27029 ;
  assign n27031 = ~n21285 & n27030 ;
  assign n27032 = ~\pi0146  & n2352 ;
  assign n27033 = ~\pi0215  & ~n27032 ;
  assign n27034 = n21285 & n27033 ;
  assign n27035 = ~n27031 & ~n27034 ;
  assign n27036 = ~n27027 & ~n27035 ;
  assign n27037 = \pi0146  & ~n21728 ;
  assign n27038 = ~n21724 & n27037 ;
  assign n27039 = \pi0299  & ~n26994 ;
  assign n27040 = ~n27038 & n27039 ;
  assign n27041 = ~n21948 & ~n27040 ;
  assign n27042 = ~n27036 & ~n27041 ;
  assign n27043 = ~n27014 & ~n27042 ;
  assign n27044 = \pi0039  & n26945 ;
  assign n27045 = ~n27043 & n27044 ;
  assign n27046 = ~n26966 & ~n27045 ;
  assign n27047 = ~\pi0146  & ~n11834 ;
  assign n27048 = ~\pi0832  & ~n27047 ;
  assign n27049 = n27046 & n27048 ;
  assign n27050 = ~n26937 & ~n27049 ;
  assign n27051 = ~\pi0770  & \pi0947  ;
  assign n27052 = \pi0726  & n26930 ;
  assign n27053 = ~n27051 & ~n27052 ;
  assign n27054 = n1689 & ~n27053 ;
  assign n27055 = ~\pi0147  & ~n1689 ;
  assign n27056 = \pi0832  & ~n27055 ;
  assign n27057 = ~n27054 & n27056 ;
  assign n27058 = ~n21690 & n26930 ;
  assign n27059 = n21688 & n27058 ;
  assign n27060 = ~n21614 & n27059 ;
  assign n27061 = n6205 & ~n27060 ;
  assign n27062 = \pi0299  & n26930 ;
  assign n27063 = ~n21205 & n27062 ;
  assign n27064 = ~n21238 & n27063 ;
  assign n27065 = ~\pi0299  & n26930 ;
  assign n27066 = ~n21740 & n27065 ;
  assign n27067 = ~n21738 & n27066 ;
  assign n27068 = ~n27064 & ~n27067 ;
  assign n27069 = ~\pi0039  & n27068 ;
  assign n27070 = ~n21285 & n26930 ;
  assign n27071 = ~\pi0215  & n2352 ;
  assign n27072 = ~n27070 & n27071 ;
  assign n27073 = \pi0299  & n27072 ;
  assign n27074 = ~n21334 & n26930 ;
  assign n27075 = n6713 & n26930 ;
  assign n27076 = ~n21329 & n27075 ;
  assign n27077 = ~n27074 & ~n27076 ;
  assign n27078 = \pi0299  & n24388 ;
  assign n27079 = n27077 & n27078 ;
  assign n27080 = ~n27073 & ~n27079 ;
  assign n27081 = n21627 & n26930 ;
  assign n27082 = ~n21726 & n27081 ;
  assign n27083 = n2259 & ~n27082 ;
  assign n27084 = n27080 & ~n27083 ;
  assign n27085 = \pi0039  & ~n27084 ;
  assign n27086 = \pi0147  & ~n27085 ;
  assign n27087 = ~n27069 & n27086 ;
  assign n27088 = ~n27061 & n27087 ;
  assign n27089 = ~\pi0038  & ~n27088 ;
  assign n27090 = ~\pi0147  & ~n21757 ;
  assign n27091 = n1689 & n26930 ;
  assign n27092 = n6784 & n27091 ;
  assign n27093 = n1266 & n27092 ;
  assign n27094 = n26939 & n27093 ;
  assign n27095 = n10323 & n27094 ;
  assign n27096 = \pi0038  & ~n27095 ;
  assign n27097 = ~n27090 & n27096 ;
  assign n27098 = \pi0770  & ~n27097 ;
  assign n27099 = ~n27089 & n27098 ;
  assign n27100 = \pi0299  & ~n26930 ;
  assign n27101 = ~n21205 & n27100 ;
  assign n27102 = ~n21238 & n27101 ;
  assign n27103 = ~\pi0299  & ~n26930 ;
  assign n27104 = ~n21740 & n27103 ;
  assign n27105 = ~n21738 & n27104 ;
  assign n27106 = ~n27102 & ~n27105 ;
  assign n27107 = ~\pi0039  & n27106 ;
  assign n27108 = ~\pi0147  & \pi0770  ;
  assign n27109 = ~n27097 & n27108 ;
  assign n27110 = n27107 & n27109 ;
  assign n27111 = \pi0215  & \pi0947  ;
  assign n27112 = \pi0299  & n27111 ;
  assign n27113 = n21627 & n27112 ;
  assign n27114 = ~n21726 & n27113 ;
  assign n27115 = \pi0215  & ~n21724 ;
  assign n27116 = \pi0299  & ~n27115 ;
  assign n27117 = ~n27114 & ~n27116 ;
  assign n27118 = \pi0947  & ~n21334 ;
  assign n27119 = \pi0947  & n6713 ;
  assign n27120 = ~n21329 & n27119 ;
  assign n27121 = ~n27118 & ~n27120 ;
  assign n27122 = ~n2352 & ~n27121 ;
  assign n27123 = ~n21698 & ~n27122 ;
  assign n27124 = n21694 & ~n27122 ;
  assign n27125 = ~n21711 & n27124 ;
  assign n27126 = ~n27123 & ~n27125 ;
  assign n27127 = n2352 & ~n26930 ;
  assign n27128 = ~n21285 & n27127 ;
  assign n27129 = ~\pi0215  & ~n27128 ;
  assign n27130 = ~n27114 & n27129 ;
  assign n27131 = ~n27126 & n27130 ;
  assign n27132 = ~n27117 & ~n27131 ;
  assign n27133 = ~\pi0039  & ~n27106 ;
  assign n27134 = ~n21690 & n27103 ;
  assign n27135 = n21688 & n27134 ;
  assign n27136 = ~n21614 & n27135 ;
  assign n27137 = ~n27133 & ~n27136 ;
  assign n27138 = n27109 & n27137 ;
  assign n27139 = ~n27132 & n27138 ;
  assign n27140 = ~n27110 & ~n27139 ;
  assign n27141 = ~n27099 & n27140 ;
  assign n27142 = n1689 & n6730 ;
  assign n27143 = n4520 & n27142 ;
  assign n27144 = n1638 & n27143 ;
  assign n27145 = ~\pi0147  & ~\pi0770  ;
  assign n27146 = ~n27144 & n27145 ;
  assign n27147 = \pi0726  & \pi0770  ;
  assign n27148 = n1689 & ~n6730 ;
  assign n27149 = n1354 & n27148 ;
  assign n27150 = n8413 & n27149 ;
  assign n27151 = n1358 & n27150 ;
  assign n27152 = \pi0038  & \pi0726  ;
  assign n27153 = ~n27151 & n27152 ;
  assign n27154 = ~n27147 & ~n27153 ;
  assign n27155 = ~n27146 & ~n27154 ;
  assign n27156 = ~n6730 & n21688 ;
  assign n27157 = ~n21690 & n27156 ;
  assign n27158 = ~n21614 & n27157 ;
  assign n27159 = n6205 & ~n27158 ;
  assign n27160 = \pi0299  & ~n6730 ;
  assign n27161 = ~n21205 & n27160 ;
  assign n27162 = ~n21238 & n27161 ;
  assign n27163 = ~\pi0299  & ~n6730 ;
  assign n27164 = ~n21740 & n27163 ;
  assign n27165 = ~n21738 & n27164 ;
  assign n27166 = ~n27162 & ~n27165 ;
  assign n27167 = ~\pi0039  & n27166 ;
  assign n27168 = n2352 & ~n6730 ;
  assign n27169 = ~n21285 & n27168 ;
  assign n27170 = ~\pi0215  & ~n27169 ;
  assign n27171 = n21703 & n27170 ;
  assign n27172 = ~n21729 & ~n27171 ;
  assign n27173 = n2297 & ~n27172 ;
  assign n27174 = \pi0147  & ~n27173 ;
  assign n27175 = ~n27167 & n27174 ;
  assign n27176 = ~n27159 & n27175 ;
  assign n27177 = ~\pi0038  & \pi0726  ;
  assign n27178 = ~n27176 & n27177 ;
  assign n27179 = ~n27155 & ~n27178 ;
  assign n27180 = ~\pi0947  & ~n6761 ;
  assign n27181 = ~\pi0947  & n21658 ;
  assign n27182 = ~n21684 & n27181 ;
  assign n27183 = ~n27180 & ~n27182 ;
  assign n27184 = n21651 & ~n27183 ;
  assign n27185 = ~n6761 & ~n26930 ;
  assign n27186 = n21658 & ~n26930 ;
  assign n27187 = ~n21684 & n27186 ;
  assign n27188 = ~n27185 & ~n27187 ;
  assign n27189 = \pi0223  & n21651 ;
  assign n27190 = ~n27188 & n27189 ;
  assign n27191 = n27184 & n27190 ;
  assign n27192 = ~\pi0299  & n27191 ;
  assign n27193 = n1281 & n2165 ;
  assign n27194 = n1260 & n27193 ;
  assign n27195 = ~n21285 & n27194 ;
  assign n27196 = n21612 & ~n27195 ;
  assign n27197 = ~n21606 & n27196 ;
  assign n27198 = n2165 & ~n2280 ;
  assign n27199 = n2165 & ~n21282 ;
  assign n27200 = ~n21281 & n27199 ;
  assign n27201 = ~n27198 & ~n27200 ;
  assign n27202 = n6730 & n27201 ;
  assign n27203 = ~n27197 & n27202 ;
  assign n27204 = \pi0223  & ~n27184 ;
  assign n27205 = n21651 & ~n27188 ;
  assign n27206 = \pi0223  & ~n27205 ;
  assign n27207 = ~n27204 & ~n27206 ;
  assign n27208 = ~\pi0299  & n27207 ;
  assign n27209 = n27203 & n27208 ;
  assign n27210 = ~n27192 & ~n27209 ;
  assign n27211 = ~n27126 & n27129 ;
  assign n27212 = \pi0299  & ~\pi0947  ;
  assign n27213 = ~n27115 & n27212 ;
  assign n27214 = ~n27211 & n27213 ;
  assign n27215 = n27210 & ~n27214 ;
  assign n27216 = \pi0039  & ~n27215 ;
  assign n27217 = ~n21238 & n26957 ;
  assign n27218 = ~\pi0299  & ~n21740 ;
  assign n27219 = ~n21738 & n27218 ;
  assign n27220 = ~n27217 & ~n27219 ;
  assign n27221 = ~\pi0039  & ~\pi0947  ;
  assign n27222 = ~\pi0907  & n27221 ;
  assign n27223 = ~n27220 & n27222 ;
  assign n27224 = ~\pi0147  & ~n27223 ;
  assign n27225 = ~n27155 & n27224 ;
  assign n27226 = ~n27216 & n27225 ;
  assign n27227 = ~n27179 & ~n27226 ;
  assign n27228 = n27141 & n27227 ;
  assign n27229 = ~\pi0147  & ~n11834 ;
  assign n27230 = ~\pi0832  & ~n27229 ;
  assign n27231 = n27228 & n27230 ;
  assign n27232 = ~\pi0947  & n25039 ;
  assign n27233 = ~n21205 & n27212 ;
  assign n27234 = ~n21238 & n27233 ;
  assign n27235 = n1288 & n27234 ;
  assign n27236 = ~\pi0299  & ~\pi0947  ;
  assign n27237 = ~n21740 & n27236 ;
  assign n27238 = ~n21738 & n27237 ;
  assign n27239 = n1288 & n27238 ;
  assign n27240 = ~n27235 & ~n27239 ;
  assign n27241 = ~\pi0039  & ~n27234 ;
  assign n27242 = ~n27238 & n27241 ;
  assign n27243 = ~\pi0038  & ~n27242 ;
  assign n27244 = ~\pi0299  & \pi0947  ;
  assign n27245 = ~n21690 & n27244 ;
  assign n27246 = n21688 & n27245 ;
  assign n27247 = ~n21614 & n27246 ;
  assign n27248 = n27243 & ~n27247 ;
  assign n27249 = n27240 & ~n27248 ;
  assign n27250 = ~n2352 & ~n27077 ;
  assign n27251 = ~n21698 & ~n27250 ;
  assign n27252 = n21694 & ~n27250 ;
  assign n27253 = ~n21711 & n27252 ;
  assign n27254 = ~n27251 & ~n27253 ;
  assign n27255 = ~\pi0947  & n2352 ;
  assign n27256 = ~n21285 & n27255 ;
  assign n27257 = ~\pi0215  & ~n27256 ;
  assign n27258 = ~n27254 & n27257 ;
  assign n27259 = \pi0215  & ~n27082 ;
  assign n27260 = ~n21724 & n27259 ;
  assign n27261 = \pi0299  & ~n27260 ;
  assign n27262 = ~n27258 & n27261 ;
  assign n27263 = ~\pi0299  & ~n21690 ;
  assign n27264 = n21688 & n27263 ;
  assign n27265 = ~n21614 & n27264 ;
  assign n27266 = n27240 & ~n27265 ;
  assign n27267 = ~n27262 & n27266 ;
  assign n27268 = ~n27249 & ~n27267 ;
  assign n27269 = ~n27232 & ~n27268 ;
  assign n27270 = ~\pi0770  & ~n27269 ;
  assign n27271 = ~\pi0038  & \pi0770  ;
  assign n27272 = \pi0770  & n21765 ;
  assign n27273 = n1638 & n27272 ;
  assign n27274 = ~n27271 & ~n27273 ;
  assign n27275 = n11834 & n27274 ;
  assign n27276 = n11834 & n21770 ;
  assign n27277 = ~n21734 & n27276 ;
  assign n27278 = ~n27275 & ~n27277 ;
  assign n27279 = ~\pi0147  & ~n27278 ;
  assign n27280 = ~n27270 & n27279 ;
  assign n27281 = \pi0147  & ~\pi0770  ;
  assign n27282 = ~\pi0726  & ~n27281 ;
  assign n27283 = \pi0947  & n21688 ;
  assign n27284 = ~n21690 & n27283 ;
  assign n27285 = ~n21614 & n27284 ;
  assign n27286 = n6205 & ~n27285 ;
  assign n27287 = n7304 & ~n21205 ;
  assign n27288 = ~n21238 & n27287 ;
  assign n27289 = ~n21740 & n27244 ;
  assign n27290 = ~n21738 & n27289 ;
  assign n27291 = ~n27288 & ~n27290 ;
  assign n27292 = ~\pi0039  & n27291 ;
  assign n27293 = ~n22124 & ~n27232 ;
  assign n27294 = ~\pi0215  & \pi0947  ;
  assign n27295 = ~n21285 & n27294 ;
  assign n27296 = ~n24388 & ~n27295 ;
  assign n27297 = ~n27121 & ~n27296 ;
  assign n27298 = n21627 & n27111 ;
  assign n27299 = ~n21726 & n27298 ;
  assign n27300 = n2352 & n27294 ;
  assign n27301 = ~n21285 & n27300 ;
  assign n27302 = \pi0299  & ~n27301 ;
  assign n27303 = ~n27299 & n27302 ;
  assign n27304 = ~n27297 & n27303 ;
  assign n27305 = \pi0039  & n27304 ;
  assign n27306 = n27293 & ~n27305 ;
  assign n27307 = ~n27292 & n27306 ;
  assign n27308 = ~n27286 & n27307 ;
  assign n27309 = \pi0038  & n22123 ;
  assign n27310 = ~n27232 & n27309 ;
  assign n27311 = ~\pi0726  & ~n27310 ;
  assign n27312 = ~n27308 & n27311 ;
  assign n27313 = ~n27282 & ~n27312 ;
  assign n27314 = n11834 & n27313 ;
  assign n27315 = n27230 & ~n27314 ;
  assign n27316 = ~n27280 & n27315 ;
  assign n27317 = ~n27231 & ~n27316 ;
  assign n27318 = ~n27057 & n27317 ;
  assign n27319 = ~\pi0749  & \pi0947  ;
  assign n27320 = n27151 & ~n27319 ;
  assign n27321 = ~\pi0148  & ~n21757 ;
  assign n27322 = ~n27320 & ~n27321 ;
  assign n27323 = \pi0038  & ~n27322 ;
  assign n27324 = \pi0706  & ~n27323 ;
  assign n27325 = ~\pi0299  & n21740 ;
  assign n27326 = ~\pi0299  & n21737 ;
  assign n27327 = n21232 & n27326 ;
  assign n27328 = ~n27325 & ~n27327 ;
  assign n27329 = ~\pi0148  & ~n27328 ;
  assign n27330 = ~\pi0148  & \pi0299  ;
  assign n27331 = n21205 & n27330 ;
  assign n27332 = n21237 & n27330 ;
  assign n27333 = n21232 & n27332 ;
  assign n27334 = ~n27331 & ~n27333 ;
  assign n27335 = ~\pi0039  & n27334 ;
  assign n27336 = ~n27329 & n27335 ;
  assign n27337 = ~n27166 & ~n27319 ;
  assign n27338 = n27336 & ~n27337 ;
  assign n27339 = ~\pi0038  & ~n27338 ;
  assign n27340 = n27324 & ~n27339 ;
  assign n27341 = ~\pi0148  & n27215 ;
  assign n27342 = ~\pi0299  & ~n27158 ;
  assign n27343 = \pi0299  & ~n27172 ;
  assign n27344 = \pi0148  & ~n27343 ;
  assign n27345 = ~n27342 & n27344 ;
  assign n27346 = \pi0749  & ~n27345 ;
  assign n27347 = ~n27341 & n27346 ;
  assign n27348 = ~n27132 & ~n27136 ;
  assign n27349 = ~\pi0749  & ~n11168 ;
  assign n27350 = ~n27348 & n27349 ;
  assign n27351 = \pi0148  & ~n27084 ;
  assign n27352 = \pi0148  & ~\pi0299  ;
  assign n27353 = ~n21692 & n27352 ;
  assign n27354 = ~n27351 & ~n27353 ;
  assign n27355 = ~\pi0749  & ~n27354 ;
  assign n27356 = ~n27350 & ~n27355 ;
  assign n27357 = ~n27347 & n27356 ;
  assign n27358 = \pi0039  & n27324 ;
  assign n27359 = ~n27357 & n27358 ;
  assign n27360 = ~n27340 & ~n27359 ;
  assign n27361 = ~\pi0299  & ~n27285 ;
  assign n27362 = ~\pi0148  & ~n21692 ;
  assign n27363 = n27361 & ~n27362 ;
  assign n27364 = \pi0749  & ~n27363 ;
  assign n27365 = \pi0749  & \pi0947  ;
  assign n27366 = \pi0299  & n27365 ;
  assign n27367 = ~n21205 & n27366 ;
  assign n27368 = ~n21238 & n27367 ;
  assign n27369 = ~\pi0299  & n27365 ;
  assign n27370 = ~n21740 & n27369 ;
  assign n27371 = ~n21738 & n27370 ;
  assign n27372 = ~n27368 & ~n27371 ;
  assign n27373 = n27336 & n27372 ;
  assign n27374 = ~\pi0038  & ~n27373 ;
  assign n27375 = ~n27304 & ~n27330 ;
  assign n27376 = ~\pi0148  & n27260 ;
  assign n27377 = ~\pi0148  & n27257 ;
  assign n27378 = ~n27254 & n27377 ;
  assign n27379 = ~n27376 & ~n27378 ;
  assign n27380 = ~n27375 & n27379 ;
  assign n27381 = n27374 & ~n27380 ;
  assign n27382 = n27364 & n27381 ;
  assign n27383 = ~\pi0148  & ~\pi0749  ;
  assign n27384 = ~\pi0299  & n27383 ;
  assign n27385 = ~n21692 & n27384 ;
  assign n27386 = \pi0039  & ~n27383 ;
  assign n27387 = ~n21733 & ~n27386 ;
  assign n27388 = ~n27385 & ~n27387 ;
  assign n27389 = n27374 & ~n27388 ;
  assign n27390 = n1689 & ~n27365 ;
  assign n27391 = n6784 & n27390 ;
  assign n27392 = n1266 & n27391 ;
  assign n27393 = n1354 & n27392 ;
  assign n27394 = n1358 & n27393 ;
  assign n27395 = \pi0038  & ~n27394 ;
  assign n27396 = ~\pi0706  & ~n27395 ;
  assign n27397 = \pi0148  & ~\pi0706  ;
  assign n27398 = ~n22123 & n27397 ;
  assign n27399 = ~n27396 & ~n27398 ;
  assign n27400 = ~n27389 & ~n27399 ;
  assign n27401 = ~n27382 & n27400 ;
  assign n27402 = n6848 & n6861 ;
  assign n27403 = \pi0057  & \pi0148  ;
  assign n27404 = ~\pi0832  & ~n27403 ;
  assign n27405 = n27402 & n27404 ;
  assign n27406 = ~n27401 & n27405 ;
  assign n27407 = n27360 & n27406 ;
  assign n27408 = ~\pi0057  & n6848 ;
  assign n27409 = n6861 & n27408 ;
  assign n27410 = ~\pi0057  & \pi0148  ;
  assign n27411 = n27404 & ~n27410 ;
  assign n27412 = ~n27409 & n27411 ;
  assign n27413 = \pi0706  & n26930 ;
  assign n27414 = n27390 & ~n27413 ;
  assign n27415 = \pi0148  & ~n1689 ;
  assign n27416 = \pi0832  & ~n27415 ;
  assign n27417 = ~n27414 & n27416 ;
  assign n27418 = ~n27412 & ~n27417 ;
  assign n27419 = ~n27407 & n27418 ;
  assign n27420 = ~\pi0149  & ~n11834 ;
  assign n27421 = ~\pi0832  & ~n27420 ;
  assign n27422 = ~\pi0755  & \pi0947  ;
  assign n27423 = ~\pi0725  & n26930 ;
  assign n27424 = ~n27422 & ~n27423 ;
  assign n27425 = n1689 & ~n27424 ;
  assign n27426 = ~\pi0149  & ~n1689 ;
  assign n27427 = \pi0832  & ~n27426 ;
  assign n27428 = ~n27425 & n27427 ;
  assign n27429 = ~n27421 & ~n27428 ;
  assign n27430 = n6784 & ~n27422 ;
  assign n27431 = n1266 & n27430 ;
  assign n27432 = n22706 & n27431 ;
  assign n27433 = n1358 & n27432 ;
  assign n27434 = ~n26930 & n27433 ;
  assign n27435 = \pi0149  & ~n21757 ;
  assign n27436 = \pi0038  & ~n27435 ;
  assign n27437 = ~n27434 & n27436 ;
  assign n27438 = ~\pi0725  & ~n27437 ;
  assign n27439 = ~\pi0149  & ~n27328 ;
  assign n27440 = n20009 & n21205 ;
  assign n27441 = n20009 & n21237 ;
  assign n27442 = n21232 & n27441 ;
  assign n27443 = ~n27440 & ~n27442 ;
  assign n27444 = ~\pi0039  & n27443 ;
  assign n27445 = ~n27439 & n27444 ;
  assign n27446 = \pi0299  & n27422 ;
  assign n27447 = ~n21205 & n27446 ;
  assign n27448 = ~n21238 & n27447 ;
  assign n27449 = ~\pi0299  & n27422 ;
  assign n27450 = ~n21740 & n27449 ;
  assign n27451 = ~n21738 & n27450 ;
  assign n27452 = ~n27448 & ~n27451 ;
  assign n27453 = n27068 & n27452 ;
  assign n27454 = n27445 & n27453 ;
  assign n27455 = ~\pi0038  & ~n27454 ;
  assign n27456 = n27438 & ~n27455 ;
  assign n27457 = ~\pi0149  & n27132 ;
  assign n27458 = \pi0149  & ~n27084 ;
  assign n27459 = \pi0149  & ~\pi0299  ;
  assign n27460 = ~n21692 & n27459 ;
  assign n27461 = ~n27458 & ~n27460 ;
  assign n27462 = ~n27136 & n27461 ;
  assign n27463 = ~n27457 & n27462 ;
  assign n27464 = \pi0755  & ~n27463 ;
  assign n27465 = ~\pi0149  & n27215 ;
  assign n27466 = \pi0149  & ~n27343 ;
  assign n27467 = ~\pi0755  & ~n27466 ;
  assign n27468 = ~\pi0299  & ~\pi0755  ;
  assign n27469 = ~n27158 & n27468 ;
  assign n27470 = ~n27467 & ~n27469 ;
  assign n27471 = ~n27465 & ~n27470 ;
  assign n27472 = ~n27464 & ~n27471 ;
  assign n27473 = \pi0039  & n27438 ;
  assign n27474 = ~n27472 & n27473 ;
  assign n27475 = ~n27456 & ~n27474 ;
  assign n27476 = n27445 & n27452 ;
  assign n27477 = ~\pi0038  & ~n27476 ;
  assign n27478 = \pi0038  & ~n27433 ;
  assign n27479 = \pi0725  & ~n27478 ;
  assign n27480 = \pi0149  & \pi0725  ;
  assign n27481 = ~n22123 & n27480 ;
  assign n27482 = ~n27479 & ~n27481 ;
  assign n27483 = ~n27477 & ~n27482 ;
  assign n27484 = ~\pi0149  & ~n21692 ;
  assign n27485 = n27361 & ~n27484 ;
  assign n27486 = ~\pi0755  & ~n27485 ;
  assign n27487 = ~n20009 & ~n27304 ;
  assign n27488 = ~\pi0149  & n27260 ;
  assign n27489 = ~\pi0149  & n27257 ;
  assign n27490 = ~n27254 & n27489 ;
  assign n27491 = ~n27488 & ~n27490 ;
  assign n27492 = ~n27487 & n27491 ;
  assign n27493 = n27486 & ~n27492 ;
  assign n27494 = ~\pi0149  & \pi0755  ;
  assign n27495 = ~\pi0299  & n27494 ;
  assign n27496 = ~n21692 & n27495 ;
  assign n27497 = \pi0039  & ~n27494 ;
  assign n27498 = ~n21733 & ~n27497 ;
  assign n27499 = ~n27496 & ~n27498 ;
  assign n27500 = ~n27482 & n27499 ;
  assign n27501 = ~n27493 & n27500 ;
  assign n27502 = ~n27483 & ~n27501 ;
  assign n27503 = n11834 & ~n27428 ;
  assign n27504 = n27502 & n27503 ;
  assign n27505 = n27475 & n27504 ;
  assign n27506 = ~n27429 & ~n27505 ;
  assign n27507 = ~\pi0751  & \pi0947  ;
  assign n27508 = ~\pi0701  & n26930 ;
  assign n27509 = ~n27507 & ~n27508 ;
  assign n27510 = n1689 & ~n27509 ;
  assign n27511 = ~\pi0150  & ~n1689 ;
  assign n27512 = \pi0832  & ~n27511 ;
  assign n27513 = ~n27510 & n27512 ;
  assign n27514 = ~\pi0150  & n27215 ;
  assign n27515 = \pi0150  & ~n27343 ;
  assign n27516 = ~\pi0751  & ~n27515 ;
  assign n27517 = ~\pi0299  & ~\pi0751  ;
  assign n27518 = ~n27158 & n27517 ;
  assign n27519 = ~n27516 & ~n27518 ;
  assign n27520 = ~n27514 & ~n27519 ;
  assign n27521 = ~\pi0150  & ~n27136 ;
  assign n27522 = ~n27132 & n27521 ;
  assign n27523 = ~\pi0299  & ~n27060 ;
  assign n27524 = \pi0150  & ~n27083 ;
  assign n27525 = n27080 & n27524 ;
  assign n27526 = ~n27523 & n27525 ;
  assign n27527 = \pi0751  & ~n27526 ;
  assign n27528 = ~n27522 & n27527 ;
  assign n27529 = \pi0039  & ~n27528 ;
  assign n27530 = ~n27520 & n27529 ;
  assign n27531 = ~n27106 & ~n27507 ;
  assign n27532 = \pi0150  & ~n27219 ;
  assign n27533 = ~n27217 & n27532 ;
  assign n27534 = ~\pi0039  & ~n27533 ;
  assign n27535 = ~n27531 & n27534 ;
  assign n27536 = ~\pi0038  & ~n27535 ;
  assign n27537 = ~n27530 & n27536 ;
  assign n27538 = \pi0150  & ~n21757 ;
  assign n27539 = n6784 & ~n27507 ;
  assign n27540 = n1266 & n27539 ;
  assign n27541 = n22706 & n27540 ;
  assign n27542 = n1358 & n27541 ;
  assign n27543 = ~n26930 & n27542 ;
  assign n27544 = ~n27538 & ~n27543 ;
  assign n27545 = \pi0038  & ~n27544 ;
  assign n27546 = ~\pi0701  & n11834 ;
  assign n27547 = ~n27545 & n27546 ;
  assign n27548 = ~n27537 & n27547 ;
  assign n27549 = ~n27262 & ~n27265 ;
  assign n27550 = ~\pi0150  & ~n27247 ;
  assign n27551 = ~n27549 & n27550 ;
  assign n27552 = \pi0150  & ~\pi0299  ;
  assign n27553 = ~n27285 & n27552 ;
  assign n27554 = \pi0150  & n27304 ;
  assign n27555 = ~\pi0751  & ~n27554 ;
  assign n27556 = ~n27553 & n27555 ;
  assign n27557 = ~n27551 & n27556 ;
  assign n27558 = \pi0299  & \pi0751  ;
  assign n27559 = ~n21205 & n27558 ;
  assign n27560 = ~n21238 & n27559 ;
  assign n27561 = ~\pi0299  & \pi0751  ;
  assign n27562 = ~n21740 & n27561 ;
  assign n27563 = ~n21738 & n27562 ;
  assign n27564 = ~n27560 & ~n27563 ;
  assign n27565 = ~n27533 & n27564 ;
  assign n27566 = n27242 & n27565 ;
  assign n27567 = ~\pi0038  & ~n27566 ;
  assign n27568 = ~\pi0150  & \pi0751  ;
  assign n27569 = ~\pi0299  & n27568 ;
  assign n27570 = ~n21692 & n27569 ;
  assign n27571 = ~n25541 & n27568 ;
  assign n27572 = ~n27570 & ~n27571 ;
  assign n27573 = n27567 & n27572 ;
  assign n27574 = ~n27557 & n27573 ;
  assign n27575 = n1288 & ~n27566 ;
  assign n27576 = \pi0038  & \pi0150  ;
  assign n27577 = ~n22123 & n27576 ;
  assign n27578 = \pi0038  & n27542 ;
  assign n27579 = \pi0701  & ~n27578 ;
  assign n27580 = ~n27577 & n27579 ;
  assign n27581 = ~n27575 & n27580 ;
  assign n27582 = n11834 & n27581 ;
  assign n27583 = ~n27574 & n27582 ;
  assign n27584 = ~\pi0150  & ~n11834 ;
  assign n27585 = ~\pi0832  & ~n27584 ;
  assign n27586 = ~n27583 & n27585 ;
  assign n27587 = ~n27548 & n27586 ;
  assign n27588 = ~n27513 & ~n27587 ;
  assign n27589 = ~\pi0745  & \pi0947  ;
  assign n27590 = ~\pi0723  & n26930 ;
  assign n27591 = ~n27589 & ~n27590 ;
  assign n27592 = n1689 & ~n27591 ;
  assign n27593 = ~\pi0151  & ~n1689 ;
  assign n27594 = \pi0832  & ~n27593 ;
  assign n27595 = ~n27592 & n27594 ;
  assign n27596 = ~\pi0039  & ~\pi0745  ;
  assign n27597 = ~n27291 & n27596 ;
  assign n27598 = ~\pi0151  & ~n27219 ;
  assign n27599 = ~\pi0039  & ~n27217 ;
  assign n27600 = n27598 & n27599 ;
  assign n27601 = ~\pi0038  & ~n27600 ;
  assign n27602 = ~n27597 & n27601 ;
  assign n27603 = \pi0038  & \pi0151  ;
  assign n27604 = ~n22123 & n27603 ;
  assign n27605 = n6784 & ~n27589 ;
  assign n27606 = n1266 & n27605 ;
  assign n27607 = n22706 & n27606 ;
  assign n27608 = n1358 & n27607 ;
  assign n27609 = \pi0038  & n27608 ;
  assign n27610 = \pi0723  & ~n27609 ;
  assign n27611 = ~n27604 & n27610 ;
  assign n27612 = ~n27602 & n27611 ;
  assign n27613 = n11834 & n27612 ;
  assign n27614 = ~\pi0745  & ~n21693 ;
  assign n27615 = ~\pi0151  & ~n25541 ;
  assign n27616 = ~\pi0151  & ~\pi0299  ;
  assign n27617 = ~n21692 & n27616 ;
  assign n27618 = ~n27615 & ~n27617 ;
  assign n27619 = ~n27614 & ~n27618 ;
  assign n27620 = ~\pi0215  & ~n27254 ;
  assign n27621 = \pi0151  & n2352 ;
  assign n27622 = n21285 & n27621 ;
  assign n27623 = ~n27256 & ~n27622 ;
  assign n27624 = ~n6730 & ~n21334 ;
  assign n27625 = n6713 & ~n6730 ;
  assign n27626 = ~n21329 & n27625 ;
  assign n27627 = ~n27624 & ~n27626 ;
  assign n27628 = \pi0151  & ~n2352 ;
  assign n27629 = n27627 & n27628 ;
  assign n27630 = ~n21698 & ~n27629 ;
  assign n27631 = n21694 & ~n27629 ;
  assign n27632 = ~n21711 & n27631 ;
  assign n27633 = ~n27630 & ~n27632 ;
  assign n27634 = n27623 & ~n27633 ;
  assign n27635 = n27620 & n27634 ;
  assign n27636 = \pi0299  & ~n27259 ;
  assign n27637 = ~\pi0151  & ~n27082 ;
  assign n27638 = ~n21724 & n27637 ;
  assign n27639 = \pi0299  & ~n21728 ;
  assign n27640 = ~n27638 & n27639 ;
  assign n27641 = ~n27636 & ~n27640 ;
  assign n27642 = ~n27635 & ~n27641 ;
  assign n27643 = ~\pi0745  & ~n27361 ;
  assign n27644 = ~n27642 & n27643 ;
  assign n27645 = ~n27619 & ~n27644 ;
  assign n27646 = \pi0039  & \pi0723  ;
  assign n27647 = ~n27609 & n27646 ;
  assign n27648 = ~n27604 & n27647 ;
  assign n27649 = n11834 & n27648 ;
  assign n27650 = ~n27645 & n27649 ;
  assign n27651 = ~n27613 & ~n27650 ;
  assign n27652 = ~\pi0151  & ~n21692 ;
  assign n27653 = ~\pi0299  & \pi0745  ;
  assign n27654 = ~n27060 & n27653 ;
  assign n27655 = ~n27652 & n27654 ;
  assign n27656 = ~\pi0215  & ~n27126 ;
  assign n27657 = ~n27128 & ~n27622 ;
  assign n27658 = ~n27299 & n27657 ;
  assign n27659 = ~n27633 & n27658 ;
  assign n27660 = n27656 & n27659 ;
  assign n27661 = \pi0215  & n21728 ;
  assign n27662 = \pi0215  & n27637 ;
  assign n27663 = ~n21724 & n27662 ;
  assign n27664 = ~n27661 & ~n27663 ;
  assign n27665 = ~n27299 & ~n27664 ;
  assign n27666 = \pi0299  & \pi0745  ;
  assign n27667 = ~n27665 & n27666 ;
  assign n27668 = ~n27660 & n27667 ;
  assign n27669 = ~n27655 & ~n27668 ;
  assign n27670 = n27203 & n27207 ;
  assign n27671 = ~\pi0299  & ~n27191 ;
  assign n27672 = ~n27670 & n27671 ;
  assign n27673 = \pi0151  & ~n27158 ;
  assign n27674 = n27672 & ~n27673 ;
  assign n27675 = \pi0299  & ~n27664 ;
  assign n27676 = ~n6730 & ~n21285 ;
  assign n27677 = ~n27657 & ~n27676 ;
  assign n27678 = ~\pi0215  & ~n27677 ;
  assign n27679 = \pi0299  & n27678 ;
  assign n27680 = ~n27633 & n27679 ;
  assign n27681 = ~n27675 & ~n27680 ;
  assign n27682 = ~\pi0745  & n27681 ;
  assign n27683 = ~n27674 & n27682 ;
  assign n27684 = n27669 & ~n27683 ;
  assign n27685 = n9627 & ~n27684 ;
  assign n27686 = ~n27217 & n27598 ;
  assign n27687 = ~\pi0745  & ~n27291 ;
  assign n27688 = ~n27686 & ~n27687 ;
  assign n27689 = ~\pi0038  & n27069 ;
  assign n27690 = n27688 & n27689 ;
  assign n27691 = \pi0151  & ~n21757 ;
  assign n27692 = ~n26930 & n27608 ;
  assign n27693 = ~n27691 & ~n27692 ;
  assign n27694 = \pi0038  & ~n27693 ;
  assign n27695 = ~\pi0723  & n11834 ;
  assign n27696 = ~n27694 & n27695 ;
  assign n27697 = ~n27690 & n27696 ;
  assign n27698 = ~n27685 & n27697 ;
  assign n27699 = n27651 & ~n27698 ;
  assign n27700 = ~\pi0151  & ~n11834 ;
  assign n27701 = ~\pi0832  & ~n27700 ;
  assign n27702 = n27699 & n27701 ;
  assign n27703 = ~n27595 & ~n27702 ;
  assign n27704 = ~\pi0152  & ~n11834 ;
  assign n27705 = ~\pi0832  & ~n27704 ;
  assign n27706 = \pi0759  & \pi0947  ;
  assign n27707 = n1689 & ~n27706 ;
  assign n27708 = \pi0696  & n26930 ;
  assign n27709 = n27707 & ~n27708 ;
  assign n27710 = ~\pi0152  & ~n1689 ;
  assign n27711 = \pi0832  & ~n27710 ;
  assign n27712 = ~n27709 & n27711 ;
  assign n27713 = ~n27705 & ~n27712 ;
  assign n27714 = \pi0152  & ~\pi0759  ;
  assign n27715 = ~n25542 & n27714 ;
  assign n27716 = \pi0039  & ~n27715 ;
  assign n27717 = \pi0759  & ~n27291 ;
  assign n27718 = \pi0152  & ~n27328 ;
  assign n27719 = \pi0152  & \pi0299  ;
  assign n27720 = n21205 & n27719 ;
  assign n27721 = n21237 & n27719 ;
  assign n27722 = n21232 & n27721 ;
  assign n27723 = ~n27720 & ~n27722 ;
  assign n27724 = ~\pi0039  & n27723 ;
  assign n27725 = ~n27718 & n27724 ;
  assign n27726 = ~n27717 & n27725 ;
  assign n27727 = ~\pi0038  & ~n27726 ;
  assign n27728 = ~n27716 & n27727 ;
  assign n27729 = n27121 & n27254 ;
  assign n27730 = n6730 & ~n21696 ;
  assign n27731 = \pi0152  & n27121 ;
  assign n27732 = ~n27730 & n27731 ;
  assign n27733 = n21694 & n27731 ;
  assign n27734 = ~n21711 & n27733 ;
  assign n27735 = ~n27732 & ~n27734 ;
  assign n27736 = ~n2352 & n27077 ;
  assign n27737 = n27121 & n27736 ;
  assign n27738 = n27735 & n27737 ;
  assign n27739 = ~n27729 & ~n27738 ;
  assign n27740 = ~\pi0152  & n2352 ;
  assign n27741 = n21285 & n27740 ;
  assign n27742 = n27257 & ~n27741 ;
  assign n27743 = n27739 & n27742 ;
  assign n27744 = \pi0152  & ~n27082 ;
  assign n27745 = \pi0215  & n27744 ;
  assign n27746 = ~n21724 & n27745 ;
  assign n27747 = \pi0299  & ~n27299 ;
  assign n27748 = ~n27746 & n27747 ;
  assign n27749 = ~n27743 & n27748 ;
  assign n27750 = ~n2165 & n21612 ;
  assign n27751 = ~n21606 & n27750 ;
  assign n27752 = \pi0947  & ~n2165 ;
  assign n27753 = ~n27751 & ~n27752 ;
  assign n27754 = ~\pi0152  & n21612 ;
  assign n27755 = ~n21606 & n27754 ;
  assign n27756 = ~\pi0223  & ~n27755 ;
  assign n27757 = ~n27753 & n27756 ;
  assign n27758 = ~\pi0152  & ~n21651 ;
  assign n27759 = ~\pi0152  & n6761 ;
  assign n27760 = ~n21685 & n27759 ;
  assign n27761 = ~n27758 & ~n27760 ;
  assign n27762 = n27204 & n27761 ;
  assign n27763 = \pi0152  & ~\pi0224  ;
  assign n27764 = ~\pi0222  & n27763 ;
  assign n27765 = n21285 & n27764 ;
  assign n27766 = \pi0947  & n2165 ;
  assign n27767 = ~n21285 & n27766 ;
  assign n27768 = ~n27765 & ~n27767 ;
  assign n27769 = ~\pi0223  & ~n27768 ;
  assign n27770 = ~\pi0299  & ~n27769 ;
  assign n27771 = ~n27762 & n27770 ;
  assign n27772 = ~n27757 & n27771 ;
  assign n27773 = \pi0759  & ~n27772 ;
  assign n27774 = n27727 & n27773 ;
  assign n27775 = ~n27749 & n27774 ;
  assign n27776 = ~n27728 & ~n27775 ;
  assign n27777 = n1354 & ~n27706 ;
  assign n27778 = n21755 & n27777 ;
  assign n27779 = n1358 & n27778 ;
  assign n27780 = \pi0038  & ~n27779 ;
  assign n27781 = ~\pi0696  & ~n27780 ;
  assign n27782 = ~\pi0152  & ~\pi0696  ;
  assign n27783 = ~n22123 & n27782 ;
  assign n27784 = ~n27781 & ~n27783 ;
  assign n27785 = n27776 & ~n27784 ;
  assign n27786 = n11834 & ~n27712 ;
  assign n27787 = n27785 & n27786 ;
  assign n27788 = n27068 & n27726 ;
  assign n27789 = ~\pi0038  & ~n27788 ;
  assign n27790 = ~n26930 & n27779 ;
  assign n27791 = ~\pi0152  & ~n21757 ;
  assign n27792 = \pi0038  & ~n27791 ;
  assign n27793 = ~n27790 & n27792 ;
  assign n27794 = ~n27789 & ~n27793 ;
  assign n27795 = ~\pi0299  & ~n27762 ;
  assign n27796 = n2165 & n6730 ;
  assign n27797 = ~\pi0223  & ~n27796 ;
  assign n27798 = ~n21285 & n27797 ;
  assign n27799 = ~\pi0152  & n2165 ;
  assign n27800 = ~\pi0223  & ~n27799 ;
  assign n27801 = n21285 & n27800 ;
  assign n27802 = ~n27798 & ~n27801 ;
  assign n27803 = ~n27755 & ~n27802 ;
  assign n27804 = ~n27753 & n27803 ;
  assign n27805 = ~n2165 & n6730 ;
  assign n27806 = ~n27802 & ~n27805 ;
  assign n27807 = ~n27751 & n27806 ;
  assign n27808 = n27206 & n27761 ;
  assign n27809 = ~n27807 & ~n27808 ;
  assign n27810 = ~n27804 & n27809 ;
  assign n27811 = n27795 & n27810 ;
  assign n27812 = ~\pi0907  & n27255 ;
  assign n27813 = ~n21285 & n27812 ;
  assign n27814 = ~n27741 & ~n27813 ;
  assign n27815 = ~\pi0215  & n27814 ;
  assign n27816 = ~\pi0152  & ~n21728 ;
  assign n27817 = \pi0215  & ~n27816 ;
  assign n27818 = ~n21724 & n27817 ;
  assign n27819 = \pi0299  & ~n27818 ;
  assign n27820 = ~n27815 & n27819 ;
  assign n27821 = n27627 & n27736 ;
  assign n27822 = n27819 & n27821 ;
  assign n27823 = n27735 & n27822 ;
  assign n27824 = ~n27820 & ~n27823 ;
  assign n27825 = \pi0759  & n27824 ;
  assign n27826 = ~n27811 & n27825 ;
  assign n27827 = ~n2165 & n26930 ;
  assign n27828 = ~n27751 & ~n27827 ;
  assign n27829 = n27756 & ~n27828 ;
  assign n27830 = n2165 & n26930 ;
  assign n27831 = ~n21285 & n27830 ;
  assign n27832 = \pi0152  & n2165 ;
  assign n27833 = n21285 & n27832 ;
  assign n27834 = ~n27831 & ~n27833 ;
  assign n27835 = ~\pi0223  & ~n27834 ;
  assign n27836 = ~\pi0299  & ~n27808 ;
  assign n27837 = ~n27835 & n27836 ;
  assign n27838 = ~n27829 & n27837 ;
  assign n27839 = ~\pi0299  & ~\pi0759  ;
  assign n27840 = ~\pi0215  & ~n26930 ;
  assign n27841 = n21727 & ~n26930 ;
  assign n27842 = ~n21726 & n27841 ;
  assign n27843 = ~n27840 & ~n27842 ;
  assign n27844 = ~\pi0759  & n27843 ;
  assign n27845 = n27818 & n27844 ;
  assign n27846 = ~n27839 & ~n27845 ;
  assign n27847 = n27735 & n27736 ;
  assign n27848 = ~\pi0215  & ~\pi0759  ;
  assign n27849 = ~n27128 & n27848 ;
  assign n27850 = n27814 & n27849 ;
  assign n27851 = ~n27847 & n27850 ;
  assign n27852 = n27846 & ~n27851 ;
  assign n27853 = ~n27838 & ~n27852 ;
  assign n27854 = ~n27826 & ~n27853 ;
  assign n27855 = \pi0039  & ~n27793 ;
  assign n27856 = n27854 & n27855 ;
  assign n27857 = ~n27794 & ~n27856 ;
  assign n27858 = \pi0696  & n27786 ;
  assign n27859 = ~n27857 & n27858 ;
  assign n27860 = ~n27787 & ~n27859 ;
  assign n27861 = ~n27713 & n27860 ;
  assign n27862 = \pi0700  & n26930 ;
  assign n27863 = \pi0766  & \pi0947  ;
  assign n27864 = n1689 & ~n27863 ;
  assign n27865 = ~n27862 & n27864 ;
  assign n27866 = \pi0153  & ~n1689 ;
  assign n27867 = \pi0832  & ~n27866 ;
  assign n27868 = ~n27865 & n27867 ;
  assign n27869 = \pi0057  & \pi0153  ;
  assign n27870 = ~\pi0832  & ~n27869 ;
  assign n27871 = ~\pi0057  & \pi0153  ;
  assign n27872 = ~n27409 & ~n27871 ;
  assign n27873 = \pi0153  & ~\pi0700  ;
  assign n27874 = ~n22123 & n27873 ;
  assign n27875 = \pi0700  & n27402 ;
  assign n27876 = n1354 & ~n27863 ;
  assign n27877 = n21755 & n27876 ;
  assign n27878 = n1358 & n27877 ;
  assign n27879 = \pi0038  & n27402 ;
  assign n27880 = ~n27878 & n27879 ;
  assign n27881 = ~n27875 & ~n27880 ;
  assign n27882 = ~n27874 & ~n27881 ;
  assign n27883 = ~\pi0153  & ~n21692 ;
  assign n27884 = n27361 & ~n27883 ;
  assign n27885 = \pi0153  & ~n21728 ;
  assign n27886 = n27259 & ~n27885 ;
  assign n27887 = ~n21724 & n27886 ;
  assign n27888 = \pi0299  & ~n27887 ;
  assign n27889 = \pi0766  & ~n27888 ;
  assign n27890 = n21694 & ~n21711 ;
  assign n27891 = n21698 & ~n27890 ;
  assign n27892 = \pi0153  & ~n2352 ;
  assign n27893 = n27627 & n27892 ;
  assign n27894 = \pi0153  & n2352 ;
  assign n27895 = n21285 & n27894 ;
  assign n27896 = ~n27256 & ~n27895 ;
  assign n27897 = \pi0766  & n27896 ;
  assign n27898 = ~n27893 & n27897 ;
  assign n27899 = ~\pi0215  & ~n27250 ;
  assign n27900 = n27898 & n27899 ;
  assign n27901 = ~n27891 & n27900 ;
  assign n27902 = ~n27889 & ~n27901 ;
  assign n27903 = ~n27884 & ~n27902 ;
  assign n27904 = ~\pi0153  & ~\pi0766  ;
  assign n27905 = ~\pi0299  & n27904 ;
  assign n27906 = ~n21692 & n27905 ;
  assign n27907 = \pi0039  & ~n27904 ;
  assign n27908 = ~n21733 & ~n27907 ;
  assign n27909 = ~n27906 & ~n27908 ;
  assign n27910 = ~n27903 & n27909 ;
  assign n27911 = ~\pi0766  & ~n21743 ;
  assign n27912 = ~n27292 & ~n27911 ;
  assign n27913 = ~\pi0153  & ~n27219 ;
  assign n27914 = ~n27217 & n27913 ;
  assign n27915 = ~n27912 & ~n27914 ;
  assign n27916 = ~\pi0038  & n27402 ;
  assign n27917 = ~n27915 & n27916 ;
  assign n27918 = ~n27910 & n27917 ;
  assign n27919 = ~n27882 & ~n27918 ;
  assign n27920 = ~n27872 & n27919 ;
  assign n27921 = n27068 & ~n27914 ;
  assign n27922 = ~n27912 & n27921 ;
  assign n27923 = ~\pi0038  & ~n27922 ;
  assign n27924 = \pi0153  & ~n27158 ;
  assign n27925 = n27672 & ~n27924 ;
  assign n27926 = ~\pi0299  & \pi0766  ;
  assign n27927 = ~n27813 & ~n27895 ;
  assign n27928 = ~\pi0215  & n27927 ;
  assign n27929 = ~n27893 & n27928 ;
  assign n27930 = ~n21698 & n27929 ;
  assign n27931 = n21694 & n27929 ;
  assign n27932 = ~n21711 & n27931 ;
  assign n27933 = ~n27930 & ~n27932 ;
  assign n27934 = \pi0215  & ~n27885 ;
  assign n27935 = ~n21724 & n27934 ;
  assign n27936 = \pi0766  & ~n27935 ;
  assign n27937 = n27933 & n27936 ;
  assign n27938 = ~n27926 & ~n27937 ;
  assign n27939 = ~n27925 & ~n27938 ;
  assign n27940 = \pi0039  & n27939 ;
  assign n27941 = ~n27128 & ~n27895 ;
  assign n27942 = ~n27893 & n27941 ;
  assign n27943 = ~n27122 & n27942 ;
  assign n27944 = ~n27891 & n27943 ;
  assign n27945 = n21948 & ~n27944 ;
  assign n27946 = n27523 & ~n27883 ;
  assign n27947 = n21724 & n21729 ;
  assign n27948 = \pi0153  & \pi0215  ;
  assign n27949 = ~n21728 & n27948 ;
  assign n27950 = ~n27299 & ~n27949 ;
  assign n27951 = ~n27947 & n27950 ;
  assign n27952 = \pi0299  & ~n27951 ;
  assign n27953 = ~n27946 & ~n27952 ;
  assign n27954 = ~n27945 & n27953 ;
  assign n27955 = \pi0039  & ~\pi0766  ;
  assign n27956 = ~n27954 & n27955 ;
  assign n27957 = ~n27940 & ~n27956 ;
  assign n27958 = n27923 & n27957 ;
  assign n27959 = ~n26930 & n27878 ;
  assign n27960 = \pi0153  & ~n21757 ;
  assign n27961 = \pi0038  & ~n27960 ;
  assign n27962 = ~n27959 & n27961 ;
  assign n27963 = \pi0700  & ~n27962 ;
  assign n27964 = ~n27872 & n27963 ;
  assign n27965 = ~n27958 & n27964 ;
  assign n27966 = ~n27920 & ~n27965 ;
  assign n27967 = n27870 & n27966 ;
  assign n27968 = ~n27868 & ~n27967 ;
  assign n27969 = ~\pi0742  & \pi0947  ;
  assign n27970 = ~\pi0704  & n26930 ;
  assign n27971 = ~n27969 & ~n27970 ;
  assign n27972 = n1689 & ~n27971 ;
  assign n27973 = ~\pi0154  & ~n1689 ;
  assign n27974 = \pi0832  & ~n27973 ;
  assign n27975 = ~n27972 & n27974 ;
  assign n27976 = ~\pi0154  & ~n27219 ;
  assign n27977 = ~n27217 & n27976 ;
  assign n27978 = n27069 & ~n27977 ;
  assign n27979 = n27166 & n27978 ;
  assign n27980 = ~\pi0154  & ~n27979 ;
  assign n27981 = n27215 & n27980 ;
  assign n27982 = \pi0039  & ~\pi0299  ;
  assign n27983 = ~n27158 & n27982 ;
  assign n27984 = \pi0154  & ~n27343 ;
  assign n27985 = \pi0039  & ~n27984 ;
  assign n27986 = ~n27983 & ~n27985 ;
  assign n27987 = ~n27979 & n27986 ;
  assign n27988 = ~\pi0038  & ~n27987 ;
  assign n27989 = ~n27981 & n27988 ;
  assign n27990 = \pi0038  & ~n27151 ;
  assign n27991 = ~\pi0154  & ~n21757 ;
  assign n27992 = n27990 & ~n27991 ;
  assign n27993 = ~\pi0742  & ~n27992 ;
  assign n27994 = ~n27989 & n27993 ;
  assign n27995 = ~\pi0154  & ~n27136 ;
  assign n27996 = ~n27132 & n27995 ;
  assign n27997 = ~n27060 & n27982 ;
  assign n27998 = \pi0154  & ~n27083 ;
  assign n27999 = n27080 & n27998 ;
  assign n28000 = \pi0039  & ~n27999 ;
  assign n28001 = ~n27997 & ~n28000 ;
  assign n28002 = ~n27996 & ~n28001 ;
  assign n28003 = n27096 & ~n27991 ;
  assign n28004 = \pi0742  & ~n28003 ;
  assign n28005 = ~n27978 & n28004 ;
  assign n28006 = ~n28002 & n28005 ;
  assign n28007 = \pi0038  & \pi0742  ;
  assign n28008 = ~n28003 & n28007 ;
  assign n28009 = ~\pi0704  & ~n28008 ;
  assign n28010 = ~n28006 & n28009 ;
  assign n28011 = ~n27994 & n28010 ;
  assign n28012 = ~\pi0154  & \pi0742  ;
  assign n28013 = n21770 & n28012 ;
  assign n28014 = ~n21734 & n28013 ;
  assign n28015 = \pi0038  & n28012 ;
  assign n28016 = ~n22123 & n28015 ;
  assign n28017 = \pi0704  & ~n28016 ;
  assign n28018 = ~n28014 & n28017 ;
  assign n28019 = n11834 & ~n28018 ;
  assign n28020 = n27292 & ~n27977 ;
  assign n28021 = ~\pi0038  & n28020 ;
  assign n28022 = \pi0154  & ~n27304 ;
  assign n28023 = ~n27361 & n28022 ;
  assign n28024 = n9627 & ~n28023 ;
  assign n28025 = ~n28021 & ~n28024 ;
  assign n28026 = \pi0038  & \pi0154  ;
  assign n28027 = ~\pi0742  & ~n28026 ;
  assign n28028 = ~\pi0742  & n21765 ;
  assign n28029 = n1638 & n28028 ;
  assign n28030 = ~n28027 & ~n28029 ;
  assign n28031 = \pi0038  & ~\pi0947  ;
  assign n28032 = n21765 & n28031 ;
  assign n28033 = n1638 & n28032 ;
  assign n28034 = n11834 & ~n28033 ;
  assign n28035 = ~n28030 & n28034 ;
  assign n28036 = n28025 & n28035 ;
  assign n28037 = ~n27247 & ~n27549 ;
  assign n28038 = ~\pi0154  & ~n28020 ;
  assign n28039 = n28035 & n28038 ;
  assign n28040 = ~n28037 & n28039 ;
  assign n28041 = ~n28036 & ~n28040 ;
  assign n28042 = ~n28019 & n28041 ;
  assign n28043 = ~n28011 & ~n28042 ;
  assign n28044 = ~\pi0154  & ~n11834 ;
  assign n28045 = ~\pi0832  & ~n28044 ;
  assign n28046 = ~n28043 & n28045 ;
  assign n28047 = ~n27975 & ~n28046 ;
  assign n28048 = \pi0038  & n27151 ;
  assign n28049 = ~n27173 & ~n27990 ;
  assign n28050 = ~n27167 & n28049 ;
  assign n28051 = ~n27159 & n28050 ;
  assign n28052 = ~n28048 & ~n28051 ;
  assign n28053 = ~\pi0686  & ~\pi0757  ;
  assign n28054 = ~n28052 & n28053 ;
  assign n28055 = \pi0038  & n27093 ;
  assign n28056 = n26939 & n28055 ;
  assign n28057 = n10323 & n28056 ;
  assign n28058 = ~n27085 & ~n27096 ;
  assign n28059 = ~n27069 & n28058 ;
  assign n28060 = ~n27061 & n28059 ;
  assign n28061 = ~n28057 & ~n28060 ;
  assign n28062 = ~\pi0686  & \pi0757  ;
  assign n28063 = ~n28061 & n28062 ;
  assign n28064 = ~n28054 & ~n28063 ;
  assign n28065 = \pi0686  & ~\pi0757  ;
  assign n28066 = ~\pi0832  & ~n28065 ;
  assign n28067 = ~\pi0832  & ~n27310 ;
  assign n28068 = ~n27308 & n28067 ;
  assign n28069 = ~n28066 & ~n28068 ;
  assign n28070 = n28064 & ~n28069 ;
  assign n28071 = ~\pi0757  & \pi0947  ;
  assign n28072 = ~\pi0686  & n26930 ;
  assign n28073 = ~n28071 & ~n28072 ;
  assign n28074 = n1689 & ~n28073 ;
  assign n28075 = ~\pi0155  & ~n1689 ;
  assign n28076 = \pi0832  & ~n28075 ;
  assign n28077 = ~n28074 & n28076 ;
  assign n28078 = ~\pi0057  & \pi0155  ;
  assign n28079 = n6848 & n28078 ;
  assign n28080 = n6861 & n28079 ;
  assign n28081 = ~\pi0832  & ~n28080 ;
  assign n28082 = ~n28077 & ~n28081 ;
  assign n28083 = ~n28070 & n28082 ;
  assign n28084 = ~n21734 & n21770 ;
  assign n28085 = \pi0757  & ~n22124 ;
  assign n28086 = ~n28084 & n28085 ;
  assign n28087 = \pi0686  & ~n28086 ;
  assign n28088 = ~\pi0057  & n27402 ;
  assign n28089 = ~n28087 & n28088 ;
  assign n28090 = ~\pi0757  & n1289 ;
  assign n28091 = n1287 & n28090 ;
  assign n28092 = n9948 & n28091 ;
  assign n28093 = ~n27269 & n28092 ;
  assign n28094 = ~n28089 & ~n28093 ;
  assign n28095 = ~\pi0155  & ~n28076 ;
  assign n28096 = ~\pi0155  & n1689 ;
  assign n28097 = ~n28073 & n28096 ;
  assign n28098 = ~n28095 & ~n28097 ;
  assign n28099 = n28094 & ~n28098 ;
  assign n28100 = ~\pi0038  & n27223 ;
  assign n28101 = n9627 & ~n27215 ;
  assign n28102 = ~n28100 & ~n28101 ;
  assign n28103 = \pi0038  & n4520 ;
  assign n28104 = n27142 & n28103 ;
  assign n28105 = n1638 & n28104 ;
  assign n28106 = n28102 & ~n28105 ;
  assign n28107 = ~\pi0757  & ~n28106 ;
  assign n28108 = ~n27132 & n27137 ;
  assign n28109 = ~\pi0038  & \pi0757  ;
  assign n28110 = ~n27107 & n28109 ;
  assign n28111 = ~n28108 & n28110 ;
  assign n28112 = n12800 & ~n26930 ;
  assign n28113 = n1689 & n28112 ;
  assign n28114 = n1259 & n28113 ;
  assign n28115 = n1249 & n28114 ;
  assign n28116 = \pi0757  & n1281 ;
  assign n28117 = n28115 & n28116 ;
  assign n28118 = ~\pi0686  & ~n28117 ;
  assign n28119 = ~n28111 & n28118 ;
  assign n28120 = ~n28098 & n28119 ;
  assign n28121 = ~n28107 & n28120 ;
  assign n28122 = ~n28099 & ~n28121 ;
  assign n28123 = ~n28083 & n28122 ;
  assign n28124 = ~\pi0741  & \pi0947  ;
  assign n28125 = ~\pi0724  & n26930 ;
  assign n28126 = ~n28124 & ~n28125 ;
  assign n28127 = n1689 & ~n28126 ;
  assign n28128 = ~\pi0156  & ~n1689 ;
  assign n28129 = \pi0832  & ~n28128 ;
  assign n28130 = ~n28127 & n28129 ;
  assign n28131 = ~\pi0724  & \pi0741  ;
  assign n28132 = ~\pi0724  & ~n28105 ;
  assign n28133 = n28102 & n28132 ;
  assign n28134 = ~n28131 & ~n28133 ;
  assign n28135 = ~\pi0038  & \pi0741  ;
  assign n28136 = ~n27107 & n28135 ;
  assign n28137 = ~n28108 & n28136 ;
  assign n28138 = \pi0741  & n1281 ;
  assign n28139 = n28115 & n28138 ;
  assign n28140 = ~\pi0156  & ~n28139 ;
  assign n28141 = ~n28137 & n28140 ;
  assign n28142 = ~n28134 & n28141 ;
  assign n28143 = ~\pi0741  & n1289 ;
  assign n28144 = n1287 & n28143 ;
  assign n28145 = n9948 & n28144 ;
  assign n28146 = ~n27269 & n28145 ;
  assign n28147 = ~\pi0156  & ~n11834 ;
  assign n28148 = \pi0741  & ~n22124 ;
  assign n28149 = ~n28084 & n28148 ;
  assign n28150 = ~\pi0156  & \pi0724  ;
  assign n28151 = ~n28149 & n28150 ;
  assign n28152 = ~n28147 & ~n28151 ;
  assign n28153 = ~n28146 & ~n28152 ;
  assign n28154 = ~\pi0057  & \pi0156  ;
  assign n28155 = n6848 & n28154 ;
  assign n28156 = n6861 & n28155 ;
  assign n28157 = ~\pi0832  & ~n28156 ;
  assign n28158 = ~\pi0724  & ~\pi0741  ;
  assign n28159 = ~n28052 & n28158 ;
  assign n28160 = ~n28061 & n28131 ;
  assign n28161 = ~n28159 & ~n28160 ;
  assign n28162 = \pi0724  & ~\pi0741  ;
  assign n28163 = ~\pi0832  & ~n28162 ;
  assign n28164 = ~n28068 & ~n28163 ;
  assign n28165 = n28161 & ~n28164 ;
  assign n28166 = ~n28157 & ~n28165 ;
  assign n28167 = ~n28153 & ~n28166 ;
  assign n28168 = ~n28142 & n28167 ;
  assign n28169 = ~n28130 & ~n28168 ;
  assign n28170 = ~\pi0157  & ~n11834 ;
  assign n28171 = ~\pi0832  & ~n28170 ;
  assign n28172 = ~\pi0760  & \pi0947  ;
  assign n28173 = \pi0299  & n28172 ;
  assign n28174 = ~n21205 & n28173 ;
  assign n28175 = ~n21238 & n28174 ;
  assign n28176 = ~\pi0299  & n28172 ;
  assign n28177 = ~n21740 & n28176 ;
  assign n28178 = ~n21738 & n28177 ;
  assign n28179 = ~n28175 & ~n28178 ;
  assign n28180 = ~\pi0157  & ~n27328 ;
  assign n28181 = n16528 & n21205 ;
  assign n28182 = n16528 & n21237 ;
  assign n28183 = n21232 & n28182 ;
  assign n28184 = ~n28181 & ~n28183 ;
  assign n28185 = ~\pi0039  & n28184 ;
  assign n28186 = ~n28180 & n28185 ;
  assign n28187 = n28179 & n28186 ;
  assign n28188 = ~\pi0038  & ~n28187 ;
  assign n28189 = n6784 & ~n28172 ;
  assign n28190 = n1266 & n28189 ;
  assign n28191 = n22706 & n28190 ;
  assign n28192 = n1358 & n28191 ;
  assign n28193 = \pi0038  & ~n28192 ;
  assign n28194 = \pi0688  & ~n28193 ;
  assign n28195 = \pi0157  & \pi0688  ;
  assign n28196 = ~n22123 & n28195 ;
  assign n28197 = ~n28194 & ~n28196 ;
  assign n28198 = ~n28188 & ~n28197 ;
  assign n28199 = ~\pi0157  & ~n21692 ;
  assign n28200 = n27361 & ~n28199 ;
  assign n28201 = ~\pi0760  & ~n28200 ;
  assign n28202 = ~n16528 & ~n27304 ;
  assign n28203 = ~\pi0157  & n27260 ;
  assign n28204 = ~\pi0157  & n27257 ;
  assign n28205 = ~n27254 & n28204 ;
  assign n28206 = ~n28203 & ~n28205 ;
  assign n28207 = ~n28202 & n28206 ;
  assign n28208 = n28201 & ~n28207 ;
  assign n28209 = ~\pi0157  & \pi0760  ;
  assign n28210 = ~\pi0299  & n28209 ;
  assign n28211 = ~n21692 & n28210 ;
  assign n28212 = \pi0039  & ~n28209 ;
  assign n28213 = ~n21733 & ~n28212 ;
  assign n28214 = ~n28211 & ~n28213 ;
  assign n28215 = ~n28197 & n28214 ;
  assign n28216 = ~n28208 & n28215 ;
  assign n28217 = ~n28198 & ~n28216 ;
  assign n28218 = n11834 & n28217 ;
  assign n28219 = n28171 & ~n28218 ;
  assign n28220 = n27068 & n28179 ;
  assign n28221 = n28186 & n28220 ;
  assign n28222 = ~\pi0038  & ~n28221 ;
  assign n28223 = ~\pi0039  & n28222 ;
  assign n28224 = ~\pi0760  & n27215 ;
  assign n28225 = \pi0760  & ~n27136 ;
  assign n28226 = ~n27132 & n28225 ;
  assign n28227 = ~\pi0157  & ~n28226 ;
  assign n28228 = ~n28224 & n28227 ;
  assign n28229 = \pi0760  & n27084 ;
  assign n28230 = ~n27523 & n28229 ;
  assign n28231 = ~\pi0760  & ~n27343 ;
  assign n28232 = \pi0157  & ~n28231 ;
  assign n28233 = \pi0157  & ~\pi0299  ;
  assign n28234 = ~n27158 & n28233 ;
  assign n28235 = ~n28232 & ~n28234 ;
  assign n28236 = ~n28230 & ~n28235 ;
  assign n28237 = n28222 & ~n28236 ;
  assign n28238 = ~n28228 & n28237 ;
  assign n28239 = ~n28223 & ~n28238 ;
  assign n28240 = ~n26930 & n28192 ;
  assign n28241 = \pi0157  & ~n21757 ;
  assign n28242 = \pi0038  & ~n28241 ;
  assign n28243 = ~n28240 & n28242 ;
  assign n28244 = ~\pi0688  & ~n28243 ;
  assign n28245 = n28171 & n28244 ;
  assign n28246 = n28239 & n28245 ;
  assign n28247 = ~n28219 & ~n28246 ;
  assign n28248 = ~\pi0688  & n26930 ;
  assign n28249 = ~n28172 & ~n28248 ;
  assign n28250 = n1689 & ~n28249 ;
  assign n28251 = ~\pi0157  & ~n1689 ;
  assign n28252 = \pi0832  & ~n28251 ;
  assign n28253 = ~n28250 & n28252 ;
  assign n28254 = n28247 & ~n28253 ;
  assign n28255 = ~\pi0753  & \pi0947  ;
  assign n28256 = ~\pi0702  & n26930 ;
  assign n28257 = ~n28255 & ~n28256 ;
  assign n28258 = n1689 & ~n28257 ;
  assign n28259 = ~\pi0158  & ~n1689 ;
  assign n28260 = \pi0832  & ~n28259 ;
  assign n28261 = ~n28258 & n28260 ;
  assign n28262 = ~\pi0158  & n27215 ;
  assign n28263 = \pi0158  & ~n27343 ;
  assign n28264 = ~\pi0753  & ~n28263 ;
  assign n28265 = ~\pi0299  & ~\pi0753  ;
  assign n28266 = ~n27158 & n28265 ;
  assign n28267 = ~n28264 & ~n28266 ;
  assign n28268 = ~n28262 & ~n28267 ;
  assign n28269 = ~\pi0158  & ~n27136 ;
  assign n28270 = ~n27132 & n28269 ;
  assign n28271 = \pi0158  & n27084 ;
  assign n28272 = ~n27523 & n28271 ;
  assign n28273 = \pi0753  & ~n28272 ;
  assign n28274 = ~n28270 & n28273 ;
  assign n28275 = \pi0039  & ~n28274 ;
  assign n28276 = ~n28268 & n28275 ;
  assign n28277 = ~n27106 & ~n28255 ;
  assign n28278 = \pi0158  & ~n27219 ;
  assign n28279 = ~n27217 & n28278 ;
  assign n28280 = ~\pi0039  & ~n28279 ;
  assign n28281 = ~n28277 & n28280 ;
  assign n28282 = ~\pi0038  & ~n28281 ;
  assign n28283 = ~n28276 & n28282 ;
  assign n28284 = \pi0158  & ~n21757 ;
  assign n28285 = n6784 & ~n28255 ;
  assign n28286 = n1266 & n28285 ;
  assign n28287 = n22706 & n28286 ;
  assign n28288 = n1358 & n28287 ;
  assign n28289 = ~n26930 & n28288 ;
  assign n28290 = ~n28284 & ~n28289 ;
  assign n28291 = \pi0038  & ~n28290 ;
  assign n28292 = ~\pi0702  & n11834 ;
  assign n28293 = ~n28291 & n28292 ;
  assign n28294 = ~n28283 & n28293 ;
  assign n28295 = \pi0299  & \pi0753  ;
  assign n28296 = ~n21205 & n28295 ;
  assign n28297 = ~n21238 & n28296 ;
  assign n28298 = ~\pi0299  & \pi0753  ;
  assign n28299 = ~n21740 & n28298 ;
  assign n28300 = ~n21738 & n28299 ;
  assign n28301 = ~n28297 & ~n28300 ;
  assign n28302 = ~n28279 & n28301 ;
  assign n28303 = n27242 & n28302 ;
  assign n28304 = n1288 & ~n28303 ;
  assign n28305 = ~\pi0038  & ~n28303 ;
  assign n28306 = ~\pi0158  & \pi0753  ;
  assign n28307 = ~\pi0299  & n28306 ;
  assign n28308 = ~n21692 & n28307 ;
  assign n28309 = ~n25541 & n28306 ;
  assign n28310 = ~n28308 & ~n28309 ;
  assign n28311 = n28305 & n28310 ;
  assign n28312 = ~n28304 & ~n28311 ;
  assign n28313 = ~\pi0158  & ~n27247 ;
  assign n28314 = ~n27549 & n28313 ;
  assign n28315 = \pi0158  & ~\pi0299  ;
  assign n28316 = ~n27285 & n28315 ;
  assign n28317 = \pi0158  & n27304 ;
  assign n28318 = ~\pi0753  & ~n28317 ;
  assign n28319 = ~n28316 & n28318 ;
  assign n28320 = ~n28304 & n28319 ;
  assign n28321 = ~n28314 & n28320 ;
  assign n28322 = ~n28312 & ~n28321 ;
  assign n28323 = \pi0038  & \pi0158  ;
  assign n28324 = ~n22123 & n28323 ;
  assign n28325 = \pi0038  & n28288 ;
  assign n28326 = \pi0702  & ~n28325 ;
  assign n28327 = ~n28324 & n28326 ;
  assign n28328 = n11834 & n28327 ;
  assign n28329 = ~n28322 & n28328 ;
  assign n28330 = ~\pi0158  & ~n11834 ;
  assign n28331 = ~\pi0832  & ~n28330 ;
  assign n28332 = ~n28329 & n28331 ;
  assign n28333 = ~n28294 & n28332 ;
  assign n28334 = ~n28261 & ~n28333 ;
  assign n28335 = ~\pi0754  & \pi0947  ;
  assign n28336 = ~\pi0709  & n26930 ;
  assign n28337 = ~n28335 & ~n28336 ;
  assign n28338 = n1689 & ~n28337 ;
  assign n28339 = ~\pi0159  & ~n1689 ;
  assign n28340 = \pi0832  & ~n28339 ;
  assign n28341 = ~n28338 & n28340 ;
  assign n28342 = ~\pi0159  & n27215 ;
  assign n28343 = \pi0159  & ~n27343 ;
  assign n28344 = ~\pi0754  & ~n28343 ;
  assign n28345 = ~\pi0299  & ~\pi0754  ;
  assign n28346 = ~n27158 & n28345 ;
  assign n28347 = ~n28344 & ~n28346 ;
  assign n28348 = ~n28342 & ~n28347 ;
  assign n28349 = ~\pi0159  & ~n27136 ;
  assign n28350 = ~n27132 & n28349 ;
  assign n28351 = \pi0159  & n27084 ;
  assign n28352 = ~n27523 & n28351 ;
  assign n28353 = \pi0754  & ~n28352 ;
  assign n28354 = ~n28350 & n28353 ;
  assign n28355 = \pi0039  & ~n28354 ;
  assign n28356 = ~n28348 & n28355 ;
  assign n28357 = ~n27106 & ~n28335 ;
  assign n28358 = \pi0159  & ~n27219 ;
  assign n28359 = ~n27217 & n28358 ;
  assign n28360 = ~\pi0039  & ~n28359 ;
  assign n28361 = ~n28357 & n28360 ;
  assign n28362 = ~\pi0038  & ~n28361 ;
  assign n28363 = ~n28356 & n28362 ;
  assign n28364 = \pi0159  & ~n21757 ;
  assign n28365 = n6784 & ~n28335 ;
  assign n28366 = n1266 & n28365 ;
  assign n28367 = n22706 & n28366 ;
  assign n28368 = n1358 & n28367 ;
  assign n28369 = ~n26930 & n28368 ;
  assign n28370 = ~n28364 & ~n28369 ;
  assign n28371 = \pi0038  & ~n28370 ;
  assign n28372 = ~\pi0709  & n11834 ;
  assign n28373 = ~n28371 & n28372 ;
  assign n28374 = ~n28363 & n28373 ;
  assign n28375 = \pi0299  & \pi0754  ;
  assign n28376 = ~n21205 & n28375 ;
  assign n28377 = ~n21238 & n28376 ;
  assign n28378 = ~\pi0299  & \pi0754  ;
  assign n28379 = ~n21740 & n28378 ;
  assign n28380 = ~n21738 & n28379 ;
  assign n28381 = ~n28377 & ~n28380 ;
  assign n28382 = ~n28359 & n28381 ;
  assign n28383 = n27242 & n28382 ;
  assign n28384 = n1288 & ~n28383 ;
  assign n28385 = ~\pi0038  & ~n28383 ;
  assign n28386 = ~\pi0159  & \pi0754  ;
  assign n28387 = ~\pi0299  & n28386 ;
  assign n28388 = ~n21692 & n28387 ;
  assign n28389 = ~n25541 & n28386 ;
  assign n28390 = ~n28388 & ~n28389 ;
  assign n28391 = n28385 & n28390 ;
  assign n28392 = ~n28384 & ~n28391 ;
  assign n28393 = ~\pi0159  & ~n27247 ;
  assign n28394 = ~n27549 & n28393 ;
  assign n28395 = \pi0159  & ~\pi0299  ;
  assign n28396 = ~n27285 & n28395 ;
  assign n28397 = \pi0159  & n27304 ;
  assign n28398 = ~\pi0754  & ~n28397 ;
  assign n28399 = ~n28396 & n28398 ;
  assign n28400 = ~n28384 & n28399 ;
  assign n28401 = ~n28394 & n28400 ;
  assign n28402 = ~n28392 & ~n28401 ;
  assign n28403 = \pi0038  & \pi0159  ;
  assign n28404 = ~n22123 & n28403 ;
  assign n28405 = \pi0038  & n28368 ;
  assign n28406 = \pi0709  & ~n28405 ;
  assign n28407 = ~n28404 & n28406 ;
  assign n28408 = n11834 & n28407 ;
  assign n28409 = ~n28402 & n28408 ;
  assign n28410 = ~\pi0159  & ~n11834 ;
  assign n28411 = ~\pi0832  & ~n28410 ;
  assign n28412 = ~n28409 & n28411 ;
  assign n28413 = ~n28374 & n28412 ;
  assign n28414 = ~n28341 & ~n28413 ;
  assign n28415 = ~\pi0756  & \pi0947  ;
  assign n28416 = ~\pi0734  & n26930 ;
  assign n28417 = ~n28415 & ~n28416 ;
  assign n28418 = n1689 & ~n28417 ;
  assign n28419 = ~\pi0160  & ~n1689 ;
  assign n28420 = \pi0832  & ~n28419 ;
  assign n28421 = ~n28418 & n28420 ;
  assign n28422 = ~\pi0160  & ~n11834 ;
  assign n28423 = ~\pi0832  & ~n28422 ;
  assign n28424 = ~n28421 & ~n28423 ;
  assign n28425 = n6784 & ~n28415 ;
  assign n28426 = n1266 & n28425 ;
  assign n28427 = n22706 & n28426 ;
  assign n28428 = n1358 & n28427 ;
  assign n28429 = ~n26930 & n28428 ;
  assign n28430 = \pi0160  & ~n21757 ;
  assign n28431 = \pi0038  & ~n28430 ;
  assign n28432 = ~n28429 & n28431 ;
  assign n28433 = ~\pi0734  & ~n28432 ;
  assign n28434 = ~\pi0160  & ~n27328 ;
  assign n28435 = ~\pi0160  & \pi0299  ;
  assign n28436 = n21205 & n28435 ;
  assign n28437 = n21237 & n28435 ;
  assign n28438 = n21232 & n28437 ;
  assign n28439 = ~n28436 & ~n28438 ;
  assign n28440 = ~\pi0039  & n28439 ;
  assign n28441 = ~n28434 & n28440 ;
  assign n28442 = \pi0299  & n28415 ;
  assign n28443 = ~n21205 & n28442 ;
  assign n28444 = ~n21238 & n28443 ;
  assign n28445 = ~\pi0299  & n28415 ;
  assign n28446 = ~n21740 & n28445 ;
  assign n28447 = ~n21738 & n28446 ;
  assign n28448 = ~n28444 & ~n28447 ;
  assign n28449 = n27068 & n28448 ;
  assign n28450 = n28441 & n28449 ;
  assign n28451 = ~\pi0038  & ~n28450 ;
  assign n28452 = n28433 & ~n28451 ;
  assign n28453 = ~\pi0160  & n27132 ;
  assign n28454 = \pi0160  & ~n27084 ;
  assign n28455 = \pi0160  & ~\pi0299  ;
  assign n28456 = ~n21692 & n28455 ;
  assign n28457 = ~n28454 & ~n28456 ;
  assign n28458 = ~n27136 & n28457 ;
  assign n28459 = ~n28453 & n28458 ;
  assign n28460 = \pi0756  & ~n28459 ;
  assign n28461 = ~\pi0160  & n27215 ;
  assign n28462 = \pi0160  & ~n27343 ;
  assign n28463 = ~\pi0756  & ~n28462 ;
  assign n28464 = ~\pi0299  & ~\pi0756  ;
  assign n28465 = ~n27158 & n28464 ;
  assign n28466 = ~n28463 & ~n28465 ;
  assign n28467 = ~n28461 & ~n28466 ;
  assign n28468 = ~n28460 & ~n28467 ;
  assign n28469 = \pi0039  & n28433 ;
  assign n28470 = ~n28468 & n28469 ;
  assign n28471 = ~n28452 & ~n28470 ;
  assign n28472 = n28441 & n28448 ;
  assign n28473 = ~\pi0038  & ~n28472 ;
  assign n28474 = \pi0038  & ~n28428 ;
  assign n28475 = \pi0734  & ~n28474 ;
  assign n28476 = \pi0160  & \pi0734  ;
  assign n28477 = ~n22123 & n28476 ;
  assign n28478 = ~n28475 & ~n28477 ;
  assign n28479 = ~n28473 & ~n28478 ;
  assign n28480 = ~\pi0160  & ~n21692 ;
  assign n28481 = n27361 & ~n28480 ;
  assign n28482 = ~\pi0756  & ~n28481 ;
  assign n28483 = ~n27304 & ~n28435 ;
  assign n28484 = ~\pi0160  & n27260 ;
  assign n28485 = ~\pi0160  & n27257 ;
  assign n28486 = ~n27254 & n28485 ;
  assign n28487 = ~n28484 & ~n28486 ;
  assign n28488 = ~n28483 & n28487 ;
  assign n28489 = n28482 & ~n28488 ;
  assign n28490 = ~\pi0160  & \pi0756  ;
  assign n28491 = ~\pi0299  & n28490 ;
  assign n28492 = ~n21692 & n28491 ;
  assign n28493 = \pi0039  & ~n28490 ;
  assign n28494 = ~n21733 & ~n28493 ;
  assign n28495 = ~n28492 & ~n28494 ;
  assign n28496 = ~n28478 & n28495 ;
  assign n28497 = ~n28489 & n28496 ;
  assign n28498 = ~n28479 & ~n28497 ;
  assign n28499 = n11834 & ~n28421 ;
  assign n28500 = n28498 & n28499 ;
  assign n28501 = n28471 & n28500 ;
  assign n28502 = ~n28424 & ~n28501 ;
  assign n28503 = ~\pi0161  & ~n11834 ;
  assign n28504 = ~\pi0832  & ~n28503 ;
  assign n28505 = \pi0758  & \pi0947  ;
  assign n28506 = n1689 & ~n28505 ;
  assign n28507 = \pi0736  & n26930 ;
  assign n28508 = n28506 & ~n28507 ;
  assign n28509 = ~\pi0161  & ~n1689 ;
  assign n28510 = \pi0832  & ~n28509 ;
  assign n28511 = ~n28508 & n28510 ;
  assign n28512 = ~n28504 & ~n28511 ;
  assign n28513 = \pi0161  & ~\pi0758  ;
  assign n28514 = ~n25542 & n28513 ;
  assign n28515 = \pi0039  & ~n28514 ;
  assign n28516 = \pi0161  & ~n27328 ;
  assign n28517 = \pi0161  & \pi0299  ;
  assign n28518 = n21205 & n28517 ;
  assign n28519 = n21237 & n28517 ;
  assign n28520 = n21232 & n28519 ;
  assign n28521 = ~n28518 & ~n28520 ;
  assign n28522 = ~\pi0039  & n28521 ;
  assign n28523 = ~n28516 & n28522 ;
  assign n28524 = \pi0299  & n28505 ;
  assign n28525 = ~n21205 & n28524 ;
  assign n28526 = ~n21238 & n28525 ;
  assign n28527 = ~\pi0299  & n28505 ;
  assign n28528 = ~n21740 & n28527 ;
  assign n28529 = ~n21738 & n28528 ;
  assign n28530 = ~n28526 & ~n28529 ;
  assign n28531 = n28523 & n28530 ;
  assign n28532 = ~\pi0038  & ~n28531 ;
  assign n28533 = ~n28515 & n28532 ;
  assign n28534 = \pi0161  & n27121 ;
  assign n28535 = ~n27730 & n28534 ;
  assign n28536 = n21694 & n28534 ;
  assign n28537 = ~n21711 & n28536 ;
  assign n28538 = ~n28535 & ~n28537 ;
  assign n28539 = n27737 & n28538 ;
  assign n28540 = ~n27729 & ~n28539 ;
  assign n28541 = ~\pi0161  & n2352 ;
  assign n28542 = n21285 & n28541 ;
  assign n28543 = n27257 & ~n28542 ;
  assign n28544 = n28540 & n28543 ;
  assign n28545 = \pi0161  & \pi0215  ;
  assign n28546 = ~n27082 & n28545 ;
  assign n28547 = ~n21724 & n28546 ;
  assign n28548 = n27747 & ~n28547 ;
  assign n28549 = ~n28544 & n28548 ;
  assign n28550 = ~\pi0161  & n21612 ;
  assign n28551 = ~n21606 & n28550 ;
  assign n28552 = ~\pi0223  & ~n28551 ;
  assign n28553 = ~n27753 & n28552 ;
  assign n28554 = ~\pi0161  & ~n21651 ;
  assign n28555 = ~\pi0161  & n6761 ;
  assign n28556 = ~n21685 & n28555 ;
  assign n28557 = ~n28554 & ~n28556 ;
  assign n28558 = n27204 & n28557 ;
  assign n28559 = ~\pi0223  & n27766 ;
  assign n28560 = ~n21285 & n28559 ;
  assign n28561 = \pi0161  & n2165 ;
  assign n28562 = ~\pi0223  & n28561 ;
  assign n28563 = n21285 & n28562 ;
  assign n28564 = ~n28560 & ~n28563 ;
  assign n28565 = ~\pi0299  & n28564 ;
  assign n28566 = ~n28558 & n28565 ;
  assign n28567 = ~n28553 & n28566 ;
  assign n28568 = \pi0758  & ~n28567 ;
  assign n28569 = n28532 & n28568 ;
  assign n28570 = ~n28549 & n28569 ;
  assign n28571 = ~n28533 & ~n28570 ;
  assign n28572 = n1354 & ~n28505 ;
  assign n28573 = n21755 & n28572 ;
  assign n28574 = n1358 & n28573 ;
  assign n28575 = \pi0038  & ~n28574 ;
  assign n28576 = ~\pi0736  & ~n28575 ;
  assign n28577 = ~\pi0161  & ~\pi0736  ;
  assign n28578 = ~n22123 & n28577 ;
  assign n28579 = ~n28576 & ~n28578 ;
  assign n28580 = n28571 & ~n28579 ;
  assign n28581 = n11834 & ~n28511 ;
  assign n28582 = n28580 & n28581 ;
  assign n28583 = n27068 & n28530 ;
  assign n28584 = n28523 & n28583 ;
  assign n28585 = ~\pi0038  & ~n28584 ;
  assign n28586 = ~n26930 & n28574 ;
  assign n28587 = ~\pi0161  & ~n21757 ;
  assign n28588 = \pi0038  & ~n28587 ;
  assign n28589 = ~n28586 & n28588 ;
  assign n28590 = ~n28585 & ~n28589 ;
  assign n28591 = ~\pi0299  & ~n28558 ;
  assign n28592 = ~\pi0161  & n2165 ;
  assign n28593 = ~\pi0223  & ~n28592 ;
  assign n28594 = n21285 & n28593 ;
  assign n28595 = ~n27798 & ~n28594 ;
  assign n28596 = ~n28551 & ~n28595 ;
  assign n28597 = ~n27753 & n28596 ;
  assign n28598 = ~n27805 & ~n28595 ;
  assign n28599 = ~n27751 & n28598 ;
  assign n28600 = n27206 & n28557 ;
  assign n28601 = ~n28599 & ~n28600 ;
  assign n28602 = ~n28597 & n28601 ;
  assign n28603 = n28591 & n28602 ;
  assign n28604 = ~n27813 & ~n28542 ;
  assign n28605 = ~\pi0215  & n28604 ;
  assign n28606 = ~\pi0161  & ~n21728 ;
  assign n28607 = \pi0215  & ~n28606 ;
  assign n28608 = ~n21724 & n28607 ;
  assign n28609 = \pi0299  & ~n28608 ;
  assign n28610 = ~n28605 & n28609 ;
  assign n28611 = n27821 & n28609 ;
  assign n28612 = n28538 & n28611 ;
  assign n28613 = ~n28610 & ~n28612 ;
  assign n28614 = \pi0758  & n28613 ;
  assign n28615 = ~n28603 & n28614 ;
  assign n28616 = ~n27828 & n28552 ;
  assign n28617 = n21285 & n28561 ;
  assign n28618 = ~n27831 & ~n28617 ;
  assign n28619 = ~\pi0223  & ~n28618 ;
  assign n28620 = ~\pi0299  & ~n28600 ;
  assign n28621 = ~n28619 & n28620 ;
  assign n28622 = ~n28616 & n28621 ;
  assign n28623 = ~\pi0758  & n27843 ;
  assign n28624 = n28608 & n28623 ;
  assign n28625 = ~n25548 & ~n28624 ;
  assign n28626 = n27736 & n28538 ;
  assign n28627 = ~\pi0215  & ~\pi0758  ;
  assign n28628 = ~n27128 & n28627 ;
  assign n28629 = n28604 & n28628 ;
  assign n28630 = ~n28626 & n28629 ;
  assign n28631 = n28625 & ~n28630 ;
  assign n28632 = ~n28622 & ~n28631 ;
  assign n28633 = ~n28615 & ~n28632 ;
  assign n28634 = \pi0039  & ~n28589 ;
  assign n28635 = n28633 & n28634 ;
  assign n28636 = ~n28590 & ~n28635 ;
  assign n28637 = \pi0736  & n28581 ;
  assign n28638 = ~n28636 & n28637 ;
  assign n28639 = ~n28582 & ~n28638 ;
  assign n28640 = ~n28512 & n28639 ;
  assign n28641 = ~\pi0761  & \pi0947  ;
  assign n28642 = ~\pi0738  & n26930 ;
  assign n28643 = ~n28641 & ~n28642 ;
  assign n28644 = n1689 & ~n28643 ;
  assign n28645 = ~\pi0162  & ~n1689 ;
  assign n28646 = \pi0832  & ~n28645 ;
  assign n28647 = ~n28644 & n28646 ;
  assign n28648 = ~\pi0162  & ~n11834 ;
  assign n28649 = ~\pi0832  & ~n28648 ;
  assign n28650 = ~n28647 & ~n28649 ;
  assign n28651 = n6784 & ~n28641 ;
  assign n28652 = n1266 & n28651 ;
  assign n28653 = n22706 & n28652 ;
  assign n28654 = n1358 & n28653 ;
  assign n28655 = ~n26930 & n28654 ;
  assign n28656 = \pi0162  & ~n21757 ;
  assign n28657 = \pi0038  & ~n28656 ;
  assign n28658 = ~n28655 & n28657 ;
  assign n28659 = ~\pi0738  & ~n28658 ;
  assign n28660 = ~\pi0162  & ~n27328 ;
  assign n28661 = ~\pi0162  & \pi0299  ;
  assign n28662 = n21205 & n28661 ;
  assign n28663 = n21237 & n28661 ;
  assign n28664 = n21232 & n28663 ;
  assign n28665 = ~n28662 & ~n28664 ;
  assign n28666 = ~\pi0039  & n28665 ;
  assign n28667 = ~n28660 & n28666 ;
  assign n28668 = \pi0299  & n28641 ;
  assign n28669 = ~n21205 & n28668 ;
  assign n28670 = ~n21238 & n28669 ;
  assign n28671 = ~\pi0299  & n28641 ;
  assign n28672 = ~n21740 & n28671 ;
  assign n28673 = ~n21738 & n28672 ;
  assign n28674 = ~n28670 & ~n28673 ;
  assign n28675 = n27068 & n28674 ;
  assign n28676 = n28667 & n28675 ;
  assign n28677 = ~\pi0038  & ~n28676 ;
  assign n28678 = n28659 & ~n28677 ;
  assign n28679 = \pi0162  & ~n27084 ;
  assign n28680 = \pi0162  & ~\pi0299  ;
  assign n28681 = ~n21692 & n28680 ;
  assign n28682 = ~n28679 & ~n28681 ;
  assign n28683 = \pi0761  & ~n28682 ;
  assign n28684 = \pi0761  & ~n18435 ;
  assign n28685 = ~n27348 & n28684 ;
  assign n28686 = ~n28683 & ~n28685 ;
  assign n28687 = ~\pi0162  & n27215 ;
  assign n28688 = \pi0162  & ~n27343 ;
  assign n28689 = ~\pi0761  & ~n28688 ;
  assign n28690 = ~\pi0299  & ~\pi0761  ;
  assign n28691 = ~n27158 & n28690 ;
  assign n28692 = ~n28689 & ~n28691 ;
  assign n28693 = ~n28687 & ~n28692 ;
  assign n28694 = n28686 & ~n28693 ;
  assign n28695 = \pi0039  & n28659 ;
  assign n28696 = ~n28694 & n28695 ;
  assign n28697 = ~n28678 & ~n28696 ;
  assign n28698 = ~n27299 & ~n27301 ;
  assign n28699 = ~n27297 & n28698 ;
  assign n28700 = n18435 & ~n28699 ;
  assign n28701 = ~\pi0761  & ~n28700 ;
  assign n28702 = ~n27247 & n28701 ;
  assign n28703 = ~n27549 & n28702 ;
  assign n28704 = \pi0162  & ~n28700 ;
  assign n28705 = ~n27247 & n28704 ;
  assign n28706 = ~\pi0761  & ~n28705 ;
  assign n28707 = ~\pi0162  & ~n28705 ;
  assign n28708 = ~n25542 & n28707 ;
  assign n28709 = ~n28706 & ~n28708 ;
  assign n28710 = ~n28703 & ~n28709 ;
  assign n28711 = \pi0038  & ~n28654 ;
  assign n28712 = \pi0738  & ~n28711 ;
  assign n28713 = \pi0162  & \pi0738  ;
  assign n28714 = ~n22123 & n28713 ;
  assign n28715 = ~n28712 & ~n28714 ;
  assign n28716 = \pi0039  & ~n28715 ;
  assign n28717 = ~n28710 & n28716 ;
  assign n28718 = \pi0038  & ~n28715 ;
  assign n28719 = n28674 & ~n28715 ;
  assign n28720 = n28667 & n28719 ;
  assign n28721 = ~n28718 & ~n28720 ;
  assign n28722 = n11834 & n28721 ;
  assign n28723 = ~n28717 & n28722 ;
  assign n28724 = ~n28647 & n28723 ;
  assign n28725 = n28697 & n28724 ;
  assign n28726 = ~n28650 & ~n28725 ;
  assign n28727 = ~\pi0163  & ~n11834 ;
  assign n28728 = ~\pi0832  & ~n28727 ;
  assign n28729 = ~\pi0777  & \pi0947  ;
  assign n28730 = ~\pi0737  & n26930 ;
  assign n28731 = ~n28729 & ~n28730 ;
  assign n28732 = n1689 & ~n28731 ;
  assign n28733 = ~\pi0163  & ~n1689 ;
  assign n28734 = \pi0832  & ~n28733 ;
  assign n28735 = ~n28732 & n28734 ;
  assign n28736 = ~n28728 & ~n28735 ;
  assign n28737 = n6784 & ~n28729 ;
  assign n28738 = n1266 & n28737 ;
  assign n28739 = n22706 & n28738 ;
  assign n28740 = n1358 & n28739 ;
  assign n28741 = ~n26930 & n28740 ;
  assign n28742 = \pi0163  & ~n21757 ;
  assign n28743 = \pi0038  & ~n28742 ;
  assign n28744 = ~n28741 & n28743 ;
  assign n28745 = ~\pi0737  & ~n28744 ;
  assign n28746 = ~\pi0163  & ~n27328 ;
  assign n28747 = n17723 & n21205 ;
  assign n28748 = n17723 & n21237 ;
  assign n28749 = n21232 & n28748 ;
  assign n28750 = ~n28747 & ~n28749 ;
  assign n28751 = ~\pi0039  & n28750 ;
  assign n28752 = ~n28746 & n28751 ;
  assign n28753 = \pi0299  & n28729 ;
  assign n28754 = ~n21205 & n28753 ;
  assign n28755 = ~n21238 & n28754 ;
  assign n28756 = ~\pi0299  & n28729 ;
  assign n28757 = ~n21740 & n28756 ;
  assign n28758 = ~n21738 & n28757 ;
  assign n28759 = ~n28755 & ~n28758 ;
  assign n28760 = n27068 & n28759 ;
  assign n28761 = n28752 & n28760 ;
  assign n28762 = ~\pi0038  & ~n28761 ;
  assign n28763 = n28745 & ~n28762 ;
  assign n28764 = ~\pi0163  & n27132 ;
  assign n28765 = \pi0163  & ~n27084 ;
  assign n28766 = \pi0163  & ~\pi0299  ;
  assign n28767 = ~n21692 & n28766 ;
  assign n28768 = ~n28765 & ~n28767 ;
  assign n28769 = ~n27136 & n28768 ;
  assign n28770 = ~n28764 & n28769 ;
  assign n28771 = \pi0777  & ~n28770 ;
  assign n28772 = ~\pi0163  & n27215 ;
  assign n28773 = \pi0163  & ~n27343 ;
  assign n28774 = ~\pi0777  & ~n28773 ;
  assign n28775 = ~\pi0299  & ~\pi0777  ;
  assign n28776 = ~n27158 & n28775 ;
  assign n28777 = ~n28774 & ~n28776 ;
  assign n28778 = ~n28772 & ~n28777 ;
  assign n28779 = ~n28771 & ~n28778 ;
  assign n28780 = \pi0039  & n28745 ;
  assign n28781 = ~n28779 & n28780 ;
  assign n28782 = ~n28763 & ~n28781 ;
  assign n28783 = n28752 & n28759 ;
  assign n28784 = ~\pi0038  & ~n28783 ;
  assign n28785 = \pi0038  & ~n28740 ;
  assign n28786 = \pi0737  & ~n28785 ;
  assign n28787 = \pi0163  & \pi0737  ;
  assign n28788 = ~n22123 & n28787 ;
  assign n28789 = ~n28786 & ~n28788 ;
  assign n28790 = ~n28784 & ~n28789 ;
  assign n28791 = ~\pi0163  & ~n21692 ;
  assign n28792 = n27361 & ~n28791 ;
  assign n28793 = ~\pi0777  & ~n28792 ;
  assign n28794 = ~n17723 & ~n27304 ;
  assign n28795 = ~\pi0163  & n27260 ;
  assign n28796 = ~\pi0163  & n27257 ;
  assign n28797 = ~n27254 & n28796 ;
  assign n28798 = ~n28795 & ~n28797 ;
  assign n28799 = ~n28794 & n28798 ;
  assign n28800 = n28793 & ~n28799 ;
  assign n28801 = ~\pi0163  & \pi0777  ;
  assign n28802 = ~\pi0299  & n28801 ;
  assign n28803 = ~n21692 & n28802 ;
  assign n28804 = \pi0039  & ~n28801 ;
  assign n28805 = ~n21733 & ~n28804 ;
  assign n28806 = ~n28803 & ~n28805 ;
  assign n28807 = ~n28789 & n28806 ;
  assign n28808 = ~n28800 & n28807 ;
  assign n28809 = ~n28790 & ~n28808 ;
  assign n28810 = n11834 & ~n28735 ;
  assign n28811 = n28809 & n28810 ;
  assign n28812 = n28782 & n28811 ;
  assign n28813 = ~n28736 & ~n28812 ;
  assign n28814 = ~\pi0752  & \pi0947  ;
  assign n28815 = \pi0703  & n26930 ;
  assign n28816 = ~n28814 & ~n28815 ;
  assign n28817 = n1689 & ~n28816 ;
  assign n28818 = ~\pi0164  & ~n1689 ;
  assign n28819 = \pi0832  & ~n28818 ;
  assign n28820 = ~n28817 & n28819 ;
  assign n28821 = ~\pi0164  & ~n11834 ;
  assign n28822 = ~\pi0832  & ~n28821 ;
  assign n28823 = ~n28820 & ~n28822 ;
  assign n28824 = n11834 & ~n28820 ;
  assign n28825 = ~n28823 & ~n28824 ;
  assign n28826 = \pi0164  & ~n27085 ;
  assign n28827 = ~n27069 & n28826 ;
  assign n28828 = ~n27061 & n28827 ;
  assign n28829 = ~\pi0038  & ~n28828 ;
  assign n28830 = ~\pi0164  & ~n21757 ;
  assign n28831 = n27096 & ~n28830 ;
  assign n28832 = \pi0752  & ~n28831 ;
  assign n28833 = ~n28829 & n28832 ;
  assign n28834 = ~\pi0164  & \pi0752  ;
  assign n28835 = ~n28831 & n28834 ;
  assign n28836 = n27107 & n28835 ;
  assign n28837 = n27137 & n28835 ;
  assign n28838 = ~n27132 & n28837 ;
  assign n28839 = ~n28836 & ~n28838 ;
  assign n28840 = ~n28833 & n28839 ;
  assign n28841 = \pi0703  & ~n28840 ;
  assign n28842 = ~\pi0164  & ~n27223 ;
  assign n28843 = ~n27216 & n28842 ;
  assign n28844 = \pi0164  & ~n27173 ;
  assign n28845 = ~n27167 & n28844 ;
  assign n28846 = ~n27159 & n28845 ;
  assign n28847 = ~\pi0038  & ~n28846 ;
  assign n28848 = ~n28843 & n28847 ;
  assign n28849 = ~\pi0752  & ~n27990 ;
  assign n28850 = ~\pi0164  & ~\pi0752  ;
  assign n28851 = ~n27144 & n28850 ;
  assign n28852 = ~n28849 & ~n28851 ;
  assign n28853 = \pi0703  & ~n28852 ;
  assign n28854 = ~n28848 & n28853 ;
  assign n28855 = ~n28841 & ~n28854 ;
  assign n28856 = ~\pi0752  & ~\pi0947  ;
  assign n28857 = n25039 & n28856 ;
  assign n28858 = ~n28850 & ~n28857 ;
  assign n28859 = ~n27269 & ~n28858 ;
  assign n28860 = ~\pi0164  & n21770 ;
  assign n28861 = ~n21734 & n28860 ;
  assign n28862 = \pi0038  & ~\pi0164  ;
  assign n28863 = ~n22123 & n28862 ;
  assign n28864 = \pi0752  & ~n28863 ;
  assign n28865 = ~n28861 & n28864 ;
  assign n28866 = \pi0164  & ~n27310 ;
  assign n28867 = ~n27308 & n28866 ;
  assign n28868 = ~\pi0703  & ~n28867 ;
  assign n28869 = ~n28865 & n28868 ;
  assign n28870 = ~n28859 & n28869 ;
  assign n28871 = ~n28823 & ~n28870 ;
  assign n28872 = n28855 & n28871 ;
  assign n28873 = ~n28825 & ~n28872 ;
  assign n28874 = ~\pi0774  & \pi0947  ;
  assign n28875 = \pi0687  & n26930 ;
  assign n28876 = ~n28874 & ~n28875 ;
  assign n28877 = n1689 & ~n28876 ;
  assign n28878 = ~\pi0165  & ~n1689 ;
  assign n28879 = \pi0832  & ~n28878 ;
  assign n28880 = ~n28877 & n28879 ;
  assign n28881 = ~\pi0165  & ~n11834 ;
  assign n28882 = ~\pi0832  & ~n28881 ;
  assign n28883 = ~n28880 & ~n28882 ;
  assign n28884 = n11834 & ~n28880 ;
  assign n28885 = ~n28883 & ~n28884 ;
  assign n28886 = \pi0165  & ~n27085 ;
  assign n28887 = ~n27069 & n28886 ;
  assign n28888 = ~n27061 & n28887 ;
  assign n28889 = ~\pi0038  & ~n28888 ;
  assign n28890 = ~\pi0165  & ~n21757 ;
  assign n28891 = n27096 & ~n28890 ;
  assign n28892 = \pi0774  & ~n28891 ;
  assign n28893 = ~n28889 & n28892 ;
  assign n28894 = ~\pi0165  & \pi0774  ;
  assign n28895 = ~n28891 & n28894 ;
  assign n28896 = n27107 & n28895 ;
  assign n28897 = n27137 & n28895 ;
  assign n28898 = ~n27132 & n28897 ;
  assign n28899 = ~n28896 & ~n28898 ;
  assign n28900 = ~n28893 & n28899 ;
  assign n28901 = \pi0687  & ~n28900 ;
  assign n28902 = ~\pi0165  & ~n27223 ;
  assign n28903 = ~n27216 & n28902 ;
  assign n28904 = \pi0165  & ~n27173 ;
  assign n28905 = ~n27167 & n28904 ;
  assign n28906 = ~n27159 & n28905 ;
  assign n28907 = ~\pi0038  & ~n28906 ;
  assign n28908 = ~n28903 & n28907 ;
  assign n28909 = ~\pi0774  & ~n27990 ;
  assign n28910 = ~\pi0165  & ~\pi0774  ;
  assign n28911 = ~n27144 & n28910 ;
  assign n28912 = ~n28909 & ~n28911 ;
  assign n28913 = \pi0687  & ~n28912 ;
  assign n28914 = ~n28908 & n28913 ;
  assign n28915 = ~n28901 & ~n28914 ;
  assign n28916 = ~\pi0774  & ~\pi0947  ;
  assign n28917 = n25039 & n28916 ;
  assign n28918 = ~n28910 & ~n28917 ;
  assign n28919 = ~n27269 & ~n28918 ;
  assign n28920 = ~\pi0165  & n21770 ;
  assign n28921 = ~n21734 & n28920 ;
  assign n28922 = \pi0038  & ~\pi0165  ;
  assign n28923 = ~n22123 & n28922 ;
  assign n28924 = \pi0774  & ~n28923 ;
  assign n28925 = ~n28921 & n28924 ;
  assign n28926 = \pi0165  & ~n27310 ;
  assign n28927 = ~n27308 & n28926 ;
  assign n28928 = ~\pi0687  & ~n28927 ;
  assign n28929 = ~n28925 & n28928 ;
  assign n28930 = ~n28919 & n28929 ;
  assign n28931 = ~n28883 & ~n28930 ;
  assign n28932 = n28915 & n28931 ;
  assign n28933 = ~n28885 & ~n28932 ;
  assign n28934 = ~\pi0166  & ~n11834 ;
  assign n28935 = ~\pi0832  & ~n28934 ;
  assign n28936 = \pi0772  & \pi0947  ;
  assign n28937 = n1689 & ~n28936 ;
  assign n28938 = \pi0727  & n26930 ;
  assign n28939 = n28937 & ~n28938 ;
  assign n28940 = ~\pi0166  & ~n1689 ;
  assign n28941 = \pi0832  & ~n28940 ;
  assign n28942 = ~n28939 & n28941 ;
  assign n28943 = ~n28935 & ~n28942 ;
  assign n28944 = \pi0166  & ~\pi0772  ;
  assign n28945 = ~n25542 & n28944 ;
  assign n28946 = \pi0039  & ~n28945 ;
  assign n28947 = \pi0166  & ~n27328 ;
  assign n28948 = \pi0166  & \pi0299  ;
  assign n28949 = n21205 & n28948 ;
  assign n28950 = n21237 & n28948 ;
  assign n28951 = n21232 & n28950 ;
  assign n28952 = ~n28949 & ~n28951 ;
  assign n28953 = ~\pi0039  & n28952 ;
  assign n28954 = ~n28947 & n28953 ;
  assign n28955 = \pi0299  & n28936 ;
  assign n28956 = ~n21205 & n28955 ;
  assign n28957 = ~n21238 & n28956 ;
  assign n28958 = ~\pi0299  & n28936 ;
  assign n28959 = ~n21740 & n28958 ;
  assign n28960 = ~n21738 & n28959 ;
  assign n28961 = ~n28957 & ~n28960 ;
  assign n28962 = n28954 & n28961 ;
  assign n28963 = ~\pi0038  & ~n28962 ;
  assign n28964 = ~n28946 & n28963 ;
  assign n28965 = \pi0166  & n27121 ;
  assign n28966 = ~n27730 & n28965 ;
  assign n28967 = n21694 & n28965 ;
  assign n28968 = ~n21711 & n28967 ;
  assign n28969 = ~n28966 & ~n28968 ;
  assign n28970 = n27737 & n28969 ;
  assign n28971 = ~n27729 & ~n28970 ;
  assign n28972 = ~\pi0166  & n2352 ;
  assign n28973 = n21285 & n28972 ;
  assign n28974 = n27257 & ~n28973 ;
  assign n28975 = n28971 & n28974 ;
  assign n28976 = \pi0166  & \pi0215  ;
  assign n28977 = ~n27082 & n28976 ;
  assign n28978 = ~n21724 & n28977 ;
  assign n28979 = n27747 & ~n28978 ;
  assign n28980 = ~n28975 & n28979 ;
  assign n28981 = ~\pi0166  & n21612 ;
  assign n28982 = ~n21606 & n28981 ;
  assign n28983 = ~\pi0223  & ~n28982 ;
  assign n28984 = ~n27753 & n28983 ;
  assign n28985 = ~\pi0166  & ~n21651 ;
  assign n28986 = ~\pi0166  & n6761 ;
  assign n28987 = ~n21685 & n28986 ;
  assign n28988 = ~n28985 & ~n28987 ;
  assign n28989 = n27204 & n28988 ;
  assign n28990 = \pi0166  & n2165 ;
  assign n28991 = ~\pi0223  & n28990 ;
  assign n28992 = n21285 & n28991 ;
  assign n28993 = ~n28560 & ~n28992 ;
  assign n28994 = ~\pi0299  & n28993 ;
  assign n28995 = ~n28989 & n28994 ;
  assign n28996 = ~n28984 & n28995 ;
  assign n28997 = \pi0772  & ~n28996 ;
  assign n28998 = n28963 & n28997 ;
  assign n28999 = ~n28980 & n28998 ;
  assign n29000 = ~n28964 & ~n28999 ;
  assign n29001 = n1354 & ~n28936 ;
  assign n29002 = n21755 & n29001 ;
  assign n29003 = n1358 & n29002 ;
  assign n29004 = \pi0038  & ~n29003 ;
  assign n29005 = ~\pi0727  & ~n29004 ;
  assign n29006 = ~\pi0166  & ~\pi0727  ;
  assign n29007 = ~n22123 & n29006 ;
  assign n29008 = ~n29005 & ~n29007 ;
  assign n29009 = n29000 & ~n29008 ;
  assign n29010 = n11834 & ~n28942 ;
  assign n29011 = n29009 & n29010 ;
  assign n29012 = n27068 & n28961 ;
  assign n29013 = n28954 & n29012 ;
  assign n29014 = ~\pi0038  & ~n29013 ;
  assign n29015 = ~n26930 & n29003 ;
  assign n29016 = ~\pi0166  & ~n21757 ;
  assign n29017 = \pi0038  & ~n29016 ;
  assign n29018 = ~n29015 & n29017 ;
  assign n29019 = ~n29014 & ~n29018 ;
  assign n29020 = ~n27751 & ~n27805 ;
  assign n29021 = ~\pi0166  & n2165 ;
  assign n29022 = ~\pi0223  & ~n29021 ;
  assign n29023 = n21285 & n29022 ;
  assign n29024 = ~n27798 & ~n29023 ;
  assign n29025 = n29020 & ~n29024 ;
  assign n29026 = ~n21606 & n21612 ;
  assign n29027 = ~n26930 & ~n29026 ;
  assign n29028 = ~n28982 & ~n29024 ;
  assign n29029 = ~n29027 & n29028 ;
  assign n29030 = ~n29025 & ~n29029 ;
  assign n29031 = ~\pi0299  & ~n28989 ;
  assign n29032 = ~n6730 & ~n6761 ;
  assign n29033 = ~n6730 & n21658 ;
  assign n29034 = ~n21684 & n29033 ;
  assign n29035 = ~n29032 & ~n29034 ;
  assign n29036 = n21651 & ~n29035 ;
  assign n29037 = ~\pi0166  & ~n29036 ;
  assign n29038 = n27206 & ~n29037 ;
  assign n29039 = n29031 & ~n29038 ;
  assign n29040 = n29030 & n29039 ;
  assign n29041 = ~n27813 & ~n28973 ;
  assign n29042 = ~\pi0215  & n29041 ;
  assign n29043 = ~\pi0166  & ~n21728 ;
  assign n29044 = \pi0215  & ~n29043 ;
  assign n29045 = ~n21724 & n29044 ;
  assign n29046 = \pi0299  & ~n29045 ;
  assign n29047 = ~n29042 & n29046 ;
  assign n29048 = n27821 & n29046 ;
  assign n29049 = n28969 & n29048 ;
  assign n29050 = ~n29047 & ~n29049 ;
  assign n29051 = \pi0772  & n29050 ;
  assign n29052 = ~n29040 & n29051 ;
  assign n29053 = ~n2165 & n28982 ;
  assign n29054 = ~n2165 & ~n26930 ;
  assign n29055 = ~n29026 & n29054 ;
  assign n29056 = ~n29053 & ~n29055 ;
  assign n29057 = ~n21285 & n27796 ;
  assign n29058 = n21285 & n29021 ;
  assign n29059 = ~n29057 & ~n29058 ;
  assign n29060 = ~\pi0223  & ~n27767 ;
  assign n29061 = n29059 & n29060 ;
  assign n29062 = n29056 & n29061 ;
  assign n29063 = ~\pi0299  & ~n29038 ;
  assign n29064 = ~n29062 & n29063 ;
  assign n29065 = ~\pi0299  & ~\pi0772  ;
  assign n29066 = ~\pi0772  & n27843 ;
  assign n29067 = n29045 & n29066 ;
  assign n29068 = ~n29065 & ~n29067 ;
  assign n29069 = n27736 & n28969 ;
  assign n29070 = ~\pi0215  & ~\pi0772  ;
  assign n29071 = ~n27128 & n29070 ;
  assign n29072 = n29041 & n29071 ;
  assign n29073 = ~n29069 & n29072 ;
  assign n29074 = n29068 & ~n29073 ;
  assign n29075 = ~n29064 & ~n29074 ;
  assign n29076 = ~n29052 & ~n29075 ;
  assign n29077 = \pi0039  & ~n29018 ;
  assign n29078 = n29076 & n29077 ;
  assign n29079 = ~n29019 & ~n29078 ;
  assign n29080 = \pi0727  & n29010 ;
  assign n29081 = ~n29079 & n29080 ;
  assign n29082 = ~n29011 & ~n29081 ;
  assign n29083 = ~n28943 & n29082 ;
  assign n29084 = \pi0167  & ~n27085 ;
  assign n29085 = ~n27069 & n29084 ;
  assign n29086 = ~n27061 & n29085 ;
  assign n29087 = ~\pi0038  & ~n29086 ;
  assign n29088 = ~\pi0167  & ~n21757 ;
  assign n29089 = n27096 & ~n29088 ;
  assign n29090 = \pi0768  & ~n29089 ;
  assign n29091 = ~n29087 & n29090 ;
  assign n29092 = ~\pi0167  & \pi0768  ;
  assign n29093 = ~n29089 & n29092 ;
  assign n29094 = n27107 & n29093 ;
  assign n29095 = n27137 & n29093 ;
  assign n29096 = ~n27132 & n29095 ;
  assign n29097 = ~n29094 & ~n29096 ;
  assign n29098 = ~n29091 & n29097 ;
  assign n29099 = \pi0705  & ~n29098 ;
  assign n29100 = ~\pi0167  & ~n27223 ;
  assign n29101 = ~n27216 & n29100 ;
  assign n29102 = \pi0167  & ~n27173 ;
  assign n29103 = ~n27167 & n29102 ;
  assign n29104 = ~n27159 & n29103 ;
  assign n29105 = ~\pi0038  & ~n29104 ;
  assign n29106 = ~n29101 & n29105 ;
  assign n29107 = ~\pi0768  & ~n27990 ;
  assign n29108 = ~\pi0167  & ~\pi0768  ;
  assign n29109 = ~n27144 & n29108 ;
  assign n29110 = ~n29107 & ~n29109 ;
  assign n29111 = \pi0705  & ~n29110 ;
  assign n29112 = ~n29106 & n29111 ;
  assign n29113 = ~n29099 & ~n29112 ;
  assign n29114 = ~\pi0167  & ~n11834 ;
  assign n29115 = ~\pi0832  & ~n29114 ;
  assign n29116 = ~\pi0768  & n28033 ;
  assign n29117 = \pi0038  & \pi0167  ;
  assign n29118 = ~\pi0768  & n29117 ;
  assign n29119 = ~n22123 & n29118 ;
  assign n29120 = ~n29116 & ~n29119 ;
  assign n29121 = n27268 & n29108 ;
  assign n29122 = n29120 & ~n29121 ;
  assign n29123 = \pi0768  & ~n22124 ;
  assign n29124 = ~n28084 & n29123 ;
  assign n29125 = ~\pi0768  & ~n27305 ;
  assign n29126 = ~n27292 & n29125 ;
  assign n29127 = ~n27286 & n29126 ;
  assign n29128 = \pi0038  & ~\pi0768  ;
  assign n29129 = \pi0167  & ~n29128 ;
  assign n29130 = ~n29127 & n29129 ;
  assign n29131 = ~\pi0705  & ~n29130 ;
  assign n29132 = ~n29124 & n29131 ;
  assign n29133 = n29122 & n29132 ;
  assign n29134 = n29115 & ~n29133 ;
  assign n29135 = n29113 & n29134 ;
  assign n29136 = ~\pi0768  & \pi0947  ;
  assign n29137 = \pi0705  & n26930 ;
  assign n29138 = ~n29136 & ~n29137 ;
  assign n29139 = n1689 & ~n29138 ;
  assign n29140 = ~\pi0167  & ~n1689 ;
  assign n29141 = \pi0832  & ~n29140 ;
  assign n29142 = ~n29139 & n29141 ;
  assign n29143 = \pi0167  & ~\pi0832  ;
  assign n29144 = ~n11834 & n29143 ;
  assign n29145 = ~n29142 & ~n29144 ;
  assign n29146 = ~n29135 & n29145 ;
  assign n29147 = \pi0699  & n26930 ;
  assign n29148 = \pi0763  & \pi0947  ;
  assign n29149 = n1689 & ~n29148 ;
  assign n29150 = ~n29147 & n29149 ;
  assign n29151 = \pi0168  & ~n1689 ;
  assign n29152 = \pi0832  & ~n29151 ;
  assign n29153 = ~n29150 & n29152 ;
  assign n29154 = \pi0057  & \pi0168  ;
  assign n29155 = ~\pi0832  & ~n29154 ;
  assign n29156 = ~\pi0057  & \pi0168  ;
  assign n29157 = ~n27409 & ~n29156 ;
  assign n29158 = \pi0168  & ~\pi0699  ;
  assign n29159 = ~n22123 & n29158 ;
  assign n29160 = \pi0699  & n27402 ;
  assign n29161 = n1354 & ~n29148 ;
  assign n29162 = n21755 & n29161 ;
  assign n29163 = n1358 & n29162 ;
  assign n29164 = n27879 & ~n29163 ;
  assign n29165 = ~n29160 & ~n29164 ;
  assign n29166 = ~n29159 & ~n29165 ;
  assign n29167 = ~\pi0168  & ~n21692 ;
  assign n29168 = n27361 & ~n29167 ;
  assign n29169 = \pi0168  & ~n21728 ;
  assign n29170 = n27259 & ~n29169 ;
  assign n29171 = ~n21724 & n29170 ;
  assign n29172 = \pi0299  & ~n29171 ;
  assign n29173 = \pi0763  & ~n29172 ;
  assign n29174 = \pi0168  & ~n2352 ;
  assign n29175 = n27627 & n29174 ;
  assign n29176 = \pi0168  & n2352 ;
  assign n29177 = n21285 & n29176 ;
  assign n29178 = ~n27256 & ~n29177 ;
  assign n29179 = \pi0763  & n29178 ;
  assign n29180 = ~n29175 & n29179 ;
  assign n29181 = n27899 & n29180 ;
  assign n29182 = ~n27891 & n29181 ;
  assign n29183 = ~n29173 & ~n29182 ;
  assign n29184 = ~n29168 & ~n29183 ;
  assign n29185 = ~\pi0168  & ~\pi0763  ;
  assign n29186 = ~\pi0299  & n29185 ;
  assign n29187 = ~n21692 & n29186 ;
  assign n29188 = \pi0039  & ~n29185 ;
  assign n29189 = ~n21733 & ~n29188 ;
  assign n29190 = ~n29187 & ~n29189 ;
  assign n29191 = ~n29184 & n29190 ;
  assign n29192 = ~\pi0763  & ~n21743 ;
  assign n29193 = ~n27292 & ~n29192 ;
  assign n29194 = ~\pi0168  & ~n27219 ;
  assign n29195 = ~n27217 & n29194 ;
  assign n29196 = ~n29193 & ~n29195 ;
  assign n29197 = n27916 & ~n29196 ;
  assign n29198 = ~n29191 & n29197 ;
  assign n29199 = ~n29166 & ~n29198 ;
  assign n29200 = ~n29157 & n29199 ;
  assign n29201 = n27068 & ~n29195 ;
  assign n29202 = ~n29193 & n29201 ;
  assign n29203 = ~\pi0038  & ~n29202 ;
  assign n29204 = \pi0168  & ~n27158 ;
  assign n29205 = n27672 & ~n29204 ;
  assign n29206 = ~\pi0299  & \pi0763  ;
  assign n29207 = ~n27813 & ~n29177 ;
  assign n29208 = ~\pi0215  & n29207 ;
  assign n29209 = ~n29175 & n29208 ;
  assign n29210 = ~n21698 & n29209 ;
  assign n29211 = n21694 & n29209 ;
  assign n29212 = ~n21711 & n29211 ;
  assign n29213 = ~n29210 & ~n29212 ;
  assign n29214 = \pi0215  & ~n29169 ;
  assign n29215 = ~n21724 & n29214 ;
  assign n29216 = \pi0763  & ~n29215 ;
  assign n29217 = n29213 & n29216 ;
  assign n29218 = ~n29206 & ~n29217 ;
  assign n29219 = ~n29205 & ~n29218 ;
  assign n29220 = \pi0039  & n29219 ;
  assign n29221 = ~n27128 & ~n29177 ;
  assign n29222 = ~n29175 & n29221 ;
  assign n29223 = ~n27122 & n29222 ;
  assign n29224 = ~n27891 & n29223 ;
  assign n29225 = n21948 & ~n29224 ;
  assign n29226 = n27523 & ~n29167 ;
  assign n29227 = \pi0168  & \pi0215  ;
  assign n29228 = ~n21728 & n29227 ;
  assign n29229 = ~n27299 & ~n29228 ;
  assign n29230 = ~n27947 & n29229 ;
  assign n29231 = \pi0299  & ~n29230 ;
  assign n29232 = ~n29226 & ~n29231 ;
  assign n29233 = ~n29225 & n29232 ;
  assign n29234 = \pi0039  & ~\pi0763  ;
  assign n29235 = ~n29233 & n29234 ;
  assign n29236 = ~n29220 & ~n29235 ;
  assign n29237 = n29203 & n29236 ;
  assign n29238 = ~n26930 & n29163 ;
  assign n29239 = \pi0168  & ~n21757 ;
  assign n29240 = \pi0038  & ~n29239 ;
  assign n29241 = ~n29238 & n29240 ;
  assign n29242 = \pi0699  & ~n29241 ;
  assign n29243 = ~n29157 & n29242 ;
  assign n29244 = ~n29237 & n29243 ;
  assign n29245 = ~n29200 & ~n29244 ;
  assign n29246 = n29155 & n29245 ;
  assign n29247 = ~n29153 & ~n29246 ;
  assign n29248 = \pi0729  & n26930 ;
  assign n29249 = \pi0746  & \pi0947  ;
  assign n29250 = n1689 & ~n29249 ;
  assign n29251 = ~n29248 & n29250 ;
  assign n29252 = \pi0169  & ~n1689 ;
  assign n29253 = \pi0832  & ~n29252 ;
  assign n29254 = ~n29251 & n29253 ;
  assign n29255 = \pi0057  & \pi0169  ;
  assign n29256 = ~\pi0832  & ~n29255 ;
  assign n29257 = ~\pi0057  & \pi0169  ;
  assign n29258 = ~n27409 & ~n29257 ;
  assign n29259 = \pi0169  & ~\pi0729  ;
  assign n29260 = ~n22123 & n29259 ;
  assign n29261 = \pi0729  & n27402 ;
  assign n29262 = n1354 & ~n29249 ;
  assign n29263 = n21755 & n29262 ;
  assign n29264 = n1358 & n29263 ;
  assign n29265 = n27879 & ~n29264 ;
  assign n29266 = ~n29261 & ~n29265 ;
  assign n29267 = ~n29260 & ~n29266 ;
  assign n29268 = ~\pi0169  & ~n21692 ;
  assign n29269 = n27361 & ~n29268 ;
  assign n29270 = \pi0169  & ~n21728 ;
  assign n29271 = n27259 & ~n29270 ;
  assign n29272 = ~n21724 & n29271 ;
  assign n29273 = \pi0299  & ~n29272 ;
  assign n29274 = \pi0746  & ~n29273 ;
  assign n29275 = \pi0169  & ~n2352 ;
  assign n29276 = n27627 & n29275 ;
  assign n29277 = \pi0169  & n2352 ;
  assign n29278 = n21285 & n29277 ;
  assign n29279 = ~n27256 & ~n29278 ;
  assign n29280 = \pi0746  & n29279 ;
  assign n29281 = ~n29276 & n29280 ;
  assign n29282 = n27899 & n29281 ;
  assign n29283 = ~n27891 & n29282 ;
  assign n29284 = ~n29274 & ~n29283 ;
  assign n29285 = ~n29269 & ~n29284 ;
  assign n29286 = ~\pi0169  & ~\pi0746  ;
  assign n29287 = ~\pi0299  & n29286 ;
  assign n29288 = ~n21692 & n29287 ;
  assign n29289 = \pi0039  & ~n29286 ;
  assign n29290 = ~n21733 & ~n29289 ;
  assign n29291 = ~n29288 & ~n29290 ;
  assign n29292 = ~n29285 & n29291 ;
  assign n29293 = ~\pi0746  & ~n21743 ;
  assign n29294 = ~n27292 & ~n29293 ;
  assign n29295 = ~\pi0169  & ~n27219 ;
  assign n29296 = ~n27217 & n29295 ;
  assign n29297 = ~n29294 & ~n29296 ;
  assign n29298 = n27916 & ~n29297 ;
  assign n29299 = ~n29292 & n29298 ;
  assign n29300 = ~n29267 & ~n29299 ;
  assign n29301 = ~n29258 & n29300 ;
  assign n29302 = n27068 & ~n29296 ;
  assign n29303 = ~n29294 & n29302 ;
  assign n29304 = ~\pi0038  & ~n29303 ;
  assign n29305 = \pi0169  & ~n27158 ;
  assign n29306 = n27672 & ~n29305 ;
  assign n29307 = ~\pi0299  & \pi0746  ;
  assign n29308 = ~n27813 & ~n29278 ;
  assign n29309 = ~\pi0215  & n29308 ;
  assign n29310 = ~n29276 & n29309 ;
  assign n29311 = ~n21698 & n29310 ;
  assign n29312 = n21694 & n29310 ;
  assign n29313 = ~n21711 & n29312 ;
  assign n29314 = ~n29311 & ~n29313 ;
  assign n29315 = \pi0215  & ~n29270 ;
  assign n29316 = ~n21724 & n29315 ;
  assign n29317 = \pi0746  & ~n29316 ;
  assign n29318 = n29314 & n29317 ;
  assign n29319 = ~n29307 & ~n29318 ;
  assign n29320 = ~n29306 & ~n29319 ;
  assign n29321 = \pi0039  & n29320 ;
  assign n29322 = ~n27128 & ~n29278 ;
  assign n29323 = ~n29276 & n29322 ;
  assign n29324 = ~n27122 & n29323 ;
  assign n29325 = ~n27891 & n29324 ;
  assign n29326 = n21948 & ~n29325 ;
  assign n29327 = n27523 & ~n29268 ;
  assign n29328 = \pi0169  & \pi0215  ;
  assign n29329 = ~n21728 & n29328 ;
  assign n29330 = ~n27299 & ~n29329 ;
  assign n29331 = ~n27947 & n29330 ;
  assign n29332 = \pi0299  & ~n29331 ;
  assign n29333 = ~n29327 & ~n29332 ;
  assign n29334 = ~n29326 & n29333 ;
  assign n29335 = \pi0039  & ~\pi0746  ;
  assign n29336 = ~n29334 & n29335 ;
  assign n29337 = ~n29321 & ~n29336 ;
  assign n29338 = n29304 & n29337 ;
  assign n29339 = ~n26930 & n29264 ;
  assign n29340 = \pi0169  & ~n21757 ;
  assign n29341 = \pi0038  & ~n29340 ;
  assign n29342 = ~n29339 & n29341 ;
  assign n29343 = \pi0729  & ~n29342 ;
  assign n29344 = ~n29258 & n29343 ;
  assign n29345 = ~n29338 & n29344 ;
  assign n29346 = ~n29301 & ~n29345 ;
  assign n29347 = n29256 & n29346 ;
  assign n29348 = ~n29254 & ~n29347 ;
  assign n29349 = \pi0730  & n26930 ;
  assign n29350 = \pi0748  & \pi0947  ;
  assign n29351 = n1689 & ~n29350 ;
  assign n29352 = ~n29349 & n29351 ;
  assign n29353 = \pi0170  & ~n1689 ;
  assign n29354 = \pi0832  & ~n29353 ;
  assign n29355 = ~n29352 & n29354 ;
  assign n29356 = \pi0057  & \pi0170  ;
  assign n29357 = ~\pi0832  & ~n29356 ;
  assign n29358 = ~n29355 & ~n29357 ;
  assign n29359 = ~\pi0170  & ~n27219 ;
  assign n29360 = ~n27217 & n29359 ;
  assign n29361 = n1288 & n27068 ;
  assign n29362 = ~n29360 & n29361 ;
  assign n29363 = ~n9627 & ~n29362 ;
  assign n29364 = \pi0170  & \pi0215  ;
  assign n29365 = ~n21728 & n29364 ;
  assign n29366 = ~n27299 & ~n29365 ;
  assign n29367 = ~n27947 & n29366 ;
  assign n29368 = \pi0299  & ~n29367 ;
  assign n29369 = ~\pi0170  & ~n21692 ;
  assign n29370 = n27523 & ~n29369 ;
  assign n29371 = ~n29368 & ~n29370 ;
  assign n29372 = \pi0170  & ~n2352 ;
  assign n29373 = n27627 & n29372 ;
  assign n29374 = \pi0170  & n2352 ;
  assign n29375 = n21285 & n29374 ;
  assign n29376 = ~n27128 & ~n29375 ;
  assign n29377 = ~n29373 & n29376 ;
  assign n29378 = ~n27122 & n29377 ;
  assign n29379 = ~n27891 & n29378 ;
  assign n29380 = n21948 & ~n29379 ;
  assign n29381 = ~n29362 & ~n29380 ;
  assign n29382 = n29371 & n29381 ;
  assign n29383 = ~n29363 & ~n29382 ;
  assign n29384 = ~\pi0170  & ~n21757 ;
  assign n29385 = n27096 & ~n29384 ;
  assign n29386 = ~\pi0748  & ~n29385 ;
  assign n29387 = ~n29383 & n29386 ;
  assign n29388 = n27990 & ~n29384 ;
  assign n29389 = \pi0748  & ~n29388 ;
  assign n29390 = \pi0730  & ~n29389 ;
  assign n29391 = \pi0170  & ~n27158 ;
  assign n29392 = n27167 & ~n29360 ;
  assign n29393 = ~n29391 & ~n29392 ;
  assign n29394 = n27672 & n29393 ;
  assign n29395 = ~n27813 & ~n29375 ;
  assign n29396 = ~\pi0215  & n29395 ;
  assign n29397 = ~n29373 & n29396 ;
  assign n29398 = ~n21698 & n29397 ;
  assign n29399 = n21694 & n29397 ;
  assign n29400 = ~n21711 & n29399 ;
  assign n29401 = ~n29398 & ~n29400 ;
  assign n29402 = \pi0170  & ~n21728 ;
  assign n29403 = \pi0215  & ~n29402 ;
  assign n29404 = ~n21724 & n29403 ;
  assign n29405 = \pi0039  & ~n29404 ;
  assign n29406 = n29401 & n29405 ;
  assign n29407 = ~n6205 & ~n29406 ;
  assign n29408 = ~n29392 & n29407 ;
  assign n29409 = ~\pi0038  & \pi0730  ;
  assign n29410 = ~n29408 & n29409 ;
  assign n29411 = ~n29394 & n29410 ;
  assign n29412 = ~n29390 & ~n29411 ;
  assign n29413 = ~n29387 & ~n29412 ;
  assign n29414 = ~\pi0170  & ~\pi0748  ;
  assign n29415 = n21770 & n29414 ;
  assign n29416 = ~n21734 & n29415 ;
  assign n29417 = \pi0038  & n29414 ;
  assign n29418 = ~n22123 & n29417 ;
  assign n29419 = ~\pi0730  & ~n29418 ;
  assign n29420 = ~n29416 & n29419 ;
  assign n29421 = ~n27256 & ~n29375 ;
  assign n29422 = ~n29373 & n29421 ;
  assign n29423 = n27899 & n29422 ;
  assign n29424 = ~n27891 & n29423 ;
  assign n29425 = n27259 & ~n29402 ;
  assign n29426 = ~n21724 & n29425 ;
  assign n29427 = \pi0299  & ~n29426 ;
  assign n29428 = ~n29424 & n29427 ;
  assign n29429 = n27361 & ~n29369 ;
  assign n29430 = ~n29428 & ~n29429 ;
  assign n29431 = n9627 & ~n29430 ;
  assign n29432 = n1288 & n27291 ;
  assign n29433 = ~n29360 & n29432 ;
  assign n29434 = \pi0038  & \pi0170  ;
  assign n29435 = \pi0748  & ~n29434 ;
  assign n29436 = \pi0748  & n21765 ;
  assign n29437 = n1638 & n29436 ;
  assign n29438 = ~n29435 & ~n29437 ;
  assign n29439 = ~n28033 & ~n29438 ;
  assign n29440 = ~n29433 & n29439 ;
  assign n29441 = ~n29431 & n29440 ;
  assign n29442 = n29420 & ~n29441 ;
  assign n29443 = n27402 & ~n29442 ;
  assign n29444 = ~n29413 & n29443 ;
  assign n29445 = ~\pi0057  & \pi0170  ;
  assign n29446 = ~n27409 & ~n29445 ;
  assign n29447 = ~n29355 & ~n29446 ;
  assign n29448 = ~n29444 & n29447 ;
  assign n29449 = ~n29358 & ~n29448 ;
  assign n29450 = \pi0691  & n26930 ;
  assign n29451 = \pi0764  & \pi0947  ;
  assign n29452 = n1689 & ~n29451 ;
  assign n29453 = ~n29450 & n29452 ;
  assign n29454 = \pi0171  & ~n1689 ;
  assign n29455 = \pi0832  & ~n29454 ;
  assign n29456 = ~n29453 & n29455 ;
  assign n29457 = \pi0057  & \pi0171  ;
  assign n29458 = ~\pi0832  & ~n29457 ;
  assign n29459 = ~\pi0057  & \pi0171  ;
  assign n29460 = ~n27409 & ~n29459 ;
  assign n29461 = \pi0171  & ~\pi0691  ;
  assign n29462 = ~n22123 & n29461 ;
  assign n29463 = \pi0691  & n27402 ;
  assign n29464 = n1354 & ~n29451 ;
  assign n29465 = n21755 & n29464 ;
  assign n29466 = n1358 & n29465 ;
  assign n29467 = n27879 & ~n29466 ;
  assign n29468 = ~n29463 & ~n29467 ;
  assign n29469 = ~n29462 & ~n29468 ;
  assign n29470 = ~\pi0171  & ~n21692 ;
  assign n29471 = n27361 & ~n29470 ;
  assign n29472 = \pi0171  & ~n21728 ;
  assign n29473 = n27259 & ~n29472 ;
  assign n29474 = ~n21724 & n29473 ;
  assign n29475 = \pi0299  & ~n29474 ;
  assign n29476 = \pi0764  & ~n29475 ;
  assign n29477 = \pi0171  & ~n2352 ;
  assign n29478 = n27627 & n29477 ;
  assign n29479 = \pi0171  & n2352 ;
  assign n29480 = n21285 & n29479 ;
  assign n29481 = ~n27256 & ~n29480 ;
  assign n29482 = \pi0764  & n29481 ;
  assign n29483 = ~n29478 & n29482 ;
  assign n29484 = n27899 & n29483 ;
  assign n29485 = ~n27891 & n29484 ;
  assign n29486 = ~n29476 & ~n29485 ;
  assign n29487 = ~n29471 & ~n29486 ;
  assign n29488 = ~\pi0171  & ~\pi0764  ;
  assign n29489 = ~\pi0299  & n29488 ;
  assign n29490 = ~n21692 & n29489 ;
  assign n29491 = \pi0039  & ~n29488 ;
  assign n29492 = ~n21733 & ~n29491 ;
  assign n29493 = ~n29490 & ~n29492 ;
  assign n29494 = ~n29487 & n29493 ;
  assign n29495 = ~\pi0764  & ~n21743 ;
  assign n29496 = ~n27292 & ~n29495 ;
  assign n29497 = ~\pi0171  & ~n27219 ;
  assign n29498 = ~n27217 & n29497 ;
  assign n29499 = ~n29496 & ~n29498 ;
  assign n29500 = n27916 & ~n29499 ;
  assign n29501 = ~n29494 & n29500 ;
  assign n29502 = ~n29469 & ~n29501 ;
  assign n29503 = ~n29460 & n29502 ;
  assign n29504 = n27068 & ~n29498 ;
  assign n29505 = ~n29496 & n29504 ;
  assign n29506 = ~\pi0038  & ~n29505 ;
  assign n29507 = \pi0171  & ~n27158 ;
  assign n29508 = n27672 & ~n29507 ;
  assign n29509 = ~\pi0299  & \pi0764  ;
  assign n29510 = ~n27813 & ~n29480 ;
  assign n29511 = ~\pi0215  & n29510 ;
  assign n29512 = ~n29478 & n29511 ;
  assign n29513 = ~n21698 & n29512 ;
  assign n29514 = n21694 & n29512 ;
  assign n29515 = ~n21711 & n29514 ;
  assign n29516 = ~n29513 & ~n29515 ;
  assign n29517 = \pi0215  & ~n29472 ;
  assign n29518 = ~n21724 & n29517 ;
  assign n29519 = \pi0764  & ~n29518 ;
  assign n29520 = n29516 & n29519 ;
  assign n29521 = ~n29509 & ~n29520 ;
  assign n29522 = ~n29508 & ~n29521 ;
  assign n29523 = \pi0039  & n29522 ;
  assign n29524 = ~n27128 & ~n29480 ;
  assign n29525 = ~n29478 & n29524 ;
  assign n29526 = ~n27122 & n29525 ;
  assign n29527 = ~n27891 & n29526 ;
  assign n29528 = n21948 & ~n29527 ;
  assign n29529 = n27523 & ~n29470 ;
  assign n29530 = \pi0171  & \pi0215  ;
  assign n29531 = ~n21728 & n29530 ;
  assign n29532 = ~n27299 & ~n29531 ;
  assign n29533 = ~n27947 & n29532 ;
  assign n29534 = \pi0299  & ~n29533 ;
  assign n29535 = ~n29529 & ~n29534 ;
  assign n29536 = ~n29528 & n29535 ;
  assign n29537 = \pi0039  & ~\pi0764  ;
  assign n29538 = ~n29536 & n29537 ;
  assign n29539 = ~n29523 & ~n29538 ;
  assign n29540 = n29506 & n29539 ;
  assign n29541 = ~n26930 & n29466 ;
  assign n29542 = \pi0171  & ~n21757 ;
  assign n29543 = \pi0038  & ~n29542 ;
  assign n29544 = ~n29541 & n29543 ;
  assign n29545 = \pi0691  & ~n29544 ;
  assign n29546 = ~n29460 & n29545 ;
  assign n29547 = ~n29540 & n29546 ;
  assign n29548 = ~n29503 & ~n29547 ;
  assign n29549 = n29458 & n29548 ;
  assign n29550 = ~n29456 & ~n29549 ;
  assign n29551 = \pi0690  & n26930 ;
  assign n29552 = \pi0739  & \pi0947  ;
  assign n29553 = n1689 & ~n29552 ;
  assign n29554 = ~n29551 & n29553 ;
  assign n29555 = \pi0172  & ~n1689 ;
  assign n29556 = \pi0832  & ~n29555 ;
  assign n29557 = ~n29554 & n29556 ;
  assign n29558 = \pi0057  & \pi0172  ;
  assign n29559 = ~\pi0832  & ~n29558 ;
  assign n29560 = ~\pi0057  & \pi0172  ;
  assign n29561 = ~n27409 & ~n29560 ;
  assign n29562 = \pi0172  & ~\pi0690  ;
  assign n29563 = ~n22123 & n29562 ;
  assign n29564 = \pi0690  & n27402 ;
  assign n29565 = n1354 & ~n29552 ;
  assign n29566 = n21755 & n29565 ;
  assign n29567 = n1358 & n29566 ;
  assign n29568 = n27879 & ~n29567 ;
  assign n29569 = ~n29564 & ~n29568 ;
  assign n29570 = ~n29563 & ~n29569 ;
  assign n29571 = ~\pi0172  & ~n21692 ;
  assign n29572 = n27361 & ~n29571 ;
  assign n29573 = \pi0172  & ~n21728 ;
  assign n29574 = n27259 & ~n29573 ;
  assign n29575 = ~n21724 & n29574 ;
  assign n29576 = \pi0299  & ~n29575 ;
  assign n29577 = \pi0739  & ~n29576 ;
  assign n29578 = \pi0172  & ~n2352 ;
  assign n29579 = n27627 & n29578 ;
  assign n29580 = \pi0172  & n2352 ;
  assign n29581 = n21285 & n29580 ;
  assign n29582 = ~n27256 & ~n29581 ;
  assign n29583 = \pi0739  & n29582 ;
  assign n29584 = ~n29579 & n29583 ;
  assign n29585 = n27899 & n29584 ;
  assign n29586 = ~n27891 & n29585 ;
  assign n29587 = ~n29577 & ~n29586 ;
  assign n29588 = ~n29572 & ~n29587 ;
  assign n29589 = ~\pi0172  & ~\pi0739  ;
  assign n29590 = ~\pi0299  & n29589 ;
  assign n29591 = ~n21692 & n29590 ;
  assign n29592 = \pi0039  & ~n29589 ;
  assign n29593 = ~n21733 & ~n29592 ;
  assign n29594 = ~n29591 & ~n29593 ;
  assign n29595 = ~n29588 & n29594 ;
  assign n29596 = ~\pi0172  & ~n27328 ;
  assign n29597 = ~\pi0172  & \pi0299  ;
  assign n29598 = n21205 & n29597 ;
  assign n29599 = n21237 & n29597 ;
  assign n29600 = n21232 & n29599 ;
  assign n29601 = ~n29598 & ~n29600 ;
  assign n29602 = ~\pi0039  & n29601 ;
  assign n29603 = ~n29596 & n29602 ;
  assign n29604 = \pi0299  & n29552 ;
  assign n29605 = ~n21205 & n29604 ;
  assign n29606 = ~n21238 & n29605 ;
  assign n29607 = ~\pi0299  & n29552 ;
  assign n29608 = ~n21740 & n29607 ;
  assign n29609 = ~n21738 & n29608 ;
  assign n29610 = ~n29606 & ~n29609 ;
  assign n29611 = n29603 & n29610 ;
  assign n29612 = n27916 & ~n29611 ;
  assign n29613 = ~n29595 & n29612 ;
  assign n29614 = ~n29570 & ~n29613 ;
  assign n29615 = ~n29561 & n29614 ;
  assign n29616 = n27068 & n29610 ;
  assign n29617 = n29603 & n29616 ;
  assign n29618 = ~\pi0038  & ~n29617 ;
  assign n29619 = \pi0172  & \pi0215  ;
  assign n29620 = ~n21728 & n29619 ;
  assign n29621 = ~n27299 & ~n29620 ;
  assign n29622 = ~n27947 & n29621 ;
  assign n29623 = \pi0299  & ~n29622 ;
  assign n29624 = ~n27128 & ~n29581 ;
  assign n29625 = ~n29579 & n29624 ;
  assign n29626 = ~n27122 & n29625 ;
  assign n29627 = ~n27891 & n29626 ;
  assign n29628 = n21948 & ~n29627 ;
  assign n29629 = ~n29623 & ~n29628 ;
  assign n29630 = n27523 & ~n29571 ;
  assign n29631 = ~\pi0739  & ~n29630 ;
  assign n29632 = n29629 & n29631 ;
  assign n29633 = \pi0172  & ~n27158 ;
  assign n29634 = \pi0739  & ~n29633 ;
  assign n29635 = n27672 & n29634 ;
  assign n29636 = \pi0215  & ~n29573 ;
  assign n29637 = ~n21724 & n29636 ;
  assign n29638 = ~n27813 & ~n29581 ;
  assign n29639 = ~\pi0215  & n29638 ;
  assign n29640 = ~n29579 & n29639 ;
  assign n29641 = ~n21698 & n29640 ;
  assign n29642 = n21694 & n29640 ;
  assign n29643 = ~n21711 & n29642 ;
  assign n29644 = ~n29641 & ~n29643 ;
  assign n29645 = ~n29637 & n29644 ;
  assign n29646 = \pi0299  & \pi0739  ;
  assign n29647 = ~n29645 & n29646 ;
  assign n29648 = \pi0039  & ~n29647 ;
  assign n29649 = ~n29635 & n29648 ;
  assign n29650 = ~n29632 & n29649 ;
  assign n29651 = n29618 & ~n29650 ;
  assign n29652 = ~n26930 & n29567 ;
  assign n29653 = \pi0172  & ~n21757 ;
  assign n29654 = \pi0038  & ~n29653 ;
  assign n29655 = ~n29652 & n29654 ;
  assign n29656 = \pi0690  & ~n29655 ;
  assign n29657 = ~n29561 & n29656 ;
  assign n29658 = ~n29651 & n29657 ;
  assign n29659 = ~n29615 & ~n29658 ;
  assign n29660 = n29559 & n29659 ;
  assign n29661 = ~n29557 & ~n29660 ;
  assign n29662 = \pi0173  & ~\pi0832  ;
  assign n29663 = ~n21132 & ~n29662 ;
  assign n29664 = ~\pi0173  & \pi0788  ;
  assign n29665 = ~n1689 & n29664 ;
  assign n29666 = ~n20778 & n29665 ;
  assign n29667 = ~\pi0745  & n1689 ;
  assign n29668 = n20784 & n29667 ;
  assign n29669 = n22767 & n29668 ;
  assign n29670 = ~\pi0173  & ~n1689 ;
  assign n29671 = ~n29668 & ~n29670 ;
  assign n29672 = ~n20792 & ~n29671 ;
  assign n29673 = ~n29669 & n29672 ;
  assign n29674 = n20801 & ~n29673 ;
  assign n29675 = ~\pi1155  & ~n29670 ;
  assign n29676 = \pi0785  & n29675 ;
  assign n29677 = ~n29669 & n29676 ;
  assign n29678 = ~\pi0785  & ~n29670 ;
  assign n29679 = ~n29668 & n29678 ;
  assign n29680 = ~n20804 & ~n29679 ;
  assign n29681 = n20877 & ~n21032 ;
  assign n29682 = ~n20812 & ~n29681 ;
  assign n29683 = n29680 & n29682 ;
  assign n29684 = ~n29677 & n29683 ;
  assign n29685 = ~n29674 & n29684 ;
  assign n29686 = n20816 & n29685 ;
  assign n29687 = ~n29666 & ~n29686 ;
  assign n29688 = ~\pi0788  & n29685 ;
  assign n29689 = ~\pi0723  & n1689 ;
  assign n29690 = n20855 & n29689 ;
  assign n29691 = ~n29670 & ~n29690 ;
  assign n29692 = ~\pi0778  & ~n29691 ;
  assign n29693 = ~\pi0625  & ~\pi0723  ;
  assign n29694 = n1689 & n29693 ;
  assign n29695 = n20855 & n29694 ;
  assign n29696 = \pi1153  & n29695 ;
  assign n29697 = \pi1153  & ~n29670 ;
  assign n29698 = ~n29690 & n29697 ;
  assign n29699 = ~n29696 & ~n29698 ;
  assign n29700 = ~\pi1153  & ~n29670 ;
  assign n29701 = ~n29695 & n29700 ;
  assign n29702 = \pi0778  & ~n29701 ;
  assign n29703 = n29699 & n29702 ;
  assign n29704 = ~n29692 & ~n29703 ;
  assign n29705 = n26485 & ~n29704 ;
  assign n29706 = ~\pi0629  & ~n29705 ;
  assign n29707 = ~n29688 & n29706 ;
  assign n29708 = n29687 & n29707 ;
  assign n29709 = ~\pi0629  & ~n20887 ;
  assign n29710 = ~n29705 & n29709 ;
  assign n29711 = \pi0792  & ~n29710 ;
  assign n29712 = ~n29708 & n29711 ;
  assign n29713 = n26474 & ~n29704 ;
  assign n29714 = \pi0629  & ~n20886 ;
  assign n29715 = ~n29713 & n29714 ;
  assign n29716 = \pi0629  & ~n29713 ;
  assign n29717 = ~n29688 & n29716 ;
  assign n29718 = n29687 & n29717 ;
  assign n29719 = ~n29715 & ~n29718 ;
  assign n29720 = n29712 & n29719 ;
  assign n29721 = ~n21067 & ~n29720 ;
  assign n29722 = ~\pi0787  & ~n24761 ;
  assign n29723 = ~\pi0173  & \pi0792  ;
  assign n29724 = ~n1689 & n29723 ;
  assign n29725 = ~n20845 & n29724 ;
  assign n29726 = ~n20910 & ~n29725 ;
  assign n29727 = n20846 & n29726 ;
  assign n29728 = ~n29688 & n29726 ;
  assign n29729 = n29687 & n29728 ;
  assign n29730 = ~n29727 & ~n29729 ;
  assign n29731 = n20850 & ~n29670 ;
  assign n29732 = n26333 & ~n29704 ;
  assign n29733 = n20852 & ~n29732 ;
  assign n29734 = ~n29731 & ~n29733 ;
  assign n29735 = n26319 & ~n29704 ;
  assign n29736 = ~\pi0173  & \pi0647  ;
  assign n29737 = ~n1689 & n29736 ;
  assign n29738 = n20897 & ~n29737 ;
  assign n29739 = ~n29735 & n29738 ;
  assign n29740 = ~n24761 & ~n29739 ;
  assign n29741 = n29734 & n29740 ;
  assign n29742 = n29730 & n29741 ;
  assign n29743 = ~n29722 & ~n29742 ;
  assign n29744 = ~n29721 & ~n29743 ;
  assign n29745 = \pi0608  & ~n29701 ;
  assign n29746 = ~n29668 & n29697 ;
  assign n29747 = \pi0778  & ~n29746 ;
  assign n29748 = n26421 & ~n29691 ;
  assign n29749 = ~n29747 & ~n29748 ;
  assign n29750 = n29745 & ~n29749 ;
  assign n29751 = n26147 & ~n29691 ;
  assign n29752 = ~\pi0723  & ~n20784 ;
  assign n29753 = n22113 & n29752 ;
  assign n29754 = n29671 & ~n29753 ;
  assign n29755 = ~n29751 & ~n29754 ;
  assign n29756 = n29700 & ~n29755 ;
  assign n29757 = n26415 & n29699 ;
  assign n29758 = ~n29756 & n29757 ;
  assign n29759 = ~n29750 & ~n29758 ;
  assign n29760 = ~\pi1155  & ~n29692 ;
  assign n29761 = ~n29703 & n29760 ;
  assign n29762 = ~n20999 & ~n29761 ;
  assign n29763 = ~\pi0778  & ~n29754 ;
  assign n29764 = ~n29762 & ~n29763 ;
  assign n29765 = n29759 & n29764 ;
  assign n29766 = \pi0609  & ~\pi1155  ;
  assign n29767 = ~n29692 & n29766 ;
  assign n29768 = ~n29703 & n29767 ;
  assign n29769 = \pi1155  & ~n29673 ;
  assign n29770 = ~\pi0660  & ~n29769 ;
  assign n29771 = ~n29768 & n29770 ;
  assign n29772 = ~n29765 & n29771 ;
  assign n29773 = \pi0785  & ~n29772 ;
  assign n29774 = n1689 & ~n20811 ;
  assign n29775 = n20871 & ~n29774 ;
  assign n29776 = n29680 & n29775 ;
  assign n29777 = ~n29677 & n29776 ;
  assign n29778 = ~n29674 & n29777 ;
  assign n29779 = ~n20868 & n23667 ;
  assign n29780 = ~n29704 & n29779 ;
  assign n29781 = ~n29778 & ~n29780 ;
  assign n29782 = \pi0781  & ~n29781 ;
  assign n29783 = \pi1155  & ~n29692 ;
  assign n29784 = ~n29703 & n29783 ;
  assign n29785 = ~n21774 & ~n29784 ;
  assign n29786 = ~n29763 & ~n29785 ;
  assign n29787 = n29759 & n29786 ;
  assign n29788 = n26121 & ~n29692 ;
  assign n29789 = ~n29703 & n29788 ;
  assign n29790 = \pi0660  & ~n29675 ;
  assign n29791 = \pi0660  & n29668 ;
  assign n29792 = n22767 & n29791 ;
  assign n29793 = ~n29790 & ~n29792 ;
  assign n29794 = ~n29789 & ~n29793 ;
  assign n29795 = ~n29787 & n29794 ;
  assign n29796 = ~n29782 & ~n29795 ;
  assign n29797 = n29773 & n29796 ;
  assign n29798 = ~\pi0785  & ~n29763 ;
  assign n29799 = ~n29750 & n29798 ;
  assign n29800 = ~n29758 & n29799 ;
  assign n29801 = n21022 & ~n29800 ;
  assign n29802 = ~n29782 & ~n29801 ;
  assign n29803 = ~n21034 & ~n21038 ;
  assign n29804 = ~n29802 & n29803 ;
  assign n29805 = ~n29797 & n29804 ;
  assign n29806 = n1689 & ~n21032 ;
  assign n29807 = ~n20876 & ~n29806 ;
  assign n29808 = ~n20812 & n29807 ;
  assign n29809 = n29680 & n29808 ;
  assign n29810 = ~n29677 & n29809 ;
  assign n29811 = ~n29674 & n29810 ;
  assign n29812 = \pi0648  & n20828 ;
  assign n29813 = ~\pi0648  & n21031 ;
  assign n29814 = ~n29812 & ~n29813 ;
  assign n29815 = n20873 & ~n29814 ;
  assign n29816 = ~n29704 & n29815 ;
  assign n29817 = ~n29811 & ~n29816 ;
  assign n29818 = \pi0789  & ~n21038 ;
  assign n29819 = ~n29817 & n29818 ;
  assign n29820 = n20947 & n29685 ;
  assign n29821 = n26458 & ~n29704 ;
  assign n29822 = ~n20778 & n29670 ;
  assign n29823 = ~n20883 & n29822 ;
  assign n29824 = ~n29821 & ~n29823 ;
  assign n29825 = ~n29820 & n29824 ;
  assign n29826 = \pi0788  & ~n29825 ;
  assign n29827 = ~n29819 & ~n29826 ;
  assign n29828 = ~n29805 & n29827 ;
  assign n29829 = ~n23856 & ~n29743 ;
  assign n29830 = ~n29828 & n29829 ;
  assign n29831 = ~n29744 & ~n29830 ;
  assign n29832 = n20923 & ~n29670 ;
  assign n29833 = n20925 & ~n29732 ;
  assign n29834 = ~n29832 & ~n29833 ;
  assign n29835 = ~\pi1157  & ~n29737 ;
  assign n29836 = ~n29735 & n29835 ;
  assign n29837 = n29834 & ~n29836 ;
  assign n29838 = \pi0787  & ~n29837 ;
  assign n29839 = ~\pi0787  & ~n29732 ;
  assign n29840 = \pi0790  & ~n29839 ;
  assign n29841 = n23518 & n29840 ;
  assign n29842 = ~n29838 & n29841 ;
  assign n29843 = ~n23414 & n29670 ;
  assign n29844 = ~n24886 & n29843 ;
  assign n29845 = ~n29688 & ~n29844 ;
  assign n29846 = n29687 & n29845 ;
  assign n29847 = ~n23415 & ~n29670 ;
  assign n29848 = n20846 & ~n29670 ;
  assign n29849 = ~n23414 & ~n29848 ;
  assign n29850 = ~n29847 & n29849 ;
  assign n29851 = \pi0790  & n29850 ;
  assign n29852 = ~n29846 & n29851 ;
  assign n29853 = \pi0832  & ~n29852 ;
  assign n29854 = ~n29842 & n29853 ;
  assign n29855 = n29831 & n29854 ;
  assign n29856 = n29663 & ~n29855 ;
  assign n29857 = n21749 & n29667 ;
  assign n29858 = n1354 & n29857 ;
  assign n29859 = n8413 & n29858 ;
  assign n29860 = n1358 & n29859 ;
  assign n29861 = \pi0038  & ~\pi0173  ;
  assign n29862 = ~n21757 & n29861 ;
  assign n29863 = ~n29860 & ~n29862 ;
  assign n29864 = \pi0038  & n29863 ;
  assign n29865 = ~\pi0173  & ~n21467 ;
  assign n29866 = ~\pi0039  & ~\pi0173  ;
  assign n29867 = n21272 & n29866 ;
  assign n29868 = ~n29865 & ~n29867 ;
  assign n29869 = ~\pi0173  & ~\pi0745  ;
  assign n29870 = ~\pi0745  & ~n21566 ;
  assign n29871 = n21484 & n29870 ;
  assign n29872 = ~n29869 & ~n29871 ;
  assign n29873 = n29868 & ~n29872 ;
  assign n29874 = ~\pi0173  & \pi0745  ;
  assign n29875 = n21743 & n29874 ;
  assign n29876 = ~n21734 & n29875 ;
  assign n29877 = n29863 & ~n29876 ;
  assign n29878 = ~n29873 & n29877 ;
  assign n29879 = ~n29864 & ~n29878 ;
  assign n29880 = \pi0723  & n29879 ;
  assign n29881 = ~\pi0173  & ~\pi0778  ;
  assign n29882 = ~n23622 & ~n29881 ;
  assign n29883 = n29880 & ~n29882 ;
  assign n29884 = ~\pi0173  & n23548 ;
  assign n29885 = ~n26540 & n29884 ;
  assign n29886 = ~\pi0745  & ~n23558 ;
  assign n29887 = n23557 & n29886 ;
  assign n29888 = ~n29869 & ~n29887 ;
  assign n29889 = ~n29885 & ~n29888 ;
  assign n29890 = ~\pi0038  & ~n29889 ;
  assign n29891 = ~\pi0173  & ~n23567 ;
  assign n29892 = n23565 & n29891 ;
  assign n29893 = \pi0745  & n23575 ;
  assign n29894 = n23572 & n29893 ;
  assign n29895 = ~n29874 & ~n29894 ;
  assign n29896 = ~n29892 & ~n29895 ;
  assign n29897 = n6861 & ~n29896 ;
  assign n29898 = n29890 & n29897 ;
  assign n29899 = \pi0173  & \pi0603  ;
  assign n29900 = ~n20783 & n29899 ;
  assign n29901 = n29667 & n29900 ;
  assign n29902 = \pi0173  & ~n20784 ;
  assign n29903 = n22113 & n29902 ;
  assign n29904 = ~n29901 & ~n29903 ;
  assign n29905 = n26554 & ~n29904 ;
  assign n29906 = n1358 & n29905 ;
  assign n29907 = \pi0038  & ~n29906 ;
  assign n29908 = ~\pi0723  & ~n29907 ;
  assign n29909 = ~\pi0173  & ~\pi0723  ;
  assign n29910 = ~n26566 & n29909 ;
  assign n29911 = ~\pi0745  & n29909 ;
  assign n29912 = ~n22536 & n29911 ;
  assign n29913 = ~n29910 & ~n29912 ;
  assign n29914 = ~n29908 & n29913 ;
  assign n29915 = n6861 & n29914 ;
  assign n29916 = ~n29882 & ~n29915 ;
  assign n29917 = ~n29898 & n29916 ;
  assign n29918 = ~n29883 & ~n29917 ;
  assign n29919 = \pi0609  & ~n29918 ;
  assign n29920 = ~\pi0173  & ~\pi0625  ;
  assign n29921 = ~n22734 & ~n29920 ;
  assign n29922 = n29880 & ~n29921 ;
  assign n29923 = ~n29915 & ~n29921 ;
  assign n29924 = ~n29898 & n29923 ;
  assign n29925 = ~n29922 & ~n29924 ;
  assign n29926 = n6861 & ~n29879 ;
  assign n29927 = ~\pi0173  & \pi0625  ;
  assign n29928 = ~n22727 & ~n29927 ;
  assign n29929 = ~n29926 & ~n29928 ;
  assign n29930 = ~\pi1153  & ~n29929 ;
  assign n29931 = n29925 & n29930 ;
  assign n29932 = ~\pi0074  & ~\pi0723  ;
  assign n29933 = ~\pi0100  & n29932 ;
  assign n29934 = n1287 & n29933 ;
  assign n29935 = ~\pi0173  & ~n29934 ;
  assign n29936 = n21768 & n29935 ;
  assign n29937 = n21770 & n29935 ;
  assign n29938 = ~n21734 & n29937 ;
  assign n29939 = ~n29936 & ~n29938 ;
  assign n29940 = \pi0625  & ~n29939 ;
  assign n29941 = ~\pi0038  & ~\pi0173  ;
  assign n29942 = n6861 & ~n29941 ;
  assign n29943 = ~n22109 & n29942 ;
  assign n29944 = ~\pi0173  & ~n22017 ;
  assign n29945 = ~n21994 & n29944 ;
  assign n29946 = ~n29943 & ~n29945 ;
  assign n29947 = ~\pi0173  & ~n21757 ;
  assign n29948 = n22117 & ~n29947 ;
  assign n29949 = ~\pi0723  & ~n29948 ;
  assign n29950 = \pi0625  & n29949 ;
  assign n29951 = ~n29946 & n29950 ;
  assign n29952 = ~n29940 & ~n29951 ;
  assign n29953 = n21768 & n29920 ;
  assign n29954 = n21770 & n29920 ;
  assign n29955 = ~n21734 & n29954 ;
  assign n29956 = ~n29953 & ~n29955 ;
  assign n29957 = \pi1153  & n29956 ;
  assign n29958 = n29952 & n29957 ;
  assign n29959 = ~\pi0608  & ~n29958 ;
  assign n29960 = ~n29931 & n29959 ;
  assign n29961 = n29880 & ~n29928 ;
  assign n29962 = ~n29915 & ~n29928 ;
  assign n29963 = ~n29898 & n29962 ;
  assign n29964 = ~n29961 & ~n29963 ;
  assign n29965 = \pi1153  & n29921 ;
  assign n29966 = n23606 & ~n29879 ;
  assign n29967 = ~n29965 & ~n29966 ;
  assign n29968 = n29964 & ~n29967 ;
  assign n29969 = ~\pi0625  & ~n29939 ;
  assign n29970 = ~\pi0625  & n29949 ;
  assign n29971 = ~n29946 & n29970 ;
  assign n29972 = ~n29969 & ~n29971 ;
  assign n29973 = n21768 & n29927 ;
  assign n29974 = n21770 & n29927 ;
  assign n29975 = ~n21734 & n29974 ;
  assign n29976 = ~n29973 & ~n29975 ;
  assign n29977 = ~\pi1153  & n29976 ;
  assign n29978 = n29972 & n29977 ;
  assign n29979 = \pi0608  & ~n29978 ;
  assign n29980 = ~n29968 & n29979 ;
  assign n29981 = ~n29960 & ~n29980 ;
  assign n29982 = n23638 & ~n29981 ;
  assign n29983 = ~n29919 & ~n29982 ;
  assign n29984 = \pi0173  & ~n6861 ;
  assign n29985 = ~n20985 & n29984 ;
  assign n29986 = n21774 & n29985 ;
  assign n29987 = n26646 & ~n29879 ;
  assign n29988 = ~n29986 & ~n29987 ;
  assign n29989 = ~\pi0173  & n21768 ;
  assign n29990 = ~\pi0173  & n21770 ;
  assign n29991 = ~n21734 & n29990 ;
  assign n29992 = ~n29989 & ~n29991 ;
  assign n29993 = n26653 & n29992 ;
  assign n29994 = ~\pi0660  & ~n29993 ;
  assign n29995 = n29988 & n29994 ;
  assign n29996 = ~n29946 & n29949 ;
  assign n29997 = ~\pi0778  & n29939 ;
  assign n29998 = ~n29996 & n29997 ;
  assign n29999 = ~\pi0609  & ~n29998 ;
  assign n30000 = \pi1155  & ~n29999 ;
  assign n30001 = ~n29958 & ~n29978 ;
  assign n30002 = n22722 & ~n30001 ;
  assign n30003 = ~n30000 & ~n30002 ;
  assign n30004 = ~n29995 & ~n30003 ;
  assign n30005 = n29983 & n30004 ;
  assign n30006 = \pi0778  & ~n29981 ;
  assign n30007 = \pi0778  & ~n30001 ;
  assign n30008 = \pi0609  & ~n29998 ;
  assign n30009 = ~n30007 & n30008 ;
  assign n30010 = ~\pi1155  & n29985 ;
  assign n30011 = n26672 & ~n29879 ;
  assign n30012 = ~n30010 & ~n30011 ;
  assign n30013 = ~\pi0609  & ~n30012 ;
  assign n30014 = n26676 & n29992 ;
  assign n30015 = ~n22787 & ~n30014 ;
  assign n30016 = ~n30013 & n30015 ;
  assign n30017 = ~n30009 & ~n30016 ;
  assign n30018 = \pi0785  & ~n30017 ;
  assign n30019 = n29918 & ~n30018 ;
  assign n30020 = ~n30006 & n30019 ;
  assign n30021 = n20999 & n29985 ;
  assign n30022 = n26685 & ~n29879 ;
  assign n30023 = ~n30021 & ~n30022 ;
  assign n30024 = \pi0660  & ~n30014 ;
  assign n30025 = n30023 & n30024 ;
  assign n30026 = ~n29995 & ~n30025 ;
  assign n30027 = \pi0609  & ~n30015 ;
  assign n30028 = n29998 & n30027 ;
  assign n30029 = \pi0778  & n30027 ;
  assign n30030 = ~n30001 & n30029 ;
  assign n30031 = ~n30028 & ~n30030 ;
  assign n30032 = ~n30026 & n30031 ;
  assign n30033 = ~n30020 & n30032 ;
  assign n30034 = ~n30005 & n30033 ;
  assign n30035 = ~\pi0785  & ~n30020 ;
  assign n30036 = n26700 & ~n30035 ;
  assign n30037 = ~n30034 & n30036 ;
  assign n30038 = n23456 & ~n29879 ;
  assign n30039 = n21777 & n29984 ;
  assign n30040 = ~n21777 & n29992 ;
  assign n30041 = n20811 & ~n30040 ;
  assign n30042 = ~n30039 & n30041 ;
  assign n30043 = ~n30038 & n30042 ;
  assign n30044 = ~\pi0173  & ~n20811 ;
  assign n30045 = n21768 & n30044 ;
  assign n30046 = n21770 & n30044 ;
  assign n30047 = ~n21734 & n30046 ;
  assign n30048 = ~n30045 & ~n30047 ;
  assign n30049 = n22155 & n30048 ;
  assign n30050 = ~n30043 & n30049 ;
  assign n30051 = ~n22147 & ~n29998 ;
  assign n30052 = n22147 & ~n29992 ;
  assign n30053 = n23666 & n23830 ;
  assign n30054 = ~n30052 & n30053 ;
  assign n30055 = ~n30051 & n30054 ;
  assign n30056 = \pi0778  & n30054 ;
  assign n30057 = ~n30001 & n30056 ;
  assign n30058 = ~n30055 & ~n30057 ;
  assign n30059 = ~n30050 & n30058 ;
  assign n30060 = ~n21034 & ~n30059 ;
  assign n30061 = ~\pi0173  & ~n20778 ;
  assign n30062 = n21768 & n30061 ;
  assign n30063 = n21770 & n30061 ;
  assign n30064 = ~n21734 & n30063 ;
  assign n30065 = ~n30062 & ~n30064 ;
  assign n30066 = \pi0788  & ~n30065 ;
  assign n30067 = ~\pi0781  & ~n30040 ;
  assign n30068 = ~n23423 & ~n30039 ;
  assign n30069 = n30067 & n30068 ;
  assign n30070 = ~n30038 & n30069 ;
  assign n30071 = n23423 & ~n29992 ;
  assign n30072 = ~n30070 & ~n30071 ;
  assign n30073 = n20816 & ~n30072 ;
  assign n30074 = ~n30043 & n30048 ;
  assign n30075 = n26728 & ~n30074 ;
  assign n30076 = ~n30073 & ~n30075 ;
  assign n30077 = ~n30066 & n30076 ;
  assign n30078 = ~\pi0788  & ~n30072 ;
  assign n30079 = n26733 & ~n30074 ;
  assign n30080 = ~n30078 & ~n30079 ;
  assign n30081 = n24691 & n30080 ;
  assign n30082 = n30077 & n30081 ;
  assign n30083 = n26065 & ~n30001 ;
  assign n30084 = n26739 & n29939 ;
  assign n30085 = ~n29996 & n30084 ;
  assign n30086 = ~n23885 & n29992 ;
  assign n30087 = ~\pi0628  & ~n30086 ;
  assign n30088 = ~n30085 & n30087 ;
  assign n30089 = ~n30083 & n30088 ;
  assign n30090 = ~\pi0173  & \pi0628  ;
  assign n30091 = n21768 & n30090 ;
  assign n30092 = n21770 & n30090 ;
  assign n30093 = ~n21734 & n30092 ;
  assign n30094 = ~n30091 & ~n30093 ;
  assign n30095 = n20844 & n30094 ;
  assign n30096 = ~n30089 & n30095 ;
  assign n30097 = \pi0628  & ~n30086 ;
  assign n30098 = ~n30085 & n30097 ;
  assign n30099 = ~n30083 & n30098 ;
  assign n30100 = ~\pi0173  & ~\pi0628  ;
  assign n30101 = n21768 & n30100 ;
  assign n30102 = n21770 & n30100 ;
  assign n30103 = ~n21734 & n30102 ;
  assign n30104 = ~n30101 & ~n30103 ;
  assign n30105 = n20843 & n30104 ;
  assign n30106 = ~n30099 & n30105 ;
  assign n30107 = ~n30096 & ~n30106 ;
  assign n30108 = ~n30082 & n30107 ;
  assign n30109 = \pi0792  & ~n30108 ;
  assign n30110 = n23380 & ~n29998 ;
  assign n30111 = ~\pi0173  & ~n26770 ;
  assign n30112 = n21050 & ~n30111 ;
  assign n30113 = ~n30110 & n30112 ;
  assign n30114 = \pi0778  & n30112 ;
  assign n30115 = ~n30001 & n30114 ;
  assign n30116 = ~n30113 & ~n30115 ;
  assign n30117 = \pi0789  & ~n30116 ;
  assign n30118 = n23683 & ~n30074 ;
  assign n30119 = n21032 & ~n30039 ;
  assign n30120 = n30067 & n30119 ;
  assign n30121 = ~n30038 & n30120 ;
  assign n30122 = ~n21032 & ~n29992 ;
  assign n30123 = ~n20876 & ~n30122 ;
  assign n30124 = ~n30121 & n30123 ;
  assign n30125 = \pi0789  & n30124 ;
  assign n30126 = ~n30118 & n30125 ;
  assign n30127 = ~n30117 & ~n30126 ;
  assign n30128 = ~n21038 & n30127 ;
  assign n30129 = ~n30109 & n30128 ;
  assign n30130 = ~n30060 & n30129 ;
  assign n30131 = ~n30037 & n30130 ;
  assign n30132 = ~n20883 & ~n30065 ;
  assign n30133 = n20947 & ~n30072 ;
  assign n30134 = n26806 & ~n30074 ;
  assign n30135 = ~n30133 & ~n30134 ;
  assign n30136 = ~n30132 & n30135 ;
  assign n30137 = ~n22160 & ~n30111 ;
  assign n30138 = ~n30110 & n30137 ;
  assign n30139 = \pi0778  & n30137 ;
  assign n30140 = ~n30001 & n30139 ;
  assign n30141 = ~n30138 & ~n30140 ;
  assign n30142 = n20951 & ~n29992 ;
  assign n30143 = ~n23838 & ~n30142 ;
  assign n30144 = n30141 & ~n30143 ;
  assign n30145 = ~n23856 & ~n30144 ;
  assign n30146 = n30136 & n30145 ;
  assign n30147 = ~n26803 & ~n30146 ;
  assign n30148 = ~n30109 & n30147 ;
  assign n30149 = ~n21067 & ~n30148 ;
  assign n30150 = ~n30131 & n30149 ;
  assign n30151 = n21092 & n30080 ;
  assign n30152 = n30077 & n30151 ;
  assign n30153 = ~n21092 & n29992 ;
  assign n30154 = n26824 & ~n30153 ;
  assign n30155 = ~n30152 & n30154 ;
  assign n30156 = ~\pi0173  & ~\pi0644  ;
  assign n30157 = n21768 & n30156 ;
  assign n30158 = n21770 & n30156 ;
  assign n30159 = ~n21734 & n30158 ;
  assign n30160 = ~n30157 & ~n30159 ;
  assign n30161 = ~\pi0715  & n30160 ;
  assign n30162 = n26824 & ~n30161 ;
  assign n30163 = \pi0790  & ~n30162 ;
  assign n30164 = ~n30155 & n30163 ;
  assign n30165 = ~n30085 & ~n30086 ;
  assign n30166 = ~n30083 & n30165 ;
  assign n30167 = ~\pi0792  & ~n30166 ;
  assign n30168 = ~\pi0647  & ~n30167 ;
  assign n30169 = n21768 & n29736 ;
  assign n30170 = n21770 & n29736 ;
  assign n30171 = ~n21734 & n30170 ;
  assign n30172 = ~n30169 & ~n30171 ;
  assign n30173 = n20897 & n30172 ;
  assign n30174 = ~n30168 & n30173 ;
  assign n30175 = \pi1156  & n30104 ;
  assign n30176 = ~n30099 & n30175 ;
  assign n30177 = ~\pi1156  & n30094 ;
  assign n30178 = ~n30089 & n30177 ;
  assign n30179 = ~n30176 & ~n30178 ;
  assign n30180 = \pi0792  & n30173 ;
  assign n30181 = ~n30179 & n30180 ;
  assign n30182 = ~n30174 & ~n30181 ;
  assign n30183 = n20846 & ~n29992 ;
  assign n30184 = ~n20910 & ~n30183 ;
  assign n30185 = n20846 & n30184 ;
  assign n30186 = n30080 & n30184 ;
  assign n30187 = n30077 & n30186 ;
  assign n30188 = ~n30185 & ~n30187 ;
  assign n30189 = \pi0647  & ~n30167 ;
  assign n30190 = ~\pi0173  & ~\pi0647  ;
  assign n30191 = n21768 & n30190 ;
  assign n30192 = n21770 & n30190 ;
  assign n30193 = ~n21734 & n30192 ;
  assign n30194 = ~n30191 & ~n30193 ;
  assign n30195 = n20849 & n30194 ;
  assign n30196 = ~n30189 & n30195 ;
  assign n30197 = \pi0792  & n30195 ;
  assign n30198 = ~n30179 & n30197 ;
  assign n30199 = ~n30196 & ~n30198 ;
  assign n30200 = n30188 & n30199 ;
  assign n30201 = n30182 & n30200 ;
  assign n30202 = \pi0787  & ~n30201 ;
  assign n30203 = ~n30164 & ~n30202 ;
  assign n30204 = ~n30150 & n30203 ;
  assign n30205 = n9948 & ~n29855 ;
  assign n30206 = n30204 & n30205 ;
  assign n30207 = ~\pi0787  & n30167 ;
  assign n30208 = n23011 & ~n30179 ;
  assign n30209 = ~n30207 & ~n30208 ;
  assign n30210 = \pi0644  & ~n30209 ;
  assign n30211 = \pi1157  & n30194 ;
  assign n30212 = ~n30189 & n30211 ;
  assign n30213 = \pi0792  & n30211 ;
  assign n30214 = ~n30179 & n30213 ;
  assign n30215 = ~n30212 & ~n30214 ;
  assign n30216 = ~\pi1157  & n30172 ;
  assign n30217 = ~n30168 & n30216 ;
  assign n30218 = \pi0792  & n30216 ;
  assign n30219 = ~n30179 & n30218 ;
  assign n30220 = ~n30217 & ~n30219 ;
  assign n30221 = n30215 & n30220 ;
  assign n30222 = n23074 & ~n30221 ;
  assign n30223 = ~n30210 & ~n30222 ;
  assign n30224 = \pi0644  & n30223 ;
  assign n30225 = ~n30202 & n30223 ;
  assign n30226 = ~n30150 & n30225 ;
  assign n30227 = ~n30224 & ~n30226 ;
  assign n30228 = n23316 & ~n30227 ;
  assign n30229 = ~\pi0173  & \pi0715  ;
  assign n30230 = n21768 & n30229 ;
  assign n30231 = n21770 & n30229 ;
  assign n30232 = ~n21734 & n30231 ;
  assign n30233 = ~n30230 & ~n30232 ;
  assign n30234 = ~n23313 & n30233 ;
  assign n30235 = ~\pi1160  & ~n30153 ;
  assign n30236 = ~n30152 & n30235 ;
  assign n30237 = ~n26911 & ~n30236 ;
  assign n30238 = ~n30234 & ~n30237 ;
  assign n30239 = ~\pi0644  & n30209 ;
  assign n30240 = \pi0715  & ~n30239 ;
  assign n30241 = n26918 & ~n30221 ;
  assign n30242 = ~n30240 & ~n30241 ;
  assign n30243 = \pi1160  & ~n30161 ;
  assign n30244 = ~n30155 & ~n30243 ;
  assign n30245 = n30242 & ~n30244 ;
  assign n30246 = ~n30238 & ~n30245 ;
  assign n30247 = ~n30228 & n30246 ;
  assign n30248 = \pi0790  & n30205 ;
  assign n30249 = ~n30247 & n30248 ;
  assign n30250 = ~n30206 & ~n30249 ;
  assign n30251 = ~n29856 & n30250 ;
  assign n30252 = ~\pi0174  & ~n6848 ;
  assign n30253 = ~\pi0057  & ~n30252 ;
  assign n30254 = \pi0057  & \pi0174  ;
  assign n30255 = ~n30253 & ~n30254 ;
  assign n30256 = \pi0174  & n21768 ;
  assign n30257 = \pi0174  & n21770 ;
  assign n30258 = ~n21734 & n30257 ;
  assign n30259 = ~n30256 & ~n30258 ;
  assign n30260 = ~\pi0074  & \pi0696  ;
  assign n30261 = ~\pi0100  & n30260 ;
  assign n30262 = n1287 & n30261 ;
  assign n30263 = n30259 & ~n30262 ;
  assign n30264 = \pi0174  & n22017 ;
  assign n30265 = \pi0039  & \pi0174  ;
  assign n30266 = ~n21993 & n30265 ;
  assign n30267 = ~n30264 & ~n30266 ;
  assign n30268 = ~\pi0174  & ~n22107 ;
  assign n30269 = n22089 & n30268 ;
  assign n30270 = ~\pi0038  & ~n30269 ;
  assign n30271 = n30267 & n30270 ;
  assign n30272 = ~\pi0174  & ~n21757 ;
  assign n30273 = n25669 & ~n30272 ;
  assign n30274 = n30262 & ~n30273 ;
  assign n30275 = ~n30271 & n30274 ;
  assign n30276 = ~n30263 & ~n30275 ;
  assign n30277 = ~\pi0778  & n30276 ;
  assign n30278 = n23380 & ~n30277 ;
  assign n30279 = ~n23380 & n30259 ;
  assign n30280 = ~n30278 & ~n30279 ;
  assign n30281 = \pi0625  & ~n30276 ;
  assign n30282 = \pi0174  & \pi1153  ;
  assign n30283 = n21768 & n30282 ;
  assign n30284 = n21770 & n30282 ;
  assign n30285 = ~n21734 & n30284 ;
  assign n30286 = ~n30283 & ~n30285 ;
  assign n30287 = ~n24550 & n30286 ;
  assign n30288 = ~n30281 & ~n30287 ;
  assign n30289 = ~\pi0625  & ~n30276 ;
  assign n30290 = \pi0174  & ~\pi1153  ;
  assign n30291 = n21768 & n30290 ;
  assign n30292 = n21770 & n30290 ;
  assign n30293 = ~n21734 & n30292 ;
  assign n30294 = ~n30291 & ~n30293 ;
  assign n30295 = ~n24561 & n30294 ;
  assign n30296 = ~n30289 & ~n30295 ;
  assign n30297 = ~n30288 & ~n30296 ;
  assign n30298 = \pi0778  & ~n30279 ;
  assign n30299 = ~n30297 & n30298 ;
  assign n30300 = ~n30280 & ~n30299 ;
  assign n30301 = n22162 & n30300 ;
  assign n30302 = ~n22162 & n30259 ;
  assign n30303 = ~\pi0792  & ~n30302 ;
  assign n30304 = ~n30301 & n30303 ;
  assign n30305 = ~\pi0647  & ~n30304 ;
  assign n30306 = \pi0647  & n30259 ;
  assign n30307 = n20897 & ~n30306 ;
  assign n30308 = ~n30305 & n30307 ;
  assign n30309 = \pi0628  & n30302 ;
  assign n30310 = \pi0628  & n22162 ;
  assign n30311 = n30300 & n30310 ;
  assign n30312 = ~n30309 & ~n30311 ;
  assign n30313 = ~\pi0628  & n30259 ;
  assign n30314 = \pi1156  & ~n30313 ;
  assign n30315 = n30312 & n30314 ;
  assign n30316 = ~\pi0628  & n30302 ;
  assign n30317 = ~\pi0628  & n22162 ;
  assign n30318 = n30300 & n30317 ;
  assign n30319 = ~n30316 & ~n30318 ;
  assign n30320 = \pi0628  & n30259 ;
  assign n30321 = ~\pi1156  & ~n30320 ;
  assign n30322 = n30319 & n30321 ;
  assign n30323 = ~n30315 & ~n30322 ;
  assign n30324 = \pi0792  & n30307 ;
  assign n30325 = ~n30323 & n30324 ;
  assign n30326 = ~n30308 & ~n30325 ;
  assign n30327 = \pi0299  & ~\pi0759  ;
  assign n30328 = ~n21205 & n30327 ;
  assign n30329 = ~n21238 & n30328 ;
  assign n30330 = ~n21740 & n27839 ;
  assign n30331 = ~n21738 & n30330 ;
  assign n30332 = ~n30329 & ~n30331 ;
  assign n30333 = ~\pi0039  & n30332 ;
  assign n30334 = ~\pi0299  & \pi0759  ;
  assign n30335 = ~n25554 & n30334 ;
  assign n30336 = ~n30333 & ~n30335 ;
  assign n30337 = \pi0759  & ~n30335 ;
  assign n30338 = n21272 & n30337 ;
  assign n30339 = ~n30336 & ~n30338 ;
  assign n30340 = ~\pi0759  & ~n25542 ;
  assign n30341 = \pi0299  & \pi0759  ;
  assign n30342 = ~n25557 & n30341 ;
  assign n30343 = ~n30340 & ~n30342 ;
  assign n30344 = ~n30339 & n30343 ;
  assign n30345 = ~\pi0039  & ~n30332 ;
  assign n30346 = ~\pi0039  & \pi0759  ;
  assign n30347 = n21272 & n30346 ;
  assign n30348 = ~n30345 & ~n30347 ;
  assign n30349 = ~\pi0038  & \pi0174  ;
  assign n30350 = n30348 & n30349 ;
  assign n30351 = ~n30344 & n30350 ;
  assign n30352 = ~\pi0174  & \pi0759  ;
  assign n30353 = ~\pi0038  & n30352 ;
  assign n30354 = n25023 & n30353 ;
  assign n30355 = \pi0174  & ~n6861 ;
  assign n30356 = \pi0603  & \pi0759  ;
  assign n30357 = ~n20783 & n30356 ;
  assign n30358 = n1689 & ~n30357 ;
  assign n30359 = n1354 & n30358 ;
  assign n30360 = n8413 & n30359 ;
  assign n30361 = n1358 & n30360 ;
  assign n30362 = \pi0038  & ~n30361 ;
  assign n30363 = ~n30272 & n30362 ;
  assign n30364 = ~n30355 & ~n30363 ;
  assign n30365 = ~n30354 & n30364 ;
  assign n30366 = ~n30351 & n30365 ;
  assign n30367 = ~\pi0174  & ~n6861 ;
  assign n30368 = ~n20985 & ~n30367 ;
  assign n30369 = ~n30366 & n30368 ;
  assign n30370 = n20985 & ~n30259 ;
  assign n30371 = ~n25588 & ~n30370 ;
  assign n30372 = ~n30369 & n30371 ;
  assign n30373 = n21776 & n30259 ;
  assign n30374 = n23831 & ~n30373 ;
  assign n30375 = ~n30372 & n30374 ;
  assign n30376 = ~n20846 & ~n23880 ;
  assign n30377 = ~n23831 & ~n30259 ;
  assign n30378 = n30376 & ~n30377 ;
  assign n30379 = ~n30375 & n30378 ;
  assign n30380 = n30259 & ~n30376 ;
  assign n30381 = ~n20910 & ~n30380 ;
  assign n30382 = ~n30379 & n30381 ;
  assign n30383 = ~n20849 & ~n30382 ;
  assign n30384 = \pi0647  & n30304 ;
  assign n30385 = n22956 & ~n30323 ;
  assign n30386 = ~n30384 & ~n30385 ;
  assign n30387 = \pi0174  & ~\pi0647  ;
  assign n30388 = n21768 & n30387 ;
  assign n30389 = n21770 & n30387 ;
  assign n30390 = ~n21734 & n30389 ;
  assign n30391 = ~n30388 & ~n30390 ;
  assign n30392 = ~n30382 & n30391 ;
  assign n30393 = n30386 & n30392 ;
  assign n30394 = ~n30383 & ~n30393 ;
  assign n30395 = n30326 & ~n30394 ;
  assign n30396 = \pi0787  & ~n30395 ;
  assign n30397 = n23413 & n30259 ;
  assign n30398 = ~n24781 & ~n30397 ;
  assign n30399 = ~n30380 & ~n30397 ;
  assign n30400 = ~n30379 & n30399 ;
  assign n30401 = ~n30398 & ~n30400 ;
  assign n30402 = n24777 & n30259 ;
  assign n30403 = \pi0790  & ~n30402 ;
  assign n30404 = \pi0644  & n30403 ;
  assign n30405 = ~n30401 & n30404 ;
  assign n30406 = n23412 & n30259 ;
  assign n30407 = ~n24766 & ~n30406 ;
  assign n30408 = ~n30380 & ~n30406 ;
  assign n30409 = ~n30379 & n30408 ;
  assign n30410 = ~n30407 & ~n30409 ;
  assign n30411 = ~\pi0644  & n30403 ;
  assign n30412 = ~n30410 & n30411 ;
  assign n30413 = ~n30405 & ~n30412 ;
  assign n30414 = \pi0790  & n30413 ;
  assign n30415 = \pi0787  & ~n30306 ;
  assign n30416 = ~n30305 & n30415 ;
  assign n30417 = \pi0792  & n30415 ;
  assign n30418 = ~n30323 & n30417 ;
  assign n30419 = ~n30416 & ~n30418 ;
  assign n30420 = ~n24994 & n30419 ;
  assign n30421 = \pi1157  & n30391 ;
  assign n30422 = n30386 & n30421 ;
  assign n30423 = ~n30420 & ~n30422 ;
  assign n30424 = n23011 & ~n30323 ;
  assign n30425 = ~\pi0787  & ~\pi0792  ;
  assign n30426 = ~n30302 & n30425 ;
  assign n30427 = ~n30301 & n30426 ;
  assign n30428 = n23518 & ~n30427 ;
  assign n30429 = ~n30424 & n30428 ;
  assign n30430 = \pi0790  & n30429 ;
  assign n30431 = ~n30423 & n30430 ;
  assign n30432 = ~n30414 & ~n30431 ;
  assign n30433 = n30396 & n30432 ;
  assign n30434 = n21034 & ~n21038 ;
  assign n30435 = ~n30364 & ~n30367 ;
  assign n30436 = \pi0038  & ~n25217 ;
  assign n30437 = \pi0174  & ~\pi0299  ;
  assign n30438 = n22407 & n30437 ;
  assign n30439 = \pi0174  & \pi0299  ;
  assign n30440 = n22291 & n30439 ;
  assign n30441 = ~n30438 & ~n30440 ;
  assign n30442 = \pi0299  & ~n22431 ;
  assign n30443 = ~\pi0174  & ~n22379 ;
  assign n30444 = ~n30442 & n30443 ;
  assign n30445 = n30441 & ~n30444 ;
  assign n30446 = ~\pi0759  & n30445 ;
  assign n30447 = \pi0299  & ~n22530 ;
  assign n30448 = n22487 & ~n22509 ;
  assign n30449 = ~\pi0174  & n22468 ;
  assign n30450 = ~n30448 & n30449 ;
  assign n30451 = ~n30447 & n30450 ;
  assign n30452 = n22601 & n30437 ;
  assign n30453 = n22630 & n30439 ;
  assign n30454 = \pi0759  & ~n30453 ;
  assign n30455 = ~n30452 & n30454 ;
  assign n30456 = ~n30451 & n30455 ;
  assign n30457 = \pi0039  & ~n30456 ;
  assign n30458 = ~n30446 & n30457 ;
  assign n30459 = \pi0174  & n22643 ;
  assign n30460 = ~n22652 & n30459 ;
  assign n30461 = ~\pi0174  & ~\pi0299  ;
  assign n30462 = n22676 & n30461 ;
  assign n30463 = ~\pi0174  & \pi0299  ;
  assign n30464 = ~n22657 & n30463 ;
  assign n30465 = ~n22660 & n30464 ;
  assign n30466 = n22664 & n30465 ;
  assign n30467 = ~\pi0759  & ~n30466 ;
  assign n30468 = ~n30462 & n30467 ;
  assign n30469 = ~n30460 & n30468 ;
  assign n30470 = \pi0759  & n21272 ;
  assign n30471 = n22006 & n30439 ;
  assign n30472 = n22649 & n30437 ;
  assign n30473 = ~n30471 & ~n30472 ;
  assign n30474 = n30470 & ~n30473 ;
  assign n30475 = n22693 & n30352 ;
  assign n30476 = ~\pi0039  & ~n30475 ;
  assign n30477 = ~n30474 & n30476 ;
  assign n30478 = ~n30469 & n30477 ;
  assign n30479 = \pi0696  & ~n25217 ;
  assign n30480 = ~n30478 & n30479 ;
  assign n30481 = ~n30458 & n30480 ;
  assign n30482 = ~n30436 & ~n30481 ;
  assign n30483 = ~\pi0696  & ~n30354 ;
  assign n30484 = ~n30351 & n30483 ;
  assign n30485 = ~n30367 & ~n30484 ;
  assign n30486 = n30482 & n30485 ;
  assign n30487 = ~n30435 & ~n30486 ;
  assign n30488 = \pi0608  & \pi0625  ;
  assign n30489 = n30295 & n30488 ;
  assign n30490 = n30487 & n30489 ;
  assign n30491 = ~\pi0608  & ~\pi0625  ;
  assign n30492 = n30287 & n30491 ;
  assign n30493 = n30487 & n30492 ;
  assign n30494 = ~\pi1153  & ~n30367 ;
  assign n30495 = ~n30366 & n30494 ;
  assign n30496 = ~n24561 & ~n30495 ;
  assign n30497 = ~\pi0608  & n30287 ;
  assign n30498 = n22755 & ~n30276 ;
  assign n30499 = ~n30497 & ~n30498 ;
  assign n30500 = n30496 & ~n30499 ;
  assign n30501 = \pi0608  & n30295 ;
  assign n30502 = n22740 & ~n30276 ;
  assign n30503 = ~n30501 & ~n30502 ;
  assign n30504 = \pi1153  & ~n30367 ;
  assign n30505 = ~n30366 & n30504 ;
  assign n30506 = ~n24550 & ~n30505 ;
  assign n30507 = ~n30503 & n30506 ;
  assign n30508 = ~n30500 & ~n30507 ;
  assign n30509 = ~n30493 & n30508 ;
  assign n30510 = ~n30490 & n30509 ;
  assign n30511 = \pi0778  & ~n30510 ;
  assign n30512 = ~\pi0778  & n30487 ;
  assign n30513 = ~n23808 & ~n30512 ;
  assign n30514 = n21022 & n30513 ;
  assign n30515 = ~n30511 & n30514 ;
  assign n30516 = n20811 & n30373 ;
  assign n30517 = n20811 & n30371 ;
  assign n30518 = ~n30369 & n30517 ;
  assign n30519 = ~n30516 & ~n30518 ;
  assign n30520 = n20811 & n20871 ;
  assign n30521 = \pi0174  & n20871 ;
  assign n30522 = n21768 & n30521 ;
  assign n30523 = n21770 & n30521 ;
  assign n30524 = ~n21734 & n30523 ;
  assign n30525 = ~n30522 & ~n30524 ;
  assign n30526 = ~n30520 & n30525 ;
  assign n30527 = \pi0781  & ~n30526 ;
  assign n30528 = n30519 & n30527 ;
  assign n30529 = n22148 & ~n30297 ;
  assign n30530 = n22151 & n30276 ;
  assign n30531 = n22147 & ~n30259 ;
  assign n30532 = ~n30530 & ~n30531 ;
  assign n30533 = ~n30529 & n30532 ;
  assign n30534 = n30053 & ~n30533 ;
  assign n30535 = ~n30528 & ~n30534 ;
  assign n30536 = n26125 & n30276 ;
  assign n30537 = ~n26119 & ~n30297 ;
  assign n30538 = ~n30536 & ~n30537 ;
  assign n30539 = ~\pi0609  & ~n30370 ;
  assign n30540 = ~n30369 & n30539 ;
  assign n30541 = \pi0609  & n30259 ;
  assign n30542 = n20865 & ~n30541 ;
  assign n30543 = ~n30540 & n30542 ;
  assign n30544 = \pi0609  & ~n30370 ;
  assign n30545 = ~n30369 & n30544 ;
  assign n30546 = ~\pi0609  & n30259 ;
  assign n30547 = n20864 & ~n30546 ;
  assign n30548 = ~n30545 & n30547 ;
  assign n30549 = ~n30543 & ~n30548 ;
  assign n30550 = n30538 & n30549 ;
  assign n30551 = n21023 & ~n30550 ;
  assign n30552 = n30535 & ~n30551 ;
  assign n30553 = ~n21038 & n30552 ;
  assign n30554 = ~n30515 & n30553 ;
  assign n30555 = ~n30434 & ~n30554 ;
  assign n30556 = n21050 & ~n30300 ;
  assign n30557 = ~\pi0619  & ~n23830 ;
  assign n30558 = n30373 & n30557 ;
  assign n30559 = n30371 & n30557 ;
  assign n30560 = ~n30369 & n30559 ;
  assign n30561 = ~n30558 & ~n30560 ;
  assign n30562 = n20874 & ~n30259 ;
  assign n30563 = ~\pi0619  & n20874 ;
  assign n30564 = ~n23830 & n30563 ;
  assign n30565 = ~n30562 & ~n30564 ;
  assign n30566 = n30561 & ~n30565 ;
  assign n30567 = \pi0619  & ~n23830 ;
  assign n30568 = n30373 & n30567 ;
  assign n30569 = n30371 & n30567 ;
  assign n30570 = ~n30369 & n30569 ;
  assign n30571 = ~n30568 & ~n30570 ;
  assign n30572 = \pi0619  & n23830 ;
  assign n30573 = n30259 & n30572 ;
  assign n30574 = ~\pi0619  & n30259 ;
  assign n30575 = n20875 & ~n30574 ;
  assign n30576 = ~n30573 & n30575 ;
  assign n30577 = n30571 & n30576 ;
  assign n30578 = ~n30566 & ~n30577 ;
  assign n30579 = ~n30556 & n30578 ;
  assign n30580 = \pi0789  & ~n30579 ;
  assign n30581 = \pi0628  & ~n30580 ;
  assign n30582 = ~n30555 & n30581 ;
  assign n30583 = n22160 & n30259 ;
  assign n30584 = \pi0641  & ~n30583 ;
  assign n30585 = \pi0174  & ~\pi0641  ;
  assign n30586 = n21768 & n30585 ;
  assign n30587 = n21770 & n30585 ;
  assign n30588 = ~n21734 & n30587 ;
  assign n30589 = ~n30586 & ~n30588 ;
  assign n30590 = ~n30584 & n30589 ;
  assign n30591 = ~n22160 & n30589 ;
  assign n30592 = n30300 & n30591 ;
  assign n30593 = ~n30590 & ~n30592 ;
  assign n30594 = n20776 & ~n30593 ;
  assign n30595 = ~\pi0641  & ~n30583 ;
  assign n30596 = \pi0174  & \pi0641  ;
  assign n30597 = n21768 & n30596 ;
  assign n30598 = n21770 & n30596 ;
  assign n30599 = ~n21734 & n30598 ;
  assign n30600 = ~n30597 & ~n30599 ;
  assign n30601 = n20777 & n30600 ;
  assign n30602 = ~n30595 & n30601 ;
  assign n30603 = ~n22160 & n30601 ;
  assign n30604 = n30300 & n30603 ;
  assign n30605 = ~n30602 & ~n30604 ;
  assign n30606 = ~n20883 & ~n20950 ;
  assign n30607 = ~n30377 & n30606 ;
  assign n30608 = ~n30375 & n30607 ;
  assign n30609 = n30605 & ~n30608 ;
  assign n30610 = ~n30594 & n30609 ;
  assign n30611 = \pi0628  & \pi0788  ;
  assign n30612 = ~n30610 & n30611 ;
  assign n30613 = n23880 & ~n30259 ;
  assign n30614 = ~\pi0628  & ~n30613 ;
  assign n30615 = n23880 & n30614 ;
  assign n30616 = ~n30377 & n30614 ;
  assign n30617 = ~n30375 & n30616 ;
  assign n30618 = ~n30615 & ~n30617 ;
  assign n30619 = \pi1156  & n30618 ;
  assign n30620 = ~n30612 & n30619 ;
  assign n30621 = ~n30582 & n30620 ;
  assign n30622 = \pi0629  & ~n30322 ;
  assign n30623 = ~n30621 & n30622 ;
  assign n30624 = ~\pi0628  & ~n30580 ;
  assign n30625 = ~n30555 & n30624 ;
  assign n30626 = ~\pi0628  & \pi0788  ;
  assign n30627 = ~n30610 & n30626 ;
  assign n30628 = \pi0628  & ~n30613 ;
  assign n30629 = n23880 & n30628 ;
  assign n30630 = ~n30377 & n30628 ;
  assign n30631 = ~n30375 & n30630 ;
  assign n30632 = ~n30629 & ~n30631 ;
  assign n30633 = ~\pi1156  & n30632 ;
  assign n30634 = ~n30627 & n30633 ;
  assign n30635 = ~n30625 & n30634 ;
  assign n30636 = ~\pi0629  & ~n30315 ;
  assign n30637 = ~n30635 & n30636 ;
  assign n30638 = ~n30623 & ~n30637 ;
  assign n30639 = \pi0792  & ~n30638 ;
  assign n30640 = ~\pi0792  & ~n30580 ;
  assign n30641 = ~n30555 & n30640 ;
  assign n30642 = n23263 & ~n30610 ;
  assign n30643 = ~n21067 & ~n30642 ;
  assign n30644 = ~n30641 & n30643 ;
  assign n30645 = n30432 & n30644 ;
  assign n30646 = ~n30639 & n30645 ;
  assign n30647 = ~n30433 & ~n30646 ;
  assign n30648 = ~n30423 & n30429 ;
  assign n30649 = ~n23318 & ~n30413 ;
  assign n30650 = ~n30648 & n30649 ;
  assign n30651 = n6848 & ~n30650 ;
  assign n30652 = ~n30254 & n30651 ;
  assign n30653 = n30647 & n30652 ;
  assign n30654 = ~n30255 & ~n30653 ;
  assign n30655 = ~\pi0832  & ~n30654 ;
  assign n30656 = \pi0696  & n1689 ;
  assign n30657 = n20855 & n30656 ;
  assign n30658 = \pi0174  & ~n1689 ;
  assign n30659 = ~n30657 & ~n30658 ;
  assign n30660 = ~\pi0778  & ~n30659 ;
  assign n30661 = n23885 & n30660 ;
  assign n30662 = \pi0625  & \pi0696  ;
  assign n30663 = n1689 & n30662 ;
  assign n30664 = n20855 & n30663 ;
  assign n30665 = ~n30658 & ~n30664 ;
  assign n30666 = \pi1153  & ~n30665 ;
  assign n30667 = ~\pi1153  & ~n30664 ;
  assign n30668 = ~n30659 & n30667 ;
  assign n30669 = ~n30666 & ~n30668 ;
  assign n30670 = n26065 & ~n30669 ;
  assign n30671 = ~n30661 & ~n30670 ;
  assign n30672 = n26069 & ~n30671 ;
  assign n30673 = n26080 & n30658 ;
  assign n30674 = \pi0759  & n1689 ;
  assign n30675 = n20784 & n30674 ;
  assign n30676 = ~n23880 & n30675 ;
  assign n30677 = ~n20846 & n30676 ;
  assign n30678 = n23832 & n30677 ;
  assign n30679 = n26082 & n30678 ;
  assign n30680 = ~n30673 & ~n30679 ;
  assign n30681 = n26076 & n30658 ;
  assign n30682 = n26078 & n30678 ;
  assign n30683 = ~n30681 & ~n30682 ;
  assign n30684 = n30680 & n30683 ;
  assign n30685 = ~n30672 & n30684 ;
  assign n30686 = \pi0790  & ~n30685 ;
  assign n30687 = \pi0832  & ~n30686 ;
  assign n30688 = \pi0629  & ~n23880 ;
  assign n30689 = n30675 & n30688 ;
  assign n30690 = n23832 & n30689 ;
  assign n30691 = n20886 & ~n30690 ;
  assign n30692 = n24724 & n30691 ;
  assign n30693 = n20843 & ~n30690 ;
  assign n30694 = n24724 & n30693 ;
  assign n30695 = n30671 & n30694 ;
  assign n30696 = ~n30692 & ~n30695 ;
  assign n30697 = ~\pi0628  & ~n30671 ;
  assign n30698 = ~\pi0629  & n30676 ;
  assign n30699 = n23832 & n30698 ;
  assign n30700 = ~n25956 & ~n30699 ;
  assign n30701 = ~n21067 & n26218 ;
  assign n30702 = n30700 & n30701 ;
  assign n30703 = ~n30697 & n30702 ;
  assign n30704 = n30696 & ~n30703 ;
  assign n30705 = ~n30658 & ~n30704 ;
  assign n30706 = n21064 & ~n30678 ;
  assign n30707 = n20897 & ~n23920 ;
  assign n30708 = n20897 & ~n30661 ;
  assign n30709 = ~n30670 & n30708 ;
  assign n30710 = ~n30707 & ~n30709 ;
  assign n30711 = ~n30706 & n30710 ;
  assign n30712 = \pi0630  & \pi0647  ;
  assign n30713 = ~n23908 & ~n30712 ;
  assign n30714 = ~n30661 & ~n30712 ;
  assign n30715 = ~n30670 & n30714 ;
  assign n30716 = ~n30713 & ~n30715 ;
  assign n30717 = \pi0630  & ~n20846 ;
  assign n30718 = n30676 & n30717 ;
  assign n30719 = n23832 & n30718 ;
  assign n30720 = \pi1157  & ~n30719 ;
  assign n30721 = ~n30716 & n30720 ;
  assign n30722 = n30711 & ~n30721 ;
  assign n30723 = \pi0787  & ~n30658 ;
  assign n30724 = ~n30722 & n30723 ;
  assign n30725 = ~n30705 & ~n30724 ;
  assign n30726 = n23846 & n30660 ;
  assign n30727 = \pi0778  & n23846 ;
  assign n30728 = ~n30669 & n30727 ;
  assign n30729 = ~n30726 & ~n30728 ;
  assign n30730 = ~\pi0627  & \pi1154  ;
  assign n30731 = n30675 & n30730 ;
  assign n30732 = n21777 & n30731 ;
  assign n30733 = \pi0174  & ~\pi1154  ;
  assign n30734 = ~n1689 & n30733 ;
  assign n30735 = ~n30732 & ~n30734 ;
  assign n30736 = \pi0618  & ~n30735 ;
  assign n30737 = ~n20869 & ~n23849 ;
  assign n30738 = n30658 & n30737 ;
  assign n30739 = \pi0627  & n25612 ;
  assign n30740 = n30675 & n30739 ;
  assign n30741 = n21777 & n30740 ;
  assign n30742 = ~n30738 & ~n30741 ;
  assign n30743 = ~n30736 & n30742 ;
  assign n30744 = n30729 & n30743 ;
  assign n30745 = \pi0781  & ~n30744 ;
  assign n30746 = ~n26119 & ~n30669 ;
  assign n30747 = n26125 & ~n30659 ;
  assign n30748 = ~n20866 & n30658 ;
  assign n30749 = ~n20866 & n30675 ;
  assign n30750 = n26128 & n30749 ;
  assign n30751 = ~n30748 & ~n30750 ;
  assign n30752 = ~n30747 & n30751 ;
  assign n30753 = ~n30746 & n30752 ;
  assign n30754 = n21023 & ~n30753 ;
  assign n30755 = \pi0608  & n30664 ;
  assign n30756 = \pi0608  & ~n30658 ;
  assign n30757 = ~n30657 & n30756 ;
  assign n30758 = ~n30755 & ~n30757 ;
  assign n30759 = n26147 & n30657 ;
  assign n30760 = ~\pi1153  & ~n30759 ;
  assign n30761 = n30758 & n30760 ;
  assign n30762 = ~\pi0625  & ~n30675 ;
  assign n30763 = \pi0608  & \pi1153  ;
  assign n30764 = ~n30762 & n30763 ;
  assign n30765 = \pi0778  & ~\pi1153  ;
  assign n30766 = \pi0778  & ~n30658 ;
  assign n30767 = ~n30664 & n30766 ;
  assign n30768 = ~n30765 & ~n30767 ;
  assign n30769 = ~n30764 & ~n30768 ;
  assign n30770 = ~n30761 & n30769 ;
  assign n30771 = ~n20986 & n30657 ;
  assign n30772 = ~n30658 & ~n30675 ;
  assign n30773 = ~n30771 & n30772 ;
  assign n30774 = n21022 & ~n23808 ;
  assign n30775 = ~n30773 & n30774 ;
  assign n30776 = ~n30770 & n30775 ;
  assign n30777 = ~n21034 & ~n30776 ;
  assign n30778 = ~n30754 & n30777 ;
  assign n30779 = ~n30745 & n30778 ;
  assign n30780 = \pi0778  & n23380 ;
  assign n30781 = ~n30669 & n30780 ;
  assign n30782 = n23380 & n30660 ;
  assign n30783 = \pi0789  & ~n30658 ;
  assign n30784 = ~n29814 & n30783 ;
  assign n30785 = ~n30782 & n30784 ;
  assign n30786 = ~n30781 & n30785 ;
  assign n30787 = n26177 & n30675 ;
  assign n30788 = n22160 & ~n30658 ;
  assign n30789 = ~n30787 & n30788 ;
  assign n30790 = ~n21038 & ~n30789 ;
  assign n30791 = ~n30786 & n30790 ;
  assign n30792 = ~n30779 & n30791 ;
  assign n30793 = n20777 & ~n22160 ;
  assign n30794 = n30782 & n30793 ;
  assign n30795 = n30780 & n30793 ;
  assign n30796 = ~n30669 & n30795 ;
  assign n30797 = ~n30794 & ~n30796 ;
  assign n30798 = n20777 & n30658 ;
  assign n30799 = ~\pi0641  & ~n30658 ;
  assign n30800 = ~n22899 & ~n30799 ;
  assign n30801 = n26196 & n30674 ;
  assign n30802 = ~n22899 & n30801 ;
  assign n30803 = n23832 & n30802 ;
  assign n30804 = ~n30800 & ~n30803 ;
  assign n30805 = ~n30798 & n30804 ;
  assign n30806 = n30797 & n30805 ;
  assign n30807 = n20776 & ~n22160 ;
  assign n30808 = n30782 & n30807 ;
  assign n30809 = n30780 & n30807 ;
  assign n30810 = ~n30669 & n30809 ;
  assign n30811 = ~n30808 & ~n30810 ;
  assign n30812 = n20776 & n30658 ;
  assign n30813 = \pi0641  & ~n30658 ;
  assign n30814 = ~n22884 & ~n30813 ;
  assign n30815 = n26205 & n30674 ;
  assign n30816 = ~n22884 & n30815 ;
  assign n30817 = n23832 & n30816 ;
  assign n30818 = ~n30814 & ~n30817 ;
  assign n30819 = ~n30812 & n30818 ;
  assign n30820 = n30811 & n30819 ;
  assign n30821 = ~n30806 & ~n30820 ;
  assign n30822 = \pi0788  & n30821 ;
  assign n30823 = ~n21067 & ~n23856 ;
  assign n30824 = ~n30822 & n30823 ;
  assign n30825 = ~n30792 & n30824 ;
  assign n30826 = ~n24761 & ~n30825 ;
  assign n30827 = n30725 & n30826 ;
  assign n30828 = n30687 & ~n30827 ;
  assign n30829 = ~n30655 & ~n30828 ;
  assign n30830 = \pi0766  & n1689 ;
  assign n30831 = n20784 & n30830 ;
  assign n30832 = n22767 & n30831 ;
  assign n30833 = ~\pi0175  & ~n1689 ;
  assign n30834 = ~n30831 & ~n30833 ;
  assign n30835 = ~n20792 & ~n30834 ;
  assign n30836 = ~n30832 & n30835 ;
  assign n30837 = n20801 & ~n30836 ;
  assign n30838 = ~\pi1155  & ~n30833 ;
  assign n30839 = \pi0785  & n30838 ;
  assign n30840 = ~n30832 & n30839 ;
  assign n30841 = ~\pi0785  & ~n30833 ;
  assign n30842 = ~n30831 & n30841 ;
  assign n30843 = ~n20804 & ~n30842 ;
  assign n30844 = n29682 & n30843 ;
  assign n30845 = ~n30840 & n30844 ;
  assign n30846 = ~n30837 & n30845 ;
  assign n30847 = n20886 & ~n23880 ;
  assign n30848 = n30846 & n30847 ;
  assign n30849 = \pi0700  & n1689 ;
  assign n30850 = n20855 & n30849 ;
  assign n30851 = ~n30833 & ~n30850 ;
  assign n30852 = ~\pi0778  & ~n30851 ;
  assign n30853 = ~\pi0625  & \pi0700  ;
  assign n30854 = n1689 & n30853 ;
  assign n30855 = n20855 & n30854 ;
  assign n30856 = \pi1153  & n30855 ;
  assign n30857 = \pi1153  & ~n30833 ;
  assign n30858 = ~n30850 & n30857 ;
  assign n30859 = ~n30856 & ~n30858 ;
  assign n30860 = ~\pi1153  & ~n30833 ;
  assign n30861 = ~n30855 & n30860 ;
  assign n30862 = \pi0778  & ~n30861 ;
  assign n30863 = n30859 & n30862 ;
  assign n30864 = ~n30852 & ~n30863 ;
  assign n30865 = n26474 & ~n30864 ;
  assign n30866 = ~\pi0175  & \pi0788  ;
  assign n30867 = ~n1689 & n30866 ;
  assign n30868 = ~n20778 & n30867 ;
  assign n30869 = n20886 & n30868 ;
  assign n30870 = \pi0629  & ~n30869 ;
  assign n30871 = ~n30865 & n30870 ;
  assign n30872 = ~n30848 & n30871 ;
  assign n30873 = n20887 & ~n23880 ;
  assign n30874 = n30846 & n30873 ;
  assign n30875 = n26485 & ~n30864 ;
  assign n30876 = n20887 & n30868 ;
  assign n30877 = ~\pi0629  & ~n30876 ;
  assign n30878 = ~n30875 & n30877 ;
  assign n30879 = ~n30874 & n30878 ;
  assign n30880 = \pi0792  & ~n30879 ;
  assign n30881 = ~n30872 & n30880 ;
  assign n30882 = ~n21067 & ~n30881 ;
  assign n30883 = n26325 & ~n30864 ;
  assign n30884 = ~\pi0175  & ~\pi0647  ;
  assign n30885 = ~n1689 & n30884 ;
  assign n30886 = n20849 & ~n30885 ;
  assign n30887 = ~n30883 & n30886 ;
  assign n30888 = n26319 & ~n30864 ;
  assign n30889 = ~\pi0175  & \pi0647  ;
  assign n30890 = ~n1689 & n30889 ;
  assign n30891 = n20897 & ~n30890 ;
  assign n30892 = ~n30888 & n30891 ;
  assign n30893 = ~n30887 & ~n30892 ;
  assign n30894 = \pi0787  & ~n30893 ;
  assign n30895 = n30376 & n30846 ;
  assign n30896 = ~n20846 & n30868 ;
  assign n30897 = ~\pi0175  & \pi0792  ;
  assign n30898 = ~n1689 & n30897 ;
  assign n30899 = ~n20845 & n30898 ;
  assign n30900 = ~n24996 & ~n30899 ;
  assign n30901 = ~n30896 & n30900 ;
  assign n30902 = ~n30895 & n30901 ;
  assign n30903 = ~n24761 & ~n30902 ;
  assign n30904 = ~n30894 & n30903 ;
  assign n30905 = ~n30882 & n30904 ;
  assign n30906 = \pi0608  & ~n30861 ;
  assign n30907 = ~n30831 & n30857 ;
  assign n30908 = \pi0778  & ~n30907 ;
  assign n30909 = n26421 & ~n30851 ;
  assign n30910 = ~n30908 & ~n30909 ;
  assign n30911 = n30906 & ~n30910 ;
  assign n30912 = n26147 & ~n30851 ;
  assign n30913 = \pi0700  & ~n20784 ;
  assign n30914 = n22113 & n30913 ;
  assign n30915 = n30834 & ~n30914 ;
  assign n30916 = ~n30912 & ~n30915 ;
  assign n30917 = n30860 & ~n30916 ;
  assign n30918 = n26415 & n30859 ;
  assign n30919 = ~n30917 & n30918 ;
  assign n30920 = ~n30911 & ~n30919 ;
  assign n30921 = ~\pi1155  & ~n30852 ;
  assign n30922 = ~n30863 & n30921 ;
  assign n30923 = ~n20999 & ~n30922 ;
  assign n30924 = ~\pi0778  & ~n30915 ;
  assign n30925 = ~n30923 & ~n30924 ;
  assign n30926 = n30920 & n30925 ;
  assign n30927 = n29766 & ~n30852 ;
  assign n30928 = ~n30863 & n30927 ;
  assign n30929 = \pi1155  & ~n30836 ;
  assign n30930 = ~\pi0660  & ~n30929 ;
  assign n30931 = ~n30928 & n30930 ;
  assign n30932 = ~n30926 & n30931 ;
  assign n30933 = \pi0785  & ~n30932 ;
  assign n30934 = n29775 & n30843 ;
  assign n30935 = ~n30840 & n30934 ;
  assign n30936 = ~n30837 & n30935 ;
  assign n30937 = n29779 & ~n30864 ;
  assign n30938 = ~n30936 & ~n30937 ;
  assign n30939 = \pi0781  & ~n30938 ;
  assign n30940 = \pi1155  & ~n30852 ;
  assign n30941 = ~n30863 & n30940 ;
  assign n30942 = ~n21774 & ~n30941 ;
  assign n30943 = ~n30924 & ~n30942 ;
  assign n30944 = n30920 & n30943 ;
  assign n30945 = n26121 & ~n30852 ;
  assign n30946 = ~n30863 & n30945 ;
  assign n30947 = \pi0660  & ~n30838 ;
  assign n30948 = \pi0660  & n30831 ;
  assign n30949 = n22767 & n30948 ;
  assign n30950 = ~n30947 & ~n30949 ;
  assign n30951 = ~n30946 & ~n30950 ;
  assign n30952 = ~n30944 & n30951 ;
  assign n30953 = ~n30939 & ~n30952 ;
  assign n30954 = n30933 & n30953 ;
  assign n30955 = ~\pi0785  & ~n30924 ;
  assign n30956 = ~n30911 & n30955 ;
  assign n30957 = ~n30919 & n30956 ;
  assign n30958 = n21022 & ~n30957 ;
  assign n30959 = ~n30939 & ~n30958 ;
  assign n30960 = n29803 & ~n30959 ;
  assign n30961 = ~n30954 & n30960 ;
  assign n30962 = n29808 & n30843 ;
  assign n30963 = ~n30840 & n30962 ;
  assign n30964 = ~n30837 & n30963 ;
  assign n30965 = ~n20872 & ~n29814 ;
  assign n30966 = ~n20868 & n30965 ;
  assign n30967 = ~n30864 & n30966 ;
  assign n30968 = ~n30964 & ~n30967 ;
  assign n30969 = n29818 & ~n30968 ;
  assign n30970 = \pi0626  & ~n30846 ;
  assign n30971 = ~\pi0626  & ~n30833 ;
  assign n30972 = n20881 & ~n30971 ;
  assign n30973 = ~n30970 & n30972 ;
  assign n30974 = n26458 & ~n30864 ;
  assign n30975 = ~\pi0626  & ~n30846 ;
  assign n30976 = \pi0626  & ~n30833 ;
  assign n30977 = n20882 & ~n30976 ;
  assign n30978 = ~n30975 & n30977 ;
  assign n30979 = ~n30974 & ~n30978 ;
  assign n30980 = ~n30973 & n30979 ;
  assign n30981 = \pi0788  & ~n30980 ;
  assign n30982 = ~n30969 & ~n30981 ;
  assign n30983 = ~n30961 & n30982 ;
  assign n30984 = ~n23856 & n30904 ;
  assign n30985 = ~n30983 & n30984 ;
  assign n30986 = ~n30905 & ~n30985 ;
  assign n30987 = \pi1160  & ~n21088 ;
  assign n30988 = n30896 & n30987 ;
  assign n30989 = n30376 & n30987 ;
  assign n30990 = n30846 & n30989 ;
  assign n30991 = ~n30988 & ~n30990 ;
  assign n30992 = n23312 & ~n30991 ;
  assign n30993 = \pi1157  & ~n30885 ;
  assign n30994 = ~n30883 & n30993 ;
  assign n30995 = ~\pi1157  & ~n30890 ;
  assign n30996 = ~n30888 & n30995 ;
  assign n30997 = ~n30994 & ~n30996 ;
  assign n30998 = \pi0787  & ~n30997 ;
  assign n30999 = n26333 & ~n30864 ;
  assign n31000 = ~\pi0787  & ~n30999 ;
  assign n31001 = ~\pi1160  & ~n31000 ;
  assign n31002 = n23312 & n31001 ;
  assign n31003 = ~n30998 & n31002 ;
  assign n31004 = ~n30992 & ~n31003 ;
  assign n31005 = \pi0790  & ~n31004 ;
  assign n31006 = \pi1160  & ~n31000 ;
  assign n31007 = ~n30998 & n31006 ;
  assign n31008 = ~n23414 & n30833 ;
  assign n31009 = ~n24886 & n31008 ;
  assign n31010 = ~\pi1160  & ~n21088 ;
  assign n31011 = n30896 & n31010 ;
  assign n31012 = n30376 & n31010 ;
  assign n31013 = n30846 & n31012 ;
  assign n31014 = ~n31011 & ~n31013 ;
  assign n31015 = ~n31009 & n31014 ;
  assign n31016 = ~n31007 & n31015 ;
  assign n31017 = ~n23313 & ~n31008 ;
  assign n31018 = ~n20846 & ~n23313 ;
  assign n31019 = n23415 & n31018 ;
  assign n31020 = ~n31017 & ~n31019 ;
  assign n31021 = \pi0790  & n31020 ;
  assign n31022 = ~n31016 & n31021 ;
  assign n31023 = ~n31005 & ~n31022 ;
  assign n31024 = \pi0832  & n31023 ;
  assign n31025 = n30986 & n31024 ;
  assign n31026 = ~\pi0175  & \pi0766  ;
  assign n31027 = ~n21467 & n31026 ;
  assign n31028 = ~\pi0039  & n31026 ;
  assign n31029 = n21272 & n31028 ;
  assign n31030 = ~n31027 & ~n31029 ;
  assign n31031 = \pi0766  & n21484 ;
  assign n31032 = ~\pi0175  & n21743 ;
  assign n31033 = ~n31026 & ~n31032 ;
  assign n31034 = ~n31031 & n31033 ;
  assign n31035 = n31030 & ~n31034 ;
  assign n31036 = ~\pi0038  & ~n31035 ;
  assign n31037 = ~\pi0766  & ~n21731 ;
  assign n31038 = n21714 & n31037 ;
  assign n31039 = ~n21693 & n31038 ;
  assign n31040 = \pi0175  & ~n21543 ;
  assign n31041 = \pi0175  & n21562 ;
  assign n31042 = ~n21552 & n31041 ;
  assign n31043 = ~n31040 & ~n31042 ;
  assign n31044 = ~n21536 & ~n31043 ;
  assign n31045 = ~n31039 & ~n31044 ;
  assign n31046 = n9627 & ~n31045 ;
  assign n31047 = \pi0175  & ~n6861 ;
  assign n31048 = ~\pi0175  & ~n21757 ;
  assign n31049 = n8413 & n30831 ;
  assign n31050 = n1354 & n31049 ;
  assign n31051 = n1358 & n31050 ;
  assign n31052 = \pi0038  & ~n31051 ;
  assign n31053 = ~n31048 & n31052 ;
  assign n31054 = ~n31047 & ~n31053 ;
  assign n31055 = ~n31046 & n31054 ;
  assign n31056 = ~n31036 & n31055 ;
  assign n31057 = ~\pi0175  & ~n6861 ;
  assign n31058 = n22767 & ~n31057 ;
  assign n31059 = ~n31056 & n31058 ;
  assign n31060 = ~\pi0175  & n21768 ;
  assign n31061 = ~\pi0175  & n21770 ;
  assign n31062 = ~n21734 & n31061 ;
  assign n31063 = ~n31060 & ~n31062 ;
  assign n31064 = ~n22767 & n31063 ;
  assign n31065 = \pi0660  & ~n31064 ;
  assign n31066 = ~n31059 & n31065 ;
  assign n31067 = n29766 & ~n31066 ;
  assign n31068 = ~\pi0175  & ~\pi0700  ;
  assign n31069 = n21770 & n31068 ;
  assign n31070 = ~n21734 & n31069 ;
  assign n31071 = \pi0038  & n31068 ;
  assign n31072 = ~n22123 & n31071 ;
  assign n31073 = n6861 & ~n31072 ;
  assign n31074 = ~n31070 & n31073 ;
  assign n31075 = ~n31047 & ~n31074 ;
  assign n31076 = ~\pi0175  & ~n22017 ;
  assign n31077 = ~n21994 & n31076 ;
  assign n31078 = ~\pi0038  & ~\pi0175  ;
  assign n31079 = ~n22109 & ~n31078 ;
  assign n31080 = ~n31077 & ~n31079 ;
  assign n31081 = n22117 & ~n31048 ;
  assign n31082 = \pi0700  & ~n31047 ;
  assign n31083 = ~n31081 & n31082 ;
  assign n31084 = ~n31080 & n31083 ;
  assign n31085 = ~n31075 & ~n31084 ;
  assign n31086 = ~\pi0778  & n31085 ;
  assign n31087 = \pi0785  & n31086 ;
  assign n31088 = \pi0625  & ~n31085 ;
  assign n31089 = ~\pi0175  & ~\pi0625  ;
  assign n31090 = n21768 & n31089 ;
  assign n31091 = n21770 & n31089 ;
  assign n31092 = ~n21734 & n31091 ;
  assign n31093 = ~n31090 & ~n31092 ;
  assign n31094 = \pi1153  & n31093 ;
  assign n31095 = ~n31088 & n31094 ;
  assign n31096 = ~\pi0625  & ~n31085 ;
  assign n31097 = ~\pi0175  & \pi0625  ;
  assign n31098 = n21768 & n31097 ;
  assign n31099 = n21770 & n31097 ;
  assign n31100 = ~n21734 & n31099 ;
  assign n31101 = ~n31098 & ~n31100 ;
  assign n31102 = ~\pi1153  & n31101 ;
  assign n31103 = ~n31096 & n31102 ;
  assign n31104 = ~n31095 & ~n31103 ;
  assign n31105 = \pi0778  & \pi0785  ;
  assign n31106 = ~n31104 & n31105 ;
  assign n31107 = ~n31087 & ~n31106 ;
  assign n31108 = n31067 & ~n31107 ;
  assign n31109 = \pi0778  & n26121 ;
  assign n31110 = ~n31104 & n31109 ;
  assign n31111 = ~n22766 & ~n31066 ;
  assign n31112 = ~\pi0778  & n26121 ;
  assign n31113 = n31085 & n31112 ;
  assign n31114 = ~n31111 & ~n31113 ;
  assign n31115 = ~n31110 & n31114 ;
  assign n31116 = n22788 & ~n31057 ;
  assign n31117 = ~n31056 & n31116 ;
  assign n31118 = ~n22788 & n31063 ;
  assign n31119 = ~\pi0660  & ~n31118 ;
  assign n31120 = ~n31117 & n31119 ;
  assign n31121 = \pi0785  & ~n22787 ;
  assign n31122 = ~n31120 & n31121 ;
  assign n31123 = ~n31115 & n31122 ;
  assign n31124 = ~n31108 & ~n31123 ;
  assign n31125 = n26700 & ~n31124 ;
  assign n31126 = ~\pi1155  & ~n31066 ;
  assign n31127 = \pi0778  & ~n31104 ;
  assign n31128 = \pi0609  & ~n31086 ;
  assign n31129 = ~n31127 & n31128 ;
  assign n31130 = n31126 & ~n31129 ;
  assign n31131 = n21774 & ~n22787 ;
  assign n31132 = ~n31120 & n31131 ;
  assign n31133 = \pi0785  & ~n31132 ;
  assign n31134 = ~n31130 & n31133 ;
  assign n31135 = ~\pi0700  & ~n31053 ;
  assign n31136 = ~n31046 & n31135 ;
  assign n31137 = ~n31036 & n31136 ;
  assign n31138 = n6861 & ~n31137 ;
  assign n31139 = ~n22734 & ~n31089 ;
  assign n31140 = ~n31138 & ~n31139 ;
  assign n31141 = ~\pi0039  & ~\pi0175  ;
  assign n31142 = ~n22683 & n31141 ;
  assign n31143 = ~\pi0175  & ~n23548 ;
  assign n31144 = \pi0766  & ~n31143 ;
  assign n31145 = ~n31142 & n31144 ;
  assign n31146 = \pi0175  & ~n23558 ;
  assign n31147 = n23557 & n31146 ;
  assign n31148 = ~\pi0038  & ~n31147 ;
  assign n31149 = n31145 & n31148 ;
  assign n31150 = ~\pi0175  & ~n23568 ;
  assign n31151 = \pi0175  & n23575 ;
  assign n31152 = n23572 & n31151 ;
  assign n31153 = ~\pi0038  & ~\pi0766  ;
  assign n31154 = ~n31152 & n31153 ;
  assign n31155 = ~n31150 & n31154 ;
  assign n31156 = ~n31149 & ~n31155 ;
  assign n31157 = \pi0175  & \pi0603  ;
  assign n31158 = ~n20783 & n31157 ;
  assign n31159 = n30830 & n31158 ;
  assign n31160 = \pi0175  & ~n20784 ;
  assign n31161 = n22113 & n31160 ;
  assign n31162 = ~n31159 & ~n31161 ;
  assign n31163 = n26554 & ~n31162 ;
  assign n31164 = n1358 & n31163 ;
  assign n31165 = \pi0038  & ~n31164 ;
  assign n31166 = \pi0700  & ~n31165 ;
  assign n31167 = \pi0766  & ~n22317 ;
  assign n31168 = \pi0680  & ~n20854 ;
  assign n31169 = ~n20784 & n31168 ;
  assign n31170 = ~\pi0039  & ~n31169 ;
  assign n31171 = ~n31167 & n31170 ;
  assign n31172 = n21289 & n31171 ;
  assign n31173 = ~\pi0175  & \pi0700  ;
  assign n31174 = ~n31172 & n31173 ;
  assign n31175 = ~n31166 & ~n31174 ;
  assign n31176 = ~n31139 & ~n31175 ;
  assign n31177 = n31156 & n31176 ;
  assign n31178 = ~n31140 & ~n31177 ;
  assign n31179 = ~\pi1153  & ~n31057 ;
  assign n31180 = ~n31056 & n31179 ;
  assign n31181 = ~n24561 & ~n31180 ;
  assign n31182 = n31178 & ~n31181 ;
  assign n31183 = ~\pi0608  & ~n31094 ;
  assign n31184 = n22755 & ~n31085 ;
  assign n31185 = ~n31183 & ~n31184 ;
  assign n31186 = ~n31182 & ~n31185 ;
  assign n31187 = ~n22727 & ~n31097 ;
  assign n31188 = ~n31138 & ~n31187 ;
  assign n31189 = ~n31175 & ~n31187 ;
  assign n31190 = n31156 & n31189 ;
  assign n31191 = ~n31188 & ~n31190 ;
  assign n31192 = \pi1153  & ~n31057 ;
  assign n31193 = ~n31056 & n31192 ;
  assign n31194 = ~n24550 & ~n31193 ;
  assign n31195 = n31191 & ~n31194 ;
  assign n31196 = \pi0608  & ~n31102 ;
  assign n31197 = n22740 & ~n31085 ;
  assign n31198 = ~n31196 & ~n31197 ;
  assign n31199 = ~n31195 & ~n31198 ;
  assign n31200 = ~n31186 & ~n31199 ;
  assign n31201 = \pi0778  & ~n31200 ;
  assign n31202 = ~n31134 & ~n31201 ;
  assign n31203 = ~\pi0175  & ~\pi0778  ;
  assign n31204 = ~n23622 & ~n31203 ;
  assign n31205 = ~n31138 & ~n31204 ;
  assign n31206 = ~n31175 & ~n31204 ;
  assign n31207 = n31156 & n31206 ;
  assign n31208 = ~n31205 & ~n31207 ;
  assign n31209 = n26700 & n31208 ;
  assign n31210 = n31202 & n31209 ;
  assign n31211 = ~n31125 & ~n31210 ;
  assign n31212 = n26065 & ~n31104 ;
  assign n31213 = n26739 & n31085 ;
  assign n31214 = ~n23885 & n31063 ;
  assign n31215 = ~\pi0628  & ~n31214 ;
  assign n31216 = ~n31213 & n31215 ;
  assign n31217 = ~n31212 & n31216 ;
  assign n31218 = ~\pi0175  & \pi0628  ;
  assign n31219 = n21768 & n31218 ;
  assign n31220 = n21770 & n31218 ;
  assign n31221 = ~n21734 & n31220 ;
  assign n31222 = ~n31219 & ~n31221 ;
  assign n31223 = n20844 & n31222 ;
  assign n31224 = ~n31217 & n31223 ;
  assign n31225 = ~\pi0175  & ~n20811 ;
  assign n31226 = n21768 & n31225 ;
  assign n31227 = n21770 & n31225 ;
  assign n31228 = ~n21734 & n31227 ;
  assign n31229 = ~n31226 & ~n31228 ;
  assign n31230 = n23424 & ~n31229 ;
  assign n31231 = n21777 & ~n31057 ;
  assign n31232 = ~n31056 & n31231 ;
  assign n31233 = ~n21777 & n31063 ;
  assign n31234 = n20811 & ~n31233 ;
  assign n31235 = n23424 & n31234 ;
  assign n31236 = ~n31232 & n31235 ;
  assign n31237 = ~n31230 & ~n31236 ;
  assign n31238 = ~\pi0781  & ~n31233 ;
  assign n31239 = ~n23423 & n31238 ;
  assign n31240 = ~n31232 & n31239 ;
  assign n31241 = n23423 & ~n31063 ;
  assign n31242 = ~n31240 & ~n31241 ;
  assign n31243 = n31237 & n31242 ;
  assign n31244 = ~n23880 & ~n31243 ;
  assign n31245 = n23880 & ~n31063 ;
  assign n31246 = n24691 & ~n31245 ;
  assign n31247 = ~n31244 & n31246 ;
  assign n31248 = \pi0628  & ~n31214 ;
  assign n31249 = ~n31213 & n31248 ;
  assign n31250 = ~n31212 & n31249 ;
  assign n31251 = ~\pi0175  & ~\pi0628  ;
  assign n31252 = n21768 & n31251 ;
  assign n31253 = n21770 & n31251 ;
  assign n31254 = ~n21734 & n31253 ;
  assign n31255 = ~n31252 & ~n31254 ;
  assign n31256 = n20843 & n31255 ;
  assign n31257 = ~n31250 & n31256 ;
  assign n31258 = ~n31247 & ~n31257 ;
  assign n31259 = ~n31224 & n31258 ;
  assign n31260 = \pi0792  & ~n31259 ;
  assign n31261 = ~n31232 & n31234 ;
  assign n31262 = n22155 & n31229 ;
  assign n31263 = ~n31261 & n31262 ;
  assign n31264 = ~n22147 & ~n31086 ;
  assign n31265 = n22147 & ~n31063 ;
  assign n31266 = n30053 & ~n31265 ;
  assign n31267 = ~n31264 & n31266 ;
  assign n31268 = \pi0778  & n31266 ;
  assign n31269 = ~n31104 & n31268 ;
  assign n31270 = ~n31267 & ~n31269 ;
  assign n31271 = ~n31263 & n31270 ;
  assign n31272 = ~n21034 & ~n31271 ;
  assign n31273 = n30780 & ~n31104 ;
  assign n31274 = ~\pi0778  & n23380 ;
  assign n31275 = n31085 & n31274 ;
  assign n31276 = ~n23380 & n31063 ;
  assign n31277 = ~n31275 & ~n31276 ;
  assign n31278 = ~n31273 & n31277 ;
  assign n31279 = \pi0789  & ~\pi1159  ;
  assign n31280 = n21029 & n31279 ;
  assign n31281 = \pi0789  & \pi1159  ;
  assign n31282 = n21028 & n31281 ;
  assign n31283 = ~n31280 & ~n31282 ;
  assign n31284 = ~n31278 & ~n31283 ;
  assign n31285 = n23683 & ~n31229 ;
  assign n31286 = n23683 & n31234 ;
  assign n31287 = ~n31232 & n31286 ;
  assign n31288 = ~n31285 & ~n31287 ;
  assign n31289 = n21032 & n31238 ;
  assign n31290 = ~n31232 & n31289 ;
  assign n31291 = ~n21032 & ~n31063 ;
  assign n31292 = ~n20876 & ~n31291 ;
  assign n31293 = \pi0789  & n31292 ;
  assign n31294 = ~n31290 & n31293 ;
  assign n31295 = n31288 & n31294 ;
  assign n31296 = ~n21038 & ~n31295 ;
  assign n31297 = ~n31284 & n31296 ;
  assign n31298 = ~n31272 & n31297 ;
  assign n31299 = ~n31260 & n31298 ;
  assign n31300 = n31211 & n31299 ;
  assign n31301 = n23380 & n23838 ;
  assign n31302 = n20951 & ~n31063 ;
  assign n31303 = ~n31301 & ~n31302 ;
  assign n31304 = ~n31275 & ~n31303 ;
  assign n31305 = ~n31273 & n31304 ;
  assign n31306 = n20951 & n22160 ;
  assign n31307 = ~n31063 & n31306 ;
  assign n31308 = ~n23856 & ~n31307 ;
  assign n31309 = ~n31305 & n31308 ;
  assign n31310 = \pi0626  & ~n31241 ;
  assign n31311 = ~n31240 & n31310 ;
  assign n31312 = n31237 & n31311 ;
  assign n31313 = ~\pi0626  & n31063 ;
  assign n31314 = n20881 & ~n31313 ;
  assign n31315 = ~n31312 & n31314 ;
  assign n31316 = ~\pi0626  & ~n31241 ;
  assign n31317 = ~n31240 & n31316 ;
  assign n31318 = n31237 & n31317 ;
  assign n31319 = \pi0626  & n31063 ;
  assign n31320 = n20882 & ~n31319 ;
  assign n31321 = ~n31318 & n31320 ;
  assign n31322 = ~n31315 & ~n31321 ;
  assign n31323 = n31309 & n31322 ;
  assign n31324 = ~n26803 & ~n31323 ;
  assign n31325 = ~n31260 & n31324 ;
  assign n31326 = ~n21067 & ~n31325 ;
  assign n31327 = ~n31300 & n31326 ;
  assign n31328 = ~n20846 & n31245 ;
  assign n31329 = n30376 & ~n31243 ;
  assign n31330 = ~n31328 & ~n31329 ;
  assign n31331 = n20846 & ~n31063 ;
  assign n31332 = ~n20910 & ~n31331 ;
  assign n31333 = n31330 & n31332 ;
  assign n31334 = n21768 & n30889 ;
  assign n31335 = n21770 & n30889 ;
  assign n31336 = ~n21734 & n31335 ;
  assign n31337 = ~n31334 & ~n31336 ;
  assign n31338 = \pi0647  & n20897 ;
  assign n31339 = n31337 & n31338 ;
  assign n31340 = ~n23907 & ~n31214 ;
  assign n31341 = ~n31213 & n31340 ;
  assign n31342 = ~n31212 & n31341 ;
  assign n31343 = n23907 & ~n31063 ;
  assign n31344 = n20897 & n31337 ;
  assign n31345 = ~n31343 & n31344 ;
  assign n31346 = ~n31342 & n31345 ;
  assign n31347 = ~n31339 & ~n31346 ;
  assign n31348 = n21768 & n30884 ;
  assign n31349 = n21770 & n30884 ;
  assign n31350 = ~n21734 & n31349 ;
  assign n31351 = ~n31348 & ~n31350 ;
  assign n31352 = n20850 & n31351 ;
  assign n31353 = n20849 & n31351 ;
  assign n31354 = ~n31343 & n31353 ;
  assign n31355 = ~n31342 & n31354 ;
  assign n31356 = ~n31352 & ~n31355 ;
  assign n31357 = n31347 & n31356 ;
  assign n31358 = ~n31333 & n31357 ;
  assign n31359 = \pi0787  & ~n31358 ;
  assign n31360 = ~\pi0175  & \pi0644  ;
  assign n31361 = n21768 & n31360 ;
  assign n31362 = n21770 & n31360 ;
  assign n31363 = ~n21734 & n31362 ;
  assign n31364 = ~n31361 & ~n31363 ;
  assign n31365 = n23939 & n31364 ;
  assign n31366 = \pi0715  & n31364 ;
  assign n31367 = n21092 & ~n23880 ;
  assign n31368 = ~\pi0175  & ~n31367 ;
  assign n31369 = n21768 & n31368 ;
  assign n31370 = n21770 & n31368 ;
  assign n31371 = ~n21734 & n31370 ;
  assign n31372 = ~n31369 & ~n31371 ;
  assign n31373 = n31366 & n31372 ;
  assign n31374 = ~n31365 & ~n31373 ;
  assign n31375 = ~n31365 & n31367 ;
  assign n31376 = ~n31243 & n31375 ;
  assign n31377 = ~n31374 & ~n31376 ;
  assign n31378 = ~\pi0644  & ~\pi1160  ;
  assign n31379 = ~n31377 & n31378 ;
  assign n31380 = ~\pi0715  & n31372 ;
  assign n31381 = ~n23958 & ~n31380 ;
  assign n31382 = ~n23958 & n31367 ;
  assign n31383 = ~n31243 & n31382 ;
  assign n31384 = ~n31381 & ~n31383 ;
  assign n31385 = n26824 & ~n31384 ;
  assign n31386 = \pi0790  & ~n31385 ;
  assign n31387 = ~n31379 & n31386 ;
  assign n31388 = n9948 & ~n31387 ;
  assign n31389 = ~n31359 & n31388 ;
  assign n31390 = ~n31327 & n31389 ;
  assign n31391 = n23942 & n31063 ;
  assign n31392 = \pi0644  & ~n31391 ;
  assign n31393 = ~\pi0715  & ~n31392 ;
  assign n31394 = ~n23942 & ~n31343 ;
  assign n31395 = ~\pi0715  & n31394 ;
  assign n31396 = ~n31342 & n31395 ;
  assign n31397 = ~n31393 & ~n31396 ;
  assign n31398 = ~\pi1160  & ~n31377 ;
  assign n31399 = n31397 & n31398 ;
  assign n31400 = n9948 & n31399 ;
  assign n31401 = ~\pi0175  & ~\pi0644  ;
  assign n31402 = n21768 & n31401 ;
  assign n31403 = n21770 & n31401 ;
  assign n31404 = ~n21734 & n31403 ;
  assign n31405 = ~n31402 & ~n31404 ;
  assign n31406 = n31384 & n31405 ;
  assign n31407 = ~\pi0644  & ~n31391 ;
  assign n31408 = \pi0715  & ~n31407 ;
  assign n31409 = \pi0715  & n31394 ;
  assign n31410 = ~n31342 & n31409 ;
  assign n31411 = ~n31408 & ~n31410 ;
  assign n31412 = ~n31406 & n31411 ;
  assign n31413 = \pi1160  & n9948 ;
  assign n31414 = n31412 & n31413 ;
  assign n31415 = ~n31400 & ~n31414 ;
  assign n31416 = \pi0790  & ~n31415 ;
  assign n31417 = \pi0175  & ~\pi0832  ;
  assign n31418 = ~n21132 & ~n31417 ;
  assign n31419 = ~n31416 & ~n31418 ;
  assign n31420 = ~n31390 & n31419 ;
  assign n31421 = ~n31025 & ~n31420 ;
  assign n31422 = ~\pi0704  & n1689 ;
  assign n31423 = n20855 & n31422 ;
  assign n31424 = ~n20861 & n31423 ;
  assign n31425 = ~\pi0176  & ~n1689 ;
  assign n31426 = ~n31424 & ~n31425 ;
  assign n31427 = n20879 & ~n31426 ;
  assign n31428 = n20938 & n31427 ;
  assign n31429 = n29714 & ~n31428 ;
  assign n31430 = ~n21032 & ~n31425 ;
  assign n31431 = \pi0789  & n31430 ;
  assign n31432 = n23423 & ~n31431 ;
  assign n31433 = ~\pi0742  & n1689 ;
  assign n31434 = n20784 & n31433 ;
  assign n31435 = ~n31425 & ~n31434 ;
  assign n31436 = n20794 & ~n31435 ;
  assign n31437 = n20796 & ~n31436 ;
  assign n31438 = n20799 & ~n31435 ;
  assign n31439 = n20801 & ~n31438 ;
  assign n31440 = ~n31437 & ~n31439 ;
  assign n31441 = ~\pi0785  & ~n31425 ;
  assign n31442 = ~n31434 & n31441 ;
  assign n31443 = ~n20804 & ~n31442 ;
  assign n31444 = ~n20812 & n31443 ;
  assign n31445 = ~n31431 & n31444 ;
  assign n31446 = n31440 & n31445 ;
  assign n31447 = ~n31432 & ~n31446 ;
  assign n31448 = ~n23880 & ~n31447 ;
  assign n31449 = n21077 & n31427 ;
  assign n31450 = n29709 & ~n31449 ;
  assign n31451 = \pi0792  & ~n31450 ;
  assign n31452 = n31448 & n31451 ;
  assign n31453 = ~\pi0176  & \pi0788  ;
  assign n31454 = ~n1689 & n31453 ;
  assign n31455 = ~n20778 & n31454 ;
  assign n31456 = \pi0629  & ~n31455 ;
  assign n31457 = ~n31428 & n31456 ;
  assign n31458 = ~\pi0629  & ~n31455 ;
  assign n31459 = ~n31449 & n31458 ;
  assign n31460 = ~n31457 & ~n31459 ;
  assign n31461 = n31451 & n31460 ;
  assign n31462 = ~n31452 & ~n31461 ;
  assign n31463 = ~n31429 & ~n31462 ;
  assign n31464 = ~n21067 & ~n31463 ;
  assign n31465 = ~\pi0176  & \pi0792  ;
  assign n31466 = ~n1689 & n31465 ;
  assign n31467 = ~n20845 & n31466 ;
  assign n31468 = ~n20910 & ~n31467 ;
  assign n31469 = n20846 & n31468 ;
  assign n31470 = n20895 & n31427 ;
  assign n31471 = ~\pi0176  & \pi0647  ;
  assign n31472 = ~n1689 & n31471 ;
  assign n31473 = n20897 & ~n31472 ;
  assign n31474 = ~n31470 & n31473 ;
  assign n31475 = ~\pi0176  & ~\pi0647  ;
  assign n31476 = ~n1689 & n31475 ;
  assign n31477 = n20849 & ~n31476 ;
  assign n31478 = ~n24761 & ~n31477 ;
  assign n31479 = ~n24761 & n24830 ;
  assign n31480 = n31427 & n31479 ;
  assign n31481 = ~n31478 & ~n31480 ;
  assign n31482 = ~n31474 & ~n31481 ;
  assign n31483 = ~n31469 & n31482 ;
  assign n31484 = ~n29722 & ~n31483 ;
  assign n31485 = ~n31455 & n31468 ;
  assign n31486 = ~n29722 & n31485 ;
  assign n31487 = ~n31448 & n31486 ;
  assign n31488 = ~n31484 & ~n31487 ;
  assign n31489 = ~n31464 & n31488 ;
  assign n31490 = ~\pi0626  & n31447 ;
  assign n31491 = \pi0626  & ~n31425 ;
  assign n31492 = n20882 & ~n31491 ;
  assign n31493 = ~n31490 & n31492 ;
  assign n31494 = n23170 & ~n31426 ;
  assign n31495 = ~\pi0626  & ~n31425 ;
  assign n31496 = n20881 & ~n31495 ;
  assign n31497 = ~n31494 & ~n31496 ;
  assign n31498 = \pi0626  & ~n31494 ;
  assign n31499 = n31447 & n31498 ;
  assign n31500 = ~n31497 & ~n31499 ;
  assign n31501 = ~n31493 & ~n31500 ;
  assign n31502 = \pi0788  & ~n31501 ;
  assign n31503 = ~\pi0704  & ~n20784 ;
  assign n31504 = ~\pi0704  & ~n20790 ;
  assign n31505 = n20789 & n31504 ;
  assign n31506 = ~n31503 & ~n31505 ;
  assign n31507 = n24915 & ~n31506 ;
  assign n31508 = \pi0603  & ~\pi0742  ;
  assign n31509 = ~n20783 & n31508 ;
  assign n31510 = ~n20985 & n31509 ;
  assign n31511 = ~n31425 & ~n31510 ;
  assign n31512 = ~n31507 & n31511 ;
  assign n31513 = \pi0176  & ~n1689 ;
  assign n31514 = ~\pi0609  & ~n31513 ;
  assign n31515 = ~n31512 & n31514 ;
  assign n31516 = ~\pi1155  & ~n31425 ;
  assign n31517 = ~n31424 & n31516 ;
  assign n31518 = ~n20999 & ~n31517 ;
  assign n31519 = ~n31515 & ~n31518 ;
  assign n31520 = \pi1155  & ~n31438 ;
  assign n31521 = ~\pi0660  & ~n31520 ;
  assign n31522 = ~n31519 & n31521 ;
  assign n31523 = ~n21007 & ~n31437 ;
  assign n31524 = \pi0609  & ~n31513 ;
  assign n31525 = ~n31512 & n31524 ;
  assign n31526 = \pi1155  & ~n31425 ;
  assign n31527 = ~n31424 & n31526 ;
  assign n31528 = ~n21774 & ~n31527 ;
  assign n31529 = \pi0785  & ~n31528 ;
  assign n31530 = ~n31525 & n31529 ;
  assign n31531 = n31523 & ~n31530 ;
  assign n31532 = ~n31522 & ~n31531 ;
  assign n31533 = ~n31512 & ~n31513 ;
  assign n31534 = ~\pi0785  & ~n31533 ;
  assign n31535 = n21022 & ~n31534 ;
  assign n31536 = ~n31532 & n31535 ;
  assign n31537 = n20964 & n31443 ;
  assign n31538 = n31440 & n31537 ;
  assign n31539 = \pi0627  & ~n31425 ;
  assign n31540 = ~n31424 & n31539 ;
  assign n31541 = ~n20968 & ~n31540 ;
  assign n31542 = ~n31538 & ~n31541 ;
  assign n31543 = ~\pi0627  & ~n31425 ;
  assign n31544 = ~n31424 & n31543 ;
  assign n31545 = ~n20978 & ~n31544 ;
  assign n31546 = \pi0781  & n31545 ;
  assign n31547 = n20974 & n31443 ;
  assign n31548 = \pi0781  & n31547 ;
  assign n31549 = n31440 & n31548 ;
  assign n31550 = ~n31546 & ~n31549 ;
  assign n31551 = ~n31542 & ~n31550 ;
  assign n31552 = ~n21034 & ~n31551 ;
  assign n31553 = ~n31536 & n31552 ;
  assign n31554 = n21050 & ~n31425 ;
  assign n31555 = ~n31424 & n31554 ;
  assign n31556 = ~n21051 & ~n31555 ;
  assign n31557 = ~n20876 & n31430 ;
  assign n31558 = ~n21038 & ~n31557 ;
  assign n31559 = n31556 & n31558 ;
  assign n31560 = ~n23177 & ~n31559 ;
  assign n31561 = n31440 & n31444 ;
  assign n31562 = ~n23177 & n24969 ;
  assign n31563 = ~n31561 & n31562 ;
  assign n31564 = ~n31560 & ~n31563 ;
  assign n31565 = ~n31553 & n31564 ;
  assign n31566 = ~n31502 & ~n31565 ;
  assign n31567 = ~n23856 & n31488 ;
  assign n31568 = ~n31566 & n31567 ;
  assign n31569 = ~n31489 & ~n31568 ;
  assign n31570 = n24830 & n31427 ;
  assign n31571 = \pi1157  & ~n31476 ;
  assign n31572 = ~n31570 & n31571 ;
  assign n31573 = ~\pi1157  & ~n31472 ;
  assign n31574 = ~n31470 & n31573 ;
  assign n31575 = ~n31572 & ~n31574 ;
  assign n31576 = \pi0787  & ~n31575 ;
  assign n31577 = n24844 & n31427 ;
  assign n31578 = ~n24843 & ~n31577 ;
  assign n31579 = ~n31576 & ~n31578 ;
  assign n31580 = ~n20846 & n31010 ;
  assign n31581 = n31455 & n31580 ;
  assign n31582 = ~n23880 & n31580 ;
  assign n31583 = ~n31447 & n31582 ;
  assign n31584 = ~n31581 & ~n31583 ;
  assign n31585 = ~n31579 & n31584 ;
  assign n31586 = n23313 & ~n31585 ;
  assign n31587 = \pi0790  & n31586 ;
  assign n31588 = ~n20846 & n30987 ;
  assign n31589 = n31455 & n31588 ;
  assign n31590 = ~n23880 & n31588 ;
  assign n31591 = ~n31447 & n31590 ;
  assign n31592 = ~n31589 & ~n31591 ;
  assign n31593 = ~n23414 & n31425 ;
  assign n31594 = ~n24886 & n31593 ;
  assign n31595 = n20891 & n31427 ;
  assign n31596 = ~\pi0787  & ~n31595 ;
  assign n31597 = ~\pi1160  & ~n31596 ;
  assign n31598 = ~n31576 & n31597 ;
  assign n31599 = ~n31594 & ~n31598 ;
  assign n31600 = n31592 & n31599 ;
  assign n31601 = ~n23312 & ~n31593 ;
  assign n31602 = ~n20846 & ~n23312 ;
  assign n31603 = n23415 & n31602 ;
  assign n31604 = ~n31601 & ~n31603 ;
  assign n31605 = \pi0790  & n31604 ;
  assign n31606 = ~n31600 & n31605 ;
  assign n31607 = ~n31587 & ~n31606 ;
  assign n31608 = \pi0832  & n31607 ;
  assign n31609 = n31569 & n31608 ;
  assign n31610 = \pi0176  & ~\pi0832  ;
  assign n31611 = ~n21132 & ~n31610 ;
  assign n31612 = ~n31609 & n31611 ;
  assign n31613 = ~\pi0176  & n21770 ;
  assign n31614 = ~n21734 & n31613 ;
  assign n31615 = ~\pi0176  & n21768 ;
  assign n31616 = ~n31614 & ~n31615 ;
  assign n31617 = n23942 & n31616 ;
  assign n31618 = \pi0644  & ~n31617 ;
  assign n31619 = ~\pi0715  & ~n31618 ;
  assign n31620 = ~\pi0176  & n22124 ;
  assign n31621 = ~n31614 & ~n31620 ;
  assign n31622 = \pi0704  & n6861 ;
  assign n31623 = n31621 & n31622 ;
  assign n31624 = ~\pi0038  & ~n22017 ;
  assign n31625 = ~n21994 & n31624 ;
  assign n31626 = ~\pi0176  & ~n25669 ;
  assign n31627 = ~n31625 & n31626 ;
  assign n31628 = ~\pi0704  & n6861 ;
  assign n31629 = n31627 & n31628 ;
  assign n31630 = ~n31623 & ~n31629 ;
  assign n31631 = n6861 & ~n22117 ;
  assign n31632 = ~n22109 & n31631 ;
  assign n31633 = \pi0176  & ~n31632 ;
  assign n31634 = \pi0625  & ~n31633 ;
  assign n31635 = n31630 & n31634 ;
  assign n31636 = ~\pi0176  & ~\pi0625  ;
  assign n31637 = n21768 & n31636 ;
  assign n31638 = n21770 & n31636 ;
  assign n31639 = ~n21734 & n31638 ;
  assign n31640 = ~n31637 & ~n31639 ;
  assign n31641 = \pi1153  & n31640 ;
  assign n31642 = ~n31635 & n31641 ;
  assign n31643 = ~\pi0625  & ~n31633 ;
  assign n31644 = n31630 & n31643 ;
  assign n31645 = ~\pi0176  & \pi0625  ;
  assign n31646 = n21768 & n31645 ;
  assign n31647 = n21770 & n31645 ;
  assign n31648 = ~n21734 & n31647 ;
  assign n31649 = ~n31646 & ~n31648 ;
  assign n31650 = ~\pi1153  & n31649 ;
  assign n31651 = ~n31644 & n31650 ;
  assign n31652 = ~n31642 & ~n31651 ;
  assign n31653 = n26065 & ~n31652 ;
  assign n31654 = n31630 & ~n31633 ;
  assign n31655 = n26739 & ~n31654 ;
  assign n31656 = ~n23885 & n31616 ;
  assign n31657 = ~n23907 & ~n31656 ;
  assign n31658 = ~n31655 & n31657 ;
  assign n31659 = ~n31653 & n31658 ;
  assign n31660 = n23907 & ~n31616 ;
  assign n31661 = ~n23942 & ~n31660 ;
  assign n31662 = ~\pi0715  & n31661 ;
  assign n31663 = ~n31659 & n31662 ;
  assign n31664 = ~n31619 & ~n31663 ;
  assign n31665 = ~\pi0176  & \pi0644  ;
  assign n31666 = n21768 & n31665 ;
  assign n31667 = n21770 & n31665 ;
  assign n31668 = ~n21734 & n31667 ;
  assign n31669 = ~n31666 & ~n31668 ;
  assign n31670 = n23939 & n31669 ;
  assign n31671 = \pi0715  & n31669 ;
  assign n31672 = ~\pi0176  & ~n31367 ;
  assign n31673 = n21768 & n31672 ;
  assign n31674 = n21770 & n31672 ;
  assign n31675 = ~n21734 & n31674 ;
  assign n31676 = ~n31673 & ~n31675 ;
  assign n31677 = n31671 & n31676 ;
  assign n31678 = ~n31670 & ~n31677 ;
  assign n31679 = ~\pi0176  & ~n20811 ;
  assign n31680 = n21768 & n31679 ;
  assign n31681 = n21770 & n31679 ;
  assign n31682 = ~n21734 & n31681 ;
  assign n31683 = ~n31680 & ~n31682 ;
  assign n31684 = ~n21777 & n31616 ;
  assign n31685 = n20811 & ~n31684 ;
  assign n31686 = n31683 & ~n31685 ;
  assign n31687 = ~\pi0176  & ~n25033 ;
  assign n31688 = ~n25028 & n31687 ;
  assign n31689 = \pi0176  & ~n25040 ;
  assign n31690 = ~n25024 & n31689 ;
  assign n31691 = ~n31688 & ~n31690 ;
  assign n31692 = ~\pi0742  & n6861 ;
  assign n31693 = ~n31691 & n31692 ;
  assign n31694 = \pi0176  & ~n6861 ;
  assign n31695 = \pi0742  & n1289 ;
  assign n31696 = n1287 & n31695 ;
  assign n31697 = n31621 & n31696 ;
  assign n31698 = ~n31694 & ~n31697 ;
  assign n31699 = ~n31693 & n31698 ;
  assign n31700 = n21777 & n31683 ;
  assign n31701 = ~n31699 & n31700 ;
  assign n31702 = ~n31686 & ~n31701 ;
  assign n31703 = n23424 & n31702 ;
  assign n31704 = n21777 & ~n31699 ;
  assign n31705 = ~\pi0781  & ~n31684 ;
  assign n31706 = ~n23423 & n31705 ;
  assign n31707 = ~n31704 & n31706 ;
  assign n31708 = n23423 & ~n31616 ;
  assign n31709 = ~n31707 & ~n31708 ;
  assign n31710 = ~n31703 & n31709 ;
  assign n31711 = n31367 & ~n31670 ;
  assign n31712 = ~n31710 & n31711 ;
  assign n31713 = ~n31678 & ~n31712 ;
  assign n31714 = ~\pi1160  & ~n31713 ;
  assign n31715 = n31664 & n31714 ;
  assign n31716 = ~\pi0715  & n31676 ;
  assign n31717 = ~n23958 & ~n31716 ;
  assign n31718 = n31382 & ~n31710 ;
  assign n31719 = ~n31717 & ~n31718 ;
  assign n31720 = ~\pi0176  & ~\pi0644  ;
  assign n31721 = n21768 & n31720 ;
  assign n31722 = n21770 & n31720 ;
  assign n31723 = ~n21734 & n31722 ;
  assign n31724 = ~n31721 & ~n31723 ;
  assign n31725 = n31719 & n31724 ;
  assign n31726 = ~\pi0644  & ~n31617 ;
  assign n31727 = \pi0715  & ~n31726 ;
  assign n31728 = \pi0715  & n31661 ;
  assign n31729 = ~n31659 & n31728 ;
  assign n31730 = ~n31727 & ~n31729 ;
  assign n31731 = \pi1160  & n31730 ;
  assign n31732 = ~n31725 & n31731 ;
  assign n31733 = ~n31715 & ~n31732 ;
  assign n31734 = \pi0790  & ~n31733 ;
  assign n31735 = ~n31609 & n31734 ;
  assign n31736 = \pi0038  & \pi0176  ;
  assign n31737 = ~n22708 & n31736 ;
  assign n31738 = ~\pi0038  & \pi0176  ;
  assign n31739 = ~n31737 & ~n31738 ;
  assign n31740 = ~n23558 & ~n31737 ;
  assign n31741 = n23557 & n31740 ;
  assign n31742 = ~n31739 & ~n31741 ;
  assign n31743 = ~\pi0176  & n23548 ;
  assign n31744 = ~n25191 & n31743 ;
  assign n31745 = ~n25190 & n31744 ;
  assign n31746 = ~\pi0704  & ~\pi0742  ;
  assign n31747 = ~n31745 & n31746 ;
  assign n31748 = ~n31742 & n31747 ;
  assign n31749 = ~n25204 & ~n25209 ;
  assign n31750 = ~\pi0176  & ~n31749 ;
  assign n31751 = \pi0176  & ~n25217 ;
  assign n31752 = \pi0742  & ~n31751 ;
  assign n31753 = ~\pi0038  & n23575 ;
  assign n31754 = \pi0742  & n31753 ;
  assign n31755 = n23572 & n31754 ;
  assign n31756 = ~n31752 & ~n31755 ;
  assign n31757 = ~\pi0704  & ~n31756 ;
  assign n31758 = ~n31750 & n31757 ;
  assign n31759 = ~n31748 & ~n31758 ;
  assign n31760 = \pi0742  & n31621 ;
  assign n31761 = \pi0704  & \pi0742  ;
  assign n31762 = \pi0704  & ~n31690 ;
  assign n31763 = ~n31688 & n31762 ;
  assign n31764 = ~n31761 & ~n31763 ;
  assign n31765 = ~n31760 & ~n31764 ;
  assign n31766 = n6861 & ~n31765 ;
  assign n31767 = n31759 & n31766 ;
  assign n31768 = ~n22734 & ~n31636 ;
  assign n31769 = ~n31767 & ~n31768 ;
  assign n31770 = ~n22727 & ~n31645 ;
  assign n31771 = ~n31697 & ~n31770 ;
  assign n31772 = ~n31693 & n31771 ;
  assign n31773 = ~\pi1153  & ~n31772 ;
  assign n31774 = ~n31769 & n31773 ;
  assign n31775 = ~\pi0608  & ~n31642 ;
  assign n31776 = ~n31774 & n31775 ;
  assign n31777 = ~n31767 & ~n31770 ;
  assign n31778 = ~n31697 & ~n31768 ;
  assign n31779 = ~n31693 & n31778 ;
  assign n31780 = \pi1153  & ~n31779 ;
  assign n31781 = ~n31777 & n31780 ;
  assign n31782 = \pi0608  & ~n31651 ;
  assign n31783 = ~n31781 & n31782 ;
  assign n31784 = ~n31776 & ~n31783 ;
  assign n31785 = n23638 & ~n31784 ;
  assign n31786 = \pi0778  & ~n31652 ;
  assign n31787 = ~\pi0609  & ~n31633 ;
  assign n31788 = n31630 & n31787 ;
  assign n31789 = ~n23613 & ~n31788 ;
  assign n31790 = ~n31786 & ~n31789 ;
  assign n31791 = ~\pi0176  & ~\pi0778  ;
  assign n31792 = ~n23622 & ~n31791 ;
  assign n31793 = \pi0609  & ~n31792 ;
  assign n31794 = ~n31767 & n31793 ;
  assign n31795 = ~n22788 & n31616 ;
  assign n31796 = ~\pi0660  & ~n31795 ;
  assign n31797 = \pi1155  & ~n31796 ;
  assign n31798 = \pi1155  & n22788 ;
  assign n31799 = ~n31699 & n31798 ;
  assign n31800 = ~n31797 & ~n31799 ;
  assign n31801 = ~n31794 & ~n31800 ;
  assign n31802 = ~n31790 & n31801 ;
  assign n31803 = ~n31785 & n31802 ;
  assign n31804 = n23613 & ~n31784 ;
  assign n31805 = \pi0609  & ~n31633 ;
  assign n31806 = n31630 & n31805 ;
  assign n31807 = ~n23638 & ~n31806 ;
  assign n31808 = ~n31786 & ~n31807 ;
  assign n31809 = ~n22767 & n31616 ;
  assign n31810 = \pi0660  & ~n31809 ;
  assign n31811 = ~\pi1155  & ~n31810 ;
  assign n31812 = ~\pi1155  & n22767 ;
  assign n31813 = ~n31699 & n31812 ;
  assign n31814 = ~n31811 & ~n31813 ;
  assign n31815 = ~\pi0609  & ~n31792 ;
  assign n31816 = ~n31767 & n31815 ;
  assign n31817 = ~n31814 & ~n31816 ;
  assign n31818 = ~n31808 & n31817 ;
  assign n31819 = ~n31804 & n31818 ;
  assign n31820 = ~n31803 & ~n31819 ;
  assign n31821 = ~n22766 & ~n31810 ;
  assign n31822 = ~n22766 & n22767 ;
  assign n31823 = ~n31699 & n31822 ;
  assign n31824 = ~n31821 & ~n31823 ;
  assign n31825 = n22788 & ~n31699 ;
  assign n31826 = n31796 & ~n31825 ;
  assign n31827 = ~n31824 & ~n31826 ;
  assign n31828 = ~n22787 & n31827 ;
  assign n31829 = \pi0785  & ~n31828 ;
  assign n31830 = n31820 & n31829 ;
  assign n31831 = ~\pi0785  & ~n31792 ;
  assign n31832 = ~n31767 & n31831 ;
  assign n31833 = n23673 & ~n31784 ;
  assign n31834 = ~n31832 & ~n31833 ;
  assign n31835 = n26700 & n31834 ;
  assign n31836 = ~n31830 & n31835 ;
  assign n31837 = n22155 & ~n31702 ;
  assign n31838 = ~n22147 & ~n31633 ;
  assign n31839 = n31630 & n31838 ;
  assign n31840 = ~n22148 & ~n31839 ;
  assign n31841 = n22147 & ~n31616 ;
  assign n31842 = n30053 & ~n31841 ;
  assign n31843 = n31840 & n31842 ;
  assign n31844 = \pi0778  & n31842 ;
  assign n31845 = ~n31652 & n31844 ;
  assign n31846 = ~n31843 & ~n31845 ;
  assign n31847 = ~n31837 & n31846 ;
  assign n31848 = ~n21034 & ~n31847 ;
  assign n31849 = ~n23880 & ~n31710 ;
  assign n31850 = n23880 & ~n31616 ;
  assign n31851 = n24691 & ~n31850 ;
  assign n31852 = ~n31849 & n31851 ;
  assign n31853 = \pi0628  & ~n31656 ;
  assign n31854 = ~n31655 & n31853 ;
  assign n31855 = ~n31653 & n31854 ;
  assign n31856 = ~\pi0176  & ~\pi0628  ;
  assign n31857 = n21768 & n31856 ;
  assign n31858 = n21770 & n31856 ;
  assign n31859 = ~n21734 & n31858 ;
  assign n31860 = ~n31857 & ~n31859 ;
  assign n31861 = n20843 & n31860 ;
  assign n31862 = ~n31855 & n31861 ;
  assign n31863 = ~\pi0628  & ~n31656 ;
  assign n31864 = ~n31655 & n31863 ;
  assign n31865 = ~n31653 & n31864 ;
  assign n31866 = ~\pi0176  & \pi0628  ;
  assign n31867 = n21768 & n31866 ;
  assign n31868 = n21770 & n31866 ;
  assign n31869 = ~n21734 & n31868 ;
  assign n31870 = ~n31867 & ~n31869 ;
  assign n31871 = n20844 & n31870 ;
  assign n31872 = ~n31865 & n31871 ;
  assign n31873 = ~n31862 & ~n31872 ;
  assign n31874 = ~n31852 & n31873 ;
  assign n31875 = \pi0792  & ~n31874 ;
  assign n31876 = n30780 & ~n31652 ;
  assign n31877 = n31274 & ~n31654 ;
  assign n31878 = ~n23380 & n31616 ;
  assign n31879 = ~n31877 & ~n31878 ;
  assign n31880 = ~n31876 & n31879 ;
  assign n31881 = ~n31283 & ~n31880 ;
  assign n31882 = n23683 & n31702 ;
  assign n31883 = n21032 & n31705 ;
  assign n31884 = ~n31704 & n31883 ;
  assign n31885 = ~n21032 & ~n31616 ;
  assign n31886 = ~n20876 & ~n31885 ;
  assign n31887 = \pi0789  & n31886 ;
  assign n31888 = ~n31884 & n31887 ;
  assign n31889 = ~n31882 & n31888 ;
  assign n31890 = ~n21038 & ~n31889 ;
  assign n31891 = ~n31881 & n31890 ;
  assign n31892 = ~n31875 & n31891 ;
  assign n31893 = ~n31848 & n31892 ;
  assign n31894 = ~n31836 & n31893 ;
  assign n31895 = \pi0626  & n31616 ;
  assign n31896 = n20882 & ~n31895 ;
  assign n31897 = ~\pi0626  & ~n31708 ;
  assign n31898 = ~n31707 & n31897 ;
  assign n31899 = ~n31703 & n31898 ;
  assign n31900 = n31896 & ~n31899 ;
  assign n31901 = \pi0626  & ~n31708 ;
  assign n31902 = ~n31707 & n31901 ;
  assign n31903 = ~n31703 & n31902 ;
  assign n31904 = ~\pi0626  & n31616 ;
  assign n31905 = n20881 & ~n31904 ;
  assign n31906 = ~n31903 & n31905 ;
  assign n31907 = ~n31900 & ~n31906 ;
  assign n31908 = n20951 & ~n31616 ;
  assign n31909 = ~n31301 & ~n31908 ;
  assign n31910 = ~n31877 & ~n31909 ;
  assign n31911 = ~n31876 & n31910 ;
  assign n31912 = n31306 & ~n31616 ;
  assign n31913 = ~n23856 & ~n31912 ;
  assign n31914 = ~n31911 & n31913 ;
  assign n31915 = n31907 & n31914 ;
  assign n31916 = ~n26803 & ~n31915 ;
  assign n31917 = ~n31875 & n31916 ;
  assign n31918 = ~n21067 & ~n31917 ;
  assign n31919 = ~n31894 & n31918 ;
  assign n31920 = n30376 & ~n31710 ;
  assign n31921 = ~n20846 & n23880 ;
  assign n31922 = ~n31616 & n31921 ;
  assign n31923 = n20846 & ~n31616 ;
  assign n31924 = ~n20910 & ~n31923 ;
  assign n31925 = ~n31922 & n31924 ;
  assign n31926 = ~n31920 & n31925 ;
  assign n31927 = n21768 & n31475 ;
  assign n31928 = n21770 & n31475 ;
  assign n31929 = ~n21734 & n31928 ;
  assign n31930 = ~n31927 & ~n31929 ;
  assign n31931 = n20850 & n31930 ;
  assign n31932 = n20849 & n31930 ;
  assign n31933 = ~n31660 & n31932 ;
  assign n31934 = ~n31659 & n31933 ;
  assign n31935 = ~n31931 & ~n31934 ;
  assign n31936 = n21768 & n31471 ;
  assign n31937 = n21770 & n31471 ;
  assign n31938 = ~n21734 & n31937 ;
  assign n31939 = ~n31936 & ~n31938 ;
  assign n31940 = n31338 & n31939 ;
  assign n31941 = n20897 & n31939 ;
  assign n31942 = ~n31660 & n31941 ;
  assign n31943 = ~n31659 & n31942 ;
  assign n31944 = ~n31940 & ~n31943 ;
  assign n31945 = n31935 & n31944 ;
  assign n31946 = ~n31926 & n31945 ;
  assign n31947 = \pi0787  & ~n31946 ;
  assign n31948 = n31378 & ~n31713 ;
  assign n31949 = n26824 & ~n31719 ;
  assign n31950 = \pi0790  & ~n31949 ;
  assign n31951 = ~n31948 & n31950 ;
  assign n31952 = ~n31947 & ~n31951 ;
  assign n31953 = ~n31609 & n31952 ;
  assign n31954 = ~n31919 & n31953 ;
  assign n31955 = ~n31735 & ~n31954 ;
  assign n31956 = n9948 & ~n31955 ;
  assign n31957 = ~n31612 & ~n31956 ;
  assign n31958 = \pi0177  & ~\pi0832  ;
  assign n31959 = ~n21132 & ~n31958 ;
  assign n31960 = ~\pi0177  & n21768 ;
  assign n31961 = ~\pi0177  & n21770 ;
  assign n31962 = ~n21734 & n31961 ;
  assign n31963 = ~n31960 & ~n31962 ;
  assign n31964 = ~n21777 & n31963 ;
  assign n31965 = ~\pi0781  & ~n31964 ;
  assign n31966 = ~\pi0789  & ~n31965 ;
  assign n31967 = ~\pi0177  & ~n25033 ;
  assign n31968 = ~n25040 & n31967 ;
  assign n31969 = ~n25028 & n31968 ;
  assign n31970 = \pi0177  & ~n25040 ;
  assign n31971 = ~n25024 & n31970 ;
  assign n31972 = ~n31969 & ~n31971 ;
  assign n31973 = ~\pi0757  & n6861 ;
  assign n31974 = ~n31972 & n31973 ;
  assign n31975 = \pi0177  & ~n6861 ;
  assign n31976 = ~\pi0177  & n22124 ;
  assign n31977 = ~n31962 & ~n31976 ;
  assign n31978 = \pi0757  & n1289 ;
  assign n31979 = n1287 & n31978 ;
  assign n31980 = n31977 & n31979 ;
  assign n31981 = ~n31975 & ~n31980 ;
  assign n31982 = ~n31974 & n31981 ;
  assign n31983 = ~\pi0789  & n21777 ;
  assign n31984 = ~n31982 & n31983 ;
  assign n31985 = ~n31966 & ~n31984 ;
  assign n31986 = ~n23880 & n31985 ;
  assign n31987 = ~\pi0177  & ~n20811 ;
  assign n31988 = n21768 & n31987 ;
  assign n31989 = n21770 & n31987 ;
  assign n31990 = ~n21734 & n31989 ;
  assign n31991 = ~n31988 & ~n31990 ;
  assign n31992 = n20811 & ~n31964 ;
  assign n31993 = n31991 & ~n31992 ;
  assign n31994 = n21777 & n31991 ;
  assign n31995 = ~n31982 & n31994 ;
  assign n31996 = ~n31993 & ~n31995 ;
  assign n31997 = \pi0781  & ~n23880 ;
  assign n31998 = n31996 & n31997 ;
  assign n31999 = ~n31986 & ~n31998 ;
  assign n32000 = n23880 & ~n31963 ;
  assign n32001 = n24691 & ~n32000 ;
  assign n32002 = n31999 & n32001 ;
  assign n32003 = n22869 & n31996 ;
  assign n32004 = n21777 & ~n31982 ;
  assign n32005 = ~\pi0619  & n31965 ;
  assign n32006 = ~n32004 & n32005 ;
  assign n32007 = ~\pi0177  & \pi0619  ;
  assign n32008 = n21768 & n32007 ;
  assign n32009 = n21770 & n32007 ;
  assign n32010 = ~n21734 & n32009 ;
  assign n32011 = ~n32008 & ~n32010 ;
  assign n32012 = ~\pi1159  & n32011 ;
  assign n32013 = ~n32006 & n32012 ;
  assign n32014 = ~n32003 & n32013 ;
  assign n32015 = n22859 & n31996 ;
  assign n32016 = \pi0619  & n31965 ;
  assign n32017 = ~n32004 & n32016 ;
  assign n32018 = ~\pi0177  & ~\pi0619  ;
  assign n32019 = n21768 & n32018 ;
  assign n32020 = n21770 & n32018 ;
  assign n32021 = ~n21734 & n32020 ;
  assign n32022 = ~n32019 & ~n32021 ;
  assign n32023 = \pi1159  & n32022 ;
  assign n32024 = ~n32017 & n32023 ;
  assign n32025 = ~n32015 & n32024 ;
  assign n32026 = ~n32014 & ~n32025 ;
  assign n32027 = \pi0789  & n32001 ;
  assign n32028 = ~n32026 & n32027 ;
  assign n32029 = ~n32002 & ~n32028 ;
  assign n32030 = ~n23380 & n31963 ;
  assign n32031 = ~\pi0778  & n31975 ;
  assign n32032 = ~\pi0177  & ~n22017 ;
  assign n32033 = ~n21994 & n32032 ;
  assign n32034 = ~\pi0038  & ~\pi0177  ;
  assign n32035 = ~n22109 & ~n32034 ;
  assign n32036 = ~n32033 & ~n32035 ;
  assign n32037 = ~\pi0177  & ~n21757 ;
  assign n32038 = n22117 & ~n32037 ;
  assign n32039 = ~\pi0686  & ~n32038 ;
  assign n32040 = ~n32036 & n32039 ;
  assign n32041 = \pi0686  & ~n31977 ;
  assign n32042 = ~n32040 & ~n32041 ;
  assign n32043 = n25171 & n32042 ;
  assign n32044 = ~n32031 & ~n32043 ;
  assign n32045 = ~n22147 & ~n32044 ;
  assign n32046 = ~n22155 & n32045 ;
  assign n32047 = ~\pi0177  & \pi0625  ;
  assign n32048 = ~n22727 & ~n32047 ;
  assign n32049 = ~\pi0177  & ~\pi0625  ;
  assign n32050 = n21768 & n32049 ;
  assign n32051 = n21770 & n32049 ;
  assign n32052 = ~n21734 & n32051 ;
  assign n32053 = ~n32050 & ~n32052 ;
  assign n32054 = \pi1153  & n32053 ;
  assign n32055 = n32048 & n32054 ;
  assign n32056 = n6861 & n32054 ;
  assign n32057 = n32042 & n32056 ;
  assign n32058 = ~n32055 & ~n32057 ;
  assign n32059 = ~n22734 & ~n32049 ;
  assign n32060 = n21768 & n32047 ;
  assign n32061 = n21770 & n32047 ;
  assign n32062 = ~n21734 & n32061 ;
  assign n32063 = ~n32060 & ~n32062 ;
  assign n32064 = ~\pi1153  & n32063 ;
  assign n32065 = n32059 & n32064 ;
  assign n32066 = n6861 & n32064 ;
  assign n32067 = n32042 & n32066 ;
  assign n32068 = ~n32065 & ~n32067 ;
  assign n32069 = n32058 & n32068 ;
  assign n32070 = n23697 & ~n32069 ;
  assign n32071 = ~n32046 & ~n32070 ;
  assign n32072 = ~n32030 & n32071 ;
  assign n32073 = n22162 & ~n32072 ;
  assign n32074 = ~n22162 & n31963 ;
  assign n32075 = ~\pi0628  & ~n32074 ;
  assign n32076 = ~n32073 & n32075 ;
  assign n32077 = ~\pi0177  & \pi0628  ;
  assign n32078 = n21768 & n32077 ;
  assign n32079 = n21770 & n32077 ;
  assign n32080 = ~n21734 & n32079 ;
  assign n32081 = ~n32078 & ~n32080 ;
  assign n32082 = n20844 & n32081 ;
  assign n32083 = ~n32076 & n32082 ;
  assign n32084 = \pi0628  & ~n32074 ;
  assign n32085 = ~n32073 & n32084 ;
  assign n32086 = ~\pi0177  & ~\pi0628  ;
  assign n32087 = n21768 & n32086 ;
  assign n32088 = n21770 & n32086 ;
  assign n32089 = ~n21734 & n32088 ;
  assign n32090 = ~n32087 & ~n32089 ;
  assign n32091 = n20843 & n32090 ;
  assign n32092 = ~n32085 & n32091 ;
  assign n32093 = ~n32083 & ~n32092 ;
  assign n32094 = n32029 & n32093 ;
  assign n32095 = \pi0792  & ~n32094 ;
  assign n32096 = ~n21067 & n32095 ;
  assign n32097 = \pi0619  & ~n32030 ;
  assign n32098 = n32071 & n32097 ;
  assign n32099 = ~\pi1159  & ~n32098 ;
  assign n32100 = ~\pi0648  & ~n32025 ;
  assign n32101 = ~n32099 & n32100 ;
  assign n32102 = ~\pi0619  & ~n32030 ;
  assign n32103 = n32071 & n32102 ;
  assign n32104 = \pi1159  & ~n32103 ;
  assign n32105 = \pi0648  & ~n32014 ;
  assign n32106 = ~n32104 & n32105 ;
  assign n32107 = ~n32101 & ~n32106 ;
  assign n32108 = n29818 & ~n32107 ;
  assign n32109 = n22148 & ~n32069 ;
  assign n32110 = ~n32045 & ~n32109 ;
  assign n32111 = n20871 & ~n31996 ;
  assign n32112 = n22147 & n31963 ;
  assign n32113 = ~n32111 & ~n32112 ;
  assign n32114 = n32110 & n32113 ;
  assign n32115 = n22155 & ~n31996 ;
  assign n32116 = ~n24348 & ~n32115 ;
  assign n32117 = ~n32114 & ~n32116 ;
  assign n32118 = n20828 & n32022 ;
  assign n32119 = ~n32017 & n32118 ;
  assign n32120 = ~n32015 & n32119 ;
  assign n32121 = \pi0619  & \pi0648  ;
  assign n32122 = ~n32011 & n32121 ;
  assign n32123 = ~\pi0619  & ~\pi0648  ;
  assign n32124 = \pi1159  & n32121 ;
  assign n32125 = ~n32123 & ~n32124 ;
  assign n32126 = ~n32122 & n32125 ;
  assign n32127 = ~n32120 & ~n32126 ;
  assign n32128 = \pi0789  & ~n32127 ;
  assign n32129 = ~n32117 & ~n32128 ;
  assign n32130 = ~n21038 & n32129 ;
  assign n32131 = ~n32108 & ~n32130 ;
  assign n32132 = \pi0177  & ~n23558 ;
  assign n32133 = n23557 & n32132 ;
  assign n32134 = ~\pi0039  & ~\pi0177  ;
  assign n32135 = ~n22683 & n32134 ;
  assign n32136 = ~\pi0177  & ~n23548 ;
  assign n32137 = ~\pi0038  & ~n32136 ;
  assign n32138 = ~n32135 & n32137 ;
  assign n32139 = ~n32133 & n32138 ;
  assign n32140 = n25195 & ~n32037 ;
  assign n32141 = ~\pi0757  & ~n32140 ;
  assign n32142 = ~n32139 & n32141 ;
  assign n32143 = n23587 & ~n32037 ;
  assign n32144 = ~\pi0177  & \pi0757  ;
  assign n32145 = ~n32143 & n32144 ;
  assign n32146 = ~n23568 & n32145 ;
  assign n32147 = \pi0757  & ~n32143 ;
  assign n32148 = \pi0038  & n32147 ;
  assign n32149 = \pi0177  & n23575 ;
  assign n32150 = n32147 & n32149 ;
  assign n32151 = n23572 & n32150 ;
  assign n32152 = ~n32148 & ~n32151 ;
  assign n32153 = ~n32146 & n32152 ;
  assign n32154 = ~n32142 & n32153 ;
  assign n32155 = ~\pi0686  & ~n32154 ;
  assign n32156 = \pi0757  & n31977 ;
  assign n32157 = \pi0686  & \pi0757  ;
  assign n32158 = \pi0686  & ~n31971 ;
  assign n32159 = ~n31969 & n32158 ;
  assign n32160 = ~n32157 & ~n32159 ;
  assign n32161 = ~n32156 & ~n32160 ;
  assign n32162 = n6861 & ~n32161 ;
  assign n32163 = ~n32155 & n32162 ;
  assign n32164 = ~n32059 & ~n32163 ;
  assign n32165 = ~n31980 & ~n32048 ;
  assign n32166 = ~n31974 & n32165 ;
  assign n32167 = ~\pi1153  & ~n32166 ;
  assign n32168 = ~n32164 & n32167 ;
  assign n32169 = ~\pi0608  & n32058 ;
  assign n32170 = ~n32168 & n32169 ;
  assign n32171 = ~n32048 & ~n32163 ;
  assign n32172 = ~n31980 & ~n32059 ;
  assign n32173 = ~n31974 & n32172 ;
  assign n32174 = \pi1153  & ~n32173 ;
  assign n32175 = ~n32171 & n32174 ;
  assign n32176 = \pi0608  & n32068 ;
  assign n32177 = ~n32175 & n32176 ;
  assign n32178 = ~n32170 & ~n32177 ;
  assign n32179 = n23638 & ~n32178 ;
  assign n32180 = \pi0778  & ~n32069 ;
  assign n32181 = ~\pi0609  & n32044 ;
  assign n32182 = ~n32180 & n32181 ;
  assign n32183 = ~\pi0177  & ~\pi0778  ;
  assign n32184 = ~n23622 & ~n32183 ;
  assign n32185 = \pi0609  & ~n32184 ;
  assign n32186 = ~n32163 & n32185 ;
  assign n32187 = ~n22788 & n31963 ;
  assign n32188 = ~\pi0660  & ~n32187 ;
  assign n32189 = \pi1155  & ~n32188 ;
  assign n32190 = n31798 & ~n31982 ;
  assign n32191 = ~n32189 & ~n32190 ;
  assign n32192 = ~n32186 & ~n32191 ;
  assign n32193 = ~n32182 & n32192 ;
  assign n32194 = ~n32179 & n32193 ;
  assign n32195 = n23613 & ~n32178 ;
  assign n32196 = \pi0609  & n32044 ;
  assign n32197 = ~n32180 & n32196 ;
  assign n32198 = ~n22767 & n31963 ;
  assign n32199 = \pi0660  & ~n32198 ;
  assign n32200 = ~\pi1155  & ~n32199 ;
  assign n32201 = n31812 & ~n31982 ;
  assign n32202 = ~n32200 & ~n32201 ;
  assign n32203 = ~\pi0609  & ~n32184 ;
  assign n32204 = ~n32163 & n32203 ;
  assign n32205 = ~n32202 & ~n32204 ;
  assign n32206 = ~n32197 & n32205 ;
  assign n32207 = ~n32195 & n32206 ;
  assign n32208 = ~n32194 & ~n32207 ;
  assign n32209 = ~n22766 & ~n32199 ;
  assign n32210 = n31822 & ~n31982 ;
  assign n32211 = ~n32209 & ~n32210 ;
  assign n32212 = n22788 & ~n31982 ;
  assign n32213 = n32188 & ~n32212 ;
  assign n32214 = ~n32211 & ~n32213 ;
  assign n32215 = ~n22787 & n32214 ;
  assign n32216 = \pi0785  & ~n32215 ;
  assign n32217 = n32208 & n32216 ;
  assign n32218 = n23673 & ~n32178 ;
  assign n32219 = ~\pi0785  & ~n32184 ;
  assign n32220 = ~n32163 & n32219 ;
  assign n32221 = n21022 & ~n32220 ;
  assign n32222 = ~n32218 & n32221 ;
  assign n32223 = ~n32108 & n32222 ;
  assign n32224 = ~n32217 & n32223 ;
  assign n32225 = ~n32131 & ~n32224 ;
  assign n32226 = \pi0789  & ~n32026 ;
  assign n32227 = \pi0781  & n31996 ;
  assign n32228 = ~n31985 & ~n32227 ;
  assign n32229 = n30606 & ~n32228 ;
  assign n32230 = ~n32226 & n32229 ;
  assign n32231 = ~\pi0641  & n31963 ;
  assign n32232 = n20776 & ~n32231 ;
  assign n32233 = ~n22160 & ~n32030 ;
  assign n32234 = n32071 & n32233 ;
  assign n32235 = ~\pi0177  & \pi0789  ;
  assign n32236 = ~n20876 & n32235 ;
  assign n32237 = n21768 & n32236 ;
  assign n32238 = n21770 & n32236 ;
  assign n32239 = ~n21734 & n32238 ;
  assign n32240 = ~n32237 & ~n32239 ;
  assign n32241 = \pi0641  & n32240 ;
  assign n32242 = ~n32234 & n32241 ;
  assign n32243 = n32232 & ~n32242 ;
  assign n32244 = ~n32230 & ~n32243 ;
  assign n32245 = \pi0641  & n31963 ;
  assign n32246 = n20777 & ~n32245 ;
  assign n32247 = ~n23856 & ~n32246 ;
  assign n32248 = ~\pi0641  & n32240 ;
  assign n32249 = ~n23856 & n32248 ;
  assign n32250 = ~n32234 & n32249 ;
  assign n32251 = ~n32247 & ~n32250 ;
  assign n32252 = n32244 & ~n32251 ;
  assign n32253 = ~n26803 & ~n32252 ;
  assign n32254 = ~n21067 & ~n32253 ;
  assign n32255 = ~n32225 & n32254 ;
  assign n32256 = ~n32096 & ~n32255 ;
  assign n32257 = ~n24761 & ~n32256 ;
  assign n32258 = ~\pi0792  & n32074 ;
  assign n32259 = ~\pi0792  & n22162 ;
  assign n32260 = ~n32072 & n32259 ;
  assign n32261 = ~n32258 & ~n32260 ;
  assign n32262 = \pi0647  & n32261 ;
  assign n32263 = ~\pi0177  & ~\pi0647  ;
  assign n32264 = n21768 & n32263 ;
  assign n32265 = n21770 & n32263 ;
  assign n32266 = ~n21734 & n32265 ;
  assign n32267 = ~n32264 & ~n32266 ;
  assign n32268 = n20849 & n32267 ;
  assign n32269 = ~n32262 & n32268 ;
  assign n32270 = \pi1156  & n32090 ;
  assign n32271 = ~n32085 & n32270 ;
  assign n32272 = ~\pi1156  & n32081 ;
  assign n32273 = ~n32076 & n32272 ;
  assign n32274 = ~n32271 & ~n32273 ;
  assign n32275 = \pi0792  & n32268 ;
  assign n32276 = ~n32274 & n32275 ;
  assign n32277 = ~n32269 & ~n32276 ;
  assign n32278 = ~\pi0647  & n32261 ;
  assign n32279 = ~\pi0177  & \pi0647  ;
  assign n32280 = n21768 & n32279 ;
  assign n32281 = n21770 & n32279 ;
  assign n32282 = ~n21734 & n32281 ;
  assign n32283 = ~n32280 & ~n32282 ;
  assign n32284 = n20897 & n32283 ;
  assign n32285 = ~n32278 & n32284 ;
  assign n32286 = \pi0792  & n32284 ;
  assign n32287 = ~n32274 & n32286 ;
  assign n32288 = ~n32285 & ~n32287 ;
  assign n32289 = n30376 & n32228 ;
  assign n32290 = \pi0789  & n30376 ;
  assign n32291 = ~n32026 & n32290 ;
  assign n32292 = ~n32289 & ~n32291 ;
  assign n32293 = ~n30376 & n31963 ;
  assign n32294 = n32292 & ~n32293 ;
  assign n32295 = ~n20910 & ~n32294 ;
  assign n32296 = n32288 & ~n32295 ;
  assign n32297 = n32277 & n32296 ;
  assign n32298 = \pi0787  & ~n24761 ;
  assign n32299 = ~n32297 & n32298 ;
  assign n32300 = n9948 & ~n32299 ;
  assign n32301 = ~n32257 & n32300 ;
  assign n32302 = ~n31959 & ~n32301 ;
  assign n32303 = ~\pi1157  & n32283 ;
  assign n32304 = ~n32278 & n32303 ;
  assign n32305 = \pi0792  & n32303 ;
  assign n32306 = ~n32274 & n32305 ;
  assign n32307 = ~n32304 & ~n32306 ;
  assign n32308 = \pi1157  & n32267 ;
  assign n32309 = ~n32262 & n32308 ;
  assign n32310 = \pi0792  & n32308 ;
  assign n32311 = ~n32274 & n32310 ;
  assign n32312 = ~n32309 & ~n32311 ;
  assign n32313 = n32307 & n32312 ;
  assign n32314 = \pi0787  & n23313 ;
  assign n32315 = ~n32313 & n32314 ;
  assign n32316 = ~\pi0787  & ~n32261 ;
  assign n32317 = n23011 & ~n32274 ;
  assign n32318 = ~n32316 & ~n32317 ;
  assign n32319 = n23313 & ~n32318 ;
  assign n32320 = ~\pi0177  & ~\pi0644  ;
  assign n32321 = n21768 & n32320 ;
  assign n32322 = n21770 & n32320 ;
  assign n32323 = ~n21734 & n32322 ;
  assign n32324 = ~n32321 & ~n32323 ;
  assign n32325 = ~\pi0715  & n32324 ;
  assign n32326 = \pi1160  & ~n32325 ;
  assign n32327 = n21092 & n31999 ;
  assign n32328 = \pi0789  & n21092 ;
  assign n32329 = ~n32026 & n32328 ;
  assign n32330 = ~n32327 & ~n32329 ;
  assign n32331 = ~n32000 & ~n32330 ;
  assign n32332 = ~n21092 & n31963 ;
  assign n32333 = n26824 & ~n32332 ;
  assign n32334 = ~n32331 & n32333 ;
  assign n32335 = ~n32326 & ~n32334 ;
  assign n32336 = ~n32319 & ~n32335 ;
  assign n32337 = ~n32315 & n32336 ;
  assign n32338 = \pi0790  & ~n32337 ;
  assign n32339 = \pi0787  & n23312 ;
  assign n32340 = ~n32313 & n32339 ;
  assign n32341 = n23312 & ~n32318 ;
  assign n32342 = ~\pi0177  & \pi0644  ;
  assign n32343 = n21768 & n32342 ;
  assign n32344 = n21770 & n32342 ;
  assign n32345 = ~n21734 & n32344 ;
  assign n32346 = ~n32343 & ~n32345 ;
  assign n32347 = \pi0715  & n32346 ;
  assign n32348 = ~\pi1160  & ~n32347 ;
  assign n32349 = n31378 & ~n32332 ;
  assign n32350 = ~n32331 & n32349 ;
  assign n32351 = ~n32348 & ~n32350 ;
  assign n32352 = ~n32341 & ~n32351 ;
  assign n32353 = ~n32340 & n32352 ;
  assign n32354 = ~n31959 & ~n32353 ;
  assign n32355 = n32338 & n32354 ;
  assign n32356 = ~\pi0686  & n1689 ;
  assign n32357 = n20855 & n32356 ;
  assign n32358 = ~n20861 & n32357 ;
  assign n32359 = ~\pi0177  & ~n1689 ;
  assign n32360 = ~n32358 & ~n32359 ;
  assign n32361 = n20879 & ~n32360 ;
  assign n32362 = n20938 & n32361 ;
  assign n32363 = n29714 & ~n32362 ;
  assign n32364 = ~n21032 & ~n32359 ;
  assign n32365 = \pi0789  & n32364 ;
  assign n32366 = n23423 & ~n32365 ;
  assign n32367 = ~\pi0757  & n1689 ;
  assign n32368 = n20784 & n32367 ;
  assign n32369 = ~n32359 & ~n32368 ;
  assign n32370 = n20794 & ~n32369 ;
  assign n32371 = n20796 & ~n32370 ;
  assign n32372 = n20799 & ~n32369 ;
  assign n32373 = n20801 & ~n32372 ;
  assign n32374 = ~n32371 & ~n32373 ;
  assign n32375 = ~\pi0785  & ~n32359 ;
  assign n32376 = ~n32368 & n32375 ;
  assign n32377 = ~n20804 & ~n32376 ;
  assign n32378 = ~n20812 & n32377 ;
  assign n32379 = ~n32365 & n32378 ;
  assign n32380 = n32374 & n32379 ;
  assign n32381 = ~n32366 & ~n32380 ;
  assign n32382 = ~n23880 & ~n32381 ;
  assign n32383 = n21077 & n32361 ;
  assign n32384 = n29709 & ~n32383 ;
  assign n32385 = \pi0792  & ~n32384 ;
  assign n32386 = n32382 & n32385 ;
  assign n32387 = ~\pi0177  & \pi0788  ;
  assign n32388 = ~n1689 & n32387 ;
  assign n32389 = ~n20778 & n32388 ;
  assign n32390 = \pi0629  & ~n32389 ;
  assign n32391 = ~n32362 & n32390 ;
  assign n32392 = ~\pi0629  & ~n32389 ;
  assign n32393 = ~n32383 & n32392 ;
  assign n32394 = ~n32391 & ~n32393 ;
  assign n32395 = n32385 & n32394 ;
  assign n32396 = ~n32386 & ~n32395 ;
  assign n32397 = ~n32363 & ~n32396 ;
  assign n32398 = ~n21067 & ~n32397 ;
  assign n32399 = ~\pi0177  & \pi0792  ;
  assign n32400 = ~n1689 & n32399 ;
  assign n32401 = ~n20845 & n32400 ;
  assign n32402 = ~n20910 & ~n32401 ;
  assign n32403 = n20846 & n32402 ;
  assign n32404 = n20895 & n32361 ;
  assign n32405 = ~n1689 & n32279 ;
  assign n32406 = n20897 & ~n32405 ;
  assign n32407 = ~n32404 & n32406 ;
  assign n32408 = ~n1689 & n32263 ;
  assign n32409 = n20849 & ~n32408 ;
  assign n32410 = ~n24761 & ~n32409 ;
  assign n32411 = n31479 & n32361 ;
  assign n32412 = ~n32410 & ~n32411 ;
  assign n32413 = ~n32407 & ~n32412 ;
  assign n32414 = ~n32403 & n32413 ;
  assign n32415 = ~n29722 & ~n32414 ;
  assign n32416 = ~n32389 & n32402 ;
  assign n32417 = ~n29722 & n32416 ;
  assign n32418 = ~n32382 & n32417 ;
  assign n32419 = ~n32415 & ~n32418 ;
  assign n32420 = ~n32398 & n32419 ;
  assign n32421 = ~\pi0626  & n32381 ;
  assign n32422 = \pi0626  & ~n32359 ;
  assign n32423 = n20882 & ~n32422 ;
  assign n32424 = ~n32421 & n32423 ;
  assign n32425 = n23170 & ~n32360 ;
  assign n32426 = ~\pi0626  & ~n32359 ;
  assign n32427 = n20881 & ~n32426 ;
  assign n32428 = ~n32425 & ~n32427 ;
  assign n32429 = \pi0626  & ~n32425 ;
  assign n32430 = n32381 & n32429 ;
  assign n32431 = ~n32428 & ~n32430 ;
  assign n32432 = ~n32424 & ~n32431 ;
  assign n32433 = \pi0788  & ~n32432 ;
  assign n32434 = ~\pi0686  & ~n20784 ;
  assign n32435 = ~\pi0686  & ~n20790 ;
  assign n32436 = n20789 & n32435 ;
  assign n32437 = ~n32434 & ~n32436 ;
  assign n32438 = n24915 & ~n32437 ;
  assign n32439 = \pi0603  & ~\pi0757  ;
  assign n32440 = ~n20783 & n32439 ;
  assign n32441 = ~n20985 & n32440 ;
  assign n32442 = ~n32359 & ~n32441 ;
  assign n32443 = ~n32438 & n32442 ;
  assign n32444 = \pi0177  & ~n1689 ;
  assign n32445 = ~\pi0609  & ~n32444 ;
  assign n32446 = ~n32443 & n32445 ;
  assign n32447 = ~\pi1155  & ~n32359 ;
  assign n32448 = ~n32358 & n32447 ;
  assign n32449 = ~n20999 & ~n32448 ;
  assign n32450 = ~n32446 & ~n32449 ;
  assign n32451 = \pi1155  & ~n32372 ;
  assign n32452 = ~\pi0660  & ~n32451 ;
  assign n32453 = ~n32450 & n32452 ;
  assign n32454 = ~n21007 & ~n32371 ;
  assign n32455 = \pi0609  & ~n32444 ;
  assign n32456 = ~n32443 & n32455 ;
  assign n32457 = \pi1155  & ~n32359 ;
  assign n32458 = ~n32358 & n32457 ;
  assign n32459 = ~n21774 & ~n32458 ;
  assign n32460 = \pi0785  & ~n32459 ;
  assign n32461 = ~n32456 & n32460 ;
  assign n32462 = n32454 & ~n32461 ;
  assign n32463 = ~n32453 & ~n32462 ;
  assign n32464 = n21022 & ~n32444 ;
  assign n32465 = ~n32443 & n32464 ;
  assign n32466 = ~n21023 & ~n32465 ;
  assign n32467 = ~n32463 & ~n32466 ;
  assign n32468 = n20964 & n32377 ;
  assign n32469 = n32374 & n32468 ;
  assign n32470 = \pi0627  & ~n32359 ;
  assign n32471 = ~n32358 & n32470 ;
  assign n32472 = ~n20968 & ~n32471 ;
  assign n32473 = ~n32469 & ~n32472 ;
  assign n32474 = ~\pi0627  & ~n32359 ;
  assign n32475 = ~n32358 & n32474 ;
  assign n32476 = ~n20978 & ~n32475 ;
  assign n32477 = \pi0781  & n32476 ;
  assign n32478 = n20974 & n32377 ;
  assign n32479 = \pi0781  & n32478 ;
  assign n32480 = n32374 & n32479 ;
  assign n32481 = ~n32477 & ~n32480 ;
  assign n32482 = ~n32473 & ~n32481 ;
  assign n32483 = ~n21034 & ~n32482 ;
  assign n32484 = ~n32467 & n32483 ;
  assign n32485 = n21050 & ~n32359 ;
  assign n32486 = ~n32358 & n32485 ;
  assign n32487 = ~n21051 & ~n32486 ;
  assign n32488 = ~n20876 & n32364 ;
  assign n32489 = ~n21038 & ~n32488 ;
  assign n32490 = n32487 & n32489 ;
  assign n32491 = ~n23177 & ~n32490 ;
  assign n32492 = n32374 & n32378 ;
  assign n32493 = n31562 & ~n32492 ;
  assign n32494 = ~n32491 & ~n32493 ;
  assign n32495 = ~n32484 & n32494 ;
  assign n32496 = ~n32433 & ~n32495 ;
  assign n32497 = ~n23856 & n32419 ;
  assign n32498 = ~n32496 & n32497 ;
  assign n32499 = ~n32420 & ~n32498 ;
  assign n32500 = n24830 & n32361 ;
  assign n32501 = \pi1157  & ~n32408 ;
  assign n32502 = ~n32500 & n32501 ;
  assign n32503 = ~\pi1157  & ~n32405 ;
  assign n32504 = ~n32404 & n32503 ;
  assign n32505 = ~n32502 & ~n32504 ;
  assign n32506 = \pi0787  & ~n32505 ;
  assign n32507 = n24844 & n32361 ;
  assign n32508 = ~n24843 & ~n32507 ;
  assign n32509 = ~n32506 & ~n32508 ;
  assign n32510 = n31580 & n32389 ;
  assign n32511 = n31582 & ~n32381 ;
  assign n32512 = ~n32510 & ~n32511 ;
  assign n32513 = ~n32509 & n32512 ;
  assign n32514 = n23313 & ~n32513 ;
  assign n32515 = \pi0790  & n32514 ;
  assign n32516 = n31588 & n32389 ;
  assign n32517 = n31590 & ~n32381 ;
  assign n32518 = ~n32516 & ~n32517 ;
  assign n32519 = ~n23414 & n32359 ;
  assign n32520 = ~n24886 & n32519 ;
  assign n32521 = n20891 & n32361 ;
  assign n32522 = ~\pi0787  & ~n32521 ;
  assign n32523 = ~\pi1160  & ~n32522 ;
  assign n32524 = ~n32506 & n32523 ;
  assign n32525 = ~n32520 & ~n32524 ;
  assign n32526 = n32518 & n32525 ;
  assign n32527 = ~n23312 & ~n32519 ;
  assign n32528 = ~n31603 & ~n32527 ;
  assign n32529 = \pi0790  & n32528 ;
  assign n32530 = ~n32526 & n32529 ;
  assign n32531 = ~n32515 & ~n32530 ;
  assign n32532 = \pi0832  & n32531 ;
  assign n32533 = n32499 & n32532 ;
  assign n32534 = ~n32355 & ~n32533 ;
  assign n32535 = ~n32302 & n32534 ;
  assign n32536 = ~\pi0178  & \pi0788  ;
  assign n32537 = ~n1689 & n32536 ;
  assign n32538 = ~n20778 & n32537 ;
  assign n32539 = n20886 & n32538 ;
  assign n32540 = ~\pi0760  & n1689 ;
  assign n32541 = n20784 & n32540 ;
  assign n32542 = n22767 & n32541 ;
  assign n32543 = ~\pi0178  & ~n1689 ;
  assign n32544 = ~n32541 & ~n32543 ;
  assign n32545 = ~n20792 & ~n32544 ;
  assign n32546 = ~n32542 & n32545 ;
  assign n32547 = n20801 & ~n32546 ;
  assign n32548 = ~\pi1155  & ~n32543 ;
  assign n32549 = \pi0785  & n32548 ;
  assign n32550 = ~n32542 & n32549 ;
  assign n32551 = ~\pi0785  & ~n32543 ;
  assign n32552 = ~n32541 & n32551 ;
  assign n32553 = ~n20804 & ~n32552 ;
  assign n32554 = n29682 & n32553 ;
  assign n32555 = ~n32550 & n32554 ;
  assign n32556 = ~n32547 & n32555 ;
  assign n32557 = n30847 & n32556 ;
  assign n32558 = ~n32539 & ~n32557 ;
  assign n32559 = ~\pi0688  & n1689 ;
  assign n32560 = n20855 & n32559 ;
  assign n32561 = ~n32543 & ~n32560 ;
  assign n32562 = ~\pi0778  & ~n32561 ;
  assign n32563 = ~\pi0625  & ~\pi0688  ;
  assign n32564 = n1689 & n32563 ;
  assign n32565 = n20855 & n32564 ;
  assign n32566 = \pi1153  & n32565 ;
  assign n32567 = \pi1153  & ~n32543 ;
  assign n32568 = ~n32560 & n32567 ;
  assign n32569 = ~n32566 & ~n32568 ;
  assign n32570 = ~\pi1153  & ~n32543 ;
  assign n32571 = ~n32565 & n32570 ;
  assign n32572 = \pi0778  & ~n32571 ;
  assign n32573 = n32569 & n32572 ;
  assign n32574 = ~n32562 & ~n32573 ;
  assign n32575 = n26474 & ~n32574 ;
  assign n32576 = \pi0629  & ~n32575 ;
  assign n32577 = n32558 & n32576 ;
  assign n32578 = n20887 & n32538 ;
  assign n32579 = n20887 & ~n23880 ;
  assign n32580 = n32556 & n32579 ;
  assign n32581 = ~n32578 & ~n32580 ;
  assign n32582 = n26485 & ~n32574 ;
  assign n32583 = ~\pi0629  & ~n32582 ;
  assign n32584 = n32581 & n32583 ;
  assign n32585 = \pi0792  & ~n32584 ;
  assign n32586 = ~n32577 & n32585 ;
  assign n32587 = ~n21067 & ~n32586 ;
  assign n32588 = n26325 & ~n32574 ;
  assign n32589 = ~\pi0178  & ~\pi0647  ;
  assign n32590 = ~n1689 & n32589 ;
  assign n32591 = n20849 & ~n32590 ;
  assign n32592 = ~n32588 & n32591 ;
  assign n32593 = n26319 & ~n32574 ;
  assign n32594 = ~\pi0178  & \pi0647  ;
  assign n32595 = ~n1689 & n32594 ;
  assign n32596 = n20897 & ~n32595 ;
  assign n32597 = ~n32593 & n32596 ;
  assign n32598 = ~n32592 & ~n32597 ;
  assign n32599 = \pi0787  & ~n32598 ;
  assign n32600 = ~n20846 & n32538 ;
  assign n32601 = n30376 & n32556 ;
  assign n32602 = ~n32600 & ~n32601 ;
  assign n32603 = ~\pi0178  & \pi0792  ;
  assign n32604 = ~n1689 & n32603 ;
  assign n32605 = ~n20845 & n32604 ;
  assign n32606 = \pi0787  & ~n20910 ;
  assign n32607 = ~n32605 & n32606 ;
  assign n32608 = n32602 & n32607 ;
  assign n32609 = ~n32599 & ~n32608 ;
  assign n32610 = ~n24761 & n32609 ;
  assign n32611 = ~n32587 & n32610 ;
  assign n32612 = \pi0608  & ~n32571 ;
  assign n32613 = ~n32541 & n32567 ;
  assign n32614 = \pi0778  & ~n32613 ;
  assign n32615 = n26421 & ~n32561 ;
  assign n32616 = ~n32614 & ~n32615 ;
  assign n32617 = n32612 & ~n32616 ;
  assign n32618 = n26147 & ~n32561 ;
  assign n32619 = ~\pi0688  & ~n20784 ;
  assign n32620 = n22113 & n32619 ;
  assign n32621 = n32544 & ~n32620 ;
  assign n32622 = ~n32618 & ~n32621 ;
  assign n32623 = n32570 & ~n32622 ;
  assign n32624 = n26415 & n32569 ;
  assign n32625 = ~n32623 & n32624 ;
  assign n32626 = ~n32617 & ~n32625 ;
  assign n32627 = ~\pi1155  & ~n32562 ;
  assign n32628 = ~n32573 & n32627 ;
  assign n32629 = ~n20999 & ~n32628 ;
  assign n32630 = ~\pi0778  & ~n32621 ;
  assign n32631 = ~n32629 & ~n32630 ;
  assign n32632 = n32626 & n32631 ;
  assign n32633 = n29766 & ~n32562 ;
  assign n32634 = ~n32573 & n32633 ;
  assign n32635 = \pi1155  & ~n32546 ;
  assign n32636 = ~\pi0660  & ~n32635 ;
  assign n32637 = ~n32634 & n32636 ;
  assign n32638 = ~n32632 & n32637 ;
  assign n32639 = \pi0785  & ~n32638 ;
  assign n32640 = n29775 & n32553 ;
  assign n32641 = ~n32550 & n32640 ;
  assign n32642 = ~n32547 & n32641 ;
  assign n32643 = n29779 & ~n32574 ;
  assign n32644 = ~n32642 & ~n32643 ;
  assign n32645 = \pi0781  & ~n32644 ;
  assign n32646 = \pi1155  & ~n32562 ;
  assign n32647 = ~n32573 & n32646 ;
  assign n32648 = ~n21774 & ~n32647 ;
  assign n32649 = ~n32630 & ~n32648 ;
  assign n32650 = n32626 & n32649 ;
  assign n32651 = n26121 & ~n32562 ;
  assign n32652 = ~n32573 & n32651 ;
  assign n32653 = \pi0660  & ~n32548 ;
  assign n32654 = \pi0660  & n32541 ;
  assign n32655 = n22767 & n32654 ;
  assign n32656 = ~n32653 & ~n32655 ;
  assign n32657 = ~n32652 & ~n32656 ;
  assign n32658 = ~n32650 & n32657 ;
  assign n32659 = ~n32645 & ~n32658 ;
  assign n32660 = n32639 & n32659 ;
  assign n32661 = ~\pi0785  & ~n32630 ;
  assign n32662 = ~n32617 & n32661 ;
  assign n32663 = ~n32625 & n32662 ;
  assign n32664 = n21022 & ~n32663 ;
  assign n32665 = ~n32645 & ~n32664 ;
  assign n32666 = n29803 & ~n32665 ;
  assign n32667 = ~n32660 & n32666 ;
  assign n32668 = n29808 & n32553 ;
  assign n32669 = ~n32550 & n32668 ;
  assign n32670 = ~n32547 & n32669 ;
  assign n32671 = n30966 & ~n32574 ;
  assign n32672 = ~n32670 & ~n32671 ;
  assign n32673 = n29818 & ~n32672 ;
  assign n32674 = \pi0626  & ~n32556 ;
  assign n32675 = ~\pi0626  & ~n32543 ;
  assign n32676 = n20881 & ~n32675 ;
  assign n32677 = ~n32674 & n32676 ;
  assign n32678 = n26458 & ~n32574 ;
  assign n32679 = ~\pi0626  & ~n32556 ;
  assign n32680 = \pi0626  & ~n32543 ;
  assign n32681 = n20882 & ~n32680 ;
  assign n32682 = ~n32679 & n32681 ;
  assign n32683 = ~n32678 & ~n32682 ;
  assign n32684 = ~n32677 & n32683 ;
  assign n32685 = \pi0788  & ~n32684 ;
  assign n32686 = ~n32673 & ~n32685 ;
  assign n32687 = ~n32667 & n32686 ;
  assign n32688 = ~n23856 & n32610 ;
  assign n32689 = ~n32687 & n32688 ;
  assign n32690 = ~n32611 & ~n32689 ;
  assign n32691 = n30987 & ~n32602 ;
  assign n32692 = n23312 & n32691 ;
  assign n32693 = \pi1157  & ~n32590 ;
  assign n32694 = ~n32588 & n32693 ;
  assign n32695 = ~\pi1157  & ~n32595 ;
  assign n32696 = ~n32593 & n32695 ;
  assign n32697 = ~n32694 & ~n32696 ;
  assign n32698 = \pi0787  & ~n32697 ;
  assign n32699 = n26333 & ~n32574 ;
  assign n32700 = ~\pi0787  & ~n32699 ;
  assign n32701 = ~\pi1160  & ~n32700 ;
  assign n32702 = n23312 & n32701 ;
  assign n32703 = ~n32698 & n32702 ;
  assign n32704 = ~n32692 & ~n32703 ;
  assign n32705 = \pi0790  & ~n32704 ;
  assign n32706 = \pi1160  & ~n32700 ;
  assign n32707 = ~n32698 & n32706 ;
  assign n32708 = ~n23414 & n32543 ;
  assign n32709 = ~n24886 & n32708 ;
  assign n32710 = n31010 & ~n32602 ;
  assign n32711 = ~n32709 & ~n32710 ;
  assign n32712 = ~n32707 & n32711 ;
  assign n32713 = ~n23313 & ~n32708 ;
  assign n32714 = ~n31019 & ~n32713 ;
  assign n32715 = \pi0790  & n32714 ;
  assign n32716 = ~n32712 & n32715 ;
  assign n32717 = ~n32705 & ~n32716 ;
  assign n32718 = \pi0832  & n32717 ;
  assign n32719 = n32690 & n32718 ;
  assign n32720 = \pi0178  & ~\pi0832  ;
  assign n32721 = ~n21132 & ~n32720 ;
  assign n32722 = ~n32719 & n32721 ;
  assign n32723 = n9948 & ~n32719 ;
  assign n32724 = ~n32722 & ~n32723 ;
  assign n32725 = \pi0178  & ~n6861 ;
  assign n32726 = ~n20985 & n32725 ;
  assign n32727 = n21774 & n32726 ;
  assign n32728 = \pi0038  & n32541 ;
  assign n32729 = n8413 & n32728 ;
  assign n32730 = n1354 & n32729 ;
  assign n32731 = n1358 & n32730 ;
  assign n32732 = \pi0038  & ~\pi0178  ;
  assign n32733 = ~n21757 & n32732 ;
  assign n32734 = ~n32731 & ~n32733 ;
  assign n32735 = \pi0038  & n32734 ;
  assign n32736 = ~\pi0178  & ~n21467 ;
  assign n32737 = ~\pi0039  & ~\pi0178  ;
  assign n32738 = n21272 & n32737 ;
  assign n32739 = ~n32736 & ~n32738 ;
  assign n32740 = ~\pi0178  & ~\pi0760  ;
  assign n32741 = ~\pi0760  & ~n21566 ;
  assign n32742 = n21484 & n32741 ;
  assign n32743 = ~n32740 & ~n32742 ;
  assign n32744 = n32739 & ~n32743 ;
  assign n32745 = ~\pi0178  & \pi0760  ;
  assign n32746 = n21743 & n32745 ;
  assign n32747 = ~n21734 & n32746 ;
  assign n32748 = n32734 & ~n32747 ;
  assign n32749 = ~n32744 & n32748 ;
  assign n32750 = ~n32735 & ~n32749 ;
  assign n32751 = n26646 & ~n32750 ;
  assign n32752 = ~n32727 & ~n32751 ;
  assign n32753 = ~\pi0178  & n21768 ;
  assign n32754 = ~\pi0178  & n21770 ;
  assign n32755 = ~n21734 & n32754 ;
  assign n32756 = ~n32753 & ~n32755 ;
  assign n32757 = \pi1155  & ~n20790 ;
  assign n32758 = n20789 & n32757 ;
  assign n32759 = ~n26121 & ~n32758 ;
  assign n32760 = n32756 & ~n32759 ;
  assign n32761 = ~\pi0660  & ~n32760 ;
  assign n32762 = n32752 & n32761 ;
  assign n32763 = n20999 & n32726 ;
  assign n32764 = n26685 & ~n32750 ;
  assign n32765 = ~n32763 & ~n32764 ;
  assign n32766 = ~\pi1155  & ~n20790 ;
  assign n32767 = n20789 & n32766 ;
  assign n32768 = ~n29766 & ~n32767 ;
  assign n32769 = n32756 & ~n32768 ;
  assign n32770 = \pi0660  & ~n32769 ;
  assign n32771 = n32765 & n32770 ;
  assign n32772 = ~n32762 & ~n32771 ;
  assign n32773 = \pi0688  & n32750 ;
  assign n32774 = ~\pi0178  & ~\pi0625  ;
  assign n32775 = ~n22734 & ~n32774 ;
  assign n32776 = n32773 & ~n32775 ;
  assign n32777 = ~\pi0178  & n23548 ;
  assign n32778 = ~\pi0760  & ~n32777 ;
  assign n32779 = ~\pi0039  & ~\pi0760  ;
  assign n32780 = ~n22683 & n32779 ;
  assign n32781 = ~n32778 & ~n32780 ;
  assign n32782 = ~\pi0038  & n32781 ;
  assign n32783 = ~\pi0038  & \pi0178  ;
  assign n32784 = ~n26538 & n32783 ;
  assign n32785 = ~n32782 & ~n32784 ;
  assign n32786 = ~\pi0178  & ~n23567 ;
  assign n32787 = n23565 & n32786 ;
  assign n32788 = \pi0760  & n23575 ;
  assign n32789 = n23572 & n32788 ;
  assign n32790 = ~n32745 & ~n32789 ;
  assign n32791 = ~n32787 & ~n32790 ;
  assign n32792 = ~n32785 & ~n32791 ;
  assign n32793 = n6861 & n32792 ;
  assign n32794 = ~\pi0178  & ~\pi0688  ;
  assign n32795 = ~n26566 & n32794 ;
  assign n32796 = ~\pi0760  & n32794 ;
  assign n32797 = ~n22536 & n32796 ;
  assign n32798 = ~n32795 & ~n32797 ;
  assign n32799 = \pi0688  & n6861 ;
  assign n32800 = \pi0178  & ~\pi0760  ;
  assign n32801 = n1689 & n32800 ;
  assign n32802 = n20784 & n32801 ;
  assign n32803 = \pi0178  & ~n20784 ;
  assign n32804 = n22113 & n32803 ;
  assign n32805 = ~n32802 & ~n32804 ;
  assign n32806 = n26554 & ~n32805 ;
  assign n32807 = n1358 & n32806 ;
  assign n32808 = \pi0038  & n6861 ;
  assign n32809 = ~n32807 & n32808 ;
  assign n32810 = ~n32799 & ~n32809 ;
  assign n32811 = n32798 & ~n32810 ;
  assign n32812 = ~n32775 & ~n32811 ;
  assign n32813 = ~n32793 & n32812 ;
  assign n32814 = ~n32776 & ~n32813 ;
  assign n32815 = n6861 & ~n32750 ;
  assign n32816 = ~\pi0178  & \pi0625  ;
  assign n32817 = ~n22727 & ~n32816 ;
  assign n32818 = ~n32815 & ~n32817 ;
  assign n32819 = ~\pi1153  & ~n32818 ;
  assign n32820 = n32814 & n32819 ;
  assign n32821 = ~\pi0074  & ~\pi0688  ;
  assign n32822 = ~\pi0100  & n32821 ;
  assign n32823 = n1287 & n32822 ;
  assign n32824 = ~\pi0178  & ~n32823 ;
  assign n32825 = n21768 & n32824 ;
  assign n32826 = n21770 & n32824 ;
  assign n32827 = ~n21734 & n32826 ;
  assign n32828 = ~n32825 & ~n32827 ;
  assign n32829 = \pi0625  & ~n32828 ;
  assign n32830 = ~\pi0038  & ~\pi0178  ;
  assign n32831 = n6861 & ~n32830 ;
  assign n32832 = ~n22109 & n32831 ;
  assign n32833 = ~\pi0178  & ~n22017 ;
  assign n32834 = ~n21994 & n32833 ;
  assign n32835 = ~n32832 & ~n32834 ;
  assign n32836 = ~\pi0178  & ~n21757 ;
  assign n32837 = n22117 & ~n32836 ;
  assign n32838 = ~\pi0688  & ~n32837 ;
  assign n32839 = \pi0625  & n32838 ;
  assign n32840 = ~n32835 & n32839 ;
  assign n32841 = ~n32829 & ~n32840 ;
  assign n32842 = n21768 & n32774 ;
  assign n32843 = n21770 & n32774 ;
  assign n32844 = ~n21734 & n32843 ;
  assign n32845 = ~n32842 & ~n32844 ;
  assign n32846 = \pi1153  & n32845 ;
  assign n32847 = n32841 & n32846 ;
  assign n32848 = ~\pi0608  & ~n32847 ;
  assign n32849 = ~n32820 & n32848 ;
  assign n32850 = n32773 & ~n32817 ;
  assign n32851 = ~n32811 & ~n32817 ;
  assign n32852 = ~n32793 & n32851 ;
  assign n32853 = ~n32850 & ~n32852 ;
  assign n32854 = \pi1153  & n32775 ;
  assign n32855 = n23606 & ~n32750 ;
  assign n32856 = ~n32854 & ~n32855 ;
  assign n32857 = n32853 & ~n32856 ;
  assign n32858 = ~\pi0625  & ~n32828 ;
  assign n32859 = ~\pi0625  & n32838 ;
  assign n32860 = ~n32835 & n32859 ;
  assign n32861 = ~n32858 & ~n32860 ;
  assign n32862 = n21768 & n32816 ;
  assign n32863 = n21770 & n32816 ;
  assign n32864 = ~n21734 & n32863 ;
  assign n32865 = ~n32862 & ~n32864 ;
  assign n32866 = ~\pi1153  & n32865 ;
  assign n32867 = n32861 & n32866 ;
  assign n32868 = \pi0608  & ~n32867 ;
  assign n32869 = ~n32857 & n32868 ;
  assign n32870 = ~n32849 & ~n32869 ;
  assign n32871 = n23638 & ~n32870 ;
  assign n32872 = ~\pi0178  & ~\pi0778  ;
  assign n32873 = ~n23622 & ~n32872 ;
  assign n32874 = n32773 & ~n32873 ;
  assign n32875 = ~n32811 & ~n32873 ;
  assign n32876 = ~n32793 & n32875 ;
  assign n32877 = ~n32874 & ~n32876 ;
  assign n32878 = \pi0609  & ~n32877 ;
  assign n32879 = ~n32835 & n32838 ;
  assign n32880 = ~\pi0778  & n32828 ;
  assign n32881 = ~n32879 & n32880 ;
  assign n32882 = ~\pi0609  & ~n32881 ;
  assign n32883 = \pi1155  & ~n32882 ;
  assign n32884 = ~n32847 & ~n32867 ;
  assign n32885 = n22722 & ~n32884 ;
  assign n32886 = ~n32883 & ~n32885 ;
  assign n32887 = ~n32762 & ~n32886 ;
  assign n32888 = ~n32878 & n32887 ;
  assign n32889 = ~n32871 & n32888 ;
  assign n32890 = ~n32772 & ~n32889 ;
  assign n32891 = \pi0778  & ~n32870 ;
  assign n32892 = \pi0778  & ~n32884 ;
  assign n32893 = \pi0609  & ~n32881 ;
  assign n32894 = ~n32892 & n32893 ;
  assign n32895 = ~\pi1155  & n32726 ;
  assign n32896 = n26672 & ~n32750 ;
  assign n32897 = ~n32895 & ~n32896 ;
  assign n32898 = ~\pi0609  & ~n32897 ;
  assign n32899 = ~n22787 & ~n32769 ;
  assign n32900 = ~n32898 & n32899 ;
  assign n32901 = ~n32894 & ~n32900 ;
  assign n32902 = \pi0785  & ~n32901 ;
  assign n32903 = n32877 & ~n32902 ;
  assign n32904 = ~n32891 & n32903 ;
  assign n32905 = \pi0609  & ~n32899 ;
  assign n32906 = n32881 & n32905 ;
  assign n32907 = \pi0778  & n32905 ;
  assign n32908 = ~n32884 & n32907 ;
  assign n32909 = ~n32906 & ~n32908 ;
  assign n32910 = ~n32904 & n32909 ;
  assign n32911 = n32890 & n32910 ;
  assign n32912 = ~\pi0785  & ~n32904 ;
  assign n32913 = n26700 & ~n32912 ;
  assign n32914 = ~n32911 & n32913 ;
  assign n32915 = n23456 & ~n32750 ;
  assign n32916 = n21777 & n32725 ;
  assign n32917 = ~n21777 & n32756 ;
  assign n32918 = n20811 & ~n32917 ;
  assign n32919 = ~n32916 & n32918 ;
  assign n32920 = ~n32915 & n32919 ;
  assign n32921 = ~n20811 & ~n32756 ;
  assign n32922 = n22155 & ~n32921 ;
  assign n32923 = ~n32920 & n32922 ;
  assign n32924 = ~n21034 & n32923 ;
  assign n32925 = ~n22147 & ~n32881 ;
  assign n32926 = ~n32892 & n32925 ;
  assign n32927 = n22147 & ~n32756 ;
  assign n32928 = n24348 & ~n32927 ;
  assign n32929 = ~n21034 & n32928 ;
  assign n32930 = ~n32926 & n32929 ;
  assign n32931 = ~n32924 & ~n32930 ;
  assign n32932 = ~n32920 & ~n32921 ;
  assign n32933 = n23424 & ~n32932 ;
  assign n32934 = ~\pi0781  & ~n32917 ;
  assign n32935 = ~n23423 & ~n32916 ;
  assign n32936 = n32934 & n32935 ;
  assign n32937 = ~n32915 & n32936 ;
  assign n32938 = n23423 & ~n32756 ;
  assign n32939 = ~n32937 & ~n32938 ;
  assign n32940 = ~n32933 & n32939 ;
  assign n32941 = ~n23880 & ~n32940 ;
  assign n32942 = n23880 & ~n32756 ;
  assign n32943 = n24691 & ~n32942 ;
  assign n32944 = ~n32941 & n32943 ;
  assign n32945 = n26065 & ~n32884 ;
  assign n32946 = n26739 & n32828 ;
  assign n32947 = ~n32879 & n32946 ;
  assign n32948 = ~n23885 & n32756 ;
  assign n32949 = \pi0628  & ~n32948 ;
  assign n32950 = ~n32947 & n32949 ;
  assign n32951 = ~n32945 & n32950 ;
  assign n32952 = ~\pi0178  & ~\pi0628  ;
  assign n32953 = n21768 & n32952 ;
  assign n32954 = n21770 & n32952 ;
  assign n32955 = ~n21734 & n32954 ;
  assign n32956 = ~n32953 & ~n32955 ;
  assign n32957 = \pi1156  & n32956 ;
  assign n32958 = ~\pi0629  & n32957 ;
  assign n32959 = ~n32951 & n32958 ;
  assign n32960 = ~\pi0628  & ~n32948 ;
  assign n32961 = ~n32947 & n32960 ;
  assign n32962 = ~n32945 & n32961 ;
  assign n32963 = ~\pi0178  & \pi0628  ;
  assign n32964 = n21768 & n32963 ;
  assign n32965 = n21770 & n32963 ;
  assign n32966 = ~n21734 & n32965 ;
  assign n32967 = ~n32964 & ~n32966 ;
  assign n32968 = ~\pi1156  & n32967 ;
  assign n32969 = \pi0629  & n32968 ;
  assign n32970 = ~n32962 & n32969 ;
  assign n32971 = ~n32959 & ~n32970 ;
  assign n32972 = ~n32944 & n32971 ;
  assign n32973 = \pi0792  & ~n32972 ;
  assign n32974 = n23380 & ~n32881 ;
  assign n32975 = ~n23380 & ~n32756 ;
  assign n32976 = n21050 & ~n32975 ;
  assign n32977 = ~n32974 & n32976 ;
  assign n32978 = \pi0778  & n32976 ;
  assign n32979 = ~n32884 & n32978 ;
  assign n32980 = ~n32977 & ~n32979 ;
  assign n32981 = \pi0789  & ~n32980 ;
  assign n32982 = n23683 & ~n32932 ;
  assign n32983 = n21032 & ~n32916 ;
  assign n32984 = n32934 & n32983 ;
  assign n32985 = ~n32915 & n32984 ;
  assign n32986 = ~n21032 & ~n32756 ;
  assign n32987 = ~n20876 & ~n32986 ;
  assign n32988 = ~n32985 & n32987 ;
  assign n32989 = \pi0789  & n32988 ;
  assign n32990 = ~n32982 & n32989 ;
  assign n32991 = ~n32981 & ~n32990 ;
  assign n32992 = ~n21038 & n32991 ;
  assign n32993 = ~n32973 & n32992 ;
  assign n32994 = n32931 & n32993 ;
  assign n32995 = ~n32914 & n32994 ;
  assign n32996 = ~n22160 & ~n32975 ;
  assign n32997 = ~n32974 & n32996 ;
  assign n32998 = \pi0778  & n32996 ;
  assign n32999 = ~n32884 & n32998 ;
  assign n33000 = ~n32997 & ~n32999 ;
  assign n33001 = n22160 & n32756 ;
  assign n33002 = n20951 & ~n33001 ;
  assign n33003 = n33000 & n33002 ;
  assign n33004 = ~\pi0626  & ~n32938 ;
  assign n33005 = ~n32937 & n33004 ;
  assign n33006 = ~n32933 & n33005 ;
  assign n33007 = \pi0626  & n32756 ;
  assign n33008 = n20882 & ~n33007 ;
  assign n33009 = ~n33006 & n33008 ;
  assign n33010 = ~n33003 & ~n33009 ;
  assign n33011 = \pi0626  & ~n32938 ;
  assign n33012 = ~n32937 & n33011 ;
  assign n33013 = ~n32933 & n33012 ;
  assign n33014 = ~\pi0626  & n32756 ;
  assign n33015 = n20881 & ~n33014 ;
  assign n33016 = ~n33013 & n33015 ;
  assign n33017 = ~n23856 & ~n33016 ;
  assign n33018 = n33010 & n33017 ;
  assign n33019 = ~n26803 & ~n33018 ;
  assign n33020 = ~n32973 & n33019 ;
  assign n33021 = ~n21067 & ~n33020 ;
  assign n33022 = ~n32995 & n33021 ;
  assign n33023 = ~n31367 & ~n32756 ;
  assign n33024 = ~\pi0715  & ~n33023 ;
  assign n33025 = ~n23958 & ~n33024 ;
  assign n33026 = n31382 & ~n32940 ;
  assign n33027 = ~n33025 & ~n33026 ;
  assign n33028 = n26824 & ~n33027 ;
  assign n33029 = ~\pi0178  & \pi0644  ;
  assign n33030 = n21768 & n33029 ;
  assign n33031 = n21770 & n33029 ;
  assign n33032 = ~n21734 & n33031 ;
  assign n33033 = ~n33030 & ~n33032 ;
  assign n33034 = n23939 & n33033 ;
  assign n33035 = \pi0715  & n33033 ;
  assign n33036 = ~n33023 & n33035 ;
  assign n33037 = ~n33034 & ~n33036 ;
  assign n33038 = n31367 & ~n33034 ;
  assign n33039 = ~n32940 & n33038 ;
  assign n33040 = ~n33037 & ~n33039 ;
  assign n33041 = n31378 & ~n33040 ;
  assign n33042 = \pi0790  & ~n33041 ;
  assign n33043 = ~n33028 & n33042 ;
  assign n33044 = ~n32947 & ~n32948 ;
  assign n33045 = ~n32945 & n33044 ;
  assign n33046 = ~\pi0792  & ~n33045 ;
  assign n33047 = \pi0647  & ~n33046 ;
  assign n33048 = n21768 & n32589 ;
  assign n33049 = n21770 & n32589 ;
  assign n33050 = ~n21734 & n33049 ;
  assign n33051 = ~n33048 & ~n33050 ;
  assign n33052 = \pi1157  & n33051 ;
  assign n33053 = ~n33047 & n33052 ;
  assign n33054 = ~n32951 & n32957 ;
  assign n33055 = ~n32962 & n32968 ;
  assign n33056 = ~n33054 & ~n33055 ;
  assign n33057 = \pi0792  & n33052 ;
  assign n33058 = ~n33056 & n33057 ;
  assign n33059 = ~n33053 & ~n33058 ;
  assign n33060 = ~\pi0630  & ~n33059 ;
  assign n33061 = ~\pi0647  & ~n33046 ;
  assign n33062 = n21768 & n32594 ;
  assign n33063 = n21770 & n32594 ;
  assign n33064 = ~n21734 & n33063 ;
  assign n33065 = ~n33062 & ~n33064 ;
  assign n33066 = ~\pi1157  & n33065 ;
  assign n33067 = ~n33061 & n33066 ;
  assign n33068 = \pi0792  & n33066 ;
  assign n33069 = ~n33056 & n33068 ;
  assign n33070 = ~n33067 & ~n33069 ;
  assign n33071 = \pi0630  & ~n33070 ;
  assign n33072 = ~n20846 & n32942 ;
  assign n33073 = n30376 & ~n32940 ;
  assign n33074 = ~n33072 & ~n33073 ;
  assign n33075 = n20846 & ~n32756 ;
  assign n33076 = ~n20910 & ~n33075 ;
  assign n33077 = n33074 & n33076 ;
  assign n33078 = ~n33071 & ~n33077 ;
  assign n33079 = ~n33060 & n33078 ;
  assign n33080 = \pi0787  & ~n33079 ;
  assign n33081 = ~n33043 & ~n33080 ;
  assign n33082 = ~n33022 & n33081 ;
  assign n33083 = ~\pi0787  & n33046 ;
  assign n33084 = ~\pi0787  & \pi0792  ;
  assign n33085 = ~n33056 & n33084 ;
  assign n33086 = ~n33083 & ~n33085 ;
  assign n33087 = ~\pi0644  & n33086 ;
  assign n33088 = \pi0715  & ~n33087 ;
  assign n33089 = n33059 & n33070 ;
  assign n33090 = n26918 & ~n33089 ;
  assign n33091 = ~n33088 & ~n33090 ;
  assign n33092 = ~\pi0644  & ~n32756 ;
  assign n33093 = n33027 & ~n33092 ;
  assign n33094 = \pi1160  & ~n33093 ;
  assign n33095 = n33091 & n33094 ;
  assign n33096 = \pi0644  & n33086 ;
  assign n33097 = ~\pi0715  & ~n33096 ;
  assign n33098 = ~\pi0715  & \pi0787  ;
  assign n33099 = ~n33089 & n33098 ;
  assign n33100 = ~n33097 & ~n33099 ;
  assign n33101 = ~\pi1160  & ~n33040 ;
  assign n33102 = n33100 & n33101 ;
  assign n33103 = ~n33095 & ~n33102 ;
  assign n33104 = \pi0790  & ~n33103 ;
  assign n33105 = ~n32722 & ~n33104 ;
  assign n33106 = ~n33082 & n33105 ;
  assign n33107 = ~n32724 & ~n33106 ;
  assign n33108 = ~\pi0179  & ~n1689 ;
  assign n33109 = ~n21032 & ~n33108 ;
  assign n33110 = \pi0789  & n33109 ;
  assign n33111 = ~n23880 & ~n33110 ;
  assign n33112 = n23423 & n33111 ;
  assign n33113 = ~\pi0741  & n1689 ;
  assign n33114 = n20784 & n33113 ;
  assign n33115 = ~n33108 & ~n33114 ;
  assign n33116 = n20794 & ~n33115 ;
  assign n33117 = n20796 & ~n33116 ;
  assign n33118 = n20799 & ~n33115 ;
  assign n33119 = n20801 & ~n33118 ;
  assign n33120 = ~n33117 & ~n33119 ;
  assign n33121 = ~\pi0785  & ~n33108 ;
  assign n33122 = ~n33114 & n33121 ;
  assign n33123 = ~n20804 & ~n33122 ;
  assign n33124 = ~n20812 & n33123 ;
  assign n33125 = n33111 & n33124 ;
  assign n33126 = n33120 & n33125 ;
  assign n33127 = ~n33112 & ~n33126 ;
  assign n33128 = ~\pi0179  & \pi0788  ;
  assign n33129 = ~n1689 & n33128 ;
  assign n33130 = ~n20778 & n33129 ;
  assign n33131 = ~\pi0179  & \pi0792  ;
  assign n33132 = ~n1689 & n33131 ;
  assign n33133 = ~n20845 & n33132 ;
  assign n33134 = ~n20910 & ~n33133 ;
  assign n33135 = ~n33130 & n33134 ;
  assign n33136 = n33127 & n33135 ;
  assign n33137 = n20846 & n33134 ;
  assign n33138 = ~\pi0724  & n1689 ;
  assign n33139 = n20855 & n33138 ;
  assign n33140 = ~n20861 & n33139 ;
  assign n33141 = ~n33108 & ~n33140 ;
  assign n33142 = n20879 & ~n33141 ;
  assign n33143 = n20895 & n33142 ;
  assign n33144 = ~\pi0179  & \pi0647  ;
  assign n33145 = ~n1689 & n33144 ;
  assign n33146 = n20897 & ~n33145 ;
  assign n33147 = ~n33143 & n33146 ;
  assign n33148 = ~\pi0179  & ~\pi0647  ;
  assign n33149 = ~n1689 & n33148 ;
  assign n33150 = n20849 & ~n33149 ;
  assign n33151 = ~n24761 & ~n33150 ;
  assign n33152 = n31479 & n33142 ;
  assign n33153 = ~n33151 & ~n33152 ;
  assign n33154 = ~n33147 & ~n33153 ;
  assign n33155 = ~n33137 & n33154 ;
  assign n33156 = ~n33136 & n33155 ;
  assign n33157 = ~n29722 & ~n33156 ;
  assign n33158 = n23423 & ~n33110 ;
  assign n33159 = ~n33110 & n33124 ;
  assign n33160 = n33120 & n33159 ;
  assign n33161 = ~n33158 & ~n33160 ;
  assign n33162 = ~\pi0626  & n33161 ;
  assign n33163 = \pi0626  & ~n33108 ;
  assign n33164 = n20882 & ~n33163 ;
  assign n33165 = ~n33162 & n33164 ;
  assign n33166 = n23170 & ~n33141 ;
  assign n33167 = ~\pi0626  & ~n33108 ;
  assign n33168 = n20881 & ~n33167 ;
  assign n33169 = ~n33166 & ~n33168 ;
  assign n33170 = \pi0626  & ~n33166 ;
  assign n33171 = n33161 & n33170 ;
  assign n33172 = ~n33169 & ~n33171 ;
  assign n33173 = ~n33165 & ~n33172 ;
  assign n33174 = \pi0788  & ~n33173 ;
  assign n33175 = ~n23856 & n33174 ;
  assign n33176 = ~\pi0724  & n20855 ;
  assign n33177 = ~n20861 & n33176 ;
  assign n33178 = ~n20986 & n33177 ;
  assign n33179 = ~\pi0741  & n20784 ;
  assign n33180 = ~n20985 & n33179 ;
  assign n33181 = ~n33108 & ~n33180 ;
  assign n33182 = ~n33178 & n33181 ;
  assign n33183 = \pi0179  & ~n1689 ;
  assign n33184 = ~\pi0609  & ~n33183 ;
  assign n33185 = ~n33182 & n33184 ;
  assign n33186 = ~\pi1155  & ~n33108 ;
  assign n33187 = ~n33140 & n33186 ;
  assign n33188 = ~n20999 & ~n33187 ;
  assign n33189 = ~n33185 & ~n33188 ;
  assign n33190 = \pi1155  & ~n33118 ;
  assign n33191 = ~\pi0660  & ~n33190 ;
  assign n33192 = ~n33189 & n33191 ;
  assign n33193 = ~n21007 & ~n33117 ;
  assign n33194 = \pi0609  & ~n33183 ;
  assign n33195 = ~n33182 & n33194 ;
  assign n33196 = \pi1155  & ~n33108 ;
  assign n33197 = ~n33140 & n33196 ;
  assign n33198 = ~n21774 & ~n33197 ;
  assign n33199 = \pi0785  & ~n33198 ;
  assign n33200 = ~n33195 & n33199 ;
  assign n33201 = n33193 & ~n33200 ;
  assign n33202 = ~n33192 & ~n33201 ;
  assign n33203 = ~n33182 & ~n33183 ;
  assign n33204 = ~\pi0785  & ~n33203 ;
  assign n33205 = n21022 & ~n33204 ;
  assign n33206 = ~n33202 & n33205 ;
  assign n33207 = n20964 & n33123 ;
  assign n33208 = n33120 & n33207 ;
  assign n33209 = \pi0627  & ~n33108 ;
  assign n33210 = ~n33140 & n33209 ;
  assign n33211 = ~n20968 & ~n33210 ;
  assign n33212 = ~n33208 & ~n33211 ;
  assign n33213 = n20974 & n33123 ;
  assign n33214 = n33120 & n33213 ;
  assign n33215 = ~\pi0627  & ~n33108 ;
  assign n33216 = ~n33140 & n33215 ;
  assign n33217 = ~n20978 & ~n33216 ;
  assign n33218 = ~n33214 & ~n33217 ;
  assign n33219 = ~n33212 & ~n33218 ;
  assign n33220 = \pi0781  & n33219 ;
  assign n33221 = ~n21034 & ~n33220 ;
  assign n33222 = ~n33206 & n33221 ;
  assign n33223 = ~n20876 & n33109 ;
  assign n33224 = ~n24969 & ~n33223 ;
  assign n33225 = n33124 & ~n33223 ;
  assign n33226 = n33120 & n33225 ;
  assign n33227 = ~n33224 & ~n33226 ;
  assign n33228 = n21050 & ~n33108 ;
  assign n33229 = ~n33140 & n33228 ;
  assign n33230 = ~n21051 & ~n33229 ;
  assign n33231 = ~n21038 & n33230 ;
  assign n33232 = ~n33227 & n33231 ;
  assign n33233 = ~n23177 & ~n33232 ;
  assign n33234 = ~n23856 & ~n33233 ;
  assign n33235 = ~n33222 & n33234 ;
  assign n33236 = ~n33175 & ~n33235 ;
  assign n33237 = ~n33157 & ~n33236 ;
  assign n33238 = n24830 & n33142 ;
  assign n33239 = \pi1157  & ~n33149 ;
  assign n33240 = ~n33238 & n33239 ;
  assign n33241 = ~\pi1157  & ~n33145 ;
  assign n33242 = ~n33143 & n33241 ;
  assign n33243 = ~n33240 & ~n33242 ;
  assign n33244 = \pi0787  & ~n33243 ;
  assign n33245 = n24844 & n33142 ;
  assign n33246 = ~n24843 & ~n33245 ;
  assign n33247 = ~n33244 & ~n33246 ;
  assign n33248 = n33127 & ~n33130 ;
  assign n33249 = n31580 & ~n33248 ;
  assign n33250 = ~n33247 & ~n33249 ;
  assign n33251 = n23313 & ~n33250 ;
  assign n33252 = \pi0790  & n33251 ;
  assign n33253 = n31588 & ~n33248 ;
  assign n33254 = ~n23414 & n33108 ;
  assign n33255 = ~n24886 & n33254 ;
  assign n33256 = n20891 & n33142 ;
  assign n33257 = ~\pi0787  & ~n33256 ;
  assign n33258 = ~\pi1160  & ~n33257 ;
  assign n33259 = ~n33244 & n33258 ;
  assign n33260 = ~n33255 & ~n33259 ;
  assign n33261 = ~n33253 & n33260 ;
  assign n33262 = ~n23312 & ~n33254 ;
  assign n33263 = ~n31603 & ~n33262 ;
  assign n33264 = \pi0790  & n33263 ;
  assign n33265 = ~n33261 & n33264 ;
  assign n33266 = ~n33252 & ~n33265 ;
  assign n33267 = n20938 & n33142 ;
  assign n33268 = \pi0629  & ~n33130 ;
  assign n33269 = ~n33267 & n33268 ;
  assign n33270 = n33127 & n33269 ;
  assign n33271 = n21077 & n33142 ;
  assign n33272 = ~\pi0629  & ~n33130 ;
  assign n33273 = ~n33271 & n33272 ;
  assign n33274 = n33127 & n33273 ;
  assign n33275 = n29714 & ~n33267 ;
  assign n33276 = n29709 & ~n33271 ;
  assign n33277 = \pi0792  & ~n33276 ;
  assign n33278 = ~n33275 & n33277 ;
  assign n33279 = ~n33274 & n33278 ;
  assign n33280 = ~n33270 & n33279 ;
  assign n33281 = ~n21067 & ~n33280 ;
  assign n33282 = ~n33157 & ~n33281 ;
  assign n33283 = \pi0832  & ~n33282 ;
  assign n33284 = n33266 & n33283 ;
  assign n33285 = ~n33237 & n33284 ;
  assign n33286 = \pi0179  & ~\pi0832  ;
  assign n33287 = ~n21132 & ~n33286 ;
  assign n33288 = ~n33285 & n33287 ;
  assign n33289 = ~\pi0179  & n21768 ;
  assign n33290 = ~\pi0179  & n21770 ;
  assign n33291 = ~n21734 & n33290 ;
  assign n33292 = ~n33289 & ~n33291 ;
  assign n33293 = ~n22849 & n33292 ;
  assign n33294 = ~n22161 & ~n23907 ;
  assign n33295 = n33293 & n33294 ;
  assign n33296 = ~\pi0074  & ~\pi0724  ;
  assign n33297 = ~\pi0100  & n33296 ;
  assign n33298 = n1287 & n33297 ;
  assign n33299 = ~\pi0179  & ~n33298 ;
  assign n33300 = n21768 & n33299 ;
  assign n33301 = n21770 & n33299 ;
  assign n33302 = ~n21734 & n33301 ;
  assign n33303 = ~n33300 & ~n33302 ;
  assign n33304 = ~\pi0625  & ~n33303 ;
  assign n33305 = ~\pi0179  & ~n22017 ;
  assign n33306 = ~n21994 & n33305 ;
  assign n33307 = ~\pi0038  & ~\pi0179  ;
  assign n33308 = n6861 & ~n33307 ;
  assign n33309 = ~n22109 & n33308 ;
  assign n33310 = ~n33306 & ~n33309 ;
  assign n33311 = ~\pi0179  & ~n21757 ;
  assign n33312 = n22117 & ~n33311 ;
  assign n33313 = ~\pi0724  & ~n33312 ;
  assign n33314 = ~\pi0625  & n33313 ;
  assign n33315 = ~n33310 & n33314 ;
  assign n33316 = ~n33304 & ~n33315 ;
  assign n33317 = ~\pi0179  & \pi0625  ;
  assign n33318 = n21768 & n33317 ;
  assign n33319 = n21770 & n33317 ;
  assign n33320 = ~n21734 & n33319 ;
  assign n33321 = ~n33318 & ~n33320 ;
  assign n33322 = ~\pi1153  & n33321 ;
  assign n33323 = n33316 & n33322 ;
  assign n33324 = \pi0625  & ~n33303 ;
  assign n33325 = \pi0625  & n33313 ;
  assign n33326 = ~n33310 & n33325 ;
  assign n33327 = ~n33324 & ~n33326 ;
  assign n33328 = ~\pi0179  & ~\pi0625  ;
  assign n33329 = n21768 & n33328 ;
  assign n33330 = n21770 & n33328 ;
  assign n33331 = ~n21734 & n33330 ;
  assign n33332 = ~n33329 & ~n33331 ;
  assign n33333 = \pi1153  & n33332 ;
  assign n33334 = n33327 & n33333 ;
  assign n33335 = ~n33323 & ~n33334 ;
  assign n33336 = n22148 & ~n33335 ;
  assign n33337 = ~n33310 & n33313 ;
  assign n33338 = n22151 & n33303 ;
  assign n33339 = ~n33337 & n33338 ;
  assign n33340 = n22147 & n33292 ;
  assign n33341 = ~n33339 & ~n33340 ;
  assign n33342 = ~n33336 & n33341 ;
  assign n33343 = n22849 & n33294 ;
  assign n33344 = ~n33342 & n33343 ;
  assign n33345 = ~n33295 & ~n33344 ;
  assign n33346 = n33292 & ~n33294 ;
  assign n33347 = \pi0644  & ~n33346 ;
  assign n33348 = n33345 & n33347 ;
  assign n33349 = ~n23074 & ~n33348 ;
  assign n33350 = ~\pi0715  & n33349 ;
  assign n33351 = \pi0647  & ~n33346 ;
  assign n33352 = n33345 & n33351 ;
  assign n33353 = n21768 & n33148 ;
  assign n33354 = n21770 & n33148 ;
  assign n33355 = ~n21734 & n33354 ;
  assign n33356 = ~n33353 & ~n33355 ;
  assign n33357 = \pi1157  & n33356 ;
  assign n33358 = ~n33352 & n33357 ;
  assign n33359 = ~\pi0647  & ~n33346 ;
  assign n33360 = n33345 & n33359 ;
  assign n33361 = n21768 & n33144 ;
  assign n33362 = n21770 & n33144 ;
  assign n33363 = ~n21734 & n33362 ;
  assign n33364 = ~n33361 & ~n33363 ;
  assign n33365 = ~\pi1157  & n33364 ;
  assign n33366 = ~n33360 & n33365 ;
  assign n33367 = ~n33358 & ~n33366 ;
  assign n33368 = n33098 & ~n33367 ;
  assign n33369 = ~n33350 & ~n33368 ;
  assign n33370 = ~\pi0179  & \pi0644  ;
  assign n33371 = n21768 & n33370 ;
  assign n33372 = n21770 & n33370 ;
  assign n33373 = ~n21734 & n33372 ;
  assign n33374 = ~n33371 & ~n33373 ;
  assign n33375 = \pi0715  & n33374 ;
  assign n33376 = ~\pi1160  & ~n33375 ;
  assign n33377 = n23880 & ~n33292 ;
  assign n33378 = ~\pi0179  & \pi0618  ;
  assign n33379 = n21768 & n33378 ;
  assign n33380 = n21770 & n33378 ;
  assign n33381 = ~n21734 & n33380 ;
  assign n33382 = ~n33379 & ~n33381 ;
  assign n33383 = ~\pi1154  & n33382 ;
  assign n33384 = \pi0781  & ~n33383 ;
  assign n33385 = \pi0179  & ~n6861 ;
  assign n33386 = n21777 & n33385 ;
  assign n33387 = ~n23456 & ~n33386 ;
  assign n33388 = \pi0179  & \pi0741  ;
  assign n33389 = \pi0179  & ~n25040 ;
  assign n33390 = ~n33388 & ~n33389 ;
  assign n33391 = ~\pi0038  & ~n33388 ;
  assign n33392 = n25023 & n33391 ;
  assign n33393 = ~n33390 & ~n33392 ;
  assign n33394 = ~\pi0179  & ~\pi0741  ;
  assign n33395 = ~n25033 & n33394 ;
  assign n33396 = ~n25040 & n33395 ;
  assign n33397 = ~n25028 & n33396 ;
  assign n33398 = ~n33393 & ~n33397 ;
  assign n33399 = ~n28149 & ~n33386 ;
  assign n33400 = n33398 & n33399 ;
  assign n33401 = ~n33387 & ~n33400 ;
  assign n33402 = ~n21777 & n33292 ;
  assign n33403 = ~\pi0618  & ~n33402 ;
  assign n33404 = \pi0781  & n33403 ;
  assign n33405 = ~n33401 & n33404 ;
  assign n33406 = ~n33384 & ~n33405 ;
  assign n33407 = \pi0618  & ~n33402 ;
  assign n33408 = ~n33401 & n33407 ;
  assign n33409 = ~\pi0179  & ~\pi0618  ;
  assign n33410 = n21768 & n33409 ;
  assign n33411 = n21770 & n33409 ;
  assign n33412 = ~n21734 & n33411 ;
  assign n33413 = ~n33410 & ~n33412 ;
  assign n33414 = \pi1154  & n33413 ;
  assign n33415 = ~n33408 & n33414 ;
  assign n33416 = ~n33406 & ~n33415 ;
  assign n33417 = ~\pi0781  & ~n33402 ;
  assign n33418 = ~n33401 & n33417 ;
  assign n33419 = ~\pi0789  & ~n33418 ;
  assign n33420 = ~n33416 & n33419 ;
  assign n33421 = ~n23880 & ~n33420 ;
  assign n33422 = n21092 & ~n33421 ;
  assign n33423 = ~\pi0619  & ~n33414 ;
  assign n33424 = ~\pi0619  & n33407 ;
  assign n33425 = ~n33401 & n33424 ;
  assign n33426 = ~n33423 & ~n33425 ;
  assign n33427 = ~n33406 & ~n33426 ;
  assign n33428 = ~\pi0619  & n33417 ;
  assign n33429 = ~n33401 & n33428 ;
  assign n33430 = ~\pi0179  & \pi0619  ;
  assign n33431 = n21768 & n33430 ;
  assign n33432 = n21770 & n33430 ;
  assign n33433 = ~n21734 & n33432 ;
  assign n33434 = ~n33431 & ~n33433 ;
  assign n33435 = ~\pi1159  & n33434 ;
  assign n33436 = ~n33429 & n33435 ;
  assign n33437 = ~n33427 & n33436 ;
  assign n33438 = ~\pi0179  & ~\pi0619  ;
  assign n33439 = n21768 & n33438 ;
  assign n33440 = n21770 & n33438 ;
  assign n33441 = ~n21734 & n33440 ;
  assign n33442 = ~n33439 & ~n33441 ;
  assign n33443 = \pi1159  & n33442 ;
  assign n33444 = ~\pi0619  & n33443 ;
  assign n33445 = ~n33418 & n33443 ;
  assign n33446 = ~n33416 & n33445 ;
  assign n33447 = ~n33444 & ~n33446 ;
  assign n33448 = ~n33437 & n33447 ;
  assign n33449 = n32328 & ~n33448 ;
  assign n33450 = ~n33422 & ~n33449 ;
  assign n33451 = ~n33377 & ~n33450 ;
  assign n33452 = ~n21092 & n33292 ;
  assign n33453 = n31378 & ~n33452 ;
  assign n33454 = ~n33451 & n33453 ;
  assign n33455 = ~n33376 & ~n33454 ;
  assign n33456 = n33369 & ~n33455 ;
  assign n33457 = \pi0644  & ~n33452 ;
  assign n33458 = ~n33451 & n33457 ;
  assign n33459 = ~\pi0179  & ~\pi0644  ;
  assign n33460 = n21768 & n33459 ;
  assign n33461 = n21770 & n33459 ;
  assign n33462 = ~n21734 & n33461 ;
  assign n33463 = ~n33460 & ~n33462 ;
  assign n33464 = ~\pi0715  & n33463 ;
  assign n33465 = ~n33458 & n33464 ;
  assign n33466 = ~\pi0644  & ~n33346 ;
  assign n33467 = n33345 & n33466 ;
  assign n33468 = ~n23021 & ~n33467 ;
  assign n33469 = \pi0715  & n33468 ;
  assign n33470 = n26918 & ~n33367 ;
  assign n33471 = ~n33469 & ~n33470 ;
  assign n33472 = \pi1160  & n33471 ;
  assign n33473 = ~n33465 & n33472 ;
  assign n33474 = ~n33456 & ~n33473 ;
  assign n33475 = \pi0790  & ~n33474 ;
  assign n33476 = n31378 & ~n33375 ;
  assign n33477 = ~n33454 & ~n33476 ;
  assign n33478 = n26824 & ~n33452 ;
  assign n33479 = ~n33451 & n33478 ;
  assign n33480 = \pi0715  & n26824 ;
  assign n33481 = \pi0790  & ~n33480 ;
  assign n33482 = ~n33479 & n33481 ;
  assign n33483 = n33477 & n33482 ;
  assign n33484 = \pi0619  & \pi1159  ;
  assign n33485 = ~n22155 & ~n33340 ;
  assign n33486 = ~n33339 & n33485 ;
  assign n33487 = ~n33336 & n33486 ;
  assign n33488 = n22155 & ~n33292 ;
  assign n33489 = \pi1159  & ~n33488 ;
  assign n33490 = ~n33487 & n33489 ;
  assign n33491 = ~n33484 & ~n33490 ;
  assign n33492 = \pi0648  & ~n33437 ;
  assign n33493 = n33491 & n33492 ;
  assign n33494 = \pi0789  & n33493 ;
  assign n33495 = ~\pi0648  & n33447 ;
  assign n33496 = ~\pi1159  & ~n33488 ;
  assign n33497 = ~n33487 & n33496 ;
  assign n33498 = ~n22872 & ~n33497 ;
  assign n33499 = \pi0789  & n33498 ;
  assign n33500 = n33495 & n33499 ;
  assign n33501 = ~n33494 & ~n33500 ;
  assign n33502 = ~\pi0618  & ~n33340 ;
  assign n33503 = ~n33339 & n33502 ;
  assign n33504 = ~n33336 & n33503 ;
  assign n33505 = \pi1154  & ~n33504 ;
  assign n33506 = \pi0627  & ~n33383 ;
  assign n33507 = \pi0627  & n33403 ;
  assign n33508 = ~n33401 & n33507 ;
  assign n33509 = ~n33506 & ~n33508 ;
  assign n33510 = ~n33505 & ~n33509 ;
  assign n33511 = \pi0618  & ~n33340 ;
  assign n33512 = ~n33339 & n33511 ;
  assign n33513 = ~n33336 & n33512 ;
  assign n33514 = ~\pi1154  & ~n33513 ;
  assign n33515 = ~\pi0627  & ~n33414 ;
  assign n33516 = ~\pi0627  & n33407 ;
  assign n33517 = ~n33401 & n33516 ;
  assign n33518 = ~n33515 & ~n33517 ;
  assign n33519 = ~n33514 & ~n33518 ;
  assign n33520 = ~n33510 & ~n33519 ;
  assign n33521 = n32123 & ~n33443 ;
  assign n33522 = \pi0789  & ~n32121 ;
  assign n33523 = n31279 & n33434 ;
  assign n33524 = ~n33522 & ~n33523 ;
  assign n33525 = ~n33521 & ~n33524 ;
  assign n33526 = \pi0781  & ~n33525 ;
  assign n33527 = ~n33520 & n33526 ;
  assign n33528 = n33501 & ~n33527 ;
  assign n33529 = ~n21038 & ~n33528 ;
  assign n33530 = \pi0724  & ~n33393 ;
  assign n33531 = ~n33397 & n33530 ;
  assign n33532 = ~n28149 & n33531 ;
  assign n33533 = n6861 & ~n33532 ;
  assign n33534 = ~n22727 & ~n33317 ;
  assign n33535 = ~n33533 & ~n33534 ;
  assign n33536 = n23587 & ~n33311 ;
  assign n33537 = \pi0741  & ~n33536 ;
  assign n33538 = \pi0038  & n33537 ;
  assign n33539 = \pi0179  & n23575 ;
  assign n33540 = ~n23571 & n33539 ;
  assign n33541 = ~n23570 & n33537 ;
  assign n33542 = n33540 & n33541 ;
  assign n33543 = ~n33538 & ~n33542 ;
  assign n33544 = ~\pi0179  & \pi0741  ;
  assign n33545 = ~n33536 & n33544 ;
  assign n33546 = ~n23568 & n33545 ;
  assign n33547 = n33543 & ~n33546 ;
  assign n33548 = \pi0038  & \pi0179  ;
  assign n33549 = ~n22708 & n33548 ;
  assign n33550 = ~\pi0038  & \pi0179  ;
  assign n33551 = ~n33549 & ~n33550 ;
  assign n33552 = ~n23558 & ~n33549 ;
  assign n33553 = n23557 & n33552 ;
  assign n33554 = ~n33551 & ~n33553 ;
  assign n33555 = ~\pi0179  & n23548 ;
  assign n33556 = ~n25191 & n33555 ;
  assign n33557 = ~n25190 & n33556 ;
  assign n33558 = ~\pi0741  & ~n33557 ;
  assign n33559 = ~n33554 & n33558 ;
  assign n33560 = n33547 & ~n33559 ;
  assign n33561 = ~\pi0724  & ~n33534 ;
  assign n33562 = ~n33560 & n33561 ;
  assign n33563 = ~n33535 & ~n33562 ;
  assign n33564 = ~n22734 & ~n33328 ;
  assign n33565 = ~n6861 & ~n33564 ;
  assign n33566 = ~n28149 & ~n33564 ;
  assign n33567 = n33398 & n33566 ;
  assign n33568 = ~n33565 & ~n33567 ;
  assign n33569 = \pi1153  & n33568 ;
  assign n33570 = n33563 & n33569 ;
  assign n33571 = \pi0608  & ~n33323 ;
  assign n33572 = ~n33570 & n33571 ;
  assign n33573 = ~n33533 & ~n33564 ;
  assign n33574 = ~\pi0724  & ~n33564 ;
  assign n33575 = ~n33560 & n33574 ;
  assign n33576 = ~n33573 & ~n33575 ;
  assign n33577 = ~n6861 & ~n33534 ;
  assign n33578 = ~n28149 & ~n33534 ;
  assign n33579 = n33398 & n33578 ;
  assign n33580 = ~n33577 & ~n33579 ;
  assign n33581 = ~\pi1153  & n33580 ;
  assign n33582 = n33576 & n33581 ;
  assign n33583 = ~\pi0608  & ~n33334 ;
  assign n33584 = ~n33582 & n33583 ;
  assign n33585 = ~n33572 & ~n33584 ;
  assign n33586 = n23613 & ~n33585 ;
  assign n33587 = \pi0778  & ~n33335 ;
  assign n33588 = ~\pi0778  & n33303 ;
  assign n33589 = ~n33337 & n33588 ;
  assign n33590 = \pi0609  & ~n33589 ;
  assign n33591 = ~n33587 & n33590 ;
  assign n33592 = ~\pi0179  & ~\pi0778  ;
  assign n33593 = ~n23622 & ~n33592 ;
  assign n33594 = ~n33533 & ~n33593 ;
  assign n33595 = ~\pi0724  & ~n33593 ;
  assign n33596 = ~n33560 & n33595 ;
  assign n33597 = ~n33594 & ~n33596 ;
  assign n33598 = ~\pi0609  & ~n33597 ;
  assign n33599 = ~\pi1155  & ~n33598 ;
  assign n33600 = ~n33591 & n33599 ;
  assign n33601 = ~n33586 & n33600 ;
  assign n33602 = ~n20985 & n33385 ;
  assign n33603 = ~n26645 & ~n33602 ;
  assign n33604 = ~n28149 & ~n33602 ;
  assign n33605 = n33398 & n33604 ;
  assign n33606 = ~n33603 & ~n33605 ;
  assign n33607 = n21774 & n33606 ;
  assign n33608 = ~n32759 & n33292 ;
  assign n33609 = ~\pi0660  & ~n33608 ;
  assign n33610 = ~n33607 & n33609 ;
  assign n33611 = ~n33601 & n33610 ;
  assign n33612 = n20999 & n33606 ;
  assign n33613 = ~n32768 & n33292 ;
  assign n33614 = \pi0660  & ~n33613 ;
  assign n33615 = ~n33612 & n33614 ;
  assign n33616 = \pi0785  & ~n33615 ;
  assign n33617 = \pi0609  & ~n33597 ;
  assign n33618 = ~\pi0609  & ~n33589 ;
  assign n33619 = \pi1155  & ~n33618 ;
  assign n33620 = n22722 & ~n33335 ;
  assign n33621 = ~n33619 & ~n33620 ;
  assign n33622 = \pi0785  & ~n33621 ;
  assign n33623 = ~n33617 & n33622 ;
  assign n33624 = ~n33616 & ~n33623 ;
  assign n33625 = n23638 & ~n33616 ;
  assign n33626 = ~n33585 & n33625 ;
  assign n33627 = ~n33624 & ~n33626 ;
  assign n33628 = ~n33611 & n33627 ;
  assign n33629 = n21019 & ~n33383 ;
  assign n33630 = \pi0781  & ~n21016 ;
  assign n33631 = n21020 & n33413 ;
  assign n33632 = ~n33630 & ~n33631 ;
  assign n33633 = ~n33629 & ~n33632 ;
  assign n33634 = ~\pi0785  & n33597 ;
  assign n33635 = ~n33525 & ~n33634 ;
  assign n33636 = \pi0778  & ~n33525 ;
  assign n33637 = ~n33585 & n33636 ;
  assign n33638 = ~n33635 & ~n33637 ;
  assign n33639 = ~n33633 & ~n33638 ;
  assign n33640 = ~n21038 & n33639 ;
  assign n33641 = ~n33628 & n33640 ;
  assign n33642 = ~n33529 & ~n33641 ;
  assign n33643 = ~\pi0789  & ~n33420 ;
  assign n33644 = ~n33420 & ~n33437 ;
  assign n33645 = n33447 & n33644 ;
  assign n33646 = ~n33643 & ~n33645 ;
  assign n33647 = n30606 & ~n33646 ;
  assign n33648 = ~\pi0641  & n33293 ;
  assign n33649 = ~\pi0641  & n22849 ;
  assign n33650 = ~n33342 & n33649 ;
  assign n33651 = ~n33648 & ~n33650 ;
  assign n33652 = \pi0641  & n33292 ;
  assign n33653 = n20777 & ~n33652 ;
  assign n33654 = n33651 & n33653 ;
  assign n33655 = \pi0641  & n33293 ;
  assign n33656 = \pi0641  & n22849 ;
  assign n33657 = ~n33342 & n33656 ;
  assign n33658 = ~n33655 & ~n33657 ;
  assign n33659 = ~\pi0641  & n33292 ;
  assign n33660 = n20776 & ~n33659 ;
  assign n33661 = n33658 & n33660 ;
  assign n33662 = ~n23856 & ~n33661 ;
  assign n33663 = ~n33654 & n33662 ;
  assign n33664 = ~n33647 & n33663 ;
  assign n33665 = ~n26803 & ~n33664 ;
  assign n33666 = ~n21067 & ~n33665 ;
  assign n33667 = n33642 & n33666 ;
  assign n33668 = ~n30376 & n33292 ;
  assign n33669 = ~n20910 & n33668 ;
  assign n33670 = ~n20910 & n30376 ;
  assign n33671 = n33646 & n33670 ;
  assign n33672 = ~n33669 & ~n33671 ;
  assign n33673 = ~\pi0630  & n33357 ;
  assign n33674 = ~n33352 & n33673 ;
  assign n33675 = \pi0630  & n33365 ;
  assign n33676 = ~n33360 & n33675 ;
  assign n33677 = ~n33674 & ~n33676 ;
  assign n33678 = n33672 & n33677 ;
  assign n33679 = \pi0787  & ~n33678 ;
  assign n33680 = ~n33377 & ~n33421 ;
  assign n33681 = \pi0789  & ~n33377 ;
  assign n33682 = ~n33448 & n33681 ;
  assign n33683 = ~n33680 & ~n33682 ;
  assign n33684 = n24691 & ~n33683 ;
  assign n33685 = n22162 & ~n33488 ;
  assign n33686 = ~n33487 & n33685 ;
  assign n33687 = ~n22162 & n33292 ;
  assign n33688 = \pi0628  & ~n33687 ;
  assign n33689 = ~n33686 & n33688 ;
  assign n33690 = ~\pi0179  & ~\pi0628  ;
  assign n33691 = n21768 & n33690 ;
  assign n33692 = n21770 & n33690 ;
  assign n33693 = ~n21734 & n33692 ;
  assign n33694 = ~n33691 & ~n33693 ;
  assign n33695 = n20843 & n33694 ;
  assign n33696 = ~n33689 & n33695 ;
  assign n33697 = ~\pi0628  & ~n33687 ;
  assign n33698 = ~n33686 & n33697 ;
  assign n33699 = ~\pi0179  & \pi0628  ;
  assign n33700 = n21768 & n33699 ;
  assign n33701 = n21770 & n33699 ;
  assign n33702 = ~n21734 & n33701 ;
  assign n33703 = ~n33700 & ~n33702 ;
  assign n33704 = n20844 & n33703 ;
  assign n33705 = ~n33698 & n33704 ;
  assign n33706 = ~n33696 & ~n33705 ;
  assign n33707 = ~n33684 & n33706 ;
  assign n33708 = n24724 & ~n33707 ;
  assign n33709 = ~n33679 & ~n33708 ;
  assign n33710 = ~n33667 & n33709 ;
  assign n33711 = ~n33483 & n33710 ;
  assign n33712 = ~n33475 & ~n33711 ;
  assign n33713 = n9948 & ~n33285 ;
  assign n33714 = ~n33712 & n33713 ;
  assign n33715 = ~n33288 & ~n33714 ;
  assign n33716 = ~\pi0180  & \pi0788  ;
  assign n33717 = ~n1689 & n33716 ;
  assign n33718 = ~n20778 & n33717 ;
  assign n33719 = n20886 & n33718 ;
  assign n33720 = ~\pi0753  & n1689 ;
  assign n33721 = n20784 & n33720 ;
  assign n33722 = n22767 & n33721 ;
  assign n33723 = ~\pi0180  & ~n1689 ;
  assign n33724 = ~n33721 & ~n33723 ;
  assign n33725 = ~n20792 & ~n33724 ;
  assign n33726 = ~n33722 & n33725 ;
  assign n33727 = n20801 & ~n33726 ;
  assign n33728 = ~\pi1155  & ~n33723 ;
  assign n33729 = \pi0785  & n33728 ;
  assign n33730 = ~n33722 & n33729 ;
  assign n33731 = ~\pi0785  & ~n33723 ;
  assign n33732 = ~n33721 & n33731 ;
  assign n33733 = ~n20804 & ~n33732 ;
  assign n33734 = n29682 & n33733 ;
  assign n33735 = ~n33730 & n33734 ;
  assign n33736 = ~n33727 & n33735 ;
  assign n33737 = n30847 & n33736 ;
  assign n33738 = ~n33719 & ~n33737 ;
  assign n33739 = ~\pi0702  & n1689 ;
  assign n33740 = n20855 & n33739 ;
  assign n33741 = ~n33723 & ~n33740 ;
  assign n33742 = ~\pi0778  & ~n33741 ;
  assign n33743 = ~\pi0625  & ~\pi0702  ;
  assign n33744 = n1689 & n33743 ;
  assign n33745 = n20855 & n33744 ;
  assign n33746 = \pi1153  & n33745 ;
  assign n33747 = \pi1153  & ~n33723 ;
  assign n33748 = ~n33740 & n33747 ;
  assign n33749 = ~n33746 & ~n33748 ;
  assign n33750 = ~\pi1153  & ~n33723 ;
  assign n33751 = ~n33745 & n33750 ;
  assign n33752 = \pi0778  & ~n33751 ;
  assign n33753 = n33749 & n33752 ;
  assign n33754 = ~n33742 & ~n33753 ;
  assign n33755 = n26474 & ~n33754 ;
  assign n33756 = \pi0629  & ~n33755 ;
  assign n33757 = n33738 & n33756 ;
  assign n33758 = n20887 & n33718 ;
  assign n33759 = n32579 & n33736 ;
  assign n33760 = ~n33758 & ~n33759 ;
  assign n33761 = n26485 & ~n33754 ;
  assign n33762 = ~\pi0629  & ~n33761 ;
  assign n33763 = n33760 & n33762 ;
  assign n33764 = ~n33757 & ~n33763 ;
  assign n33765 = \pi0792  & n33764 ;
  assign n33766 = ~n21067 & ~n33765 ;
  assign n33767 = n26325 & ~n33754 ;
  assign n33768 = ~\pi0180  & ~\pi0647  ;
  assign n33769 = ~n1689 & n33768 ;
  assign n33770 = n20849 & ~n33769 ;
  assign n33771 = ~n33767 & n33770 ;
  assign n33772 = n26319 & ~n33754 ;
  assign n33773 = ~\pi0180  & \pi0647  ;
  assign n33774 = ~n1689 & n33773 ;
  assign n33775 = n20897 & ~n33774 ;
  assign n33776 = ~n33772 & n33775 ;
  assign n33777 = ~n33771 & ~n33776 ;
  assign n33778 = \pi0787  & ~n33777 ;
  assign n33779 = ~n20846 & n33718 ;
  assign n33780 = n30376 & n33736 ;
  assign n33781 = ~n33779 & ~n33780 ;
  assign n33782 = ~\pi0180  & \pi0792  ;
  assign n33783 = ~n1689 & n33782 ;
  assign n33784 = ~n20845 & n33783 ;
  assign n33785 = n32606 & ~n33784 ;
  assign n33786 = n33781 & n33785 ;
  assign n33787 = ~n33778 & ~n33786 ;
  assign n33788 = ~n24761 & n33787 ;
  assign n33789 = ~n33766 & n33788 ;
  assign n33790 = \pi0608  & ~n33751 ;
  assign n33791 = ~n33721 & n33747 ;
  assign n33792 = \pi0778  & ~n33791 ;
  assign n33793 = n26421 & ~n33741 ;
  assign n33794 = ~n33792 & ~n33793 ;
  assign n33795 = n33790 & ~n33794 ;
  assign n33796 = n26147 & ~n33741 ;
  assign n33797 = ~\pi0702  & ~n20784 ;
  assign n33798 = n22113 & n33797 ;
  assign n33799 = n33724 & ~n33798 ;
  assign n33800 = ~n33796 & ~n33799 ;
  assign n33801 = n33750 & ~n33800 ;
  assign n33802 = n26415 & n33749 ;
  assign n33803 = ~n33801 & n33802 ;
  assign n33804 = ~n33795 & ~n33803 ;
  assign n33805 = ~\pi1155  & ~n33742 ;
  assign n33806 = ~n33753 & n33805 ;
  assign n33807 = ~n20999 & ~n33806 ;
  assign n33808 = ~\pi0778  & ~n33799 ;
  assign n33809 = ~n33807 & ~n33808 ;
  assign n33810 = n33804 & n33809 ;
  assign n33811 = n29766 & ~n33742 ;
  assign n33812 = ~n33753 & n33811 ;
  assign n33813 = \pi1155  & ~n33726 ;
  assign n33814 = ~\pi0660  & ~n33813 ;
  assign n33815 = ~n33812 & n33814 ;
  assign n33816 = ~n33810 & n33815 ;
  assign n33817 = \pi0785  & ~n33816 ;
  assign n33818 = n29775 & n33733 ;
  assign n33819 = ~n33730 & n33818 ;
  assign n33820 = ~n33727 & n33819 ;
  assign n33821 = n29779 & ~n33754 ;
  assign n33822 = ~n33820 & ~n33821 ;
  assign n33823 = \pi0781  & ~n33822 ;
  assign n33824 = \pi1155  & ~n33742 ;
  assign n33825 = ~n33753 & n33824 ;
  assign n33826 = ~n21774 & ~n33825 ;
  assign n33827 = ~n33808 & ~n33826 ;
  assign n33828 = n33804 & n33827 ;
  assign n33829 = n26121 & ~n33742 ;
  assign n33830 = ~n33753 & n33829 ;
  assign n33831 = \pi0660  & ~n33728 ;
  assign n33832 = \pi0660  & n33721 ;
  assign n33833 = n22767 & n33832 ;
  assign n33834 = ~n33831 & ~n33833 ;
  assign n33835 = ~n33830 & ~n33834 ;
  assign n33836 = ~n33828 & n33835 ;
  assign n33837 = ~n33823 & ~n33836 ;
  assign n33838 = n33817 & n33837 ;
  assign n33839 = ~\pi0785  & ~n33808 ;
  assign n33840 = ~n33795 & n33839 ;
  assign n33841 = ~n33803 & n33840 ;
  assign n33842 = n21022 & ~n33841 ;
  assign n33843 = ~n33823 & ~n33842 ;
  assign n33844 = n29803 & ~n33843 ;
  assign n33845 = ~n33838 & n33844 ;
  assign n33846 = n29808 & n33733 ;
  assign n33847 = ~n33730 & n33846 ;
  assign n33848 = ~n33727 & n33847 ;
  assign n33849 = n30966 & ~n33754 ;
  assign n33850 = ~n33848 & ~n33849 ;
  assign n33851 = n29818 & ~n33850 ;
  assign n33852 = \pi0626  & ~n33736 ;
  assign n33853 = ~\pi0626  & ~n33723 ;
  assign n33854 = n20881 & ~n33853 ;
  assign n33855 = ~n33852 & n33854 ;
  assign n33856 = n26458 & ~n33754 ;
  assign n33857 = ~\pi0626  & ~n33736 ;
  assign n33858 = \pi0626  & ~n33723 ;
  assign n33859 = n20882 & ~n33858 ;
  assign n33860 = ~n33857 & n33859 ;
  assign n33861 = ~n33856 & ~n33860 ;
  assign n33862 = ~n33855 & n33861 ;
  assign n33863 = \pi0788  & ~n33862 ;
  assign n33864 = ~n33851 & ~n33863 ;
  assign n33865 = ~n33845 & n33864 ;
  assign n33866 = ~n23856 & n33788 ;
  assign n33867 = ~n33865 & n33866 ;
  assign n33868 = ~n33789 & ~n33867 ;
  assign n33869 = n30987 & ~n33781 ;
  assign n33870 = n23312 & n33869 ;
  assign n33871 = \pi1157  & ~n33769 ;
  assign n33872 = ~n33767 & n33871 ;
  assign n33873 = ~\pi1157  & ~n33774 ;
  assign n33874 = ~n33772 & n33873 ;
  assign n33875 = ~n33872 & ~n33874 ;
  assign n33876 = \pi0787  & ~n33875 ;
  assign n33877 = n26333 & ~n33754 ;
  assign n33878 = ~\pi0787  & ~n33877 ;
  assign n33879 = ~\pi1160  & ~n33878 ;
  assign n33880 = n23312 & n33879 ;
  assign n33881 = ~n33876 & n33880 ;
  assign n33882 = ~n33870 & ~n33881 ;
  assign n33883 = \pi0790  & ~n33882 ;
  assign n33884 = \pi1160  & ~n33878 ;
  assign n33885 = ~n33876 & n33884 ;
  assign n33886 = ~n23414 & n33723 ;
  assign n33887 = ~n24886 & n33886 ;
  assign n33888 = n31010 & ~n33781 ;
  assign n33889 = ~n33887 & ~n33888 ;
  assign n33890 = ~n33885 & n33889 ;
  assign n33891 = ~n23313 & ~n33886 ;
  assign n33892 = ~n31019 & ~n33891 ;
  assign n33893 = \pi0790  & n33892 ;
  assign n33894 = ~n33890 & n33893 ;
  assign n33895 = ~n33883 & ~n33894 ;
  assign n33896 = \pi0832  & n33895 ;
  assign n33897 = n33868 & n33896 ;
  assign n33898 = \pi0180  & ~\pi0832  ;
  assign n33899 = ~n21132 & ~n33898 ;
  assign n33900 = ~n33897 & n33899 ;
  assign n33901 = n9948 & ~n33897 ;
  assign n33902 = ~n33900 & ~n33901 ;
  assign n33903 = \pi0038  & n33721 ;
  assign n33904 = n8413 & n33903 ;
  assign n33905 = n1354 & n33904 ;
  assign n33906 = n1358 & n33905 ;
  assign n33907 = \pi0038  & ~\pi0180  ;
  assign n33908 = ~n21757 & n33907 ;
  assign n33909 = ~n33906 & ~n33908 ;
  assign n33910 = ~\pi0180  & \pi0753  ;
  assign n33911 = n21743 & n33910 ;
  assign n33912 = ~n21734 & n33911 ;
  assign n33913 = ~\pi0038  & n33912 ;
  assign n33914 = \pi0180  & ~n25023 ;
  assign n33915 = ~\pi0180  & ~n21467 ;
  assign n33916 = ~\pi0753  & ~n33915 ;
  assign n33917 = ~n33914 & n33916 ;
  assign n33918 = ~\pi0039  & ~\pi0180  ;
  assign n33919 = n21272 & n33918 ;
  assign n33920 = ~\pi0038  & ~n33919 ;
  assign n33921 = n33917 & n33920 ;
  assign n33922 = ~n33913 & ~n33921 ;
  assign n33923 = n33909 & n33922 ;
  assign n33924 = \pi0702  & ~n33923 ;
  assign n33925 = ~\pi0180  & ~\pi0778  ;
  assign n33926 = ~n23622 & ~n33925 ;
  assign n33927 = n33924 & ~n33926 ;
  assign n33928 = ~\pi0180  & n23548 ;
  assign n33929 = ~\pi0753  & ~n33928 ;
  assign n33930 = ~\pi0039  & ~\pi0753  ;
  assign n33931 = ~n22683 & n33930 ;
  assign n33932 = ~n33929 & ~n33931 ;
  assign n33933 = ~\pi0038  & n33932 ;
  assign n33934 = ~\pi0038  & \pi0180  ;
  assign n33935 = ~n26538 & n33934 ;
  assign n33936 = ~n33933 & ~n33935 ;
  assign n33937 = ~\pi0180  & ~n23567 ;
  assign n33938 = n23565 & n33937 ;
  assign n33939 = \pi0753  & n23575 ;
  assign n33940 = n23572 & n33939 ;
  assign n33941 = ~n33910 & ~n33940 ;
  assign n33942 = ~n33938 & ~n33941 ;
  assign n33943 = ~n33936 & ~n33942 ;
  assign n33944 = n6861 & n33943 ;
  assign n33945 = \pi0180  & ~\pi0753  ;
  assign n33946 = n1689 & n33945 ;
  assign n33947 = n20784 & n33946 ;
  assign n33948 = \pi0180  & ~n20784 ;
  assign n33949 = n22113 & n33948 ;
  assign n33950 = ~n33947 & ~n33949 ;
  assign n33951 = n26554 & ~n33950 ;
  assign n33952 = n1358 & n33951 ;
  assign n33953 = \pi0038  & ~n33952 ;
  assign n33954 = ~\pi0702  & ~n33953 ;
  assign n33955 = ~\pi0180  & ~\pi0702  ;
  assign n33956 = ~n26566 & n33955 ;
  assign n33957 = ~\pi0753  & n33955 ;
  assign n33958 = ~n22536 & n33957 ;
  assign n33959 = ~n33956 & ~n33958 ;
  assign n33960 = ~n33954 & n33959 ;
  assign n33961 = n6861 & n33960 ;
  assign n33962 = ~n33926 & ~n33961 ;
  assign n33963 = ~n33944 & n33962 ;
  assign n33964 = ~n33927 & ~n33963 ;
  assign n33965 = \pi0609  & ~n33964 ;
  assign n33966 = ~\pi0180  & ~\pi0625  ;
  assign n33967 = ~n22734 & ~n33966 ;
  assign n33968 = n33924 & ~n33967 ;
  assign n33969 = ~n33961 & ~n33967 ;
  assign n33970 = ~n33944 & n33969 ;
  assign n33971 = ~n33968 & ~n33970 ;
  assign n33972 = n6861 & n33909 ;
  assign n33973 = n33922 & n33972 ;
  assign n33974 = ~\pi0180  & \pi0625  ;
  assign n33975 = ~n22727 & ~n33974 ;
  assign n33976 = ~n33973 & ~n33975 ;
  assign n33977 = ~\pi1153  & ~n33976 ;
  assign n33978 = n33971 & n33977 ;
  assign n33979 = ~\pi0074  & ~\pi0702  ;
  assign n33980 = ~\pi0100  & n33979 ;
  assign n33981 = n1287 & n33980 ;
  assign n33982 = ~\pi0180  & ~n33981 ;
  assign n33983 = n21768 & n33982 ;
  assign n33984 = n21770 & n33982 ;
  assign n33985 = ~n21734 & n33984 ;
  assign n33986 = ~n33983 & ~n33985 ;
  assign n33987 = \pi0625  & ~n33986 ;
  assign n33988 = ~\pi0180  & ~n22017 ;
  assign n33989 = ~n21994 & n33988 ;
  assign n33990 = ~\pi0038  & ~\pi0180  ;
  assign n33991 = n6861 & ~n33990 ;
  assign n33992 = ~n22109 & n33991 ;
  assign n33993 = ~n33989 & ~n33992 ;
  assign n33994 = ~\pi0180  & ~n21757 ;
  assign n33995 = n22117 & ~n33994 ;
  assign n33996 = ~\pi0702  & ~n33995 ;
  assign n33997 = \pi0625  & n33996 ;
  assign n33998 = ~n33993 & n33997 ;
  assign n33999 = ~n33987 & ~n33998 ;
  assign n34000 = n21768 & n33966 ;
  assign n34001 = n21770 & n33966 ;
  assign n34002 = ~n21734 & n34001 ;
  assign n34003 = ~n34000 & ~n34002 ;
  assign n34004 = \pi1153  & n34003 ;
  assign n34005 = n33999 & n34004 ;
  assign n34006 = ~\pi0608  & ~n34005 ;
  assign n34007 = ~n33978 & n34006 ;
  assign n34008 = n33924 & ~n33975 ;
  assign n34009 = ~n33961 & ~n33975 ;
  assign n34010 = ~n33944 & n34009 ;
  assign n34011 = ~n34008 & ~n34010 ;
  assign n34012 = ~n33967 & ~n33973 ;
  assign n34013 = \pi1153  & ~n34012 ;
  assign n34014 = n34011 & n34013 ;
  assign n34015 = ~\pi0625  & ~n33986 ;
  assign n34016 = ~\pi0625  & n33996 ;
  assign n34017 = ~n33993 & n34016 ;
  assign n34018 = ~n34015 & ~n34017 ;
  assign n34019 = n21768 & n33974 ;
  assign n34020 = n21770 & n33974 ;
  assign n34021 = ~n21734 & n34020 ;
  assign n34022 = ~n34019 & ~n34021 ;
  assign n34023 = ~\pi1153  & n34022 ;
  assign n34024 = n34018 & n34023 ;
  assign n34025 = \pi0608  & ~n34024 ;
  assign n34026 = ~n34014 & n34025 ;
  assign n34027 = ~n34007 & ~n34026 ;
  assign n34028 = n23638 & ~n34027 ;
  assign n34029 = ~n33965 & ~n34028 ;
  assign n34030 = ~\pi0180  & n21768 ;
  assign n34031 = ~\pi0180  & n21770 ;
  assign n34032 = ~n21734 & n34031 ;
  assign n34033 = ~n34030 & ~n34032 ;
  assign n34034 = ~n32759 & n34033 ;
  assign n34035 = ~\pi0660  & ~n21774 ;
  assign n34036 = n26645 & n33909 ;
  assign n34037 = n33922 & n34036 ;
  assign n34038 = \pi0180  & ~n6861 ;
  assign n34039 = ~n20985 & n34038 ;
  assign n34040 = ~\pi0660  & ~n34039 ;
  assign n34041 = ~n34037 & n34040 ;
  assign n34042 = ~n34035 & ~n34041 ;
  assign n34043 = ~n34034 & ~n34042 ;
  assign n34044 = ~n33993 & n33996 ;
  assign n34045 = ~\pi0778  & n33986 ;
  assign n34046 = ~n34044 & n34045 ;
  assign n34047 = ~\pi0609  & ~n34046 ;
  assign n34048 = \pi1155  & ~n34047 ;
  assign n34049 = ~n34005 & ~n34024 ;
  assign n34050 = n22722 & ~n34049 ;
  assign n34051 = ~n34048 & ~n34050 ;
  assign n34052 = ~n34043 & ~n34051 ;
  assign n34053 = n34029 & n34052 ;
  assign n34054 = \pi0778  & ~n34027 ;
  assign n34055 = ~n34037 & ~n34039 ;
  assign n34056 = n20999 & ~n34055 ;
  assign n34057 = ~n32768 & n34033 ;
  assign n34058 = ~n22787 & ~n34057 ;
  assign n34059 = ~n34056 & n34058 ;
  assign n34060 = \pi0785  & n34059 ;
  assign n34061 = \pi0778  & ~n34049 ;
  assign n34062 = \pi0609  & ~n34046 ;
  assign n34063 = \pi0785  & n34062 ;
  assign n34064 = ~n34061 & n34063 ;
  assign n34065 = ~n34060 & ~n34064 ;
  assign n34066 = n33964 & n34065 ;
  assign n34067 = ~n34054 & n34066 ;
  assign n34068 = \pi0660  & ~n34057 ;
  assign n34069 = ~n34056 & n34068 ;
  assign n34070 = ~n34043 & ~n34069 ;
  assign n34071 = \pi0609  & ~n34058 ;
  assign n34072 = n34046 & n34071 ;
  assign n34073 = \pi0778  & n34071 ;
  assign n34074 = ~n34049 & n34073 ;
  assign n34075 = ~n34072 & ~n34074 ;
  assign n34076 = ~n34070 & n34075 ;
  assign n34077 = ~n34067 & n34076 ;
  assign n34078 = ~n34053 & n34077 ;
  assign n34079 = ~\pi0785  & ~n34067 ;
  assign n34080 = n26700 & ~n34079 ;
  assign n34081 = ~n34078 & n34080 ;
  assign n34082 = n23456 & n33909 ;
  assign n34083 = n33922 & n34082 ;
  assign n34084 = ~n21777 & n34033 ;
  assign n34085 = n21777 & n34038 ;
  assign n34086 = n20811 & ~n34085 ;
  assign n34087 = ~n34084 & n34086 ;
  assign n34088 = ~n34083 & n34087 ;
  assign n34089 = ~\pi0180  & ~n20811 ;
  assign n34090 = n21768 & n34089 ;
  assign n34091 = n21770 & n34089 ;
  assign n34092 = ~n21734 & n34091 ;
  assign n34093 = ~n34090 & ~n34092 ;
  assign n34094 = n22155 & n34093 ;
  assign n34095 = ~n34088 & n34094 ;
  assign n34096 = ~n21034 & n34095 ;
  assign n34097 = ~n22147 & ~n34046 ;
  assign n34098 = ~n34061 & n34097 ;
  assign n34099 = n22147 & ~n34033 ;
  assign n34100 = n24348 & ~n34099 ;
  assign n34101 = ~n21034 & n34100 ;
  assign n34102 = ~n34098 & n34101 ;
  assign n34103 = ~n34096 & ~n34102 ;
  assign n34104 = ~n34088 & n34093 ;
  assign n34105 = n23424 & ~n34104 ;
  assign n34106 = ~\pi0781  & ~n34085 ;
  assign n34107 = ~n34084 & n34106 ;
  assign n34108 = ~n34083 & n34107 ;
  assign n34109 = ~n23423 & n34108 ;
  assign n34110 = n23423 & ~n34033 ;
  assign n34111 = ~n34109 & ~n34110 ;
  assign n34112 = ~n34105 & n34111 ;
  assign n34113 = ~n23880 & ~n34112 ;
  assign n34114 = n23880 & ~n34033 ;
  assign n34115 = n24691 & ~n34114 ;
  assign n34116 = ~n34113 & n34115 ;
  assign n34117 = n26065 & ~n34049 ;
  assign n34118 = n26739 & n33986 ;
  assign n34119 = ~n34044 & n34118 ;
  assign n34120 = ~n23885 & n34033 ;
  assign n34121 = \pi0628  & ~n34120 ;
  assign n34122 = ~n34119 & n34121 ;
  assign n34123 = ~n34117 & n34122 ;
  assign n34124 = ~\pi0180  & ~\pi0628  ;
  assign n34125 = n21768 & n34124 ;
  assign n34126 = n21770 & n34124 ;
  assign n34127 = ~n21734 & n34126 ;
  assign n34128 = ~n34125 & ~n34127 ;
  assign n34129 = \pi1156  & n34128 ;
  assign n34130 = ~\pi0629  & n34129 ;
  assign n34131 = ~n34123 & n34130 ;
  assign n34132 = ~\pi0628  & ~n34120 ;
  assign n34133 = ~n34119 & n34132 ;
  assign n34134 = ~n34117 & n34133 ;
  assign n34135 = ~\pi0180  & \pi0628  ;
  assign n34136 = n21768 & n34135 ;
  assign n34137 = n21770 & n34135 ;
  assign n34138 = ~n21734 & n34137 ;
  assign n34139 = ~n34136 & ~n34138 ;
  assign n34140 = ~\pi1156  & n34139 ;
  assign n34141 = \pi0629  & n34140 ;
  assign n34142 = ~n34134 & n34141 ;
  assign n34143 = ~n34131 & ~n34142 ;
  assign n34144 = ~n34116 & n34143 ;
  assign n34145 = \pi0792  & ~n34144 ;
  assign n34146 = n23380 & ~n34046 ;
  assign n34147 = ~\pi0180  & ~n23380 ;
  assign n34148 = n21768 & n34147 ;
  assign n34149 = n21770 & n34147 ;
  assign n34150 = ~n21734 & n34149 ;
  assign n34151 = ~n34148 & ~n34150 ;
  assign n34152 = n21050 & n34151 ;
  assign n34153 = ~n34146 & n34152 ;
  assign n34154 = \pi0778  & n34152 ;
  assign n34155 = ~n34049 & n34154 ;
  assign n34156 = ~n34153 & ~n34155 ;
  assign n34157 = n23683 & ~n34104 ;
  assign n34158 = n21032 & n34108 ;
  assign n34159 = ~n21032 & ~n34033 ;
  assign n34160 = ~n20876 & ~n34159 ;
  assign n34161 = ~n34158 & n34160 ;
  assign n34162 = ~n34157 & n34161 ;
  assign n34163 = n34156 & ~n34162 ;
  assign n34164 = \pi0789  & ~n34163 ;
  assign n34165 = ~n21038 & ~n34164 ;
  assign n34166 = ~n34145 & n34165 ;
  assign n34167 = n34103 & n34166 ;
  assign n34168 = ~n34081 & n34167 ;
  assign n34169 = ~n22160 & n34151 ;
  assign n34170 = ~n34146 & n34169 ;
  assign n34171 = \pi0778  & n34169 ;
  assign n34172 = ~n34049 & n34171 ;
  assign n34173 = ~n34170 & ~n34172 ;
  assign n34174 = n22160 & n34033 ;
  assign n34175 = n20951 & ~n34174 ;
  assign n34176 = n34173 & n34175 ;
  assign n34177 = ~\pi0626  & ~n34110 ;
  assign n34178 = ~n34109 & n34177 ;
  assign n34179 = ~n34105 & n34178 ;
  assign n34180 = \pi0626  & n34033 ;
  assign n34181 = n20882 & ~n34180 ;
  assign n34182 = ~n34179 & n34181 ;
  assign n34183 = ~n34176 & ~n34182 ;
  assign n34184 = \pi0626  & ~n34110 ;
  assign n34185 = ~n34109 & n34184 ;
  assign n34186 = ~n34105 & n34185 ;
  assign n34187 = ~\pi0626  & n34033 ;
  assign n34188 = n20881 & ~n34187 ;
  assign n34189 = ~n34186 & n34188 ;
  assign n34190 = ~n23856 & ~n34189 ;
  assign n34191 = n34183 & n34190 ;
  assign n34192 = ~n26803 & ~n34191 ;
  assign n34193 = ~n34145 & n34192 ;
  assign n34194 = ~n21067 & ~n34193 ;
  assign n34195 = ~n34168 & n34194 ;
  assign n34196 = ~\pi0180  & \pi0644  ;
  assign n34197 = n21768 & n34196 ;
  assign n34198 = n21770 & n34196 ;
  assign n34199 = ~n21734 & n34198 ;
  assign n34200 = ~n34197 & ~n34199 ;
  assign n34201 = \pi0715  & n34200 ;
  assign n34202 = ~\pi0180  & ~n31367 ;
  assign n34203 = n21768 & n34202 ;
  assign n34204 = n21770 & n34202 ;
  assign n34205 = ~n21734 & n34204 ;
  assign n34206 = ~n34203 & ~n34205 ;
  assign n34207 = ~\pi0644  & ~n34206 ;
  assign n34208 = ~\pi0644  & n31367 ;
  assign n34209 = ~n34112 & n34208 ;
  assign n34210 = ~n34207 & ~n34209 ;
  assign n34211 = n34201 & n34210 ;
  assign n34212 = n31378 & ~n34211 ;
  assign n34213 = ~\pi0715  & n34206 ;
  assign n34214 = ~n23958 & ~n34213 ;
  assign n34215 = n31382 & ~n34112 ;
  assign n34216 = ~n34214 & ~n34215 ;
  assign n34217 = n26824 & ~n34216 ;
  assign n34218 = \pi0790  & ~n34217 ;
  assign n34219 = ~n34212 & n34218 ;
  assign n34220 = ~n34119 & ~n34120 ;
  assign n34221 = ~n34117 & n34220 ;
  assign n34222 = ~\pi0792  & ~n34221 ;
  assign n34223 = ~\pi0647  & ~n34222 ;
  assign n34224 = n21768 & n33773 ;
  assign n34225 = n21770 & n33773 ;
  assign n34226 = ~n21734 & n34225 ;
  assign n34227 = ~n34224 & ~n34226 ;
  assign n34228 = ~\pi1157  & n34227 ;
  assign n34229 = ~n34223 & n34228 ;
  assign n34230 = ~n34123 & n34129 ;
  assign n34231 = ~n34134 & n34140 ;
  assign n34232 = ~n34230 & ~n34231 ;
  assign n34233 = \pi0792  & n34228 ;
  assign n34234 = ~n34232 & n34233 ;
  assign n34235 = ~n34229 & ~n34234 ;
  assign n34236 = ~n20846 & n34114 ;
  assign n34237 = n30376 & ~n34112 ;
  assign n34238 = ~n34236 & ~n34237 ;
  assign n34239 = n20846 & ~n34033 ;
  assign n34240 = ~n20910 & ~n34239 ;
  assign n34241 = n34238 & n34240 ;
  assign n34242 = \pi0630  & ~n34241 ;
  assign n34243 = n34235 & n34242 ;
  assign n34244 = \pi0647  & ~n34222 ;
  assign n34245 = n21768 & n33768 ;
  assign n34246 = n21770 & n33768 ;
  assign n34247 = ~n21734 & n34246 ;
  assign n34248 = ~n34245 & ~n34247 ;
  assign n34249 = \pi1157  & n34248 ;
  assign n34250 = ~n34244 & n34249 ;
  assign n34251 = \pi0792  & n34249 ;
  assign n34252 = ~n34232 & n34251 ;
  assign n34253 = ~n34250 & ~n34252 ;
  assign n34254 = ~\pi0630  & ~n34241 ;
  assign n34255 = n34253 & n34254 ;
  assign n34256 = ~n34243 & ~n34255 ;
  assign n34257 = \pi0787  & n34256 ;
  assign n34258 = ~n34219 & ~n34257 ;
  assign n34259 = ~n34195 & n34258 ;
  assign n34260 = ~\pi0787  & n34222 ;
  assign n34261 = n33084 & ~n34232 ;
  assign n34262 = ~n34260 & ~n34261 ;
  assign n34263 = ~\pi0644  & n34262 ;
  assign n34264 = \pi0715  & ~n34263 ;
  assign n34265 = n34235 & n34253 ;
  assign n34266 = n26918 & ~n34265 ;
  assign n34267 = ~n34264 & ~n34266 ;
  assign n34268 = ~\pi0180  & ~\pi0644  ;
  assign n34269 = n21768 & n34268 ;
  assign n34270 = n21770 & n34268 ;
  assign n34271 = ~n21734 & n34270 ;
  assign n34272 = ~n34269 & ~n34271 ;
  assign n34273 = n34216 & n34272 ;
  assign n34274 = \pi1160  & ~n34273 ;
  assign n34275 = n34267 & n34274 ;
  assign n34276 = \pi0644  & n34262 ;
  assign n34277 = ~\pi0715  & ~n34276 ;
  assign n34278 = n33098 & ~n34265 ;
  assign n34279 = ~n34277 & ~n34278 ;
  assign n34280 = ~\pi1160  & ~n34211 ;
  assign n34281 = n34279 & n34280 ;
  assign n34282 = ~n34275 & ~n34281 ;
  assign n34283 = \pi0790  & ~n34282 ;
  assign n34284 = ~n33900 & ~n34283 ;
  assign n34285 = ~n34259 & n34284 ;
  assign n34286 = ~n33902 & ~n34285 ;
  assign n34287 = ~\pi0181  & \pi0788  ;
  assign n34288 = ~n1689 & n34287 ;
  assign n34289 = ~n20778 & n34288 ;
  assign n34290 = n20886 & n34289 ;
  assign n34291 = ~\pi0754  & n1689 ;
  assign n34292 = n20784 & n34291 ;
  assign n34293 = n22767 & n34292 ;
  assign n34294 = ~\pi0181  & ~n1689 ;
  assign n34295 = ~n34292 & ~n34294 ;
  assign n34296 = ~n20792 & ~n34295 ;
  assign n34297 = ~n34293 & n34296 ;
  assign n34298 = n20801 & ~n34297 ;
  assign n34299 = ~\pi1155  & ~n34294 ;
  assign n34300 = \pi0785  & n34299 ;
  assign n34301 = ~n34293 & n34300 ;
  assign n34302 = ~\pi0785  & ~n34294 ;
  assign n34303 = ~n34292 & n34302 ;
  assign n34304 = ~n20804 & ~n34303 ;
  assign n34305 = n29682 & n34304 ;
  assign n34306 = ~n34301 & n34305 ;
  assign n34307 = ~n34298 & n34306 ;
  assign n34308 = n30847 & n34307 ;
  assign n34309 = ~n34290 & ~n34308 ;
  assign n34310 = ~\pi0709  & n1689 ;
  assign n34311 = n20855 & n34310 ;
  assign n34312 = ~n34294 & ~n34311 ;
  assign n34313 = ~\pi0778  & ~n34312 ;
  assign n34314 = ~\pi0625  & ~\pi0709  ;
  assign n34315 = n1689 & n34314 ;
  assign n34316 = n20855 & n34315 ;
  assign n34317 = \pi1153  & n34316 ;
  assign n34318 = \pi1153  & ~n34294 ;
  assign n34319 = ~n34311 & n34318 ;
  assign n34320 = ~n34317 & ~n34319 ;
  assign n34321 = ~\pi1153  & ~n34294 ;
  assign n34322 = ~n34316 & n34321 ;
  assign n34323 = \pi0778  & ~n34322 ;
  assign n34324 = n34320 & n34323 ;
  assign n34325 = ~n34313 & ~n34324 ;
  assign n34326 = n26474 & ~n34325 ;
  assign n34327 = \pi0629  & ~n34326 ;
  assign n34328 = n34309 & n34327 ;
  assign n34329 = n20887 & n34289 ;
  assign n34330 = n32579 & n34307 ;
  assign n34331 = ~n34329 & ~n34330 ;
  assign n34332 = n26485 & ~n34325 ;
  assign n34333 = ~\pi0629  & ~n34332 ;
  assign n34334 = n34331 & n34333 ;
  assign n34335 = ~n34328 & ~n34334 ;
  assign n34336 = \pi0792  & n34335 ;
  assign n34337 = ~n21067 & ~n34336 ;
  assign n34338 = n26325 & ~n34325 ;
  assign n34339 = ~\pi0181  & ~\pi0647  ;
  assign n34340 = ~n1689 & n34339 ;
  assign n34341 = n20849 & ~n34340 ;
  assign n34342 = ~n34338 & n34341 ;
  assign n34343 = n26319 & ~n34325 ;
  assign n34344 = ~\pi0181  & \pi0647  ;
  assign n34345 = ~n1689 & n34344 ;
  assign n34346 = n20897 & ~n34345 ;
  assign n34347 = ~n34343 & n34346 ;
  assign n34348 = ~n34342 & ~n34347 ;
  assign n34349 = \pi0787  & ~n34348 ;
  assign n34350 = ~n20846 & n34289 ;
  assign n34351 = n30376 & n34307 ;
  assign n34352 = ~n34350 & ~n34351 ;
  assign n34353 = ~\pi0181  & \pi0792  ;
  assign n34354 = ~n1689 & n34353 ;
  assign n34355 = ~n20845 & n34354 ;
  assign n34356 = n32606 & ~n34355 ;
  assign n34357 = n34352 & n34356 ;
  assign n34358 = ~n34349 & ~n34357 ;
  assign n34359 = ~n24761 & n34358 ;
  assign n34360 = ~n34337 & n34359 ;
  assign n34361 = \pi0608  & ~n34322 ;
  assign n34362 = ~n34292 & n34318 ;
  assign n34363 = \pi0778  & ~n34362 ;
  assign n34364 = n26421 & ~n34312 ;
  assign n34365 = ~n34363 & ~n34364 ;
  assign n34366 = n34361 & ~n34365 ;
  assign n34367 = n26147 & ~n34312 ;
  assign n34368 = ~\pi0709  & ~n20784 ;
  assign n34369 = n22113 & n34368 ;
  assign n34370 = n34295 & ~n34369 ;
  assign n34371 = ~n34367 & ~n34370 ;
  assign n34372 = n34321 & ~n34371 ;
  assign n34373 = n26415 & n34320 ;
  assign n34374 = ~n34372 & n34373 ;
  assign n34375 = ~n34366 & ~n34374 ;
  assign n34376 = ~\pi1155  & ~n34313 ;
  assign n34377 = ~n34324 & n34376 ;
  assign n34378 = ~n20999 & ~n34377 ;
  assign n34379 = ~\pi0778  & ~n34370 ;
  assign n34380 = ~n34378 & ~n34379 ;
  assign n34381 = n34375 & n34380 ;
  assign n34382 = n29766 & ~n34313 ;
  assign n34383 = ~n34324 & n34382 ;
  assign n34384 = \pi1155  & ~n34297 ;
  assign n34385 = ~\pi0660  & ~n34384 ;
  assign n34386 = ~n34383 & n34385 ;
  assign n34387 = ~n34381 & n34386 ;
  assign n34388 = \pi0785  & ~n34387 ;
  assign n34389 = n29775 & n34304 ;
  assign n34390 = ~n34301 & n34389 ;
  assign n34391 = ~n34298 & n34390 ;
  assign n34392 = n29779 & ~n34325 ;
  assign n34393 = ~n34391 & ~n34392 ;
  assign n34394 = \pi0781  & ~n34393 ;
  assign n34395 = \pi1155  & ~n34313 ;
  assign n34396 = ~n34324 & n34395 ;
  assign n34397 = ~n21774 & ~n34396 ;
  assign n34398 = ~n34379 & ~n34397 ;
  assign n34399 = n34375 & n34398 ;
  assign n34400 = n26121 & ~n34313 ;
  assign n34401 = ~n34324 & n34400 ;
  assign n34402 = \pi0660  & ~n34299 ;
  assign n34403 = \pi0660  & n34292 ;
  assign n34404 = n22767 & n34403 ;
  assign n34405 = ~n34402 & ~n34404 ;
  assign n34406 = ~n34401 & ~n34405 ;
  assign n34407 = ~n34399 & n34406 ;
  assign n34408 = ~n34394 & ~n34407 ;
  assign n34409 = n34388 & n34408 ;
  assign n34410 = ~\pi0785  & ~n34379 ;
  assign n34411 = ~n34366 & n34410 ;
  assign n34412 = ~n34374 & n34411 ;
  assign n34413 = n21022 & ~n34412 ;
  assign n34414 = ~n34394 & ~n34413 ;
  assign n34415 = n29803 & ~n34414 ;
  assign n34416 = ~n34409 & n34415 ;
  assign n34417 = n29808 & n34304 ;
  assign n34418 = ~n34301 & n34417 ;
  assign n34419 = ~n34298 & n34418 ;
  assign n34420 = n30966 & ~n34325 ;
  assign n34421 = ~n34419 & ~n34420 ;
  assign n34422 = n29818 & ~n34421 ;
  assign n34423 = \pi0626  & ~n34307 ;
  assign n34424 = ~\pi0626  & ~n34294 ;
  assign n34425 = n20881 & ~n34424 ;
  assign n34426 = ~n34423 & n34425 ;
  assign n34427 = n26458 & ~n34325 ;
  assign n34428 = ~\pi0626  & ~n34307 ;
  assign n34429 = \pi0626  & ~n34294 ;
  assign n34430 = n20882 & ~n34429 ;
  assign n34431 = ~n34428 & n34430 ;
  assign n34432 = ~n34427 & ~n34431 ;
  assign n34433 = ~n34426 & n34432 ;
  assign n34434 = \pi0788  & ~n34433 ;
  assign n34435 = ~n34422 & ~n34434 ;
  assign n34436 = ~n34416 & n34435 ;
  assign n34437 = ~n23856 & n34359 ;
  assign n34438 = ~n34436 & n34437 ;
  assign n34439 = ~n34360 & ~n34438 ;
  assign n34440 = n30987 & ~n34352 ;
  assign n34441 = n23312 & n34440 ;
  assign n34442 = \pi1157  & ~n34340 ;
  assign n34443 = ~n34338 & n34442 ;
  assign n34444 = ~\pi1157  & ~n34345 ;
  assign n34445 = ~n34343 & n34444 ;
  assign n34446 = ~n34443 & ~n34445 ;
  assign n34447 = \pi0787  & ~n34446 ;
  assign n34448 = n26333 & ~n34325 ;
  assign n34449 = ~\pi0787  & ~n34448 ;
  assign n34450 = ~\pi1160  & ~n34449 ;
  assign n34451 = n23312 & n34450 ;
  assign n34452 = ~n34447 & n34451 ;
  assign n34453 = ~n34441 & ~n34452 ;
  assign n34454 = \pi0790  & ~n34453 ;
  assign n34455 = \pi1160  & ~n34449 ;
  assign n34456 = ~n34447 & n34455 ;
  assign n34457 = ~n23414 & n34294 ;
  assign n34458 = ~n24886 & n34457 ;
  assign n34459 = n31010 & ~n34352 ;
  assign n34460 = ~n34458 & ~n34459 ;
  assign n34461 = ~n34456 & n34460 ;
  assign n34462 = ~n23313 & ~n34457 ;
  assign n34463 = ~n31019 & ~n34462 ;
  assign n34464 = \pi0790  & n34463 ;
  assign n34465 = ~n34461 & n34464 ;
  assign n34466 = ~n34454 & ~n34465 ;
  assign n34467 = \pi0832  & n34466 ;
  assign n34468 = n34439 & n34467 ;
  assign n34469 = \pi0181  & ~\pi0832  ;
  assign n34470 = ~n21132 & ~n34469 ;
  assign n34471 = ~n34468 & n34470 ;
  assign n34472 = ~\pi0074  & ~\pi0709  ;
  assign n34473 = ~\pi0100  & n34472 ;
  assign n34474 = n1287 & n34473 ;
  assign n34475 = ~\pi0181  & ~n34474 ;
  assign n34476 = n21768 & n34475 ;
  assign n34477 = n21770 & n34475 ;
  assign n34478 = ~n21734 & n34477 ;
  assign n34479 = ~n34476 & ~n34478 ;
  assign n34480 = \pi0625  & ~n34479 ;
  assign n34481 = ~\pi0181  & ~n22017 ;
  assign n34482 = ~n21994 & n34481 ;
  assign n34483 = ~\pi0038  & ~\pi0181  ;
  assign n34484 = n6861 & ~n34483 ;
  assign n34485 = ~n22109 & n34484 ;
  assign n34486 = ~n34482 & ~n34485 ;
  assign n34487 = ~\pi0181  & ~n21757 ;
  assign n34488 = n22117 & ~n34487 ;
  assign n34489 = ~\pi0709  & ~n34488 ;
  assign n34490 = \pi0625  & n34489 ;
  assign n34491 = ~n34486 & n34490 ;
  assign n34492 = ~n34480 & ~n34491 ;
  assign n34493 = ~\pi0181  & ~\pi0625  ;
  assign n34494 = n21768 & n34493 ;
  assign n34495 = n21770 & n34493 ;
  assign n34496 = ~n21734 & n34495 ;
  assign n34497 = ~n34494 & ~n34496 ;
  assign n34498 = \pi1153  & n34497 ;
  assign n34499 = n34492 & n34498 ;
  assign n34500 = ~\pi0625  & ~n34479 ;
  assign n34501 = ~\pi0625  & n34489 ;
  assign n34502 = ~n34486 & n34501 ;
  assign n34503 = ~n34500 & ~n34502 ;
  assign n34504 = ~\pi0181  & \pi0625  ;
  assign n34505 = n21768 & n34504 ;
  assign n34506 = n21770 & n34504 ;
  assign n34507 = ~n21734 & n34506 ;
  assign n34508 = ~n34505 & ~n34507 ;
  assign n34509 = ~\pi1153  & n34508 ;
  assign n34510 = n34503 & n34509 ;
  assign n34511 = ~n34499 & ~n34510 ;
  assign n34512 = n26065 & ~n34511 ;
  assign n34513 = ~n34486 & n34489 ;
  assign n34514 = n26739 & n34479 ;
  assign n34515 = ~n34513 & n34514 ;
  assign n34516 = ~\pi0181  & n21768 ;
  assign n34517 = ~\pi0181  & n21770 ;
  assign n34518 = ~n21734 & n34517 ;
  assign n34519 = ~n34516 & ~n34518 ;
  assign n34520 = ~n23885 & n34519 ;
  assign n34521 = ~n34515 & ~n34520 ;
  assign n34522 = ~n34512 & n34521 ;
  assign n34523 = ~\pi0792  & ~n34522 ;
  assign n34524 = ~\pi0787  & n34523 ;
  assign n34525 = \pi0628  & ~n34520 ;
  assign n34526 = ~n34515 & n34525 ;
  assign n34527 = ~n34512 & n34526 ;
  assign n34528 = ~\pi0181  & ~\pi0628  ;
  assign n34529 = n21768 & n34528 ;
  assign n34530 = n21770 & n34528 ;
  assign n34531 = ~n21734 & n34530 ;
  assign n34532 = ~n34529 & ~n34531 ;
  assign n34533 = \pi1156  & n34532 ;
  assign n34534 = ~n34527 & n34533 ;
  assign n34535 = ~\pi0628  & ~n34520 ;
  assign n34536 = ~n34515 & n34535 ;
  assign n34537 = ~n34512 & n34536 ;
  assign n34538 = ~\pi0181  & \pi0628  ;
  assign n34539 = n21768 & n34538 ;
  assign n34540 = n21770 & n34538 ;
  assign n34541 = ~n21734 & n34540 ;
  assign n34542 = ~n34539 & ~n34541 ;
  assign n34543 = ~\pi1156  & n34542 ;
  assign n34544 = ~n34537 & n34543 ;
  assign n34545 = ~n34534 & ~n34544 ;
  assign n34546 = n33084 & ~n34545 ;
  assign n34547 = ~n34524 & ~n34546 ;
  assign n34548 = ~\pi0644  & n34547 ;
  assign n34549 = \pi0715  & ~n34548 ;
  assign n34550 = \pi0647  & ~n34523 ;
  assign n34551 = n21768 & n34339 ;
  assign n34552 = n21770 & n34339 ;
  assign n34553 = ~n21734 & n34552 ;
  assign n34554 = ~n34551 & ~n34553 ;
  assign n34555 = \pi1157  & n34554 ;
  assign n34556 = ~n34550 & n34555 ;
  assign n34557 = \pi0792  & n34555 ;
  assign n34558 = ~n34545 & n34557 ;
  assign n34559 = ~n34556 & ~n34558 ;
  assign n34560 = ~\pi0647  & ~n34523 ;
  assign n34561 = n21768 & n34344 ;
  assign n34562 = n21770 & n34344 ;
  assign n34563 = ~n21734 & n34562 ;
  assign n34564 = ~n34561 & ~n34563 ;
  assign n34565 = ~\pi1157  & n34564 ;
  assign n34566 = ~n34560 & n34565 ;
  assign n34567 = \pi0792  & n34565 ;
  assign n34568 = ~n34545 & n34567 ;
  assign n34569 = ~n34566 & ~n34568 ;
  assign n34570 = n34559 & n34569 ;
  assign n34571 = n26918 & ~n34570 ;
  assign n34572 = ~n34549 & ~n34571 ;
  assign n34573 = ~\pi0181  & ~n31367 ;
  assign n34574 = n21768 & n34573 ;
  assign n34575 = n21770 & n34573 ;
  assign n34576 = ~n21734 & n34575 ;
  assign n34577 = ~n34574 & ~n34576 ;
  assign n34578 = ~\pi0715  & n34577 ;
  assign n34579 = ~n23958 & ~n34578 ;
  assign n34580 = ~\pi0181  & ~n20811 ;
  assign n34581 = n21768 & n34580 ;
  assign n34582 = n21770 & n34580 ;
  assign n34583 = ~n21734 & n34582 ;
  assign n34584 = ~n34581 & ~n34583 ;
  assign n34585 = ~\pi0181  & \pi0754  ;
  assign n34586 = n21743 & n34585 ;
  assign n34587 = ~n21734 & n34586 ;
  assign n34588 = ~\pi0038  & n34587 ;
  assign n34589 = \pi0181  & ~n25023 ;
  assign n34590 = ~\pi0181  & ~n21467 ;
  assign n34591 = ~\pi0754  & ~n34590 ;
  assign n34592 = ~n34589 & n34591 ;
  assign n34593 = ~\pi0039  & ~\pi0181  ;
  assign n34594 = n21272 & n34593 ;
  assign n34595 = ~\pi0038  & ~n34594 ;
  assign n34596 = n34592 & n34595 ;
  assign n34597 = ~n34588 & ~n34596 ;
  assign n34598 = \pi0038  & n34292 ;
  assign n34599 = n8413 & n34598 ;
  assign n34600 = n1354 & n34599 ;
  assign n34601 = n1358 & n34600 ;
  assign n34602 = \pi0038  & ~\pi0181  ;
  assign n34603 = ~n21757 & n34602 ;
  assign n34604 = ~n34601 & ~n34603 ;
  assign n34605 = n23456 & n34604 ;
  assign n34606 = n34597 & n34605 ;
  assign n34607 = ~n21777 & n34519 ;
  assign n34608 = \pi0181  & ~n6861 ;
  assign n34609 = n21777 & n34608 ;
  assign n34610 = n20811 & ~n34609 ;
  assign n34611 = ~n34607 & n34610 ;
  assign n34612 = ~n34606 & n34611 ;
  assign n34613 = n34584 & ~n34612 ;
  assign n34614 = n23424 & ~n34613 ;
  assign n34615 = ~\pi0781  & ~n34609 ;
  assign n34616 = ~n34607 & n34615 ;
  assign n34617 = ~n34606 & n34616 ;
  assign n34618 = ~n23423 & n34617 ;
  assign n34619 = n23423 & ~n34519 ;
  assign n34620 = ~n34618 & ~n34619 ;
  assign n34621 = ~n34614 & n34620 ;
  assign n34622 = n31382 & ~n34621 ;
  assign n34623 = ~n34579 & ~n34622 ;
  assign n34624 = ~\pi0181  & ~\pi0644  ;
  assign n34625 = n21768 & n34624 ;
  assign n34626 = n21770 & n34624 ;
  assign n34627 = ~n21734 & n34626 ;
  assign n34628 = ~n34625 & ~n34627 ;
  assign n34629 = n34623 & n34628 ;
  assign n34630 = \pi1160  & ~n34629 ;
  assign n34631 = n34572 & n34630 ;
  assign n34632 = \pi0644  & n34547 ;
  assign n34633 = ~\pi0715  & ~n34632 ;
  assign n34634 = n33098 & ~n34570 ;
  assign n34635 = ~n34633 & ~n34634 ;
  assign n34636 = ~\pi0181  & \pi0644  ;
  assign n34637 = n21768 & n34636 ;
  assign n34638 = n21770 & n34636 ;
  assign n34639 = ~n21734 & n34638 ;
  assign n34640 = ~n34637 & ~n34639 ;
  assign n34641 = \pi0715  & n34640 ;
  assign n34642 = ~\pi0644  & ~n34577 ;
  assign n34643 = n34208 & ~n34621 ;
  assign n34644 = ~n34642 & ~n34643 ;
  assign n34645 = n34641 & n34644 ;
  assign n34646 = ~\pi1160  & ~n34645 ;
  assign n34647 = n34635 & n34646 ;
  assign n34648 = ~n34631 & ~n34647 ;
  assign n34649 = \pi0790  & ~n34648 ;
  assign n34650 = n9948 & ~n34468 ;
  assign n34651 = n34649 & n34650 ;
  assign n34652 = ~n23880 & ~n34621 ;
  assign n34653 = n23880 & ~n34519 ;
  assign n34654 = n24691 & ~n34653 ;
  assign n34655 = ~n34652 & n34654 ;
  assign n34656 = ~\pi0629  & n34533 ;
  assign n34657 = ~n34527 & n34656 ;
  assign n34658 = \pi0629  & n34543 ;
  assign n34659 = ~n34537 & n34658 ;
  assign n34660 = ~n34657 & ~n34659 ;
  assign n34661 = ~n34655 & n34660 ;
  assign n34662 = \pi0792  & ~n34661 ;
  assign n34663 = ~\pi0778  & n34479 ;
  assign n34664 = ~n34513 & n34663 ;
  assign n34665 = n23380 & ~n34664 ;
  assign n34666 = ~\pi0181  & ~n23380 ;
  assign n34667 = n21768 & n34666 ;
  assign n34668 = n21770 & n34666 ;
  assign n34669 = ~n21734 & n34668 ;
  assign n34670 = ~n34667 & ~n34669 ;
  assign n34671 = ~n22160 & n34670 ;
  assign n34672 = ~n34665 & n34671 ;
  assign n34673 = \pi0778  & n34671 ;
  assign n34674 = ~n34511 & n34673 ;
  assign n34675 = ~n34672 & ~n34674 ;
  assign n34676 = n22160 & n34519 ;
  assign n34677 = n20951 & ~n34676 ;
  assign n34678 = n34675 & n34677 ;
  assign n34679 = ~\pi0626  & ~n34619 ;
  assign n34680 = ~n34618 & n34679 ;
  assign n34681 = ~n34614 & n34680 ;
  assign n34682 = \pi0626  & n34519 ;
  assign n34683 = n20882 & ~n34682 ;
  assign n34684 = ~n34681 & n34683 ;
  assign n34685 = ~n34678 & ~n34684 ;
  assign n34686 = \pi0626  & ~n34619 ;
  assign n34687 = ~n34618 & n34686 ;
  assign n34688 = ~n34614 & n34687 ;
  assign n34689 = ~\pi0626  & n34519 ;
  assign n34690 = n20881 & ~n34689 ;
  assign n34691 = ~n34688 & n34690 ;
  assign n34692 = ~n23856 & ~n34691 ;
  assign n34693 = n34685 & n34692 ;
  assign n34694 = ~n26803 & ~n34693 ;
  assign n34695 = ~n34662 & n34694 ;
  assign n34696 = ~n21067 & ~n34695 ;
  assign n34697 = ~n20846 & n34653 ;
  assign n34698 = n30376 & ~n34621 ;
  assign n34699 = ~n34697 & ~n34698 ;
  assign n34700 = ~n20845 & n21768 ;
  assign n34701 = ~n20845 & n21770 ;
  assign n34702 = ~n21734 & n34701 ;
  assign n34703 = ~n34700 & ~n34702 ;
  assign n34704 = n34353 & ~n34703 ;
  assign n34705 = ~n20910 & ~n34704 ;
  assign n34706 = n34699 & n34705 ;
  assign n34707 = \pi0630  & ~n34706 ;
  assign n34708 = n34569 & n34707 ;
  assign n34709 = ~\pi0630  & ~n34706 ;
  assign n34710 = n34559 & n34709 ;
  assign n34711 = ~n34708 & ~n34710 ;
  assign n34712 = \pi0787  & n34711 ;
  assign n34713 = ~n34696 & ~n34712 ;
  assign n34714 = n34597 & n34604 ;
  assign n34715 = \pi0709  & ~n34714 ;
  assign n34716 = ~\pi0181  & ~\pi0778  ;
  assign n34717 = ~n23622 & ~n34716 ;
  assign n34718 = n34715 & ~n34717 ;
  assign n34719 = ~\pi0181  & n23548 ;
  assign n34720 = ~\pi0754  & ~n34719 ;
  assign n34721 = ~\pi0039  & ~\pi0754  ;
  assign n34722 = ~n22683 & n34721 ;
  assign n34723 = ~n34720 & ~n34722 ;
  assign n34724 = ~\pi0038  & n34723 ;
  assign n34725 = ~\pi0038  & \pi0181  ;
  assign n34726 = ~n26538 & n34725 ;
  assign n34727 = ~n34724 & ~n34726 ;
  assign n34728 = ~\pi0181  & ~n23567 ;
  assign n34729 = n23565 & n34728 ;
  assign n34730 = \pi0754  & n23575 ;
  assign n34731 = n23572 & n34730 ;
  assign n34732 = ~n34585 & ~n34731 ;
  assign n34733 = ~n34729 & ~n34732 ;
  assign n34734 = ~n34727 & ~n34733 ;
  assign n34735 = n6861 & n34734 ;
  assign n34736 = \pi0181  & ~\pi0754  ;
  assign n34737 = n1689 & n34736 ;
  assign n34738 = n20784 & n34737 ;
  assign n34739 = \pi0181  & ~n20784 ;
  assign n34740 = n22113 & n34739 ;
  assign n34741 = ~n34738 & ~n34740 ;
  assign n34742 = n26554 & ~n34741 ;
  assign n34743 = n1358 & n34742 ;
  assign n34744 = \pi0038  & ~n34743 ;
  assign n34745 = ~\pi0709  & ~n34744 ;
  assign n34746 = ~\pi0181  & ~\pi0709  ;
  assign n34747 = ~n26566 & n34746 ;
  assign n34748 = ~\pi0754  & n34746 ;
  assign n34749 = ~n22536 & n34748 ;
  assign n34750 = ~n34747 & ~n34749 ;
  assign n34751 = ~n34745 & n34750 ;
  assign n34752 = n6861 & n34751 ;
  assign n34753 = ~n34717 & ~n34752 ;
  assign n34754 = ~n34735 & n34753 ;
  assign n34755 = ~n34718 & ~n34754 ;
  assign n34756 = \pi0609  & ~n34755 ;
  assign n34757 = ~n22734 & ~n34493 ;
  assign n34758 = n34715 & ~n34757 ;
  assign n34759 = ~n34752 & ~n34757 ;
  assign n34760 = ~n34735 & n34759 ;
  assign n34761 = ~n34758 & ~n34760 ;
  assign n34762 = n6861 & n34604 ;
  assign n34763 = n34597 & n34762 ;
  assign n34764 = ~n22727 & ~n34504 ;
  assign n34765 = ~n34763 & ~n34764 ;
  assign n34766 = ~\pi1153  & ~n34765 ;
  assign n34767 = n34761 & n34766 ;
  assign n34768 = ~\pi0608  & ~n34499 ;
  assign n34769 = ~n34767 & n34768 ;
  assign n34770 = n34715 & ~n34764 ;
  assign n34771 = ~n34752 & ~n34764 ;
  assign n34772 = ~n34735 & n34771 ;
  assign n34773 = ~n34770 & ~n34772 ;
  assign n34774 = ~n34757 & ~n34763 ;
  assign n34775 = \pi1153  & ~n34774 ;
  assign n34776 = n34773 & n34775 ;
  assign n34777 = \pi0608  & ~n34510 ;
  assign n34778 = ~n34776 & n34777 ;
  assign n34779 = ~n34769 & ~n34778 ;
  assign n34780 = n23638 & ~n34779 ;
  assign n34781 = ~n34756 & ~n34780 ;
  assign n34782 = ~n32759 & n34519 ;
  assign n34783 = n26645 & n34604 ;
  assign n34784 = n34597 & n34783 ;
  assign n34785 = ~n20985 & n34608 ;
  assign n34786 = ~\pi0660  & ~n34785 ;
  assign n34787 = ~n34784 & n34786 ;
  assign n34788 = ~n34035 & ~n34787 ;
  assign n34789 = ~n34782 & ~n34788 ;
  assign n34790 = ~\pi0609  & ~n34664 ;
  assign n34791 = \pi1155  & ~n34790 ;
  assign n34792 = n22722 & ~n34511 ;
  assign n34793 = ~n34791 & ~n34792 ;
  assign n34794 = ~n34789 & ~n34793 ;
  assign n34795 = n34781 & n34794 ;
  assign n34796 = \pi0778  & ~n34779 ;
  assign n34797 = ~n34784 & ~n34785 ;
  assign n34798 = n20999 & ~n34797 ;
  assign n34799 = ~n32768 & n34519 ;
  assign n34800 = ~n22787 & ~n34799 ;
  assign n34801 = ~n34798 & n34800 ;
  assign n34802 = \pi0785  & n34801 ;
  assign n34803 = \pi0778  & ~n34511 ;
  assign n34804 = \pi0609  & ~n34664 ;
  assign n34805 = \pi0785  & n34804 ;
  assign n34806 = ~n34803 & n34805 ;
  assign n34807 = ~n34802 & ~n34806 ;
  assign n34808 = n34755 & n34807 ;
  assign n34809 = ~n34796 & n34808 ;
  assign n34810 = \pi0660  & ~n34799 ;
  assign n34811 = ~n34798 & n34810 ;
  assign n34812 = ~n34789 & ~n34811 ;
  assign n34813 = \pi0609  & ~n34800 ;
  assign n34814 = n34664 & n34813 ;
  assign n34815 = \pi0778  & n34813 ;
  assign n34816 = ~n34511 & n34815 ;
  assign n34817 = ~n34814 & ~n34816 ;
  assign n34818 = ~n34812 & n34817 ;
  assign n34819 = ~n34809 & n34818 ;
  assign n34820 = ~n34795 & n34819 ;
  assign n34821 = ~\pi0785  & ~n34809 ;
  assign n34822 = n26700 & ~n34821 ;
  assign n34823 = ~n34820 & n34822 ;
  assign n34824 = n21050 & n34670 ;
  assign n34825 = ~n34665 & n34824 ;
  assign n34826 = \pi0778  & n34824 ;
  assign n34827 = ~n34511 & n34826 ;
  assign n34828 = ~n34825 & ~n34827 ;
  assign n34829 = n23683 & ~n34613 ;
  assign n34830 = n21032 & n34617 ;
  assign n34831 = ~\pi0181  & ~n21032 ;
  assign n34832 = n21768 & n34831 ;
  assign n34833 = n21770 & n34831 ;
  assign n34834 = ~n21734 & n34833 ;
  assign n34835 = ~n34832 & ~n34834 ;
  assign n34836 = ~n20876 & n34835 ;
  assign n34837 = ~n34830 & n34836 ;
  assign n34838 = ~n34829 & n34837 ;
  assign n34839 = n34828 & ~n34838 ;
  assign n34840 = \pi0789  & ~n34839 ;
  assign n34841 = n22155 & n34584 ;
  assign n34842 = ~n34612 & n34841 ;
  assign n34843 = ~n21034 & n34842 ;
  assign n34844 = ~n22147 & ~n34664 ;
  assign n34845 = ~n34803 & n34844 ;
  assign n34846 = n22147 & ~n34519 ;
  assign n34847 = n24348 & ~n34846 ;
  assign n34848 = ~n21034 & n34847 ;
  assign n34849 = ~n34845 & n34848 ;
  assign n34850 = ~n34843 & ~n34849 ;
  assign n34851 = ~n21038 & n34850 ;
  assign n34852 = ~n34840 & n34851 ;
  assign n34853 = ~n34662 & n34852 ;
  assign n34854 = ~n34712 & n34853 ;
  assign n34855 = ~n34823 & n34854 ;
  assign n34856 = ~n34713 & ~n34855 ;
  assign n34857 = n31378 & ~n34645 ;
  assign n34858 = n26824 & ~n34623 ;
  assign n34859 = \pi0790  & ~n34858 ;
  assign n34860 = ~n34857 & n34859 ;
  assign n34861 = n34650 & ~n34860 ;
  assign n34862 = ~n34856 & n34861 ;
  assign n34863 = ~n34651 & ~n34862 ;
  assign n34864 = ~n34471 & n34863 ;
  assign n34865 = ~\pi0182  & \pi0788  ;
  assign n34866 = ~n1689 & n34865 ;
  assign n34867 = ~n20778 & n34866 ;
  assign n34868 = n20886 & n34867 ;
  assign n34869 = ~\pi0756  & n1689 ;
  assign n34870 = n20784 & n34869 ;
  assign n34871 = n22767 & n34870 ;
  assign n34872 = ~\pi0182  & ~n1689 ;
  assign n34873 = ~n34870 & ~n34872 ;
  assign n34874 = ~n20792 & ~n34873 ;
  assign n34875 = ~n34871 & n34874 ;
  assign n34876 = n20801 & ~n34875 ;
  assign n34877 = ~\pi1155  & ~n34872 ;
  assign n34878 = \pi0785  & n34877 ;
  assign n34879 = ~n34871 & n34878 ;
  assign n34880 = ~\pi0785  & ~n34872 ;
  assign n34881 = ~n34870 & n34880 ;
  assign n34882 = ~n20804 & ~n34881 ;
  assign n34883 = n29682 & n34882 ;
  assign n34884 = ~n34879 & n34883 ;
  assign n34885 = ~n34876 & n34884 ;
  assign n34886 = n30847 & n34885 ;
  assign n34887 = ~n34868 & ~n34886 ;
  assign n34888 = ~\pi0734  & n1689 ;
  assign n34889 = n20855 & n34888 ;
  assign n34890 = ~n34872 & ~n34889 ;
  assign n34891 = ~\pi0778  & ~n34890 ;
  assign n34892 = ~\pi0625  & ~\pi0734  ;
  assign n34893 = n1689 & n34892 ;
  assign n34894 = n20855 & n34893 ;
  assign n34895 = \pi1153  & n34894 ;
  assign n34896 = \pi1153  & ~n34872 ;
  assign n34897 = ~n34889 & n34896 ;
  assign n34898 = ~n34895 & ~n34897 ;
  assign n34899 = ~\pi1153  & ~n34872 ;
  assign n34900 = ~n34894 & n34899 ;
  assign n34901 = \pi0778  & ~n34900 ;
  assign n34902 = n34898 & n34901 ;
  assign n34903 = ~n34891 & ~n34902 ;
  assign n34904 = n26474 & ~n34903 ;
  assign n34905 = \pi0629  & ~n34904 ;
  assign n34906 = n34887 & n34905 ;
  assign n34907 = n20887 & n34867 ;
  assign n34908 = n32579 & n34885 ;
  assign n34909 = ~n34907 & ~n34908 ;
  assign n34910 = n26485 & ~n34903 ;
  assign n34911 = ~\pi0629  & ~n34910 ;
  assign n34912 = n34909 & n34911 ;
  assign n34913 = ~n34906 & ~n34912 ;
  assign n34914 = \pi0792  & n34913 ;
  assign n34915 = ~n21067 & ~n34914 ;
  assign n34916 = n26325 & ~n34903 ;
  assign n34917 = ~\pi0182  & ~\pi0647  ;
  assign n34918 = ~n1689 & n34917 ;
  assign n34919 = n20849 & ~n34918 ;
  assign n34920 = ~n34916 & n34919 ;
  assign n34921 = n26319 & ~n34903 ;
  assign n34922 = ~\pi0182  & \pi0647  ;
  assign n34923 = ~n1689 & n34922 ;
  assign n34924 = n20897 & ~n34923 ;
  assign n34925 = ~n34921 & n34924 ;
  assign n34926 = ~n34920 & ~n34925 ;
  assign n34927 = \pi0787  & ~n34926 ;
  assign n34928 = ~n20846 & n34867 ;
  assign n34929 = n30376 & n34885 ;
  assign n34930 = ~n34928 & ~n34929 ;
  assign n34931 = ~\pi0182  & \pi0792  ;
  assign n34932 = ~n1689 & n34931 ;
  assign n34933 = ~n20845 & n34932 ;
  assign n34934 = n32606 & ~n34933 ;
  assign n34935 = n34930 & n34934 ;
  assign n34936 = ~n34927 & ~n34935 ;
  assign n34937 = ~n24761 & n34936 ;
  assign n34938 = ~n34915 & n34937 ;
  assign n34939 = \pi0608  & ~n34900 ;
  assign n34940 = ~n34870 & n34896 ;
  assign n34941 = \pi0778  & ~n34940 ;
  assign n34942 = n26421 & ~n34890 ;
  assign n34943 = ~n34941 & ~n34942 ;
  assign n34944 = n34939 & ~n34943 ;
  assign n34945 = n26147 & ~n34890 ;
  assign n34946 = ~\pi0734  & ~n20784 ;
  assign n34947 = n22113 & n34946 ;
  assign n34948 = n34873 & ~n34947 ;
  assign n34949 = ~n34945 & ~n34948 ;
  assign n34950 = n34899 & ~n34949 ;
  assign n34951 = n26415 & n34898 ;
  assign n34952 = ~n34950 & n34951 ;
  assign n34953 = ~n34944 & ~n34952 ;
  assign n34954 = ~\pi1155  & ~n34891 ;
  assign n34955 = ~n34902 & n34954 ;
  assign n34956 = ~n20999 & ~n34955 ;
  assign n34957 = ~\pi0778  & ~n34948 ;
  assign n34958 = ~n34956 & ~n34957 ;
  assign n34959 = n34953 & n34958 ;
  assign n34960 = n29766 & ~n34891 ;
  assign n34961 = ~n34902 & n34960 ;
  assign n34962 = \pi1155  & ~n34875 ;
  assign n34963 = ~\pi0660  & ~n34962 ;
  assign n34964 = ~n34961 & n34963 ;
  assign n34965 = ~n34959 & n34964 ;
  assign n34966 = \pi0785  & ~n34965 ;
  assign n34967 = n29775 & n34882 ;
  assign n34968 = ~n34879 & n34967 ;
  assign n34969 = ~n34876 & n34968 ;
  assign n34970 = n29779 & ~n34903 ;
  assign n34971 = ~n34969 & ~n34970 ;
  assign n34972 = \pi0781  & ~n34971 ;
  assign n34973 = \pi1155  & ~n34891 ;
  assign n34974 = ~n34902 & n34973 ;
  assign n34975 = ~n21774 & ~n34974 ;
  assign n34976 = ~n34957 & ~n34975 ;
  assign n34977 = n34953 & n34976 ;
  assign n34978 = n26121 & ~n34891 ;
  assign n34979 = ~n34902 & n34978 ;
  assign n34980 = \pi0660  & ~n34877 ;
  assign n34981 = \pi0660  & n34870 ;
  assign n34982 = n22767 & n34981 ;
  assign n34983 = ~n34980 & ~n34982 ;
  assign n34984 = ~n34979 & ~n34983 ;
  assign n34985 = ~n34977 & n34984 ;
  assign n34986 = ~n34972 & ~n34985 ;
  assign n34987 = n34966 & n34986 ;
  assign n34988 = ~\pi0785  & ~n34957 ;
  assign n34989 = ~n34944 & n34988 ;
  assign n34990 = ~n34952 & n34989 ;
  assign n34991 = n21022 & ~n34990 ;
  assign n34992 = ~n34972 & ~n34991 ;
  assign n34993 = n29803 & ~n34992 ;
  assign n34994 = ~n34987 & n34993 ;
  assign n34995 = n29808 & n34882 ;
  assign n34996 = ~n34879 & n34995 ;
  assign n34997 = ~n34876 & n34996 ;
  assign n34998 = n30966 & ~n34903 ;
  assign n34999 = ~n34997 & ~n34998 ;
  assign n35000 = n29818 & ~n34999 ;
  assign n35001 = \pi0626  & ~n34885 ;
  assign n35002 = ~\pi0626  & ~n34872 ;
  assign n35003 = n20881 & ~n35002 ;
  assign n35004 = ~n35001 & n35003 ;
  assign n35005 = n26458 & ~n34903 ;
  assign n35006 = ~\pi0626  & ~n34885 ;
  assign n35007 = \pi0626  & ~n34872 ;
  assign n35008 = n20882 & ~n35007 ;
  assign n35009 = ~n35006 & n35008 ;
  assign n35010 = ~n35005 & ~n35009 ;
  assign n35011 = ~n35004 & n35010 ;
  assign n35012 = \pi0788  & ~n35011 ;
  assign n35013 = ~n35000 & ~n35012 ;
  assign n35014 = ~n34994 & n35013 ;
  assign n35015 = ~n23856 & n34937 ;
  assign n35016 = ~n35014 & n35015 ;
  assign n35017 = ~n34938 & ~n35016 ;
  assign n35018 = n30987 & ~n34930 ;
  assign n35019 = n23312 & n35018 ;
  assign n35020 = \pi1157  & ~n34918 ;
  assign n35021 = ~n34916 & n35020 ;
  assign n35022 = ~\pi1157  & ~n34923 ;
  assign n35023 = ~n34921 & n35022 ;
  assign n35024 = ~n35021 & ~n35023 ;
  assign n35025 = \pi0787  & ~n35024 ;
  assign n35026 = n26333 & ~n34903 ;
  assign n35027 = ~\pi0787  & ~n35026 ;
  assign n35028 = ~\pi1160  & ~n35027 ;
  assign n35029 = n23312 & n35028 ;
  assign n35030 = ~n35025 & n35029 ;
  assign n35031 = ~n35019 & ~n35030 ;
  assign n35032 = \pi0790  & ~n35031 ;
  assign n35033 = \pi1160  & ~n35027 ;
  assign n35034 = ~n35025 & n35033 ;
  assign n35035 = ~n23414 & n34872 ;
  assign n35036 = ~n24886 & n35035 ;
  assign n35037 = n31010 & ~n34930 ;
  assign n35038 = ~n35036 & ~n35037 ;
  assign n35039 = ~n35034 & n35038 ;
  assign n35040 = ~n23313 & ~n35035 ;
  assign n35041 = ~n31019 & ~n35040 ;
  assign n35042 = \pi0790  & n35041 ;
  assign n35043 = ~n35039 & n35042 ;
  assign n35044 = ~n35032 & ~n35043 ;
  assign n35045 = \pi0832  & n35044 ;
  assign n35046 = n35017 & n35045 ;
  assign n35047 = \pi0182  & ~\pi0832  ;
  assign n35048 = ~n21132 & ~n35047 ;
  assign n35049 = ~n35046 & n35048 ;
  assign n35050 = ~\pi0074  & ~\pi0734  ;
  assign n35051 = ~\pi0100  & n35050 ;
  assign n35052 = n1287 & n35051 ;
  assign n35053 = ~\pi0182  & ~n35052 ;
  assign n35054 = n21768 & n35053 ;
  assign n35055 = n21770 & n35053 ;
  assign n35056 = ~n21734 & n35055 ;
  assign n35057 = ~n35054 & ~n35056 ;
  assign n35058 = \pi0625  & ~n35057 ;
  assign n35059 = ~\pi0182  & ~n22017 ;
  assign n35060 = ~n21994 & n35059 ;
  assign n35061 = ~\pi0038  & ~\pi0182  ;
  assign n35062 = n6861 & ~n35061 ;
  assign n35063 = ~n22109 & n35062 ;
  assign n35064 = ~n35060 & ~n35063 ;
  assign n35065 = ~\pi0182  & ~n21757 ;
  assign n35066 = n22117 & ~n35065 ;
  assign n35067 = ~\pi0734  & ~n35066 ;
  assign n35068 = \pi0625  & n35067 ;
  assign n35069 = ~n35064 & n35068 ;
  assign n35070 = ~n35058 & ~n35069 ;
  assign n35071 = ~\pi0182  & ~\pi0625  ;
  assign n35072 = n21768 & n35071 ;
  assign n35073 = n21770 & n35071 ;
  assign n35074 = ~n21734 & n35073 ;
  assign n35075 = ~n35072 & ~n35074 ;
  assign n35076 = \pi1153  & n35075 ;
  assign n35077 = n35070 & n35076 ;
  assign n35078 = ~\pi0625  & ~n35057 ;
  assign n35079 = ~\pi0625  & n35067 ;
  assign n35080 = ~n35064 & n35079 ;
  assign n35081 = ~n35078 & ~n35080 ;
  assign n35082 = ~\pi0182  & \pi0625  ;
  assign n35083 = n21768 & n35082 ;
  assign n35084 = n21770 & n35082 ;
  assign n35085 = ~n21734 & n35084 ;
  assign n35086 = ~n35083 & ~n35085 ;
  assign n35087 = ~\pi1153  & n35086 ;
  assign n35088 = n35081 & n35087 ;
  assign n35089 = ~n35077 & ~n35088 ;
  assign n35090 = n26065 & ~n35089 ;
  assign n35091 = ~n35064 & n35067 ;
  assign n35092 = n26739 & n35057 ;
  assign n35093 = ~n35091 & n35092 ;
  assign n35094 = ~\pi0182  & n21768 ;
  assign n35095 = ~\pi0182  & n21770 ;
  assign n35096 = ~n21734 & n35095 ;
  assign n35097 = ~n35094 & ~n35096 ;
  assign n35098 = ~n23885 & n35097 ;
  assign n35099 = ~n35093 & ~n35098 ;
  assign n35100 = ~n35090 & n35099 ;
  assign n35101 = ~\pi0792  & ~n35100 ;
  assign n35102 = ~\pi0787  & n35101 ;
  assign n35103 = \pi0628  & ~n35098 ;
  assign n35104 = ~n35093 & n35103 ;
  assign n35105 = ~n35090 & n35104 ;
  assign n35106 = ~\pi0182  & ~\pi0628  ;
  assign n35107 = n21768 & n35106 ;
  assign n35108 = n21770 & n35106 ;
  assign n35109 = ~n21734 & n35108 ;
  assign n35110 = ~n35107 & ~n35109 ;
  assign n35111 = \pi1156  & n35110 ;
  assign n35112 = ~n35105 & n35111 ;
  assign n35113 = ~\pi0628  & ~n35098 ;
  assign n35114 = ~n35093 & n35113 ;
  assign n35115 = ~n35090 & n35114 ;
  assign n35116 = ~\pi0182  & \pi0628  ;
  assign n35117 = n21768 & n35116 ;
  assign n35118 = n21770 & n35116 ;
  assign n35119 = ~n21734 & n35118 ;
  assign n35120 = ~n35117 & ~n35119 ;
  assign n35121 = ~\pi1156  & n35120 ;
  assign n35122 = ~n35115 & n35121 ;
  assign n35123 = ~n35112 & ~n35122 ;
  assign n35124 = n33084 & ~n35123 ;
  assign n35125 = ~n35102 & ~n35124 ;
  assign n35126 = ~\pi0644  & n35125 ;
  assign n35127 = \pi0715  & ~n35126 ;
  assign n35128 = \pi0647  & ~n35101 ;
  assign n35129 = n21768 & n34917 ;
  assign n35130 = n21770 & n34917 ;
  assign n35131 = ~n21734 & n35130 ;
  assign n35132 = ~n35129 & ~n35131 ;
  assign n35133 = \pi1157  & n35132 ;
  assign n35134 = ~n35128 & n35133 ;
  assign n35135 = \pi0792  & n35133 ;
  assign n35136 = ~n35123 & n35135 ;
  assign n35137 = ~n35134 & ~n35136 ;
  assign n35138 = ~\pi0647  & ~n35101 ;
  assign n35139 = n21768 & n34922 ;
  assign n35140 = n21770 & n34922 ;
  assign n35141 = ~n21734 & n35140 ;
  assign n35142 = ~n35139 & ~n35141 ;
  assign n35143 = ~\pi1157  & n35142 ;
  assign n35144 = ~n35138 & n35143 ;
  assign n35145 = \pi0792  & n35143 ;
  assign n35146 = ~n35123 & n35145 ;
  assign n35147 = ~n35144 & ~n35146 ;
  assign n35148 = n35137 & n35147 ;
  assign n35149 = n26918 & ~n35148 ;
  assign n35150 = ~n35127 & ~n35149 ;
  assign n35151 = ~\pi0182  & ~n31367 ;
  assign n35152 = n21768 & n35151 ;
  assign n35153 = n21770 & n35151 ;
  assign n35154 = ~n21734 & n35153 ;
  assign n35155 = ~n35152 & ~n35154 ;
  assign n35156 = ~\pi0715  & n35155 ;
  assign n35157 = ~n23958 & ~n35156 ;
  assign n35158 = ~\pi0182  & ~n20811 ;
  assign n35159 = n21768 & n35158 ;
  assign n35160 = n21770 & n35158 ;
  assign n35161 = ~n21734 & n35160 ;
  assign n35162 = ~n35159 & ~n35161 ;
  assign n35163 = ~\pi0182  & \pi0756  ;
  assign n35164 = n21743 & n35163 ;
  assign n35165 = ~n21734 & n35164 ;
  assign n35166 = ~\pi0038  & n35165 ;
  assign n35167 = \pi0182  & ~n25023 ;
  assign n35168 = ~\pi0182  & ~n21467 ;
  assign n35169 = ~\pi0756  & ~n35168 ;
  assign n35170 = ~n35167 & n35169 ;
  assign n35171 = ~\pi0039  & ~\pi0182  ;
  assign n35172 = n21272 & n35171 ;
  assign n35173 = ~\pi0038  & ~n35172 ;
  assign n35174 = n35170 & n35173 ;
  assign n35175 = ~n35166 & ~n35174 ;
  assign n35176 = \pi0038  & n34870 ;
  assign n35177 = n8413 & n35176 ;
  assign n35178 = n1354 & n35177 ;
  assign n35179 = n1358 & n35178 ;
  assign n35180 = \pi0038  & ~\pi0182  ;
  assign n35181 = ~n21757 & n35180 ;
  assign n35182 = ~n35179 & ~n35181 ;
  assign n35183 = n23456 & n35182 ;
  assign n35184 = n35175 & n35183 ;
  assign n35185 = ~n21777 & n35097 ;
  assign n35186 = \pi0182  & ~n6861 ;
  assign n35187 = n21777 & n35186 ;
  assign n35188 = n20811 & ~n35187 ;
  assign n35189 = ~n35185 & n35188 ;
  assign n35190 = ~n35184 & n35189 ;
  assign n35191 = n35162 & ~n35190 ;
  assign n35192 = n23424 & ~n35191 ;
  assign n35193 = ~\pi0781  & ~n35187 ;
  assign n35194 = ~n35185 & n35193 ;
  assign n35195 = ~n35184 & n35194 ;
  assign n35196 = ~n23423 & n35195 ;
  assign n35197 = n23423 & ~n35097 ;
  assign n35198 = ~n35196 & ~n35197 ;
  assign n35199 = ~n35192 & n35198 ;
  assign n35200 = n31382 & ~n35199 ;
  assign n35201 = ~n35157 & ~n35200 ;
  assign n35202 = ~\pi0182  & ~\pi0644  ;
  assign n35203 = n21768 & n35202 ;
  assign n35204 = n21770 & n35202 ;
  assign n35205 = ~n21734 & n35204 ;
  assign n35206 = ~n35203 & ~n35205 ;
  assign n35207 = n35201 & n35206 ;
  assign n35208 = \pi1160  & ~n35207 ;
  assign n35209 = n35150 & n35208 ;
  assign n35210 = \pi0644  & n35125 ;
  assign n35211 = ~\pi0715  & ~n35210 ;
  assign n35212 = n33098 & ~n35148 ;
  assign n35213 = ~n35211 & ~n35212 ;
  assign n35214 = ~\pi0182  & \pi0644  ;
  assign n35215 = n21768 & n35214 ;
  assign n35216 = n21770 & n35214 ;
  assign n35217 = ~n21734 & n35216 ;
  assign n35218 = ~n35215 & ~n35217 ;
  assign n35219 = \pi0715  & n35218 ;
  assign n35220 = ~\pi0644  & ~n35155 ;
  assign n35221 = n34208 & ~n35199 ;
  assign n35222 = ~n35220 & ~n35221 ;
  assign n35223 = n35219 & n35222 ;
  assign n35224 = ~\pi1160  & ~n35223 ;
  assign n35225 = n35213 & n35224 ;
  assign n35226 = ~n35209 & ~n35225 ;
  assign n35227 = \pi0790  & ~n35226 ;
  assign n35228 = n35175 & n35182 ;
  assign n35229 = \pi0734  & ~n35228 ;
  assign n35230 = ~\pi0182  & ~\pi0778  ;
  assign n35231 = ~n23622 & ~n35230 ;
  assign n35232 = n35229 & ~n35231 ;
  assign n35233 = ~\pi0182  & n23548 ;
  assign n35234 = ~\pi0756  & ~n35233 ;
  assign n35235 = ~\pi0039  & ~\pi0756  ;
  assign n35236 = ~n22683 & n35235 ;
  assign n35237 = ~n35234 & ~n35236 ;
  assign n35238 = ~\pi0038  & n35237 ;
  assign n35239 = ~\pi0038  & \pi0182  ;
  assign n35240 = ~n26538 & n35239 ;
  assign n35241 = ~n35238 & ~n35240 ;
  assign n35242 = ~\pi0182  & ~n23567 ;
  assign n35243 = n23565 & n35242 ;
  assign n35244 = n6861 & n35243 ;
  assign n35245 = \pi0756  & n23575 ;
  assign n35246 = n23572 & n35245 ;
  assign n35247 = n6861 & ~n35163 ;
  assign n35248 = ~n35246 & n35247 ;
  assign n35249 = ~n35244 & ~n35248 ;
  assign n35250 = ~n35241 & ~n35249 ;
  assign n35251 = \pi0182  & ~\pi0756  ;
  assign n35252 = n1689 & n35251 ;
  assign n35253 = n20784 & n35252 ;
  assign n35254 = \pi0182  & ~n20784 ;
  assign n35255 = n22113 & n35254 ;
  assign n35256 = ~n35253 & ~n35255 ;
  assign n35257 = n26554 & ~n35256 ;
  assign n35258 = n1358 & n35257 ;
  assign n35259 = \pi0038  & ~n35258 ;
  assign n35260 = ~\pi0734  & ~n35259 ;
  assign n35261 = ~\pi0182  & ~\pi0734  ;
  assign n35262 = ~n26566 & n35261 ;
  assign n35263 = ~\pi0756  & n35261 ;
  assign n35264 = ~n22536 & n35263 ;
  assign n35265 = ~n35262 & ~n35264 ;
  assign n35266 = ~n35260 & n35265 ;
  assign n35267 = n6861 & n35266 ;
  assign n35268 = ~n35231 & ~n35267 ;
  assign n35269 = ~n35250 & n35268 ;
  assign n35270 = ~n35232 & ~n35269 ;
  assign n35271 = \pi0609  & ~n35270 ;
  assign n35272 = ~n22734 & ~n35071 ;
  assign n35273 = n35229 & ~n35272 ;
  assign n35274 = ~n35267 & ~n35272 ;
  assign n35275 = ~n35250 & n35274 ;
  assign n35276 = ~n35273 & ~n35275 ;
  assign n35277 = n6861 & n35182 ;
  assign n35278 = n35175 & n35277 ;
  assign n35279 = ~n22727 & ~n35082 ;
  assign n35280 = ~n35278 & ~n35279 ;
  assign n35281 = ~\pi1153  & ~n35280 ;
  assign n35282 = n35276 & n35281 ;
  assign n35283 = ~\pi0608  & ~n35077 ;
  assign n35284 = ~n35282 & n35283 ;
  assign n35285 = n35229 & ~n35279 ;
  assign n35286 = ~n35267 & ~n35279 ;
  assign n35287 = ~n35250 & n35286 ;
  assign n35288 = ~n35285 & ~n35287 ;
  assign n35289 = ~n35272 & ~n35278 ;
  assign n35290 = \pi1153  & ~n35289 ;
  assign n35291 = n35288 & n35290 ;
  assign n35292 = \pi0608  & ~n35088 ;
  assign n35293 = ~n35291 & n35292 ;
  assign n35294 = ~n35284 & ~n35293 ;
  assign n35295 = n23638 & ~n35294 ;
  assign n35296 = ~n35271 & ~n35295 ;
  assign n35297 = ~n32759 & n35097 ;
  assign n35298 = n26645 & n35182 ;
  assign n35299 = n35175 & n35298 ;
  assign n35300 = ~n20985 & n35186 ;
  assign n35301 = ~\pi0660  & ~n35300 ;
  assign n35302 = ~n35299 & n35301 ;
  assign n35303 = ~n34035 & ~n35302 ;
  assign n35304 = ~n35297 & ~n35303 ;
  assign n35305 = ~\pi0778  & n35057 ;
  assign n35306 = ~n35091 & n35305 ;
  assign n35307 = ~\pi0609  & ~n35306 ;
  assign n35308 = \pi1155  & ~n35307 ;
  assign n35309 = n22722 & ~n35089 ;
  assign n35310 = ~n35308 & ~n35309 ;
  assign n35311 = ~n35304 & ~n35310 ;
  assign n35312 = n35296 & n35311 ;
  assign n35313 = \pi0778  & ~n35294 ;
  assign n35314 = ~n35299 & ~n35300 ;
  assign n35315 = n20999 & ~n35314 ;
  assign n35316 = ~n32768 & n35097 ;
  assign n35317 = ~n22787 & ~n35316 ;
  assign n35318 = ~n35315 & n35317 ;
  assign n35319 = \pi0785  & n35318 ;
  assign n35320 = \pi0778  & ~n35089 ;
  assign n35321 = \pi0609  & ~n35306 ;
  assign n35322 = \pi0785  & n35321 ;
  assign n35323 = ~n35320 & n35322 ;
  assign n35324 = ~n35319 & ~n35323 ;
  assign n35325 = n35270 & n35324 ;
  assign n35326 = ~n35313 & n35325 ;
  assign n35327 = \pi0660  & ~n35316 ;
  assign n35328 = ~n35315 & n35327 ;
  assign n35329 = ~n35304 & ~n35328 ;
  assign n35330 = \pi0609  & ~n35317 ;
  assign n35331 = n35306 & n35330 ;
  assign n35332 = \pi0778  & n35330 ;
  assign n35333 = ~n35089 & n35332 ;
  assign n35334 = ~n35331 & ~n35333 ;
  assign n35335 = ~n35329 & n35334 ;
  assign n35336 = ~n35326 & n35335 ;
  assign n35337 = ~n35312 & n35336 ;
  assign n35338 = ~\pi0785  & ~n35326 ;
  assign n35339 = n26700 & ~n35338 ;
  assign n35340 = ~n35337 & n35339 ;
  assign n35341 = n22155 & n35162 ;
  assign n35342 = ~n35190 & n35341 ;
  assign n35343 = ~n21034 & n35342 ;
  assign n35344 = ~n22147 & ~n35306 ;
  assign n35345 = ~n35320 & n35344 ;
  assign n35346 = n22147 & ~n35097 ;
  assign n35347 = n24348 & ~n35346 ;
  assign n35348 = ~n21034 & n35347 ;
  assign n35349 = ~n35345 & n35348 ;
  assign n35350 = ~n35343 & ~n35349 ;
  assign n35351 = ~n23880 & ~n35199 ;
  assign n35352 = n23880 & ~n35097 ;
  assign n35353 = n24691 & ~n35352 ;
  assign n35354 = ~n35351 & n35353 ;
  assign n35355 = ~\pi0629  & n35111 ;
  assign n35356 = ~n35105 & n35355 ;
  assign n35357 = \pi0629  & n35121 ;
  assign n35358 = ~n35115 & n35357 ;
  assign n35359 = ~n35356 & ~n35358 ;
  assign n35360 = ~n35354 & n35359 ;
  assign n35361 = \pi0792  & ~n35360 ;
  assign n35362 = n23380 & ~n35306 ;
  assign n35363 = ~\pi0182  & ~n23380 ;
  assign n35364 = n21768 & n35363 ;
  assign n35365 = n21770 & n35363 ;
  assign n35366 = ~n21734 & n35365 ;
  assign n35367 = ~n35364 & ~n35366 ;
  assign n35368 = n21050 & n35367 ;
  assign n35369 = ~n35362 & n35368 ;
  assign n35370 = \pi0778  & n35368 ;
  assign n35371 = ~n35089 & n35370 ;
  assign n35372 = ~n35369 & ~n35371 ;
  assign n35373 = n23683 & ~n35191 ;
  assign n35374 = n21032 & n35195 ;
  assign n35375 = ~\pi0182  & ~n21032 ;
  assign n35376 = n21768 & n35375 ;
  assign n35377 = n21770 & n35375 ;
  assign n35378 = ~n21734 & n35377 ;
  assign n35379 = ~n35376 & ~n35378 ;
  assign n35380 = ~n20876 & n35379 ;
  assign n35381 = ~n35374 & n35380 ;
  assign n35382 = ~n35373 & n35381 ;
  assign n35383 = n35372 & ~n35382 ;
  assign n35384 = \pi0789  & ~n35383 ;
  assign n35385 = ~n21038 & ~n35384 ;
  assign n35386 = ~n35361 & n35385 ;
  assign n35387 = n35350 & n35386 ;
  assign n35388 = ~n35340 & n35387 ;
  assign n35389 = ~n22160 & n35367 ;
  assign n35390 = ~n35362 & n35389 ;
  assign n35391 = \pi0778  & n35389 ;
  assign n35392 = ~n35089 & n35391 ;
  assign n35393 = ~n35390 & ~n35392 ;
  assign n35394 = n22160 & n35097 ;
  assign n35395 = n20951 & ~n35394 ;
  assign n35396 = n35393 & n35395 ;
  assign n35397 = ~\pi0626  & ~n35197 ;
  assign n35398 = ~n35196 & n35397 ;
  assign n35399 = ~n35192 & n35398 ;
  assign n35400 = \pi0626  & n35097 ;
  assign n35401 = n20882 & ~n35400 ;
  assign n35402 = ~n35399 & n35401 ;
  assign n35403 = ~n35396 & ~n35402 ;
  assign n35404 = \pi0626  & ~n35197 ;
  assign n35405 = ~n35196 & n35404 ;
  assign n35406 = ~n35192 & n35405 ;
  assign n35407 = ~\pi0626  & n35097 ;
  assign n35408 = n20881 & ~n35407 ;
  assign n35409 = ~n35406 & n35408 ;
  assign n35410 = ~n23856 & ~n35409 ;
  assign n35411 = n35403 & n35410 ;
  assign n35412 = ~n26803 & ~n35411 ;
  assign n35413 = ~n35361 & n35412 ;
  assign n35414 = ~n21067 & ~n35413 ;
  assign n35415 = ~n35388 & n35414 ;
  assign n35416 = n26824 & ~n35201 ;
  assign n35417 = \pi0790  & ~n31378 ;
  assign n35418 = \pi0790  & n35219 ;
  assign n35419 = n35222 & n35418 ;
  assign n35420 = ~n35417 & ~n35419 ;
  assign n35421 = ~n35416 & ~n35420 ;
  assign n35422 = ~\pi0630  & ~n35128 ;
  assign n35423 = ~\pi0630  & \pi0792  ;
  assign n35424 = ~n35123 & n35423 ;
  assign n35425 = ~n35422 & ~n35424 ;
  assign n35426 = n35133 & ~n35425 ;
  assign n35427 = \pi0630  & ~n35147 ;
  assign n35428 = ~n20846 & n35352 ;
  assign n35429 = n30376 & ~n35199 ;
  assign n35430 = ~n35428 & ~n35429 ;
  assign n35431 = ~n34703 & n34931 ;
  assign n35432 = ~n20910 & ~n35431 ;
  assign n35433 = n35430 & n35432 ;
  assign n35434 = ~n35427 & ~n35433 ;
  assign n35435 = ~n35426 & n35434 ;
  assign n35436 = \pi0787  & ~n35435 ;
  assign n35437 = ~n35421 & ~n35436 ;
  assign n35438 = ~n35415 & n35437 ;
  assign n35439 = ~n35227 & ~n35438 ;
  assign n35440 = n9948 & ~n35046 ;
  assign n35441 = ~n35439 & n35440 ;
  assign n35442 = ~n35049 & ~n35441 ;
  assign n35443 = \pi0183  & ~\pi0832  ;
  assign n35444 = ~n21132 & ~n35443 ;
  assign n35445 = ~\pi0183  & \pi0788  ;
  assign n35446 = ~n1689 & n35445 ;
  assign n35447 = ~n20778 & n35446 ;
  assign n35448 = n20886 & n35447 ;
  assign n35449 = ~\pi0755  & n1689 ;
  assign n35450 = n20784 & n35449 ;
  assign n35451 = n22767 & n35450 ;
  assign n35452 = ~\pi0183  & ~n1689 ;
  assign n35453 = ~n35450 & ~n35452 ;
  assign n35454 = ~n20792 & ~n35453 ;
  assign n35455 = ~n35451 & n35454 ;
  assign n35456 = n20801 & ~n35455 ;
  assign n35457 = ~\pi1155  & ~n35452 ;
  assign n35458 = \pi0785  & n35457 ;
  assign n35459 = ~n35451 & n35458 ;
  assign n35460 = ~\pi0785  & ~n35452 ;
  assign n35461 = ~n35450 & n35460 ;
  assign n35462 = ~n20804 & ~n35461 ;
  assign n35463 = n29682 & n35462 ;
  assign n35464 = ~n35459 & n35463 ;
  assign n35465 = ~n35456 & n35464 ;
  assign n35466 = n30847 & n35465 ;
  assign n35467 = ~n35448 & ~n35466 ;
  assign n35468 = ~\pi0725  & n1689 ;
  assign n35469 = n20855 & n35468 ;
  assign n35470 = ~n35452 & ~n35469 ;
  assign n35471 = ~\pi0778  & ~n35470 ;
  assign n35472 = ~\pi0625  & ~\pi0725  ;
  assign n35473 = n1689 & n35472 ;
  assign n35474 = n20855 & n35473 ;
  assign n35475 = \pi1153  & n35474 ;
  assign n35476 = \pi1153  & ~n35452 ;
  assign n35477 = ~n35469 & n35476 ;
  assign n35478 = ~n35475 & ~n35477 ;
  assign n35479 = ~\pi1153  & ~n35452 ;
  assign n35480 = ~n35474 & n35479 ;
  assign n35481 = \pi0778  & ~n35480 ;
  assign n35482 = n35478 & n35481 ;
  assign n35483 = ~n35471 & ~n35482 ;
  assign n35484 = n26474 & ~n35483 ;
  assign n35485 = \pi0629  & ~n35484 ;
  assign n35486 = n35467 & n35485 ;
  assign n35487 = n20887 & n35447 ;
  assign n35488 = n32579 & n35465 ;
  assign n35489 = ~n35487 & ~n35488 ;
  assign n35490 = n26485 & ~n35483 ;
  assign n35491 = ~\pi0629  & ~n35490 ;
  assign n35492 = n35489 & n35491 ;
  assign n35493 = \pi0792  & ~n35492 ;
  assign n35494 = ~n35486 & n35493 ;
  assign n35495 = ~n21067 & ~n35494 ;
  assign n35496 = n26325 & ~n35483 ;
  assign n35497 = ~\pi0183  & ~\pi0647  ;
  assign n35498 = ~n1689 & n35497 ;
  assign n35499 = n20849 & ~n35498 ;
  assign n35500 = ~n35496 & n35499 ;
  assign n35501 = n26319 & ~n35483 ;
  assign n35502 = ~\pi0183  & \pi0647  ;
  assign n35503 = ~n1689 & n35502 ;
  assign n35504 = n20897 & ~n35503 ;
  assign n35505 = ~n35501 & n35504 ;
  assign n35506 = ~n35500 & ~n35505 ;
  assign n35507 = \pi0787  & ~n35506 ;
  assign n35508 = ~n20846 & n35447 ;
  assign n35509 = n30376 & n35465 ;
  assign n35510 = ~n35508 & ~n35509 ;
  assign n35511 = ~\pi0183  & \pi0792  ;
  assign n35512 = ~n1689 & n35511 ;
  assign n35513 = ~n20845 & n35512 ;
  assign n35514 = n32606 & ~n35513 ;
  assign n35515 = n35510 & n35514 ;
  assign n35516 = ~n35507 & ~n35515 ;
  assign n35517 = ~n24761 & n35516 ;
  assign n35518 = ~n35495 & n35517 ;
  assign n35519 = \pi0608  & ~n35480 ;
  assign n35520 = ~n35450 & n35476 ;
  assign n35521 = \pi0778  & ~n35520 ;
  assign n35522 = n26421 & ~n35470 ;
  assign n35523 = ~n35521 & ~n35522 ;
  assign n35524 = n35519 & ~n35523 ;
  assign n35525 = n26147 & ~n35470 ;
  assign n35526 = ~\pi0725  & ~n20784 ;
  assign n35527 = n22113 & n35526 ;
  assign n35528 = n35453 & ~n35527 ;
  assign n35529 = ~n35525 & ~n35528 ;
  assign n35530 = n35479 & ~n35529 ;
  assign n35531 = n26415 & n35478 ;
  assign n35532 = ~n35530 & n35531 ;
  assign n35533 = ~n35524 & ~n35532 ;
  assign n35534 = ~\pi1155  & ~n35471 ;
  assign n35535 = ~n35482 & n35534 ;
  assign n35536 = ~n20999 & ~n35535 ;
  assign n35537 = ~\pi0778  & ~n35528 ;
  assign n35538 = ~n35536 & ~n35537 ;
  assign n35539 = n35533 & n35538 ;
  assign n35540 = n29766 & ~n35471 ;
  assign n35541 = ~n35482 & n35540 ;
  assign n35542 = \pi1155  & ~n35455 ;
  assign n35543 = ~\pi0660  & ~n35542 ;
  assign n35544 = ~n35541 & n35543 ;
  assign n35545 = ~n35539 & n35544 ;
  assign n35546 = \pi0785  & ~n35545 ;
  assign n35547 = n29775 & n35462 ;
  assign n35548 = ~n35459 & n35547 ;
  assign n35549 = ~n35456 & n35548 ;
  assign n35550 = n29779 & ~n35483 ;
  assign n35551 = ~n35549 & ~n35550 ;
  assign n35552 = \pi0781  & ~n35551 ;
  assign n35553 = \pi1155  & ~n35471 ;
  assign n35554 = ~n35482 & n35553 ;
  assign n35555 = ~n21774 & ~n35554 ;
  assign n35556 = ~n35537 & ~n35555 ;
  assign n35557 = n35533 & n35556 ;
  assign n35558 = n26121 & ~n35471 ;
  assign n35559 = ~n35482 & n35558 ;
  assign n35560 = \pi0660  & ~n35457 ;
  assign n35561 = \pi0660  & n35450 ;
  assign n35562 = n22767 & n35561 ;
  assign n35563 = ~n35560 & ~n35562 ;
  assign n35564 = ~n35559 & ~n35563 ;
  assign n35565 = ~n35557 & n35564 ;
  assign n35566 = ~n35552 & ~n35565 ;
  assign n35567 = n35546 & n35566 ;
  assign n35568 = ~\pi0785  & ~n35537 ;
  assign n35569 = ~n35524 & n35568 ;
  assign n35570 = ~n35532 & n35569 ;
  assign n35571 = n21022 & ~n35570 ;
  assign n35572 = ~n35552 & ~n35571 ;
  assign n35573 = n29803 & ~n35572 ;
  assign n35574 = ~n35567 & n35573 ;
  assign n35575 = n29808 & n35462 ;
  assign n35576 = ~n35459 & n35575 ;
  assign n35577 = ~n35456 & n35576 ;
  assign n35578 = n30966 & ~n35483 ;
  assign n35579 = ~n35577 & ~n35578 ;
  assign n35580 = n29818 & ~n35579 ;
  assign n35581 = \pi0626  & ~n35465 ;
  assign n35582 = ~\pi0626  & ~n35452 ;
  assign n35583 = n20881 & ~n35582 ;
  assign n35584 = ~n35581 & n35583 ;
  assign n35585 = n26458 & ~n35483 ;
  assign n35586 = ~\pi0626  & ~n35465 ;
  assign n35587 = \pi0626  & ~n35452 ;
  assign n35588 = n20882 & ~n35587 ;
  assign n35589 = ~n35586 & n35588 ;
  assign n35590 = ~n35585 & ~n35589 ;
  assign n35591 = ~n35584 & n35590 ;
  assign n35592 = \pi0788  & ~n35591 ;
  assign n35593 = ~n35580 & ~n35592 ;
  assign n35594 = ~n35574 & n35593 ;
  assign n35595 = ~n23856 & n35517 ;
  assign n35596 = ~n35594 & n35595 ;
  assign n35597 = ~n35518 & ~n35596 ;
  assign n35598 = n30987 & ~n35510 ;
  assign n35599 = n23312 & n35598 ;
  assign n35600 = \pi1157  & ~n35498 ;
  assign n35601 = ~n35496 & n35600 ;
  assign n35602 = ~\pi1157  & ~n35503 ;
  assign n35603 = ~n35501 & n35602 ;
  assign n35604 = ~n35601 & ~n35603 ;
  assign n35605 = \pi0787  & ~n35604 ;
  assign n35606 = n26333 & ~n35483 ;
  assign n35607 = ~\pi0787  & ~n35606 ;
  assign n35608 = ~\pi1160  & ~n35607 ;
  assign n35609 = n23312 & n35608 ;
  assign n35610 = ~n35605 & n35609 ;
  assign n35611 = ~n35599 & ~n35610 ;
  assign n35612 = ~n23414 & n35452 ;
  assign n35613 = ~n24886 & n35612 ;
  assign n35614 = ~n23313 & ~n35613 ;
  assign n35615 = \pi1160  & ~n35607 ;
  assign n35616 = ~n35605 & n35615 ;
  assign n35617 = n31010 & ~n35510 ;
  assign n35618 = ~n35613 & ~n35617 ;
  assign n35619 = ~n35616 & n35618 ;
  assign n35620 = ~n35614 & ~n35619 ;
  assign n35621 = n35611 & ~n35620 ;
  assign n35622 = \pi0790  & ~n35621 ;
  assign n35623 = \pi0832  & ~n35622 ;
  assign n35624 = n35597 & n35623 ;
  assign n35625 = n35444 & ~n35624 ;
  assign n35626 = ~\pi0074  & ~\pi0725  ;
  assign n35627 = ~\pi0100  & n35626 ;
  assign n35628 = n1287 & n35627 ;
  assign n35629 = ~\pi0183  & ~n35628 ;
  assign n35630 = n21768 & n35629 ;
  assign n35631 = n21770 & n35629 ;
  assign n35632 = ~n21734 & n35631 ;
  assign n35633 = ~n35630 & ~n35632 ;
  assign n35634 = \pi0625  & ~n35633 ;
  assign n35635 = ~\pi0183  & ~n22017 ;
  assign n35636 = ~n21994 & n35635 ;
  assign n35637 = ~\pi0038  & ~\pi0183  ;
  assign n35638 = n6861 & ~n35637 ;
  assign n35639 = ~n22109 & n35638 ;
  assign n35640 = ~n35636 & ~n35639 ;
  assign n35641 = ~\pi0183  & ~n21757 ;
  assign n35642 = n22117 & ~n35641 ;
  assign n35643 = ~\pi0725  & ~n35642 ;
  assign n35644 = \pi0625  & n35643 ;
  assign n35645 = ~n35640 & n35644 ;
  assign n35646 = ~n35634 & ~n35645 ;
  assign n35647 = ~\pi0183  & ~\pi0625  ;
  assign n35648 = n21768 & n35647 ;
  assign n35649 = n21770 & n35647 ;
  assign n35650 = ~n21734 & n35649 ;
  assign n35651 = ~n35648 & ~n35650 ;
  assign n35652 = \pi1153  & n35651 ;
  assign n35653 = n35646 & n35652 ;
  assign n35654 = ~\pi0625  & ~n35633 ;
  assign n35655 = ~\pi0625  & n35643 ;
  assign n35656 = ~n35640 & n35655 ;
  assign n35657 = ~n35654 & ~n35656 ;
  assign n35658 = ~\pi0183  & \pi0625  ;
  assign n35659 = n21768 & n35658 ;
  assign n35660 = n21770 & n35658 ;
  assign n35661 = ~n21734 & n35660 ;
  assign n35662 = ~n35659 & ~n35661 ;
  assign n35663 = ~\pi1153  & n35662 ;
  assign n35664 = n35657 & n35663 ;
  assign n35665 = ~n35653 & ~n35664 ;
  assign n35666 = n26065 & ~n35665 ;
  assign n35667 = ~n35640 & n35643 ;
  assign n35668 = n26739 & n35633 ;
  assign n35669 = ~n35667 & n35668 ;
  assign n35670 = ~\pi0183  & n21768 ;
  assign n35671 = ~\pi0183  & n21770 ;
  assign n35672 = ~n21734 & n35671 ;
  assign n35673 = ~n35670 & ~n35672 ;
  assign n35674 = ~n23885 & n35673 ;
  assign n35675 = ~n35669 & ~n35674 ;
  assign n35676 = ~n35666 & n35675 ;
  assign n35677 = ~\pi0792  & ~n35676 ;
  assign n35678 = ~\pi0787  & n35677 ;
  assign n35679 = \pi0628  & ~n35674 ;
  assign n35680 = ~n35669 & n35679 ;
  assign n35681 = ~n35666 & n35680 ;
  assign n35682 = ~\pi0183  & ~\pi0628  ;
  assign n35683 = n21768 & n35682 ;
  assign n35684 = n21770 & n35682 ;
  assign n35685 = ~n21734 & n35684 ;
  assign n35686 = ~n35683 & ~n35685 ;
  assign n35687 = \pi1156  & n35686 ;
  assign n35688 = ~n35681 & n35687 ;
  assign n35689 = ~\pi0628  & ~n35674 ;
  assign n35690 = ~n35669 & n35689 ;
  assign n35691 = ~n35666 & n35690 ;
  assign n35692 = ~\pi0183  & \pi0628  ;
  assign n35693 = n21768 & n35692 ;
  assign n35694 = n21770 & n35692 ;
  assign n35695 = ~n21734 & n35694 ;
  assign n35696 = ~n35693 & ~n35695 ;
  assign n35697 = ~\pi1156  & n35696 ;
  assign n35698 = ~n35691 & n35697 ;
  assign n35699 = ~n35688 & ~n35698 ;
  assign n35700 = n33084 & ~n35699 ;
  assign n35701 = ~n35678 & ~n35700 ;
  assign n35702 = ~\pi0644  & n35701 ;
  assign n35703 = \pi0715  & ~n35702 ;
  assign n35704 = \pi0647  & ~n35677 ;
  assign n35705 = n21768 & n35497 ;
  assign n35706 = n21770 & n35497 ;
  assign n35707 = ~n21734 & n35706 ;
  assign n35708 = ~n35705 & ~n35707 ;
  assign n35709 = \pi1157  & n35708 ;
  assign n35710 = ~n35704 & n35709 ;
  assign n35711 = \pi0792  & n35709 ;
  assign n35712 = ~n35699 & n35711 ;
  assign n35713 = ~n35710 & ~n35712 ;
  assign n35714 = ~\pi0647  & ~n35677 ;
  assign n35715 = n21768 & n35502 ;
  assign n35716 = n21770 & n35502 ;
  assign n35717 = ~n21734 & n35716 ;
  assign n35718 = ~n35715 & ~n35717 ;
  assign n35719 = ~\pi1157  & n35718 ;
  assign n35720 = ~n35714 & n35719 ;
  assign n35721 = \pi0792  & n35719 ;
  assign n35722 = ~n35699 & n35721 ;
  assign n35723 = ~n35720 & ~n35722 ;
  assign n35724 = n35713 & n35723 ;
  assign n35725 = n26918 & ~n35724 ;
  assign n35726 = ~n35703 & ~n35725 ;
  assign n35727 = ~\pi0183  & ~n31367 ;
  assign n35728 = n21768 & n35727 ;
  assign n35729 = n21770 & n35727 ;
  assign n35730 = ~n21734 & n35729 ;
  assign n35731 = ~n35728 & ~n35730 ;
  assign n35732 = ~\pi0715  & n35731 ;
  assign n35733 = ~n23958 & ~n35732 ;
  assign n35734 = ~\pi0183  & ~n20811 ;
  assign n35735 = n21768 & n35734 ;
  assign n35736 = n21770 & n35734 ;
  assign n35737 = ~n21734 & n35736 ;
  assign n35738 = ~n35735 & ~n35737 ;
  assign n35739 = ~\pi0183  & \pi0755  ;
  assign n35740 = n21743 & n35739 ;
  assign n35741 = ~n21734 & n35740 ;
  assign n35742 = ~\pi0038  & n35741 ;
  assign n35743 = \pi0183  & ~n25023 ;
  assign n35744 = ~\pi0183  & ~n21467 ;
  assign n35745 = ~\pi0755  & ~n35744 ;
  assign n35746 = ~n35743 & n35745 ;
  assign n35747 = ~\pi0039  & ~\pi0183  ;
  assign n35748 = n21272 & n35747 ;
  assign n35749 = ~\pi0038  & ~n35748 ;
  assign n35750 = n35746 & n35749 ;
  assign n35751 = ~n35742 & ~n35750 ;
  assign n35752 = \pi0038  & n35450 ;
  assign n35753 = n8413 & n35752 ;
  assign n35754 = n1354 & n35753 ;
  assign n35755 = n1358 & n35754 ;
  assign n35756 = \pi0038  & ~\pi0183  ;
  assign n35757 = ~n21757 & n35756 ;
  assign n35758 = ~n35755 & ~n35757 ;
  assign n35759 = n23456 & n35758 ;
  assign n35760 = n35751 & n35759 ;
  assign n35761 = ~n21777 & n35673 ;
  assign n35762 = \pi0183  & ~n6861 ;
  assign n35763 = n21777 & n35762 ;
  assign n35764 = n20811 & ~n35763 ;
  assign n35765 = ~n35761 & n35764 ;
  assign n35766 = ~n35760 & n35765 ;
  assign n35767 = n35738 & ~n35766 ;
  assign n35768 = n23424 & ~n35767 ;
  assign n35769 = ~\pi0781  & ~n35763 ;
  assign n35770 = ~n35761 & n35769 ;
  assign n35771 = ~n35760 & n35770 ;
  assign n35772 = ~n23423 & n35771 ;
  assign n35773 = n23423 & ~n35673 ;
  assign n35774 = ~n35772 & ~n35773 ;
  assign n35775 = ~n35768 & n35774 ;
  assign n35776 = n31382 & ~n35775 ;
  assign n35777 = ~n35733 & ~n35776 ;
  assign n35778 = ~\pi0183  & ~\pi0644  ;
  assign n35779 = n21768 & n35778 ;
  assign n35780 = n21770 & n35778 ;
  assign n35781 = ~n21734 & n35780 ;
  assign n35782 = ~n35779 & ~n35781 ;
  assign n35783 = n35777 & n35782 ;
  assign n35784 = \pi1160  & ~n35783 ;
  assign n35785 = n35726 & n35784 ;
  assign n35786 = \pi0644  & n35701 ;
  assign n35787 = ~\pi0715  & ~n35786 ;
  assign n35788 = n33098 & ~n35724 ;
  assign n35789 = ~n35787 & ~n35788 ;
  assign n35790 = ~\pi0183  & \pi0644  ;
  assign n35791 = n21768 & n35790 ;
  assign n35792 = n21770 & n35790 ;
  assign n35793 = ~n21734 & n35792 ;
  assign n35794 = ~n35791 & ~n35793 ;
  assign n35795 = \pi0715  & n35794 ;
  assign n35796 = ~\pi0644  & ~n35731 ;
  assign n35797 = n34208 & ~n35775 ;
  assign n35798 = ~n35796 & ~n35797 ;
  assign n35799 = n35795 & n35798 ;
  assign n35800 = ~\pi1160  & ~n35799 ;
  assign n35801 = n35789 & n35800 ;
  assign n35802 = ~n35785 & ~n35801 ;
  assign n35803 = \pi0790  & ~n35802 ;
  assign n35804 = n9948 & ~n35624 ;
  assign n35805 = n35803 & n35804 ;
  assign n35806 = n35751 & n35758 ;
  assign n35807 = \pi0725  & ~n35806 ;
  assign n35808 = ~\pi0183  & ~\pi0778  ;
  assign n35809 = ~n23622 & ~n35808 ;
  assign n35810 = n35807 & ~n35809 ;
  assign n35811 = ~\pi0183  & n23548 ;
  assign n35812 = ~\pi0755  & ~n35811 ;
  assign n35813 = ~\pi0039  & ~\pi0755  ;
  assign n35814 = ~n22683 & n35813 ;
  assign n35815 = ~n35812 & ~n35814 ;
  assign n35816 = ~\pi0038  & n35815 ;
  assign n35817 = ~\pi0038  & \pi0183  ;
  assign n35818 = ~n26538 & n35817 ;
  assign n35819 = ~n35816 & ~n35818 ;
  assign n35820 = ~\pi0183  & ~n23567 ;
  assign n35821 = n23565 & n35820 ;
  assign n35822 = \pi0755  & n23575 ;
  assign n35823 = n23572 & n35822 ;
  assign n35824 = ~n35739 & ~n35823 ;
  assign n35825 = ~n35821 & ~n35824 ;
  assign n35826 = ~n35819 & ~n35825 ;
  assign n35827 = n6861 & n35826 ;
  assign n35828 = \pi0183  & ~\pi0755  ;
  assign n35829 = n1689 & n35828 ;
  assign n35830 = n20784 & n35829 ;
  assign n35831 = \pi0183  & \pi0680  ;
  assign n35832 = ~n20854 & n35831 ;
  assign n35833 = ~n20784 & n35832 ;
  assign n35834 = n1689 & n35833 ;
  assign n35835 = ~n35830 & ~n35834 ;
  assign n35836 = n26554 & ~n35835 ;
  assign n35837 = n1358 & n35836 ;
  assign n35838 = \pi0038  & ~n35837 ;
  assign n35839 = ~\pi0725  & ~n35838 ;
  assign n35840 = ~\pi0183  & ~\pi0725  ;
  assign n35841 = ~n26566 & n35840 ;
  assign n35842 = ~\pi0755  & n35840 ;
  assign n35843 = ~n22536 & n35842 ;
  assign n35844 = ~n35841 & ~n35843 ;
  assign n35845 = ~n35839 & n35844 ;
  assign n35846 = n6861 & n35845 ;
  assign n35847 = ~n35809 & ~n35846 ;
  assign n35848 = ~n35827 & n35847 ;
  assign n35849 = ~n35810 & ~n35848 ;
  assign n35850 = \pi0609  & ~n35849 ;
  assign n35851 = ~n22734 & ~n35647 ;
  assign n35852 = n35807 & ~n35851 ;
  assign n35853 = ~n35846 & ~n35851 ;
  assign n35854 = ~n35827 & n35853 ;
  assign n35855 = ~n35852 & ~n35854 ;
  assign n35856 = n6861 & n35758 ;
  assign n35857 = n35751 & n35856 ;
  assign n35858 = ~n22727 & ~n35658 ;
  assign n35859 = ~n35857 & ~n35858 ;
  assign n35860 = ~\pi1153  & ~n35859 ;
  assign n35861 = n35855 & n35860 ;
  assign n35862 = ~\pi0608  & ~n35653 ;
  assign n35863 = ~n35861 & n35862 ;
  assign n35864 = n35807 & ~n35858 ;
  assign n35865 = ~n35846 & ~n35858 ;
  assign n35866 = ~n35827 & n35865 ;
  assign n35867 = ~n35864 & ~n35866 ;
  assign n35868 = ~n35851 & ~n35857 ;
  assign n35869 = \pi1153  & ~n35868 ;
  assign n35870 = n35867 & n35869 ;
  assign n35871 = \pi0608  & ~n35664 ;
  assign n35872 = ~n35870 & n35871 ;
  assign n35873 = ~n35863 & ~n35872 ;
  assign n35874 = n23638 & ~n35873 ;
  assign n35875 = ~n35850 & ~n35874 ;
  assign n35876 = ~n32759 & n35673 ;
  assign n35877 = n26645 & n35758 ;
  assign n35878 = n35751 & n35877 ;
  assign n35879 = ~n20985 & n35762 ;
  assign n35880 = ~\pi0660  & ~n35879 ;
  assign n35881 = ~n35878 & n35880 ;
  assign n35882 = ~n34035 & ~n35881 ;
  assign n35883 = ~n35876 & ~n35882 ;
  assign n35884 = ~\pi0778  & n35633 ;
  assign n35885 = ~n35667 & n35884 ;
  assign n35886 = ~\pi0609  & ~n35885 ;
  assign n35887 = \pi1155  & ~n35886 ;
  assign n35888 = n22722 & ~n35665 ;
  assign n35889 = ~n35887 & ~n35888 ;
  assign n35890 = ~n35883 & ~n35889 ;
  assign n35891 = n35875 & n35890 ;
  assign n35892 = \pi0778  & ~n35873 ;
  assign n35893 = ~n35878 & ~n35879 ;
  assign n35894 = n20999 & ~n35893 ;
  assign n35895 = ~n32768 & n35673 ;
  assign n35896 = ~n22787 & ~n35895 ;
  assign n35897 = ~n35894 & n35896 ;
  assign n35898 = \pi0785  & n35897 ;
  assign n35899 = \pi0778  & ~n35665 ;
  assign n35900 = \pi0609  & ~n35885 ;
  assign n35901 = \pi0785  & n35900 ;
  assign n35902 = ~n35899 & n35901 ;
  assign n35903 = ~n35898 & ~n35902 ;
  assign n35904 = n35849 & n35903 ;
  assign n35905 = ~n35892 & n35904 ;
  assign n35906 = \pi0660  & ~n35895 ;
  assign n35907 = ~n35894 & n35906 ;
  assign n35908 = ~n35883 & ~n35907 ;
  assign n35909 = \pi0609  & ~n35896 ;
  assign n35910 = n35885 & n35909 ;
  assign n35911 = \pi0778  & n35909 ;
  assign n35912 = ~n35665 & n35911 ;
  assign n35913 = ~n35910 & ~n35912 ;
  assign n35914 = ~n35908 & n35913 ;
  assign n35915 = ~n35905 & n35914 ;
  assign n35916 = ~n35891 & n35915 ;
  assign n35917 = ~\pi0785  & ~n35905 ;
  assign n35918 = n26700 & ~n35917 ;
  assign n35919 = ~n35916 & n35918 ;
  assign n35920 = ~n23880 & ~n35775 ;
  assign n35921 = n23880 & ~n35673 ;
  assign n35922 = n24691 & ~n35921 ;
  assign n35923 = ~n35920 & n35922 ;
  assign n35924 = ~\pi0629  & n35687 ;
  assign n35925 = ~n35681 & n35924 ;
  assign n35926 = \pi0629  & n35697 ;
  assign n35927 = ~n35691 & n35926 ;
  assign n35928 = ~n35925 & ~n35927 ;
  assign n35929 = ~n35923 & n35928 ;
  assign n35930 = \pi0792  & ~n35929 ;
  assign n35931 = n23380 & ~n35885 ;
  assign n35932 = ~\pi0183  & ~n23380 ;
  assign n35933 = n21768 & n35932 ;
  assign n35934 = n21770 & n35932 ;
  assign n35935 = ~n21734 & n35934 ;
  assign n35936 = ~n35933 & ~n35935 ;
  assign n35937 = n21050 & n35936 ;
  assign n35938 = ~n35931 & n35937 ;
  assign n35939 = \pi0778  & n35937 ;
  assign n35940 = ~n35665 & n35939 ;
  assign n35941 = ~n35938 & ~n35940 ;
  assign n35942 = n23683 & ~n35767 ;
  assign n35943 = n21032 & n35771 ;
  assign n35944 = ~n21032 & ~n35673 ;
  assign n35945 = ~n20876 & ~n35944 ;
  assign n35946 = ~n35943 & n35945 ;
  assign n35947 = ~n35942 & n35946 ;
  assign n35948 = n35941 & ~n35947 ;
  assign n35949 = \pi0789  & ~n35948 ;
  assign n35950 = n22155 & n35738 ;
  assign n35951 = ~n35766 & n35950 ;
  assign n35952 = ~n21034 & n35951 ;
  assign n35953 = ~n22147 & ~n35885 ;
  assign n35954 = ~n35899 & n35953 ;
  assign n35955 = n22147 & ~n35673 ;
  assign n35956 = n24348 & ~n35955 ;
  assign n35957 = ~n21034 & n35956 ;
  assign n35958 = ~n35954 & n35957 ;
  assign n35959 = ~n35952 & ~n35958 ;
  assign n35960 = ~n21038 & n35959 ;
  assign n35961 = ~n35949 & n35960 ;
  assign n35962 = ~n35930 & n35961 ;
  assign n35963 = ~n35919 & n35962 ;
  assign n35964 = ~n22160 & n35936 ;
  assign n35965 = ~n35931 & n35964 ;
  assign n35966 = \pi0778  & n35964 ;
  assign n35967 = ~n35665 & n35966 ;
  assign n35968 = ~n35965 & ~n35967 ;
  assign n35969 = n22160 & n35673 ;
  assign n35970 = n20951 & ~n35969 ;
  assign n35971 = n35968 & n35970 ;
  assign n35972 = ~\pi0626  & ~n35773 ;
  assign n35973 = ~n35772 & n35972 ;
  assign n35974 = ~n35768 & n35973 ;
  assign n35975 = \pi0626  & n35673 ;
  assign n35976 = n20882 & ~n35975 ;
  assign n35977 = ~n35974 & n35976 ;
  assign n35978 = ~n35971 & ~n35977 ;
  assign n35979 = \pi0626  & ~n35773 ;
  assign n35980 = ~n35772 & n35979 ;
  assign n35981 = ~n35768 & n35980 ;
  assign n35982 = ~\pi0626  & n35673 ;
  assign n35983 = n20881 & ~n35982 ;
  assign n35984 = ~n35981 & n35983 ;
  assign n35985 = ~n23856 & ~n35984 ;
  assign n35986 = n35978 & n35985 ;
  assign n35987 = ~n26803 & ~n35986 ;
  assign n35988 = ~n35930 & n35987 ;
  assign n35989 = ~n21067 & ~n35988 ;
  assign n35990 = ~n35963 & n35989 ;
  assign n35991 = ~n35714 & n35718 ;
  assign n35992 = \pi0792  & n35718 ;
  assign n35993 = ~n35699 & n35992 ;
  assign n35994 = ~n35991 & ~n35993 ;
  assign n35995 = n20897 & ~n35994 ;
  assign n35996 = ~n20846 & n35921 ;
  assign n35997 = n30376 & ~n35775 ;
  assign n35998 = ~n35996 & ~n35997 ;
  assign n35999 = ~n34703 & n35511 ;
  assign n36000 = ~n20910 & ~n35999 ;
  assign n36001 = n35998 & n36000 ;
  assign n36002 = n20849 & n35708 ;
  assign n36003 = ~n35704 & n36002 ;
  assign n36004 = \pi0792  & n36002 ;
  assign n36005 = ~n35699 & n36004 ;
  assign n36006 = ~n36003 & ~n36005 ;
  assign n36007 = ~n36001 & n36006 ;
  assign n36008 = ~n35995 & n36007 ;
  assign n36009 = \pi0787  & ~n36008 ;
  assign n36010 = n26824 & ~n35777 ;
  assign n36011 = \pi0790  & n35795 ;
  assign n36012 = n35798 & n36011 ;
  assign n36013 = ~n35417 & ~n36012 ;
  assign n36014 = ~n36010 & ~n36013 ;
  assign n36015 = ~n36009 & ~n36014 ;
  assign n36016 = n35804 & n36015 ;
  assign n36017 = ~n35990 & n36016 ;
  assign n36018 = ~n35805 & ~n36017 ;
  assign n36019 = ~n35625 & n36018 ;
  assign n36020 = ~\pi0184  & \pi0788  ;
  assign n36021 = ~n1689 & n36020 ;
  assign n36022 = ~n20778 & n36021 ;
  assign n36023 = n20886 & n36022 ;
  assign n36024 = ~\pi0777  & n1689 ;
  assign n36025 = n20784 & n36024 ;
  assign n36026 = n22767 & n36025 ;
  assign n36027 = ~\pi0184  & ~n1689 ;
  assign n36028 = ~n36025 & ~n36027 ;
  assign n36029 = ~n20792 & ~n36028 ;
  assign n36030 = ~n36026 & n36029 ;
  assign n36031 = n20801 & ~n36030 ;
  assign n36032 = ~\pi1155  & ~n36027 ;
  assign n36033 = \pi0785  & n36032 ;
  assign n36034 = ~n36026 & n36033 ;
  assign n36035 = ~\pi0785  & ~n36027 ;
  assign n36036 = ~n36025 & n36035 ;
  assign n36037 = ~n20804 & ~n36036 ;
  assign n36038 = n29682 & n36037 ;
  assign n36039 = ~n36034 & n36038 ;
  assign n36040 = ~n36031 & n36039 ;
  assign n36041 = n30847 & n36040 ;
  assign n36042 = ~n36023 & ~n36041 ;
  assign n36043 = ~\pi0737  & n1689 ;
  assign n36044 = n20855 & n36043 ;
  assign n36045 = ~n36027 & ~n36044 ;
  assign n36046 = ~\pi0778  & ~n36045 ;
  assign n36047 = ~\pi0625  & ~\pi0737  ;
  assign n36048 = n1689 & n36047 ;
  assign n36049 = n20855 & n36048 ;
  assign n36050 = \pi1153  & n36049 ;
  assign n36051 = \pi1153  & ~n36027 ;
  assign n36052 = ~n36044 & n36051 ;
  assign n36053 = ~n36050 & ~n36052 ;
  assign n36054 = ~\pi1153  & ~n36027 ;
  assign n36055 = ~n36049 & n36054 ;
  assign n36056 = \pi0778  & ~n36055 ;
  assign n36057 = n36053 & n36056 ;
  assign n36058 = ~n36046 & ~n36057 ;
  assign n36059 = n26474 & ~n36058 ;
  assign n36060 = \pi0629  & ~n36059 ;
  assign n36061 = n36042 & n36060 ;
  assign n36062 = n20887 & n36022 ;
  assign n36063 = n32579 & n36040 ;
  assign n36064 = ~n36062 & ~n36063 ;
  assign n36065 = n26485 & ~n36058 ;
  assign n36066 = ~\pi0629  & ~n36065 ;
  assign n36067 = n36064 & n36066 ;
  assign n36068 = ~n36061 & ~n36067 ;
  assign n36069 = \pi0792  & n36068 ;
  assign n36070 = ~n21067 & ~n36069 ;
  assign n36071 = n26325 & ~n36058 ;
  assign n36072 = ~\pi0184  & ~\pi0647  ;
  assign n36073 = ~n1689 & n36072 ;
  assign n36074 = n20849 & ~n36073 ;
  assign n36075 = ~n36071 & n36074 ;
  assign n36076 = n26319 & ~n36058 ;
  assign n36077 = ~\pi0184  & \pi0647  ;
  assign n36078 = ~n1689 & n36077 ;
  assign n36079 = n20897 & ~n36078 ;
  assign n36080 = ~n36076 & n36079 ;
  assign n36081 = ~n36075 & ~n36080 ;
  assign n36082 = \pi0787  & ~n36081 ;
  assign n36083 = ~n20846 & n36022 ;
  assign n36084 = n30376 & n36040 ;
  assign n36085 = ~n36083 & ~n36084 ;
  assign n36086 = ~\pi0184  & \pi0792  ;
  assign n36087 = ~n1689 & n36086 ;
  assign n36088 = ~n20845 & n36087 ;
  assign n36089 = n32606 & ~n36088 ;
  assign n36090 = n36085 & n36089 ;
  assign n36091 = ~n36082 & ~n36090 ;
  assign n36092 = ~n24761 & n36091 ;
  assign n36093 = ~n36070 & n36092 ;
  assign n36094 = \pi0608  & ~n36055 ;
  assign n36095 = ~n36025 & n36051 ;
  assign n36096 = \pi0778  & ~n36095 ;
  assign n36097 = n26421 & ~n36045 ;
  assign n36098 = ~n36096 & ~n36097 ;
  assign n36099 = n36094 & ~n36098 ;
  assign n36100 = n26147 & ~n36045 ;
  assign n36101 = ~\pi0737  & ~n20784 ;
  assign n36102 = n22113 & n36101 ;
  assign n36103 = n36028 & ~n36102 ;
  assign n36104 = ~n36100 & ~n36103 ;
  assign n36105 = n36054 & ~n36104 ;
  assign n36106 = n26415 & n36053 ;
  assign n36107 = ~n36105 & n36106 ;
  assign n36108 = ~n36099 & ~n36107 ;
  assign n36109 = ~\pi1155  & ~n36046 ;
  assign n36110 = ~n36057 & n36109 ;
  assign n36111 = ~n20999 & ~n36110 ;
  assign n36112 = ~\pi0778  & ~n36103 ;
  assign n36113 = ~n36111 & ~n36112 ;
  assign n36114 = n36108 & n36113 ;
  assign n36115 = n29766 & ~n36046 ;
  assign n36116 = ~n36057 & n36115 ;
  assign n36117 = \pi1155  & ~n36030 ;
  assign n36118 = ~\pi0660  & ~n36117 ;
  assign n36119 = ~n36116 & n36118 ;
  assign n36120 = ~n36114 & n36119 ;
  assign n36121 = \pi0785  & ~n36120 ;
  assign n36122 = n29775 & n36037 ;
  assign n36123 = ~n36034 & n36122 ;
  assign n36124 = ~n36031 & n36123 ;
  assign n36125 = n29779 & ~n36058 ;
  assign n36126 = ~n36124 & ~n36125 ;
  assign n36127 = \pi0781  & ~n36126 ;
  assign n36128 = \pi1155  & ~n36046 ;
  assign n36129 = ~n36057 & n36128 ;
  assign n36130 = ~n21774 & ~n36129 ;
  assign n36131 = ~n36112 & ~n36130 ;
  assign n36132 = n36108 & n36131 ;
  assign n36133 = n26121 & ~n36046 ;
  assign n36134 = ~n36057 & n36133 ;
  assign n36135 = \pi0660  & ~n36032 ;
  assign n36136 = \pi0660  & n36025 ;
  assign n36137 = n22767 & n36136 ;
  assign n36138 = ~n36135 & ~n36137 ;
  assign n36139 = ~n36134 & ~n36138 ;
  assign n36140 = ~n36132 & n36139 ;
  assign n36141 = ~n36127 & ~n36140 ;
  assign n36142 = n36121 & n36141 ;
  assign n36143 = ~\pi0785  & ~n36112 ;
  assign n36144 = ~n36099 & n36143 ;
  assign n36145 = ~n36107 & n36144 ;
  assign n36146 = n21022 & ~n36145 ;
  assign n36147 = ~n36127 & ~n36146 ;
  assign n36148 = n29803 & ~n36147 ;
  assign n36149 = ~n36142 & n36148 ;
  assign n36150 = n29808 & n36037 ;
  assign n36151 = ~n36034 & n36150 ;
  assign n36152 = ~n36031 & n36151 ;
  assign n36153 = n30966 & ~n36058 ;
  assign n36154 = ~n36152 & ~n36153 ;
  assign n36155 = \pi0789  & ~n21038 ;
  assign n36156 = ~n36154 & n36155 ;
  assign n36157 = \pi0626  & ~n36040 ;
  assign n36158 = ~\pi0626  & ~n36027 ;
  assign n36159 = n20881 & ~n36158 ;
  assign n36160 = ~n36157 & n36159 ;
  assign n36161 = n26458 & ~n36058 ;
  assign n36162 = ~\pi0626  & ~n36040 ;
  assign n36163 = \pi0626  & ~n36027 ;
  assign n36164 = n20882 & ~n36163 ;
  assign n36165 = ~n36162 & n36164 ;
  assign n36166 = ~n36161 & ~n36165 ;
  assign n36167 = ~n36160 & n36166 ;
  assign n36168 = \pi0788  & ~n36167 ;
  assign n36169 = ~n36156 & ~n36168 ;
  assign n36170 = ~n36149 & n36169 ;
  assign n36171 = ~n23856 & n36092 ;
  assign n36172 = ~n36170 & n36171 ;
  assign n36173 = ~n36093 & ~n36172 ;
  assign n36174 = n30987 & ~n36085 ;
  assign n36175 = n23312 & n36174 ;
  assign n36176 = \pi1157  & ~n36073 ;
  assign n36177 = ~n36071 & n36176 ;
  assign n36178 = ~\pi1157  & ~n36078 ;
  assign n36179 = ~n36076 & n36178 ;
  assign n36180 = ~n36177 & ~n36179 ;
  assign n36181 = \pi0787  & ~n36180 ;
  assign n36182 = n26333 & ~n36058 ;
  assign n36183 = ~\pi0787  & ~n36182 ;
  assign n36184 = ~\pi1160  & ~n36183 ;
  assign n36185 = n23312 & n36184 ;
  assign n36186 = ~n36181 & n36185 ;
  assign n36187 = ~n36175 & ~n36186 ;
  assign n36188 = ~n23414 & n36027 ;
  assign n36189 = ~n24886 & n36188 ;
  assign n36190 = ~n23313 & ~n36189 ;
  assign n36191 = \pi1160  & ~n36183 ;
  assign n36192 = ~n36181 & n36191 ;
  assign n36193 = n31010 & ~n36085 ;
  assign n36194 = ~n36189 & ~n36193 ;
  assign n36195 = ~n36192 & n36194 ;
  assign n36196 = ~n36190 & ~n36195 ;
  assign n36197 = n36187 & ~n36196 ;
  assign n36198 = \pi0790  & ~n36197 ;
  assign n36199 = \pi0832  & ~n36198 ;
  assign n36200 = n36173 & n36199 ;
  assign n36201 = \pi0184  & ~\pi0832  ;
  assign n36202 = ~n21132 & ~n36201 ;
  assign n36203 = ~n36200 & n36202 ;
  assign n36204 = ~\pi0074  & ~\pi0737  ;
  assign n36205 = ~\pi0100  & n36204 ;
  assign n36206 = n1287 & n36205 ;
  assign n36207 = ~\pi0184  & ~n36206 ;
  assign n36208 = n21768 & n36207 ;
  assign n36209 = n21770 & n36207 ;
  assign n36210 = ~n21734 & n36209 ;
  assign n36211 = ~n36208 & ~n36210 ;
  assign n36212 = \pi0625  & ~n36211 ;
  assign n36213 = ~\pi0184  & ~n22017 ;
  assign n36214 = ~n21994 & n36213 ;
  assign n36215 = ~\pi0038  & ~\pi0184  ;
  assign n36216 = n6861 & ~n36215 ;
  assign n36217 = ~n22109 & n36216 ;
  assign n36218 = ~n36214 & ~n36217 ;
  assign n36219 = ~\pi0184  & ~n21757 ;
  assign n36220 = n22117 & ~n36219 ;
  assign n36221 = ~\pi0737  & ~n36220 ;
  assign n36222 = \pi0625  & n36221 ;
  assign n36223 = ~n36218 & n36222 ;
  assign n36224 = ~n36212 & ~n36223 ;
  assign n36225 = ~\pi0184  & ~\pi0625  ;
  assign n36226 = n21768 & n36225 ;
  assign n36227 = n21770 & n36225 ;
  assign n36228 = ~n21734 & n36227 ;
  assign n36229 = ~n36226 & ~n36228 ;
  assign n36230 = \pi1153  & n36229 ;
  assign n36231 = n36224 & n36230 ;
  assign n36232 = ~\pi0625  & ~n36211 ;
  assign n36233 = ~\pi0625  & n36221 ;
  assign n36234 = ~n36218 & n36233 ;
  assign n36235 = ~n36232 & ~n36234 ;
  assign n36236 = ~\pi0184  & \pi0625  ;
  assign n36237 = n21768 & n36236 ;
  assign n36238 = n21770 & n36236 ;
  assign n36239 = ~n21734 & n36238 ;
  assign n36240 = ~n36237 & ~n36239 ;
  assign n36241 = ~\pi1153  & n36240 ;
  assign n36242 = n36235 & n36241 ;
  assign n36243 = ~n36231 & ~n36242 ;
  assign n36244 = n26065 & ~n36243 ;
  assign n36245 = ~n36218 & n36221 ;
  assign n36246 = n26739 & n36211 ;
  assign n36247 = ~n36245 & n36246 ;
  assign n36248 = ~\pi0184  & n21768 ;
  assign n36249 = ~\pi0184  & n21770 ;
  assign n36250 = ~n21734 & n36249 ;
  assign n36251 = ~n36248 & ~n36250 ;
  assign n36252 = ~n23885 & n36251 ;
  assign n36253 = ~n36247 & ~n36252 ;
  assign n36254 = ~n36244 & n36253 ;
  assign n36255 = ~\pi0792  & ~n36254 ;
  assign n36256 = ~\pi0787  & n36255 ;
  assign n36257 = \pi0628  & ~n36252 ;
  assign n36258 = ~n36247 & n36257 ;
  assign n36259 = ~n36244 & n36258 ;
  assign n36260 = ~\pi0184  & ~\pi0628  ;
  assign n36261 = n21768 & n36260 ;
  assign n36262 = n21770 & n36260 ;
  assign n36263 = ~n21734 & n36262 ;
  assign n36264 = ~n36261 & ~n36263 ;
  assign n36265 = \pi1156  & n36264 ;
  assign n36266 = ~n36259 & n36265 ;
  assign n36267 = ~\pi0628  & ~n36252 ;
  assign n36268 = ~n36247 & n36267 ;
  assign n36269 = ~n36244 & n36268 ;
  assign n36270 = ~\pi0184  & \pi0628  ;
  assign n36271 = n21768 & n36270 ;
  assign n36272 = n21770 & n36270 ;
  assign n36273 = ~n21734 & n36272 ;
  assign n36274 = ~n36271 & ~n36273 ;
  assign n36275 = ~\pi1156  & n36274 ;
  assign n36276 = ~n36269 & n36275 ;
  assign n36277 = ~n36266 & ~n36276 ;
  assign n36278 = n33084 & ~n36277 ;
  assign n36279 = ~n36256 & ~n36278 ;
  assign n36280 = ~\pi0644  & n36279 ;
  assign n36281 = \pi0715  & ~n36280 ;
  assign n36282 = \pi0647  & ~n36255 ;
  assign n36283 = n21768 & n36072 ;
  assign n36284 = n21770 & n36072 ;
  assign n36285 = ~n21734 & n36284 ;
  assign n36286 = ~n36283 & ~n36285 ;
  assign n36287 = \pi1157  & n36286 ;
  assign n36288 = ~n36282 & n36287 ;
  assign n36289 = \pi0792  & n36287 ;
  assign n36290 = ~n36277 & n36289 ;
  assign n36291 = ~n36288 & ~n36290 ;
  assign n36292 = ~\pi0647  & ~n36255 ;
  assign n36293 = n21768 & n36077 ;
  assign n36294 = n21770 & n36077 ;
  assign n36295 = ~n21734 & n36294 ;
  assign n36296 = ~n36293 & ~n36295 ;
  assign n36297 = ~\pi1157  & n36296 ;
  assign n36298 = ~n36292 & n36297 ;
  assign n36299 = \pi0792  & n36297 ;
  assign n36300 = ~n36277 & n36299 ;
  assign n36301 = ~n36298 & ~n36300 ;
  assign n36302 = n36291 & n36301 ;
  assign n36303 = n26918 & ~n36302 ;
  assign n36304 = ~n36281 & ~n36303 ;
  assign n36305 = ~\pi0184  & ~n31367 ;
  assign n36306 = n21768 & n36305 ;
  assign n36307 = n21770 & n36305 ;
  assign n36308 = ~n21734 & n36307 ;
  assign n36309 = ~n36306 & ~n36308 ;
  assign n36310 = ~\pi0715  & n36309 ;
  assign n36311 = ~n23958 & ~n36310 ;
  assign n36312 = ~\pi0184  & ~n20811 ;
  assign n36313 = n21768 & n36312 ;
  assign n36314 = n21770 & n36312 ;
  assign n36315 = ~n21734 & n36314 ;
  assign n36316 = ~n36313 & ~n36315 ;
  assign n36317 = ~\pi0184  & \pi0777  ;
  assign n36318 = n21743 & n36317 ;
  assign n36319 = ~n21734 & n36318 ;
  assign n36320 = ~\pi0038  & n36319 ;
  assign n36321 = \pi0184  & ~n25023 ;
  assign n36322 = ~\pi0184  & ~n21467 ;
  assign n36323 = ~\pi0777  & ~n36322 ;
  assign n36324 = ~n36321 & n36323 ;
  assign n36325 = ~\pi0039  & ~\pi0184  ;
  assign n36326 = n21272 & n36325 ;
  assign n36327 = ~\pi0038  & ~n36326 ;
  assign n36328 = n36324 & n36327 ;
  assign n36329 = ~n36320 & ~n36328 ;
  assign n36330 = \pi0038  & n36025 ;
  assign n36331 = n8413 & n36330 ;
  assign n36332 = n1354 & n36331 ;
  assign n36333 = n1358 & n36332 ;
  assign n36334 = \pi0038  & ~\pi0184  ;
  assign n36335 = ~n21757 & n36334 ;
  assign n36336 = ~n36333 & ~n36335 ;
  assign n36337 = n23456 & n36336 ;
  assign n36338 = n36329 & n36337 ;
  assign n36339 = ~n21777 & n36251 ;
  assign n36340 = \pi0184  & ~n6861 ;
  assign n36341 = n21777 & n36340 ;
  assign n36342 = n20811 & ~n36341 ;
  assign n36343 = ~n36339 & n36342 ;
  assign n36344 = ~n36338 & n36343 ;
  assign n36345 = n36316 & ~n36344 ;
  assign n36346 = n23424 & ~n36345 ;
  assign n36347 = ~\pi0781  & ~n36341 ;
  assign n36348 = ~n36339 & n36347 ;
  assign n36349 = ~n36338 & n36348 ;
  assign n36350 = ~n23423 & n36349 ;
  assign n36351 = n23423 & ~n36251 ;
  assign n36352 = ~n36350 & ~n36351 ;
  assign n36353 = ~n36346 & n36352 ;
  assign n36354 = n31382 & ~n36353 ;
  assign n36355 = ~n36311 & ~n36354 ;
  assign n36356 = ~\pi0184  & ~\pi0644  ;
  assign n36357 = n21768 & n36356 ;
  assign n36358 = n21770 & n36356 ;
  assign n36359 = ~n21734 & n36358 ;
  assign n36360 = ~n36357 & ~n36359 ;
  assign n36361 = n36355 & n36360 ;
  assign n36362 = \pi1160  & ~n36361 ;
  assign n36363 = n36304 & n36362 ;
  assign n36364 = \pi0644  & n36279 ;
  assign n36365 = ~\pi0715  & ~n36364 ;
  assign n36366 = n33098 & ~n36302 ;
  assign n36367 = ~n36365 & ~n36366 ;
  assign n36368 = ~\pi0184  & \pi0644  ;
  assign n36369 = n21768 & n36368 ;
  assign n36370 = n21770 & n36368 ;
  assign n36371 = ~n21734 & n36370 ;
  assign n36372 = ~n36369 & ~n36371 ;
  assign n36373 = \pi0715  & n36372 ;
  assign n36374 = ~\pi0644  & ~n36309 ;
  assign n36375 = n34208 & ~n36353 ;
  assign n36376 = ~n36374 & ~n36375 ;
  assign n36377 = n36373 & n36376 ;
  assign n36378 = ~\pi1160  & ~n36377 ;
  assign n36379 = n36367 & n36378 ;
  assign n36380 = ~n36363 & ~n36379 ;
  assign n36381 = \pi0790  & ~n36380 ;
  assign n36382 = n9948 & ~n36200 ;
  assign n36383 = n36381 & n36382 ;
  assign n36384 = n36329 & n36336 ;
  assign n36385 = \pi0737  & ~n36384 ;
  assign n36386 = ~\pi0184  & ~\pi0778  ;
  assign n36387 = ~n23622 & ~n36386 ;
  assign n36388 = n36385 & ~n36387 ;
  assign n36389 = ~\pi0184  & n23548 ;
  assign n36390 = ~\pi0777  & ~n36389 ;
  assign n36391 = ~\pi0039  & ~\pi0777  ;
  assign n36392 = ~n22683 & n36391 ;
  assign n36393 = ~n36390 & ~n36392 ;
  assign n36394 = ~\pi0038  & n36393 ;
  assign n36395 = ~\pi0038  & \pi0184  ;
  assign n36396 = ~n26538 & n36395 ;
  assign n36397 = ~n36394 & ~n36396 ;
  assign n36398 = ~\pi0184  & ~n23567 ;
  assign n36399 = n23565 & n36398 ;
  assign n36400 = \pi0777  & n23575 ;
  assign n36401 = n23572 & n36400 ;
  assign n36402 = ~n36317 & ~n36401 ;
  assign n36403 = ~n36399 & ~n36402 ;
  assign n36404 = ~n36397 & ~n36403 ;
  assign n36405 = n6861 & n36404 ;
  assign n36406 = \pi0184  & \pi0603  ;
  assign n36407 = ~n20783 & n36406 ;
  assign n36408 = n36024 & n36407 ;
  assign n36409 = \pi0184  & \pi0680  ;
  assign n36410 = ~n20854 & n36409 ;
  assign n36411 = ~n20784 & n36410 ;
  assign n36412 = n1689 & n36411 ;
  assign n36413 = ~n36408 & ~n36412 ;
  assign n36414 = n26554 & ~n36413 ;
  assign n36415 = n1358 & n36414 ;
  assign n36416 = \pi0038  & ~n36415 ;
  assign n36417 = ~\pi0737  & ~n36416 ;
  assign n36418 = ~\pi0184  & ~\pi0737  ;
  assign n36419 = ~n26566 & n36418 ;
  assign n36420 = ~\pi0777  & n36418 ;
  assign n36421 = ~n22536 & n36420 ;
  assign n36422 = ~n36419 & ~n36421 ;
  assign n36423 = ~n36417 & n36422 ;
  assign n36424 = n6861 & n36423 ;
  assign n36425 = ~n36387 & ~n36424 ;
  assign n36426 = ~n36405 & n36425 ;
  assign n36427 = ~n36388 & ~n36426 ;
  assign n36428 = \pi0609  & ~n36427 ;
  assign n36429 = ~n22734 & ~n36225 ;
  assign n36430 = n36385 & ~n36429 ;
  assign n36431 = ~n36424 & ~n36429 ;
  assign n36432 = ~n36405 & n36431 ;
  assign n36433 = ~n36430 & ~n36432 ;
  assign n36434 = n6861 & n36336 ;
  assign n36435 = n36329 & n36434 ;
  assign n36436 = ~n22727 & ~n36236 ;
  assign n36437 = ~n36435 & ~n36436 ;
  assign n36438 = ~\pi1153  & ~n36437 ;
  assign n36439 = n36433 & n36438 ;
  assign n36440 = ~\pi0608  & ~n36231 ;
  assign n36441 = ~n36439 & n36440 ;
  assign n36442 = n36385 & ~n36436 ;
  assign n36443 = ~n36424 & ~n36436 ;
  assign n36444 = ~n36405 & n36443 ;
  assign n36445 = ~n36442 & ~n36444 ;
  assign n36446 = ~n36429 & ~n36435 ;
  assign n36447 = \pi1153  & ~n36446 ;
  assign n36448 = n36445 & n36447 ;
  assign n36449 = \pi0608  & ~n36242 ;
  assign n36450 = ~n36448 & n36449 ;
  assign n36451 = ~n36441 & ~n36450 ;
  assign n36452 = n23638 & ~n36451 ;
  assign n36453 = ~n36428 & ~n36452 ;
  assign n36454 = n26653 & n36251 ;
  assign n36455 = n26645 & n36336 ;
  assign n36456 = n36329 & n36455 ;
  assign n36457 = ~n20985 & n36340 ;
  assign n36458 = ~\pi0660  & ~n36457 ;
  assign n36459 = ~n36456 & n36458 ;
  assign n36460 = ~n34035 & ~n36459 ;
  assign n36461 = ~n36454 & ~n36460 ;
  assign n36462 = ~\pi0778  & n36211 ;
  assign n36463 = ~n36245 & n36462 ;
  assign n36464 = ~\pi0609  & ~n36463 ;
  assign n36465 = \pi1155  & ~n36464 ;
  assign n36466 = n22722 & ~n36243 ;
  assign n36467 = ~n36465 & ~n36466 ;
  assign n36468 = ~n36461 & ~n36467 ;
  assign n36469 = n36453 & n36468 ;
  assign n36470 = \pi0778  & ~n36451 ;
  assign n36471 = ~n36456 & ~n36457 ;
  assign n36472 = n20999 & ~n36471 ;
  assign n36473 = ~n32768 & n36251 ;
  assign n36474 = ~n22787 & ~n36473 ;
  assign n36475 = ~n36472 & n36474 ;
  assign n36476 = \pi0785  & n36475 ;
  assign n36477 = \pi0778  & ~n36243 ;
  assign n36478 = \pi0609  & ~n36463 ;
  assign n36479 = \pi0785  & n36478 ;
  assign n36480 = ~n36477 & n36479 ;
  assign n36481 = ~n36476 & ~n36480 ;
  assign n36482 = n36427 & n36481 ;
  assign n36483 = ~n36470 & n36482 ;
  assign n36484 = \pi0660  & ~n36473 ;
  assign n36485 = ~n36472 & n36484 ;
  assign n36486 = ~n36461 & ~n36485 ;
  assign n36487 = \pi0609  & ~n36474 ;
  assign n36488 = n36463 & n36487 ;
  assign n36489 = \pi0778  & n36487 ;
  assign n36490 = ~n36243 & n36489 ;
  assign n36491 = ~n36488 & ~n36490 ;
  assign n36492 = ~n36486 & n36491 ;
  assign n36493 = ~n36483 & n36492 ;
  assign n36494 = ~n36469 & n36493 ;
  assign n36495 = ~\pi0785  & ~n36483 ;
  assign n36496 = n26700 & ~n36495 ;
  assign n36497 = ~n36494 & n36496 ;
  assign n36498 = ~n23880 & ~n36353 ;
  assign n36499 = n23880 & ~n36251 ;
  assign n36500 = n24691 & ~n36499 ;
  assign n36501 = ~n36498 & n36500 ;
  assign n36502 = ~\pi0629  & n36265 ;
  assign n36503 = ~n36259 & n36502 ;
  assign n36504 = \pi0629  & n36275 ;
  assign n36505 = ~n36269 & n36504 ;
  assign n36506 = ~n36503 & ~n36505 ;
  assign n36507 = ~n36501 & n36506 ;
  assign n36508 = \pi0792  & ~n36507 ;
  assign n36509 = n23380 & ~n36463 ;
  assign n36510 = ~\pi0184  & ~n23380 ;
  assign n36511 = n21768 & n36510 ;
  assign n36512 = n21770 & n36510 ;
  assign n36513 = ~n21734 & n36512 ;
  assign n36514 = ~n36511 & ~n36513 ;
  assign n36515 = n21050 & n36514 ;
  assign n36516 = ~n36509 & n36515 ;
  assign n36517 = \pi0778  & n36515 ;
  assign n36518 = ~n36243 & n36517 ;
  assign n36519 = ~n36516 & ~n36518 ;
  assign n36520 = n23683 & ~n36345 ;
  assign n36521 = n21032 & n36349 ;
  assign n36522 = ~n21032 & ~n36251 ;
  assign n36523 = ~n20876 & ~n36522 ;
  assign n36524 = ~n36521 & n36523 ;
  assign n36525 = ~n36520 & n36524 ;
  assign n36526 = n36519 & ~n36525 ;
  assign n36527 = \pi0789  & ~n36526 ;
  assign n36528 = n22155 & n36316 ;
  assign n36529 = ~n36344 & n36528 ;
  assign n36530 = ~n21034 & n36529 ;
  assign n36531 = ~n22147 & ~n36463 ;
  assign n36532 = ~n36477 & n36531 ;
  assign n36533 = n22147 & ~n36251 ;
  assign n36534 = n24348 & ~n36533 ;
  assign n36535 = ~n21034 & n36534 ;
  assign n36536 = ~n36532 & n36535 ;
  assign n36537 = ~n36530 & ~n36536 ;
  assign n36538 = ~n21038 & n36537 ;
  assign n36539 = ~n36527 & n36538 ;
  assign n36540 = ~n36508 & n36539 ;
  assign n36541 = ~n36497 & n36540 ;
  assign n36542 = ~n22160 & n36514 ;
  assign n36543 = ~n36509 & n36542 ;
  assign n36544 = \pi0778  & n36542 ;
  assign n36545 = ~n36243 & n36544 ;
  assign n36546 = ~n36543 & ~n36545 ;
  assign n36547 = n22160 & n36251 ;
  assign n36548 = n20951 & ~n36547 ;
  assign n36549 = n36546 & n36548 ;
  assign n36550 = ~\pi0626  & ~n36351 ;
  assign n36551 = ~n36350 & n36550 ;
  assign n36552 = ~n36346 & n36551 ;
  assign n36553 = \pi0626  & n36251 ;
  assign n36554 = n20882 & ~n36553 ;
  assign n36555 = ~n36552 & n36554 ;
  assign n36556 = ~n36549 & ~n36555 ;
  assign n36557 = \pi0626  & ~n36351 ;
  assign n36558 = ~n36350 & n36557 ;
  assign n36559 = ~n36346 & n36558 ;
  assign n36560 = ~\pi0626  & n36251 ;
  assign n36561 = n20881 & ~n36560 ;
  assign n36562 = ~n36559 & n36561 ;
  assign n36563 = ~n23856 & ~n36562 ;
  assign n36564 = n36556 & n36563 ;
  assign n36565 = ~n26803 & ~n36564 ;
  assign n36566 = ~n36508 & n36565 ;
  assign n36567 = ~n21067 & ~n36566 ;
  assign n36568 = ~n36541 & n36567 ;
  assign n36569 = \pi0630  & ~n36301 ;
  assign n36570 = ~n20846 & n36499 ;
  assign n36571 = n30376 & ~n36353 ;
  assign n36572 = ~n36570 & ~n36571 ;
  assign n36573 = ~n34703 & n36086 ;
  assign n36574 = ~n20910 & ~n36573 ;
  assign n36575 = n36572 & n36574 ;
  assign n36576 = n20849 & n36286 ;
  assign n36577 = ~n36282 & n36576 ;
  assign n36578 = \pi0792  & n36576 ;
  assign n36579 = ~n36277 & n36578 ;
  assign n36580 = ~n36577 & ~n36579 ;
  assign n36581 = ~n36575 & n36580 ;
  assign n36582 = ~n36569 & n36581 ;
  assign n36583 = \pi0787  & ~n36582 ;
  assign n36584 = n26824 & ~n36355 ;
  assign n36585 = \pi0790  & n36373 ;
  assign n36586 = n36376 & n36585 ;
  assign n36587 = ~n35417 & ~n36586 ;
  assign n36588 = ~n36584 & ~n36587 ;
  assign n36589 = ~n36583 & ~n36588 ;
  assign n36590 = n36382 & n36589 ;
  assign n36591 = ~n36568 & n36590 ;
  assign n36592 = ~n36383 & ~n36591 ;
  assign n36593 = ~n36203 & n36592 ;
  assign n36594 = ~\pi0185  & \pi0788  ;
  assign n36595 = ~n1689 & n36594 ;
  assign n36596 = ~n20778 & n36595 ;
  assign n36597 = n20886 & n36596 ;
  assign n36598 = ~\pi0751  & n1689 ;
  assign n36599 = n20784 & n36598 ;
  assign n36600 = n22767 & n36599 ;
  assign n36601 = ~\pi0185  & ~n1689 ;
  assign n36602 = ~n36599 & ~n36601 ;
  assign n36603 = ~n20792 & ~n36602 ;
  assign n36604 = ~n36600 & n36603 ;
  assign n36605 = n20801 & ~n36604 ;
  assign n36606 = ~\pi1155  & ~n36601 ;
  assign n36607 = \pi0785  & n36606 ;
  assign n36608 = ~n36600 & n36607 ;
  assign n36609 = ~\pi0785  & ~n36601 ;
  assign n36610 = ~n36599 & n36609 ;
  assign n36611 = ~n20804 & ~n36610 ;
  assign n36612 = n29682 & n36611 ;
  assign n36613 = ~n36608 & n36612 ;
  assign n36614 = ~n36605 & n36613 ;
  assign n36615 = n30847 & n36614 ;
  assign n36616 = ~n36597 & ~n36615 ;
  assign n36617 = ~\pi0701  & n1689 ;
  assign n36618 = n20855 & n36617 ;
  assign n36619 = ~n36601 & ~n36618 ;
  assign n36620 = ~\pi0778  & ~n36619 ;
  assign n36621 = ~\pi0625  & ~\pi0701  ;
  assign n36622 = n1689 & n36621 ;
  assign n36623 = n20855 & n36622 ;
  assign n36624 = \pi1153  & n36623 ;
  assign n36625 = \pi1153  & ~n36601 ;
  assign n36626 = ~n36618 & n36625 ;
  assign n36627 = ~n36624 & ~n36626 ;
  assign n36628 = ~\pi1153  & ~n36601 ;
  assign n36629 = ~n36623 & n36628 ;
  assign n36630 = \pi0778  & ~n36629 ;
  assign n36631 = n36627 & n36630 ;
  assign n36632 = ~n36620 & ~n36631 ;
  assign n36633 = n26474 & ~n36632 ;
  assign n36634 = \pi0629  & ~n36633 ;
  assign n36635 = n36616 & n36634 ;
  assign n36636 = n20887 & n36596 ;
  assign n36637 = n32579 & n36614 ;
  assign n36638 = ~n36636 & ~n36637 ;
  assign n36639 = n26485 & ~n36632 ;
  assign n36640 = ~\pi0629  & ~n36639 ;
  assign n36641 = n36638 & n36640 ;
  assign n36642 = ~n36635 & ~n36641 ;
  assign n36643 = \pi0792  & n36642 ;
  assign n36644 = ~n21067 & ~n36643 ;
  assign n36645 = n26325 & ~n36632 ;
  assign n36646 = ~\pi0185  & ~\pi0647  ;
  assign n36647 = ~n1689 & n36646 ;
  assign n36648 = n20849 & ~n36647 ;
  assign n36649 = ~n36645 & n36648 ;
  assign n36650 = n26319 & ~n36632 ;
  assign n36651 = ~\pi0185  & \pi0647  ;
  assign n36652 = ~n1689 & n36651 ;
  assign n36653 = n20897 & ~n36652 ;
  assign n36654 = ~n36650 & n36653 ;
  assign n36655 = ~n36649 & ~n36654 ;
  assign n36656 = \pi0787  & ~n36655 ;
  assign n36657 = ~n20846 & n36596 ;
  assign n36658 = n30376 & n36614 ;
  assign n36659 = ~n36657 & ~n36658 ;
  assign n36660 = ~\pi0185  & \pi0792  ;
  assign n36661 = ~n1689 & n36660 ;
  assign n36662 = ~n20845 & n36661 ;
  assign n36663 = n32606 & ~n36662 ;
  assign n36664 = n36659 & n36663 ;
  assign n36665 = ~n36656 & ~n36664 ;
  assign n36666 = ~n24761 & n36665 ;
  assign n36667 = ~n36644 & n36666 ;
  assign n36668 = \pi0608  & ~n36629 ;
  assign n36669 = ~n36599 & n36625 ;
  assign n36670 = \pi0778  & ~n36669 ;
  assign n36671 = n26421 & ~n36619 ;
  assign n36672 = ~n36670 & ~n36671 ;
  assign n36673 = n36668 & ~n36672 ;
  assign n36674 = n26147 & ~n36619 ;
  assign n36675 = ~\pi0701  & ~n20784 ;
  assign n36676 = n22113 & n36675 ;
  assign n36677 = n36602 & ~n36676 ;
  assign n36678 = ~n36674 & ~n36677 ;
  assign n36679 = n36628 & ~n36678 ;
  assign n36680 = n26415 & n36627 ;
  assign n36681 = ~n36679 & n36680 ;
  assign n36682 = ~n36673 & ~n36681 ;
  assign n36683 = ~\pi1155  & ~n36620 ;
  assign n36684 = ~n36631 & n36683 ;
  assign n36685 = ~n20999 & ~n36684 ;
  assign n36686 = ~\pi0778  & ~n36677 ;
  assign n36687 = ~n36685 & ~n36686 ;
  assign n36688 = n36682 & n36687 ;
  assign n36689 = n29766 & ~n36620 ;
  assign n36690 = ~n36631 & n36689 ;
  assign n36691 = \pi1155  & ~n36604 ;
  assign n36692 = ~\pi0660  & ~n36691 ;
  assign n36693 = ~n36690 & n36692 ;
  assign n36694 = ~n36688 & n36693 ;
  assign n36695 = \pi0785  & ~n36694 ;
  assign n36696 = n29775 & n36611 ;
  assign n36697 = ~n36608 & n36696 ;
  assign n36698 = ~n36605 & n36697 ;
  assign n36699 = n29779 & ~n36632 ;
  assign n36700 = ~n36698 & ~n36699 ;
  assign n36701 = \pi0781  & ~n36700 ;
  assign n36702 = \pi1155  & ~n36620 ;
  assign n36703 = ~n36631 & n36702 ;
  assign n36704 = ~n21774 & ~n36703 ;
  assign n36705 = ~n36686 & ~n36704 ;
  assign n36706 = n36682 & n36705 ;
  assign n36707 = n26121 & ~n36620 ;
  assign n36708 = ~n36631 & n36707 ;
  assign n36709 = \pi0660  & ~n36606 ;
  assign n36710 = \pi0660  & n36599 ;
  assign n36711 = n22767 & n36710 ;
  assign n36712 = ~n36709 & ~n36711 ;
  assign n36713 = ~n36708 & ~n36712 ;
  assign n36714 = ~n36706 & n36713 ;
  assign n36715 = ~n36701 & ~n36714 ;
  assign n36716 = n36695 & n36715 ;
  assign n36717 = ~\pi0785  & ~n36686 ;
  assign n36718 = ~n36673 & n36717 ;
  assign n36719 = ~n36681 & n36718 ;
  assign n36720 = n21022 & ~n36719 ;
  assign n36721 = ~n36701 & ~n36720 ;
  assign n36722 = n29803 & ~n36721 ;
  assign n36723 = ~n36716 & n36722 ;
  assign n36724 = n29808 & n36611 ;
  assign n36725 = ~n36608 & n36724 ;
  assign n36726 = ~n36605 & n36725 ;
  assign n36727 = n30966 & ~n36632 ;
  assign n36728 = ~n36726 & ~n36727 ;
  assign n36729 = n36155 & ~n36728 ;
  assign n36730 = \pi0626  & ~n36614 ;
  assign n36731 = ~\pi0626  & ~n36601 ;
  assign n36732 = n20881 & ~n36731 ;
  assign n36733 = ~n36730 & n36732 ;
  assign n36734 = n26458 & ~n36632 ;
  assign n36735 = ~\pi0626  & ~n36614 ;
  assign n36736 = \pi0626  & ~n36601 ;
  assign n36737 = n20882 & ~n36736 ;
  assign n36738 = ~n36735 & n36737 ;
  assign n36739 = ~n36734 & ~n36738 ;
  assign n36740 = ~n36733 & n36739 ;
  assign n36741 = \pi0788  & ~n36740 ;
  assign n36742 = ~n36729 & ~n36741 ;
  assign n36743 = ~n36723 & n36742 ;
  assign n36744 = ~n23856 & n36666 ;
  assign n36745 = ~n36743 & n36744 ;
  assign n36746 = ~n36667 & ~n36745 ;
  assign n36747 = n30987 & ~n36659 ;
  assign n36748 = n23312 & n36747 ;
  assign n36749 = \pi1157  & ~n36647 ;
  assign n36750 = ~n36645 & n36749 ;
  assign n36751 = ~\pi1157  & ~n36652 ;
  assign n36752 = ~n36650 & n36751 ;
  assign n36753 = ~n36750 & ~n36752 ;
  assign n36754 = \pi0787  & ~n36753 ;
  assign n36755 = n26333 & ~n36632 ;
  assign n36756 = ~\pi0787  & ~n36755 ;
  assign n36757 = ~\pi1160  & ~n36756 ;
  assign n36758 = n23312 & n36757 ;
  assign n36759 = ~n36754 & n36758 ;
  assign n36760 = ~n36748 & ~n36759 ;
  assign n36761 = ~n23414 & n36601 ;
  assign n36762 = ~n24886 & n36761 ;
  assign n36763 = ~n23313 & ~n36762 ;
  assign n36764 = \pi1160  & ~n36756 ;
  assign n36765 = ~n36754 & n36764 ;
  assign n36766 = n31010 & ~n36659 ;
  assign n36767 = ~n36762 & ~n36766 ;
  assign n36768 = ~n36765 & n36767 ;
  assign n36769 = ~n36763 & ~n36768 ;
  assign n36770 = n36760 & ~n36769 ;
  assign n36771 = \pi0790  & ~n36770 ;
  assign n36772 = \pi0832  & ~n36771 ;
  assign n36773 = n36746 & n36772 ;
  assign n36774 = \pi0185  & ~\pi0832  ;
  assign n36775 = ~n21132 & ~n36774 ;
  assign n36776 = ~n36773 & n36775 ;
  assign n36777 = n9948 & ~n36773 ;
  assign n36778 = ~n36776 & ~n36777 ;
  assign n36779 = \pi0038  & n36599 ;
  assign n36780 = n8413 & n36779 ;
  assign n36781 = n1354 & n36780 ;
  assign n36782 = n1358 & n36781 ;
  assign n36783 = \pi0038  & ~\pi0185  ;
  assign n36784 = ~n21757 & n36783 ;
  assign n36785 = ~n36782 & ~n36784 ;
  assign n36786 = ~\pi0185  & \pi0751  ;
  assign n36787 = n21743 & n36786 ;
  assign n36788 = ~n21734 & n36787 ;
  assign n36789 = ~\pi0038  & n36788 ;
  assign n36790 = \pi0185  & ~n25023 ;
  assign n36791 = ~\pi0185  & ~n21467 ;
  assign n36792 = ~\pi0751  & ~n36791 ;
  assign n36793 = ~n36790 & n36792 ;
  assign n36794 = ~\pi0039  & ~\pi0185  ;
  assign n36795 = n21272 & n36794 ;
  assign n36796 = ~\pi0038  & ~n36795 ;
  assign n36797 = n36793 & n36796 ;
  assign n36798 = ~n36789 & ~n36797 ;
  assign n36799 = n36785 & n36798 ;
  assign n36800 = \pi0701  & ~n36799 ;
  assign n36801 = ~\pi0185  & ~\pi0778  ;
  assign n36802 = ~n23622 & ~n36801 ;
  assign n36803 = n36800 & ~n36802 ;
  assign n36804 = ~\pi0185  & n23548 ;
  assign n36805 = ~\pi0751  & ~n36804 ;
  assign n36806 = ~\pi0039  & ~\pi0751  ;
  assign n36807 = ~n22683 & n36806 ;
  assign n36808 = ~n36805 & ~n36807 ;
  assign n36809 = ~\pi0038  & n36808 ;
  assign n36810 = ~\pi0038  & \pi0185  ;
  assign n36811 = ~n26538 & n36810 ;
  assign n36812 = ~n36809 & ~n36811 ;
  assign n36813 = ~\pi0185  & ~n23567 ;
  assign n36814 = n23565 & n36813 ;
  assign n36815 = \pi0751  & n23575 ;
  assign n36816 = n23572 & n36815 ;
  assign n36817 = ~n36786 & ~n36816 ;
  assign n36818 = ~n36814 & ~n36817 ;
  assign n36819 = ~n36812 & ~n36818 ;
  assign n36820 = n6861 & n36819 ;
  assign n36821 = \pi0185  & \pi0603  ;
  assign n36822 = ~n20783 & n36821 ;
  assign n36823 = n36598 & n36822 ;
  assign n36824 = \pi0185  & \pi0680  ;
  assign n36825 = ~n20854 & n36824 ;
  assign n36826 = ~n20784 & n36825 ;
  assign n36827 = n1689 & n36826 ;
  assign n36828 = ~n36823 & ~n36827 ;
  assign n36829 = n26554 & ~n36828 ;
  assign n36830 = n1358 & n36829 ;
  assign n36831 = \pi0038  & ~n36830 ;
  assign n36832 = ~\pi0701  & ~n36831 ;
  assign n36833 = ~\pi0185  & ~\pi0701  ;
  assign n36834 = ~n26566 & n36833 ;
  assign n36835 = ~\pi0751  & n36833 ;
  assign n36836 = ~n22536 & n36835 ;
  assign n36837 = ~n36834 & ~n36836 ;
  assign n36838 = ~n36832 & n36837 ;
  assign n36839 = n6861 & n36838 ;
  assign n36840 = ~n36802 & ~n36839 ;
  assign n36841 = ~n36820 & n36840 ;
  assign n36842 = ~n36803 & ~n36841 ;
  assign n36843 = \pi0609  & ~n36842 ;
  assign n36844 = ~\pi0185  & ~\pi0625  ;
  assign n36845 = ~n22734 & ~n36844 ;
  assign n36846 = n36800 & ~n36845 ;
  assign n36847 = ~n36839 & ~n36845 ;
  assign n36848 = ~n36820 & n36847 ;
  assign n36849 = ~n36846 & ~n36848 ;
  assign n36850 = n6861 & n36785 ;
  assign n36851 = n36798 & n36850 ;
  assign n36852 = ~\pi0185  & \pi0625  ;
  assign n36853 = ~n22727 & ~n36852 ;
  assign n36854 = ~n36851 & ~n36853 ;
  assign n36855 = ~\pi1153  & ~n36854 ;
  assign n36856 = n36849 & n36855 ;
  assign n36857 = ~\pi0074  & ~\pi0701  ;
  assign n36858 = ~\pi0100  & n36857 ;
  assign n36859 = n1287 & n36858 ;
  assign n36860 = ~\pi0185  & ~n36859 ;
  assign n36861 = n21768 & n36860 ;
  assign n36862 = n21770 & n36860 ;
  assign n36863 = ~n21734 & n36862 ;
  assign n36864 = ~n36861 & ~n36863 ;
  assign n36865 = \pi0625  & ~n36864 ;
  assign n36866 = ~\pi0185  & ~n22017 ;
  assign n36867 = ~n21994 & n36866 ;
  assign n36868 = ~\pi0038  & ~\pi0185  ;
  assign n36869 = n6861 & ~n36868 ;
  assign n36870 = ~n22109 & n36869 ;
  assign n36871 = ~n36867 & ~n36870 ;
  assign n36872 = ~\pi0185  & ~n21757 ;
  assign n36873 = n22117 & ~n36872 ;
  assign n36874 = ~\pi0701  & ~n36873 ;
  assign n36875 = \pi0625  & n36874 ;
  assign n36876 = ~n36871 & n36875 ;
  assign n36877 = ~n36865 & ~n36876 ;
  assign n36878 = n21768 & n36844 ;
  assign n36879 = n21770 & n36844 ;
  assign n36880 = ~n21734 & n36879 ;
  assign n36881 = ~n36878 & ~n36880 ;
  assign n36882 = \pi1153  & n36881 ;
  assign n36883 = n36877 & n36882 ;
  assign n36884 = ~\pi0608  & ~n36883 ;
  assign n36885 = ~n36856 & n36884 ;
  assign n36886 = n36800 & ~n36853 ;
  assign n36887 = ~n36839 & ~n36853 ;
  assign n36888 = ~n36820 & n36887 ;
  assign n36889 = ~n36886 & ~n36888 ;
  assign n36890 = ~n36845 & ~n36851 ;
  assign n36891 = \pi1153  & ~n36890 ;
  assign n36892 = n36889 & n36891 ;
  assign n36893 = ~\pi0625  & ~n36864 ;
  assign n36894 = ~\pi0625  & n36874 ;
  assign n36895 = ~n36871 & n36894 ;
  assign n36896 = ~n36893 & ~n36895 ;
  assign n36897 = n21768 & n36852 ;
  assign n36898 = n21770 & n36852 ;
  assign n36899 = ~n21734 & n36898 ;
  assign n36900 = ~n36897 & ~n36899 ;
  assign n36901 = ~\pi1153  & n36900 ;
  assign n36902 = n36896 & n36901 ;
  assign n36903 = \pi0608  & ~n36902 ;
  assign n36904 = ~n36892 & n36903 ;
  assign n36905 = ~n36885 & ~n36904 ;
  assign n36906 = n23638 & ~n36905 ;
  assign n36907 = ~n36843 & ~n36906 ;
  assign n36908 = ~\pi0185  & n21768 ;
  assign n36909 = ~\pi0185  & n21770 ;
  assign n36910 = ~n21734 & n36909 ;
  assign n36911 = ~n36908 & ~n36910 ;
  assign n36912 = n26653 & n36911 ;
  assign n36913 = n26645 & n36785 ;
  assign n36914 = n36798 & n36913 ;
  assign n36915 = \pi0185  & ~n6861 ;
  assign n36916 = ~n20985 & n36915 ;
  assign n36917 = ~\pi0660  & ~n36916 ;
  assign n36918 = ~n36914 & n36917 ;
  assign n36919 = ~n34035 & ~n36918 ;
  assign n36920 = ~n36912 & ~n36919 ;
  assign n36921 = ~n36871 & n36874 ;
  assign n36922 = ~\pi0778  & n36864 ;
  assign n36923 = ~n36921 & n36922 ;
  assign n36924 = ~\pi0609  & ~n36923 ;
  assign n36925 = \pi1155  & ~n36924 ;
  assign n36926 = ~n36883 & ~n36902 ;
  assign n36927 = n22722 & ~n36926 ;
  assign n36928 = ~n36925 & ~n36927 ;
  assign n36929 = ~n36920 & ~n36928 ;
  assign n36930 = n36907 & n36929 ;
  assign n36931 = \pi0778  & ~n36905 ;
  assign n36932 = ~n36914 & ~n36916 ;
  assign n36933 = n20999 & ~n36932 ;
  assign n36934 = ~n32768 & n36911 ;
  assign n36935 = ~n22787 & ~n36934 ;
  assign n36936 = ~n36933 & n36935 ;
  assign n36937 = \pi0785  & n36936 ;
  assign n36938 = \pi0778  & ~n36926 ;
  assign n36939 = \pi0609  & ~n36923 ;
  assign n36940 = \pi0785  & n36939 ;
  assign n36941 = ~n36938 & n36940 ;
  assign n36942 = ~n36937 & ~n36941 ;
  assign n36943 = n36842 & n36942 ;
  assign n36944 = ~n36931 & n36943 ;
  assign n36945 = \pi0660  & ~n36934 ;
  assign n36946 = ~n36933 & n36945 ;
  assign n36947 = ~n36920 & ~n36946 ;
  assign n36948 = \pi0609  & ~n36935 ;
  assign n36949 = n36923 & n36948 ;
  assign n36950 = \pi0778  & n36948 ;
  assign n36951 = ~n36926 & n36950 ;
  assign n36952 = ~n36949 & ~n36951 ;
  assign n36953 = ~n36947 & n36952 ;
  assign n36954 = ~n36944 & n36953 ;
  assign n36955 = ~n36930 & n36954 ;
  assign n36956 = ~\pi0785  & ~n36944 ;
  assign n36957 = n26700 & ~n36956 ;
  assign n36958 = ~n36955 & n36957 ;
  assign n36959 = ~\pi0185  & ~n20811 ;
  assign n36960 = n21768 & n36959 ;
  assign n36961 = n21770 & n36959 ;
  assign n36962 = ~n21734 & n36961 ;
  assign n36963 = ~n36960 & ~n36962 ;
  assign n36964 = n23456 & n36785 ;
  assign n36965 = n36798 & n36964 ;
  assign n36966 = ~n21777 & n36911 ;
  assign n36967 = n21777 & n36915 ;
  assign n36968 = n20811 & ~n36967 ;
  assign n36969 = ~n36966 & n36968 ;
  assign n36970 = ~n36965 & n36969 ;
  assign n36971 = n36963 & ~n36970 ;
  assign n36972 = n23424 & ~n36971 ;
  assign n36973 = ~\pi0781  & ~n36967 ;
  assign n36974 = ~n36966 & n36973 ;
  assign n36975 = ~n36965 & n36974 ;
  assign n36976 = ~n23423 & n36975 ;
  assign n36977 = n23423 & ~n36911 ;
  assign n36978 = ~n36976 & ~n36977 ;
  assign n36979 = ~n36972 & n36978 ;
  assign n36980 = ~n23880 & ~n36979 ;
  assign n36981 = n23880 & ~n36911 ;
  assign n36982 = n24691 & ~n36981 ;
  assign n36983 = ~n36980 & n36982 ;
  assign n36984 = n26065 & ~n36926 ;
  assign n36985 = n26739 & n36864 ;
  assign n36986 = ~n36921 & n36985 ;
  assign n36987 = ~n23885 & n36911 ;
  assign n36988 = \pi0628  & ~n36987 ;
  assign n36989 = ~n36986 & n36988 ;
  assign n36990 = ~n36984 & n36989 ;
  assign n36991 = ~\pi0185  & ~\pi0628  ;
  assign n36992 = n21768 & n36991 ;
  assign n36993 = n21770 & n36991 ;
  assign n36994 = ~n21734 & n36993 ;
  assign n36995 = ~n36992 & ~n36994 ;
  assign n36996 = \pi1156  & n36995 ;
  assign n36997 = ~\pi0629  & n36996 ;
  assign n36998 = ~n36990 & n36997 ;
  assign n36999 = ~\pi0628  & ~n36987 ;
  assign n37000 = ~n36986 & n36999 ;
  assign n37001 = ~n36984 & n37000 ;
  assign n37002 = ~\pi0185  & \pi0628  ;
  assign n37003 = n21768 & n37002 ;
  assign n37004 = n21770 & n37002 ;
  assign n37005 = ~n21734 & n37004 ;
  assign n37006 = ~n37003 & ~n37005 ;
  assign n37007 = ~\pi1156  & n37006 ;
  assign n37008 = \pi0629  & n37007 ;
  assign n37009 = ~n37001 & n37008 ;
  assign n37010 = ~n36998 & ~n37009 ;
  assign n37011 = ~n36983 & n37010 ;
  assign n37012 = \pi0792  & ~n37011 ;
  assign n37013 = n23380 & ~n36923 ;
  assign n37014 = ~\pi0185  & ~n23380 ;
  assign n37015 = n21768 & n37014 ;
  assign n37016 = n21770 & n37014 ;
  assign n37017 = ~n21734 & n37016 ;
  assign n37018 = ~n37015 & ~n37017 ;
  assign n37019 = n21050 & n37018 ;
  assign n37020 = ~n37013 & n37019 ;
  assign n37021 = \pi0778  & n37019 ;
  assign n37022 = ~n36926 & n37021 ;
  assign n37023 = ~n37020 & ~n37022 ;
  assign n37024 = n23683 & ~n36971 ;
  assign n37025 = n21032 & n36975 ;
  assign n37026 = ~n21032 & ~n36911 ;
  assign n37027 = ~n20876 & ~n37026 ;
  assign n37028 = ~n37025 & n37027 ;
  assign n37029 = ~n37024 & n37028 ;
  assign n37030 = n37023 & ~n37029 ;
  assign n37031 = \pi0789  & ~n37030 ;
  assign n37032 = n22155 & n36963 ;
  assign n37033 = ~n36970 & n37032 ;
  assign n37034 = ~n21034 & n37033 ;
  assign n37035 = ~n22147 & ~n36923 ;
  assign n37036 = ~n36938 & n37035 ;
  assign n37037 = n22147 & ~n36911 ;
  assign n37038 = n24348 & ~n37037 ;
  assign n37039 = ~n21034 & n37038 ;
  assign n37040 = ~n37036 & n37039 ;
  assign n37041 = ~n37034 & ~n37040 ;
  assign n37042 = ~n21038 & n37041 ;
  assign n37043 = ~n37031 & n37042 ;
  assign n37044 = ~n37012 & n37043 ;
  assign n37045 = ~n36958 & n37044 ;
  assign n37046 = ~n22160 & n37018 ;
  assign n37047 = ~n37013 & n37046 ;
  assign n37048 = \pi0778  & n37046 ;
  assign n37049 = ~n36926 & n37048 ;
  assign n37050 = ~n37047 & ~n37049 ;
  assign n37051 = n22160 & n36911 ;
  assign n37052 = n20951 & ~n37051 ;
  assign n37053 = n37050 & n37052 ;
  assign n37054 = ~\pi0626  & ~n36977 ;
  assign n37055 = ~n36976 & n37054 ;
  assign n37056 = ~n36972 & n37055 ;
  assign n37057 = \pi0626  & n36911 ;
  assign n37058 = n20882 & ~n37057 ;
  assign n37059 = ~n37056 & n37058 ;
  assign n37060 = ~n37053 & ~n37059 ;
  assign n37061 = \pi0626  & ~n36977 ;
  assign n37062 = ~n36976 & n37061 ;
  assign n37063 = ~n36972 & n37062 ;
  assign n37064 = ~\pi0626  & n36911 ;
  assign n37065 = n20881 & ~n37064 ;
  assign n37066 = ~n37063 & n37065 ;
  assign n37067 = ~n23856 & ~n37066 ;
  assign n37068 = n37060 & n37067 ;
  assign n37069 = ~n26803 & ~n37068 ;
  assign n37070 = ~n37012 & n37069 ;
  assign n37071 = ~n21067 & ~n37070 ;
  assign n37072 = ~n37045 & n37071 ;
  assign n37073 = ~\pi0185  & \pi0644  ;
  assign n37074 = n21768 & n37073 ;
  assign n37075 = n21770 & n37073 ;
  assign n37076 = ~n21734 & n37075 ;
  assign n37077 = ~n37074 & ~n37076 ;
  assign n37078 = \pi0715  & n37077 ;
  assign n37079 = ~\pi0185  & ~n31367 ;
  assign n37080 = n21768 & n37079 ;
  assign n37081 = n21770 & n37079 ;
  assign n37082 = ~n21734 & n37081 ;
  assign n37083 = ~n37080 & ~n37082 ;
  assign n37084 = ~\pi0644  & ~n37083 ;
  assign n37085 = n34208 & ~n36979 ;
  assign n37086 = ~n37084 & ~n37085 ;
  assign n37087 = n37078 & n37086 ;
  assign n37088 = n31378 & ~n37087 ;
  assign n37089 = ~\pi0715  & n37083 ;
  assign n37090 = ~n23958 & ~n37089 ;
  assign n37091 = n31382 & ~n36979 ;
  assign n37092 = ~n37090 & ~n37091 ;
  assign n37093 = n26824 & ~n37092 ;
  assign n37094 = \pi0790  & ~n37093 ;
  assign n37095 = ~n37088 & n37094 ;
  assign n37096 = ~n36986 & ~n36987 ;
  assign n37097 = ~n36984 & n37096 ;
  assign n37098 = ~\pi0792  & ~n37097 ;
  assign n37099 = ~\pi0647  & ~n37098 ;
  assign n37100 = n21768 & n36651 ;
  assign n37101 = n21770 & n36651 ;
  assign n37102 = ~n21734 & n37101 ;
  assign n37103 = ~n37100 & ~n37102 ;
  assign n37104 = ~\pi1157  & n37103 ;
  assign n37105 = ~n37099 & n37104 ;
  assign n37106 = ~n36990 & n36996 ;
  assign n37107 = ~n37001 & n37007 ;
  assign n37108 = ~n37106 & ~n37107 ;
  assign n37109 = \pi0792  & n37104 ;
  assign n37110 = ~n37108 & n37109 ;
  assign n37111 = ~n37105 & ~n37110 ;
  assign n37112 = ~n20846 & n36981 ;
  assign n37113 = n30376 & ~n36979 ;
  assign n37114 = ~n37112 & ~n37113 ;
  assign n37115 = ~n34703 & n36660 ;
  assign n37116 = ~n20910 & ~n37115 ;
  assign n37117 = n37114 & n37116 ;
  assign n37118 = \pi0630  & ~n37117 ;
  assign n37119 = n37111 & n37118 ;
  assign n37120 = \pi0647  & ~n37098 ;
  assign n37121 = n21768 & n36646 ;
  assign n37122 = n21770 & n36646 ;
  assign n37123 = ~n21734 & n37122 ;
  assign n37124 = ~n37121 & ~n37123 ;
  assign n37125 = \pi1157  & n37124 ;
  assign n37126 = ~n37120 & n37125 ;
  assign n37127 = \pi0792  & n37125 ;
  assign n37128 = ~n37108 & n37127 ;
  assign n37129 = ~n37126 & ~n37128 ;
  assign n37130 = ~\pi0630  & ~n37117 ;
  assign n37131 = n37129 & n37130 ;
  assign n37132 = ~n37119 & ~n37131 ;
  assign n37133 = \pi0787  & n37132 ;
  assign n37134 = ~n37095 & ~n37133 ;
  assign n37135 = ~n37072 & n37134 ;
  assign n37136 = ~\pi0787  & n37098 ;
  assign n37137 = n33084 & ~n37108 ;
  assign n37138 = ~n37136 & ~n37137 ;
  assign n37139 = ~\pi0644  & n37138 ;
  assign n37140 = \pi0715  & ~n37139 ;
  assign n37141 = n37111 & n37129 ;
  assign n37142 = n26918 & ~n37141 ;
  assign n37143 = ~n37140 & ~n37142 ;
  assign n37144 = ~\pi0185  & ~\pi0644  ;
  assign n37145 = n21768 & n37144 ;
  assign n37146 = n21770 & n37144 ;
  assign n37147 = ~n21734 & n37146 ;
  assign n37148 = ~n37145 & ~n37147 ;
  assign n37149 = n37092 & n37148 ;
  assign n37150 = \pi1160  & ~n37149 ;
  assign n37151 = n37143 & n37150 ;
  assign n37152 = \pi0644  & n37138 ;
  assign n37153 = ~\pi0715  & ~n37152 ;
  assign n37154 = n33098 & ~n37141 ;
  assign n37155 = ~n37153 & ~n37154 ;
  assign n37156 = ~\pi1160  & ~n37087 ;
  assign n37157 = n37155 & n37156 ;
  assign n37158 = ~n37151 & ~n37157 ;
  assign n37159 = \pi0790  & ~n37158 ;
  assign n37160 = ~n36776 & ~n37159 ;
  assign n37161 = ~n37135 & n37160 ;
  assign n37162 = ~n36778 & ~n37161 ;
  assign n37163 = ~\pi0186  & ~n1689 ;
  assign n37164 = ~n21032 & ~n37163 ;
  assign n37165 = \pi0789  & n37164 ;
  assign n37166 = ~n23880 & ~n37165 ;
  assign n37167 = n23423 & n37166 ;
  assign n37168 = ~\pi0752  & n1689 ;
  assign n37169 = n20784 & n37168 ;
  assign n37170 = ~n37163 & ~n37169 ;
  assign n37171 = n20794 & ~n37170 ;
  assign n37172 = n20796 & ~n37171 ;
  assign n37173 = n20799 & ~n37170 ;
  assign n37174 = n20801 & ~n37173 ;
  assign n37175 = ~n37172 & ~n37174 ;
  assign n37176 = ~\pi0785  & ~n37163 ;
  assign n37177 = ~n37169 & n37176 ;
  assign n37178 = ~n20804 & ~n37177 ;
  assign n37179 = ~n20812 & n37178 ;
  assign n37180 = n37166 & n37179 ;
  assign n37181 = n37175 & n37180 ;
  assign n37182 = ~n37167 & ~n37181 ;
  assign n37183 = ~\pi0186  & \pi0792  ;
  assign n37184 = ~n1689 & n37183 ;
  assign n37185 = ~n20845 & n37184 ;
  assign n37186 = ~n20910 & ~n37185 ;
  assign n37187 = ~\pi0186  & \pi0788  ;
  assign n37188 = ~n1689 & n37187 ;
  assign n37189 = ~n20778 & n37188 ;
  assign n37190 = n37186 & ~n37189 ;
  assign n37191 = n37182 & n37190 ;
  assign n37192 = n20846 & n37186 ;
  assign n37193 = \pi0703  & n1689 ;
  assign n37194 = n20855 & n37193 ;
  assign n37195 = ~n20861 & n37194 ;
  assign n37196 = ~n37163 & ~n37195 ;
  assign n37197 = n20879 & ~n37196 ;
  assign n37198 = n20895 & n37197 ;
  assign n37199 = ~\pi0186  & \pi0647  ;
  assign n37200 = ~n1689 & n37199 ;
  assign n37201 = n20897 & ~n37200 ;
  assign n37202 = ~n37198 & n37201 ;
  assign n37203 = ~\pi0186  & ~\pi0647  ;
  assign n37204 = ~n1689 & n37203 ;
  assign n37205 = n20849 & ~n37204 ;
  assign n37206 = ~n24761 & ~n37205 ;
  assign n37207 = n31479 & n37197 ;
  assign n37208 = ~n37206 & ~n37207 ;
  assign n37209 = ~n37202 & ~n37208 ;
  assign n37210 = ~n37192 & n37209 ;
  assign n37211 = ~n37191 & n37210 ;
  assign n37212 = ~n29722 & ~n37211 ;
  assign n37213 = n20938 & n37197 ;
  assign n37214 = \pi0629  & ~n37189 ;
  assign n37215 = ~n37213 & n37214 ;
  assign n37216 = n37182 & n37215 ;
  assign n37217 = n21077 & n37197 ;
  assign n37218 = ~\pi0629  & ~n37189 ;
  assign n37219 = ~n37217 & n37218 ;
  assign n37220 = n37182 & n37219 ;
  assign n37221 = n29714 & ~n37213 ;
  assign n37222 = n29709 & ~n37217 ;
  assign n37223 = \pi0792  & ~n37222 ;
  assign n37224 = ~n37221 & n37223 ;
  assign n37225 = ~n37220 & n37224 ;
  assign n37226 = ~n37216 & n37225 ;
  assign n37227 = ~n21067 & ~n37226 ;
  assign n37228 = n23423 & ~n37165 ;
  assign n37229 = ~n37165 & n37179 ;
  assign n37230 = n37175 & n37229 ;
  assign n37231 = ~n37228 & ~n37230 ;
  assign n37232 = ~\pi0626  & n37231 ;
  assign n37233 = \pi0626  & ~n37163 ;
  assign n37234 = n20882 & ~n37233 ;
  assign n37235 = ~n37232 & n37234 ;
  assign n37236 = n23170 & ~n37196 ;
  assign n37237 = ~\pi0626  & ~n37163 ;
  assign n37238 = n20881 & ~n37237 ;
  assign n37239 = ~n37236 & ~n37238 ;
  assign n37240 = \pi0626  & ~n37236 ;
  assign n37241 = n37231 & n37240 ;
  assign n37242 = ~n37239 & ~n37241 ;
  assign n37243 = ~n37235 & ~n37242 ;
  assign n37244 = \pi0788  & ~n37243 ;
  assign n37245 = ~n23856 & n37244 ;
  assign n37246 = n20964 & n37178 ;
  assign n37247 = n37175 & n37246 ;
  assign n37248 = \pi0627  & ~n37163 ;
  assign n37249 = ~n37195 & n37248 ;
  assign n37250 = ~n20968 & ~n37249 ;
  assign n37251 = ~n37247 & ~n37250 ;
  assign n37252 = n20974 & n37178 ;
  assign n37253 = n37175 & n37252 ;
  assign n37254 = ~\pi0627  & ~n37163 ;
  assign n37255 = ~n37195 & n37254 ;
  assign n37256 = ~n20978 & ~n37255 ;
  assign n37257 = ~n37253 & ~n37256 ;
  assign n37258 = ~n37251 & ~n37257 ;
  assign n37259 = \pi0781  & n37258 ;
  assign n37260 = \pi0680  & \pi0703  ;
  assign n37261 = ~n20854 & n37260 ;
  assign n37262 = ~n20861 & n37261 ;
  assign n37263 = ~n20986 & n37262 ;
  assign n37264 = \pi0603  & ~\pi0752  ;
  assign n37265 = ~n20783 & n37264 ;
  assign n37266 = ~n20985 & n37265 ;
  assign n37267 = ~n37163 & ~n37266 ;
  assign n37268 = ~n37263 & n37267 ;
  assign n37269 = \pi0186  & ~n1689 ;
  assign n37270 = ~\pi0609  & ~n37269 ;
  assign n37271 = ~n37268 & n37270 ;
  assign n37272 = ~\pi1155  & ~n37163 ;
  assign n37273 = ~n37195 & n37272 ;
  assign n37274 = ~n20999 & ~n37273 ;
  assign n37275 = ~n37271 & ~n37274 ;
  assign n37276 = \pi1155  & ~n37173 ;
  assign n37277 = ~\pi0660  & ~n37276 ;
  assign n37278 = ~n37275 & n37277 ;
  assign n37279 = ~n21007 & ~n37172 ;
  assign n37280 = \pi0609  & ~n37269 ;
  assign n37281 = ~n37268 & n37280 ;
  assign n37282 = \pi1155  & ~n37163 ;
  assign n37283 = ~n37195 & n37282 ;
  assign n37284 = ~n21774 & ~n37283 ;
  assign n37285 = \pi0785  & ~n37284 ;
  assign n37286 = ~n37281 & n37285 ;
  assign n37287 = n37279 & ~n37286 ;
  assign n37288 = ~n37278 & ~n37287 ;
  assign n37289 = ~n37268 & ~n37269 ;
  assign n37290 = ~\pi0785  & ~n37289 ;
  assign n37291 = n21022 & ~n37290 ;
  assign n37292 = ~n37288 & n37291 ;
  assign n37293 = ~n21034 & ~n37292 ;
  assign n37294 = ~n37259 & n37293 ;
  assign n37295 = ~n20876 & n37164 ;
  assign n37296 = ~n24969 & ~n37295 ;
  assign n37297 = n37179 & ~n37295 ;
  assign n37298 = n37175 & n37297 ;
  assign n37299 = ~n37296 & ~n37298 ;
  assign n37300 = n21050 & ~n37163 ;
  assign n37301 = ~n37195 & n37300 ;
  assign n37302 = ~n21051 & ~n37301 ;
  assign n37303 = ~n21038 & n37302 ;
  assign n37304 = ~n37299 & n37303 ;
  assign n37305 = ~n23177 & ~n37304 ;
  assign n37306 = ~n23856 & ~n37305 ;
  assign n37307 = ~n37294 & n37306 ;
  assign n37308 = ~n37245 & ~n37307 ;
  assign n37309 = n37227 & n37308 ;
  assign n37310 = ~n37212 & ~n37309 ;
  assign n37311 = n24830 & n37197 ;
  assign n37312 = \pi1157  & ~n37204 ;
  assign n37313 = ~n37311 & n37312 ;
  assign n37314 = ~\pi1157  & ~n37200 ;
  assign n37315 = ~n37198 & n37314 ;
  assign n37316 = ~n37313 & ~n37315 ;
  assign n37317 = \pi0787  & ~n37316 ;
  assign n37318 = n24844 & n37197 ;
  assign n37319 = ~n24843 & ~n37318 ;
  assign n37320 = ~n37317 & ~n37319 ;
  assign n37321 = n37182 & ~n37189 ;
  assign n37322 = n31580 & ~n37321 ;
  assign n37323 = ~n37320 & ~n37322 ;
  assign n37324 = n23313 & ~n37323 ;
  assign n37325 = \pi0790  & n37324 ;
  assign n37326 = n31588 & ~n37321 ;
  assign n37327 = ~n23414 & n37163 ;
  assign n37328 = ~n24886 & n37327 ;
  assign n37329 = n20891 & n37197 ;
  assign n37330 = ~\pi0787  & ~n37329 ;
  assign n37331 = ~\pi1160  & ~n37330 ;
  assign n37332 = ~n37317 & n37331 ;
  assign n37333 = ~n37328 & ~n37332 ;
  assign n37334 = ~n37326 & n37333 ;
  assign n37335 = ~n23312 & ~n37328 ;
  assign n37336 = \pi0790  & ~n37335 ;
  assign n37337 = ~n37334 & n37336 ;
  assign n37338 = ~n37325 & ~n37337 ;
  assign n37339 = \pi0832  & n37338 ;
  assign n37340 = ~n37310 & n37339 ;
  assign n37341 = \pi0186  & ~\pi0832  ;
  assign n37342 = ~n21132 & ~n37341 ;
  assign n37343 = ~n37340 & n37342 ;
  assign n37344 = \pi0186  & ~n25024 ;
  assign n37345 = ~\pi0186  & ~\pi0752  ;
  assign n37346 = ~n25033 & n37345 ;
  assign n37347 = ~n25028 & n37346 ;
  assign n37348 = ~n37344 & ~n37347 ;
  assign n37349 = n25041 & ~n37348 ;
  assign n37350 = \pi0186  & ~n6861 ;
  assign n37351 = ~\pi0186  & n22124 ;
  assign n37352 = ~\pi0186  & n21770 ;
  assign n37353 = ~n21734 & n37352 ;
  assign n37354 = ~n37351 & ~n37353 ;
  assign n37355 = \pi0752  & n1289 ;
  assign n37356 = n1287 & n37355 ;
  assign n37357 = n37354 & n37356 ;
  assign n37358 = ~n37350 & ~n37357 ;
  assign n37359 = ~n37349 & n37358 ;
  assign n37360 = n21777 & ~n37359 ;
  assign n37361 = ~\pi0186  & n21768 ;
  assign n37362 = ~n37353 & ~n37361 ;
  assign n37363 = ~n21777 & n37362 ;
  assign n37364 = ~\pi0781  & ~n37363 ;
  assign n37365 = ~n37360 & n37364 ;
  assign n37366 = \pi0619  & n37365 ;
  assign n37367 = ~\pi0618  & ~n37363 ;
  assign n37368 = ~\pi0186  & \pi0618  ;
  assign n37369 = n21768 & n37368 ;
  assign n37370 = n21770 & n37368 ;
  assign n37371 = ~n21734 & n37370 ;
  assign n37372 = ~n37369 & ~n37371 ;
  assign n37373 = ~\pi1154  & n37372 ;
  assign n37374 = ~n37367 & n37373 ;
  assign n37375 = n21777 & n37373 ;
  assign n37376 = ~n37359 & n37375 ;
  assign n37377 = ~n37374 & ~n37376 ;
  assign n37378 = \pi0781  & n37377 ;
  assign n37379 = \pi0618  & ~n37363 ;
  assign n37380 = ~\pi0186  & ~\pi0618  ;
  assign n37381 = n21768 & n37380 ;
  assign n37382 = n21770 & n37380 ;
  assign n37383 = ~n21734 & n37382 ;
  assign n37384 = ~n37381 & ~n37383 ;
  assign n37385 = \pi1154  & n37384 ;
  assign n37386 = ~n37379 & n37385 ;
  assign n37387 = n21777 & n37385 ;
  assign n37388 = ~n37359 & n37387 ;
  assign n37389 = ~n37386 & ~n37388 ;
  assign n37390 = \pi0619  & n37389 ;
  assign n37391 = n37378 & n37390 ;
  assign n37392 = ~n37366 & ~n37391 ;
  assign n37393 = ~\pi0186  & ~\pi0619  ;
  assign n37394 = n21768 & n37393 ;
  assign n37395 = n21770 & n37393 ;
  assign n37396 = ~n21734 & n37395 ;
  assign n37397 = ~n37394 & ~n37396 ;
  assign n37398 = \pi1159  & n37397 ;
  assign n37399 = n37392 & n37398 ;
  assign n37400 = \pi0789  & ~n37399 ;
  assign n37401 = ~\pi0619  & n37365 ;
  assign n37402 = ~\pi0619  & n37389 ;
  assign n37403 = n37378 & n37402 ;
  assign n37404 = ~n37401 & ~n37403 ;
  assign n37405 = ~\pi0186  & \pi0619  ;
  assign n37406 = n21768 & n37405 ;
  assign n37407 = n21770 & n37405 ;
  assign n37408 = ~n21734 & n37407 ;
  assign n37409 = ~n37406 & ~n37408 ;
  assign n37410 = ~\pi1159  & n37409 ;
  assign n37411 = n37404 & n37410 ;
  assign n37412 = ~n23880 & ~n37411 ;
  assign n37413 = n37400 & n37412 ;
  assign n37414 = ~\pi0789  & n37364 ;
  assign n37415 = ~n37360 & n37414 ;
  assign n37416 = ~\pi0789  & n37389 ;
  assign n37417 = n37378 & n37416 ;
  assign n37418 = ~n37415 & ~n37417 ;
  assign n37419 = ~n23880 & ~n37418 ;
  assign n37420 = n23880 & ~n37362 ;
  assign n37421 = n21092 & ~n37420 ;
  assign n37422 = ~n37419 & n37421 ;
  assign n37423 = ~n37413 & n37422 ;
  assign n37424 = ~n21092 & n37362 ;
  assign n37425 = \pi0644  & ~n37424 ;
  assign n37426 = ~n37423 & n37425 ;
  assign n37427 = ~\pi0186  & ~\pi0644  ;
  assign n37428 = n21768 & n37427 ;
  assign n37429 = n21770 & n37427 ;
  assign n37430 = ~n21734 & n37429 ;
  assign n37431 = ~n37428 & ~n37430 ;
  assign n37432 = n23412 & n37431 ;
  assign n37433 = ~n37426 & n37432 ;
  assign n37434 = ~\pi0644  & ~n37424 ;
  assign n37435 = ~n37423 & n37434 ;
  assign n37436 = ~\pi0186  & \pi0644  ;
  assign n37437 = n21768 & n37436 ;
  assign n37438 = n21770 & n37436 ;
  assign n37439 = ~n21734 & n37438 ;
  assign n37440 = ~n37437 & ~n37439 ;
  assign n37441 = n23413 & n37440 ;
  assign n37442 = ~n37435 & n37441 ;
  assign n37443 = ~n37433 & ~n37442 ;
  assign n37444 = \pi0790  & ~n37443 ;
  assign n37445 = ~\pi0186  & ~\pi0625  ;
  assign n37446 = ~n22734 & ~n37445 ;
  assign n37447 = ~\pi0186  & \pi0625  ;
  assign n37448 = n21768 & n37447 ;
  assign n37449 = n21770 & n37447 ;
  assign n37450 = ~n21734 & n37449 ;
  assign n37451 = ~n37448 & ~n37450 ;
  assign n37452 = ~\pi1153  & n37451 ;
  assign n37453 = n37446 & n37452 ;
  assign n37454 = ~\pi0703  & ~n37354 ;
  assign n37455 = n6861 & ~n37454 ;
  assign n37456 = ~\pi0186  & ~n22017 ;
  assign n37457 = ~n21994 & n37456 ;
  assign n37458 = ~\pi0038  & ~\pi0186  ;
  assign n37459 = ~n22109 & ~n37458 ;
  assign n37460 = ~n37457 & ~n37459 ;
  assign n37461 = ~\pi0186  & ~n21757 ;
  assign n37462 = n22117 & ~n37461 ;
  assign n37463 = \pi0703  & ~n37462 ;
  assign n37464 = ~n37460 & n37463 ;
  assign n37465 = n37452 & ~n37464 ;
  assign n37466 = n37455 & n37465 ;
  assign n37467 = ~n37453 & ~n37466 ;
  assign n37468 = ~n22727 & ~n37447 ;
  assign n37469 = n21768 & n37445 ;
  assign n37470 = n21770 & n37445 ;
  assign n37471 = ~n21734 & n37470 ;
  assign n37472 = ~n37469 & ~n37471 ;
  assign n37473 = \pi1153  & n37472 ;
  assign n37474 = n37468 & n37473 ;
  assign n37475 = ~n37464 & n37473 ;
  assign n37476 = n37455 & n37475 ;
  assign n37477 = ~n37474 & ~n37476 ;
  assign n37478 = n37467 & n37477 ;
  assign n37479 = n22148 & ~n37478 ;
  assign n37480 = ~\pi0778  & n37350 ;
  assign n37481 = ~\pi0778  & ~n37464 ;
  assign n37482 = n37455 & n37481 ;
  assign n37483 = ~n37480 & ~n37482 ;
  assign n37484 = ~n22147 & ~n37483 ;
  assign n37485 = n22147 & n37362 ;
  assign n37486 = ~n22155 & ~n37485 ;
  assign n37487 = ~n37484 & n37486 ;
  assign n37488 = ~n37479 & n37487 ;
  assign n37489 = n22155 & ~n37362 ;
  assign n37490 = n22162 & ~n37489 ;
  assign n37491 = ~n37488 & n37490 ;
  assign n37492 = ~n22162 & n37362 ;
  assign n37493 = ~\pi0647  & ~n37492 ;
  assign n37494 = ~n37491 & n37493 ;
  assign n37495 = ~n22913 & ~n37494 ;
  assign n37496 = n21768 & n37199 ;
  assign n37497 = n21770 & n37199 ;
  assign n37498 = ~n21734 & n37497 ;
  assign n37499 = ~n37496 & ~n37498 ;
  assign n37500 = ~\pi1157  & n37499 ;
  assign n37501 = n37495 & n37500 ;
  assign n37502 = \pi0628  & ~n37492 ;
  assign n37503 = ~n37491 & n37502 ;
  assign n37504 = ~\pi0186  & ~\pi0628  ;
  assign n37505 = n21768 & n37504 ;
  assign n37506 = n21770 & n37504 ;
  assign n37507 = ~n21734 & n37506 ;
  assign n37508 = ~n37505 & ~n37507 ;
  assign n37509 = \pi1156  & n37508 ;
  assign n37510 = ~n37503 & n37509 ;
  assign n37511 = ~\pi0628  & ~n37492 ;
  assign n37512 = ~n37491 & n37511 ;
  assign n37513 = ~\pi0186  & \pi0628  ;
  assign n37514 = n21768 & n37513 ;
  assign n37515 = n21770 & n37513 ;
  assign n37516 = ~n21734 & n37515 ;
  assign n37517 = ~n37514 & ~n37516 ;
  assign n37518 = ~\pi1156  & n37517 ;
  assign n37519 = ~n37512 & n37518 ;
  assign n37520 = ~n37510 & ~n37519 ;
  assign n37521 = \pi0792  & n37500 ;
  assign n37522 = ~n37520 & n37521 ;
  assign n37523 = ~n37501 & ~n37522 ;
  assign n37524 = \pi0647  & ~n37492 ;
  assign n37525 = ~n37491 & n37524 ;
  assign n37526 = ~n22956 & ~n37525 ;
  assign n37527 = n21768 & n37203 ;
  assign n37528 = n21770 & n37203 ;
  assign n37529 = ~n21734 & n37528 ;
  assign n37530 = ~n37527 & ~n37529 ;
  assign n37531 = \pi1157  & n37530 ;
  assign n37532 = n37526 & n37531 ;
  assign n37533 = \pi0792  & n37531 ;
  assign n37534 = ~n37520 & n37533 ;
  assign n37535 = ~n37532 & ~n37534 ;
  assign n37536 = n37523 & n37535 ;
  assign n37537 = \pi0787  & n37536 ;
  assign n37538 = ~\pi0787  & ~n37492 ;
  assign n37539 = ~n37491 & n37538 ;
  assign n37540 = ~n33084 & ~n37539 ;
  assign n37541 = n23518 & n37540 ;
  assign n37542 = \pi0792  & n23518 ;
  assign n37543 = ~n37520 & n37542 ;
  assign n37544 = ~n37541 & ~n37543 ;
  assign n37545 = \pi0790  & ~n37544 ;
  assign n37546 = ~n37537 & n37545 ;
  assign n37547 = ~n37444 & ~n37546 ;
  assign n37548 = n9948 & n37547 ;
  assign n37549 = n24691 & ~n37420 ;
  assign n37550 = ~n37419 & n37549 ;
  assign n37551 = ~n37413 & n37550 ;
  assign n37552 = ~\pi0629  & n37509 ;
  assign n37553 = ~n37503 & n37552 ;
  assign n37554 = \pi0629  & n37518 ;
  assign n37555 = ~n37512 & n37554 ;
  assign n37556 = ~n37553 & ~n37555 ;
  assign n37557 = ~n37551 & n37556 ;
  assign n37558 = n24724 & ~n37557 ;
  assign n37559 = \pi1159  & ~n37489 ;
  assign n37560 = ~n37488 & n37559 ;
  assign n37561 = \pi0648  & ~n20830 ;
  assign n37562 = ~n37560 & n37561 ;
  assign n37563 = ~n37411 & n37562 ;
  assign n37564 = ~\pi1159  & ~n37489 ;
  assign n37565 = ~n37488 & n37564 ;
  assign n37566 = ~\pi0648  & ~n22872 ;
  assign n37567 = ~n37565 & n37566 ;
  assign n37568 = ~n37399 & n37567 ;
  assign n37569 = ~n37563 & ~n37568 ;
  assign n37570 = \pi0789  & ~n37569 ;
  assign n37571 = ~\pi0618  & ~n37485 ;
  assign n37572 = ~n37484 & n37571 ;
  assign n37573 = ~n37479 & n37572 ;
  assign n37574 = \pi1154  & ~n37573 ;
  assign n37575 = \pi0627  & n37377 ;
  assign n37576 = ~n37574 & n37575 ;
  assign n37577 = \pi0618  & ~n37485 ;
  assign n37578 = ~n37484 & n37577 ;
  assign n37579 = ~n37479 & n37578 ;
  assign n37580 = ~\pi1154  & ~n37579 ;
  assign n37581 = ~\pi0627  & n37389 ;
  assign n37582 = ~n37580 & n37581 ;
  assign n37583 = ~n37576 & ~n37582 ;
  assign n37584 = n32123 & ~n37398 ;
  assign n37585 = n31279 & n37409 ;
  assign n37586 = ~n33522 & ~n37585 ;
  assign n37587 = ~n37584 & ~n37586 ;
  assign n37588 = \pi0781  & ~n37587 ;
  assign n37589 = ~n37583 & n37588 ;
  assign n37590 = ~n37570 & ~n37589 ;
  assign n37591 = ~n21038 & ~n37590 ;
  assign n37592 = \pi0038  & \pi0186  ;
  assign n37593 = ~n22708 & n37592 ;
  assign n37594 = ~\pi0038  & \pi0186  ;
  assign n37595 = ~n37593 & ~n37594 ;
  assign n37596 = ~n23558 & ~n37593 ;
  assign n37597 = n23557 & n37596 ;
  assign n37598 = ~n37595 & ~n37597 ;
  assign n37599 = ~\pi0186  & n23548 ;
  assign n37600 = ~n25191 & n37599 ;
  assign n37601 = ~n25190 & n37600 ;
  assign n37602 = \pi0703  & ~\pi0752  ;
  assign n37603 = ~n37601 & n37602 ;
  assign n37604 = ~n37598 & n37603 ;
  assign n37605 = ~\pi0186  & ~n25209 ;
  assign n37606 = ~n25204 & n37605 ;
  assign n37607 = n23575 & n37594 ;
  assign n37608 = n23572 & n37607 ;
  assign n37609 = ~n25217 & ~n37608 ;
  assign n37610 = ~n37606 & n37609 ;
  assign n37611 = \pi0703  & \pi0752  ;
  assign n37612 = ~n37610 & n37611 ;
  assign n37613 = ~n37604 & ~n37612 ;
  assign n37614 = \pi0752  & n37354 ;
  assign n37615 = ~\pi0703  & n25040 ;
  assign n37616 = ~\pi0703  & ~n37344 ;
  assign n37617 = ~n37347 & n37616 ;
  assign n37618 = ~n37615 & ~n37617 ;
  assign n37619 = ~n37614 & ~n37618 ;
  assign n37620 = n6861 & ~n37619 ;
  assign n37621 = n37613 & n37620 ;
  assign n37622 = ~n37468 & ~n37621 ;
  assign n37623 = ~n37357 & ~n37446 ;
  assign n37624 = ~n37349 & n37623 ;
  assign n37625 = \pi1153  & ~n37624 ;
  assign n37626 = ~n37622 & n37625 ;
  assign n37627 = \pi0608  & n37467 ;
  assign n37628 = ~n37626 & n37627 ;
  assign n37629 = ~n37446 & ~n37621 ;
  assign n37630 = ~n37357 & ~n37468 ;
  assign n37631 = ~n37349 & n37630 ;
  assign n37632 = ~\pi1153  & ~n37631 ;
  assign n37633 = ~n37629 & n37632 ;
  assign n37634 = ~\pi0608  & n37477 ;
  assign n37635 = ~n37633 & n37634 ;
  assign n37636 = ~n37628 & ~n37635 ;
  assign n37637 = n23613 & ~n37636 ;
  assign n37638 = \pi0778  & ~n37478 ;
  assign n37639 = \pi0609  & n37483 ;
  assign n37640 = ~n37638 & n37639 ;
  assign n37641 = ~\pi0186  & ~\pi0778  ;
  assign n37642 = ~n23622 & ~n37641 ;
  assign n37643 = ~\pi0609  & ~n37642 ;
  assign n37644 = ~n37621 & n37643 ;
  assign n37645 = ~\pi1155  & ~n37644 ;
  assign n37646 = ~n37640 & n37645 ;
  assign n37647 = ~n37637 & n37646 ;
  assign n37648 = ~n22788 & n37362 ;
  assign n37649 = ~\pi0660  & ~n37648 ;
  assign n37650 = ~n22787 & ~n37649 ;
  assign n37651 = ~n22787 & n22788 ;
  assign n37652 = ~n37359 & n37651 ;
  assign n37653 = ~n37650 & ~n37652 ;
  assign n37654 = ~n37647 & n37653 ;
  assign n37655 = ~n22767 & n37362 ;
  assign n37656 = \pi0660  & ~n37655 ;
  assign n37657 = ~n22766 & ~n37656 ;
  assign n37658 = n31822 & ~n37359 ;
  assign n37659 = ~n37657 & ~n37658 ;
  assign n37660 = \pi0785  & ~n37659 ;
  assign n37661 = ~\pi0609  & n37483 ;
  assign n37662 = \pi1155  & ~n37661 ;
  assign n37663 = n22722 & ~n37478 ;
  assign n37664 = ~n37662 & ~n37663 ;
  assign n37665 = \pi0609  & ~n37642 ;
  assign n37666 = ~n37621 & n37665 ;
  assign n37667 = \pi0785  & ~n37666 ;
  assign n37668 = ~n37664 & n37667 ;
  assign n37669 = ~n37660 & ~n37668 ;
  assign n37670 = n23638 & ~n37660 ;
  assign n37671 = ~n37636 & n37670 ;
  assign n37672 = ~n37669 & ~n37671 ;
  assign n37673 = ~n37654 & n37672 ;
  assign n37674 = n21019 & ~n37373 ;
  assign n37675 = n21020 & n37384 ;
  assign n37676 = ~n33630 & ~n37675 ;
  assign n37677 = ~n37674 & ~n37676 ;
  assign n37678 = ~n37621 & ~n37642 ;
  assign n37679 = ~\pi0785  & ~n37678 ;
  assign n37680 = ~n37587 & ~n37679 ;
  assign n37681 = \pi0778  & ~n37587 ;
  assign n37682 = ~n37636 & n37681 ;
  assign n37683 = ~n37680 & ~n37682 ;
  assign n37684 = ~n37677 & ~n37683 ;
  assign n37685 = ~n21038 & n37684 ;
  assign n37686 = ~n37673 & n37685 ;
  assign n37687 = ~n37591 & ~n37686 ;
  assign n37688 = n30606 & ~n37418 ;
  assign n37689 = n30606 & ~n37411 ;
  assign n37690 = n37400 & n37689 ;
  assign n37691 = ~n37688 & ~n37690 ;
  assign n37692 = ~n22849 & n37362 ;
  assign n37693 = \pi0641  & n37692 ;
  assign n37694 = ~n37484 & ~n37485 ;
  assign n37695 = ~n37479 & n37694 ;
  assign n37696 = n33656 & ~n37695 ;
  assign n37697 = ~n37693 & ~n37696 ;
  assign n37698 = ~\pi0641  & n37362 ;
  assign n37699 = n20776 & ~n37698 ;
  assign n37700 = n37697 & n37699 ;
  assign n37701 = ~\pi0641  & n37692 ;
  assign n37702 = n33649 & ~n37695 ;
  assign n37703 = ~n37701 & ~n37702 ;
  assign n37704 = \pi0641  & n37362 ;
  assign n37705 = n20777 & ~n37704 ;
  assign n37706 = n37703 & n37705 ;
  assign n37707 = ~n23856 & ~n37706 ;
  assign n37708 = ~n37700 & n37707 ;
  assign n37709 = n37691 & n37708 ;
  assign n37710 = ~n26803 & ~n37709 ;
  assign n37711 = ~n21067 & ~n37710 ;
  assign n37712 = n37687 & n37711 ;
  assign n37713 = ~n37558 & ~n37712 ;
  assign n37714 = ~n24761 & ~n37713 ;
  assign n37715 = \pi0630  & ~n37523 ;
  assign n37716 = ~\pi0630  & ~n37535 ;
  assign n37717 = n37400 & ~n37411 ;
  assign n37718 = n30376 & n37418 ;
  assign n37719 = ~n37717 & n37718 ;
  assign n37720 = ~n30376 & n37362 ;
  assign n37721 = ~n37719 & ~n37720 ;
  assign n37722 = ~n20910 & ~n37721 ;
  assign n37723 = ~n37716 & ~n37722 ;
  assign n37724 = ~n37715 & n37723 ;
  assign n37725 = n32298 & ~n37724 ;
  assign n37726 = ~n37340 & ~n37725 ;
  assign n37727 = ~n37714 & n37726 ;
  assign n37728 = n37548 & n37727 ;
  assign n37729 = ~n37343 & ~n37728 ;
  assign n37730 = ~\pi0187  & ~n1689 ;
  assign n37731 = ~n21032 & ~n37730 ;
  assign n37732 = \pi0789  & n37731 ;
  assign n37733 = ~n23880 & ~n37732 ;
  assign n37734 = n23423 & n37733 ;
  assign n37735 = ~\pi0770  & n1689 ;
  assign n37736 = n20784 & n37735 ;
  assign n37737 = ~n37730 & ~n37736 ;
  assign n37738 = n20794 & ~n37737 ;
  assign n37739 = n20796 & ~n37738 ;
  assign n37740 = n20799 & ~n37737 ;
  assign n37741 = n20801 & ~n37740 ;
  assign n37742 = ~n37739 & ~n37741 ;
  assign n37743 = ~\pi0785  & ~n37730 ;
  assign n37744 = ~n37736 & n37743 ;
  assign n37745 = ~n20804 & ~n37744 ;
  assign n37746 = ~n20812 & n37745 ;
  assign n37747 = n37733 & n37746 ;
  assign n37748 = n37742 & n37747 ;
  assign n37749 = ~n37734 & ~n37748 ;
  assign n37750 = ~\pi0187  & \pi0792  ;
  assign n37751 = ~n1689 & n37750 ;
  assign n37752 = ~n20845 & n37751 ;
  assign n37753 = ~n20910 & ~n37752 ;
  assign n37754 = ~\pi0187  & \pi0788  ;
  assign n37755 = ~n1689 & n37754 ;
  assign n37756 = ~n20778 & n37755 ;
  assign n37757 = n37753 & ~n37756 ;
  assign n37758 = n37749 & n37757 ;
  assign n37759 = n20846 & n37753 ;
  assign n37760 = \pi0726  & n1689 ;
  assign n37761 = n20855 & n37760 ;
  assign n37762 = ~n20861 & n37761 ;
  assign n37763 = ~n37730 & ~n37762 ;
  assign n37764 = n20879 & ~n37763 ;
  assign n37765 = n20895 & n37764 ;
  assign n37766 = ~\pi0187  & \pi0647  ;
  assign n37767 = ~n1689 & n37766 ;
  assign n37768 = n20897 & ~n37767 ;
  assign n37769 = ~n37765 & n37768 ;
  assign n37770 = ~\pi0187  & ~\pi0647  ;
  assign n37771 = ~n1689 & n37770 ;
  assign n37772 = n20849 & ~n37771 ;
  assign n37773 = ~n24761 & ~n37772 ;
  assign n37774 = n31479 & n37764 ;
  assign n37775 = ~n37773 & ~n37774 ;
  assign n37776 = ~n37769 & ~n37775 ;
  assign n37777 = ~n37759 & n37776 ;
  assign n37778 = ~n37758 & n37777 ;
  assign n37779 = ~n29722 & ~n37778 ;
  assign n37780 = n20938 & n37764 ;
  assign n37781 = \pi0629  & ~n37756 ;
  assign n37782 = ~n37780 & n37781 ;
  assign n37783 = n37749 & n37782 ;
  assign n37784 = n21077 & n37764 ;
  assign n37785 = ~\pi0629  & ~n37756 ;
  assign n37786 = ~n37784 & n37785 ;
  assign n37787 = n37749 & n37786 ;
  assign n37788 = n29714 & ~n37780 ;
  assign n37789 = n29709 & ~n37784 ;
  assign n37790 = \pi0792  & ~n37789 ;
  assign n37791 = ~n37788 & n37790 ;
  assign n37792 = ~n37787 & n37791 ;
  assign n37793 = ~n37783 & n37792 ;
  assign n37794 = ~n21067 & ~n37793 ;
  assign n37795 = n23423 & ~n37732 ;
  assign n37796 = ~n37732 & n37746 ;
  assign n37797 = n37742 & n37796 ;
  assign n37798 = ~n37795 & ~n37797 ;
  assign n37799 = ~\pi0626  & n37798 ;
  assign n37800 = \pi0626  & ~n37730 ;
  assign n37801 = n20882 & ~n37800 ;
  assign n37802 = ~n37799 & n37801 ;
  assign n37803 = n23170 & ~n37763 ;
  assign n37804 = ~\pi0626  & ~n37730 ;
  assign n37805 = n20881 & ~n37804 ;
  assign n37806 = ~n37803 & ~n37805 ;
  assign n37807 = \pi0626  & ~n37803 ;
  assign n37808 = n37798 & n37807 ;
  assign n37809 = ~n37806 & ~n37808 ;
  assign n37810 = ~n37802 & ~n37809 ;
  assign n37811 = \pi0788  & ~n37810 ;
  assign n37812 = ~n23856 & n37811 ;
  assign n37813 = n20964 & n37745 ;
  assign n37814 = n37742 & n37813 ;
  assign n37815 = \pi0627  & ~n37730 ;
  assign n37816 = ~n37762 & n37815 ;
  assign n37817 = ~n20968 & ~n37816 ;
  assign n37818 = ~n37814 & ~n37817 ;
  assign n37819 = n20974 & n37745 ;
  assign n37820 = n37742 & n37819 ;
  assign n37821 = ~\pi0627  & ~n37730 ;
  assign n37822 = ~n37762 & n37821 ;
  assign n37823 = ~n20978 & ~n37822 ;
  assign n37824 = ~n37820 & ~n37823 ;
  assign n37825 = ~n37818 & ~n37824 ;
  assign n37826 = \pi0781  & n37825 ;
  assign n37827 = \pi0680  & \pi0726  ;
  assign n37828 = ~n20854 & n37827 ;
  assign n37829 = ~n20861 & n37828 ;
  assign n37830 = ~n20986 & n37829 ;
  assign n37831 = \pi0603  & ~\pi0770  ;
  assign n37832 = ~n20783 & n37831 ;
  assign n37833 = ~n20985 & n37832 ;
  assign n37834 = ~n37730 & ~n37833 ;
  assign n37835 = ~n37830 & n37834 ;
  assign n37836 = \pi0187  & ~n1689 ;
  assign n37837 = ~\pi0609  & ~n37836 ;
  assign n37838 = ~n37835 & n37837 ;
  assign n37839 = ~\pi1155  & ~n37730 ;
  assign n37840 = ~n37762 & n37839 ;
  assign n37841 = ~n20999 & ~n37840 ;
  assign n37842 = ~n37838 & ~n37841 ;
  assign n37843 = \pi1155  & ~n37740 ;
  assign n37844 = ~\pi0660  & ~n37843 ;
  assign n37845 = ~n37842 & n37844 ;
  assign n37846 = ~n21007 & ~n37739 ;
  assign n37847 = \pi0609  & ~n37836 ;
  assign n37848 = ~n37835 & n37847 ;
  assign n37849 = \pi1155  & ~n37730 ;
  assign n37850 = ~n37762 & n37849 ;
  assign n37851 = ~n21774 & ~n37850 ;
  assign n37852 = \pi0785  & ~n37851 ;
  assign n37853 = ~n37848 & n37852 ;
  assign n37854 = n37846 & ~n37853 ;
  assign n37855 = ~n37845 & ~n37854 ;
  assign n37856 = ~n37835 & ~n37836 ;
  assign n37857 = ~\pi0785  & ~n37856 ;
  assign n37858 = n21022 & ~n37857 ;
  assign n37859 = ~n37855 & n37858 ;
  assign n37860 = ~n21034 & ~n37859 ;
  assign n37861 = ~n37826 & n37860 ;
  assign n37862 = ~n20876 & n37731 ;
  assign n37863 = ~n24969 & ~n37862 ;
  assign n37864 = n37746 & ~n37862 ;
  assign n37865 = n37742 & n37864 ;
  assign n37866 = ~n37863 & ~n37865 ;
  assign n37867 = n21050 & ~n37730 ;
  assign n37868 = ~n37762 & n37867 ;
  assign n37869 = ~n21051 & ~n37868 ;
  assign n37870 = ~n21038 & n37869 ;
  assign n37871 = ~n37866 & n37870 ;
  assign n37872 = ~n23177 & ~n37871 ;
  assign n37873 = ~n23856 & ~n37872 ;
  assign n37874 = ~n37861 & n37873 ;
  assign n37875 = ~n37812 & ~n37874 ;
  assign n37876 = n37794 & n37875 ;
  assign n37877 = ~n37779 & ~n37876 ;
  assign n37878 = n24830 & n37764 ;
  assign n37879 = \pi1157  & ~n37771 ;
  assign n37880 = ~n37878 & n37879 ;
  assign n37881 = ~\pi1157  & ~n37767 ;
  assign n37882 = ~n37765 & n37881 ;
  assign n37883 = ~n37880 & ~n37882 ;
  assign n37884 = \pi0787  & ~n37883 ;
  assign n37885 = n24844 & n37764 ;
  assign n37886 = ~n24843 & ~n37885 ;
  assign n37887 = ~n37884 & ~n37886 ;
  assign n37888 = n37749 & ~n37756 ;
  assign n37889 = n31580 & ~n37888 ;
  assign n37890 = ~n37887 & ~n37889 ;
  assign n37891 = n23313 & ~n37890 ;
  assign n37892 = \pi0790  & n37891 ;
  assign n37893 = n31588 & ~n37888 ;
  assign n37894 = ~n23414 & n37730 ;
  assign n37895 = ~n24886 & n37894 ;
  assign n37896 = n20891 & n37764 ;
  assign n37897 = ~\pi0787  & ~n37896 ;
  assign n37898 = ~\pi1160  & ~n37897 ;
  assign n37899 = ~n37884 & n37898 ;
  assign n37900 = ~n37895 & ~n37899 ;
  assign n37901 = ~n37893 & n37900 ;
  assign n37902 = ~n23312 & ~n37895 ;
  assign n37903 = \pi0790  & ~n37902 ;
  assign n37904 = ~n37901 & n37903 ;
  assign n37905 = ~n37892 & ~n37904 ;
  assign n37906 = \pi0832  & n37905 ;
  assign n37907 = ~n37877 & n37906 ;
  assign n37908 = \pi0187  & ~\pi0832  ;
  assign n37909 = ~n21132 & ~n37908 ;
  assign n37910 = ~n37907 & n37909 ;
  assign n37911 = ~\pi0187  & n21768 ;
  assign n37912 = ~\pi0187  & n21770 ;
  assign n37913 = ~n21734 & n37912 ;
  assign n37914 = ~n37911 & ~n37913 ;
  assign n37915 = n23880 & ~n37914 ;
  assign n37916 = ~\pi0187  & \pi0618  ;
  assign n37917 = n21768 & n37916 ;
  assign n37918 = n21770 & n37916 ;
  assign n37919 = ~n21734 & n37918 ;
  assign n37920 = ~n37917 & ~n37919 ;
  assign n37921 = ~\pi1154  & n37920 ;
  assign n37922 = \pi0781  & ~n37921 ;
  assign n37923 = \pi0187  & ~n6861 ;
  assign n37924 = n21777 & n37923 ;
  assign n37925 = ~n23456 & ~n37924 ;
  assign n37926 = \pi0187  & \pi0770  ;
  assign n37927 = \pi0187  & ~n25040 ;
  assign n37928 = ~n37926 & ~n37927 ;
  assign n37929 = ~\pi0038  & ~n37926 ;
  assign n37930 = n25023 & n37929 ;
  assign n37931 = ~n37928 & ~n37930 ;
  assign n37932 = ~\pi0187  & ~\pi0770  ;
  assign n37933 = ~n25040 & n37932 ;
  assign n37934 = ~n25033 & n37933 ;
  assign n37935 = ~n25028 & n37934 ;
  assign n37936 = ~n37931 & ~n37935 ;
  assign n37937 = ~n27274 & ~n28084 ;
  assign n37938 = ~n37924 & ~n37937 ;
  assign n37939 = n37936 & n37938 ;
  assign n37940 = ~n37925 & ~n37939 ;
  assign n37941 = ~n21777 & n37914 ;
  assign n37942 = ~\pi0618  & ~n37941 ;
  assign n37943 = \pi0781  & n37942 ;
  assign n37944 = ~n37940 & n37943 ;
  assign n37945 = ~n37922 & ~n37944 ;
  assign n37946 = \pi0618  & ~n37941 ;
  assign n37947 = ~n37940 & n37946 ;
  assign n37948 = ~\pi0187  & ~\pi0618  ;
  assign n37949 = n21768 & n37948 ;
  assign n37950 = n21770 & n37948 ;
  assign n37951 = ~n21734 & n37950 ;
  assign n37952 = ~n37949 & ~n37951 ;
  assign n37953 = \pi1154  & n37952 ;
  assign n37954 = ~n37947 & n37953 ;
  assign n37955 = ~n37945 & ~n37954 ;
  assign n37956 = ~\pi0781  & ~n37941 ;
  assign n37957 = ~n37940 & n37956 ;
  assign n37958 = ~\pi0789  & ~n37957 ;
  assign n37959 = ~n37955 & n37958 ;
  assign n37960 = ~n23880 & ~n37959 ;
  assign n37961 = n21092 & ~n37960 ;
  assign n37962 = ~\pi0619  & ~n37953 ;
  assign n37963 = ~\pi0619  & n37946 ;
  assign n37964 = ~n37940 & n37963 ;
  assign n37965 = ~n37962 & ~n37964 ;
  assign n37966 = ~n37945 & ~n37965 ;
  assign n37967 = ~\pi0619  & n37956 ;
  assign n37968 = ~n37940 & n37967 ;
  assign n37969 = ~\pi0187  & \pi0619  ;
  assign n37970 = n21768 & n37969 ;
  assign n37971 = n21770 & n37969 ;
  assign n37972 = ~n21734 & n37971 ;
  assign n37973 = ~n37970 & ~n37972 ;
  assign n37974 = ~\pi1159  & n37973 ;
  assign n37975 = ~n37968 & n37974 ;
  assign n37976 = ~n37966 & n37975 ;
  assign n37977 = ~\pi0187  & ~\pi0619  ;
  assign n37978 = n21768 & n37977 ;
  assign n37979 = n21770 & n37977 ;
  assign n37980 = ~n21734 & n37979 ;
  assign n37981 = ~n37978 & ~n37980 ;
  assign n37982 = \pi1159  & n37981 ;
  assign n37983 = ~\pi0619  & n37982 ;
  assign n37984 = ~n37957 & n37982 ;
  assign n37985 = ~n37955 & n37984 ;
  assign n37986 = ~n37983 & ~n37985 ;
  assign n37987 = ~n37976 & n37986 ;
  assign n37988 = n32328 & ~n37987 ;
  assign n37989 = ~n37961 & ~n37988 ;
  assign n37990 = ~n37915 & ~n37989 ;
  assign n37991 = ~n21092 & n37914 ;
  assign n37992 = ~\pi0644  & ~n37991 ;
  assign n37993 = ~n37990 & n37992 ;
  assign n37994 = ~\pi0187  & \pi0644  ;
  assign n37995 = n21768 & n37994 ;
  assign n37996 = n21770 & n37994 ;
  assign n37997 = ~n21734 & n37996 ;
  assign n37998 = ~n37995 & ~n37997 ;
  assign n37999 = n23413 & n37998 ;
  assign n38000 = ~n37993 & n37999 ;
  assign n38001 = \pi0644  & ~n37991 ;
  assign n38002 = ~n37990 & n38001 ;
  assign n38003 = ~\pi0187  & ~\pi0644  ;
  assign n38004 = n21768 & n38003 ;
  assign n38005 = n21770 & n38003 ;
  assign n38006 = ~n21734 & n38005 ;
  assign n38007 = ~n38004 & ~n38006 ;
  assign n38008 = n23412 & n38007 ;
  assign n38009 = ~n38002 & n38008 ;
  assign n38010 = ~n38000 & ~n38009 ;
  assign n38011 = \pi0790  & ~n38010 ;
  assign n38012 = ~\pi0187  & ~\pi0726  ;
  assign n38013 = ~\pi0038  & n38012 ;
  assign n38014 = n21743 & n38013 ;
  assign n38015 = ~n21734 & n38014 ;
  assign n38016 = \pi0038  & n38012 ;
  assign n38017 = ~n22123 & n38016 ;
  assign n38018 = n6861 & ~n38017 ;
  assign n38019 = ~n38015 & n38018 ;
  assign n38020 = ~n37923 & ~n38019 ;
  assign n38021 = ~\pi0187  & ~n22017 ;
  assign n38022 = ~n21994 & n38021 ;
  assign n38023 = ~\pi0038  & ~\pi0187  ;
  assign n38024 = ~n22109 & ~n38023 ;
  assign n38025 = ~n38022 & ~n38024 ;
  assign n38026 = ~\pi0187  & ~n21757 ;
  assign n38027 = n22117 & ~n38026 ;
  assign n38028 = \pi0726  & ~n37923 ;
  assign n38029 = ~n38027 & n38028 ;
  assign n38030 = ~n38025 & n38029 ;
  assign n38031 = ~n38020 & ~n38030 ;
  assign n38032 = \pi0625  & ~n38031 ;
  assign n38033 = ~\pi0187  & ~\pi0625  ;
  assign n38034 = n21768 & n38033 ;
  assign n38035 = n21770 & n38033 ;
  assign n38036 = ~n21734 & n38035 ;
  assign n38037 = ~n38034 & ~n38036 ;
  assign n38038 = \pi1153  & n38037 ;
  assign n38039 = ~n38032 & n38038 ;
  assign n38040 = ~\pi0625  & ~n38031 ;
  assign n38041 = ~\pi0187  & \pi0625  ;
  assign n38042 = n21768 & n38041 ;
  assign n38043 = n21770 & n38041 ;
  assign n38044 = ~n21734 & n38043 ;
  assign n38045 = ~n38042 & ~n38044 ;
  assign n38046 = ~\pi1153  & n38045 ;
  assign n38047 = ~n38040 & n38046 ;
  assign n38048 = ~n38039 & ~n38047 ;
  assign n38049 = n22148 & ~n38048 ;
  assign n38050 = n22151 & n38031 ;
  assign n38051 = n22147 & n37914 ;
  assign n38052 = ~n22155 & ~n38051 ;
  assign n38053 = ~n38050 & n38052 ;
  assign n38054 = ~n38049 & n38053 ;
  assign n38055 = n22155 & ~n37914 ;
  assign n38056 = n22162 & ~n38055 ;
  assign n38057 = ~n38054 & n38056 ;
  assign n38058 = ~n22162 & n37914 ;
  assign n38059 = ~\pi0647  & ~n38058 ;
  assign n38060 = ~n38057 & n38059 ;
  assign n38061 = ~n22913 & ~n38060 ;
  assign n38062 = n21768 & n37766 ;
  assign n38063 = n21770 & n37766 ;
  assign n38064 = ~n21734 & n38063 ;
  assign n38065 = ~n38062 & ~n38064 ;
  assign n38066 = ~\pi1157  & n38065 ;
  assign n38067 = n38061 & n38066 ;
  assign n38068 = \pi0628  & ~n38058 ;
  assign n38069 = ~n38057 & n38068 ;
  assign n38070 = ~\pi0187  & ~\pi0628  ;
  assign n38071 = n21768 & n38070 ;
  assign n38072 = n21770 & n38070 ;
  assign n38073 = ~n21734 & n38072 ;
  assign n38074 = ~n38071 & ~n38073 ;
  assign n38075 = \pi1156  & n38074 ;
  assign n38076 = ~n38069 & n38075 ;
  assign n38077 = ~\pi0628  & ~n38058 ;
  assign n38078 = ~n38057 & n38077 ;
  assign n38079 = ~\pi0187  & \pi0628  ;
  assign n38080 = n21768 & n38079 ;
  assign n38081 = n21770 & n38079 ;
  assign n38082 = ~n21734 & n38081 ;
  assign n38083 = ~n38080 & ~n38082 ;
  assign n38084 = ~\pi1156  & n38083 ;
  assign n38085 = ~n38078 & n38084 ;
  assign n38086 = ~n38076 & ~n38085 ;
  assign n38087 = \pi0792  & n38066 ;
  assign n38088 = ~n38086 & n38087 ;
  assign n38089 = ~n38067 & ~n38088 ;
  assign n38090 = \pi0787  & n38089 ;
  assign n38091 = \pi0647  & ~n38058 ;
  assign n38092 = ~n38057 & n38091 ;
  assign n38093 = ~n22956 & ~n38092 ;
  assign n38094 = n21768 & n37770 ;
  assign n38095 = n21770 & n37770 ;
  assign n38096 = ~n21734 & n38095 ;
  assign n38097 = ~n38094 & ~n38096 ;
  assign n38098 = \pi1157  & n38097 ;
  assign n38099 = n38093 & n38098 ;
  assign n38100 = \pi0792  & n38098 ;
  assign n38101 = ~n38086 & n38100 ;
  assign n38102 = ~n38099 & ~n38101 ;
  assign n38103 = n38090 & n38102 ;
  assign n38104 = ~\pi0787  & ~n38058 ;
  assign n38105 = ~n38057 & n38104 ;
  assign n38106 = ~n33084 & ~n38105 ;
  assign n38107 = n23518 & n38106 ;
  assign n38108 = n37542 & ~n38086 ;
  assign n38109 = ~n38107 & ~n38108 ;
  assign n38110 = \pi0790  & ~n38109 ;
  assign n38111 = ~n38103 & n38110 ;
  assign n38112 = ~n38011 & ~n38111 ;
  assign n38113 = n9948 & n38112 ;
  assign n38114 = n24691 & ~n37915 ;
  assign n38115 = ~n37960 & n38114 ;
  assign n38116 = \pi0789  & n38114 ;
  assign n38117 = ~n37987 & n38116 ;
  assign n38118 = ~n38115 & ~n38117 ;
  assign n38119 = ~\pi0629  & n38075 ;
  assign n38120 = ~n38069 & n38119 ;
  assign n38121 = \pi0629  & n38084 ;
  assign n38122 = ~n38078 & n38121 ;
  assign n38123 = ~n38120 & ~n38122 ;
  assign n38124 = n38118 & n38123 ;
  assign n38125 = n24724 & ~n38124 ;
  assign n38126 = ~n21067 & n26803 ;
  assign n38127 = \pi0789  & ~n37987 ;
  assign n38128 = n30606 & ~n37959 ;
  assign n38129 = ~n38127 & n38128 ;
  assign n38130 = ~n22849 & n37914 ;
  assign n38131 = \pi0641  & n38130 ;
  assign n38132 = ~n38050 & ~n38051 ;
  assign n38133 = ~n38049 & n38132 ;
  assign n38134 = n33656 & ~n38133 ;
  assign n38135 = ~n38131 & ~n38134 ;
  assign n38136 = ~\pi0641  & n37914 ;
  assign n38137 = n20776 & ~n38136 ;
  assign n38138 = n38135 & n38137 ;
  assign n38139 = ~n38129 & ~n38138 ;
  assign n38140 = ~\pi0641  & n38130 ;
  assign n38141 = n33649 & ~n38133 ;
  assign n38142 = ~n38140 & ~n38141 ;
  assign n38143 = \pi0641  & n37914 ;
  assign n38144 = n20777 & ~n38143 ;
  assign n38145 = n38142 & n38144 ;
  assign n38146 = ~n23856 & ~n38145 ;
  assign n38147 = ~n21067 & n38146 ;
  assign n38148 = n38139 & n38147 ;
  assign n38149 = ~n38126 & ~n38148 ;
  assign n38150 = ~n38125 & n38149 ;
  assign n38151 = ~n22734 & ~n38033 ;
  assign n38152 = ~n6861 & ~n38151 ;
  assign n38153 = ~n37937 & ~n38151 ;
  assign n38154 = n37936 & n38153 ;
  assign n38155 = ~n38152 & ~n38154 ;
  assign n38156 = \pi1153  & n38155 ;
  assign n38157 = \pi0608  & ~n38046 ;
  assign n38158 = n22740 & ~n38031 ;
  assign n38159 = ~n38157 & ~n38158 ;
  assign n38160 = ~n38156 & ~n38159 ;
  assign n38161 = \pi0038  & \pi0187  ;
  assign n38162 = ~n22708 & n38161 ;
  assign n38163 = ~\pi0038  & \pi0187  ;
  assign n38164 = ~n38162 & ~n38163 ;
  assign n38165 = ~n23558 & ~n38162 ;
  assign n38166 = n23557 & n38165 ;
  assign n38167 = ~n38164 & ~n38166 ;
  assign n38168 = ~\pi0187  & n23548 ;
  assign n38169 = ~n25191 & n38168 ;
  assign n38170 = ~n25190 & n38169 ;
  assign n38171 = \pi0726  & ~\pi0770  ;
  assign n38172 = ~n38170 & n38171 ;
  assign n38173 = ~n38167 & n38172 ;
  assign n38174 = ~\pi0187  & ~n25209 ;
  assign n38175 = ~n25204 & n38174 ;
  assign n38176 = n23575 & n38163 ;
  assign n38177 = n23572 & n38176 ;
  assign n38178 = ~n25217 & ~n38177 ;
  assign n38179 = ~n38175 & n38178 ;
  assign n38180 = n27147 & ~n38179 ;
  assign n38181 = ~n38173 & ~n38180 ;
  assign n38182 = ~\pi0726  & ~n37931 ;
  assign n38183 = ~n37935 & n38182 ;
  assign n38184 = ~n37937 & n38183 ;
  assign n38185 = n6861 & ~n38184 ;
  assign n38186 = n38181 & n38185 ;
  assign n38187 = ~n22727 & ~n38041 ;
  assign n38188 = ~n38159 & ~n38187 ;
  assign n38189 = ~n38186 & n38188 ;
  assign n38190 = ~n38160 & ~n38189 ;
  assign n38191 = n23613 & ~n38190 ;
  assign n38192 = ~n6861 & ~n38187 ;
  assign n38193 = ~n37937 & ~n38187 ;
  assign n38194 = n37936 & n38193 ;
  assign n38195 = ~n38192 & ~n38194 ;
  assign n38196 = n38151 & n38195 ;
  assign n38197 = n38185 & n38195 ;
  assign n38198 = n38181 & n38197 ;
  assign n38199 = ~n38196 & ~n38198 ;
  assign n38200 = ~\pi1153  & ~n38199 ;
  assign n38201 = ~\pi0608  & ~n38038 ;
  assign n38202 = n22755 & ~n38031 ;
  assign n38203 = ~n38201 & ~n38202 ;
  assign n38204 = n23613 & ~n38203 ;
  assign n38205 = ~n38200 & n38204 ;
  assign n38206 = ~n38191 & ~n38205 ;
  assign n38207 = \pi0778  & ~n38048 ;
  assign n38208 = ~\pi0778  & n38031 ;
  assign n38209 = \pi0609  & ~n38208 ;
  assign n38210 = ~n38207 & n38209 ;
  assign n38211 = ~\pi0187  & ~\pi0778  ;
  assign n38212 = ~n23622 & ~n38211 ;
  assign n38213 = ~\pi0609  & ~n38212 ;
  assign n38214 = ~n38186 & n38213 ;
  assign n38215 = ~\pi1155  & ~n38214 ;
  assign n38216 = ~n38210 & n38215 ;
  assign n38217 = n38206 & n38216 ;
  assign n38218 = ~n20985 & n37923 ;
  assign n38219 = ~n26645 & ~n38218 ;
  assign n38220 = ~n37937 & ~n38218 ;
  assign n38221 = n37936 & n38220 ;
  assign n38222 = ~n38219 & ~n38221 ;
  assign n38223 = n21774 & n38222 ;
  assign n38224 = n26653 & n37914 ;
  assign n38225 = ~\pi0660  & ~n38224 ;
  assign n38226 = ~n38223 & n38225 ;
  assign n38227 = ~n38217 & n38226 ;
  assign n38228 = n20999 & n38222 ;
  assign n38229 = ~n32768 & n37914 ;
  assign n38230 = \pi0660  & ~n38229 ;
  assign n38231 = ~n38228 & n38230 ;
  assign n38232 = \pi0785  & ~n38231 ;
  assign n38233 = n23638 & ~n38190 ;
  assign n38234 = n23638 & ~n38203 ;
  assign n38235 = ~n38200 & n38234 ;
  assign n38236 = ~n38233 & ~n38235 ;
  assign n38237 = ~\pi0609  & ~n38208 ;
  assign n38238 = \pi1155  & ~n38237 ;
  assign n38239 = n22722 & ~n38048 ;
  assign n38240 = ~n38238 & ~n38239 ;
  assign n38241 = \pi0609  & ~n38212 ;
  assign n38242 = ~n38186 & n38241 ;
  assign n38243 = \pi0785  & ~n38242 ;
  assign n38244 = ~n38240 & n38243 ;
  assign n38245 = n38236 & n38244 ;
  assign n38246 = ~n38232 & ~n38245 ;
  assign n38247 = ~n38227 & ~n38246 ;
  assign n38248 = n21019 & ~n37921 ;
  assign n38249 = n21020 & n37952 ;
  assign n38250 = ~n33630 & ~n38249 ;
  assign n38251 = ~n38248 & ~n38250 ;
  assign n38252 = n20828 & n37981 ;
  assign n38253 = ~\pi0619  & n38252 ;
  assign n38254 = ~n37957 & n38252 ;
  assign n38255 = ~n37955 & n38254 ;
  assign n38256 = ~n38253 & ~n38255 ;
  assign n38257 = n32121 & ~n37973 ;
  assign n38258 = n32125 & ~n38257 ;
  assign n38259 = n38256 & ~n38258 ;
  assign n38260 = \pi0789  & ~n38259 ;
  assign n38261 = \pi0778  & ~n38190 ;
  assign n38262 = \pi0778  & ~n38203 ;
  assign n38263 = ~n38200 & n38262 ;
  assign n38264 = ~n38261 & ~n38263 ;
  assign n38265 = ~\pi0785  & n38212 ;
  assign n38266 = ~\pi0785  & n38185 ;
  assign n38267 = n38181 & n38266 ;
  assign n38268 = ~n38265 & ~n38267 ;
  assign n38269 = n38264 & ~n38268 ;
  assign n38270 = ~n38260 & ~n38269 ;
  assign n38271 = ~n38251 & n38270 ;
  assign n38272 = ~n38247 & n38271 ;
  assign n38273 = ~\pi1159  & ~n38055 ;
  assign n38274 = ~n38054 & n38273 ;
  assign n38275 = ~n22872 & ~n38274 ;
  assign n38276 = ~\pi0648  & n37986 ;
  assign n38277 = n38275 & n38276 ;
  assign n38278 = \pi1159  & ~n38055 ;
  assign n38279 = ~n38054 & n38278 ;
  assign n38280 = n37561 & ~n37976 ;
  assign n38281 = ~n38279 & n38280 ;
  assign n38282 = ~n38277 & ~n38281 ;
  assign n38283 = \pi0789  & ~n38282 ;
  assign n38284 = ~\pi0618  & ~n38051 ;
  assign n38285 = ~n38050 & n38284 ;
  assign n38286 = ~n38049 & n38285 ;
  assign n38287 = \pi1154  & ~n38286 ;
  assign n38288 = \pi0627  & ~n37921 ;
  assign n38289 = \pi0627  & n37942 ;
  assign n38290 = ~n37940 & n38289 ;
  assign n38291 = ~n38288 & ~n38290 ;
  assign n38292 = ~n38287 & ~n38291 ;
  assign n38293 = \pi0618  & ~n38051 ;
  assign n38294 = ~n38050 & n38293 ;
  assign n38295 = ~n38049 & n38294 ;
  assign n38296 = ~\pi1154  & ~n38295 ;
  assign n38297 = ~\pi0627  & ~n37953 ;
  assign n38298 = ~\pi0627  & n37946 ;
  assign n38299 = ~n37940 & n38298 ;
  assign n38300 = ~n38297 & ~n38299 ;
  assign n38301 = ~n38296 & ~n38300 ;
  assign n38302 = ~n38292 & ~n38301 ;
  assign n38303 = ~n38260 & ~n38302 ;
  assign n38304 = \pi0781  & n38303 ;
  assign n38305 = ~n38283 & ~n38304 ;
  assign n38306 = ~n38272 & n38305 ;
  assign n38307 = ~n21038 & ~n38125 ;
  assign n38308 = ~n38306 & n38307 ;
  assign n38309 = ~n38150 & ~n38308 ;
  assign n38310 = ~n24761 & n38309 ;
  assign n38311 = ~n30376 & n37914 ;
  assign n38312 = ~n20910 & n38311 ;
  assign n38313 = ~\pi0789  & ~n37959 ;
  assign n38314 = ~n37959 & ~n37976 ;
  assign n38315 = n37986 & n38314 ;
  assign n38316 = ~n38313 & ~n38315 ;
  assign n38317 = n33670 & n38316 ;
  assign n38318 = ~n38312 & ~n38317 ;
  assign n38319 = ~\pi0630  & n38318 ;
  assign n38320 = n38102 & n38319 ;
  assign n38321 = \pi0630  & n38318 ;
  assign n38322 = n38089 & n38321 ;
  assign n38323 = ~n38320 & ~n38322 ;
  assign n38324 = n32298 & n38323 ;
  assign n38325 = ~n37907 & ~n38324 ;
  assign n38326 = ~n38310 & n38325 ;
  assign n38327 = n38113 & n38326 ;
  assign n38328 = ~n37910 & ~n38327 ;
  assign n38329 = ~\pi0188  & ~n1689 ;
  assign n38330 = ~n21032 & ~n38329 ;
  assign n38331 = \pi0789  & n38330 ;
  assign n38332 = ~n23880 & ~n38331 ;
  assign n38333 = n23423 & n38332 ;
  assign n38334 = ~\pi0768  & n1689 ;
  assign n38335 = n20784 & n38334 ;
  assign n38336 = ~n38329 & ~n38335 ;
  assign n38337 = n20794 & ~n38336 ;
  assign n38338 = n20796 & ~n38337 ;
  assign n38339 = n20799 & ~n38336 ;
  assign n38340 = n20801 & ~n38339 ;
  assign n38341 = ~n38338 & ~n38340 ;
  assign n38342 = ~\pi0785  & ~n38329 ;
  assign n38343 = ~n38335 & n38342 ;
  assign n38344 = ~n20804 & ~n38343 ;
  assign n38345 = ~n20812 & n38344 ;
  assign n38346 = n38332 & n38345 ;
  assign n38347 = n38341 & n38346 ;
  assign n38348 = ~n38333 & ~n38347 ;
  assign n38349 = ~\pi0188  & \pi0792  ;
  assign n38350 = ~n1689 & n38349 ;
  assign n38351 = ~n20845 & n38350 ;
  assign n38352 = ~n20910 & ~n38351 ;
  assign n38353 = ~\pi0188  & \pi0788  ;
  assign n38354 = ~n1689 & n38353 ;
  assign n38355 = ~n20778 & n38354 ;
  assign n38356 = n38352 & ~n38355 ;
  assign n38357 = n38348 & n38356 ;
  assign n38358 = n20846 & n38352 ;
  assign n38359 = \pi0705  & n1689 ;
  assign n38360 = n20855 & n38359 ;
  assign n38361 = ~n20861 & n38360 ;
  assign n38362 = ~n38329 & ~n38361 ;
  assign n38363 = n20879 & ~n38362 ;
  assign n38364 = n20895 & n38363 ;
  assign n38365 = ~\pi0188  & \pi0647  ;
  assign n38366 = ~n1689 & n38365 ;
  assign n38367 = n20897 & ~n38366 ;
  assign n38368 = ~n38364 & n38367 ;
  assign n38369 = ~\pi0188  & ~\pi0647  ;
  assign n38370 = ~n1689 & n38369 ;
  assign n38371 = n20849 & ~n38370 ;
  assign n38372 = ~n24761 & ~n38371 ;
  assign n38373 = n31479 & n38363 ;
  assign n38374 = ~n38372 & ~n38373 ;
  assign n38375 = ~n38368 & ~n38374 ;
  assign n38376 = ~n38358 & n38375 ;
  assign n38377 = ~n38357 & n38376 ;
  assign n38378 = ~n29722 & ~n38377 ;
  assign n38379 = n20938 & n38363 ;
  assign n38380 = \pi0629  & ~n38355 ;
  assign n38381 = ~n38379 & n38380 ;
  assign n38382 = n38348 & n38381 ;
  assign n38383 = n21077 & n38363 ;
  assign n38384 = ~\pi0629  & ~n38355 ;
  assign n38385 = ~n38383 & n38384 ;
  assign n38386 = n38348 & n38385 ;
  assign n38387 = n29714 & ~n38379 ;
  assign n38388 = n29709 & ~n38383 ;
  assign n38389 = \pi0792  & ~n38388 ;
  assign n38390 = ~n38387 & n38389 ;
  assign n38391 = ~n38386 & n38390 ;
  assign n38392 = ~n38382 & n38391 ;
  assign n38393 = ~n21067 & ~n38392 ;
  assign n38394 = n23423 & ~n38331 ;
  assign n38395 = ~n38331 & n38345 ;
  assign n38396 = n38341 & n38395 ;
  assign n38397 = ~n38394 & ~n38396 ;
  assign n38398 = ~\pi0626  & n38397 ;
  assign n38399 = \pi0626  & ~n38329 ;
  assign n38400 = n20882 & ~n38399 ;
  assign n38401 = ~n38398 & n38400 ;
  assign n38402 = n23170 & ~n38362 ;
  assign n38403 = ~\pi0626  & ~n38329 ;
  assign n38404 = n20881 & ~n38403 ;
  assign n38405 = ~n38402 & ~n38404 ;
  assign n38406 = \pi0626  & ~n38402 ;
  assign n38407 = n38397 & n38406 ;
  assign n38408 = ~n38405 & ~n38407 ;
  assign n38409 = ~n38401 & ~n38408 ;
  assign n38410 = \pi0788  & ~n38409 ;
  assign n38411 = ~n23856 & n38410 ;
  assign n38412 = n20964 & n38344 ;
  assign n38413 = n38341 & n38412 ;
  assign n38414 = \pi0627  & ~n38329 ;
  assign n38415 = ~n38361 & n38414 ;
  assign n38416 = ~n20968 & ~n38415 ;
  assign n38417 = ~n38413 & ~n38416 ;
  assign n38418 = n20974 & n38344 ;
  assign n38419 = n38341 & n38418 ;
  assign n38420 = ~\pi0627  & ~n38329 ;
  assign n38421 = ~n38361 & n38420 ;
  assign n38422 = ~n20978 & ~n38421 ;
  assign n38423 = ~n38419 & ~n38422 ;
  assign n38424 = ~n38417 & ~n38423 ;
  assign n38425 = \pi0781  & n38424 ;
  assign n38426 = \pi0680  & \pi0705  ;
  assign n38427 = ~n20854 & n38426 ;
  assign n38428 = ~n20861 & n38427 ;
  assign n38429 = ~n20986 & n38428 ;
  assign n38430 = \pi0603  & ~\pi0768  ;
  assign n38431 = ~n20783 & n38430 ;
  assign n38432 = ~n20985 & n38431 ;
  assign n38433 = ~n38329 & ~n38432 ;
  assign n38434 = ~n38429 & n38433 ;
  assign n38435 = \pi0188  & ~n1689 ;
  assign n38436 = ~\pi0609  & ~n38435 ;
  assign n38437 = ~n38434 & n38436 ;
  assign n38438 = ~\pi1155  & ~n38329 ;
  assign n38439 = ~n38361 & n38438 ;
  assign n38440 = ~n20999 & ~n38439 ;
  assign n38441 = ~n38437 & ~n38440 ;
  assign n38442 = \pi1155  & ~n38339 ;
  assign n38443 = ~\pi0660  & ~n38442 ;
  assign n38444 = ~n38441 & n38443 ;
  assign n38445 = ~n21007 & ~n38338 ;
  assign n38446 = \pi0609  & ~n38435 ;
  assign n38447 = ~n38434 & n38446 ;
  assign n38448 = \pi1155  & ~n38329 ;
  assign n38449 = ~n38361 & n38448 ;
  assign n38450 = ~n21774 & ~n38449 ;
  assign n38451 = \pi0785  & ~n38450 ;
  assign n38452 = ~n38447 & n38451 ;
  assign n38453 = n38445 & ~n38452 ;
  assign n38454 = ~n38444 & ~n38453 ;
  assign n38455 = ~n38434 & ~n38435 ;
  assign n38456 = ~\pi0785  & ~n38455 ;
  assign n38457 = n21022 & ~n38456 ;
  assign n38458 = ~n38454 & n38457 ;
  assign n38459 = ~n21034 & ~n38458 ;
  assign n38460 = ~n38425 & n38459 ;
  assign n38461 = ~n20876 & n38330 ;
  assign n38462 = ~n24969 & ~n38461 ;
  assign n38463 = n38345 & ~n38461 ;
  assign n38464 = n38341 & n38463 ;
  assign n38465 = ~n38462 & ~n38464 ;
  assign n38466 = n21050 & ~n38329 ;
  assign n38467 = ~n38361 & n38466 ;
  assign n38468 = ~n21051 & ~n38467 ;
  assign n38469 = ~n21038 & n38468 ;
  assign n38470 = ~n38465 & n38469 ;
  assign n38471 = ~n23177 & ~n38470 ;
  assign n38472 = ~n23856 & ~n38471 ;
  assign n38473 = ~n38460 & n38472 ;
  assign n38474 = ~n38411 & ~n38473 ;
  assign n38475 = n38393 & n38474 ;
  assign n38476 = ~n38378 & ~n38475 ;
  assign n38477 = n24830 & n38363 ;
  assign n38478 = \pi1157  & ~n38370 ;
  assign n38479 = ~n38477 & n38478 ;
  assign n38480 = ~\pi1157  & ~n38366 ;
  assign n38481 = ~n38364 & n38480 ;
  assign n38482 = ~n38479 & ~n38481 ;
  assign n38483 = \pi0787  & ~n38482 ;
  assign n38484 = n24844 & n38363 ;
  assign n38485 = ~n24843 & ~n38484 ;
  assign n38486 = ~n38483 & ~n38485 ;
  assign n38487 = n38348 & ~n38355 ;
  assign n38488 = n31580 & ~n38487 ;
  assign n38489 = ~n38486 & ~n38488 ;
  assign n38490 = n23313 & ~n38489 ;
  assign n38491 = \pi0790  & n38490 ;
  assign n38492 = n31588 & ~n38487 ;
  assign n38493 = ~n23414 & n38329 ;
  assign n38494 = ~n24886 & n38493 ;
  assign n38495 = n20891 & n38363 ;
  assign n38496 = ~\pi0787  & ~n38495 ;
  assign n38497 = ~\pi1160  & ~n38496 ;
  assign n38498 = ~n38483 & n38497 ;
  assign n38499 = ~n38494 & ~n38498 ;
  assign n38500 = ~n38492 & n38499 ;
  assign n38501 = ~n23312 & ~n38494 ;
  assign n38502 = \pi0790  & ~n38501 ;
  assign n38503 = ~n38500 & n38502 ;
  assign n38504 = ~n38491 & ~n38503 ;
  assign n38505 = \pi0832  & n38504 ;
  assign n38506 = ~n38476 & n38505 ;
  assign n38507 = \pi0188  & ~\pi0832  ;
  assign n38508 = ~n21132 & ~n38507 ;
  assign n38509 = ~n38506 & n38508 ;
  assign n38510 = ~\pi0188  & n21768 ;
  assign n38511 = ~\pi0188  & n21770 ;
  assign n38512 = ~n21734 & n38511 ;
  assign n38513 = ~n38510 & ~n38512 ;
  assign n38514 = n23880 & ~n38513 ;
  assign n38515 = ~\pi0188  & \pi0618  ;
  assign n38516 = n21768 & n38515 ;
  assign n38517 = n21770 & n38515 ;
  assign n38518 = ~n21734 & n38517 ;
  assign n38519 = ~n38516 & ~n38518 ;
  assign n38520 = ~\pi1154  & n38519 ;
  assign n38521 = \pi0781  & ~n38520 ;
  assign n38522 = \pi0188  & ~n6861 ;
  assign n38523 = n21777 & n38522 ;
  assign n38524 = ~n23456 & ~n38523 ;
  assign n38525 = \pi0188  & \pi0768  ;
  assign n38526 = \pi0188  & ~n25040 ;
  assign n38527 = ~n38525 & ~n38526 ;
  assign n38528 = ~\pi0038  & ~n38525 ;
  assign n38529 = n25023 & n38528 ;
  assign n38530 = ~n38527 & ~n38529 ;
  assign n38531 = ~\pi0188  & ~\pi0768  ;
  assign n38532 = ~n25040 & n38531 ;
  assign n38533 = ~n25033 & n38532 ;
  assign n38534 = ~n25028 & n38533 ;
  assign n38535 = ~n38530 & ~n38534 ;
  assign n38536 = ~n29124 & ~n38523 ;
  assign n38537 = n38535 & n38536 ;
  assign n38538 = ~n38524 & ~n38537 ;
  assign n38539 = ~n21777 & n38513 ;
  assign n38540 = ~\pi0618  & ~n38539 ;
  assign n38541 = \pi0781  & n38540 ;
  assign n38542 = ~n38538 & n38541 ;
  assign n38543 = ~n38521 & ~n38542 ;
  assign n38544 = \pi0618  & ~n38539 ;
  assign n38545 = ~n38538 & n38544 ;
  assign n38546 = ~\pi0188  & ~\pi0618  ;
  assign n38547 = n21768 & n38546 ;
  assign n38548 = n21770 & n38546 ;
  assign n38549 = ~n21734 & n38548 ;
  assign n38550 = ~n38547 & ~n38549 ;
  assign n38551 = \pi1154  & n38550 ;
  assign n38552 = ~n38545 & n38551 ;
  assign n38553 = ~n38543 & ~n38552 ;
  assign n38554 = ~\pi0781  & ~n38539 ;
  assign n38555 = ~n38538 & n38554 ;
  assign n38556 = ~\pi0789  & ~n38555 ;
  assign n38557 = ~n38553 & n38556 ;
  assign n38558 = ~n23880 & ~n38557 ;
  assign n38559 = n21092 & ~n38558 ;
  assign n38560 = ~\pi0619  & ~n38551 ;
  assign n38561 = ~\pi0619  & n38544 ;
  assign n38562 = ~n38538 & n38561 ;
  assign n38563 = ~n38560 & ~n38562 ;
  assign n38564 = ~n38543 & ~n38563 ;
  assign n38565 = ~\pi0619  & n38554 ;
  assign n38566 = ~n38538 & n38565 ;
  assign n38567 = ~\pi0188  & \pi0619  ;
  assign n38568 = n21768 & n38567 ;
  assign n38569 = n21770 & n38567 ;
  assign n38570 = ~n21734 & n38569 ;
  assign n38571 = ~n38568 & ~n38570 ;
  assign n38572 = ~\pi1159  & n38571 ;
  assign n38573 = ~n38566 & n38572 ;
  assign n38574 = ~n38564 & n38573 ;
  assign n38575 = ~\pi0188  & ~\pi0619  ;
  assign n38576 = n21768 & n38575 ;
  assign n38577 = n21770 & n38575 ;
  assign n38578 = ~n21734 & n38577 ;
  assign n38579 = ~n38576 & ~n38578 ;
  assign n38580 = \pi1159  & n38579 ;
  assign n38581 = ~\pi0619  & n38580 ;
  assign n38582 = ~n38555 & n38580 ;
  assign n38583 = ~n38553 & n38582 ;
  assign n38584 = ~n38581 & ~n38583 ;
  assign n38585 = ~n38574 & n38584 ;
  assign n38586 = n32328 & ~n38585 ;
  assign n38587 = ~n38559 & ~n38586 ;
  assign n38588 = ~n38514 & ~n38587 ;
  assign n38589 = ~n21092 & n38513 ;
  assign n38590 = ~\pi0644  & ~n38589 ;
  assign n38591 = ~n38588 & n38590 ;
  assign n38592 = ~\pi0188  & \pi0644  ;
  assign n38593 = n21768 & n38592 ;
  assign n38594 = n21770 & n38592 ;
  assign n38595 = ~n21734 & n38594 ;
  assign n38596 = ~n38593 & ~n38595 ;
  assign n38597 = n23413 & n38596 ;
  assign n38598 = ~n38591 & n38597 ;
  assign n38599 = \pi0644  & ~n38589 ;
  assign n38600 = ~n38588 & n38599 ;
  assign n38601 = ~\pi0188  & ~\pi0644  ;
  assign n38602 = n21768 & n38601 ;
  assign n38603 = n21770 & n38601 ;
  assign n38604 = ~n21734 & n38603 ;
  assign n38605 = ~n38602 & ~n38604 ;
  assign n38606 = n23412 & n38605 ;
  assign n38607 = ~n38600 & n38606 ;
  assign n38608 = ~n38598 & ~n38607 ;
  assign n38609 = \pi0790  & ~n38608 ;
  assign n38610 = ~\pi0188  & ~\pi0705  ;
  assign n38611 = ~\pi0038  & n38610 ;
  assign n38612 = n21743 & n38611 ;
  assign n38613 = ~n21734 & n38612 ;
  assign n38614 = \pi0038  & n38610 ;
  assign n38615 = ~n22123 & n38614 ;
  assign n38616 = n6861 & ~n38615 ;
  assign n38617 = ~n38613 & n38616 ;
  assign n38618 = ~n38522 & ~n38617 ;
  assign n38619 = ~\pi0188  & ~n22017 ;
  assign n38620 = ~n21994 & n38619 ;
  assign n38621 = ~\pi0038  & ~\pi0188  ;
  assign n38622 = ~n22109 & ~n38621 ;
  assign n38623 = ~n38620 & ~n38622 ;
  assign n38624 = ~\pi0188  & ~n21757 ;
  assign n38625 = n22117 & ~n38624 ;
  assign n38626 = \pi0705  & ~n38522 ;
  assign n38627 = ~n38625 & n38626 ;
  assign n38628 = ~n38623 & n38627 ;
  assign n38629 = ~n38618 & ~n38628 ;
  assign n38630 = \pi0625  & ~n38629 ;
  assign n38631 = ~\pi0188  & ~\pi0625  ;
  assign n38632 = n21768 & n38631 ;
  assign n38633 = n21770 & n38631 ;
  assign n38634 = ~n21734 & n38633 ;
  assign n38635 = ~n38632 & ~n38634 ;
  assign n38636 = \pi1153  & n38635 ;
  assign n38637 = ~n38630 & n38636 ;
  assign n38638 = ~\pi0625  & ~n38629 ;
  assign n38639 = ~\pi0188  & \pi0625  ;
  assign n38640 = n21768 & n38639 ;
  assign n38641 = n21770 & n38639 ;
  assign n38642 = ~n21734 & n38641 ;
  assign n38643 = ~n38640 & ~n38642 ;
  assign n38644 = ~\pi1153  & n38643 ;
  assign n38645 = ~n38638 & n38644 ;
  assign n38646 = ~n38637 & ~n38645 ;
  assign n38647 = n22148 & ~n38646 ;
  assign n38648 = n22151 & n38629 ;
  assign n38649 = n22147 & n38513 ;
  assign n38650 = ~n22155 & ~n38649 ;
  assign n38651 = ~n38648 & n38650 ;
  assign n38652 = ~n38647 & n38651 ;
  assign n38653 = n22155 & ~n38513 ;
  assign n38654 = n22162 & ~n38653 ;
  assign n38655 = ~n38652 & n38654 ;
  assign n38656 = ~n22162 & n38513 ;
  assign n38657 = ~\pi0647  & ~n38656 ;
  assign n38658 = ~n38655 & n38657 ;
  assign n38659 = ~n22913 & ~n38658 ;
  assign n38660 = n21768 & n38365 ;
  assign n38661 = n21770 & n38365 ;
  assign n38662 = ~n21734 & n38661 ;
  assign n38663 = ~n38660 & ~n38662 ;
  assign n38664 = ~\pi1157  & n38663 ;
  assign n38665 = n38659 & n38664 ;
  assign n38666 = \pi0628  & ~n38656 ;
  assign n38667 = ~n38655 & n38666 ;
  assign n38668 = ~\pi0188  & ~\pi0628  ;
  assign n38669 = n21768 & n38668 ;
  assign n38670 = n21770 & n38668 ;
  assign n38671 = ~n21734 & n38670 ;
  assign n38672 = ~n38669 & ~n38671 ;
  assign n38673 = \pi1156  & n38672 ;
  assign n38674 = ~n38667 & n38673 ;
  assign n38675 = ~\pi0628  & ~n38656 ;
  assign n38676 = ~n38655 & n38675 ;
  assign n38677 = ~\pi0188  & \pi0628  ;
  assign n38678 = n21768 & n38677 ;
  assign n38679 = n21770 & n38677 ;
  assign n38680 = ~n21734 & n38679 ;
  assign n38681 = ~n38678 & ~n38680 ;
  assign n38682 = ~\pi1156  & n38681 ;
  assign n38683 = ~n38676 & n38682 ;
  assign n38684 = ~n38674 & ~n38683 ;
  assign n38685 = \pi0792  & n38664 ;
  assign n38686 = ~n38684 & n38685 ;
  assign n38687 = ~n38665 & ~n38686 ;
  assign n38688 = \pi0787  & n38687 ;
  assign n38689 = \pi0647  & ~n38656 ;
  assign n38690 = ~n38655 & n38689 ;
  assign n38691 = ~n22956 & ~n38690 ;
  assign n38692 = n21768 & n38369 ;
  assign n38693 = n21770 & n38369 ;
  assign n38694 = ~n21734 & n38693 ;
  assign n38695 = ~n38692 & ~n38694 ;
  assign n38696 = \pi1157  & n38695 ;
  assign n38697 = n38691 & n38696 ;
  assign n38698 = \pi0792  & n38696 ;
  assign n38699 = ~n38684 & n38698 ;
  assign n38700 = ~n38697 & ~n38699 ;
  assign n38701 = n38688 & n38700 ;
  assign n38702 = ~\pi0787  & ~n38656 ;
  assign n38703 = ~n38655 & n38702 ;
  assign n38704 = ~n33084 & ~n38703 ;
  assign n38705 = n23518 & n38704 ;
  assign n38706 = n37542 & ~n38684 ;
  assign n38707 = ~n38705 & ~n38706 ;
  assign n38708 = \pi0790  & ~n38707 ;
  assign n38709 = ~n38701 & n38708 ;
  assign n38710 = ~n38609 & ~n38709 ;
  assign n38711 = n9948 & n38710 ;
  assign n38712 = n24691 & ~n38514 ;
  assign n38713 = ~n38558 & n38712 ;
  assign n38714 = \pi0789  & n38712 ;
  assign n38715 = ~n38585 & n38714 ;
  assign n38716 = ~n38713 & ~n38715 ;
  assign n38717 = ~\pi0629  & n38673 ;
  assign n38718 = ~n38667 & n38717 ;
  assign n38719 = \pi0629  & n38682 ;
  assign n38720 = ~n38676 & n38719 ;
  assign n38721 = ~n38718 & ~n38720 ;
  assign n38722 = n38716 & n38721 ;
  assign n38723 = n24724 & ~n38722 ;
  assign n38724 = \pi0789  & ~n38585 ;
  assign n38725 = n30606 & ~n38557 ;
  assign n38726 = ~n38724 & n38725 ;
  assign n38727 = ~n22849 & n38513 ;
  assign n38728 = \pi0641  & n38727 ;
  assign n38729 = ~n38648 & ~n38649 ;
  assign n38730 = ~n38647 & n38729 ;
  assign n38731 = n33656 & ~n38730 ;
  assign n38732 = ~n38728 & ~n38731 ;
  assign n38733 = ~\pi0641  & n38513 ;
  assign n38734 = n20776 & ~n38733 ;
  assign n38735 = n38732 & n38734 ;
  assign n38736 = ~n38726 & ~n38735 ;
  assign n38737 = ~\pi0641  & n38727 ;
  assign n38738 = n33649 & ~n38730 ;
  assign n38739 = ~n38737 & ~n38738 ;
  assign n38740 = \pi0641  & n38513 ;
  assign n38741 = n20777 & ~n38740 ;
  assign n38742 = n38739 & n38741 ;
  assign n38743 = ~n23856 & ~n38742 ;
  assign n38744 = ~n21067 & n38743 ;
  assign n38745 = n38736 & n38744 ;
  assign n38746 = ~n38126 & ~n38745 ;
  assign n38747 = ~n38723 & n38746 ;
  assign n38748 = ~n22734 & ~n38631 ;
  assign n38749 = ~n6861 & ~n38748 ;
  assign n38750 = ~n29124 & ~n38748 ;
  assign n38751 = n38535 & n38750 ;
  assign n38752 = ~n38749 & ~n38751 ;
  assign n38753 = \pi1153  & n38752 ;
  assign n38754 = \pi0608  & ~n38644 ;
  assign n38755 = n22740 & ~n38629 ;
  assign n38756 = ~n38754 & ~n38755 ;
  assign n38757 = ~n38753 & ~n38756 ;
  assign n38758 = \pi0038  & \pi0188  ;
  assign n38759 = ~n22708 & n38758 ;
  assign n38760 = ~\pi0038  & \pi0188  ;
  assign n38761 = ~n38759 & ~n38760 ;
  assign n38762 = ~n23558 & ~n38759 ;
  assign n38763 = n23557 & n38762 ;
  assign n38764 = ~n38761 & ~n38763 ;
  assign n38765 = ~\pi0188  & n23548 ;
  assign n38766 = ~n25191 & n38765 ;
  assign n38767 = ~n25190 & n38766 ;
  assign n38768 = \pi0705  & ~\pi0768  ;
  assign n38769 = ~n38767 & n38768 ;
  assign n38770 = ~n38764 & n38769 ;
  assign n38771 = ~\pi0188  & ~n25209 ;
  assign n38772 = ~n25204 & n38771 ;
  assign n38773 = n23575 & n38760 ;
  assign n38774 = n23572 & n38773 ;
  assign n38775 = ~n25217 & ~n38774 ;
  assign n38776 = ~n38772 & n38775 ;
  assign n38777 = \pi0705  & \pi0768  ;
  assign n38778 = ~n38776 & n38777 ;
  assign n38779 = ~n38770 & ~n38778 ;
  assign n38780 = ~\pi0705  & ~n38530 ;
  assign n38781 = ~n38534 & n38780 ;
  assign n38782 = ~n29124 & n38781 ;
  assign n38783 = n6861 & ~n38782 ;
  assign n38784 = n38779 & n38783 ;
  assign n38785 = ~n22727 & ~n38639 ;
  assign n38786 = ~n38756 & ~n38785 ;
  assign n38787 = ~n38784 & n38786 ;
  assign n38788 = ~n38757 & ~n38787 ;
  assign n38789 = n23613 & ~n38788 ;
  assign n38790 = ~n6861 & ~n38785 ;
  assign n38791 = ~n29124 & ~n38785 ;
  assign n38792 = n38535 & n38791 ;
  assign n38793 = ~n38790 & ~n38792 ;
  assign n38794 = n38748 & n38793 ;
  assign n38795 = n38783 & n38793 ;
  assign n38796 = n38779 & n38795 ;
  assign n38797 = ~n38794 & ~n38796 ;
  assign n38798 = ~\pi1153  & ~n38797 ;
  assign n38799 = ~\pi0608  & ~n38636 ;
  assign n38800 = n22755 & ~n38629 ;
  assign n38801 = ~n38799 & ~n38800 ;
  assign n38802 = n23613 & ~n38801 ;
  assign n38803 = ~n38798 & n38802 ;
  assign n38804 = ~n38789 & ~n38803 ;
  assign n38805 = \pi0778  & ~n38646 ;
  assign n38806 = ~\pi0778  & n38629 ;
  assign n38807 = \pi0609  & ~n38806 ;
  assign n38808 = ~n38805 & n38807 ;
  assign n38809 = ~\pi0188  & ~\pi0778  ;
  assign n38810 = ~n23622 & ~n38809 ;
  assign n38811 = ~\pi0609  & ~n38810 ;
  assign n38812 = ~n38784 & n38811 ;
  assign n38813 = ~\pi1155  & ~n38812 ;
  assign n38814 = ~n38808 & n38813 ;
  assign n38815 = n38804 & n38814 ;
  assign n38816 = ~n20985 & n38522 ;
  assign n38817 = ~n26645 & ~n38816 ;
  assign n38818 = ~n29124 & ~n38816 ;
  assign n38819 = n38535 & n38818 ;
  assign n38820 = ~n38817 & ~n38819 ;
  assign n38821 = n21774 & n38820 ;
  assign n38822 = n26653 & n38513 ;
  assign n38823 = ~\pi0660  & ~n38822 ;
  assign n38824 = ~n38821 & n38823 ;
  assign n38825 = ~n38815 & n38824 ;
  assign n38826 = n20999 & n38820 ;
  assign n38827 = ~n32768 & n38513 ;
  assign n38828 = \pi0660  & ~n38827 ;
  assign n38829 = ~n38826 & n38828 ;
  assign n38830 = \pi0785  & ~n38829 ;
  assign n38831 = n23638 & ~n38788 ;
  assign n38832 = n23638 & ~n38801 ;
  assign n38833 = ~n38798 & n38832 ;
  assign n38834 = ~n38831 & ~n38833 ;
  assign n38835 = ~\pi0609  & ~n38806 ;
  assign n38836 = \pi1155  & ~n38835 ;
  assign n38837 = n22722 & ~n38646 ;
  assign n38838 = ~n38836 & ~n38837 ;
  assign n38839 = \pi0609  & ~n38810 ;
  assign n38840 = ~n38784 & n38839 ;
  assign n38841 = \pi0785  & ~n38840 ;
  assign n38842 = ~n38838 & n38841 ;
  assign n38843 = n38834 & n38842 ;
  assign n38844 = ~n38830 & ~n38843 ;
  assign n38845 = ~n38825 & ~n38844 ;
  assign n38846 = n21019 & ~n38520 ;
  assign n38847 = n21020 & n38550 ;
  assign n38848 = ~n33630 & ~n38847 ;
  assign n38849 = ~n38846 & ~n38848 ;
  assign n38850 = n20828 & n38579 ;
  assign n38851 = ~\pi0619  & n38850 ;
  assign n38852 = ~n38555 & n38850 ;
  assign n38853 = ~n38553 & n38852 ;
  assign n38854 = ~n38851 & ~n38853 ;
  assign n38855 = n32121 & ~n38571 ;
  assign n38856 = n32125 & ~n38855 ;
  assign n38857 = n38854 & ~n38856 ;
  assign n38858 = \pi0789  & ~n38857 ;
  assign n38859 = \pi0778  & ~n38788 ;
  assign n38860 = \pi0778  & ~n38801 ;
  assign n38861 = ~n38798 & n38860 ;
  assign n38862 = ~n38859 & ~n38861 ;
  assign n38863 = ~\pi0785  & n38810 ;
  assign n38864 = ~\pi0785  & n38783 ;
  assign n38865 = n38779 & n38864 ;
  assign n38866 = ~n38863 & ~n38865 ;
  assign n38867 = n38862 & ~n38866 ;
  assign n38868 = ~n38858 & ~n38867 ;
  assign n38869 = ~n38849 & n38868 ;
  assign n38870 = ~n38845 & n38869 ;
  assign n38871 = ~\pi1159  & ~n38653 ;
  assign n38872 = ~n38652 & n38871 ;
  assign n38873 = ~n22872 & ~n38872 ;
  assign n38874 = ~\pi0648  & n38584 ;
  assign n38875 = n38873 & n38874 ;
  assign n38876 = \pi1159  & ~n38653 ;
  assign n38877 = ~n38652 & n38876 ;
  assign n38878 = n37561 & ~n38574 ;
  assign n38879 = ~n38877 & n38878 ;
  assign n38880 = ~n38875 & ~n38879 ;
  assign n38881 = \pi0789  & ~n38880 ;
  assign n38882 = ~\pi0618  & ~n38649 ;
  assign n38883 = ~n38648 & n38882 ;
  assign n38884 = ~n38647 & n38883 ;
  assign n38885 = \pi1154  & ~n38884 ;
  assign n38886 = \pi0627  & ~n38520 ;
  assign n38887 = \pi0627  & n38540 ;
  assign n38888 = ~n38538 & n38887 ;
  assign n38889 = ~n38886 & ~n38888 ;
  assign n38890 = ~n38885 & ~n38889 ;
  assign n38891 = \pi0618  & ~n38649 ;
  assign n38892 = ~n38648 & n38891 ;
  assign n38893 = ~n38647 & n38892 ;
  assign n38894 = ~\pi1154  & ~n38893 ;
  assign n38895 = ~\pi0627  & ~n38551 ;
  assign n38896 = ~\pi0627  & n38544 ;
  assign n38897 = ~n38538 & n38896 ;
  assign n38898 = ~n38895 & ~n38897 ;
  assign n38899 = ~n38894 & ~n38898 ;
  assign n38900 = ~n38890 & ~n38899 ;
  assign n38901 = ~n38858 & ~n38900 ;
  assign n38902 = \pi0781  & n38901 ;
  assign n38903 = ~n38881 & ~n38902 ;
  assign n38904 = ~n38870 & n38903 ;
  assign n38905 = ~n21038 & ~n38723 ;
  assign n38906 = ~n38904 & n38905 ;
  assign n38907 = ~n38747 & ~n38906 ;
  assign n38908 = ~n24761 & n38907 ;
  assign n38909 = ~n30376 & n38513 ;
  assign n38910 = ~n20910 & n38909 ;
  assign n38911 = ~\pi0789  & ~n38557 ;
  assign n38912 = ~n38557 & ~n38574 ;
  assign n38913 = n38584 & n38912 ;
  assign n38914 = ~n38911 & ~n38913 ;
  assign n38915 = n33670 & n38914 ;
  assign n38916 = ~n38910 & ~n38915 ;
  assign n38917 = ~\pi0630  & n38916 ;
  assign n38918 = n38700 & n38917 ;
  assign n38919 = \pi0630  & n38916 ;
  assign n38920 = n38687 & n38919 ;
  assign n38921 = ~n38918 & ~n38920 ;
  assign n38922 = n32298 & n38921 ;
  assign n38923 = ~n38506 & ~n38922 ;
  assign n38924 = ~n38908 & n38923 ;
  assign n38925 = n38711 & n38924 ;
  assign n38926 = ~n38509 & ~n38925 ;
  assign n38927 = \pi0189  & ~n1689 ;
  assign n38928 = \pi0727  & n1689 ;
  assign n38929 = n20855 & n38928 ;
  assign n38930 = ~n38927 & ~n38929 ;
  assign n38931 = ~\pi0778  & ~n38930 ;
  assign n38932 = n23846 & n38931 ;
  assign n38933 = \pi0625  & \pi0727  ;
  assign n38934 = n1689 & n38933 ;
  assign n38935 = n20855 & n38934 ;
  assign n38936 = ~n38927 & ~n38935 ;
  assign n38937 = \pi1153  & ~n38936 ;
  assign n38938 = ~\pi1153  & ~n38935 ;
  assign n38939 = ~n38930 & n38938 ;
  assign n38940 = ~n38937 & ~n38939 ;
  assign n38941 = n30727 & ~n38940 ;
  assign n38942 = ~n38932 & ~n38941 ;
  assign n38943 = \pi0772  & n1689 ;
  assign n38944 = n20784 & n38943 ;
  assign n38945 = n30730 & n38944 ;
  assign n38946 = n21777 & n38945 ;
  assign n38947 = \pi0189  & ~\pi1154  ;
  assign n38948 = ~n1689 & n38947 ;
  assign n38949 = ~n38946 & ~n38948 ;
  assign n38950 = \pi0618  & ~n38949 ;
  assign n38951 = n30737 & n38927 ;
  assign n38952 = n30739 & n38944 ;
  assign n38953 = n21777 & n38952 ;
  assign n38954 = ~n38951 & ~n38953 ;
  assign n38955 = ~n38950 & n38954 ;
  assign n38956 = n38942 & n38955 ;
  assign n38957 = \pi0781  & ~n38956 ;
  assign n38958 = ~n26119 & ~n38940 ;
  assign n38959 = n26125 & ~n38930 ;
  assign n38960 = ~n20866 & n38927 ;
  assign n38961 = ~n20866 & n38944 ;
  assign n38962 = n26128 & n38961 ;
  assign n38963 = ~n38960 & ~n38962 ;
  assign n38964 = ~n38959 & n38963 ;
  assign n38965 = ~n38958 & n38964 ;
  assign n38966 = n21023 & ~n38965 ;
  assign n38967 = \pi0608  & n38935 ;
  assign n38968 = \pi0608  & ~n38927 ;
  assign n38969 = ~n38929 & n38968 ;
  assign n38970 = ~n38967 & ~n38969 ;
  assign n38971 = n26147 & n38929 ;
  assign n38972 = ~\pi1153  & ~n38971 ;
  assign n38973 = n38970 & n38972 ;
  assign n38974 = ~\pi0625  & ~n38944 ;
  assign n38975 = n30763 & ~n38974 ;
  assign n38976 = \pi0778  & ~n38927 ;
  assign n38977 = ~n38935 & n38976 ;
  assign n38978 = ~n30765 & ~n38977 ;
  assign n38979 = ~n38975 & ~n38978 ;
  assign n38980 = ~n38973 & n38979 ;
  assign n38981 = n20784 & ~n38927 ;
  assign n38982 = ~n20985 & n38981 ;
  assign n38983 = ~n38930 & ~n38982 ;
  assign n38984 = ~n38944 & ~n38983 ;
  assign n38985 = n30774 & ~n38984 ;
  assign n38986 = ~n38980 & n38985 ;
  assign n38987 = ~n21034 & ~n38986 ;
  assign n38988 = ~n38966 & n38987 ;
  assign n38989 = ~n38957 & n38988 ;
  assign n38990 = n30780 & ~n38940 ;
  assign n38991 = n23380 & n38931 ;
  assign n38992 = \pi0789  & ~n38927 ;
  assign n38993 = ~n29814 & n38992 ;
  assign n38994 = ~n38991 & n38993 ;
  assign n38995 = ~n38990 & n38994 ;
  assign n38996 = n26177 & n38944 ;
  assign n38997 = ~n20876 & n38992 ;
  assign n38998 = ~n38996 & n38997 ;
  assign n38999 = ~n21038 & ~n38998 ;
  assign n39000 = ~n38995 & n38999 ;
  assign n39001 = ~n38989 & n39000 ;
  assign n39002 = n30793 & n38991 ;
  assign n39003 = n30795 & ~n38940 ;
  assign n39004 = ~n39002 & ~n39003 ;
  assign n39005 = n20777 & n38927 ;
  assign n39006 = ~\pi0641  & ~n38927 ;
  assign n39007 = ~n22899 & ~n39006 ;
  assign n39008 = \pi0603  & \pi0626  ;
  assign n39009 = ~n20783 & n39008 ;
  assign n39010 = n38943 & n39009 ;
  assign n39011 = ~n22899 & n39010 ;
  assign n39012 = n23832 & n39011 ;
  assign n39013 = ~n39007 & ~n39012 ;
  assign n39014 = ~n39005 & n39013 ;
  assign n39015 = n39004 & n39014 ;
  assign n39016 = n30807 & n38991 ;
  assign n39017 = n30809 & ~n38940 ;
  assign n39018 = ~n39016 & ~n39017 ;
  assign n39019 = n20776 & n38927 ;
  assign n39020 = \pi0641  & ~n38927 ;
  assign n39021 = ~n22884 & ~n39020 ;
  assign n39022 = n26205 & n38943 ;
  assign n39023 = ~n22884 & n39022 ;
  assign n39024 = n23832 & n39023 ;
  assign n39025 = ~n39021 & ~n39024 ;
  assign n39026 = ~n39019 & n39025 ;
  assign n39027 = n39018 & n39026 ;
  assign n39028 = ~n39015 & ~n39027 ;
  assign n39029 = \pi0788  & n39028 ;
  assign n39030 = n30823 & ~n39029 ;
  assign n39031 = ~n39001 & n39030 ;
  assign n39032 = ~n23880 & n38944 ;
  assign n39033 = ~n20846 & n39032 ;
  assign n39034 = n23832 & n39033 ;
  assign n39035 = n21064 & ~n39034 ;
  assign n39036 = n20897 & ~n23920 ;
  assign n39037 = n26065 & ~n38940 ;
  assign n39038 = n23885 & n38931 ;
  assign n39039 = n20897 & ~n39038 ;
  assign n39040 = ~n39037 & n39039 ;
  assign n39041 = ~n39036 & ~n39040 ;
  assign n39042 = ~n39035 & n39041 ;
  assign n39043 = ~n30712 & ~n39038 ;
  assign n39044 = ~n39037 & n39043 ;
  assign n39045 = ~n30713 & ~n39044 ;
  assign n39046 = n30717 & n39032 ;
  assign n39047 = n23832 & n39046 ;
  assign n39048 = \pi1157  & ~n39047 ;
  assign n39049 = ~n39045 & n39048 ;
  assign n39050 = n39042 & ~n39049 ;
  assign n39051 = \pi0787  & ~n38927 ;
  assign n39052 = ~n39050 & n39051 ;
  assign n39053 = n30688 & n38944 ;
  assign n39054 = n23832 & n39053 ;
  assign n39055 = n20886 & ~n39054 ;
  assign n39056 = n24724 & n39055 ;
  assign n39057 = ~n39037 & ~n39038 ;
  assign n39058 = ~\pi0629  & \pi1156  ;
  assign n39059 = ~n39054 & n39058 ;
  assign n39060 = n24724 & n39059 ;
  assign n39061 = n39057 & n39060 ;
  assign n39062 = ~n39056 & ~n39061 ;
  assign n39063 = ~\pi0628  & ~n39057 ;
  assign n39064 = ~\pi0629  & n39032 ;
  assign n39065 = n23832 & n39064 ;
  assign n39066 = ~n25956 & ~n39065 ;
  assign n39067 = n30701 & n39066 ;
  assign n39068 = ~n39063 & n39067 ;
  assign n39069 = n39062 & ~n39068 ;
  assign n39070 = ~n38927 & ~n39069 ;
  assign n39071 = ~n24761 & ~n39070 ;
  assign n39072 = ~n39052 & n39071 ;
  assign n39073 = ~n39031 & n39072 ;
  assign n39074 = n26069 & ~n39057 ;
  assign n39075 = n26080 & n38927 ;
  assign n39076 = n26082 & n39034 ;
  assign n39077 = ~n39075 & ~n39076 ;
  assign n39078 = n26076 & n38927 ;
  assign n39079 = n26078 & n39034 ;
  assign n39080 = ~n39078 & ~n39079 ;
  assign n39081 = n39077 & n39080 ;
  assign n39082 = ~n39074 & n39081 ;
  assign n39083 = \pi0790  & ~n39082 ;
  assign n39084 = \pi0832  & ~n39083 ;
  assign n39085 = ~n39073 & n39084 ;
  assign n39086 = ~\pi0189  & ~n6848 ;
  assign n39087 = ~\pi0057  & ~n39086 ;
  assign n39088 = \pi0189  & n21768 ;
  assign n39089 = \pi0189  & n21770 ;
  assign n39090 = ~n21734 & n39089 ;
  assign n39091 = ~n39088 & ~n39090 ;
  assign n39092 = ~\pi0074  & \pi0727  ;
  assign n39093 = ~\pi0100  & n39092 ;
  assign n39094 = n1287 & n39093 ;
  assign n39095 = n39091 & ~n39094 ;
  assign n39096 = ~\pi0189  & ~n22107 ;
  assign n39097 = n22089 & n39096 ;
  assign n39098 = ~\pi0038  & ~n39097 ;
  assign n39099 = \pi0039  & \pi0189  ;
  assign n39100 = ~n21993 & n39099 ;
  assign n39101 = \pi0189  & n22017 ;
  assign n39102 = ~n39100 & ~n39101 ;
  assign n39103 = n39098 & n39102 ;
  assign n39104 = ~\pi0189  & ~n21757 ;
  assign n39105 = n25669 & ~n39104 ;
  assign n39106 = n39094 & ~n39105 ;
  assign n39107 = ~n39103 & n39106 ;
  assign n39108 = ~n39095 & ~n39107 ;
  assign n39109 = ~\pi0778  & n39108 ;
  assign n39110 = n23380 & ~n39109 ;
  assign n39111 = ~n23380 & n39091 ;
  assign n39112 = ~n22160 & ~n39111 ;
  assign n39113 = ~n39110 & n39112 ;
  assign n39114 = \pi0625  & ~n39108 ;
  assign n39115 = ~\pi0625  & n39091 ;
  assign n39116 = \pi1153  & ~n39115 ;
  assign n39117 = ~n39114 & n39116 ;
  assign n39118 = ~\pi0625  & ~n39108 ;
  assign n39119 = \pi0625  & n39091 ;
  assign n39120 = ~\pi1153  & ~n39119 ;
  assign n39121 = ~n39118 & n39120 ;
  assign n39122 = ~n39117 & ~n39121 ;
  assign n39123 = \pi0778  & n39112 ;
  assign n39124 = ~n39122 & n39123 ;
  assign n39125 = ~n39113 & ~n39124 ;
  assign n39126 = n22160 & ~n39091 ;
  assign n39127 = \pi0628  & ~n22161 ;
  assign n39128 = ~n39126 & n39127 ;
  assign n39129 = n39125 & n39128 ;
  assign n39130 = n39091 & ~n39127 ;
  assign n39131 = n20843 & ~n39130 ;
  assign n39132 = ~n39129 & n39131 ;
  assign n39133 = \pi0792  & n39132 ;
  assign n39134 = ~n22162 & n39091 ;
  assign n39135 = ~\pi0628  & n39134 ;
  assign n39136 = ~n39110 & ~n39111 ;
  assign n39137 = \pi0778  & ~n39111 ;
  assign n39138 = ~n39122 & n39137 ;
  assign n39139 = ~n39136 & ~n39138 ;
  assign n39140 = n30317 & n39139 ;
  assign n39141 = ~n39135 & ~n39140 ;
  assign n39142 = \pi0628  & n39091 ;
  assign n39143 = n20844 & ~n39142 ;
  assign n39144 = \pi0792  & n39143 ;
  assign n39145 = n39141 & n39144 ;
  assign n39146 = ~n39133 & ~n39145 ;
  assign n39147 = ~n21067 & ~n39146 ;
  assign n39148 = n21776 & n39091 ;
  assign n39149 = ~\pi0781  & ~n39148 ;
  assign n39150 = ~\pi0619  & ~n39149 ;
  assign n39151 = \pi0299  & ~\pi0772  ;
  assign n39152 = ~n21205 & n39151 ;
  assign n39153 = ~n21238 & n39152 ;
  assign n39154 = ~n21740 & n29065 ;
  assign n39155 = ~n21738 & n39154 ;
  assign n39156 = ~n39153 & ~n39155 ;
  assign n39157 = ~\pi0039  & n39156 ;
  assign n39158 = ~\pi0299  & \pi0772  ;
  assign n39159 = ~n25554 & n39158 ;
  assign n39160 = ~n39157 & ~n39159 ;
  assign n39161 = \pi0772  & ~n39159 ;
  assign n39162 = n21272 & n39161 ;
  assign n39163 = ~n39160 & ~n39162 ;
  assign n39164 = ~\pi0772  & ~n25542 ;
  assign n39165 = \pi0299  & \pi0772  ;
  assign n39166 = ~n25557 & n39165 ;
  assign n39167 = ~n39164 & ~n39166 ;
  assign n39168 = ~n39163 & n39167 ;
  assign n39169 = ~\pi0039  & ~n39156 ;
  assign n39170 = ~\pi0039  & \pi0772  ;
  assign n39171 = n21272 & n39170 ;
  assign n39172 = ~n39169 & ~n39171 ;
  assign n39173 = ~\pi0038  & \pi0189  ;
  assign n39174 = n39172 & n39173 ;
  assign n39175 = ~n39168 & n39174 ;
  assign n39176 = ~\pi0189  & \pi0772  ;
  assign n39177 = ~\pi0038  & n39176 ;
  assign n39178 = n25023 & n39177 ;
  assign n39179 = \pi0189  & ~n6861 ;
  assign n39180 = \pi0603  & \pi0772  ;
  assign n39181 = ~n20783 & n39180 ;
  assign n39182 = n6784 & ~n39181 ;
  assign n39183 = n1266 & n39182 ;
  assign n39184 = n1689 & n39183 ;
  assign n39185 = n26939 & n39184 ;
  assign n39186 = n10323 & n39185 ;
  assign n39187 = \pi0038  & ~n39186 ;
  assign n39188 = ~n39104 & n39187 ;
  assign n39189 = ~n39179 & ~n39188 ;
  assign n39190 = ~n39178 & n39189 ;
  assign n39191 = ~n39175 & n39190 ;
  assign n39192 = ~\pi0189  & ~n6861 ;
  assign n39193 = ~n20985 & ~n39192 ;
  assign n39194 = ~n39191 & n39193 ;
  assign n39195 = n20985 & ~n39091 ;
  assign n39196 = ~n25588 & ~n39195 ;
  assign n39197 = ~\pi0619  & n39196 ;
  assign n39198 = ~n39194 & n39197 ;
  assign n39199 = ~n39150 & ~n39198 ;
  assign n39200 = \pi0189  & ~\pi1159  ;
  assign n39201 = n21768 & n39200 ;
  assign n39202 = n21770 & n39200 ;
  assign n39203 = ~n21734 & n39202 ;
  assign n39204 = ~n39201 & ~n39203 ;
  assign n39205 = ~n22872 & n39204 ;
  assign n39206 = n39199 & ~n39205 ;
  assign n39207 = \pi0189  & ~n20811 ;
  assign n39208 = n21768 & n39207 ;
  assign n39209 = n21770 & n39207 ;
  assign n39210 = ~n21734 & n39209 ;
  assign n39211 = ~n39208 & ~n39210 ;
  assign n39212 = n20811 & ~n39148 ;
  assign n39213 = n39211 & ~n39212 ;
  assign n39214 = n39196 & n39211 ;
  assign n39215 = ~n39194 & n39214 ;
  assign n39216 = ~n39213 & ~n39215 ;
  assign n39217 = \pi0781  & ~n39205 ;
  assign n39218 = n39216 & n39217 ;
  assign n39219 = ~n39206 & ~n39218 ;
  assign n39220 = \pi0619  & ~n39149 ;
  assign n39221 = \pi0619  & n39196 ;
  assign n39222 = ~n39194 & n39221 ;
  assign n39223 = ~n39220 & ~n39222 ;
  assign n39224 = \pi0189  & \pi1159  ;
  assign n39225 = n21768 & n39224 ;
  assign n39226 = n21770 & n39224 ;
  assign n39227 = ~n21734 & n39226 ;
  assign n39228 = ~n39225 & ~n39227 ;
  assign n39229 = ~n20830 & n39228 ;
  assign n39230 = n39223 & ~n39229 ;
  assign n39231 = \pi0781  & ~n39229 ;
  assign n39232 = n39216 & n39231 ;
  assign n39233 = ~n39230 & ~n39232 ;
  assign n39234 = n39219 & n39233 ;
  assign n39235 = \pi0789  & ~n23880 ;
  assign n39236 = ~n39234 & n39235 ;
  assign n39237 = ~n39194 & n39196 ;
  assign n39238 = ~\pi0789  & n39149 ;
  assign n39239 = ~n39237 & n39238 ;
  assign n39240 = ~n23880 & n39239 ;
  assign n39241 = n21806 & ~n23880 ;
  assign n39242 = n39216 & n39241 ;
  assign n39243 = ~n39240 & ~n39242 ;
  assign n39244 = n23880 & ~n39091 ;
  assign n39245 = n39243 & ~n39244 ;
  assign n39246 = ~n39236 & n39245 ;
  assign n39247 = n20944 & n22166 ;
  assign n39248 = n22932 & n26218 ;
  assign n39249 = ~n39247 & ~n39248 ;
  assign n39250 = ~n21067 & ~n39249 ;
  assign n39251 = ~n39246 & n39250 ;
  assign n39252 = ~n39147 & ~n39251 ;
  assign n39253 = n20871 & n39216 ;
  assign n39254 = ~n22147 & ~n39109 ;
  assign n39255 = n23667 & ~n39091 ;
  assign n39256 = ~n23846 & ~n39255 ;
  assign n39257 = ~n39254 & ~n39256 ;
  assign n39258 = \pi0778  & ~n39256 ;
  assign n39259 = ~n39122 & n39258 ;
  assign n39260 = ~n39257 & ~n39259 ;
  assign n39261 = ~n39253 & n39260 ;
  assign n39262 = \pi0781  & ~n39261 ;
  assign n39263 = ~n21022 & ~n39262 ;
  assign n39264 = ~n39189 & ~n39192 ;
  assign n39265 = \pi0189  & ~\pi0299  ;
  assign n39266 = n22407 & n39265 ;
  assign n39267 = \pi0189  & \pi0299  ;
  assign n39268 = n22291 & n39267 ;
  assign n39269 = ~n39266 & ~n39268 ;
  assign n39270 = ~\pi0189  & ~n22379 ;
  assign n39271 = ~n30442 & n39270 ;
  assign n39272 = ~\pi0772  & ~n39271 ;
  assign n39273 = n39269 & n39272 ;
  assign n39274 = n22601 & n39265 ;
  assign n39275 = n22630 & n39267 ;
  assign n39276 = \pi0772  & ~n39275 ;
  assign n39277 = ~n39274 & n39276 ;
  assign n39278 = \pi0039  & ~n39277 ;
  assign n39279 = ~\pi0189  & n22468 ;
  assign n39280 = ~n30448 & n39279 ;
  assign n39281 = \pi0039  & n39280 ;
  assign n39282 = ~n30447 & n39281 ;
  assign n39283 = ~n39278 & ~n39282 ;
  assign n39284 = ~n39273 & ~n39283 ;
  assign n39285 = \pi0189  & n22643 ;
  assign n39286 = ~n22652 & n39285 ;
  assign n39287 = ~\pi0189  & ~\pi0299  ;
  assign n39288 = n22676 & n39287 ;
  assign n39289 = ~\pi0189  & \pi0299  ;
  assign n39290 = ~n22657 & n39289 ;
  assign n39291 = ~n22660 & n39290 ;
  assign n39292 = n22664 & n39291 ;
  assign n39293 = ~\pi0772  & ~n39292 ;
  assign n39294 = ~n39288 & n39293 ;
  assign n39295 = ~n39286 & n39294 ;
  assign n39296 = \pi0772  & n21272 ;
  assign n39297 = n22006 & n39267 ;
  assign n39298 = n22649 & n39265 ;
  assign n39299 = ~n39297 & ~n39298 ;
  assign n39300 = n39296 & ~n39299 ;
  assign n39301 = n22693 & n39176 ;
  assign n39302 = ~\pi0039  & ~n39301 ;
  assign n39303 = ~n39300 & n39302 ;
  assign n39304 = ~n39295 & n39303 ;
  assign n39305 = \pi0727  & ~n25217 ;
  assign n39306 = ~n39304 & n39305 ;
  assign n39307 = ~n39284 & n39306 ;
  assign n39308 = ~n30436 & ~n39307 ;
  assign n39309 = ~\pi0727  & ~n39178 ;
  assign n39310 = ~n39175 & n39309 ;
  assign n39311 = ~n39192 & ~n39310 ;
  assign n39312 = n39308 & n39311 ;
  assign n39313 = ~n39264 & ~n39312 ;
  assign n39314 = n30488 & n39091 ;
  assign n39315 = ~n30763 & ~n39314 ;
  assign n39316 = n22740 & ~n39108 ;
  assign n39317 = n39315 & ~n39316 ;
  assign n39318 = \pi0625  & ~n39317 ;
  assign n39319 = n39313 & n39318 ;
  assign n39320 = n30491 & ~n39116 ;
  assign n39321 = n39313 & n39320 ;
  assign n39322 = ~\pi1153  & ~n39192 ;
  assign n39323 = ~n39191 & n39322 ;
  assign n39324 = ~n24561 & ~n39323 ;
  assign n39325 = ~\pi0608  & ~n39116 ;
  assign n39326 = n22755 & ~n39108 ;
  assign n39327 = ~n39325 & ~n39326 ;
  assign n39328 = n39324 & ~n39327 ;
  assign n39329 = \pi1153  & ~n39192 ;
  assign n39330 = ~n39191 & n39329 ;
  assign n39331 = ~n24550 & ~n39330 ;
  assign n39332 = ~n39317 & n39331 ;
  assign n39333 = ~n39328 & ~n39332 ;
  assign n39334 = ~n39321 & n39333 ;
  assign n39335 = ~n39319 & n39334 ;
  assign n39336 = \pi0778  & ~n39335 ;
  assign n39337 = \pi0609  & ~n39109 ;
  assign n39338 = ~\pi1155  & ~n39337 ;
  assign n39339 = n24584 & ~n39122 ;
  assign n39340 = ~n39338 & ~n39339 ;
  assign n39341 = \pi0189  & ~\pi1155  ;
  assign n39342 = n21768 & n39341 ;
  assign n39343 = n21770 & n39341 ;
  assign n39344 = ~n21734 & n39343 ;
  assign n39345 = ~n39342 & ~n39344 ;
  assign n39346 = ~n20999 & n39345 ;
  assign n39347 = \pi0660  & n39346 ;
  assign n39348 = ~\pi0609  & ~n39195 ;
  assign n39349 = \pi0660  & n39348 ;
  assign n39350 = ~n39194 & n39349 ;
  assign n39351 = ~n39347 & ~n39350 ;
  assign n39352 = ~n39340 & n39351 ;
  assign n39353 = \pi0660  & n21774 ;
  assign n39354 = \pi0785  & ~n39353 ;
  assign n39355 = ~n21774 & n39354 ;
  assign n39356 = \pi0609  & ~n39195 ;
  assign n39357 = n39354 & n39356 ;
  assign n39358 = ~n39194 & n39357 ;
  assign n39359 = ~n39355 & ~n39358 ;
  assign n39360 = ~n39352 & ~n39359 ;
  assign n39361 = ~\pi0778  & n39313 ;
  assign n39362 = ~n39360 & ~n39361 ;
  assign n39363 = ~n39336 & n39362 ;
  assign n39364 = \pi0609  & n39351 ;
  assign n39365 = ~n39340 & n39364 ;
  assign n39366 = \pi0785  & n39365 ;
  assign n39367 = ~\pi0778  & n26121 ;
  assign n39368 = n39108 & n39367 ;
  assign n39369 = n31109 & ~n39122 ;
  assign n39370 = ~n39368 & ~n39369 ;
  assign n39371 = ~n39351 & n39370 ;
  assign n39372 = \pi0189  & \pi1155  ;
  assign n39373 = n21768 & n39372 ;
  assign n39374 = n21770 & n39372 ;
  assign n39375 = ~n21734 & n39374 ;
  assign n39376 = ~n39373 & ~n39375 ;
  assign n39377 = ~n21774 & n39376 ;
  assign n39378 = ~\pi0660  & n39377 ;
  assign n39379 = ~\pi0660  & n39356 ;
  assign n39380 = ~n39194 & n39379 ;
  assign n39381 = ~n39378 & ~n39380 ;
  assign n39382 = \pi0785  & n39381 ;
  assign n39383 = ~n39371 & n39382 ;
  assign n39384 = ~n39366 & ~n39383 ;
  assign n39385 = ~n39262 & n39384 ;
  assign n39386 = ~n39363 & n39385 ;
  assign n39387 = ~n39263 & ~n39386 ;
  assign n39388 = n32121 & n39204 ;
  assign n39389 = ~n32123 & ~n39388 ;
  assign n39390 = \pi0789  & n39389 ;
  assign n39391 = \pi0619  & n39204 ;
  assign n39392 = \pi0789  & ~n39391 ;
  assign n39393 = ~n39233 & n39392 ;
  assign n39394 = ~n39390 & ~n39393 ;
  assign n39395 = ~n21038 & n39394 ;
  assign n39396 = ~n39387 & n39395 ;
  assign n39397 = ~\pi1159  & ~n39139 ;
  assign n39398 = n37566 & ~n39397 ;
  assign n39399 = n39233 & n39398 ;
  assign n39400 = \pi1159  & ~n39139 ;
  assign n39401 = \pi0648  & ~n33484 ;
  assign n39402 = ~n39400 & n39401 ;
  assign n39403 = n39219 & n39402 ;
  assign n39404 = ~n39399 & ~n39403 ;
  assign n39405 = n36155 & ~n39404 ;
  assign n39406 = \pi0189  & ~\pi0641  ;
  assign n39407 = n21768 & n39406 ;
  assign n39408 = n21770 & n39406 ;
  assign n39409 = ~n21734 & n39408 ;
  assign n39410 = ~n39407 & ~n39409 ;
  assign n39411 = n20776 & n39410 ;
  assign n39412 = ~n39126 & n39411 ;
  assign n39413 = n39125 & n39412 ;
  assign n39414 = ~\pi0641  & n20776 ;
  assign n39415 = n39410 & n39414 ;
  assign n39416 = \pi0189  & \pi0641  ;
  assign n39417 = n21768 & n39416 ;
  assign n39418 = n21770 & n39416 ;
  assign n39419 = ~n21734 & n39418 ;
  assign n39420 = ~n39417 & ~n39419 ;
  assign n39421 = \pi0641  & n20777 ;
  assign n39422 = n39420 & n39421 ;
  assign n39423 = ~n39415 & ~n39422 ;
  assign n39424 = ~n39413 & n39423 ;
  assign n39425 = n20777 & n39420 ;
  assign n39426 = ~n39126 & n39425 ;
  assign n39427 = n39125 & n39426 ;
  assign n39428 = ~n23856 & ~n39427 ;
  assign n39429 = n39424 & n39428 ;
  assign n39430 = ~n26803 & ~n39429 ;
  assign n39431 = \pi0789  & ~n39234 ;
  assign n39432 = n21806 & n39216 ;
  assign n39433 = n30606 & ~n39239 ;
  assign n39434 = ~n39432 & n39433 ;
  assign n39435 = ~n26803 & n39434 ;
  assign n39436 = ~n39431 & n39435 ;
  assign n39437 = ~n39430 & ~n39436 ;
  assign n39438 = ~n21067 & n39437 ;
  assign n39439 = ~n39405 & n39438 ;
  assign n39440 = ~n39396 & n39439 ;
  assign n39441 = n39252 & ~n39440 ;
  assign n39442 = ~n24761 & ~n39441 ;
  assign n39443 = n6848 & ~n32298 ;
  assign n39444 = \pi1156  & ~n39130 ;
  assign n39445 = ~n39129 & n39444 ;
  assign n39446 = \pi0792  & n39445 ;
  assign n39447 = ~\pi1156  & ~n39142 ;
  assign n39448 = \pi0792  & n39447 ;
  assign n39449 = n39141 & n39448 ;
  assign n39450 = ~n39446 & ~n39449 ;
  assign n39451 = n22162 & n39139 ;
  assign n39452 = ~\pi0792  & ~n39134 ;
  assign n39453 = ~n39451 & n39452 ;
  assign n39454 = \pi0647  & ~n39453 ;
  assign n39455 = n39450 & n39454 ;
  assign n39456 = ~\pi0647  & n39091 ;
  assign n39457 = n20849 & ~n39456 ;
  assign n39458 = ~n39455 & n39457 ;
  assign n39459 = ~\pi0647  & ~n39453 ;
  assign n39460 = n39450 & n39459 ;
  assign n39461 = \pi0647  & n39091 ;
  assign n39462 = n20897 & ~n39461 ;
  assign n39463 = ~n39460 & n39462 ;
  assign n39464 = ~n39458 & ~n39463 ;
  assign n39465 = ~n39239 & ~n39432 ;
  assign n39466 = n30376 & n39465 ;
  assign n39467 = ~n39431 & n39466 ;
  assign n39468 = ~n30376 & n39091 ;
  assign n39469 = ~n20910 & ~n39468 ;
  assign n39470 = ~n39467 & n39469 ;
  assign n39471 = n6848 & ~n39470 ;
  assign n39472 = n39464 & n39471 ;
  assign n39473 = ~n39443 & ~n39472 ;
  assign n39474 = ~n39442 & ~n39473 ;
  assign n39475 = ~\pi1157  & ~n39461 ;
  assign n39476 = ~n39460 & n39475 ;
  assign n39477 = \pi1157  & ~n39456 ;
  assign n39478 = ~n39455 & n39477 ;
  assign n39479 = ~n39476 & ~n39478 ;
  assign n39480 = n32314 & ~n39479 ;
  assign n39481 = n39450 & ~n39453 ;
  assign n39482 = ~\pi0787  & n23313 ;
  assign n39483 = ~n39481 & n39482 ;
  assign n39484 = \pi0189  & ~\pi0715  ;
  assign n39485 = n21768 & n39484 ;
  assign n39486 = n21770 & n39484 ;
  assign n39487 = ~n21734 & n39486 ;
  assign n39488 = ~n39485 & ~n39487 ;
  assign n39489 = \pi1160  & ~n23312 ;
  assign n39490 = n39488 & n39489 ;
  assign n39491 = ~n26824 & ~n39490 ;
  assign n39492 = n21092 & ~n39244 ;
  assign n39493 = n39243 & n39492 ;
  assign n39494 = ~n39236 & n39493 ;
  assign n39495 = ~n21092 & n39091 ;
  assign n39496 = ~n39490 & ~n39495 ;
  assign n39497 = ~n39494 & n39496 ;
  assign n39498 = ~n39491 & ~n39497 ;
  assign n39499 = ~n39483 & n39498 ;
  assign n39500 = ~n39480 & n39499 ;
  assign n39501 = \pi0790  & ~n39500 ;
  assign n39502 = n32339 & ~n39479 ;
  assign n39503 = ~\pi0787  & n23312 ;
  assign n39504 = ~n39481 & n39503 ;
  assign n39505 = \pi0189  & \pi0715  ;
  assign n39506 = n21768 & n39505 ;
  assign n39507 = n21770 & n39505 ;
  assign n39508 = ~n21734 & n39507 ;
  assign n39509 = ~n39506 & ~n39508 ;
  assign n39510 = ~\pi1160  & ~n23313 ;
  assign n39511 = n39509 & n39510 ;
  assign n39512 = ~n31378 & ~n39511 ;
  assign n39513 = ~n39495 & ~n39511 ;
  assign n39514 = ~n39494 & n39513 ;
  assign n39515 = ~n39512 & ~n39514 ;
  assign n39516 = ~n39504 & n39515 ;
  assign n39517 = ~n39502 & n39516 ;
  assign n39518 = n39501 & ~n39517 ;
  assign n39519 = n39474 & ~n39518 ;
  assign n39520 = n39087 & ~n39519 ;
  assign n39521 = \pi0057  & \pi0189  ;
  assign n39522 = ~\pi0832  & ~n39521 ;
  assign n39523 = ~n39520 & n39522 ;
  assign n39524 = ~n39085 & ~n39523 ;
  assign n39525 = ~\pi0190  & \pi0788  ;
  assign n39526 = ~n1689 & n39525 ;
  assign n39527 = ~n20778 & n39526 ;
  assign n39528 = n20886 & n39527 ;
  assign n39529 = \pi0763  & n1689 ;
  assign n39530 = n20784 & n39529 ;
  assign n39531 = n22767 & n39530 ;
  assign n39532 = ~\pi0190  & ~n1689 ;
  assign n39533 = ~n39530 & ~n39532 ;
  assign n39534 = ~n20792 & ~n39533 ;
  assign n39535 = ~n39531 & n39534 ;
  assign n39536 = n20801 & ~n39535 ;
  assign n39537 = ~\pi1155  & ~n39532 ;
  assign n39538 = \pi0785  & n39537 ;
  assign n39539 = ~n39531 & n39538 ;
  assign n39540 = ~\pi0785  & ~n39532 ;
  assign n39541 = ~n39530 & n39540 ;
  assign n39542 = ~n20804 & ~n39541 ;
  assign n39543 = n29682 & n39542 ;
  assign n39544 = ~n39539 & n39543 ;
  assign n39545 = ~n39536 & n39544 ;
  assign n39546 = n30847 & n39545 ;
  assign n39547 = ~n39528 & ~n39546 ;
  assign n39548 = \pi0699  & n1689 ;
  assign n39549 = n20855 & n39548 ;
  assign n39550 = ~n39532 & ~n39549 ;
  assign n39551 = ~\pi0778  & ~n39550 ;
  assign n39552 = ~\pi0625  & \pi0699  ;
  assign n39553 = n1689 & n39552 ;
  assign n39554 = n20855 & n39553 ;
  assign n39555 = \pi1153  & n39554 ;
  assign n39556 = \pi1153  & ~n39532 ;
  assign n39557 = ~n39549 & n39556 ;
  assign n39558 = ~n39555 & ~n39557 ;
  assign n39559 = ~\pi1153  & ~n39532 ;
  assign n39560 = ~n39554 & n39559 ;
  assign n39561 = \pi0778  & ~n39560 ;
  assign n39562 = n39558 & n39561 ;
  assign n39563 = ~n39551 & ~n39562 ;
  assign n39564 = n26474 & ~n39563 ;
  assign n39565 = \pi0629  & ~n39564 ;
  assign n39566 = n39547 & n39565 ;
  assign n39567 = n20887 & n39527 ;
  assign n39568 = n32579 & n39545 ;
  assign n39569 = ~n39567 & ~n39568 ;
  assign n39570 = n26485 & ~n39563 ;
  assign n39571 = ~\pi0629  & ~n39570 ;
  assign n39572 = n39569 & n39571 ;
  assign n39573 = ~n39566 & ~n39572 ;
  assign n39574 = \pi0792  & n39573 ;
  assign n39575 = ~n21067 & ~n39574 ;
  assign n39576 = \pi0647  & ~n20890 ;
  assign n39577 = ~n20885 & n39576 ;
  assign n39578 = n20879 & n39577 ;
  assign n39579 = ~n39563 & n39578 ;
  assign n39580 = ~\pi0190  & ~\pi0647  ;
  assign n39581 = ~n1689 & n39580 ;
  assign n39582 = n20849 & ~n39581 ;
  assign n39583 = ~n39579 & n39582 ;
  assign n39584 = n26319 & ~n39563 ;
  assign n39585 = ~\pi0190  & \pi0647  ;
  assign n39586 = ~n1689 & n39585 ;
  assign n39587 = n20897 & ~n39586 ;
  assign n39588 = ~n39584 & n39587 ;
  assign n39589 = ~n39583 & ~n39588 ;
  assign n39590 = \pi0787  & ~n39589 ;
  assign n39591 = ~n20846 & n39527 ;
  assign n39592 = n30376 & n39545 ;
  assign n39593 = ~n39591 & ~n39592 ;
  assign n39594 = ~\pi0190  & \pi0792  ;
  assign n39595 = ~n1689 & n39594 ;
  assign n39596 = ~n20845 & n39595 ;
  assign n39597 = n32606 & ~n39596 ;
  assign n39598 = n39593 & n39597 ;
  assign n39599 = ~n39590 & ~n39598 ;
  assign n39600 = ~n24761 & n39599 ;
  assign n39601 = ~n39575 & n39600 ;
  assign n39602 = \pi0608  & ~n39560 ;
  assign n39603 = ~n39530 & n39556 ;
  assign n39604 = \pi0778  & ~n39603 ;
  assign n39605 = n26421 & ~n39550 ;
  assign n39606 = ~n39604 & ~n39605 ;
  assign n39607 = n39602 & ~n39606 ;
  assign n39608 = n26147 & ~n39550 ;
  assign n39609 = \pi0699  & ~n20784 ;
  assign n39610 = n22113 & n39609 ;
  assign n39611 = n39533 & ~n39610 ;
  assign n39612 = ~n39608 & ~n39611 ;
  assign n39613 = n39559 & ~n39612 ;
  assign n39614 = n26415 & n39558 ;
  assign n39615 = ~n39613 & n39614 ;
  assign n39616 = ~n39607 & ~n39615 ;
  assign n39617 = ~\pi1155  & ~n39551 ;
  assign n39618 = ~n39562 & n39617 ;
  assign n39619 = ~n20999 & ~n39618 ;
  assign n39620 = ~\pi0778  & ~n39611 ;
  assign n39621 = ~n39619 & ~n39620 ;
  assign n39622 = n39616 & n39621 ;
  assign n39623 = n29766 & ~n39551 ;
  assign n39624 = ~n39562 & n39623 ;
  assign n39625 = \pi1155  & ~n39535 ;
  assign n39626 = ~\pi0660  & ~n39625 ;
  assign n39627 = ~n39624 & n39626 ;
  assign n39628 = ~n39622 & n39627 ;
  assign n39629 = \pi0785  & ~n39628 ;
  assign n39630 = n29775 & n39542 ;
  assign n39631 = ~n39539 & n39630 ;
  assign n39632 = ~n39536 & n39631 ;
  assign n39633 = n29779 & ~n39563 ;
  assign n39634 = ~n39632 & ~n39633 ;
  assign n39635 = \pi0781  & ~n39634 ;
  assign n39636 = \pi1155  & ~n39551 ;
  assign n39637 = ~n39562 & n39636 ;
  assign n39638 = ~n21774 & ~n39637 ;
  assign n39639 = ~n39620 & ~n39638 ;
  assign n39640 = n39616 & n39639 ;
  assign n39641 = n26121 & ~n39551 ;
  assign n39642 = ~n39562 & n39641 ;
  assign n39643 = \pi0660  & ~n39537 ;
  assign n39644 = \pi0660  & n39530 ;
  assign n39645 = n22767 & n39644 ;
  assign n39646 = ~n39643 & ~n39645 ;
  assign n39647 = ~n39642 & ~n39646 ;
  assign n39648 = ~n39640 & n39647 ;
  assign n39649 = ~n39635 & ~n39648 ;
  assign n39650 = n39629 & n39649 ;
  assign n39651 = ~\pi0785  & ~n39620 ;
  assign n39652 = ~n39607 & n39651 ;
  assign n39653 = ~n39615 & n39652 ;
  assign n39654 = n21022 & ~n39653 ;
  assign n39655 = ~n39635 & ~n39654 ;
  assign n39656 = n29803 & ~n39655 ;
  assign n39657 = ~n39650 & n39656 ;
  assign n39658 = n29808 & n39542 ;
  assign n39659 = ~n39539 & n39658 ;
  assign n39660 = ~n39536 & n39659 ;
  assign n39661 = n30966 & ~n39563 ;
  assign n39662 = ~n39660 & ~n39661 ;
  assign n39663 = n36155 & ~n39662 ;
  assign n39664 = \pi0626  & ~n39545 ;
  assign n39665 = ~\pi0626  & ~n39532 ;
  assign n39666 = n20881 & ~n39665 ;
  assign n39667 = ~n39664 & n39666 ;
  assign n39668 = n26458 & ~n39563 ;
  assign n39669 = ~\pi0626  & ~n39545 ;
  assign n39670 = \pi0626  & ~n39532 ;
  assign n39671 = n20882 & ~n39670 ;
  assign n39672 = ~n39669 & n39671 ;
  assign n39673 = ~n39668 & ~n39672 ;
  assign n39674 = ~n39667 & n39673 ;
  assign n39675 = \pi0788  & ~n39674 ;
  assign n39676 = ~n39663 & ~n39675 ;
  assign n39677 = ~n39657 & n39676 ;
  assign n39678 = ~n23856 & n39600 ;
  assign n39679 = ~n39677 & n39678 ;
  assign n39680 = ~n39601 & ~n39679 ;
  assign n39681 = n30987 & ~n39593 ;
  assign n39682 = n23312 & n39681 ;
  assign n39683 = \pi1157  & ~n39581 ;
  assign n39684 = ~n39579 & n39683 ;
  assign n39685 = ~\pi1157  & ~n39586 ;
  assign n39686 = ~n39584 & n39685 ;
  assign n39687 = ~n39684 & ~n39686 ;
  assign n39688 = \pi0787  & ~n39687 ;
  assign n39689 = n26333 & ~n39563 ;
  assign n39690 = ~\pi0787  & ~n39689 ;
  assign n39691 = ~\pi1160  & ~n39690 ;
  assign n39692 = n23312 & n39691 ;
  assign n39693 = ~n39688 & n39692 ;
  assign n39694 = ~n39682 & ~n39693 ;
  assign n39695 = ~n23414 & n39532 ;
  assign n39696 = ~n24886 & n39695 ;
  assign n39697 = ~n23313 & ~n39696 ;
  assign n39698 = \pi1160  & ~n39690 ;
  assign n39699 = ~n39688 & n39698 ;
  assign n39700 = n31010 & ~n39593 ;
  assign n39701 = ~n39696 & ~n39700 ;
  assign n39702 = ~n39699 & n39701 ;
  assign n39703 = ~n39697 & ~n39702 ;
  assign n39704 = n39694 & ~n39703 ;
  assign n39705 = \pi0790  & ~n39704 ;
  assign n39706 = \pi0832  & ~n39705 ;
  assign n39707 = n39680 & n39706 ;
  assign n39708 = \pi0190  & ~n6861 ;
  assign n39709 = ~\pi0190  & ~\pi0699  ;
  assign n39710 = ~\pi0038  & n39709 ;
  assign n39711 = n21743 & n39710 ;
  assign n39712 = ~n21734 & n39711 ;
  assign n39713 = \pi0038  & n39709 ;
  assign n39714 = ~n22123 & n39713 ;
  assign n39715 = n6861 & ~n39714 ;
  assign n39716 = ~n39712 & n39715 ;
  assign n39717 = ~n39708 & ~n39716 ;
  assign n39718 = ~\pi0190  & ~n22017 ;
  assign n39719 = ~n21994 & n39718 ;
  assign n39720 = ~\pi0038  & ~\pi0190  ;
  assign n39721 = ~n22109 & ~n39720 ;
  assign n39722 = ~n39719 & ~n39721 ;
  assign n39723 = ~\pi0190  & ~n21757 ;
  assign n39724 = n22117 & ~n39723 ;
  assign n39725 = \pi0699  & ~n39708 ;
  assign n39726 = ~n39724 & n39725 ;
  assign n39727 = ~n39722 & n39726 ;
  assign n39728 = ~n39717 & ~n39727 ;
  assign n39729 = ~\pi0778  & n39728 ;
  assign n39730 = ~\pi0190  & \pi0763  ;
  assign n39731 = ~n21467 & n39730 ;
  assign n39732 = ~\pi0039  & n39730 ;
  assign n39733 = n21272 & n39732 ;
  assign n39734 = ~n39731 & ~n39733 ;
  assign n39735 = \pi0763  & n21484 ;
  assign n39736 = ~\pi0190  & n21743 ;
  assign n39737 = ~n39730 & ~n39736 ;
  assign n39738 = ~n39735 & n39737 ;
  assign n39739 = n39734 & ~n39738 ;
  assign n39740 = ~\pi0038  & ~n39739 ;
  assign n39741 = ~\pi0763  & ~n21731 ;
  assign n39742 = n21714 & n39741 ;
  assign n39743 = ~n21693 & n39742 ;
  assign n39744 = \pi0190  & ~n21543 ;
  assign n39745 = \pi0190  & n21562 ;
  assign n39746 = ~n21552 & n39745 ;
  assign n39747 = ~n39744 & ~n39746 ;
  assign n39748 = ~n21536 & ~n39747 ;
  assign n39749 = ~n39743 & ~n39748 ;
  assign n39750 = n9627 & ~n39749 ;
  assign n39751 = n8413 & n39530 ;
  assign n39752 = n1354 & n39751 ;
  assign n39753 = n1358 & n39752 ;
  assign n39754 = \pi0038  & ~n39753 ;
  assign n39755 = ~n39723 & n39754 ;
  assign n39756 = ~n39708 & ~n39755 ;
  assign n39757 = ~n39750 & n39756 ;
  assign n39758 = ~n39740 & n39757 ;
  assign n39759 = ~\pi0190  & ~n6861 ;
  assign n39760 = ~\pi1155  & ~n39759 ;
  assign n39761 = n22767 & n39760 ;
  assign n39762 = ~n39758 & n39761 ;
  assign n39763 = ~\pi0190  & n21768 ;
  assign n39764 = ~\pi0190  & n21770 ;
  assign n39765 = ~n21734 & n39764 ;
  assign n39766 = ~n39763 & ~n39765 ;
  assign n39767 = ~n32768 & n39766 ;
  assign n39768 = ~n22787 & ~n39767 ;
  assign n39769 = ~n39762 & n39768 ;
  assign n39770 = n39729 & ~n39769 ;
  assign n39771 = \pi0625  & ~n39728 ;
  assign n39772 = ~\pi0190  & ~\pi0625  ;
  assign n39773 = n21768 & n39772 ;
  assign n39774 = n21770 & n39772 ;
  assign n39775 = ~n21734 & n39774 ;
  assign n39776 = ~n39773 & ~n39775 ;
  assign n39777 = \pi1153  & n39776 ;
  assign n39778 = ~n39771 & n39777 ;
  assign n39779 = ~\pi0625  & ~n39728 ;
  assign n39780 = ~\pi0190  & \pi0625  ;
  assign n39781 = n21768 & n39780 ;
  assign n39782 = n21770 & n39780 ;
  assign n39783 = ~n21734 & n39782 ;
  assign n39784 = ~n39781 & ~n39783 ;
  assign n39785 = ~\pi1153  & n39784 ;
  assign n39786 = ~n39779 & n39785 ;
  assign n39787 = ~n39778 & ~n39786 ;
  assign n39788 = \pi0778  & ~n39769 ;
  assign n39789 = ~n39787 & n39788 ;
  assign n39790 = ~n39770 & ~n39789 ;
  assign n39791 = \pi0609  & \pi0785  ;
  assign n39792 = ~n39790 & n39791 ;
  assign n39793 = n31109 & ~n39787 ;
  assign n39794 = n22767 & ~n39759 ;
  assign n39795 = ~n39758 & n39794 ;
  assign n39796 = ~n22767 & n39766 ;
  assign n39797 = \pi0660  & ~n39796 ;
  assign n39798 = ~n39795 & n39797 ;
  assign n39799 = ~n22766 & ~n39798 ;
  assign n39800 = n39367 & n39728 ;
  assign n39801 = ~n39799 & ~n39800 ;
  assign n39802 = ~n39793 & n39801 ;
  assign n39803 = n22788 & ~n39759 ;
  assign n39804 = ~n39758 & n39803 ;
  assign n39805 = ~n22788 & n39766 ;
  assign n39806 = ~\pi0660  & ~n39805 ;
  assign n39807 = ~n39804 & n39806 ;
  assign n39808 = n31121 & ~n39807 ;
  assign n39809 = ~n39802 & n39808 ;
  assign n39810 = ~n39792 & ~n39809 ;
  assign n39811 = n26700 & ~n39810 ;
  assign n39812 = \pi0778  & ~n39787 ;
  assign n39813 = \pi0609  & ~n39729 ;
  assign n39814 = ~n39812 & n39813 ;
  assign n39815 = ~n39769 & ~n39814 ;
  assign n39816 = n21774 & ~n22787 ;
  assign n39817 = ~n39807 & n39816 ;
  assign n39818 = \pi0785  & ~n39817 ;
  assign n39819 = ~n39815 & n39818 ;
  assign n39820 = ~\pi0699  & ~n39755 ;
  assign n39821 = ~n39750 & n39820 ;
  assign n39822 = ~n39740 & n39821 ;
  assign n39823 = n6861 & ~n39822 ;
  assign n39824 = ~n22734 & ~n39772 ;
  assign n39825 = ~n39823 & ~n39824 ;
  assign n39826 = ~\pi0190  & ~n23568 ;
  assign n39827 = \pi0190  & n23575 ;
  assign n39828 = n23572 & n39827 ;
  assign n39829 = ~\pi0038  & ~\pi0763  ;
  assign n39830 = ~n39828 & n39829 ;
  assign n39831 = ~n39826 & n39830 ;
  assign n39832 = \pi0190  & \pi0603  ;
  assign n39833 = ~n20783 & n39832 ;
  assign n39834 = n39529 & n39833 ;
  assign n39835 = \pi0190  & \pi0680  ;
  assign n39836 = ~n20854 & n39835 ;
  assign n39837 = ~n20784 & n39836 ;
  assign n39838 = n1689 & n39837 ;
  assign n39839 = ~n39834 & ~n39838 ;
  assign n39840 = n26554 & ~n39839 ;
  assign n39841 = n1358 & n39840 ;
  assign n39842 = \pi0038  & ~n39841 ;
  assign n39843 = \pi0699  & ~n39842 ;
  assign n39844 = ~\pi0190  & \pi0699  ;
  assign n39845 = \pi0763  & ~n22317 ;
  assign n39846 = ~n31169 & ~n39845 ;
  assign n39847 = ~\pi0039  & n39846 ;
  assign n39848 = n21289 & n39847 ;
  assign n39849 = n39844 & ~n39848 ;
  assign n39850 = ~n39843 & ~n39849 ;
  assign n39851 = ~n39831 & ~n39850 ;
  assign n39852 = ~\pi0039  & ~\pi0190  ;
  assign n39853 = ~n22683 & n39852 ;
  assign n39854 = ~\pi0190  & ~n23548 ;
  assign n39855 = \pi0763  & ~n39854 ;
  assign n39856 = ~n39853 & n39855 ;
  assign n39857 = \pi0190  & ~n23558 ;
  assign n39858 = n23557 & n39857 ;
  assign n39859 = ~\pi0038  & ~n39858 ;
  assign n39860 = n39856 & n39859 ;
  assign n39861 = ~n39824 & ~n39860 ;
  assign n39862 = n39851 & n39861 ;
  assign n39863 = ~n39825 & ~n39862 ;
  assign n39864 = ~\pi1153  & ~n39759 ;
  assign n39865 = ~n39758 & n39864 ;
  assign n39866 = ~n24561 & ~n39865 ;
  assign n39867 = n39863 & ~n39866 ;
  assign n39868 = ~\pi0608  & ~n39777 ;
  assign n39869 = n22755 & ~n39728 ;
  assign n39870 = ~n39868 & ~n39869 ;
  assign n39871 = ~n39867 & ~n39870 ;
  assign n39872 = ~n22727 & ~n39780 ;
  assign n39873 = ~n39823 & ~n39872 ;
  assign n39874 = ~n39860 & ~n39872 ;
  assign n39875 = n39851 & n39874 ;
  assign n39876 = ~n39873 & ~n39875 ;
  assign n39877 = \pi1153  & ~n39759 ;
  assign n39878 = ~n39758 & n39877 ;
  assign n39879 = ~n24550 & ~n39878 ;
  assign n39880 = n39876 & ~n39879 ;
  assign n39881 = \pi0608  & ~n39785 ;
  assign n39882 = n22740 & ~n39728 ;
  assign n39883 = ~n39881 & ~n39882 ;
  assign n39884 = ~n39880 & ~n39883 ;
  assign n39885 = ~n39871 & ~n39884 ;
  assign n39886 = \pi0778  & ~n39885 ;
  assign n39887 = ~n39819 & ~n39886 ;
  assign n39888 = ~\pi0190  & ~\pi0778  ;
  assign n39889 = ~n23622 & ~n39888 ;
  assign n39890 = ~n39823 & ~n39889 ;
  assign n39891 = ~n39860 & ~n39889 ;
  assign n39892 = n39851 & n39891 ;
  assign n39893 = ~n39890 & ~n39892 ;
  assign n39894 = n26700 & n39893 ;
  assign n39895 = n39887 & n39894 ;
  assign n39896 = ~n39811 & ~n39895 ;
  assign n39897 = ~\pi0190  & ~n20811 ;
  assign n39898 = n21768 & n39897 ;
  assign n39899 = n21770 & n39897 ;
  assign n39900 = ~n21734 & n39899 ;
  assign n39901 = ~n39898 & ~n39900 ;
  assign n39902 = n23424 & ~n39901 ;
  assign n39903 = n21777 & ~n39759 ;
  assign n39904 = ~n39758 & n39903 ;
  assign n39905 = ~n21777 & n39766 ;
  assign n39906 = n20811 & ~n39905 ;
  assign n39907 = n23424 & n39906 ;
  assign n39908 = ~n39904 & n39907 ;
  assign n39909 = ~n39902 & ~n39908 ;
  assign n39910 = ~\pi0781  & ~n39905 ;
  assign n39911 = ~n23423 & n39910 ;
  assign n39912 = ~n39904 & n39911 ;
  assign n39913 = n23423 & ~n39766 ;
  assign n39914 = ~n39912 & ~n39913 ;
  assign n39915 = n39909 & n39914 ;
  assign n39916 = ~n23880 & ~n39915 ;
  assign n39917 = n23880 & ~n39766 ;
  assign n39918 = n24691 & ~n39917 ;
  assign n39919 = ~n39916 & n39918 ;
  assign n39920 = n26065 & ~n39787 ;
  assign n39921 = n26739 & n39728 ;
  assign n39922 = ~n23885 & n39766 ;
  assign n39923 = \pi0628  & ~n39922 ;
  assign n39924 = ~n39921 & n39923 ;
  assign n39925 = ~n39920 & n39924 ;
  assign n39926 = ~\pi0190  & ~\pi0628  ;
  assign n39927 = n21768 & n39926 ;
  assign n39928 = n21770 & n39926 ;
  assign n39929 = ~n21734 & n39928 ;
  assign n39930 = ~n39927 & ~n39929 ;
  assign n39931 = n20843 & n39930 ;
  assign n39932 = ~n39925 & n39931 ;
  assign n39933 = ~\pi0628  & ~n39922 ;
  assign n39934 = ~n39921 & n39933 ;
  assign n39935 = ~n39920 & n39934 ;
  assign n39936 = ~\pi0190  & \pi0628  ;
  assign n39937 = n21768 & n39936 ;
  assign n39938 = n21770 & n39936 ;
  assign n39939 = ~n21734 & n39938 ;
  assign n39940 = ~n39937 & ~n39939 ;
  assign n39941 = n20844 & n39940 ;
  assign n39942 = ~n39935 & n39941 ;
  assign n39943 = ~n39932 & ~n39942 ;
  assign n39944 = ~n39919 & n39943 ;
  assign n39945 = \pi0792  & ~n39944 ;
  assign n39946 = ~n39904 & n39906 ;
  assign n39947 = n22155 & n39901 ;
  assign n39948 = ~n39946 & n39947 ;
  assign n39949 = ~n22147 & ~n39729 ;
  assign n39950 = n22147 & ~n39766 ;
  assign n39951 = \pi0781  & n23666 ;
  assign n39952 = ~n20811 & n39951 ;
  assign n39953 = ~n39950 & n39952 ;
  assign n39954 = ~n39949 & n39953 ;
  assign n39955 = \pi0778  & n39953 ;
  assign n39956 = ~n39787 & n39955 ;
  assign n39957 = ~n39954 & ~n39956 ;
  assign n39958 = ~n39948 & n39957 ;
  assign n39959 = ~n21034 & ~n39958 ;
  assign n39960 = n30780 & ~n39787 ;
  assign n39961 = n31274 & n39728 ;
  assign n39962 = ~n23380 & n39766 ;
  assign n39963 = ~n39961 & ~n39962 ;
  assign n39964 = ~n39960 & n39963 ;
  assign n39965 = ~n31283 & ~n39964 ;
  assign n39966 = n23683 & ~n39901 ;
  assign n39967 = n23683 & n39906 ;
  assign n39968 = ~n39904 & n39967 ;
  assign n39969 = ~n39966 & ~n39968 ;
  assign n39970 = n21032 & n39910 ;
  assign n39971 = ~n39904 & n39970 ;
  assign n39972 = ~n21032 & ~n39766 ;
  assign n39973 = ~n20876 & ~n39972 ;
  assign n39974 = \pi0789  & n39973 ;
  assign n39975 = ~n39971 & n39974 ;
  assign n39976 = n39969 & n39975 ;
  assign n39977 = ~n21038 & ~n39976 ;
  assign n39978 = ~n39965 & n39977 ;
  assign n39979 = ~n39959 & n39978 ;
  assign n39980 = ~n39945 & n39979 ;
  assign n39981 = n39896 & n39980 ;
  assign n39982 = n20951 & ~n39766 ;
  assign n39983 = ~n31301 & ~n39982 ;
  assign n39984 = ~n39961 & ~n39983 ;
  assign n39985 = ~n39960 & n39984 ;
  assign n39986 = n31306 & ~n39766 ;
  assign n39987 = ~n23856 & ~n39986 ;
  assign n39988 = ~n39985 & n39987 ;
  assign n39989 = ~\pi0626  & ~n39913 ;
  assign n39990 = ~n39912 & n39989 ;
  assign n39991 = n39909 & n39990 ;
  assign n39992 = \pi0626  & n39766 ;
  assign n39993 = n20882 & ~n39992 ;
  assign n39994 = ~n39991 & n39993 ;
  assign n39995 = \pi0626  & ~n39913 ;
  assign n39996 = ~n39912 & n39995 ;
  assign n39997 = n39909 & n39996 ;
  assign n39998 = ~\pi0626  & n39766 ;
  assign n39999 = n20881 & ~n39998 ;
  assign n40000 = ~n39997 & n39999 ;
  assign n40001 = ~n39994 & ~n40000 ;
  assign n40002 = n39988 & n40001 ;
  assign n40003 = ~n26803 & ~n40002 ;
  assign n40004 = ~n21067 & ~n40003 ;
  assign n40005 = n24724 & ~n39944 ;
  assign n40006 = ~n40004 & ~n40005 ;
  assign n40007 = ~n39981 & ~n40006 ;
  assign n40008 = ~n20846 & n39917 ;
  assign n40009 = n30376 & ~n39915 ;
  assign n40010 = ~n40008 & ~n40009 ;
  assign n40011 = n20846 & ~n39766 ;
  assign n40012 = ~n20910 & ~n40011 ;
  assign n40013 = n40010 & n40012 ;
  assign n40014 = n21768 & n39585 ;
  assign n40015 = n21770 & n39585 ;
  assign n40016 = ~n21734 & n40015 ;
  assign n40017 = ~n40014 & ~n40016 ;
  assign n40018 = n31338 & n40017 ;
  assign n40019 = ~n23907 & ~n39922 ;
  assign n40020 = ~n39921 & n40019 ;
  assign n40021 = ~n39920 & n40020 ;
  assign n40022 = \pi0792  & ~n20888 ;
  assign n40023 = ~n39766 & n40022 ;
  assign n40024 = n20897 & n40017 ;
  assign n40025 = ~n40023 & n40024 ;
  assign n40026 = ~n40021 & n40025 ;
  assign n40027 = ~n40018 & ~n40026 ;
  assign n40028 = n21768 & n39580 ;
  assign n40029 = n21770 & n39580 ;
  assign n40030 = ~n21734 & n40029 ;
  assign n40031 = ~n40028 & ~n40030 ;
  assign n40032 = ~\pi0647  & n20849 ;
  assign n40033 = n40031 & n40032 ;
  assign n40034 = n20849 & n40031 ;
  assign n40035 = ~n40023 & n40034 ;
  assign n40036 = ~n40021 & n40035 ;
  assign n40037 = ~n40033 & ~n40036 ;
  assign n40038 = n40027 & n40037 ;
  assign n40039 = ~n40013 & n40038 ;
  assign n40040 = \pi0787  & ~n40039 ;
  assign n40041 = ~\pi0190  & \pi0644  ;
  assign n40042 = n21768 & n40041 ;
  assign n40043 = n21770 & n40041 ;
  assign n40044 = ~n21734 & n40043 ;
  assign n40045 = ~n40042 & ~n40044 ;
  assign n40046 = n23939 & n40045 ;
  assign n40047 = \pi0715  & n40045 ;
  assign n40048 = ~\pi0190  & ~n31367 ;
  assign n40049 = n21768 & n40048 ;
  assign n40050 = n21770 & n40048 ;
  assign n40051 = ~n21734 & n40050 ;
  assign n40052 = ~n40049 & ~n40051 ;
  assign n40053 = n40047 & n40052 ;
  assign n40054 = ~n40046 & ~n40053 ;
  assign n40055 = n31367 & ~n40046 ;
  assign n40056 = ~n39915 & n40055 ;
  assign n40057 = ~n40054 & ~n40056 ;
  assign n40058 = n31378 & ~n40057 ;
  assign n40059 = ~\pi0715  & n40052 ;
  assign n40060 = ~n23958 & ~n40059 ;
  assign n40061 = n31382 & ~n39915 ;
  assign n40062 = ~n40060 & ~n40061 ;
  assign n40063 = n26824 & ~n40062 ;
  assign n40064 = \pi0790  & ~n40063 ;
  assign n40065 = ~n40058 & n40064 ;
  assign n40066 = n9948 & ~n40065 ;
  assign n40067 = ~n40040 & n40066 ;
  assign n40068 = ~n40007 & n40067 ;
  assign n40069 = n23942 & n39766 ;
  assign n40070 = \pi0644  & ~n40069 ;
  assign n40071 = ~\pi0715  & ~n40070 ;
  assign n40072 = ~n23942 & ~n40023 ;
  assign n40073 = ~\pi0715  & n40072 ;
  assign n40074 = ~n40021 & n40073 ;
  assign n40075 = ~n40071 & ~n40074 ;
  assign n40076 = ~\pi1160  & ~n40057 ;
  assign n40077 = n40075 & n40076 ;
  assign n40078 = n9948 & n40077 ;
  assign n40079 = ~\pi0190  & ~\pi0644  ;
  assign n40080 = n21768 & n40079 ;
  assign n40081 = n21770 & n40079 ;
  assign n40082 = ~n21734 & n40081 ;
  assign n40083 = ~n40080 & ~n40082 ;
  assign n40084 = n40062 & n40083 ;
  assign n40085 = ~\pi0644  & ~n40069 ;
  assign n40086 = \pi0715  & ~n40085 ;
  assign n40087 = \pi0715  & n40072 ;
  assign n40088 = ~n40021 & n40087 ;
  assign n40089 = ~n40086 & ~n40088 ;
  assign n40090 = ~n40084 & n40089 ;
  assign n40091 = n31413 & n40090 ;
  assign n40092 = ~n40078 & ~n40091 ;
  assign n40093 = \pi0790  & ~n40092 ;
  assign n40094 = \pi0190  & ~\pi0832  ;
  assign n40095 = ~n21132 & ~n40094 ;
  assign n40096 = ~n40093 & ~n40095 ;
  assign n40097 = ~n40068 & n40096 ;
  assign n40098 = ~n39707 & ~n40097 ;
  assign n40099 = ~\pi0191  & \pi0788  ;
  assign n40100 = ~n1689 & n40099 ;
  assign n40101 = ~n20778 & n40100 ;
  assign n40102 = n20886 & n40101 ;
  assign n40103 = \pi0746  & n1689 ;
  assign n40104 = n20784 & n40103 ;
  assign n40105 = n22767 & n40104 ;
  assign n40106 = ~\pi0191  & ~n1689 ;
  assign n40107 = ~n40104 & ~n40106 ;
  assign n40108 = ~n20792 & ~n40107 ;
  assign n40109 = ~n40105 & n40108 ;
  assign n40110 = n20801 & ~n40109 ;
  assign n40111 = ~\pi1155  & ~n40106 ;
  assign n40112 = \pi0785  & n40111 ;
  assign n40113 = ~n40105 & n40112 ;
  assign n40114 = ~\pi0785  & ~n40106 ;
  assign n40115 = ~n40104 & n40114 ;
  assign n40116 = ~n20804 & ~n40115 ;
  assign n40117 = n29682 & n40116 ;
  assign n40118 = ~n40113 & n40117 ;
  assign n40119 = ~n40110 & n40118 ;
  assign n40120 = n30847 & n40119 ;
  assign n40121 = ~n40102 & ~n40120 ;
  assign n40122 = \pi0729  & n1689 ;
  assign n40123 = n20855 & n40122 ;
  assign n40124 = ~n40106 & ~n40123 ;
  assign n40125 = ~\pi0778  & ~n40124 ;
  assign n40126 = ~\pi0625  & \pi0729  ;
  assign n40127 = n1689 & n40126 ;
  assign n40128 = n20855 & n40127 ;
  assign n40129 = \pi1153  & n40128 ;
  assign n40130 = \pi1153  & ~n40106 ;
  assign n40131 = ~n40123 & n40130 ;
  assign n40132 = ~n40129 & ~n40131 ;
  assign n40133 = ~\pi1153  & ~n40106 ;
  assign n40134 = ~n40128 & n40133 ;
  assign n40135 = \pi0778  & ~n40134 ;
  assign n40136 = n40132 & n40135 ;
  assign n40137 = ~n40125 & ~n40136 ;
  assign n40138 = n26474 & ~n40137 ;
  assign n40139 = \pi0629  & ~n40138 ;
  assign n40140 = n40121 & n40139 ;
  assign n40141 = n20887 & n40101 ;
  assign n40142 = n32579 & n40119 ;
  assign n40143 = ~n40141 & ~n40142 ;
  assign n40144 = n26485 & ~n40137 ;
  assign n40145 = ~\pi0629  & ~n40144 ;
  assign n40146 = n40143 & n40145 ;
  assign n40147 = ~n40140 & ~n40146 ;
  assign n40148 = \pi0792  & n40147 ;
  assign n40149 = ~n21067 & ~n40148 ;
  assign n40150 = n39578 & ~n40137 ;
  assign n40151 = ~\pi0191  & ~\pi0647  ;
  assign n40152 = ~n1689 & n40151 ;
  assign n40153 = n20849 & ~n40152 ;
  assign n40154 = ~n40150 & n40153 ;
  assign n40155 = n26319 & ~n40137 ;
  assign n40156 = ~\pi0191  & \pi0647  ;
  assign n40157 = ~n1689 & n40156 ;
  assign n40158 = n20897 & ~n40157 ;
  assign n40159 = ~n40155 & n40158 ;
  assign n40160 = ~n40154 & ~n40159 ;
  assign n40161 = \pi0787  & ~n40160 ;
  assign n40162 = ~n20846 & n40101 ;
  assign n40163 = n30376 & n40119 ;
  assign n40164 = ~n40162 & ~n40163 ;
  assign n40165 = ~\pi0191  & \pi0792  ;
  assign n40166 = ~n1689 & n40165 ;
  assign n40167 = ~n20845 & n40166 ;
  assign n40168 = n32606 & ~n40167 ;
  assign n40169 = n40164 & n40168 ;
  assign n40170 = ~n40161 & ~n40169 ;
  assign n40171 = ~n24761 & n40170 ;
  assign n40172 = ~n40149 & n40171 ;
  assign n40173 = \pi0608  & ~n40134 ;
  assign n40174 = ~n40104 & n40130 ;
  assign n40175 = \pi0778  & ~n40174 ;
  assign n40176 = n26421 & ~n40124 ;
  assign n40177 = ~n40175 & ~n40176 ;
  assign n40178 = n40173 & ~n40177 ;
  assign n40179 = n26147 & ~n40124 ;
  assign n40180 = \pi0729  & ~n20784 ;
  assign n40181 = n22113 & n40180 ;
  assign n40182 = n40107 & ~n40181 ;
  assign n40183 = ~n40179 & ~n40182 ;
  assign n40184 = n40133 & ~n40183 ;
  assign n40185 = n26415 & n40132 ;
  assign n40186 = ~n40184 & n40185 ;
  assign n40187 = ~n40178 & ~n40186 ;
  assign n40188 = ~\pi1155  & ~n40125 ;
  assign n40189 = ~n40136 & n40188 ;
  assign n40190 = ~n20999 & ~n40189 ;
  assign n40191 = ~\pi0778  & ~n40182 ;
  assign n40192 = ~n40190 & ~n40191 ;
  assign n40193 = n40187 & n40192 ;
  assign n40194 = n29766 & ~n40125 ;
  assign n40195 = ~n40136 & n40194 ;
  assign n40196 = \pi1155  & ~n40109 ;
  assign n40197 = ~\pi0660  & ~n40196 ;
  assign n40198 = ~n40195 & n40197 ;
  assign n40199 = ~n40193 & n40198 ;
  assign n40200 = \pi0785  & ~n40199 ;
  assign n40201 = n29775 & n40116 ;
  assign n40202 = ~n40113 & n40201 ;
  assign n40203 = ~n40110 & n40202 ;
  assign n40204 = n29779 & ~n40137 ;
  assign n40205 = ~n40203 & ~n40204 ;
  assign n40206 = \pi0781  & ~n40205 ;
  assign n40207 = \pi1155  & ~n40125 ;
  assign n40208 = ~n40136 & n40207 ;
  assign n40209 = ~n21774 & ~n40208 ;
  assign n40210 = ~n40191 & ~n40209 ;
  assign n40211 = n40187 & n40210 ;
  assign n40212 = n26121 & ~n40125 ;
  assign n40213 = ~n40136 & n40212 ;
  assign n40214 = \pi0660  & ~n40111 ;
  assign n40215 = \pi0660  & n40104 ;
  assign n40216 = n22767 & n40215 ;
  assign n40217 = ~n40214 & ~n40216 ;
  assign n40218 = ~n40213 & ~n40217 ;
  assign n40219 = ~n40211 & n40218 ;
  assign n40220 = ~n40206 & ~n40219 ;
  assign n40221 = n40200 & n40220 ;
  assign n40222 = ~\pi0785  & ~n40191 ;
  assign n40223 = ~n40178 & n40222 ;
  assign n40224 = ~n40186 & n40223 ;
  assign n40225 = n21022 & ~n40224 ;
  assign n40226 = ~n40206 & ~n40225 ;
  assign n40227 = n29803 & ~n40226 ;
  assign n40228 = ~n40221 & n40227 ;
  assign n40229 = n29808 & n40116 ;
  assign n40230 = ~n40113 & n40229 ;
  assign n40231 = ~n40110 & n40230 ;
  assign n40232 = n30966 & ~n40137 ;
  assign n40233 = ~n40231 & ~n40232 ;
  assign n40234 = n36155 & ~n40233 ;
  assign n40235 = \pi0626  & ~n40119 ;
  assign n40236 = ~\pi0626  & ~n40106 ;
  assign n40237 = n20881 & ~n40236 ;
  assign n40238 = ~n40235 & n40237 ;
  assign n40239 = n26458 & ~n40137 ;
  assign n40240 = ~\pi0626  & ~n40119 ;
  assign n40241 = \pi0626  & ~n40106 ;
  assign n40242 = n20882 & ~n40241 ;
  assign n40243 = ~n40240 & n40242 ;
  assign n40244 = ~n40239 & ~n40243 ;
  assign n40245 = ~n40238 & n40244 ;
  assign n40246 = \pi0788  & ~n40245 ;
  assign n40247 = ~n40234 & ~n40246 ;
  assign n40248 = ~n40228 & n40247 ;
  assign n40249 = ~n23856 & n40171 ;
  assign n40250 = ~n40248 & n40249 ;
  assign n40251 = ~n40172 & ~n40250 ;
  assign n40252 = n30987 & ~n40164 ;
  assign n40253 = n23312 & n40252 ;
  assign n40254 = \pi1157  & ~n40152 ;
  assign n40255 = ~n40150 & n40254 ;
  assign n40256 = ~\pi1157  & ~n40157 ;
  assign n40257 = ~n40155 & n40256 ;
  assign n40258 = ~n40255 & ~n40257 ;
  assign n40259 = \pi0787  & ~n40258 ;
  assign n40260 = n26333 & ~n40137 ;
  assign n40261 = ~\pi0787  & ~n40260 ;
  assign n40262 = ~\pi1160  & ~n40261 ;
  assign n40263 = n23312 & n40262 ;
  assign n40264 = ~n40259 & n40263 ;
  assign n40265 = ~n40253 & ~n40264 ;
  assign n40266 = ~n23414 & n40106 ;
  assign n40267 = ~n24886 & n40266 ;
  assign n40268 = ~n23313 & ~n40267 ;
  assign n40269 = \pi1160  & ~n40261 ;
  assign n40270 = ~n40259 & n40269 ;
  assign n40271 = n31010 & ~n40164 ;
  assign n40272 = ~n40267 & ~n40271 ;
  assign n40273 = ~n40270 & n40272 ;
  assign n40274 = ~n40268 & ~n40273 ;
  assign n40275 = n40265 & ~n40274 ;
  assign n40276 = \pi0790  & ~n40275 ;
  assign n40277 = \pi0832  & ~n40276 ;
  assign n40278 = n40251 & n40277 ;
  assign n40279 = \pi0191  & ~n6861 ;
  assign n40280 = ~\pi0191  & ~\pi0729  ;
  assign n40281 = ~\pi0038  & n40280 ;
  assign n40282 = n21743 & n40281 ;
  assign n40283 = ~n21734 & n40282 ;
  assign n40284 = \pi0038  & n40280 ;
  assign n40285 = ~n22123 & n40284 ;
  assign n40286 = n6861 & ~n40285 ;
  assign n40287 = ~n40283 & n40286 ;
  assign n40288 = ~n40279 & ~n40287 ;
  assign n40289 = ~\pi0191  & ~n22017 ;
  assign n40290 = ~n21994 & n40289 ;
  assign n40291 = ~\pi0038  & ~\pi0191  ;
  assign n40292 = ~n22109 & ~n40291 ;
  assign n40293 = ~n40290 & ~n40292 ;
  assign n40294 = ~\pi0191  & ~n21757 ;
  assign n40295 = n22117 & ~n40294 ;
  assign n40296 = \pi0729  & ~n40279 ;
  assign n40297 = ~n40295 & n40296 ;
  assign n40298 = ~n40293 & n40297 ;
  assign n40299 = ~n40288 & ~n40298 ;
  assign n40300 = ~\pi0778  & n40299 ;
  assign n40301 = ~\pi0191  & \pi0746  ;
  assign n40302 = ~n21467 & n40301 ;
  assign n40303 = ~\pi0039  & n40301 ;
  assign n40304 = n21272 & n40303 ;
  assign n40305 = ~n40302 & ~n40304 ;
  assign n40306 = \pi0746  & n21484 ;
  assign n40307 = ~\pi0191  & n21743 ;
  assign n40308 = ~n40301 & ~n40307 ;
  assign n40309 = ~n40306 & n40308 ;
  assign n40310 = n40305 & ~n40309 ;
  assign n40311 = ~\pi0038  & ~n40310 ;
  assign n40312 = ~\pi0746  & ~n21731 ;
  assign n40313 = n21714 & n40312 ;
  assign n40314 = ~n21693 & n40313 ;
  assign n40315 = \pi0191  & ~n21543 ;
  assign n40316 = \pi0191  & n21562 ;
  assign n40317 = ~n21552 & n40316 ;
  assign n40318 = ~n40315 & ~n40317 ;
  assign n40319 = ~n21536 & ~n40318 ;
  assign n40320 = ~n40314 & ~n40319 ;
  assign n40321 = n9627 & ~n40320 ;
  assign n40322 = n8413 & n40104 ;
  assign n40323 = n1354 & n40322 ;
  assign n40324 = n1358 & n40323 ;
  assign n40325 = \pi0038  & ~n40324 ;
  assign n40326 = ~n40294 & n40325 ;
  assign n40327 = ~n40279 & ~n40326 ;
  assign n40328 = ~n40321 & n40327 ;
  assign n40329 = ~n40311 & n40328 ;
  assign n40330 = ~\pi0191  & ~n6861 ;
  assign n40331 = ~\pi1155  & ~n40330 ;
  assign n40332 = n22767 & n40331 ;
  assign n40333 = ~n40329 & n40332 ;
  assign n40334 = ~\pi0191  & n21768 ;
  assign n40335 = ~\pi0191  & n21770 ;
  assign n40336 = ~n21734 & n40335 ;
  assign n40337 = ~n40334 & ~n40336 ;
  assign n40338 = ~n32768 & n40337 ;
  assign n40339 = ~n22787 & ~n40338 ;
  assign n40340 = ~n40333 & n40339 ;
  assign n40341 = n40300 & ~n40340 ;
  assign n40342 = \pi0625  & ~n40299 ;
  assign n40343 = ~\pi0191  & ~\pi0625  ;
  assign n40344 = n21768 & n40343 ;
  assign n40345 = n21770 & n40343 ;
  assign n40346 = ~n21734 & n40345 ;
  assign n40347 = ~n40344 & ~n40346 ;
  assign n40348 = \pi1153  & n40347 ;
  assign n40349 = ~n40342 & n40348 ;
  assign n40350 = ~\pi0625  & ~n40299 ;
  assign n40351 = ~\pi0191  & \pi0625  ;
  assign n40352 = n21768 & n40351 ;
  assign n40353 = n21770 & n40351 ;
  assign n40354 = ~n21734 & n40353 ;
  assign n40355 = ~n40352 & ~n40354 ;
  assign n40356 = ~\pi1153  & n40355 ;
  assign n40357 = ~n40350 & n40356 ;
  assign n40358 = ~n40349 & ~n40357 ;
  assign n40359 = \pi0778  & ~n40340 ;
  assign n40360 = ~n40358 & n40359 ;
  assign n40361 = ~n40341 & ~n40360 ;
  assign n40362 = n39791 & ~n40361 ;
  assign n40363 = n31109 & ~n40358 ;
  assign n40364 = n22767 & ~n40330 ;
  assign n40365 = ~n40329 & n40364 ;
  assign n40366 = ~n22767 & n40337 ;
  assign n40367 = \pi0660  & ~n40366 ;
  assign n40368 = ~n40365 & n40367 ;
  assign n40369 = ~n22766 & ~n40368 ;
  assign n40370 = n39367 & n40299 ;
  assign n40371 = ~n40369 & ~n40370 ;
  assign n40372 = ~n40363 & n40371 ;
  assign n40373 = n22788 & ~n40330 ;
  assign n40374 = ~n40329 & n40373 ;
  assign n40375 = ~n22788 & n40337 ;
  assign n40376 = ~\pi0660  & ~n40375 ;
  assign n40377 = ~n40374 & n40376 ;
  assign n40378 = n31121 & ~n40377 ;
  assign n40379 = ~n40372 & n40378 ;
  assign n40380 = ~n40362 & ~n40379 ;
  assign n40381 = n26700 & ~n40380 ;
  assign n40382 = \pi0778  & ~n40358 ;
  assign n40383 = \pi0609  & ~n40300 ;
  assign n40384 = ~n40382 & n40383 ;
  assign n40385 = ~n40340 & ~n40384 ;
  assign n40386 = n39816 & ~n40377 ;
  assign n40387 = \pi0785  & ~n40386 ;
  assign n40388 = ~n40385 & n40387 ;
  assign n40389 = ~\pi0729  & ~n40326 ;
  assign n40390 = ~n40321 & n40389 ;
  assign n40391 = ~n40311 & n40390 ;
  assign n40392 = n6861 & ~n40391 ;
  assign n40393 = ~n22734 & ~n40343 ;
  assign n40394 = ~n40392 & ~n40393 ;
  assign n40395 = ~\pi0039  & ~\pi0191  ;
  assign n40396 = ~n22683 & n40395 ;
  assign n40397 = ~\pi0191  & ~n23548 ;
  assign n40398 = \pi0746  & ~n40397 ;
  assign n40399 = ~n40396 & n40398 ;
  assign n40400 = \pi0191  & ~n23558 ;
  assign n40401 = n23557 & n40400 ;
  assign n40402 = ~\pi0038  & ~n40401 ;
  assign n40403 = n40399 & n40402 ;
  assign n40404 = ~\pi0191  & ~n23568 ;
  assign n40405 = \pi0191  & n23575 ;
  assign n40406 = n23572 & n40405 ;
  assign n40407 = ~\pi0038  & ~\pi0746  ;
  assign n40408 = ~n40406 & n40407 ;
  assign n40409 = ~n40404 & n40408 ;
  assign n40410 = ~n40403 & ~n40409 ;
  assign n40411 = \pi0191  & \pi0603  ;
  assign n40412 = ~n20783 & n40411 ;
  assign n40413 = n40103 & n40412 ;
  assign n40414 = \pi0191  & \pi0680  ;
  assign n40415 = ~n20854 & n40414 ;
  assign n40416 = ~n20784 & n40415 ;
  assign n40417 = n1689 & n40416 ;
  assign n40418 = ~n40413 & ~n40417 ;
  assign n40419 = n26554 & ~n40418 ;
  assign n40420 = n1358 & n40419 ;
  assign n40421 = \pi0038  & ~n40420 ;
  assign n40422 = \pi0729  & ~n40421 ;
  assign n40423 = \pi0746  & ~n22317 ;
  assign n40424 = ~n31169 & ~n40423 ;
  assign n40425 = ~\pi0039  & n40424 ;
  assign n40426 = n21289 & n40425 ;
  assign n40427 = ~\pi0191  & \pi0729  ;
  assign n40428 = ~n40426 & n40427 ;
  assign n40429 = ~n40422 & ~n40428 ;
  assign n40430 = ~n40393 & ~n40429 ;
  assign n40431 = n40410 & n40430 ;
  assign n40432 = ~n40394 & ~n40431 ;
  assign n40433 = ~\pi1153  & ~n40330 ;
  assign n40434 = ~n40329 & n40433 ;
  assign n40435 = ~n24561 & ~n40434 ;
  assign n40436 = n40432 & ~n40435 ;
  assign n40437 = ~\pi0608  & ~n40348 ;
  assign n40438 = n22755 & ~n40299 ;
  assign n40439 = ~n40437 & ~n40438 ;
  assign n40440 = ~n40436 & ~n40439 ;
  assign n40441 = ~n22727 & ~n40351 ;
  assign n40442 = ~n40392 & ~n40441 ;
  assign n40443 = ~n40429 & ~n40441 ;
  assign n40444 = n40410 & n40443 ;
  assign n40445 = ~n40442 & ~n40444 ;
  assign n40446 = \pi1153  & ~n40330 ;
  assign n40447 = ~n40329 & n40446 ;
  assign n40448 = ~n24550 & ~n40447 ;
  assign n40449 = n40445 & ~n40448 ;
  assign n40450 = \pi0608  & ~n40356 ;
  assign n40451 = n22740 & ~n40299 ;
  assign n40452 = ~n40450 & ~n40451 ;
  assign n40453 = ~n40449 & ~n40452 ;
  assign n40454 = ~n40440 & ~n40453 ;
  assign n40455 = \pi0778  & ~n40454 ;
  assign n40456 = ~n40388 & ~n40455 ;
  assign n40457 = ~\pi0191  & ~\pi0778  ;
  assign n40458 = ~n23622 & ~n40457 ;
  assign n40459 = ~n40392 & ~n40458 ;
  assign n40460 = ~n40429 & ~n40458 ;
  assign n40461 = n40410 & n40460 ;
  assign n40462 = ~n40459 & ~n40461 ;
  assign n40463 = n26700 & n40462 ;
  assign n40464 = n40456 & n40463 ;
  assign n40465 = ~n40381 & ~n40464 ;
  assign n40466 = ~\pi0191  & ~n20811 ;
  assign n40467 = n21768 & n40466 ;
  assign n40468 = n21770 & n40466 ;
  assign n40469 = ~n21734 & n40468 ;
  assign n40470 = ~n40467 & ~n40469 ;
  assign n40471 = n23424 & ~n40470 ;
  assign n40472 = n21777 & ~n40330 ;
  assign n40473 = ~n40329 & n40472 ;
  assign n40474 = ~n21777 & n40337 ;
  assign n40475 = n20811 & ~n40474 ;
  assign n40476 = n23424 & n40475 ;
  assign n40477 = ~n40473 & n40476 ;
  assign n40478 = ~n40471 & ~n40477 ;
  assign n40479 = ~\pi0781  & ~n40474 ;
  assign n40480 = ~n23423 & n40479 ;
  assign n40481 = ~n40473 & n40480 ;
  assign n40482 = n23423 & ~n40337 ;
  assign n40483 = ~n40481 & ~n40482 ;
  assign n40484 = n40478 & n40483 ;
  assign n40485 = ~n23880 & ~n40484 ;
  assign n40486 = n23880 & ~n40337 ;
  assign n40487 = n24691 & ~n40486 ;
  assign n40488 = ~n40485 & n40487 ;
  assign n40489 = n26065 & ~n40358 ;
  assign n40490 = n26739 & n40299 ;
  assign n40491 = ~n23885 & n40337 ;
  assign n40492 = \pi0628  & ~n40491 ;
  assign n40493 = ~n40490 & n40492 ;
  assign n40494 = ~n40489 & n40493 ;
  assign n40495 = ~\pi0191  & ~\pi0628  ;
  assign n40496 = n21768 & n40495 ;
  assign n40497 = n21770 & n40495 ;
  assign n40498 = ~n21734 & n40497 ;
  assign n40499 = ~n40496 & ~n40498 ;
  assign n40500 = n20843 & n40499 ;
  assign n40501 = ~n40494 & n40500 ;
  assign n40502 = ~\pi0628  & ~n40491 ;
  assign n40503 = ~n40490 & n40502 ;
  assign n40504 = ~n40489 & n40503 ;
  assign n40505 = ~\pi0191  & \pi0628  ;
  assign n40506 = n21768 & n40505 ;
  assign n40507 = n21770 & n40505 ;
  assign n40508 = ~n21734 & n40507 ;
  assign n40509 = ~n40506 & ~n40508 ;
  assign n40510 = n20844 & n40509 ;
  assign n40511 = ~n40504 & n40510 ;
  assign n40512 = ~n40501 & ~n40511 ;
  assign n40513 = ~n40488 & n40512 ;
  assign n40514 = \pi0792  & ~n40513 ;
  assign n40515 = ~n40473 & n40475 ;
  assign n40516 = n22155 & n40470 ;
  assign n40517 = ~n40515 & n40516 ;
  assign n40518 = ~n22147 & ~n40300 ;
  assign n40519 = n22147 & ~n40337 ;
  assign n40520 = n39952 & ~n40519 ;
  assign n40521 = ~n40518 & n40520 ;
  assign n40522 = \pi0778  & n40520 ;
  assign n40523 = ~n40358 & n40522 ;
  assign n40524 = ~n40521 & ~n40523 ;
  assign n40525 = ~n40517 & n40524 ;
  assign n40526 = ~n21034 & ~n40525 ;
  assign n40527 = n30780 & ~n40358 ;
  assign n40528 = n31274 & n40299 ;
  assign n40529 = ~n23380 & n40337 ;
  assign n40530 = ~n40528 & ~n40529 ;
  assign n40531 = ~n40527 & n40530 ;
  assign n40532 = ~n31283 & ~n40531 ;
  assign n40533 = n23683 & ~n40470 ;
  assign n40534 = n23683 & n40475 ;
  assign n40535 = ~n40473 & n40534 ;
  assign n40536 = ~n40533 & ~n40535 ;
  assign n40537 = n21032 & n40479 ;
  assign n40538 = ~n40473 & n40537 ;
  assign n40539 = ~n21032 & ~n40337 ;
  assign n40540 = ~n20876 & ~n40539 ;
  assign n40541 = \pi0789  & n40540 ;
  assign n40542 = ~n40538 & n40541 ;
  assign n40543 = n40536 & n40542 ;
  assign n40544 = ~n21038 & ~n40543 ;
  assign n40545 = ~n40532 & n40544 ;
  assign n40546 = ~n40526 & n40545 ;
  assign n40547 = ~n40514 & n40546 ;
  assign n40548 = n40465 & n40547 ;
  assign n40549 = n20951 & ~n40337 ;
  assign n40550 = ~n31301 & ~n40549 ;
  assign n40551 = ~n40528 & ~n40550 ;
  assign n40552 = ~n40527 & n40551 ;
  assign n40553 = n31306 & ~n40337 ;
  assign n40554 = ~n23856 & ~n40553 ;
  assign n40555 = ~n40552 & n40554 ;
  assign n40556 = ~\pi0626  & ~n40482 ;
  assign n40557 = ~n40481 & n40556 ;
  assign n40558 = n40478 & n40557 ;
  assign n40559 = \pi0626  & n40337 ;
  assign n40560 = n20882 & ~n40559 ;
  assign n40561 = ~n40558 & n40560 ;
  assign n40562 = \pi0626  & ~n40482 ;
  assign n40563 = ~n40481 & n40562 ;
  assign n40564 = n40478 & n40563 ;
  assign n40565 = ~\pi0626  & n40337 ;
  assign n40566 = n20881 & ~n40565 ;
  assign n40567 = ~n40564 & n40566 ;
  assign n40568 = ~n40561 & ~n40567 ;
  assign n40569 = n40555 & n40568 ;
  assign n40570 = ~n26803 & ~n40569 ;
  assign n40571 = ~n21067 & ~n40570 ;
  assign n40572 = n24724 & ~n40513 ;
  assign n40573 = ~n40571 & ~n40572 ;
  assign n40574 = ~n40548 & ~n40573 ;
  assign n40575 = ~n20846 & n40486 ;
  assign n40576 = n30376 & ~n40484 ;
  assign n40577 = ~n40575 & ~n40576 ;
  assign n40578 = n20846 & ~n40337 ;
  assign n40579 = ~n20910 & ~n40578 ;
  assign n40580 = n40577 & n40579 ;
  assign n40581 = n21768 & n40156 ;
  assign n40582 = n21770 & n40156 ;
  assign n40583 = ~n21734 & n40582 ;
  assign n40584 = ~n40581 & ~n40583 ;
  assign n40585 = n31338 & n40584 ;
  assign n40586 = ~n23907 & ~n40491 ;
  assign n40587 = ~n40490 & n40586 ;
  assign n40588 = ~n40489 & n40587 ;
  assign n40589 = n40022 & ~n40337 ;
  assign n40590 = n20897 & n40584 ;
  assign n40591 = ~n40589 & n40590 ;
  assign n40592 = ~n40588 & n40591 ;
  assign n40593 = ~n40585 & ~n40592 ;
  assign n40594 = n21768 & n40151 ;
  assign n40595 = n21770 & n40151 ;
  assign n40596 = ~n21734 & n40595 ;
  assign n40597 = ~n40594 & ~n40596 ;
  assign n40598 = n40032 & n40597 ;
  assign n40599 = n20849 & n40597 ;
  assign n40600 = ~n40589 & n40599 ;
  assign n40601 = ~n40588 & n40600 ;
  assign n40602 = ~n40598 & ~n40601 ;
  assign n40603 = n40593 & n40602 ;
  assign n40604 = ~n40580 & n40603 ;
  assign n40605 = \pi0787  & ~n40604 ;
  assign n40606 = ~\pi0191  & \pi0644  ;
  assign n40607 = n21768 & n40606 ;
  assign n40608 = n21770 & n40606 ;
  assign n40609 = ~n21734 & n40608 ;
  assign n40610 = ~n40607 & ~n40609 ;
  assign n40611 = n23939 & n40610 ;
  assign n40612 = \pi0715  & n40610 ;
  assign n40613 = ~\pi0191  & ~n31367 ;
  assign n40614 = n21768 & n40613 ;
  assign n40615 = n21770 & n40613 ;
  assign n40616 = ~n21734 & n40615 ;
  assign n40617 = ~n40614 & ~n40616 ;
  assign n40618 = n40612 & n40617 ;
  assign n40619 = ~n40611 & ~n40618 ;
  assign n40620 = n31367 & ~n40611 ;
  assign n40621 = ~n40484 & n40620 ;
  assign n40622 = ~n40619 & ~n40621 ;
  assign n40623 = n31378 & ~n40622 ;
  assign n40624 = ~\pi0715  & n40617 ;
  assign n40625 = ~n23958 & ~n40624 ;
  assign n40626 = n31382 & ~n40484 ;
  assign n40627 = ~n40625 & ~n40626 ;
  assign n40628 = n26824 & ~n40627 ;
  assign n40629 = \pi0790  & ~n40628 ;
  assign n40630 = ~n40623 & n40629 ;
  assign n40631 = n9948 & ~n40630 ;
  assign n40632 = ~n40605 & n40631 ;
  assign n40633 = ~n40574 & n40632 ;
  assign n40634 = n23942 & n40337 ;
  assign n40635 = \pi0644  & ~n40634 ;
  assign n40636 = ~\pi0715  & ~n40635 ;
  assign n40637 = ~n23942 & ~n40589 ;
  assign n40638 = ~\pi0715  & n40637 ;
  assign n40639 = ~n40588 & n40638 ;
  assign n40640 = ~n40636 & ~n40639 ;
  assign n40641 = ~\pi1160  & ~n40622 ;
  assign n40642 = n40640 & n40641 ;
  assign n40643 = n9948 & n40642 ;
  assign n40644 = ~\pi0191  & ~\pi0644  ;
  assign n40645 = n21768 & n40644 ;
  assign n40646 = n21770 & n40644 ;
  assign n40647 = ~n21734 & n40646 ;
  assign n40648 = ~n40645 & ~n40647 ;
  assign n40649 = n40627 & n40648 ;
  assign n40650 = ~\pi0644  & ~n40634 ;
  assign n40651 = \pi0715  & ~n40650 ;
  assign n40652 = \pi0715  & n40637 ;
  assign n40653 = ~n40588 & n40652 ;
  assign n40654 = ~n40651 & ~n40653 ;
  assign n40655 = ~n40649 & n40654 ;
  assign n40656 = n31413 & n40655 ;
  assign n40657 = ~n40643 & ~n40656 ;
  assign n40658 = \pi0790  & ~n40657 ;
  assign n40659 = \pi0191  & ~\pi0832  ;
  assign n40660 = ~n21132 & ~n40659 ;
  assign n40661 = ~n40658 & ~n40660 ;
  assign n40662 = ~n40633 & n40661 ;
  assign n40663 = ~n40278 & ~n40662 ;
  assign n40664 = ~\pi0192  & \pi0788  ;
  assign n40665 = ~n1689 & n40664 ;
  assign n40666 = ~n20778 & n40665 ;
  assign n40667 = n20886 & n40666 ;
  assign n40668 = \pi0764  & n1689 ;
  assign n40669 = n20784 & n40668 ;
  assign n40670 = n22767 & n40669 ;
  assign n40671 = ~\pi0192  & ~n1689 ;
  assign n40672 = ~n40669 & ~n40671 ;
  assign n40673 = ~n20792 & ~n40672 ;
  assign n40674 = ~n40670 & n40673 ;
  assign n40675 = n20801 & ~n40674 ;
  assign n40676 = ~\pi1155  & ~n40671 ;
  assign n40677 = \pi0785  & n40676 ;
  assign n40678 = ~n40670 & n40677 ;
  assign n40679 = ~\pi0785  & ~n40671 ;
  assign n40680 = ~n40669 & n40679 ;
  assign n40681 = ~n20804 & ~n40680 ;
  assign n40682 = n29682 & n40681 ;
  assign n40683 = ~n40678 & n40682 ;
  assign n40684 = ~n40675 & n40683 ;
  assign n40685 = n30847 & n40684 ;
  assign n40686 = ~n40667 & ~n40685 ;
  assign n40687 = \pi0691  & n1689 ;
  assign n40688 = n20855 & n40687 ;
  assign n40689 = ~n40671 & ~n40688 ;
  assign n40690 = ~\pi0778  & ~n40689 ;
  assign n40691 = ~\pi0625  & \pi0691  ;
  assign n40692 = n1689 & n40691 ;
  assign n40693 = n20855 & n40692 ;
  assign n40694 = \pi1153  & n40693 ;
  assign n40695 = \pi1153  & ~n40671 ;
  assign n40696 = ~n40688 & n40695 ;
  assign n40697 = ~n40694 & ~n40696 ;
  assign n40698 = ~\pi1153  & ~n40671 ;
  assign n40699 = ~n40693 & n40698 ;
  assign n40700 = \pi0778  & ~n40699 ;
  assign n40701 = n40697 & n40700 ;
  assign n40702 = ~n40690 & ~n40701 ;
  assign n40703 = n26474 & ~n40702 ;
  assign n40704 = \pi0629  & ~n40703 ;
  assign n40705 = n40686 & n40704 ;
  assign n40706 = n20887 & n40666 ;
  assign n40707 = n32579 & n40684 ;
  assign n40708 = ~n40706 & ~n40707 ;
  assign n40709 = n26485 & ~n40702 ;
  assign n40710 = ~\pi0629  & ~n40709 ;
  assign n40711 = n40708 & n40710 ;
  assign n40712 = ~n40705 & ~n40711 ;
  assign n40713 = \pi0792  & n40712 ;
  assign n40714 = ~n21067 & ~n40713 ;
  assign n40715 = n39578 & ~n40702 ;
  assign n40716 = ~\pi0192  & ~\pi0647  ;
  assign n40717 = ~n1689 & n40716 ;
  assign n40718 = n20849 & ~n40717 ;
  assign n40719 = ~n40715 & n40718 ;
  assign n40720 = n26319 & ~n40702 ;
  assign n40721 = ~\pi0192  & \pi0647  ;
  assign n40722 = ~n1689 & n40721 ;
  assign n40723 = n20897 & ~n40722 ;
  assign n40724 = ~n40720 & n40723 ;
  assign n40725 = ~n40719 & ~n40724 ;
  assign n40726 = \pi0787  & ~n40725 ;
  assign n40727 = ~n20846 & n40666 ;
  assign n40728 = n30376 & n40684 ;
  assign n40729 = ~n40727 & ~n40728 ;
  assign n40730 = ~\pi0192  & \pi0792  ;
  assign n40731 = ~n1689 & n40730 ;
  assign n40732 = ~n20845 & n40731 ;
  assign n40733 = n32606 & ~n40732 ;
  assign n40734 = n40729 & n40733 ;
  assign n40735 = ~n40726 & ~n40734 ;
  assign n40736 = ~n24761 & n40735 ;
  assign n40737 = ~n40714 & n40736 ;
  assign n40738 = \pi0608  & ~n40699 ;
  assign n40739 = ~n40669 & n40695 ;
  assign n40740 = \pi0778  & ~n40739 ;
  assign n40741 = n26421 & ~n40689 ;
  assign n40742 = ~n40740 & ~n40741 ;
  assign n40743 = n40738 & ~n40742 ;
  assign n40744 = n26147 & ~n40689 ;
  assign n40745 = \pi0691  & ~n20784 ;
  assign n40746 = n22113 & n40745 ;
  assign n40747 = n40672 & ~n40746 ;
  assign n40748 = ~n40744 & ~n40747 ;
  assign n40749 = n40698 & ~n40748 ;
  assign n40750 = n26415 & n40697 ;
  assign n40751 = ~n40749 & n40750 ;
  assign n40752 = ~n40743 & ~n40751 ;
  assign n40753 = ~\pi1155  & ~n40690 ;
  assign n40754 = ~n40701 & n40753 ;
  assign n40755 = ~n20999 & ~n40754 ;
  assign n40756 = ~\pi0778  & ~n40747 ;
  assign n40757 = ~n40755 & ~n40756 ;
  assign n40758 = n40752 & n40757 ;
  assign n40759 = n29766 & ~n40690 ;
  assign n40760 = ~n40701 & n40759 ;
  assign n40761 = \pi1155  & ~n40674 ;
  assign n40762 = ~\pi0660  & ~n40761 ;
  assign n40763 = ~n40760 & n40762 ;
  assign n40764 = ~n40758 & n40763 ;
  assign n40765 = \pi0785  & ~n40764 ;
  assign n40766 = n29775 & n40681 ;
  assign n40767 = ~n40678 & n40766 ;
  assign n40768 = ~n40675 & n40767 ;
  assign n40769 = n29779 & ~n40702 ;
  assign n40770 = ~n40768 & ~n40769 ;
  assign n40771 = \pi0781  & ~n40770 ;
  assign n40772 = \pi1155  & ~n40690 ;
  assign n40773 = ~n40701 & n40772 ;
  assign n40774 = ~n21774 & ~n40773 ;
  assign n40775 = ~n40756 & ~n40774 ;
  assign n40776 = n40752 & n40775 ;
  assign n40777 = n26121 & ~n40690 ;
  assign n40778 = ~n40701 & n40777 ;
  assign n40779 = \pi0660  & ~n40676 ;
  assign n40780 = \pi0660  & n40669 ;
  assign n40781 = n22767 & n40780 ;
  assign n40782 = ~n40779 & ~n40781 ;
  assign n40783 = ~n40778 & ~n40782 ;
  assign n40784 = ~n40776 & n40783 ;
  assign n40785 = ~n40771 & ~n40784 ;
  assign n40786 = n40765 & n40785 ;
  assign n40787 = ~\pi0785  & ~n40756 ;
  assign n40788 = ~n40743 & n40787 ;
  assign n40789 = ~n40751 & n40788 ;
  assign n40790 = n21022 & ~n40789 ;
  assign n40791 = ~n40771 & ~n40790 ;
  assign n40792 = n29803 & ~n40791 ;
  assign n40793 = ~n40786 & n40792 ;
  assign n40794 = n29808 & n40681 ;
  assign n40795 = ~n40678 & n40794 ;
  assign n40796 = ~n40675 & n40795 ;
  assign n40797 = n30966 & ~n40702 ;
  assign n40798 = ~n40796 & ~n40797 ;
  assign n40799 = n36155 & ~n40798 ;
  assign n40800 = \pi0626  & ~n40684 ;
  assign n40801 = ~\pi0626  & ~n40671 ;
  assign n40802 = n20881 & ~n40801 ;
  assign n40803 = ~n40800 & n40802 ;
  assign n40804 = n26458 & ~n40702 ;
  assign n40805 = ~\pi0626  & ~n40684 ;
  assign n40806 = \pi0626  & ~n40671 ;
  assign n40807 = n20882 & ~n40806 ;
  assign n40808 = ~n40805 & n40807 ;
  assign n40809 = ~n40804 & ~n40808 ;
  assign n40810 = ~n40803 & n40809 ;
  assign n40811 = \pi0788  & ~n40810 ;
  assign n40812 = ~n40799 & ~n40811 ;
  assign n40813 = ~n40793 & n40812 ;
  assign n40814 = ~n23856 & n40736 ;
  assign n40815 = ~n40813 & n40814 ;
  assign n40816 = ~n40737 & ~n40815 ;
  assign n40817 = n30987 & ~n40729 ;
  assign n40818 = n23312 & n40817 ;
  assign n40819 = \pi1157  & ~n40717 ;
  assign n40820 = ~n40715 & n40819 ;
  assign n40821 = ~\pi1157  & ~n40722 ;
  assign n40822 = ~n40720 & n40821 ;
  assign n40823 = ~n40820 & ~n40822 ;
  assign n40824 = \pi0787  & ~n40823 ;
  assign n40825 = n26333 & ~n40702 ;
  assign n40826 = ~\pi0787  & ~n40825 ;
  assign n40827 = ~\pi1160  & ~n40826 ;
  assign n40828 = n23312 & n40827 ;
  assign n40829 = ~n40824 & n40828 ;
  assign n40830 = ~n40818 & ~n40829 ;
  assign n40831 = ~n23414 & n40671 ;
  assign n40832 = ~n24886 & n40831 ;
  assign n40833 = ~n23313 & ~n40832 ;
  assign n40834 = \pi1160  & ~n40826 ;
  assign n40835 = ~n40824 & n40834 ;
  assign n40836 = n31010 & ~n40729 ;
  assign n40837 = ~n40832 & ~n40836 ;
  assign n40838 = ~n40835 & n40837 ;
  assign n40839 = ~n40833 & ~n40838 ;
  assign n40840 = n40830 & ~n40839 ;
  assign n40841 = \pi0790  & ~n40840 ;
  assign n40842 = \pi0832  & ~n40841 ;
  assign n40843 = n40816 & n40842 ;
  assign n40844 = \pi0192  & ~n6861 ;
  assign n40845 = ~\pi0192  & ~\pi0691  ;
  assign n40846 = ~\pi0038  & n40845 ;
  assign n40847 = n21743 & n40846 ;
  assign n40848 = ~n21734 & n40847 ;
  assign n40849 = \pi0038  & n40845 ;
  assign n40850 = ~n22123 & n40849 ;
  assign n40851 = n6861 & ~n40850 ;
  assign n40852 = ~n40848 & n40851 ;
  assign n40853 = ~n40844 & ~n40852 ;
  assign n40854 = ~\pi0192  & ~n22017 ;
  assign n40855 = ~n21994 & n40854 ;
  assign n40856 = ~\pi0038  & ~\pi0192  ;
  assign n40857 = ~n22109 & ~n40856 ;
  assign n40858 = ~n40855 & ~n40857 ;
  assign n40859 = ~\pi0192  & ~n21757 ;
  assign n40860 = n22117 & ~n40859 ;
  assign n40861 = \pi0691  & ~n40844 ;
  assign n40862 = ~n40860 & n40861 ;
  assign n40863 = ~n40858 & n40862 ;
  assign n40864 = ~n40853 & ~n40863 ;
  assign n40865 = ~\pi0778  & n40864 ;
  assign n40866 = ~\pi0192  & \pi0764  ;
  assign n40867 = ~n21467 & n40866 ;
  assign n40868 = ~\pi0039  & n40866 ;
  assign n40869 = n21272 & n40868 ;
  assign n40870 = ~n40867 & ~n40869 ;
  assign n40871 = \pi0764  & n21484 ;
  assign n40872 = ~\pi0192  & n21743 ;
  assign n40873 = ~n40866 & ~n40872 ;
  assign n40874 = ~n40871 & n40873 ;
  assign n40875 = n40870 & ~n40874 ;
  assign n40876 = ~\pi0038  & ~n40875 ;
  assign n40877 = ~\pi0764  & ~n21731 ;
  assign n40878 = n21714 & n40877 ;
  assign n40879 = ~n21693 & n40878 ;
  assign n40880 = \pi0192  & ~n21543 ;
  assign n40881 = \pi0192  & n21562 ;
  assign n40882 = ~n21552 & n40881 ;
  assign n40883 = ~n40880 & ~n40882 ;
  assign n40884 = ~n21536 & ~n40883 ;
  assign n40885 = ~n40879 & ~n40884 ;
  assign n40886 = n9627 & ~n40885 ;
  assign n40887 = n8413 & n40669 ;
  assign n40888 = n1354 & n40887 ;
  assign n40889 = n1358 & n40888 ;
  assign n40890 = \pi0038  & ~n40889 ;
  assign n40891 = ~n40859 & n40890 ;
  assign n40892 = ~n40844 & ~n40891 ;
  assign n40893 = ~n40886 & n40892 ;
  assign n40894 = ~n40876 & n40893 ;
  assign n40895 = ~\pi0192  & ~n6861 ;
  assign n40896 = ~\pi1155  & ~n40895 ;
  assign n40897 = n22767 & n40896 ;
  assign n40898 = ~n40894 & n40897 ;
  assign n40899 = ~\pi0192  & n21768 ;
  assign n40900 = ~\pi0192  & n21770 ;
  assign n40901 = ~n21734 & n40900 ;
  assign n40902 = ~n40899 & ~n40901 ;
  assign n40903 = ~n32768 & n40902 ;
  assign n40904 = ~n22787 & ~n40903 ;
  assign n40905 = ~n40898 & n40904 ;
  assign n40906 = n40865 & ~n40905 ;
  assign n40907 = \pi0625  & ~n40864 ;
  assign n40908 = ~\pi0192  & ~\pi0625  ;
  assign n40909 = n21768 & n40908 ;
  assign n40910 = n21770 & n40908 ;
  assign n40911 = ~n21734 & n40910 ;
  assign n40912 = ~n40909 & ~n40911 ;
  assign n40913 = \pi1153  & n40912 ;
  assign n40914 = ~n40907 & n40913 ;
  assign n40915 = ~\pi0625  & ~n40864 ;
  assign n40916 = ~\pi0192  & \pi0625  ;
  assign n40917 = n21768 & n40916 ;
  assign n40918 = n21770 & n40916 ;
  assign n40919 = ~n21734 & n40918 ;
  assign n40920 = ~n40917 & ~n40919 ;
  assign n40921 = ~\pi1153  & n40920 ;
  assign n40922 = ~n40915 & n40921 ;
  assign n40923 = ~n40914 & ~n40922 ;
  assign n40924 = \pi0778  & ~n40905 ;
  assign n40925 = ~n40923 & n40924 ;
  assign n40926 = ~n40906 & ~n40925 ;
  assign n40927 = n39791 & ~n40926 ;
  assign n40928 = n31109 & ~n40923 ;
  assign n40929 = n22767 & ~n40895 ;
  assign n40930 = ~n40894 & n40929 ;
  assign n40931 = ~n22767 & n40902 ;
  assign n40932 = \pi0660  & ~n40931 ;
  assign n40933 = ~n40930 & n40932 ;
  assign n40934 = ~n22766 & ~n40933 ;
  assign n40935 = n39367 & n40864 ;
  assign n40936 = ~n40934 & ~n40935 ;
  assign n40937 = ~n40928 & n40936 ;
  assign n40938 = n22788 & ~n40895 ;
  assign n40939 = ~n40894 & n40938 ;
  assign n40940 = ~n22788 & n40902 ;
  assign n40941 = ~\pi0660  & ~n40940 ;
  assign n40942 = ~n40939 & n40941 ;
  assign n40943 = n31121 & ~n40942 ;
  assign n40944 = ~n40937 & n40943 ;
  assign n40945 = ~n40927 & ~n40944 ;
  assign n40946 = n26700 & ~n40945 ;
  assign n40947 = \pi0778  & ~n40923 ;
  assign n40948 = \pi0609  & ~n40865 ;
  assign n40949 = ~n40947 & n40948 ;
  assign n40950 = ~n40905 & ~n40949 ;
  assign n40951 = n39816 & ~n40942 ;
  assign n40952 = \pi0785  & ~n40951 ;
  assign n40953 = ~n40950 & n40952 ;
  assign n40954 = ~\pi0691  & ~n40891 ;
  assign n40955 = ~n40886 & n40954 ;
  assign n40956 = ~n40876 & n40955 ;
  assign n40957 = n6861 & ~n40956 ;
  assign n40958 = ~n22734 & ~n40908 ;
  assign n40959 = ~n40957 & ~n40958 ;
  assign n40960 = ~\pi0039  & ~\pi0192  ;
  assign n40961 = ~n22683 & n40960 ;
  assign n40962 = ~\pi0192  & ~n23548 ;
  assign n40963 = \pi0764  & ~n40962 ;
  assign n40964 = ~n40961 & n40963 ;
  assign n40965 = \pi0192  & ~n23558 ;
  assign n40966 = n23557 & n40965 ;
  assign n40967 = ~\pi0038  & ~n40966 ;
  assign n40968 = n40964 & n40967 ;
  assign n40969 = ~\pi0192  & ~n23568 ;
  assign n40970 = \pi0192  & n23575 ;
  assign n40971 = n23572 & n40970 ;
  assign n40972 = ~\pi0038  & ~\pi0764  ;
  assign n40973 = ~n40971 & n40972 ;
  assign n40974 = ~n40969 & n40973 ;
  assign n40975 = ~n40968 & ~n40974 ;
  assign n40976 = \pi0192  & \pi0603  ;
  assign n40977 = ~n20783 & n40976 ;
  assign n40978 = n40668 & n40977 ;
  assign n40979 = \pi0192  & \pi0680  ;
  assign n40980 = ~n20854 & n40979 ;
  assign n40981 = ~n20784 & n40980 ;
  assign n40982 = n1689 & n40981 ;
  assign n40983 = ~n40978 & ~n40982 ;
  assign n40984 = n26554 & ~n40983 ;
  assign n40985 = n1358 & n40984 ;
  assign n40986 = \pi0038  & ~n40985 ;
  assign n40987 = \pi0691  & ~n40986 ;
  assign n40988 = \pi0764  & ~n22317 ;
  assign n40989 = ~n31169 & ~n40988 ;
  assign n40990 = ~\pi0039  & n40989 ;
  assign n40991 = n21289 & n40990 ;
  assign n40992 = ~\pi0192  & \pi0691  ;
  assign n40993 = ~n40991 & n40992 ;
  assign n40994 = ~n40987 & ~n40993 ;
  assign n40995 = ~n40958 & ~n40994 ;
  assign n40996 = n40975 & n40995 ;
  assign n40997 = ~n40959 & ~n40996 ;
  assign n40998 = ~\pi1153  & ~n40895 ;
  assign n40999 = ~n40894 & n40998 ;
  assign n41000 = ~n24561 & ~n40999 ;
  assign n41001 = n40997 & ~n41000 ;
  assign n41002 = ~\pi0608  & ~n40913 ;
  assign n41003 = n22755 & ~n40864 ;
  assign n41004 = ~n41002 & ~n41003 ;
  assign n41005 = ~n41001 & ~n41004 ;
  assign n41006 = ~n22727 & ~n40916 ;
  assign n41007 = ~n40957 & ~n41006 ;
  assign n41008 = ~n40994 & ~n41006 ;
  assign n41009 = n40975 & n41008 ;
  assign n41010 = ~n41007 & ~n41009 ;
  assign n41011 = \pi1153  & ~n40895 ;
  assign n41012 = ~n40894 & n41011 ;
  assign n41013 = ~n24550 & ~n41012 ;
  assign n41014 = n41010 & ~n41013 ;
  assign n41015 = \pi0608  & ~n40921 ;
  assign n41016 = n22740 & ~n40864 ;
  assign n41017 = ~n41015 & ~n41016 ;
  assign n41018 = ~n41014 & ~n41017 ;
  assign n41019 = ~n41005 & ~n41018 ;
  assign n41020 = \pi0778  & ~n41019 ;
  assign n41021 = ~n40953 & ~n41020 ;
  assign n41022 = ~\pi0192  & ~\pi0778  ;
  assign n41023 = ~n23622 & ~n41022 ;
  assign n41024 = ~n40957 & ~n41023 ;
  assign n41025 = ~n40994 & ~n41023 ;
  assign n41026 = n40975 & n41025 ;
  assign n41027 = ~n41024 & ~n41026 ;
  assign n41028 = n26700 & n41027 ;
  assign n41029 = n41021 & n41028 ;
  assign n41030 = ~n40946 & ~n41029 ;
  assign n41031 = ~\pi0192  & ~n20811 ;
  assign n41032 = n21768 & n41031 ;
  assign n41033 = n21770 & n41031 ;
  assign n41034 = ~n21734 & n41033 ;
  assign n41035 = ~n41032 & ~n41034 ;
  assign n41036 = n23424 & ~n41035 ;
  assign n41037 = n21777 & ~n40895 ;
  assign n41038 = ~n40894 & n41037 ;
  assign n41039 = ~n21777 & n40902 ;
  assign n41040 = n20811 & ~n41039 ;
  assign n41041 = n23424 & n41040 ;
  assign n41042 = ~n41038 & n41041 ;
  assign n41043 = ~n41036 & ~n41042 ;
  assign n41044 = ~\pi0781  & ~n41039 ;
  assign n41045 = ~n23423 & n41044 ;
  assign n41046 = ~n41038 & n41045 ;
  assign n41047 = n23423 & ~n40902 ;
  assign n41048 = ~n41046 & ~n41047 ;
  assign n41049 = n41043 & n41048 ;
  assign n41050 = ~n23880 & ~n41049 ;
  assign n41051 = n23880 & ~n40902 ;
  assign n41052 = n24691 & ~n41051 ;
  assign n41053 = ~n41050 & n41052 ;
  assign n41054 = n26065 & ~n40923 ;
  assign n41055 = n26739 & n40864 ;
  assign n41056 = ~n23885 & n40902 ;
  assign n41057 = \pi0628  & ~n41056 ;
  assign n41058 = ~n41055 & n41057 ;
  assign n41059 = ~n41054 & n41058 ;
  assign n41060 = ~\pi0192  & ~\pi0628  ;
  assign n41061 = n21768 & n41060 ;
  assign n41062 = n21770 & n41060 ;
  assign n41063 = ~n21734 & n41062 ;
  assign n41064 = ~n41061 & ~n41063 ;
  assign n41065 = n20843 & n41064 ;
  assign n41066 = ~n41059 & n41065 ;
  assign n41067 = ~\pi0628  & ~n41056 ;
  assign n41068 = ~n41055 & n41067 ;
  assign n41069 = ~n41054 & n41068 ;
  assign n41070 = ~\pi0192  & \pi0628  ;
  assign n41071 = n21768 & n41070 ;
  assign n41072 = n21770 & n41070 ;
  assign n41073 = ~n21734 & n41072 ;
  assign n41074 = ~n41071 & ~n41073 ;
  assign n41075 = n20844 & n41074 ;
  assign n41076 = ~n41069 & n41075 ;
  assign n41077 = ~n41066 & ~n41076 ;
  assign n41078 = ~n41053 & n41077 ;
  assign n41079 = \pi0792  & ~n41078 ;
  assign n41080 = ~n41038 & n41040 ;
  assign n41081 = n22155 & n41035 ;
  assign n41082 = ~n41080 & n41081 ;
  assign n41083 = ~n22147 & ~n40865 ;
  assign n41084 = n22147 & ~n40902 ;
  assign n41085 = n39952 & ~n41084 ;
  assign n41086 = ~n41083 & n41085 ;
  assign n41087 = \pi0778  & n41085 ;
  assign n41088 = ~n40923 & n41087 ;
  assign n41089 = ~n41086 & ~n41088 ;
  assign n41090 = ~n41082 & n41089 ;
  assign n41091 = ~n21034 & ~n41090 ;
  assign n41092 = n30780 & ~n40923 ;
  assign n41093 = n31274 & n40864 ;
  assign n41094 = ~n23380 & n40902 ;
  assign n41095 = ~n41093 & ~n41094 ;
  assign n41096 = ~n41092 & n41095 ;
  assign n41097 = ~n31283 & ~n41096 ;
  assign n41098 = n23683 & ~n41035 ;
  assign n41099 = n23683 & n41040 ;
  assign n41100 = ~n41038 & n41099 ;
  assign n41101 = ~n41098 & ~n41100 ;
  assign n41102 = n21032 & n41044 ;
  assign n41103 = ~n41038 & n41102 ;
  assign n41104 = ~n21032 & ~n40902 ;
  assign n41105 = ~n20876 & ~n41104 ;
  assign n41106 = \pi0789  & n41105 ;
  assign n41107 = ~n41103 & n41106 ;
  assign n41108 = n41101 & n41107 ;
  assign n41109 = ~n21038 & ~n41108 ;
  assign n41110 = ~n41097 & n41109 ;
  assign n41111 = ~n41091 & n41110 ;
  assign n41112 = ~n41079 & n41111 ;
  assign n41113 = n41030 & n41112 ;
  assign n41114 = n20951 & ~n40902 ;
  assign n41115 = ~n31301 & ~n41114 ;
  assign n41116 = ~n41093 & ~n41115 ;
  assign n41117 = ~n41092 & n41116 ;
  assign n41118 = n31306 & ~n40902 ;
  assign n41119 = ~n23856 & ~n41118 ;
  assign n41120 = ~n41117 & n41119 ;
  assign n41121 = ~\pi0626  & ~n41047 ;
  assign n41122 = ~n41046 & n41121 ;
  assign n41123 = n41043 & n41122 ;
  assign n41124 = \pi0626  & n40902 ;
  assign n41125 = n20882 & ~n41124 ;
  assign n41126 = ~n41123 & n41125 ;
  assign n41127 = \pi0626  & ~n41047 ;
  assign n41128 = ~n41046 & n41127 ;
  assign n41129 = n41043 & n41128 ;
  assign n41130 = ~\pi0626  & n40902 ;
  assign n41131 = n20881 & ~n41130 ;
  assign n41132 = ~n41129 & n41131 ;
  assign n41133 = ~n41126 & ~n41132 ;
  assign n41134 = n41120 & n41133 ;
  assign n41135 = ~n26803 & ~n41134 ;
  assign n41136 = ~n21067 & ~n41135 ;
  assign n41137 = n24724 & ~n41078 ;
  assign n41138 = ~n41136 & ~n41137 ;
  assign n41139 = ~n41113 & ~n41138 ;
  assign n41140 = ~n20846 & n41051 ;
  assign n41141 = n30376 & ~n41049 ;
  assign n41142 = ~n41140 & ~n41141 ;
  assign n41143 = n20846 & ~n40902 ;
  assign n41144 = ~n20910 & ~n41143 ;
  assign n41145 = n41142 & n41144 ;
  assign n41146 = n21768 & n40721 ;
  assign n41147 = n21770 & n40721 ;
  assign n41148 = ~n21734 & n41147 ;
  assign n41149 = ~n41146 & ~n41148 ;
  assign n41150 = n31338 & n41149 ;
  assign n41151 = ~n23907 & ~n41056 ;
  assign n41152 = ~n41055 & n41151 ;
  assign n41153 = ~n41054 & n41152 ;
  assign n41154 = n40022 & ~n40902 ;
  assign n41155 = n20897 & n41149 ;
  assign n41156 = ~n41154 & n41155 ;
  assign n41157 = ~n41153 & n41156 ;
  assign n41158 = ~n41150 & ~n41157 ;
  assign n41159 = n21768 & n40716 ;
  assign n41160 = n21770 & n40716 ;
  assign n41161 = ~n21734 & n41160 ;
  assign n41162 = ~n41159 & ~n41161 ;
  assign n41163 = n40032 & n41162 ;
  assign n41164 = n20849 & n41162 ;
  assign n41165 = ~n41154 & n41164 ;
  assign n41166 = ~n41153 & n41165 ;
  assign n41167 = ~n41163 & ~n41166 ;
  assign n41168 = n41158 & n41167 ;
  assign n41169 = ~n41145 & n41168 ;
  assign n41170 = \pi0787  & ~n41169 ;
  assign n41171 = ~\pi0192  & \pi0644  ;
  assign n41172 = n21768 & n41171 ;
  assign n41173 = n21770 & n41171 ;
  assign n41174 = ~n21734 & n41173 ;
  assign n41175 = ~n41172 & ~n41174 ;
  assign n41176 = n23939 & n41175 ;
  assign n41177 = \pi0715  & n41175 ;
  assign n41178 = ~\pi0192  & ~n31367 ;
  assign n41179 = n21768 & n41178 ;
  assign n41180 = n21770 & n41178 ;
  assign n41181 = ~n21734 & n41180 ;
  assign n41182 = ~n41179 & ~n41181 ;
  assign n41183 = n41177 & n41182 ;
  assign n41184 = ~n41176 & ~n41183 ;
  assign n41185 = n31367 & ~n41176 ;
  assign n41186 = ~n41049 & n41185 ;
  assign n41187 = ~n41184 & ~n41186 ;
  assign n41188 = n31378 & ~n41187 ;
  assign n41189 = ~\pi0715  & n41182 ;
  assign n41190 = ~n23958 & ~n41189 ;
  assign n41191 = n31382 & ~n41049 ;
  assign n41192 = ~n41190 & ~n41191 ;
  assign n41193 = n26824 & ~n41192 ;
  assign n41194 = \pi0790  & ~n41193 ;
  assign n41195 = ~n41188 & n41194 ;
  assign n41196 = n9948 & ~n41195 ;
  assign n41197 = ~n41170 & n41196 ;
  assign n41198 = ~n41139 & n41197 ;
  assign n41199 = n23942 & n40902 ;
  assign n41200 = \pi0644  & ~n41199 ;
  assign n41201 = ~\pi0715  & ~n41200 ;
  assign n41202 = ~n23942 & ~n41154 ;
  assign n41203 = ~\pi0715  & n41202 ;
  assign n41204 = ~n41153 & n41203 ;
  assign n41205 = ~n41201 & ~n41204 ;
  assign n41206 = ~\pi1160  & ~n41187 ;
  assign n41207 = n41205 & n41206 ;
  assign n41208 = n9948 & n41207 ;
  assign n41209 = ~\pi0192  & ~\pi0644  ;
  assign n41210 = n21768 & n41209 ;
  assign n41211 = n21770 & n41209 ;
  assign n41212 = ~n21734 & n41211 ;
  assign n41213 = ~n41210 & ~n41212 ;
  assign n41214 = n41192 & n41213 ;
  assign n41215 = ~\pi0644  & ~n41199 ;
  assign n41216 = \pi0715  & ~n41215 ;
  assign n41217 = \pi0715  & n41202 ;
  assign n41218 = ~n41153 & n41217 ;
  assign n41219 = ~n41216 & ~n41218 ;
  assign n41220 = ~n41214 & n41219 ;
  assign n41221 = n31413 & n41220 ;
  assign n41222 = ~n41208 & ~n41221 ;
  assign n41223 = \pi0790  & ~n41222 ;
  assign n41224 = \pi0192  & ~\pi0832  ;
  assign n41225 = ~n21132 & ~n41224 ;
  assign n41226 = ~n41223 & ~n41225 ;
  assign n41227 = ~n41198 & n41226 ;
  assign n41228 = ~n40843 & ~n41227 ;
  assign n41229 = ~\pi0193  & \pi0788  ;
  assign n41230 = ~n1689 & n41229 ;
  assign n41231 = ~n20778 & n41230 ;
  assign n41232 = n20886 & n41231 ;
  assign n41233 = \pi0739  & n1689 ;
  assign n41234 = n20784 & n41233 ;
  assign n41235 = n22767 & n41234 ;
  assign n41236 = ~\pi0193  & ~n1689 ;
  assign n41237 = ~n41234 & ~n41236 ;
  assign n41238 = ~n20792 & ~n41237 ;
  assign n41239 = ~n41235 & n41238 ;
  assign n41240 = n20801 & ~n41239 ;
  assign n41241 = ~\pi1155  & ~n41236 ;
  assign n41242 = \pi0785  & n41241 ;
  assign n41243 = ~n41235 & n41242 ;
  assign n41244 = ~\pi0785  & ~n41236 ;
  assign n41245 = ~n41234 & n41244 ;
  assign n41246 = ~n20804 & ~n41245 ;
  assign n41247 = n29682 & n41246 ;
  assign n41248 = ~n41243 & n41247 ;
  assign n41249 = ~n41240 & n41248 ;
  assign n41250 = n30847 & n41249 ;
  assign n41251 = ~n41232 & ~n41250 ;
  assign n41252 = \pi0690  & n1689 ;
  assign n41253 = n20855 & n41252 ;
  assign n41254 = ~n41236 & ~n41253 ;
  assign n41255 = ~\pi0778  & ~n41254 ;
  assign n41256 = ~\pi0625  & \pi0690  ;
  assign n41257 = n1689 & n41256 ;
  assign n41258 = n20855 & n41257 ;
  assign n41259 = \pi1153  & n41258 ;
  assign n41260 = \pi1153  & ~n41236 ;
  assign n41261 = ~n41253 & n41260 ;
  assign n41262 = ~n41259 & ~n41261 ;
  assign n41263 = ~\pi1153  & ~n41236 ;
  assign n41264 = ~n41258 & n41263 ;
  assign n41265 = \pi0778  & ~n41264 ;
  assign n41266 = n41262 & n41265 ;
  assign n41267 = ~n41255 & ~n41266 ;
  assign n41268 = n26474 & ~n41267 ;
  assign n41269 = \pi0629  & ~n41268 ;
  assign n41270 = n41251 & n41269 ;
  assign n41271 = n20887 & n41231 ;
  assign n41272 = n32579 & n41249 ;
  assign n41273 = ~n41271 & ~n41272 ;
  assign n41274 = n26485 & ~n41267 ;
  assign n41275 = ~\pi0629  & ~n41274 ;
  assign n41276 = n41273 & n41275 ;
  assign n41277 = \pi0792  & ~n41276 ;
  assign n41278 = ~n41270 & n41277 ;
  assign n41279 = ~n21067 & ~n41278 ;
  assign n41280 = n39578 & ~n41267 ;
  assign n41281 = ~\pi0193  & ~\pi0647  ;
  assign n41282 = ~n1689 & n41281 ;
  assign n41283 = n20849 & ~n41282 ;
  assign n41284 = ~n41280 & n41283 ;
  assign n41285 = n26319 & ~n41267 ;
  assign n41286 = ~\pi0193  & \pi0647  ;
  assign n41287 = ~n1689 & n41286 ;
  assign n41288 = n20897 & ~n41287 ;
  assign n41289 = ~n41285 & n41288 ;
  assign n41290 = ~n41284 & ~n41289 ;
  assign n41291 = \pi0787  & ~n41290 ;
  assign n41292 = ~n20846 & n41231 ;
  assign n41293 = n30376 & n41249 ;
  assign n41294 = ~n41292 & ~n41293 ;
  assign n41295 = ~\pi0193  & \pi0792  ;
  assign n41296 = ~n1689 & n41295 ;
  assign n41297 = ~n20845 & n41296 ;
  assign n41298 = n32606 & ~n41297 ;
  assign n41299 = n41294 & n41298 ;
  assign n41300 = ~n41291 & ~n41299 ;
  assign n41301 = ~n24761 & n41300 ;
  assign n41302 = ~n41279 & n41301 ;
  assign n41303 = \pi0608  & ~n41264 ;
  assign n41304 = ~n41234 & n41260 ;
  assign n41305 = \pi0778  & ~n41304 ;
  assign n41306 = n26421 & ~n41254 ;
  assign n41307 = ~n41305 & ~n41306 ;
  assign n41308 = n41303 & ~n41307 ;
  assign n41309 = n26147 & ~n41254 ;
  assign n41310 = \pi0690  & ~n20784 ;
  assign n41311 = n22113 & n41310 ;
  assign n41312 = n41237 & ~n41311 ;
  assign n41313 = ~n41309 & ~n41312 ;
  assign n41314 = n41263 & ~n41313 ;
  assign n41315 = n26415 & n41262 ;
  assign n41316 = ~n41314 & n41315 ;
  assign n41317 = ~n41308 & ~n41316 ;
  assign n41318 = ~\pi1155  & ~n41255 ;
  assign n41319 = ~n41266 & n41318 ;
  assign n41320 = ~n20999 & ~n41319 ;
  assign n41321 = ~\pi0778  & ~n41312 ;
  assign n41322 = ~n41320 & ~n41321 ;
  assign n41323 = n41317 & n41322 ;
  assign n41324 = n29766 & ~n41255 ;
  assign n41325 = ~n41266 & n41324 ;
  assign n41326 = \pi1155  & ~n41239 ;
  assign n41327 = ~\pi0660  & ~n41326 ;
  assign n41328 = ~n41325 & n41327 ;
  assign n41329 = ~n41323 & n41328 ;
  assign n41330 = \pi0785  & ~n41329 ;
  assign n41331 = n29775 & n41246 ;
  assign n41332 = ~n41243 & n41331 ;
  assign n41333 = ~n41240 & n41332 ;
  assign n41334 = n29779 & ~n41267 ;
  assign n41335 = ~n41333 & ~n41334 ;
  assign n41336 = \pi0781  & ~n41335 ;
  assign n41337 = \pi1155  & ~n41255 ;
  assign n41338 = ~n41266 & n41337 ;
  assign n41339 = ~n21774 & ~n41338 ;
  assign n41340 = ~n41321 & ~n41339 ;
  assign n41341 = n41317 & n41340 ;
  assign n41342 = n26121 & ~n41255 ;
  assign n41343 = ~n41266 & n41342 ;
  assign n41344 = \pi0660  & ~n41241 ;
  assign n41345 = \pi0660  & n41234 ;
  assign n41346 = n22767 & n41345 ;
  assign n41347 = ~n41344 & ~n41346 ;
  assign n41348 = ~n41343 & ~n41347 ;
  assign n41349 = ~n41341 & n41348 ;
  assign n41350 = ~n41336 & ~n41349 ;
  assign n41351 = n41330 & n41350 ;
  assign n41352 = ~\pi0785  & ~n41321 ;
  assign n41353 = ~n41308 & n41352 ;
  assign n41354 = ~n41316 & n41353 ;
  assign n41355 = n21022 & ~n41354 ;
  assign n41356 = ~n41336 & ~n41355 ;
  assign n41357 = n29803 & ~n41356 ;
  assign n41358 = ~n41351 & n41357 ;
  assign n41359 = n30966 & ~n41267 ;
  assign n41360 = n29808 & n41246 ;
  assign n41361 = ~n41243 & n41360 ;
  assign n41362 = ~n41240 & n41361 ;
  assign n41363 = ~n41359 & ~n41362 ;
  assign n41364 = n36155 & ~n41363 ;
  assign n41365 = \pi0626  & ~n41249 ;
  assign n41366 = ~\pi0626  & ~n41236 ;
  assign n41367 = n20881 & ~n41366 ;
  assign n41368 = ~n41365 & n41367 ;
  assign n41369 = n26458 & ~n41267 ;
  assign n41370 = ~\pi0626  & ~n41249 ;
  assign n41371 = \pi0626  & ~n41236 ;
  assign n41372 = n20882 & ~n41371 ;
  assign n41373 = ~n41370 & n41372 ;
  assign n41374 = ~n41369 & ~n41373 ;
  assign n41375 = ~n41368 & n41374 ;
  assign n41376 = \pi0788  & ~n41375 ;
  assign n41377 = ~n41364 & ~n41376 ;
  assign n41378 = ~n41358 & n41377 ;
  assign n41379 = ~n23856 & n41301 ;
  assign n41380 = ~n41378 & n41379 ;
  assign n41381 = ~n41302 & ~n41380 ;
  assign n41382 = n30987 & ~n41294 ;
  assign n41383 = n23312 & n41382 ;
  assign n41384 = \pi1157  & ~n41282 ;
  assign n41385 = ~n41280 & n41384 ;
  assign n41386 = ~\pi1157  & ~n41287 ;
  assign n41387 = ~n41285 & n41386 ;
  assign n41388 = ~n41385 & ~n41387 ;
  assign n41389 = \pi0787  & ~n41388 ;
  assign n41390 = n26333 & ~n41267 ;
  assign n41391 = ~\pi0787  & ~n41390 ;
  assign n41392 = ~\pi1160  & ~n41391 ;
  assign n41393 = n23312 & n41392 ;
  assign n41394 = ~n41389 & n41393 ;
  assign n41395 = ~n41383 & ~n41394 ;
  assign n41396 = ~n23414 & n41236 ;
  assign n41397 = ~n24886 & n41396 ;
  assign n41398 = ~n23313 & ~n41397 ;
  assign n41399 = \pi1160  & ~n41391 ;
  assign n41400 = ~n41389 & n41399 ;
  assign n41401 = n31010 & ~n41294 ;
  assign n41402 = ~n41397 & ~n41401 ;
  assign n41403 = ~n41400 & n41402 ;
  assign n41404 = ~n41398 & ~n41403 ;
  assign n41405 = n41395 & ~n41404 ;
  assign n41406 = \pi0790  & ~n41405 ;
  assign n41407 = \pi0832  & ~n41406 ;
  assign n41408 = n41381 & n41407 ;
  assign n41409 = \pi0193  & ~\pi0832  ;
  assign n41410 = ~n21132 & ~n41409 ;
  assign n41411 = ~n41408 & n41410 ;
  assign n41412 = n9948 & ~n41408 ;
  assign n41413 = ~n41411 & ~n41412 ;
  assign n41414 = \pi0038  & n41234 ;
  assign n41415 = n8413 & n41414 ;
  assign n41416 = n1354 & n41415 ;
  assign n41417 = n1358 & n41416 ;
  assign n41418 = \pi0038  & ~\pi0193  ;
  assign n41419 = ~n21757 & n41418 ;
  assign n41420 = ~n41417 & ~n41419 ;
  assign n41421 = \pi0038  & n41420 ;
  assign n41422 = ~\pi0193  & ~n21467 ;
  assign n41423 = ~\pi0039  & ~\pi0193  ;
  assign n41424 = n21272 & n41423 ;
  assign n41425 = ~n41422 & ~n41424 ;
  assign n41426 = ~\pi0193  & \pi0739  ;
  assign n41427 = \pi0739  & n25023 ;
  assign n41428 = ~n41426 & ~n41427 ;
  assign n41429 = n41425 & ~n41428 ;
  assign n41430 = ~\pi0193  & ~\pi0739  ;
  assign n41431 = n21743 & n41430 ;
  assign n41432 = ~n21734 & n41431 ;
  assign n41433 = n41420 & ~n41432 ;
  assign n41434 = ~n41429 & n41433 ;
  assign n41435 = ~n41421 & ~n41434 ;
  assign n41436 = ~\pi0690  & n41435 ;
  assign n41437 = ~\pi0193  & ~\pi0778  ;
  assign n41438 = ~n23622 & ~n41437 ;
  assign n41439 = n41436 & ~n41438 ;
  assign n41440 = ~\pi0193  & n23548 ;
  assign n41441 = \pi0739  & ~n41440 ;
  assign n41442 = ~\pi0039  & \pi0739  ;
  assign n41443 = ~n22683 & n41442 ;
  assign n41444 = ~n41441 & ~n41443 ;
  assign n41445 = ~\pi0038  & n41444 ;
  assign n41446 = ~\pi0038  & \pi0193  ;
  assign n41447 = ~n26538 & n41446 ;
  assign n41448 = ~n41445 & ~n41447 ;
  assign n41449 = ~\pi0193  & ~n23567 ;
  assign n41450 = n23565 & n41449 ;
  assign n41451 = ~\pi0739  & n23575 ;
  assign n41452 = n23572 & n41451 ;
  assign n41453 = ~n41430 & ~n41452 ;
  assign n41454 = ~n41450 & ~n41453 ;
  assign n41455 = ~n41448 & ~n41454 ;
  assign n41456 = n6861 & n41455 ;
  assign n41457 = \pi0193  & \pi0603  ;
  assign n41458 = ~n20783 & n41457 ;
  assign n41459 = n41233 & n41458 ;
  assign n41460 = \pi0193  & \pi0680  ;
  assign n41461 = ~n20854 & n41460 ;
  assign n41462 = ~n20784 & n41461 ;
  assign n41463 = n1689 & n41462 ;
  assign n41464 = ~n41459 & ~n41463 ;
  assign n41465 = n26554 & ~n41464 ;
  assign n41466 = n1358 & n41465 ;
  assign n41467 = \pi0038  & ~n41466 ;
  assign n41468 = \pi0690  & ~n41467 ;
  assign n41469 = \pi0739  & ~n22317 ;
  assign n41470 = ~n31169 & ~n41469 ;
  assign n41471 = ~\pi0039  & n41470 ;
  assign n41472 = n21289 & n41471 ;
  assign n41473 = ~\pi0193  & \pi0690  ;
  assign n41474 = ~n41472 & n41473 ;
  assign n41475 = ~n41468 & ~n41474 ;
  assign n41476 = n6861 & n41475 ;
  assign n41477 = ~n41438 & ~n41476 ;
  assign n41478 = ~n41456 & n41477 ;
  assign n41479 = ~n41439 & ~n41478 ;
  assign n41480 = \pi0609  & ~n41479 ;
  assign n41481 = ~\pi0193  & ~\pi0625  ;
  assign n41482 = ~n22734 & ~n41481 ;
  assign n41483 = n41436 & ~n41482 ;
  assign n41484 = ~n41476 & ~n41482 ;
  assign n41485 = ~n41456 & n41484 ;
  assign n41486 = ~n41483 & ~n41485 ;
  assign n41487 = n6861 & ~n41435 ;
  assign n41488 = ~\pi0193  & \pi0625  ;
  assign n41489 = ~n22727 & ~n41488 ;
  assign n41490 = ~n41487 & ~n41489 ;
  assign n41491 = ~\pi1153  & ~n41490 ;
  assign n41492 = n41486 & n41491 ;
  assign n41493 = ~\pi0074  & \pi0690  ;
  assign n41494 = ~\pi0100  & n41493 ;
  assign n41495 = n1287 & n41494 ;
  assign n41496 = ~\pi0193  & ~n41495 ;
  assign n41497 = n21768 & n41496 ;
  assign n41498 = n21770 & n41496 ;
  assign n41499 = ~n21734 & n41498 ;
  assign n41500 = ~n41497 & ~n41499 ;
  assign n41501 = \pi0625  & ~n41500 ;
  assign n41502 = ~\pi0193  & ~n22017 ;
  assign n41503 = ~n21994 & n41502 ;
  assign n41504 = ~\pi0038  & ~\pi0193  ;
  assign n41505 = n6861 & ~n41504 ;
  assign n41506 = ~n22109 & n41505 ;
  assign n41507 = ~n41503 & ~n41506 ;
  assign n41508 = ~\pi0193  & ~n21757 ;
  assign n41509 = n22117 & ~n41508 ;
  assign n41510 = \pi0690  & ~n41509 ;
  assign n41511 = \pi0625  & n41510 ;
  assign n41512 = ~n41507 & n41511 ;
  assign n41513 = ~n41501 & ~n41512 ;
  assign n41514 = n21768 & n41481 ;
  assign n41515 = n21770 & n41481 ;
  assign n41516 = ~n21734 & n41515 ;
  assign n41517 = ~n41514 & ~n41516 ;
  assign n41518 = \pi1153  & n41517 ;
  assign n41519 = n41513 & n41518 ;
  assign n41520 = ~\pi0608  & ~n41519 ;
  assign n41521 = ~n41492 & n41520 ;
  assign n41522 = n41436 & ~n41489 ;
  assign n41523 = ~n41476 & ~n41489 ;
  assign n41524 = ~n41456 & n41523 ;
  assign n41525 = ~n41522 & ~n41524 ;
  assign n41526 = \pi1153  & n41482 ;
  assign n41527 = n23606 & ~n41435 ;
  assign n41528 = ~n41526 & ~n41527 ;
  assign n41529 = n41525 & ~n41528 ;
  assign n41530 = ~\pi0625  & ~n41500 ;
  assign n41531 = ~\pi0625  & n41510 ;
  assign n41532 = ~n41507 & n41531 ;
  assign n41533 = ~n41530 & ~n41532 ;
  assign n41534 = n21768 & n41488 ;
  assign n41535 = n21770 & n41488 ;
  assign n41536 = ~n21734 & n41535 ;
  assign n41537 = ~n41534 & ~n41536 ;
  assign n41538 = ~\pi1153  & n41537 ;
  assign n41539 = n41533 & n41538 ;
  assign n41540 = \pi0608  & ~n41539 ;
  assign n41541 = ~n41529 & n41540 ;
  assign n41542 = ~n41521 & ~n41541 ;
  assign n41543 = n23638 & ~n41542 ;
  assign n41544 = ~n41480 & ~n41543 ;
  assign n41545 = \pi0193  & ~n6861 ;
  assign n41546 = ~n20985 & n41545 ;
  assign n41547 = n21774 & n41546 ;
  assign n41548 = n26646 & ~n41435 ;
  assign n41549 = ~n41547 & ~n41548 ;
  assign n41550 = ~\pi0193  & n21768 ;
  assign n41551 = ~\pi0193  & n21770 ;
  assign n41552 = ~n21734 & n41551 ;
  assign n41553 = ~n41550 & ~n41552 ;
  assign n41554 = n26653 & n41553 ;
  assign n41555 = ~\pi0660  & ~n41554 ;
  assign n41556 = n41549 & n41555 ;
  assign n41557 = ~n41507 & n41510 ;
  assign n41558 = ~\pi0778  & n41500 ;
  assign n41559 = ~n41557 & n41558 ;
  assign n41560 = ~\pi0609  & ~n41559 ;
  assign n41561 = \pi1155  & ~n41560 ;
  assign n41562 = ~n41519 & ~n41539 ;
  assign n41563 = n22722 & ~n41562 ;
  assign n41564 = ~n41561 & ~n41563 ;
  assign n41565 = ~n41556 & ~n41564 ;
  assign n41566 = n41544 & n41565 ;
  assign n41567 = \pi0778  & ~n41542 ;
  assign n41568 = \pi0778  & ~n41562 ;
  assign n41569 = \pi0609  & ~n41559 ;
  assign n41570 = ~n41568 & n41569 ;
  assign n41571 = ~\pi1155  & n41546 ;
  assign n41572 = n26672 & ~n41435 ;
  assign n41573 = ~n41571 & ~n41572 ;
  assign n41574 = ~\pi0609  & ~n41573 ;
  assign n41575 = ~\pi1155  & ~n22767 ;
  assign n41576 = n41553 & n41575 ;
  assign n41577 = ~n22787 & ~n41576 ;
  assign n41578 = ~n41574 & n41577 ;
  assign n41579 = ~n41570 & ~n41578 ;
  assign n41580 = \pi0785  & ~n41579 ;
  assign n41581 = n41479 & ~n41580 ;
  assign n41582 = ~n41567 & n41581 ;
  assign n41583 = n20999 & n41546 ;
  assign n41584 = n26685 & ~n41435 ;
  assign n41585 = ~n41583 & ~n41584 ;
  assign n41586 = \pi0660  & ~n41576 ;
  assign n41587 = n41585 & n41586 ;
  assign n41588 = ~n41556 & ~n41587 ;
  assign n41589 = \pi0609  & ~n41577 ;
  assign n41590 = n41559 & n41589 ;
  assign n41591 = \pi0778  & n41589 ;
  assign n41592 = ~n41562 & n41591 ;
  assign n41593 = ~n41590 & ~n41592 ;
  assign n41594 = ~n41588 & n41593 ;
  assign n41595 = ~n41582 & n41594 ;
  assign n41596 = ~n41566 & n41595 ;
  assign n41597 = ~\pi0785  & ~n41582 ;
  assign n41598 = n26700 & ~n41597 ;
  assign n41599 = ~n41596 & n41598 ;
  assign n41600 = n26065 & ~n41562 ;
  assign n41601 = n26739 & n41500 ;
  assign n41602 = ~n41557 & n41601 ;
  assign n41603 = ~n23885 & n41553 ;
  assign n41604 = \pi0628  & ~n41603 ;
  assign n41605 = ~n41602 & n41604 ;
  assign n41606 = ~n41600 & n41605 ;
  assign n41607 = ~\pi0193  & ~\pi0628  ;
  assign n41608 = n21768 & n41607 ;
  assign n41609 = n21770 & n41607 ;
  assign n41610 = ~n21734 & n41609 ;
  assign n41611 = ~n41608 & ~n41610 ;
  assign n41612 = \pi1156  & n41611 ;
  assign n41613 = ~\pi0629  & n41612 ;
  assign n41614 = ~n41606 & n41613 ;
  assign n41615 = ~\pi0628  & ~n41603 ;
  assign n41616 = ~n41602 & n41615 ;
  assign n41617 = ~n41600 & n41616 ;
  assign n41618 = ~\pi0193  & \pi0628  ;
  assign n41619 = n21768 & n41618 ;
  assign n41620 = n21770 & n41618 ;
  assign n41621 = ~n21734 & n41620 ;
  assign n41622 = ~n41619 & ~n41621 ;
  assign n41623 = ~\pi1156  & n41622 ;
  assign n41624 = \pi0629  & n41623 ;
  assign n41625 = ~n41617 & n41624 ;
  assign n41626 = ~n41614 & ~n41625 ;
  assign n41627 = \pi0792  & ~n41626 ;
  assign n41628 = ~\pi0193  & ~n20811 ;
  assign n41629 = n21768 & n41628 ;
  assign n41630 = n21770 & n41628 ;
  assign n41631 = ~n21734 & n41630 ;
  assign n41632 = ~n41629 & ~n41631 ;
  assign n41633 = n23456 & ~n41435 ;
  assign n41634 = n21777 & n41545 ;
  assign n41635 = ~n21777 & n41553 ;
  assign n41636 = n20811 & ~n41635 ;
  assign n41637 = ~n41634 & n41636 ;
  assign n41638 = ~n41633 & n41637 ;
  assign n41639 = n41632 & ~n41638 ;
  assign n41640 = n23424 & ~n41639 ;
  assign n41641 = ~\pi0781  & ~n41635 ;
  assign n41642 = ~n23423 & ~n41634 ;
  assign n41643 = n41641 & n41642 ;
  assign n41644 = ~n41633 & n41643 ;
  assign n41645 = n23423 & ~n41553 ;
  assign n41646 = ~n41644 & ~n41645 ;
  assign n41647 = ~n41640 & n41646 ;
  assign n41648 = ~n23880 & ~n41647 ;
  assign n41649 = n23880 & ~n41553 ;
  assign n41650 = n24691 & ~n41649 ;
  assign n41651 = \pi0792  & n41650 ;
  assign n41652 = ~n41648 & n41651 ;
  assign n41653 = ~n41627 & ~n41652 ;
  assign n41654 = n22155 & n41632 ;
  assign n41655 = ~n41638 & n41654 ;
  assign n41656 = ~n22147 & ~n41559 ;
  assign n41657 = n22147 & ~n41553 ;
  assign n41658 = n39952 & ~n41657 ;
  assign n41659 = ~n41656 & n41658 ;
  assign n41660 = \pi0778  & n41658 ;
  assign n41661 = ~n41562 & n41660 ;
  assign n41662 = ~n41659 & ~n41661 ;
  assign n41663 = ~n41655 & n41662 ;
  assign n41664 = ~n21034 & ~n41663 ;
  assign n41665 = n23380 & ~n41559 ;
  assign n41666 = ~\pi0193  & ~n23380 ;
  assign n41667 = n21768 & n41666 ;
  assign n41668 = n21770 & n41666 ;
  assign n41669 = ~n21734 & n41668 ;
  assign n41670 = ~n41667 & ~n41669 ;
  assign n41671 = n21050 & n41670 ;
  assign n41672 = ~n41665 & n41671 ;
  assign n41673 = \pi0778  & n41671 ;
  assign n41674 = ~n41562 & n41673 ;
  assign n41675 = ~n41672 & ~n41674 ;
  assign n41676 = \pi0789  & ~n41675 ;
  assign n41677 = n23683 & ~n41639 ;
  assign n41678 = n21032 & ~n41634 ;
  assign n41679 = n41641 & n41678 ;
  assign n41680 = ~n41633 & n41679 ;
  assign n41681 = ~n21032 & ~n41553 ;
  assign n41682 = ~n20876 & ~n41681 ;
  assign n41683 = ~n41680 & n41682 ;
  assign n41684 = \pi0789  & n41683 ;
  assign n41685 = ~n41677 & n41684 ;
  assign n41686 = ~n41676 & ~n41685 ;
  assign n41687 = ~n21038 & n41686 ;
  assign n41688 = ~n41664 & n41687 ;
  assign n41689 = n41653 & n41688 ;
  assign n41690 = ~n41599 & n41689 ;
  assign n41691 = ~n22160 & n41670 ;
  assign n41692 = ~n41665 & n41691 ;
  assign n41693 = \pi0778  & n41691 ;
  assign n41694 = ~n41562 & n41693 ;
  assign n41695 = ~n41692 & ~n41694 ;
  assign n41696 = n22160 & n41553 ;
  assign n41697 = n20951 & ~n41696 ;
  assign n41698 = n41695 & n41697 ;
  assign n41699 = ~\pi0626  & ~n41645 ;
  assign n41700 = ~n41644 & n41699 ;
  assign n41701 = ~n41640 & n41700 ;
  assign n41702 = \pi0626  & n41553 ;
  assign n41703 = n20882 & ~n41702 ;
  assign n41704 = ~n41701 & n41703 ;
  assign n41705 = ~n41698 & ~n41704 ;
  assign n41706 = \pi0626  & ~n41645 ;
  assign n41707 = ~n41644 & n41706 ;
  assign n41708 = ~n41640 & n41707 ;
  assign n41709 = ~\pi0626  & n41553 ;
  assign n41710 = n20881 & ~n41709 ;
  assign n41711 = ~n41708 & n41710 ;
  assign n41712 = ~n23856 & ~n41711 ;
  assign n41713 = n41705 & n41712 ;
  assign n41714 = n41653 & ~n41713 ;
  assign n41715 = ~n26803 & n41714 ;
  assign n41716 = ~n21067 & ~n41715 ;
  assign n41717 = ~n41690 & n41716 ;
  assign n41718 = ~\pi0193  & ~n31367 ;
  assign n41719 = n21768 & n41718 ;
  assign n41720 = n21770 & n41718 ;
  assign n41721 = ~n21734 & n41720 ;
  assign n41722 = ~n41719 & ~n41721 ;
  assign n41723 = ~\pi0715  & n41722 ;
  assign n41724 = ~n23958 & ~n41723 ;
  assign n41725 = n31382 & ~n41647 ;
  assign n41726 = ~n41724 & ~n41725 ;
  assign n41727 = n26824 & ~n41726 ;
  assign n41728 = ~\pi0644  & ~n41722 ;
  assign n41729 = n34208 & ~n41647 ;
  assign n41730 = ~n41728 & ~n41729 ;
  assign n41731 = ~\pi0193  & \pi0644  ;
  assign n41732 = n21768 & n41731 ;
  assign n41733 = n21770 & n41731 ;
  assign n41734 = ~n21734 & n41733 ;
  assign n41735 = ~n41732 & ~n41734 ;
  assign n41736 = \pi0715  & n41735 ;
  assign n41737 = \pi0790  & n41736 ;
  assign n41738 = n41730 & n41737 ;
  assign n41739 = ~n35417 & ~n41738 ;
  assign n41740 = ~n41727 & ~n41739 ;
  assign n41741 = ~n41602 & ~n41603 ;
  assign n41742 = ~n41600 & n41741 ;
  assign n41743 = ~\pi0792  & ~n41742 ;
  assign n41744 = \pi0647  & ~n41743 ;
  assign n41745 = n21768 & n41281 ;
  assign n41746 = n21770 & n41281 ;
  assign n41747 = ~n21734 & n41746 ;
  assign n41748 = ~n41745 & ~n41747 ;
  assign n41749 = \pi1157  & n41748 ;
  assign n41750 = ~n41744 & n41749 ;
  assign n41751 = ~n41606 & n41612 ;
  assign n41752 = ~n41617 & n41623 ;
  assign n41753 = ~n41751 & ~n41752 ;
  assign n41754 = \pi0792  & n41749 ;
  assign n41755 = ~n41753 & n41754 ;
  assign n41756 = ~n41750 & ~n41755 ;
  assign n41757 = ~\pi0630  & ~n41756 ;
  assign n41758 = ~\pi0647  & ~n41743 ;
  assign n41759 = n21768 & n41286 ;
  assign n41760 = n21770 & n41286 ;
  assign n41761 = ~n21734 & n41760 ;
  assign n41762 = ~n41759 & ~n41761 ;
  assign n41763 = ~\pi1157  & n41762 ;
  assign n41764 = ~n41758 & n41763 ;
  assign n41765 = \pi0792  & n41763 ;
  assign n41766 = ~n41753 & n41765 ;
  assign n41767 = ~n41764 & ~n41766 ;
  assign n41768 = \pi0630  & ~n41767 ;
  assign n41769 = ~n20846 & n41649 ;
  assign n41770 = n30376 & ~n41647 ;
  assign n41771 = ~n41769 & ~n41770 ;
  assign n41772 = n20846 & ~n41553 ;
  assign n41773 = ~n20910 & ~n41772 ;
  assign n41774 = n41771 & n41773 ;
  assign n41775 = ~n41768 & ~n41774 ;
  assign n41776 = ~n41757 & n41775 ;
  assign n41777 = \pi0787  & ~n41776 ;
  assign n41778 = ~n41740 & ~n41777 ;
  assign n41779 = ~n41717 & n41778 ;
  assign n41780 = ~\pi0787  & n41743 ;
  assign n41781 = n33084 & ~n41753 ;
  assign n41782 = ~n41780 & ~n41781 ;
  assign n41783 = ~\pi0644  & n41782 ;
  assign n41784 = \pi0715  & ~n41783 ;
  assign n41785 = n41756 & n41767 ;
  assign n41786 = n26918 & ~n41785 ;
  assign n41787 = ~n41784 & ~n41786 ;
  assign n41788 = ~\pi0193  & ~\pi0644  ;
  assign n41789 = n21768 & n41788 ;
  assign n41790 = n21770 & n41788 ;
  assign n41791 = ~n21734 & n41790 ;
  assign n41792 = ~n41789 & ~n41791 ;
  assign n41793 = n41726 & n41792 ;
  assign n41794 = \pi1160  & ~n41793 ;
  assign n41795 = n41787 & n41794 ;
  assign n41796 = \pi0644  & n41782 ;
  assign n41797 = ~\pi0715  & ~n41796 ;
  assign n41798 = n33098 & ~n41785 ;
  assign n41799 = ~n41797 & ~n41798 ;
  assign n41800 = n41730 & n41736 ;
  assign n41801 = ~\pi1160  & ~n41800 ;
  assign n41802 = n41799 & n41801 ;
  assign n41803 = ~n41795 & ~n41802 ;
  assign n41804 = \pi0790  & ~n41803 ;
  assign n41805 = ~n41411 & ~n41804 ;
  assign n41806 = ~n41779 & n41805 ;
  assign n41807 = ~n41413 & ~n41806 ;
  assign n41808 = \pi0194  & ~\pi0832  ;
  assign n41809 = ~n21132 & ~n41808 ;
  assign n41810 = ~\pi0194  & ~n1689 ;
  assign n41811 = ~n21032 & ~n41810 ;
  assign n41812 = \pi0789  & n41811 ;
  assign n41813 = n23423 & ~n41812 ;
  assign n41814 = \pi0748  & n1689 ;
  assign n41815 = n20784 & n41814 ;
  assign n41816 = ~n41810 & ~n41815 ;
  assign n41817 = n20794 & ~n41816 ;
  assign n41818 = n20796 & ~n41817 ;
  assign n41819 = n20799 & ~n41816 ;
  assign n41820 = n20801 & ~n41819 ;
  assign n41821 = ~n41818 & ~n41820 ;
  assign n41822 = ~\pi0785  & ~n41810 ;
  assign n41823 = ~n41815 & n41822 ;
  assign n41824 = ~n20804 & ~n41823 ;
  assign n41825 = ~n20812 & n41824 ;
  assign n41826 = ~n41812 & n41825 ;
  assign n41827 = n41821 & n41826 ;
  assign n41828 = ~n41813 & ~n41827 ;
  assign n41829 = ~\pi0626  & n41828 ;
  assign n41830 = \pi0626  & ~n41810 ;
  assign n41831 = n20882 & ~n41830 ;
  assign n41832 = ~n41829 & n41831 ;
  assign n41833 = \pi0730  & n1689 ;
  assign n41834 = n20855 & n41833 ;
  assign n41835 = ~n20861 & n41834 ;
  assign n41836 = ~n41810 & ~n41835 ;
  assign n41837 = n23170 & ~n41836 ;
  assign n41838 = ~\pi0626  & ~n41810 ;
  assign n41839 = n20881 & ~n41838 ;
  assign n41840 = ~n41837 & ~n41839 ;
  assign n41841 = \pi0626  & ~n41837 ;
  assign n41842 = n41828 & n41841 ;
  assign n41843 = ~n41840 & ~n41842 ;
  assign n41844 = ~n41832 & ~n41843 ;
  assign n41845 = \pi0788  & ~n41844 ;
  assign n41846 = \pi0680  & \pi0730  ;
  assign n41847 = ~n20854 & n41846 ;
  assign n41848 = ~n20861 & n41847 ;
  assign n41849 = ~n20986 & n41848 ;
  assign n41850 = \pi0603  & \pi0748  ;
  assign n41851 = ~n20783 & n41850 ;
  assign n41852 = ~n20985 & n41851 ;
  assign n41853 = ~n41810 & ~n41852 ;
  assign n41854 = ~n41849 & n41853 ;
  assign n41855 = \pi0194  & ~n1689 ;
  assign n41856 = ~\pi0609  & ~n41855 ;
  assign n41857 = ~n41854 & n41856 ;
  assign n41858 = ~\pi1155  & ~n41810 ;
  assign n41859 = ~n41835 & n41858 ;
  assign n41860 = ~n20999 & ~n41859 ;
  assign n41861 = ~n41857 & ~n41860 ;
  assign n41862 = \pi1155  & ~n41819 ;
  assign n41863 = ~\pi0660  & ~n41862 ;
  assign n41864 = ~n41861 & n41863 ;
  assign n41865 = ~n21007 & ~n41818 ;
  assign n41866 = \pi0609  & ~n41855 ;
  assign n41867 = ~n41854 & n41866 ;
  assign n41868 = \pi1155  & ~n41810 ;
  assign n41869 = ~n41835 & n41868 ;
  assign n41870 = ~n21774 & ~n41869 ;
  assign n41871 = \pi0785  & ~n41870 ;
  assign n41872 = ~n41867 & n41871 ;
  assign n41873 = n41865 & ~n41872 ;
  assign n41874 = ~n41864 & ~n41873 ;
  assign n41875 = ~n41854 & ~n41855 ;
  assign n41876 = ~\pi0785  & ~n41875 ;
  assign n41877 = n21022 & ~n41876 ;
  assign n41878 = ~n41874 & n41877 ;
  assign n41879 = n20964 & n41824 ;
  assign n41880 = n41821 & n41879 ;
  assign n41881 = \pi0627  & ~n41810 ;
  assign n41882 = ~n41835 & n41881 ;
  assign n41883 = ~n20968 & ~n41882 ;
  assign n41884 = ~n41880 & ~n41883 ;
  assign n41885 = n20974 & n41824 ;
  assign n41886 = n41821 & n41885 ;
  assign n41887 = ~\pi0627  & ~n41810 ;
  assign n41888 = ~n41835 & n41887 ;
  assign n41889 = ~n20978 & ~n41888 ;
  assign n41890 = ~n41886 & ~n41889 ;
  assign n41891 = ~n41884 & ~n41890 ;
  assign n41892 = \pi0781  & n41891 ;
  assign n41893 = ~n21034 & ~n41892 ;
  assign n41894 = ~n41878 & n41893 ;
  assign n41895 = ~n20876 & n41811 ;
  assign n41896 = ~n24969 & ~n41895 ;
  assign n41897 = n41825 & ~n41895 ;
  assign n41898 = n41821 & n41897 ;
  assign n41899 = ~n41896 & ~n41898 ;
  assign n41900 = n21050 & ~n41810 ;
  assign n41901 = ~n41835 & n41900 ;
  assign n41902 = ~n21051 & ~n41901 ;
  assign n41903 = ~n21038 & n41902 ;
  assign n41904 = ~n41899 & n41903 ;
  assign n41905 = ~n23177 & ~n41904 ;
  assign n41906 = ~n41894 & ~n41905 ;
  assign n41907 = ~n41845 & ~n41906 ;
  assign n41908 = ~n23880 & ~n41812 ;
  assign n41909 = n23423 & n41908 ;
  assign n41910 = n41825 & n41908 ;
  assign n41911 = n41821 & n41910 ;
  assign n41912 = ~n41909 & ~n41911 ;
  assign n41913 = ~\pi0194  & \pi0792  ;
  assign n41914 = ~n1689 & n41913 ;
  assign n41915 = ~n20845 & n41914 ;
  assign n41916 = ~n20910 & ~n41915 ;
  assign n41917 = ~\pi0194  & \pi0788  ;
  assign n41918 = ~n1689 & n41917 ;
  assign n41919 = ~n20778 & n41918 ;
  assign n41920 = n41916 & ~n41919 ;
  assign n41921 = n41912 & n41920 ;
  assign n41922 = n20846 & n41916 ;
  assign n41923 = n20879 & ~n41836 ;
  assign n41924 = n20895 & n41923 ;
  assign n41925 = ~\pi0194  & \pi0647  ;
  assign n41926 = ~n1689 & n41925 ;
  assign n41927 = n20897 & ~n41926 ;
  assign n41928 = ~n41924 & n41927 ;
  assign n41929 = ~\pi0194  & ~\pi0647  ;
  assign n41930 = ~n1689 & n41929 ;
  assign n41931 = n20849 & ~n41930 ;
  assign n41932 = ~n24761 & ~n41931 ;
  assign n41933 = ~n24761 & n39577 ;
  assign n41934 = n41923 & n41933 ;
  assign n41935 = ~n41932 & ~n41934 ;
  assign n41936 = ~n41928 & ~n41935 ;
  assign n41937 = ~n41922 & n41936 ;
  assign n41938 = ~n41921 & n41937 ;
  assign n41939 = ~n29722 & ~n41938 ;
  assign n41940 = ~n23856 & ~n41939 ;
  assign n41941 = ~n41907 & n41940 ;
  assign n41942 = n39577 & n41923 ;
  assign n41943 = \pi1157  & ~n41930 ;
  assign n41944 = ~n41942 & n41943 ;
  assign n41945 = ~\pi1157  & ~n41926 ;
  assign n41946 = ~n41924 & n41945 ;
  assign n41947 = ~n41944 & ~n41946 ;
  assign n41948 = \pi0787  & ~n41947 ;
  assign n41949 = n24844 & n41923 ;
  assign n41950 = ~n24843 & ~n41949 ;
  assign n41951 = ~n41948 & ~n41950 ;
  assign n41952 = n41912 & ~n41919 ;
  assign n41953 = n31580 & ~n41952 ;
  assign n41954 = ~n41951 & ~n41953 ;
  assign n41955 = n23313 & ~n41954 ;
  assign n41956 = \pi0790  & n41955 ;
  assign n41957 = n31588 & ~n41952 ;
  assign n41958 = ~n23414 & n41810 ;
  assign n41959 = ~n24886 & n41958 ;
  assign n41960 = n20891 & n41923 ;
  assign n41961 = ~\pi0787  & ~n41960 ;
  assign n41962 = ~\pi1160  & ~n41961 ;
  assign n41963 = ~n41948 & n41962 ;
  assign n41964 = ~n41959 & ~n41963 ;
  assign n41965 = ~n41957 & n41964 ;
  assign n41966 = ~n23312 & ~n41959 ;
  assign n41967 = \pi0790  & ~n41966 ;
  assign n41968 = ~n41965 & n41967 ;
  assign n41969 = ~n41956 & ~n41968 ;
  assign n41970 = n20938 & n41923 ;
  assign n41971 = \pi0629  & ~n41919 ;
  assign n41972 = ~n41970 & n41971 ;
  assign n41973 = n41912 & n41972 ;
  assign n41974 = n21077 & n41923 ;
  assign n41975 = ~\pi0629  & ~n41919 ;
  assign n41976 = ~n41974 & n41975 ;
  assign n41977 = n41912 & n41976 ;
  assign n41978 = n29714 & ~n41970 ;
  assign n41979 = n29709 & ~n41974 ;
  assign n41980 = \pi0792  & ~n41979 ;
  assign n41981 = ~n41978 & n41980 ;
  assign n41982 = ~n41977 & n41981 ;
  assign n41983 = ~n41973 & n41982 ;
  assign n41984 = ~n21067 & ~n41983 ;
  assign n41985 = ~n41939 & ~n41984 ;
  assign n41986 = \pi0832  & ~n41985 ;
  assign n41987 = n41969 & n41986 ;
  assign n41988 = ~n41941 & n41987 ;
  assign n41989 = n41809 & ~n41988 ;
  assign n41990 = \pi0194  & ~n25040 ;
  assign n41991 = ~n25024 & n41990 ;
  assign n41992 = \pi0748  & n41991 ;
  assign n41993 = ~\pi0194  & ~n25033 ;
  assign n41994 = \pi0748  & n41993 ;
  assign n41995 = ~n25028 & n41994 ;
  assign n41996 = ~n41992 & ~n41995 ;
  assign n41997 = n6861 & ~n41996 ;
  assign n41998 = \pi0194  & ~n6861 ;
  assign n41999 = ~\pi0194  & n21770 ;
  assign n42000 = ~n21734 & n41999 ;
  assign n42001 = ~\pi0194  & n22124 ;
  assign n42002 = ~n42000 & ~n42001 ;
  assign n42003 = ~\pi0748  & n1289 ;
  assign n42004 = n1287 & n42003 ;
  assign n42005 = n42002 & n42004 ;
  assign n42006 = ~n41998 & ~n42005 ;
  assign n42007 = ~n41997 & n42006 ;
  assign n42008 = n21777 & ~n42007 ;
  assign n42009 = ~\pi0194  & n21768 ;
  assign n42010 = ~n42000 & ~n42009 ;
  assign n42011 = ~n21777 & n42010 ;
  assign n42012 = ~\pi0781  & ~n42011 ;
  assign n42013 = ~n42008 & n42012 ;
  assign n42014 = \pi0619  & n42013 ;
  assign n42015 = ~\pi0618  & ~n42011 ;
  assign n42016 = ~\pi0194  & \pi0618  ;
  assign n42017 = n21768 & n42016 ;
  assign n42018 = n21770 & n42016 ;
  assign n42019 = ~n21734 & n42018 ;
  assign n42020 = ~n42017 & ~n42019 ;
  assign n42021 = ~\pi1154  & n42020 ;
  assign n42022 = ~n42015 & n42021 ;
  assign n42023 = n21777 & n42021 ;
  assign n42024 = ~n42007 & n42023 ;
  assign n42025 = ~n42022 & ~n42024 ;
  assign n42026 = \pi0781  & n42025 ;
  assign n42027 = \pi0618  & ~n42011 ;
  assign n42028 = ~\pi0194  & ~\pi0618  ;
  assign n42029 = n21768 & n42028 ;
  assign n42030 = n21770 & n42028 ;
  assign n42031 = ~n21734 & n42030 ;
  assign n42032 = ~n42029 & ~n42031 ;
  assign n42033 = \pi1154  & n42032 ;
  assign n42034 = ~n42027 & n42033 ;
  assign n42035 = n21777 & n42033 ;
  assign n42036 = ~n42007 & n42035 ;
  assign n42037 = ~n42034 & ~n42036 ;
  assign n42038 = \pi0619  & n42037 ;
  assign n42039 = n42026 & n42038 ;
  assign n42040 = ~n42014 & ~n42039 ;
  assign n42041 = ~\pi0194  & ~\pi0619  ;
  assign n42042 = n21768 & n42041 ;
  assign n42043 = n21770 & n42041 ;
  assign n42044 = ~n21734 & n42043 ;
  assign n42045 = ~n42042 & ~n42044 ;
  assign n42046 = \pi1159  & n42045 ;
  assign n42047 = n42040 & n42046 ;
  assign n42048 = ~\pi0619  & n42013 ;
  assign n42049 = ~\pi0619  & n42037 ;
  assign n42050 = n42026 & n42049 ;
  assign n42051 = ~n42048 & ~n42050 ;
  assign n42052 = ~\pi0194  & \pi0619  ;
  assign n42053 = n21768 & n42052 ;
  assign n42054 = n21770 & n42052 ;
  assign n42055 = ~n21734 & n42054 ;
  assign n42056 = ~n42053 & ~n42055 ;
  assign n42057 = ~\pi1159  & n42056 ;
  assign n42058 = n42051 & n42057 ;
  assign n42059 = ~n42047 & ~n42058 ;
  assign n42060 = n39235 & n42059 ;
  assign n42061 = ~\pi0789  & n42012 ;
  assign n42062 = ~n42008 & n42061 ;
  assign n42063 = ~\pi0789  & n42037 ;
  assign n42064 = n42026 & n42063 ;
  assign n42065 = ~n42062 & ~n42064 ;
  assign n42066 = ~n23880 & ~n42065 ;
  assign n42067 = n23880 & ~n42010 ;
  assign n42068 = n21092 & ~n42067 ;
  assign n42069 = ~n42066 & n42068 ;
  assign n42070 = ~n42060 & n42069 ;
  assign n42071 = ~n21092 & n42010 ;
  assign n42072 = \pi0644  & ~n42071 ;
  assign n42073 = ~n42070 & n42072 ;
  assign n42074 = ~\pi0194  & ~\pi0644  ;
  assign n42075 = n21768 & n42074 ;
  assign n42076 = n21770 & n42074 ;
  assign n42077 = ~n21734 & n42076 ;
  assign n42078 = ~n42075 & ~n42077 ;
  assign n42079 = n23412 & n42078 ;
  assign n42080 = ~n42073 & n42079 ;
  assign n42081 = ~\pi0194  & \pi0644  ;
  assign n42082 = n21768 & n42081 ;
  assign n42083 = n21770 & n42081 ;
  assign n42084 = ~n21734 & n42083 ;
  assign n42085 = ~n42082 & ~n42084 ;
  assign n42086 = n23413 & n42085 ;
  assign n42087 = ~n22849 & n42010 ;
  assign n42088 = n33294 & n42087 ;
  assign n42089 = ~\pi0730  & n6861 ;
  assign n42090 = n42002 & n42089 ;
  assign n42091 = ~\pi0194  & ~n25669 ;
  assign n42092 = ~n31625 & n42091 ;
  assign n42093 = \pi0730  & n6861 ;
  assign n42094 = n42092 & n42093 ;
  assign n42095 = ~n42090 & ~n42094 ;
  assign n42096 = \pi0194  & ~n31632 ;
  assign n42097 = \pi0625  & ~n42096 ;
  assign n42098 = n42095 & n42097 ;
  assign n42099 = ~\pi0194  & ~\pi0625  ;
  assign n42100 = n21768 & n42099 ;
  assign n42101 = n21770 & n42099 ;
  assign n42102 = ~n21734 & n42101 ;
  assign n42103 = ~n42100 & ~n42102 ;
  assign n42104 = \pi1153  & n42103 ;
  assign n42105 = ~n42098 & n42104 ;
  assign n42106 = ~\pi0625  & ~n42096 ;
  assign n42107 = n42095 & n42106 ;
  assign n42108 = ~\pi0194  & \pi0625  ;
  assign n42109 = n21768 & n42108 ;
  assign n42110 = n21770 & n42108 ;
  assign n42111 = ~n21734 & n42110 ;
  assign n42112 = ~n42109 & ~n42111 ;
  assign n42113 = ~\pi1153  & n42112 ;
  assign n42114 = ~n42107 & n42113 ;
  assign n42115 = ~n42105 & ~n42114 ;
  assign n42116 = n22148 & ~n42115 ;
  assign n42117 = n42095 & ~n42096 ;
  assign n42118 = n22151 & ~n42117 ;
  assign n42119 = n22147 & n42010 ;
  assign n42120 = ~n42118 & ~n42119 ;
  assign n42121 = ~n42116 & n42120 ;
  assign n42122 = n33343 & ~n42121 ;
  assign n42123 = ~n42088 & ~n42122 ;
  assign n42124 = ~n33294 & n42010 ;
  assign n42125 = ~n23942 & ~n42124 ;
  assign n42126 = n42123 & n42125 ;
  assign n42127 = n23942 & ~n42010 ;
  assign n42128 = n23518 & ~n42127 ;
  assign n42129 = ~n42126 & n42128 ;
  assign n42130 = ~n42086 & ~n42129 ;
  assign n42131 = ~\pi0644  & ~n42071 ;
  assign n42132 = ~n42129 & n42131 ;
  assign n42133 = ~n42070 & n42132 ;
  assign n42134 = ~n42130 & ~n42133 ;
  assign n42135 = ~n42080 & ~n42134 ;
  assign n42136 = \pi0790  & ~n42135 ;
  assign n42137 = n24761 & ~n42136 ;
  assign n42138 = n24691 & ~n42067 ;
  assign n42139 = ~n42066 & n42138 ;
  assign n42140 = ~n42060 & n42139 ;
  assign n42141 = ~n22155 & ~n42119 ;
  assign n42142 = ~n42118 & n42141 ;
  assign n42143 = ~n42116 & n42142 ;
  assign n42144 = n22155 & ~n42010 ;
  assign n42145 = n22162 & ~n42144 ;
  assign n42146 = ~n42143 & n42145 ;
  assign n42147 = ~n22162 & n42010 ;
  assign n42148 = \pi0628  & ~n42147 ;
  assign n42149 = ~n42146 & n42148 ;
  assign n42150 = ~\pi0194  & ~\pi0628  ;
  assign n42151 = n21768 & n42150 ;
  assign n42152 = n21770 & n42150 ;
  assign n42153 = ~n21734 & n42152 ;
  assign n42154 = ~n42151 & ~n42153 ;
  assign n42155 = n20843 & n42154 ;
  assign n42156 = ~n42149 & n42155 ;
  assign n42157 = ~\pi0628  & ~n42147 ;
  assign n42158 = ~n42146 & n42157 ;
  assign n42159 = ~\pi0194  & \pi0628  ;
  assign n42160 = n21768 & n42159 ;
  assign n42161 = n21770 & n42159 ;
  assign n42162 = ~n21734 & n42161 ;
  assign n42163 = ~n42160 & ~n42162 ;
  assign n42164 = n20844 & n42163 ;
  assign n42165 = ~n42158 & n42164 ;
  assign n42166 = ~n42156 & ~n42165 ;
  assign n42167 = ~n42140 & n42166 ;
  assign n42168 = n24724 & ~n42167 ;
  assign n42169 = \pi1159  & ~n42144 ;
  assign n42170 = ~n42143 & n42169 ;
  assign n42171 = n37561 & ~n42170 ;
  assign n42172 = ~n42058 & n42171 ;
  assign n42173 = ~\pi1159  & ~n42144 ;
  assign n42174 = ~n42143 & n42173 ;
  assign n42175 = n37566 & ~n42174 ;
  assign n42176 = ~n42047 & n42175 ;
  assign n42177 = ~n42172 & ~n42176 ;
  assign n42178 = \pi0789  & ~n42177 ;
  assign n42179 = ~\pi0618  & ~n42119 ;
  assign n42180 = ~n42118 & n42179 ;
  assign n42181 = ~n42116 & n42180 ;
  assign n42182 = \pi1154  & ~n42181 ;
  assign n42183 = \pi0627  & n42025 ;
  assign n42184 = ~n42182 & n42183 ;
  assign n42185 = \pi0618  & ~n42119 ;
  assign n42186 = ~n42118 & n42185 ;
  assign n42187 = ~n42116 & n42186 ;
  assign n42188 = ~\pi1154  & ~n42187 ;
  assign n42189 = ~\pi0627  & n42037 ;
  assign n42190 = ~n42188 & n42189 ;
  assign n42191 = ~n42184 & ~n42190 ;
  assign n42192 = n32123 & ~n42046 ;
  assign n42193 = n31279 & n42056 ;
  assign n42194 = ~n33522 & ~n42193 ;
  assign n42195 = ~n42192 & ~n42194 ;
  assign n42196 = \pi0781  & ~n42195 ;
  assign n42197 = ~n42191 & n42196 ;
  assign n42198 = ~n42178 & ~n42197 ;
  assign n42199 = ~n21038 & ~n42198 ;
  assign n42200 = \pi0038  & \pi0194  ;
  assign n42201 = ~n22708 & n42200 ;
  assign n42202 = ~\pi0038  & \pi0194  ;
  assign n42203 = ~n42201 & ~n42202 ;
  assign n42204 = ~n23558 & ~n42201 ;
  assign n42205 = n23557 & n42204 ;
  assign n42206 = ~n42203 & ~n42205 ;
  assign n42207 = ~\pi0194  & n23548 ;
  assign n42208 = ~n25191 & n42207 ;
  assign n42209 = ~n25190 & n42208 ;
  assign n42210 = \pi0730  & \pi0748  ;
  assign n42211 = ~n42209 & n42210 ;
  assign n42212 = ~n42206 & n42211 ;
  assign n42213 = ~\pi0194  & ~n31749 ;
  assign n42214 = \pi0194  & ~n25217 ;
  assign n42215 = ~\pi0748  & ~n42214 ;
  assign n42216 = ~\pi0748  & n31753 ;
  assign n42217 = n23572 & n42216 ;
  assign n42218 = ~n42215 & ~n42217 ;
  assign n42219 = \pi0730  & ~n42218 ;
  assign n42220 = ~n42213 & n42219 ;
  assign n42221 = ~n42212 & ~n42220 ;
  assign n42222 = ~\pi0748  & n42002 ;
  assign n42223 = ~\pi0730  & n41996 ;
  assign n42224 = ~n42222 & n42223 ;
  assign n42225 = n6861 & ~n42224 ;
  assign n42226 = n42221 & n42225 ;
  assign n42227 = ~n22734 & ~n42099 ;
  assign n42228 = ~n42226 & ~n42227 ;
  assign n42229 = ~n22727 & ~n42108 ;
  assign n42230 = ~n42005 & ~n42229 ;
  assign n42231 = ~n41997 & n42230 ;
  assign n42232 = ~\pi1153  & ~n42231 ;
  assign n42233 = ~n42228 & n42232 ;
  assign n42234 = ~\pi0608  & ~n42105 ;
  assign n42235 = ~n42233 & n42234 ;
  assign n42236 = ~n42226 & ~n42229 ;
  assign n42237 = ~n42005 & ~n42227 ;
  assign n42238 = ~n41997 & n42237 ;
  assign n42239 = \pi1153  & ~n42238 ;
  assign n42240 = ~n42236 & n42239 ;
  assign n42241 = \pi0608  & ~n42114 ;
  assign n42242 = ~n42240 & n42241 ;
  assign n42243 = ~n42235 & ~n42242 ;
  assign n42244 = n23613 & ~n42243 ;
  assign n42245 = \pi0778  & ~n42115 ;
  assign n42246 = \pi0609  & ~n42096 ;
  assign n42247 = n42095 & n42246 ;
  assign n42248 = ~n23638 & ~n42247 ;
  assign n42249 = ~n42245 & ~n42248 ;
  assign n42250 = ~\pi0194  & ~\pi0778  ;
  assign n42251 = ~n23622 & ~n42250 ;
  assign n42252 = ~\pi0609  & ~n42251 ;
  assign n42253 = ~n42226 & n42252 ;
  assign n42254 = ~\pi1155  & ~n42253 ;
  assign n42255 = ~n42249 & n42254 ;
  assign n42256 = ~n42244 & n42255 ;
  assign n42257 = ~n22788 & n42010 ;
  assign n42258 = ~\pi0660  & ~n42257 ;
  assign n42259 = ~n22787 & ~n42258 ;
  assign n42260 = n37651 & ~n42007 ;
  assign n42261 = ~n42259 & ~n42260 ;
  assign n42262 = ~n42256 & n42261 ;
  assign n42263 = ~n22767 & n42010 ;
  assign n42264 = \pi0660  & ~n42263 ;
  assign n42265 = ~n22766 & ~n42264 ;
  assign n42266 = n31822 & ~n42007 ;
  assign n42267 = ~n42265 & ~n42266 ;
  assign n42268 = \pi0785  & ~n42267 ;
  assign n42269 = ~\pi0609  & ~n42096 ;
  assign n42270 = n42095 & n42269 ;
  assign n42271 = ~n23613 & ~n42270 ;
  assign n42272 = \pi1155  & n42271 ;
  assign n42273 = n22722 & ~n42115 ;
  assign n42274 = ~n42272 & ~n42273 ;
  assign n42275 = \pi0609  & ~n42251 ;
  assign n42276 = ~n42226 & n42275 ;
  assign n42277 = \pi0785  & ~n42276 ;
  assign n42278 = ~n42274 & n42277 ;
  assign n42279 = ~n42268 & ~n42278 ;
  assign n42280 = n23638 & ~n42268 ;
  assign n42281 = ~n42243 & n42280 ;
  assign n42282 = ~n42279 & ~n42281 ;
  assign n42283 = ~n42262 & n42282 ;
  assign n42284 = n21019 & ~n42021 ;
  assign n42285 = n21020 & n42032 ;
  assign n42286 = ~n33630 & ~n42285 ;
  assign n42287 = ~n42284 & ~n42286 ;
  assign n42288 = ~n42226 & ~n42251 ;
  assign n42289 = ~\pi0785  & ~n42288 ;
  assign n42290 = ~n42195 & ~n42289 ;
  assign n42291 = \pi0778  & ~n42195 ;
  assign n42292 = ~n42243 & n42291 ;
  assign n42293 = ~n42290 & ~n42292 ;
  assign n42294 = ~n42287 & ~n42293 ;
  assign n42295 = ~n21038 & n42294 ;
  assign n42296 = ~n42283 & n42295 ;
  assign n42297 = ~n42199 & ~n42296 ;
  assign n42298 = \pi0789  & n30606 ;
  assign n42299 = n42059 & n42298 ;
  assign n42300 = n30606 & ~n42065 ;
  assign n42301 = \pi0641  & n42087 ;
  assign n42302 = n33656 & ~n42121 ;
  assign n42303 = ~n42301 & ~n42302 ;
  assign n42304 = ~\pi0641  & n42010 ;
  assign n42305 = n20776 & ~n42304 ;
  assign n42306 = n42303 & n42305 ;
  assign n42307 = ~n42300 & ~n42306 ;
  assign n42308 = ~n42299 & n42307 ;
  assign n42309 = ~\pi0641  & n42087 ;
  assign n42310 = n33649 & ~n42121 ;
  assign n42311 = ~n42309 & ~n42310 ;
  assign n42312 = \pi0641  & n42010 ;
  assign n42313 = n20777 & ~n42312 ;
  assign n42314 = n42311 & n42313 ;
  assign n42315 = ~n23856 & ~n42314 ;
  assign n42316 = ~n21067 & n42315 ;
  assign n42317 = n42308 & n42316 ;
  assign n42318 = ~n38126 & ~n42317 ;
  assign n42319 = n42297 & ~n42318 ;
  assign n42320 = ~n42168 & ~n42319 ;
  assign n42321 = ~\pi0647  & ~n42124 ;
  assign n42322 = n42123 & n42321 ;
  assign n42323 = n21768 & n41925 ;
  assign n42324 = n21770 & n41925 ;
  assign n42325 = ~n21734 & n42324 ;
  assign n42326 = ~n42323 & ~n42325 ;
  assign n42327 = n20897 & n42326 ;
  assign n42328 = ~n42322 & n42327 ;
  assign n42329 = \pi0647  & ~n42124 ;
  assign n42330 = n42123 & n42329 ;
  assign n42331 = n21768 & n41929 ;
  assign n42332 = n21770 & n41929 ;
  assign n42333 = ~n21734 & n42332 ;
  assign n42334 = ~n42331 & ~n42333 ;
  assign n42335 = n20849 & n42334 ;
  assign n42336 = ~n42330 & n42335 ;
  assign n42337 = n20910 & ~n42336 ;
  assign n42338 = \pi0789  & ~n42047 ;
  assign n42339 = ~n42058 & n42338 ;
  assign n42340 = n30376 & n42065 ;
  assign n42341 = ~n42339 & n42340 ;
  assign n42342 = ~n30376 & n42010 ;
  assign n42343 = ~n42336 & ~n42342 ;
  assign n42344 = ~n42341 & n42343 ;
  assign n42345 = ~n42337 & ~n42344 ;
  assign n42346 = ~n42328 & ~n42345 ;
  assign n42347 = \pi0787  & ~n42346 ;
  assign n42348 = ~n42136 & ~n42347 ;
  assign n42349 = n42320 & n42348 ;
  assign n42350 = ~n42137 & ~n42349 ;
  assign n42351 = n9948 & ~n41988 ;
  assign n42352 = ~n42350 & n42351 ;
  assign n42353 = ~n41989 & ~n42352 ;
  assign n42354 = n20114 & ~n20641 ;
  assign n42355 = n20061 & ~n20739 ;
  assign n42356 = ~n42354 & ~n42355 ;
  assign n42357 = n7597 & ~n20062 ;
  assign n42358 = ~n20744 & ~n42357 ;
  assign n42359 = n13577 & ~n42358 ;
  assign n42360 = n6921 & n42359 ;
  assign n42361 = \pi0299  & ~n42360 ;
  assign n42362 = \pi0232  & ~n42361 ;
  assign n42363 = n42356 & n42362 ;
  assign n42364 = n20641 & n20642 ;
  assign n42365 = ~n20752 & ~n42364 ;
  assign n42366 = \pi0039  & n42365 ;
  assign n42367 = ~n42363 & n42366 ;
  assign n42368 = n13708 & ~n20064 ;
  assign n42369 = n10937 & n42368 ;
  assign n42370 = n10319 & n42369 ;
  assign n42371 = ~\pi0039  & ~n42370 ;
  assign n42372 = ~\pi0138  & ~\pi0196  ;
  assign n42373 = n20628 & n42372 ;
  assign n42374 = n16758 & n42373 ;
  assign n42375 = \pi0195  & ~n42374 ;
  assign n42376 = n13386 & ~n42375 ;
  assign n42377 = ~n42371 & n42376 ;
  assign n42378 = ~n42367 & n42377 ;
  assign n42379 = ~\pi0062  & n20532 ;
  assign n42380 = ~n6706 & n20061 ;
  assign n42381 = ~n11239 & n42380 ;
  assign n42382 = n6706 & n20061 ;
  assign n42383 = ~n10366 & n42382 ;
  assign n42384 = ~\pi0198  & n42382 ;
  assign n42385 = ~n10375 & n42384 ;
  assign n42386 = ~n42383 & ~n42385 ;
  assign n42387 = ~n42381 & n42386 ;
  assign n42388 = ~n10366 & n20091 ;
  assign n42389 = ~\pi0210  & n20091 ;
  assign n42390 = ~n10375 & n42389 ;
  assign n42391 = ~n42388 & ~n42390 ;
  assign n42392 = \pi0299  & ~n42391 ;
  assign n42393 = \pi0299  & ~n20091 ;
  assign n42394 = ~n10735 & n42393 ;
  assign n42395 = ~n42392 & ~n42394 ;
  assign n42396 = ~n11239 & n20114 ;
  assign n42397 = \pi0232  & ~n42396 ;
  assign n42398 = n42395 & n42397 ;
  assign n42399 = n42387 & n42398 ;
  assign n42400 = ~n20580 & ~n20582 ;
  assign n42401 = n11407 & n42400 ;
  assign n42402 = ~n42399 & n42401 ;
  assign n42403 = ~n10220 & n20061 ;
  assign n42404 = \pi0232  & n42403 ;
  assign n42405 = ~n20680 & n42404 ;
  assign n42406 = ~n6736 & n10217 ;
  assign n42407 = n10216 & n42406 ;
  assign n42408 = n10173 & n42407 ;
  assign n42409 = ~\pi0040  & ~\pi0171  ;
  assign n42410 = n1256 & n42409 ;
  assign n42411 = n7597 & n42410 ;
  assign n42412 = ~n42408 & n42411 ;
  assign n42413 = n10277 & ~n42412 ;
  assign n42414 = ~n20686 & n42413 ;
  assign n42415 = ~n42405 & ~n42414 ;
  assign n42416 = ~\pi0192  & n20565 ;
  assign n42417 = ~\pi0192  & ~n20534 ;
  assign n42418 = n20567 & n42417 ;
  assign n42419 = ~n42416 & ~n42418 ;
  assign n42420 = n42415 & n42419 ;
  assign n42421 = n2327 & n20575 ;
  assign n42422 = n42420 & n42421 ;
  assign n42423 = ~n13268 & ~n42422 ;
  assign n42424 = ~\pi0087  & n42423 ;
  assign n42425 = ~n20610 & ~n42424 ;
  assign n42426 = ~n42402 & n42425 ;
  assign n42427 = ~\pi0062  & ~\pi0092  ;
  assign n42428 = ~n42426 & n42427 ;
  assign n42429 = ~n42379 & ~n42428 ;
  assign n42430 = ~\pi0055  & ~\pi0056  ;
  assign n42431 = ~n42429 & n42430 ;
  assign n42432 = \pi0195  & n2467 ;
  assign n42433 = ~n42374 & n42432 ;
  assign n42434 = ~n11149 & n42433 ;
  assign n42435 = ~n20623 & n42434 ;
  assign n42436 = ~n42431 & n42435 ;
  assign n42437 = ~n42378 & ~n42436 ;
  assign n42438 = ~\pi0038  & ~\pi0194  ;
  assign n42439 = ~\pi0039  & n42438 ;
  assign n42440 = \pi0232  & n20565 ;
  assign n42441 = \pi0232  & ~n20534 ;
  assign n42442 = n20567 & n42441 ;
  assign n42443 = ~n42440 & ~n42442 ;
  assign n42444 = ~\pi0040  & ~\pi0170  ;
  assign n42445 = n1256 & n42444 ;
  assign n42446 = n7597 & n42445 ;
  assign n42447 = ~n42408 & n42446 ;
  assign n42448 = n10277 & ~n42447 ;
  assign n42449 = ~n20686 & n42448 ;
  assign n42450 = n42443 & ~n42449 ;
  assign n42451 = n20575 & n42438 ;
  assign n42452 = n42450 & n42451 ;
  assign n42453 = ~n42439 & ~n42452 ;
  assign n42454 = n11239 & ~n42453 ;
  assign n42455 = ~n6706 & ~n11239 ;
  assign n42456 = ~\pi0039  & n42202 ;
  assign n42457 = n10118 & ~n10220 ;
  assign n42458 = ~n20680 & n42457 ;
  assign n42459 = n20575 & ~n42458 ;
  assign n42460 = n42202 & n42450 ;
  assign n42461 = n42459 & n42460 ;
  assign n42462 = ~n42456 & ~n42461 ;
  assign n42463 = n20707 & ~n42462 ;
  assign n42464 = ~n42455 & n42463 ;
  assign n42465 = ~n42454 & ~n42464 ;
  assign n42466 = n10118 & ~n42465 ;
  assign n42467 = ~\pi0100  & ~n20610 ;
  assign n42468 = n42466 & n42467 ;
  assign n42469 = ~n10735 & ~n20191 ;
  assign n42470 = ~n10366 & n20191 ;
  assign n42471 = ~\pi0210  & n20191 ;
  assign n42472 = ~n10375 & n42471 ;
  assign n42473 = ~n42470 & ~n42472 ;
  assign n42474 = n10276 & n42473 ;
  assign n42475 = ~n42469 & n42474 ;
  assign n42476 = n42400 & ~n42475 ;
  assign n42477 = ~\pi0039  & n42476 ;
  assign n42478 = n42453 & n42462 ;
  assign n42479 = n42467 & ~n42478 ;
  assign n42480 = ~n42477 & n42479 ;
  assign n42481 = ~n42468 & ~n42480 ;
  assign n42482 = ~\pi0075  & \pi0087  ;
  assign n42483 = n2327 & n42482 ;
  assign n42484 = n10182 & n42483 ;
  assign n42485 = ~\pi0055  & ~\pi0092  ;
  assign n42486 = ~n42484 & n42485 ;
  assign n42487 = n42481 & n42486 ;
  assign n42488 = ~\pi0055  & n20532 ;
  assign n42489 = n11150 & ~n20617 ;
  assign n42490 = ~n20621 & n42489 ;
  assign n42491 = ~n42488 & n42490 ;
  assign n42492 = ~n42487 & n42491 ;
  assign n42493 = ~n1292 & n2467 ;
  assign n42494 = n10158 & n42493 ;
  assign n42495 = \pi0196  & ~n42494 ;
  assign n42496 = ~n42492 & n42495 ;
  assign n42497 = n13992 & ~n20638 ;
  assign n42498 = n8368 & ~n20641 ;
  assign n42499 = ~n42497 & ~n42498 ;
  assign n42500 = ~n6706 & ~n6713 ;
  assign n42501 = ~\pi0170  & n6706 ;
  assign n42502 = ~n6732 & n42501 ;
  assign n42503 = ~n42500 & ~n42502 ;
  assign n42504 = n11062 & ~n42503 ;
  assign n42505 = n6948 & n42504 ;
  assign n42506 = n16483 & n20646 ;
  assign n42507 = n6921 & n42506 ;
  assign n42508 = \pi0232  & ~n42507 ;
  assign n42509 = ~n42505 & n42508 ;
  assign n42510 = n42499 & ~n42509 ;
  assign n42511 = \pi0039  & \pi0194  ;
  assign n42512 = ~n42510 & n42511 ;
  assign n42513 = n13708 & n20197 ;
  assign n42514 = n10937 & n42513 ;
  assign n42515 = n10319 & n42514 ;
  assign n42516 = ~\pi0039  & \pi0194  ;
  assign n42517 = ~n42515 & n42516 ;
  assign n42518 = ~n42200 & ~n42517 ;
  assign n42519 = n11834 & n42518 ;
  assign n42520 = ~n42512 & n42519 ;
  assign n42521 = ~\pi0196  & ~n42520 ;
  assign n42522 = ~\pi0138  & n20628 ;
  assign n42523 = n16758 & n42522 ;
  assign n42524 = ~n20641 & n27982 ;
  assign n42525 = n13708 & ~n20192 ;
  assign n42526 = n10937 & n42525 ;
  assign n42527 = n10319 & n42526 ;
  assign n42528 = ~\pi0039  & ~n42527 ;
  assign n42529 = ~\pi0038  & ~n42528 ;
  assign n42530 = ~n42524 & n42529 ;
  assign n42531 = ~\pi0194  & ~\pi0196  ;
  assign n42532 = ~n42530 & n42531 ;
  assign n42533 = n2297 & n42531 ;
  assign n42534 = ~n42510 & n42533 ;
  assign n42535 = ~n42532 & ~n42534 ;
  assign n42536 = ~n42523 & n42535 ;
  assign n42537 = ~n42521 & n42536 ;
  assign n42538 = ~n42496 & n42537 ;
  assign n42539 = \pi0195  & ~\pi0196  ;
  assign n42540 = ~n42494 & n42539 ;
  assign n42541 = ~n42492 & n42540 ;
  assign n42542 = ~n42520 & ~n42539 ;
  assign n42543 = ~\pi0194  & ~n42539 ;
  assign n42544 = ~n42530 & n42543 ;
  assign n42545 = n2297 & n42543 ;
  assign n42546 = ~n42510 & n42545 ;
  assign n42547 = ~n42544 & ~n42546 ;
  assign n42548 = n42523 & n42547 ;
  assign n42549 = ~n42542 & n42548 ;
  assign n42550 = ~n42541 & n42549 ;
  assign n42551 = ~n42538 & ~n42550 ;
  assign n42552 = ~\pi0197  & ~n11834 ;
  assign n42553 = ~\pi0832  & ~n42552 ;
  assign n42554 = ~\pi0197  & \pi0767  ;
  assign n42555 = ~\pi0299  & n42554 ;
  assign n42556 = ~n21692 & n42555 ;
  assign n42557 = \pi0039  & ~n42554 ;
  assign n42558 = \pi0039  & ~n21731 ;
  assign n42559 = n21714 & n42558 ;
  assign n42560 = ~n42557 & ~n42559 ;
  assign n42561 = ~n42556 & ~n42560 ;
  assign n42562 = ~\pi0767  & \pi0947  ;
  assign n42563 = \pi0299  & n42562 ;
  assign n42564 = ~n21205 & n42563 ;
  assign n42565 = ~n21238 & n42564 ;
  assign n42566 = ~\pi0299  & n42562 ;
  assign n42567 = ~n21740 & n42566 ;
  assign n42568 = ~n21738 & n42567 ;
  assign n42569 = ~n42565 & ~n42568 ;
  assign n42570 = ~\pi0197  & ~\pi0299  ;
  assign n42571 = n21740 & n42570 ;
  assign n42572 = n21737 & n42570 ;
  assign n42573 = n21232 & n42572 ;
  assign n42574 = ~n42571 & ~n42573 ;
  assign n42575 = ~\pi0197  & \pi0299  ;
  assign n42576 = n21205 & n42575 ;
  assign n42577 = n21237 & n42575 ;
  assign n42578 = n21232 & n42577 ;
  assign n42579 = ~n42576 & ~n42578 ;
  assign n42580 = ~\pi0039  & n42579 ;
  assign n42581 = n42574 & n42580 ;
  assign n42582 = n42569 & n42581 ;
  assign n42583 = ~\pi0038  & ~n42582 ;
  assign n42584 = ~n42561 & n42583 ;
  assign n42585 = ~\pi0197  & ~n21692 ;
  assign n42586 = n27361 & ~n42585 ;
  assign n42587 = ~\pi0767  & ~n42586 ;
  assign n42588 = ~n27304 & ~n42575 ;
  assign n42589 = ~n27260 & ~n42588 ;
  assign n42590 = ~n27258 & n42589 ;
  assign n42591 = \pi0197  & n27304 ;
  assign n42592 = ~\pi0038  & ~n42591 ;
  assign n42593 = ~n42582 & n42592 ;
  assign n42594 = ~n42590 & n42593 ;
  assign n42595 = n42587 & n42594 ;
  assign n42596 = ~n42584 & ~n42595 ;
  assign n42597 = n6784 & ~n42562 ;
  assign n42598 = n1266 & n42597 ;
  assign n42599 = n22706 & n42598 ;
  assign n42600 = n1358 & n42599 ;
  assign n42601 = \pi0038  & ~n42600 ;
  assign n42602 = \pi0698  & ~n42601 ;
  assign n42603 = \pi0197  & \pi0698  ;
  assign n42604 = ~n22123 & n42603 ;
  assign n42605 = ~n42602 & ~n42604 ;
  assign n42606 = n42596 & ~n42605 ;
  assign n42607 = n11834 & ~n42606 ;
  assign n42608 = n42553 & ~n42607 ;
  assign n42609 = ~\pi0197  & ~n27215 ;
  assign n42610 = \pi0197  & ~\pi0299  ;
  assign n42611 = ~n27158 & n42610 ;
  assign n42612 = \pi0197  & \pi0299  ;
  assign n42613 = ~n27172 & n42612 ;
  assign n42614 = ~\pi0767  & ~n42613 ;
  assign n42615 = ~n42611 & n42614 ;
  assign n42616 = ~n42609 & n42615 ;
  assign n42617 = ~\pi0197  & ~n27299 ;
  assign n42618 = n27115 & n42617 ;
  assign n42619 = n27129 & n42617 ;
  assign n42620 = ~n27126 & n42619 ;
  assign n42621 = ~n42618 & ~n42620 ;
  assign n42622 = n24388 & n27077 ;
  assign n42623 = \pi0197  & ~n27072 ;
  assign n42624 = ~n42622 & n42623 ;
  assign n42625 = ~n27259 & n42624 ;
  assign n42626 = \pi0299  & ~n42625 ;
  assign n42627 = n42621 & n42626 ;
  assign n42628 = n27523 & ~n42585 ;
  assign n42629 = \pi0767  & ~n42628 ;
  assign n42630 = ~n42627 & n42629 ;
  assign n42631 = \pi0039  & ~n42630 ;
  assign n42632 = ~n42616 & n42631 ;
  assign n42633 = n27068 & n42569 ;
  assign n42634 = n42581 & n42633 ;
  assign n42635 = ~\pi0038  & ~n42634 ;
  assign n42636 = ~n42632 & n42635 ;
  assign n42637 = ~n26930 & n42600 ;
  assign n42638 = \pi0197  & ~n21757 ;
  assign n42639 = \pi0038  & ~n42638 ;
  assign n42640 = ~n42637 & n42639 ;
  assign n42641 = ~\pi0698  & ~n42640 ;
  assign n42642 = n42553 & n42641 ;
  assign n42643 = ~n42636 & n42642 ;
  assign n42644 = ~n42608 & ~n42643 ;
  assign n42645 = ~\pi0698  & n26930 ;
  assign n42646 = ~n42562 & ~n42645 ;
  assign n42647 = n1689 & ~n42646 ;
  assign n42648 = ~\pi0197  & ~n1689 ;
  assign n42649 = \pi0832  & ~n42648 ;
  assign n42650 = ~n42647 & n42649 ;
  assign n42651 = n42644 & ~n42650 ;
  assign n42652 = ~\pi0198  & ~n9948 ;
  assign n42653 = ~\pi0039  & \pi0198  ;
  assign n42654 = ~n21289 & n42653 ;
  assign n42655 = \pi0039  & \pi0198  ;
  assign n42656 = \pi0038  & ~n42655 ;
  assign n42657 = \pi0634  & \pi0680  ;
  assign n42658 = ~n20854 & n42657 ;
  assign n42659 = n1689 & n42658 ;
  assign n42660 = n1259 & n42659 ;
  assign n42661 = n1281 & n42660 ;
  assign n42662 = ~\pi0039  & n1249 ;
  assign n42663 = n42661 & n42662 ;
  assign n42664 = n42656 & ~n42663 ;
  assign n42665 = ~n42654 & n42664 ;
  assign n42666 = n6861 & ~n42665 ;
  assign n42667 = \pi0198  & n21403 ;
  assign n42668 = ~n21399 & n42667 ;
  assign n42669 = ~n6706 & n42668 ;
  assign n42670 = \pi0634  & ~n20854 ;
  assign n42671 = ~n21285 & n42670 ;
  assign n42672 = ~n6706 & n42671 ;
  assign n42673 = ~n22183 & n42672 ;
  assign n42674 = ~n42669 & ~n42673 ;
  assign n42675 = \pi0198  & n21285 ;
  assign n42676 = ~n42671 & ~n42675 ;
  assign n42677 = n6706 & ~n42676 ;
  assign n42678 = ~n21285 & ~n42670 ;
  assign n42679 = \pi0198  & \pi0634  ;
  assign n42680 = ~\pi0198  & ~n42679 ;
  assign n42681 = n21285 & n42680 ;
  assign n42682 = ~n42678 & ~n42681 ;
  assign n42683 = ~n6712 & n22180 ;
  assign n42684 = n42682 & n42683 ;
  assign n42685 = ~n42677 & ~n42684 ;
  assign n42686 = n42674 & n42685 ;
  assign n42687 = n21285 & n42679 ;
  assign n42688 = ~n42671 & ~n42687 ;
  assign n42689 = ~n6712 & ~n42675 ;
  assign n42690 = n42688 & n42689 ;
  assign n42691 = n22180 & ~n42690 ;
  assign n42692 = ~n6709 & ~n42691 ;
  assign n42693 = ~n42686 & ~n42692 ;
  assign n42694 = n21520 & n21908 ;
  assign n42695 = ~n21399 & n21420 ;
  assign n42696 = ~n42694 & ~n42695 ;
  assign n42697 = ~n21352 & ~n21405 ;
  assign n42698 = \pi0198  & ~\pi0680  ;
  assign n42699 = ~n42697 & n42698 ;
  assign n42700 = ~n42696 & n42699 ;
  assign n42701 = n6761 & ~n42700 ;
  assign n42702 = ~n42693 & n42701 ;
  assign n42703 = n6735 & ~n42682 ;
  assign n42704 = ~n22183 & n42671 ;
  assign n42705 = n6706 & ~n6712 ;
  assign n42706 = ~n42668 & n42705 ;
  assign n42707 = ~n42704 & n42706 ;
  assign n42708 = ~n42703 & ~n42707 ;
  assign n42709 = n6712 & ~n42668 ;
  assign n42710 = ~n42704 & n42709 ;
  assign n42711 = n22180 & ~n42710 ;
  assign n42712 = n42708 & n42711 ;
  assign n42713 = n42695 & n42698 ;
  assign n42714 = n21908 & n42698 ;
  assign n42715 = n21520 & n42714 ;
  assign n42716 = ~n42713 & ~n42715 ;
  assign n42717 = n6709 & n42668 ;
  assign n42718 = n6709 & n42671 ;
  assign n42719 = ~n22183 & n42718 ;
  assign n42720 = ~n42717 & ~n42719 ;
  assign n42721 = ~n6761 & n42720 ;
  assign n42722 = n42716 & n42721 ;
  assign n42723 = ~n42712 & n42722 ;
  assign n42724 = ~n42702 & ~n42723 ;
  assign n42725 = \pi0223  & n42724 ;
  assign n42726 = n2165 & ~n42658 ;
  assign n42727 = ~n21285 & n42726 ;
  assign n42728 = ~\pi0198  & n2165 ;
  assign n42729 = n21285 & n42728 ;
  assign n42730 = ~n42727 & ~n42729 ;
  assign n42731 = ~\pi0223  & n42730 ;
  assign n42732 = \pi0039  & ~n42731 ;
  assign n42733 = ~n42725 & n42732 ;
  assign n42734 = \pi0634  & ~n6706 ;
  assign n42735 = ~n22293 & n42734 ;
  assign n42736 = \pi0198  & ~n21291 ;
  assign n42737 = ~\pi0120  & \pi0198  ;
  assign n42738 = ~n21304 & n42737 ;
  assign n42739 = ~n42736 & ~n42738 ;
  assign n42740 = ~n6706 & ~n42739 ;
  assign n42741 = ~n21903 & n42740 ;
  assign n42742 = ~n42677 & ~n42741 ;
  assign n42743 = ~n42735 & n42742 ;
  assign n42744 = n6709 & ~n42743 ;
  assign n42745 = n21285 & n42698 ;
  assign n42746 = n6712 & n42698 ;
  assign n42747 = ~n42745 & ~n42746 ;
  assign n42748 = ~n22033 & ~n42747 ;
  assign n42749 = ~n42744 & ~n42748 ;
  assign n42750 = n6712 & ~n42677 ;
  assign n42751 = ~n42741 & n42750 ;
  assign n42752 = ~n42735 & n42751 ;
  assign n42753 = n42691 & ~n42752 ;
  assign n42754 = ~n2165 & ~n42753 ;
  assign n42755 = n42749 & n42754 ;
  assign n42756 = ~n21275 & ~n42755 ;
  assign n42757 = \pi0039  & ~n42725 ;
  assign n42758 = ~n6706 & ~n42682 ;
  assign n42759 = n6706 & n42739 ;
  assign n42760 = n6706 & ~n21290 ;
  assign n42761 = ~n21325 & n42760 ;
  assign n42762 = ~n42759 & ~n42761 ;
  assign n42763 = ~n42758 & n42762 ;
  assign n42764 = \pi0634  & ~n42758 ;
  assign n42765 = ~n22293 & n42764 ;
  assign n42766 = ~n42763 & ~n42765 ;
  assign n42767 = ~n6712 & n42766 ;
  assign n42768 = n6712 & n42739 ;
  assign n42769 = n6712 & ~n21290 ;
  assign n42770 = ~n21325 & n42769 ;
  assign n42771 = ~n42768 & ~n42770 ;
  assign n42772 = n22180 & n42771 ;
  assign n42773 = \pi0634  & n22180 ;
  assign n42774 = ~n22293 & n42773 ;
  assign n42775 = ~n42772 & ~n42774 ;
  assign n42776 = ~n6761 & ~n42775 ;
  assign n42777 = ~n42767 & n42776 ;
  assign n42778 = n21905 & n42698 ;
  assign n42779 = n21328 & n42714 ;
  assign n42780 = ~n42778 & ~n42779 ;
  assign n42781 = n6709 & ~n42739 ;
  assign n42782 = ~n21903 & n42781 ;
  assign n42783 = \pi0634  & n6709 ;
  assign n42784 = ~n22293 & n42783 ;
  assign n42785 = ~n42782 & ~n42784 ;
  assign n42786 = n42780 & n42785 ;
  assign n42787 = ~n6761 & ~n42786 ;
  assign n42788 = ~n42777 & ~n42787 ;
  assign n42789 = n42757 & n42788 ;
  assign n42790 = ~n42756 & n42789 ;
  assign n42791 = ~n42733 & ~n42790 ;
  assign n42792 = \pi0198  & n1686 ;
  assign n42793 = \pi0198  & \pi1093  ;
  assign n42794 = ~n21229 & n42793 ;
  assign n42795 = ~n42792 & ~n42794 ;
  assign n42796 = n21995 & ~n42795 ;
  assign n42797 = ~n22102 & n42657 ;
  assign n42798 = ~n42796 & n42797 ;
  assign n42799 = ~\pi0039  & ~n21738 ;
  assign n42800 = ~n42798 & n42799 ;
  assign n42801 = ~\pi0299  & ~n42800 ;
  assign n42802 = n42791 & n42801 ;
  assign n42803 = ~\pi0038  & ~n42802 ;
  assign n42804 = ~n2352 & ~n42753 ;
  assign n42805 = n42749 & n42804 ;
  assign n42806 = ~n21444 & ~n42805 ;
  assign n42807 = n6732 & ~n42700 ;
  assign n42808 = ~n42693 & n42807 ;
  assign n42809 = ~n6732 & n42720 ;
  assign n42810 = n42716 & n42809 ;
  assign n42811 = ~n42712 & n42810 ;
  assign n42812 = \pi0215  & ~n42811 ;
  assign n42813 = ~n42808 & n42812 ;
  assign n42814 = ~n6732 & ~n42786 ;
  assign n42815 = ~n6732 & ~n42775 ;
  assign n42816 = ~n42767 & n42815 ;
  assign n42817 = ~n42814 & ~n42816 ;
  assign n42818 = ~n42813 & n42817 ;
  assign n42819 = ~n42806 & n42818 ;
  assign n42820 = n2352 & ~n42658 ;
  assign n42821 = ~n21285 & n42820 ;
  assign n42822 = ~\pi0198  & n2352 ;
  assign n42823 = n21285 & n42822 ;
  assign n42824 = ~n42821 & ~n42823 ;
  assign n42825 = ~\pi0215  & n42824 ;
  assign n42826 = \pi0039  & n42825 ;
  assign n42827 = \pi0039  & ~n42808 ;
  assign n42828 = n42812 & n42827 ;
  assign n42829 = ~n42826 & ~n42828 ;
  assign n42830 = ~n42819 & ~n42829 ;
  assign n42831 = ~\pi0198  & ~n22097 ;
  assign n42832 = ~n22095 & n42831 ;
  assign n42833 = \pi0198  & \pi0210  ;
  assign n42834 = n22002 & n42833 ;
  assign n42835 = \pi0198  & ~\pi0210  ;
  assign n42836 = ~n21996 & n42835 ;
  assign n42837 = n42657 & ~n42836 ;
  assign n42838 = ~n42834 & n42837 ;
  assign n42839 = ~n42832 & n42838 ;
  assign n42840 = ~n21205 & ~n42657 ;
  assign n42841 = ~n21238 & n42840 ;
  assign n42842 = ~\pi0198  & ~n42657 ;
  assign n42843 = ~\pi0039  & ~n42842 ;
  assign n42844 = ~n42841 & n42843 ;
  assign n42845 = ~n42839 & n42844 ;
  assign n42846 = ~n42830 & ~n42845 ;
  assign n42847 = \pi0299  & ~n42846 ;
  assign n42848 = n42803 & ~n42847 ;
  assign n42849 = n42666 & ~n42848 ;
  assign n42850 = ~\pi0198  & \pi0625  ;
  assign n42851 = ~n22727 & ~n42850 ;
  assign n42852 = ~n42849 & ~n42851 ;
  assign n42853 = \pi0198  & ~n6732 ;
  assign n42854 = n21334 & n42853 ;
  assign n42855 = ~n21330 & n42854 ;
  assign n42856 = ~n6713 & ~n21352 ;
  assign n42857 = n21355 & n42856 ;
  assign n42858 = ~n21290 & n42856 ;
  assign n42859 = ~n21325 & n42858 ;
  assign n42860 = ~n42857 & ~n42859 ;
  assign n42861 = ~\pi0198  & ~n6713 ;
  assign n42862 = ~n6713 & n6732 ;
  assign n42863 = \pi0198  & n6732 ;
  assign n42864 = n21285 & n42863 ;
  assign n42865 = ~n42862 & ~n42864 ;
  assign n42866 = ~n42861 & ~n42865 ;
  assign n42867 = n42860 & n42866 ;
  assign n42868 = ~n2352 & ~n42867 ;
  assign n42869 = ~n42855 & n42868 ;
  assign n42870 = \pi0198  & ~\pi0215  ;
  assign n42871 = n21285 & n42870 ;
  assign n42872 = ~n24388 & ~n42871 ;
  assign n42873 = ~n42869 & ~n42872 ;
  assign n42874 = n42695 & n42853 ;
  assign n42875 = n21908 & n42853 ;
  assign n42876 = n21520 & n42875 ;
  assign n42877 = ~n42874 & ~n42876 ;
  assign n42878 = n6713 & ~n42675 ;
  assign n42879 = \pi0198  & ~n42878 ;
  assign n42880 = ~n42697 & n42879 ;
  assign n42881 = \pi0299  & ~n42880 ;
  assign n42882 = n42877 & n42881 ;
  assign n42883 = ~n21948 & ~n42882 ;
  assign n42884 = ~n42873 & ~n42883 ;
  assign n42885 = \pi0198  & ~n6761 ;
  assign n42886 = n42695 & n42885 ;
  assign n42887 = n21908 & n42885 ;
  assign n42888 = n21520 & n42887 ;
  assign n42889 = ~n42886 & ~n42888 ;
  assign n42890 = ~\pi0299  & ~n42880 ;
  assign n42891 = n42889 & n42890 ;
  assign n42892 = n2511 & n12968 ;
  assign n42893 = ~n3058 & n42892 ;
  assign n42894 = ~n42891 & n42893 ;
  assign n42895 = n21334 & n42885 ;
  assign n42896 = ~n21330 & n42895 ;
  assign n42897 = ~n6713 & n6761 ;
  assign n42898 = \pi0198  & n6761 ;
  assign n42899 = n21285 & n42898 ;
  assign n42900 = ~n42897 & ~n42899 ;
  assign n42901 = ~n42861 & ~n42900 ;
  assign n42902 = n42860 & n42901 ;
  assign n42903 = ~n2165 & ~n42902 ;
  assign n42904 = ~n42896 & n42903 ;
  assign n42905 = \pi0198  & ~\pi0223  ;
  assign n42906 = n21285 & n42905 ;
  assign n42907 = ~n22316 & ~n42906 ;
  assign n42908 = n42892 & ~n42907 ;
  assign n42909 = ~n42904 & n42908 ;
  assign n42910 = ~n42894 & ~n42909 ;
  assign n42911 = ~n42884 & ~n42910 ;
  assign n42912 = ~\pi0198  & ~n42911 ;
  assign n42913 = n1288 & ~n27217 ;
  assign n42914 = ~n27219 & n42913 ;
  assign n42915 = ~n21768 & ~n42911 ;
  assign n42916 = ~n42914 & n42915 ;
  assign n42917 = ~n42912 & ~n42916 ;
  assign n42918 = ~\pi0625  & ~n42917 ;
  assign n42919 = \pi1153  & ~n42918 ;
  assign n42920 = ~n42852 & n42919 ;
  assign n42921 = ~\pi0198  & ~\pi0625  ;
  assign n42922 = ~n22734 & ~n42921 ;
  assign n42923 = ~n42849 & ~n42922 ;
  assign n42924 = ~\pi1153  & ~n42912 ;
  assign n42925 = ~n42916 & n42924 ;
  assign n42926 = ~n24561 & ~n42925 ;
  assign n42927 = ~n42923 & ~n42926 ;
  assign n42928 = ~n42920 & ~n42927 ;
  assign n42929 = n26065 & ~n42928 ;
  assign n42930 = \pi0198  & ~n6861 ;
  assign n42931 = ~\pi0778  & n42930 ;
  assign n42932 = ~\pi0778  & n42666 ;
  assign n42933 = ~n42848 & n42932 ;
  assign n42934 = ~n42931 & ~n42933 ;
  assign n42935 = n23885 & ~n42934 ;
  assign n42936 = ~n23885 & ~n42912 ;
  assign n42937 = ~n42916 & n42936 ;
  assign n42938 = ~n42935 & ~n42937 ;
  assign n42939 = ~n42929 & n42938 ;
  assign n42940 = ~\pi0792  & ~n42939 ;
  assign n42941 = ~\pi0647  & ~n42940 ;
  assign n42942 = ~\pi1157  & ~n42912 ;
  assign n42943 = ~n42916 & n42942 ;
  assign n42944 = ~n22945 & ~n42943 ;
  assign n42945 = ~n42941 & ~n42944 ;
  assign n42946 = ~\pi0628  & ~n42937 ;
  assign n42947 = ~n42935 & n42946 ;
  assign n42948 = ~n42929 & n42947 ;
  assign n42949 = ~\pi0628  & ~\pi1156  ;
  assign n42950 = ~\pi1156  & ~n42912 ;
  assign n42951 = ~n42916 & n42950 ;
  assign n42952 = ~n42949 & ~n42951 ;
  assign n42953 = ~n42948 & ~n42952 ;
  assign n42954 = \pi0628  & ~n42937 ;
  assign n42955 = ~n42935 & n42954 ;
  assign n42956 = ~n42929 & n42955 ;
  assign n42957 = \pi0628  & \pi1156  ;
  assign n42958 = \pi1156  & ~n42912 ;
  assign n42959 = ~n42916 & n42958 ;
  assign n42960 = ~n42957 & ~n42959 ;
  assign n42961 = ~n42956 & ~n42960 ;
  assign n42962 = ~n42953 & ~n42961 ;
  assign n42963 = \pi0792  & ~n42944 ;
  assign n42964 = ~n42962 & n42963 ;
  assign n42965 = ~n42945 & ~n42964 ;
  assign n42966 = \pi0647  & ~n42940 ;
  assign n42967 = \pi1157  & ~n42912 ;
  assign n42968 = ~n42916 & n42967 ;
  assign n42969 = ~n20925 & ~n42968 ;
  assign n42970 = ~n42966 & ~n42969 ;
  assign n42971 = \pi0792  & ~n42969 ;
  assign n42972 = ~n42962 & n42971 ;
  assign n42973 = ~n42970 & ~n42972 ;
  assign n42974 = n42965 & n42973 ;
  assign n42975 = ~n20811 & ~n42917 ;
  assign n42976 = n23424 & n42975 ;
  assign n42977 = ~\pi0198  & ~n21473 ;
  assign n42978 = ~n21472 & n42977 ;
  assign n42979 = n21247 & n42833 ;
  assign n42980 = \pi0603  & \pi0633  ;
  assign n42981 = ~n21241 & n42835 ;
  assign n42982 = n42980 & ~n42981 ;
  assign n42983 = ~n42979 & n42982 ;
  assign n42984 = ~n42978 & n42983 ;
  assign n42985 = ~n21205 & ~n42980 ;
  assign n42986 = ~n21238 & n42985 ;
  assign n42987 = ~\pi0198  & ~n42980 ;
  assign n42988 = ~\pi0039  & ~n42987 ;
  assign n42989 = ~n42986 & n42988 ;
  assign n42990 = ~n42984 & n42989 ;
  assign n42991 = \pi0633  & ~n20783 ;
  assign n42992 = \pi0603  & n42991 ;
  assign n42993 = ~n21285 & n42992 ;
  assign n42994 = ~n42675 & ~n42993 ;
  assign n42995 = ~n21370 & n42994 ;
  assign n42996 = n21258 & n21285 ;
  assign n42997 = n21370 & ~n42996 ;
  assign n42998 = ~n42995 & ~n42997 ;
  assign n42999 = ~n6709 & n42998 ;
  assign n43000 = \pi0198  & ~n42697 ;
  assign n43001 = n6706 & n42991 ;
  assign n43002 = ~n21285 & n43001 ;
  assign n43003 = \pi0198  & n6706 ;
  assign n43004 = n21285 & n43003 ;
  assign n43005 = ~n43002 & ~n43004 ;
  assign n43006 = ~n21285 & n42991 ;
  assign n43007 = ~n22183 & n43006 ;
  assign n43008 = n43005 & ~n43007 ;
  assign n43009 = ~n43000 & n43008 ;
  assign n43010 = \pi0603  & ~n42995 ;
  assign n43011 = ~n6709 & n43010 ;
  assign n43012 = ~n43009 & n43011 ;
  assign n43013 = ~n42999 & ~n43012 ;
  assign n43014 = ~\pi0603  & ~n21352 ;
  assign n43015 = ~n21405 & n43014 ;
  assign n43016 = ~n21256 & ~n43015 ;
  assign n43017 = n6709 & n43016 ;
  assign n43018 = ~n43009 & n43017 ;
  assign n43019 = n6732 & ~n43018 ;
  assign n43020 = n43013 & n43019 ;
  assign n43021 = \pi0633  & n21515 ;
  assign n43022 = \pi0633  & n21516 ;
  assign n43023 = ~n21520 & n43022 ;
  assign n43024 = ~n43021 & ~n43023 ;
  assign n43025 = n21526 & ~n43024 ;
  assign n43026 = \pi0198  & ~n6709 ;
  assign n43027 = n42695 & n43026 ;
  assign n43028 = n21908 & n43026 ;
  assign n43029 = n21520 & n43028 ;
  assign n43030 = ~n43027 & ~n43029 ;
  assign n43031 = ~n43025 & n43030 ;
  assign n43032 = n6709 & n21425 ;
  assign n43033 = ~n6732 & ~n43032 ;
  assign n43034 = ~n6732 & ~n42668 ;
  assign n43035 = ~n43007 & n43034 ;
  assign n43036 = ~n43033 & ~n43035 ;
  assign n43037 = n43031 & ~n43036 ;
  assign n43038 = n23979 & ~n43037 ;
  assign n43039 = ~n43020 & n43038 ;
  assign n43040 = n2352 & n42994 ;
  assign n43041 = \pi0039  & ~\pi0215  ;
  assign n43042 = ~n43040 & n43041 ;
  assign n43043 = ~n43039 & ~n43042 ;
  assign n43044 = \pi0633  & ~n6706 ;
  assign n43045 = ~n21346 & n43044 ;
  assign n43046 = ~\pi0642  & n43005 ;
  assign n43047 = ~n42741 & n43046 ;
  assign n43048 = ~n43045 & n43047 ;
  assign n43049 = ~\pi0603  & ~\pi0642  ;
  assign n43050 = ~\pi0642  & n6711 ;
  assign n43051 = \pi0603  & n6711 ;
  assign n43052 = n42991 & n43051 ;
  assign n43053 = ~n21285 & n43052 ;
  assign n43054 = \pi0198  & n43051 ;
  assign n43055 = n21285 & n43054 ;
  assign n43056 = ~n43053 & ~n43055 ;
  assign n43057 = ~n43050 & n43056 ;
  assign n43058 = ~n43049 & ~n43057 ;
  assign n43059 = ~n43048 & n43058 ;
  assign n43060 = \pi0603  & ~n6711 ;
  assign n43061 = n42991 & n43060 ;
  assign n43062 = ~n21285 & n43061 ;
  assign n43063 = \pi0198  & n43060 ;
  assign n43064 = n21285 & n43063 ;
  assign n43065 = ~n43062 & ~n43064 ;
  assign n43066 = ~n6709 & ~n42996 ;
  assign n43067 = n43065 & n43066 ;
  assign n43068 = ~n43059 & n43067 ;
  assign n43069 = n21258 & n21359 ;
  assign n43070 = n6709 & ~n43069 ;
  assign n43071 = n6732 & ~n43070 ;
  assign n43072 = ~n42741 & n43005 ;
  assign n43073 = ~n43045 & n43072 ;
  assign n43074 = \pi0603  & n6732 ;
  assign n43075 = ~n43073 & n43074 ;
  assign n43076 = ~n43071 & ~n43075 ;
  assign n43077 = ~n43068 & ~n43076 ;
  assign n43078 = \pi0603  & ~n42739 ;
  assign n43079 = ~n21903 & n43078 ;
  assign n43080 = n21370 & n43079 ;
  assign n43081 = n21370 & n42980 ;
  assign n43082 = ~n21346 & n43081 ;
  assign n43083 = ~n43080 & ~n43082 ;
  assign n43084 = n21258 & ~n21286 ;
  assign n43085 = n21328 & n43084 ;
  assign n43086 = n43083 & ~n43085 ;
  assign n43087 = ~n6706 & ~n42991 ;
  assign n43088 = ~n21285 & n43087 ;
  assign n43089 = n10570 & n21285 ;
  assign n43090 = ~n43088 & ~n43089 ;
  assign n43091 = \pi0603  & ~n21370 ;
  assign n43092 = n43090 & n43091 ;
  assign n43093 = n42762 & n43092 ;
  assign n43094 = \pi0633  & n43092 ;
  assign n43095 = ~n21346 & n43094 ;
  assign n43096 = ~n43093 & ~n43095 ;
  assign n43097 = ~n6709 & n43096 ;
  assign n43098 = n43086 & n43097 ;
  assign n43099 = ~n21346 & n42980 ;
  assign n43100 = n6709 & n42739 ;
  assign n43101 = n6709 & ~n21290 ;
  assign n43102 = ~n21325 & n43101 ;
  assign n43103 = ~n43100 & ~n43102 ;
  assign n43104 = ~n43079 & ~n43103 ;
  assign n43105 = ~n43099 & n43104 ;
  assign n43106 = ~n6732 & ~n43105 ;
  assign n43107 = ~n43098 & n43106 ;
  assign n43108 = ~n43077 & ~n43107 ;
  assign n43109 = ~n2352 & ~n43039 ;
  assign n43110 = n43108 & n43109 ;
  assign n43111 = ~n43043 & ~n43110 ;
  assign n43112 = \pi0299  & ~n43111 ;
  assign n43113 = ~n42990 & n43112 ;
  assign n43114 = n6761 & ~n43018 ;
  assign n43115 = n43013 & n43114 ;
  assign n43116 = ~n6761 & ~n43032 ;
  assign n43117 = ~n6761 & ~n42668 ;
  assign n43118 = ~n43007 & n43117 ;
  assign n43119 = ~n43116 & ~n43118 ;
  assign n43120 = n43031 & ~n43119 ;
  assign n43121 = \pi0039  & \pi0223  ;
  assign n43122 = ~n43120 & n43121 ;
  assign n43123 = ~n43115 & n43122 ;
  assign n43124 = \pi0603  & ~n43073 ;
  assign n43125 = n43070 & ~n43124 ;
  assign n43126 = ~n43068 & ~n43125 ;
  assign n43127 = n6761 & n43126 ;
  assign n43128 = ~n6761 & ~n43105 ;
  assign n43129 = ~n43098 & n43128 ;
  assign n43130 = ~n2165 & ~n43129 ;
  assign n43131 = ~n43127 & n43130 ;
  assign n43132 = n2165 & n42994 ;
  assign n43133 = ~\pi0223  & ~n43132 ;
  assign n43134 = \pi0039  & n43133 ;
  assign n43135 = ~n43131 & n43134 ;
  assign n43136 = ~n43123 & ~n43135 ;
  assign n43137 = ~\pi0198  & \pi0633  ;
  assign n43138 = ~n21255 & n43137 ;
  assign n43139 = \pi0198  & \pi0633  ;
  assign n43140 = n21247 & n43139 ;
  assign n43141 = ~n43138 & ~n43140 ;
  assign n43142 = ~n21738 & n43141 ;
  assign n43143 = ~\pi0039  & ~n21257 ;
  assign n43144 = ~n21264 & n43143 ;
  assign n43145 = ~n43142 & n43144 ;
  assign n43146 = ~\pi0299  & ~n43145 ;
  assign n43147 = n43136 & n43146 ;
  assign n43148 = ~n43113 & ~n43147 ;
  assign n43149 = ~\pi0038  & ~\pi0198  ;
  assign n43150 = n1287 & n15409 ;
  assign n43151 = ~n43149 & ~n43150 ;
  assign n43152 = ~n43148 & ~n43151 ;
  assign n43153 = ~n20783 & n42980 ;
  assign n43154 = n1689 & n43153 ;
  assign n43155 = n1259 & n43154 ;
  assign n43156 = n1249 & n43155 ;
  assign n43157 = n24145 & n43156 ;
  assign n43158 = n42656 & ~n43157 ;
  assign n43159 = ~n42654 & n43158 ;
  assign n43160 = n6861 & ~n43159 ;
  assign n43161 = ~n42930 & ~n43160 ;
  assign n43162 = n21777 & ~n43161 ;
  assign n43163 = ~n43152 & n43162 ;
  assign n43164 = ~n21777 & ~n42912 ;
  assign n43165 = ~n42916 & n43164 ;
  assign n43166 = n20811 & ~n43165 ;
  assign n43167 = n23424 & n43166 ;
  assign n43168 = ~n43163 & n43167 ;
  assign n43169 = ~n42976 & ~n43168 ;
  assign n43170 = ~\pi0781  & ~n43165 ;
  assign n43171 = ~n23423 & n43170 ;
  assign n43172 = ~n43163 & n43171 ;
  assign n43173 = ~n26824 & ~n31378 ;
  assign n43174 = ~n23880 & ~n43173 ;
  assign n43175 = n21092 & n43174 ;
  assign n43176 = ~n23423 & n43175 ;
  assign n43177 = ~n42912 & n43175 ;
  assign n43178 = ~n42916 & n43177 ;
  assign n43179 = ~n43176 & ~n43178 ;
  assign n43180 = ~n43172 & ~n43179 ;
  assign n43181 = n43169 & n43180 ;
  assign n43182 = ~n42912 & ~n43175 ;
  assign n43183 = ~n42916 & n43182 ;
  assign n43184 = ~n23414 & ~n43183 ;
  assign n43185 = ~n43181 & n43184 ;
  assign n43186 = \pi0787  & ~n43185 ;
  assign n43187 = ~n42974 & n43186 ;
  assign n43188 = n30425 & ~n42939 ;
  assign n43189 = n23518 & ~n43188 ;
  assign n43190 = ~n43185 & ~n43189 ;
  assign n43191 = n23011 & ~n43185 ;
  assign n43192 = ~n42962 & n43191 ;
  assign n43193 = ~n43190 & ~n43192 ;
  assign n43194 = \pi0790  & n43193 ;
  assign n43195 = ~n43187 & n43194 ;
  assign n43196 = ~\pi0628  & ~n42917 ;
  assign n43197 = n20843 & ~n43196 ;
  assign n43198 = ~n42956 & n43197 ;
  assign n43199 = \pi0629  & ~n42952 ;
  assign n43200 = ~n42948 & n43199 ;
  assign n43201 = ~n43198 & ~n43200 ;
  assign n43202 = \pi0792  & ~n43201 ;
  assign n43203 = ~n23423 & ~n23880 ;
  assign n43204 = ~n23880 & ~n42912 ;
  assign n43205 = ~n42916 & n43204 ;
  assign n43206 = ~n43203 & ~n43205 ;
  assign n43207 = ~n43172 & ~n43206 ;
  assign n43208 = n43169 & n43207 ;
  assign n43209 = n23880 & ~n42912 ;
  assign n43210 = ~n42916 & n43209 ;
  assign n43211 = ~n43208 & ~n43210 ;
  assign n43212 = ~n39249 & ~n43211 ;
  assign n43213 = ~n43202 & ~n43212 ;
  assign n43214 = ~n21067 & ~n43213 ;
  assign n43215 = ~\pi0625  & n43161 ;
  assign n43216 = ~\pi0625  & ~n43151 ;
  assign n43217 = ~n43148 & n43216 ;
  assign n43218 = ~n43215 & ~n43217 ;
  assign n43219 = \pi1153  & n43218 ;
  assign n43220 = \pi0608  & n42926 ;
  assign n43221 = \pi0608  & ~n42922 ;
  assign n43222 = ~n42849 & n43221 ;
  assign n43223 = ~n43220 & ~n43222 ;
  assign n43224 = ~n43219 & ~n43223 ;
  assign n43225 = \pi0198  & ~n21289 ;
  assign n43226 = n1281 & n43156 ;
  assign n43227 = \pi0634  & n24389 ;
  assign n43228 = n1281 & n43227 ;
  assign n43229 = n1260 & n43228 ;
  assign n43230 = ~n43226 & ~n43229 ;
  assign n43231 = ~n43225 & n43230 ;
  assign n43232 = n42656 & n43231 ;
  assign n43233 = ~\pi0198  & n12883 ;
  assign n43234 = n6861 & ~n43233 ;
  assign n43235 = ~n43232 & n43234 ;
  assign n43236 = \pi0038  & n43235 ;
  assign n43237 = ~\pi0680  & ~n21257 ;
  assign n43238 = ~n21264 & n43237 ;
  assign n43239 = ~n43142 & n43238 ;
  assign n43240 = ~\pi0299  & ~n43239 ;
  assign n43241 = ~\pi0603  & ~n21738 ;
  assign n43242 = ~n42798 & n43241 ;
  assign n43243 = \pi0680  & ~n43242 ;
  assign n43244 = ~\pi0039  & ~n43243 ;
  assign n43245 = \pi0634  & ~\pi0665  ;
  assign n43246 = \pi0198  & ~\pi0633  ;
  assign n43247 = n43245 & ~n43246 ;
  assign n43248 = \pi0603  & ~n43247 ;
  assign n43249 = ~\pi0198  & \pi0603  ;
  assign n43250 = ~n21241 & n43249 ;
  assign n43251 = ~n43248 & ~n43250 ;
  assign n43252 = \pi0633  & ~n43251 ;
  assign n43253 = n22002 & n42679 ;
  assign n43254 = n21263 & n43253 ;
  assign n43255 = \pi0198  & ~\pi0634  ;
  assign n43256 = n21236 & n43255 ;
  assign n43257 = n21232 & n43256 ;
  assign n43258 = ~n43251 & ~n43257 ;
  assign n43259 = ~n43254 & n43258 ;
  assign n43260 = ~n43252 & ~n43259 ;
  assign n43261 = ~\pi0039  & n43141 ;
  assign n43262 = ~n43260 & n43261 ;
  assign n43263 = ~n43244 & ~n43262 ;
  assign n43264 = n43240 & ~n43263 ;
  assign n43265 = ~n42657 & ~n42987 ;
  assign n43266 = ~n42986 & n43265 ;
  assign n43267 = ~n42984 & n43266 ;
  assign n43268 = ~n42657 & ~n43267 ;
  assign n43269 = ~n42979 & ~n42981 ;
  assign n43270 = ~n42978 & n43269 ;
  assign n43271 = \pi0198  & ~\pi0665  ;
  assign n43272 = \pi0633  & ~n43271 ;
  assign n43273 = ~n42832 & n43272 ;
  assign n43274 = n43270 & n43273 ;
  assign n43275 = ~\pi0210  & ~n21241 ;
  assign n43276 = ~\pi0198  & ~\pi0665  ;
  assign n43277 = ~n43275 & n43276 ;
  assign n43278 = ~\pi0633  & ~n43277 ;
  assign n43279 = \pi0210  & ~\pi0633  ;
  assign n43280 = n21247 & n43279 ;
  assign n43281 = ~n43278 & ~n43280 ;
  assign n43282 = \pi0603  & n43281 ;
  assign n43283 = ~n21472 & ~n21473 ;
  assign n43284 = \pi0603  & n42836 ;
  assign n43285 = \pi0603  & n42833 ;
  assign n43286 = n22002 & n43285 ;
  assign n43287 = ~n43284 & ~n43286 ;
  assign n43288 = ~n43283 & ~n43287 ;
  assign n43289 = ~n43282 & ~n43288 ;
  assign n43290 = ~n43274 & ~n43289 ;
  assign n43291 = ~n42834 & ~n42836 ;
  assign n43292 = ~n42832 & n43291 ;
  assign n43293 = ~\pi0603  & ~n43292 ;
  assign n43294 = ~n43267 & ~n43293 ;
  assign n43295 = ~n43290 & n43294 ;
  assign n43296 = ~n43268 & ~n43295 ;
  assign n43297 = n21471 & ~n43296 ;
  assign n43298 = ~n43264 & ~n43297 ;
  assign n43299 = ~\pi0680  & n42998 ;
  assign n43300 = ~\pi0680  & n43010 ;
  assign n43301 = ~n43009 & n43300 ;
  assign n43302 = ~n43299 & ~n43301 ;
  assign n43303 = n21403 & n43255 ;
  assign n43304 = ~n21399 & n43303 ;
  assign n43305 = ~n6706 & n43304 ;
  assign n43306 = ~n6706 & n43006 ;
  assign n43307 = ~n22183 & n43306 ;
  assign n43308 = ~n43305 & ~n43307 ;
  assign n43309 = n20783 & n43271 ;
  assign n43310 = ~n21390 & n43276 ;
  assign n43311 = ~n43309 & ~n43310 ;
  assign n43312 = ~n42668 & n43311 ;
  assign n43313 = n42734 & ~n43312 ;
  assign n43314 = n43308 & ~n43313 ;
  assign n43315 = ~n42675 & ~n43006 ;
  assign n43316 = n20783 & n43245 ;
  assign n43317 = ~n21285 & n43316 ;
  assign n43318 = \pi0603  & ~n43317 ;
  assign n43319 = n43315 & n43318 ;
  assign n43320 = ~n21363 & ~n43319 ;
  assign n43321 = n43314 & ~n43320 ;
  assign n43322 = ~\pi0603  & ~n42677 ;
  assign n43323 = n42674 & n43322 ;
  assign n43324 = n6709 & ~n43323 ;
  assign n43325 = ~n43321 & n43324 ;
  assign n43326 = n43302 & ~n43325 ;
  assign n43327 = ~\pi0603  & ~n42676 ;
  assign n43328 = n21370 & ~n43327 ;
  assign n43329 = ~\pi0603  & n43328 ;
  assign n43330 = n43315 & ~n43317 ;
  assign n43331 = n6706 & ~n43330 ;
  assign n43332 = n43328 & ~n43331 ;
  assign n43333 = n43314 & n43332 ;
  assign n43334 = ~n43329 & ~n43333 ;
  assign n43335 = \pi0603  & ~n43330 ;
  assign n43336 = ~n21370 & ~n43327 ;
  assign n43337 = ~n43335 & n43336 ;
  assign n43338 = n22180 & ~n43337 ;
  assign n43339 = n43334 & n43338 ;
  assign n43340 = n6761 & ~n43339 ;
  assign n43341 = n43326 & n43340 ;
  assign n43342 = ~n6706 & ~n43317 ;
  assign n43343 = n43315 & n43342 ;
  assign n43344 = n43091 & ~n43343 ;
  assign n43345 = ~n6712 & ~n43344 ;
  assign n43346 = ~n43007 & ~n43304 ;
  assign n43347 = \pi0634  & ~n43312 ;
  assign n43348 = n43346 & ~n43347 ;
  assign n43349 = ~n43345 & ~n43348 ;
  assign n43350 = ~n6706 & n43091 ;
  assign n43351 = n43317 & n43350 ;
  assign n43352 = ~n43315 & n43350 ;
  assign n43353 = ~n43351 & ~n43352 ;
  assign n43354 = n6706 & ~n42668 ;
  assign n43355 = ~n42704 & n43354 ;
  assign n43356 = ~\pi0603  & ~n42758 ;
  assign n43357 = ~n43355 & n43356 ;
  assign n43358 = n43353 & ~n43357 ;
  assign n43359 = ~n43349 & n43358 ;
  assign n43360 = n22180 & ~n43359 ;
  assign n43361 = \pi0603  & ~n43304 ;
  assign n43362 = ~n43007 & n43361 ;
  assign n43363 = ~n43347 & n43362 ;
  assign n43364 = ~\pi0603  & ~n42668 ;
  assign n43365 = ~n42704 & n43364 ;
  assign n43366 = n6709 & ~n43365 ;
  assign n43367 = ~n43363 & n43366 ;
  assign n43368 = ~\pi0680  & ~n21525 ;
  assign n43369 = ~n43024 & n43368 ;
  assign n43370 = ~n6761 & n42716 ;
  assign n43371 = ~n43369 & n43370 ;
  assign n43372 = ~n43367 & n43371 ;
  assign n43373 = ~n43360 & n43372 ;
  assign n43374 = \pi0223  & ~\pi0299  ;
  assign n43375 = ~n43373 & n43374 ;
  assign n43376 = ~n43341 & n43375 ;
  assign n43377 = n22232 & n42670 ;
  assign n43378 = ~n21285 & n43377 ;
  assign n43379 = n22232 & n42679 ;
  assign n43380 = n21285 & n43379 ;
  assign n43381 = ~n43378 & ~n43380 ;
  assign n43382 = n42994 & n43381 ;
  assign n43383 = n2165 & n43382 ;
  assign n43384 = ~\pi0223  & ~\pi0299  ;
  assign n43385 = ~n43383 & n43384 ;
  assign n43386 = ~n43376 & ~n43385 ;
  assign n43387 = n43086 & n43096 ;
  assign n43388 = ~\pi0680  & ~n43387 ;
  assign n43389 = ~n43079 & ~n43099 ;
  assign n43390 = ~n21903 & ~n42739 ;
  assign n43391 = ~n20784 & n43390 ;
  assign n43392 = \pi0634  & ~n20784 ;
  assign n43393 = ~n22293 & n43392 ;
  assign n43394 = ~n43391 & ~n43393 ;
  assign n43395 = n43389 & n43394 ;
  assign n43396 = n6709 & ~n43395 ;
  assign n43397 = ~n43388 & ~n43396 ;
  assign n43398 = n22180 & n42762 ;
  assign n43399 = ~n42774 & ~n43398 ;
  assign n43400 = n43356 & ~n43399 ;
  assign n43401 = \pi0633  & ~n21346 ;
  assign n43402 = \pi0634  & n22297 ;
  assign n43403 = ~n43390 & ~n43402 ;
  assign n43404 = ~n43401 & n43403 ;
  assign n43405 = n43353 & n43404 ;
  assign n43406 = n22180 & ~n43345 ;
  assign n43407 = ~n43405 & n43406 ;
  assign n43408 = ~n43400 & ~n43407 ;
  assign n43409 = ~n2165 & n43408 ;
  assign n43410 = n43397 & n43409 ;
  assign n43411 = ~n21368 & ~n43410 ;
  assign n43412 = ~\pi0603  & ~n42743 ;
  assign n43413 = n21586 & ~n43412 ;
  assign n43414 = n21363 & ~n43404 ;
  assign n43415 = n21361 & ~n43330 ;
  assign n43416 = \pi0680  & ~n43415 ;
  assign n43417 = ~n43414 & n43416 ;
  assign n43418 = n43413 & n43417 ;
  assign n43419 = n43050 & n43415 ;
  assign n43420 = n21363 & n43050 ;
  assign n43421 = ~n43404 & n43420 ;
  assign n43422 = ~n43419 & ~n43421 ;
  assign n43423 = n6711 & n43327 ;
  assign n43424 = \pi0603  & \pi0642  ;
  assign n43425 = n6711 & n43424 ;
  assign n43426 = ~n43330 & n43425 ;
  assign n43427 = ~n43423 & ~n43426 ;
  assign n43428 = ~\pi0603  & ~n6711 ;
  assign n43429 = ~n42676 & n43428 ;
  assign n43430 = ~n21586 & ~n43429 ;
  assign n43431 = \pi0680  & ~n43060 ;
  assign n43432 = \pi0680  & ~n43317 ;
  assign n43433 = n43315 & n43432 ;
  assign n43434 = ~n43431 & ~n43433 ;
  assign n43435 = n43430 & ~n43434 ;
  assign n43436 = n43427 & n43435 ;
  assign n43437 = n43422 & n43436 ;
  assign n43438 = ~n43418 & ~n43437 ;
  assign n43439 = ~\pi0680  & ~n42996 ;
  assign n43440 = n43065 & n43439 ;
  assign n43441 = ~n43059 & n43440 ;
  assign n43442 = n6761 & ~n43441 ;
  assign n43443 = n43438 & n43442 ;
  assign n43444 = ~n43376 & ~n43443 ;
  assign n43445 = ~n43411 & n43444 ;
  assign n43446 = ~n43386 & ~n43445 ;
  assign n43447 = n6732 & ~n43339 ;
  assign n43448 = n43326 & n43447 ;
  assign n43449 = ~n6732 & n42716 ;
  assign n43450 = ~n43369 & n43449 ;
  assign n43451 = ~n43367 & n43450 ;
  assign n43452 = \pi0215  & ~n43451 ;
  assign n43453 = \pi0215  & n22180 ;
  assign n43454 = ~n43359 & n43453 ;
  assign n43455 = ~n43452 & ~n43454 ;
  assign n43456 = \pi0299  & ~n43455 ;
  assign n43457 = ~n43448 & n43456 ;
  assign n43458 = n2352 & n43382 ;
  assign n43459 = n21948 & ~n43458 ;
  assign n43460 = ~n43457 & ~n43459 ;
  assign n43461 = ~n2352 & n43408 ;
  assign n43462 = n43397 & n43461 ;
  assign n43463 = ~n21446 & ~n43462 ;
  assign n43464 = n6732 & ~n43441 ;
  assign n43465 = n43438 & n43464 ;
  assign n43466 = ~n43457 & ~n43465 ;
  assign n43467 = ~n43463 & n43466 ;
  assign n43468 = ~n43460 & ~n43467 ;
  assign n43469 = \pi0039  & ~n43468 ;
  assign n43470 = ~n43446 & n43469 ;
  assign n43471 = n43235 & ~n43470 ;
  assign n43472 = n43298 & n43471 ;
  assign n43473 = ~n43236 & ~n43472 ;
  assign n43474 = ~n42851 & ~n43223 ;
  assign n43475 = n43473 & n43474 ;
  assign n43476 = ~n43224 & ~n43475 ;
  assign n43477 = \pi0778  & ~n43476 ;
  assign n43478 = ~n42922 & n43473 ;
  assign n43479 = \pi0625  & n43161 ;
  assign n43480 = \pi0625  & ~n43151 ;
  assign n43481 = ~n43148 & n43480 ;
  assign n43482 = ~n43479 & ~n43481 ;
  assign n43483 = ~\pi1153  & n43482 ;
  assign n43484 = ~n43478 & n43483 ;
  assign n43485 = ~\pi0608  & ~n42920 ;
  assign n43486 = \pi0778  & n43485 ;
  assign n43487 = ~n43484 & n43486 ;
  assign n43488 = ~n43477 & ~n43487 ;
  assign n43489 = \pi0609  & n42934 ;
  assign n43490 = n31812 & ~n43161 ;
  assign n43491 = ~n43152 & n43490 ;
  assign n43492 = ~n32768 & ~n42912 ;
  assign n43493 = ~n42916 & n43492 ;
  assign n43494 = ~n22787 & ~n43493 ;
  assign n43495 = ~n43491 & n43494 ;
  assign n43496 = ~n43489 & ~n43495 ;
  assign n43497 = \pi0778  & ~n43495 ;
  assign n43498 = ~n42928 & n43497 ;
  assign n43499 = ~n43496 & ~n43498 ;
  assign n43500 = \pi0785  & n43499 ;
  assign n43501 = ~\pi0198  & ~\pi0778  ;
  assign n43502 = ~n23622 & ~n43501 ;
  assign n43503 = n43473 & ~n43502 ;
  assign n43504 = ~n43500 & ~n43503 ;
  assign n43505 = n43488 & n43504 ;
  assign n43506 = n26700 & n43505 ;
  assign n43507 = n22788 & ~n43161 ;
  assign n43508 = ~n43152 & n43507 ;
  assign n43509 = ~n22788 & ~n42912 ;
  assign n43510 = ~n42916 & n43509 ;
  assign n43511 = ~\pi0660  & ~n43510 ;
  assign n43512 = ~n43508 & n43511 ;
  assign n43513 = ~n22787 & ~n43512 ;
  assign n43514 = \pi0609  & ~n43499 ;
  assign n43515 = ~n43513 & ~n43514 ;
  assign n43516 = ~\pi0609  & n42934 ;
  assign n43517 = \pi1155  & ~n43516 ;
  assign n43518 = n22722 & ~n42928 ;
  assign n43519 = ~n43517 & ~n43518 ;
  assign n43520 = ~\pi0609  & ~n43519 ;
  assign n43521 = ~n43503 & ~n43519 ;
  assign n43522 = n43488 & n43521 ;
  assign n43523 = ~n43520 & ~n43522 ;
  assign n43524 = n22767 & ~n43161 ;
  assign n43525 = ~n43152 & n43524 ;
  assign n43526 = ~n22767 & ~n42912 ;
  assign n43527 = ~n42916 & n43526 ;
  assign n43528 = \pi0660  & ~n43527 ;
  assign n43529 = ~n43525 & n43528 ;
  assign n43530 = ~n22766 & ~n43529 ;
  assign n43531 = ~n43514 & ~n43530 ;
  assign n43532 = n43523 & n43531 ;
  assign n43533 = ~n43515 & ~n43532 ;
  assign n43534 = \pi0785  & n26700 ;
  assign n43535 = n43533 & n43534 ;
  assign n43536 = ~n43506 & ~n43535 ;
  assign n43537 = ~n43163 & n43166 ;
  assign n43538 = n22155 & ~n42975 ;
  assign n43539 = ~n43537 & n43538 ;
  assign n43540 = ~n22147 & n42934 ;
  assign n43541 = \pi0781  & ~n22147 ;
  assign n43542 = \pi0781  & ~n42912 ;
  assign n43543 = ~n42916 & n43542 ;
  assign n43544 = ~n43541 & ~n43543 ;
  assign n43545 = n23667 & ~n43544 ;
  assign n43546 = ~n43540 & n43545 ;
  assign n43547 = \pi0778  & n43545 ;
  assign n43548 = ~n42928 & n43547 ;
  assign n43549 = ~n43546 & ~n43548 ;
  assign n43550 = ~n43539 & n43549 ;
  assign n43551 = ~n21034 & ~n43550 ;
  assign n43552 = n30780 & ~n42928 ;
  assign n43553 = n23380 & ~n42934 ;
  assign n43554 = ~n23380 & ~n42912 ;
  assign n43555 = ~n42916 & n43554 ;
  assign n43556 = ~n43553 & ~n43555 ;
  assign n43557 = ~n43552 & n43556 ;
  assign n43558 = n23701 & ~n43557 ;
  assign n43559 = n23683 & n42975 ;
  assign n43560 = n23683 & n43166 ;
  assign n43561 = ~n43163 & n43560 ;
  assign n43562 = ~n43559 & ~n43561 ;
  assign n43563 = n21032 & n43170 ;
  assign n43564 = ~n43163 & n43563 ;
  assign n43565 = ~n20876 & ~n42912 ;
  assign n43566 = ~n42916 & n43565 ;
  assign n43567 = ~n24969 & ~n43566 ;
  assign n43568 = \pi0789  & ~n43567 ;
  assign n43569 = ~n43564 & n43568 ;
  assign n43570 = n43562 & n43569 ;
  assign n43571 = ~n21038 & ~n43570 ;
  assign n43572 = ~n43558 & n43571 ;
  assign n43573 = ~n43551 & n43572 ;
  assign n43574 = n43536 & n43573 ;
  assign n43575 = n22160 & ~n42912 ;
  assign n43576 = ~n42916 & n43575 ;
  assign n43577 = n20951 & ~n43576 ;
  assign n43578 = ~n43555 & n43577 ;
  assign n43579 = ~n43553 & n43578 ;
  assign n43580 = ~n43552 & n43579 ;
  assign n43581 = n31306 & ~n42917 ;
  assign n43582 = ~\pi0626  & ~n23423 ;
  assign n43583 = ~\pi0626  & ~n42912 ;
  assign n43584 = ~n42916 & n43583 ;
  assign n43585 = ~n43582 & ~n43584 ;
  assign n43586 = ~n43172 & ~n43585 ;
  assign n43587 = n43169 & n43586 ;
  assign n43588 = \pi0626  & ~n42912 ;
  assign n43589 = ~n42916 & n43588 ;
  assign n43590 = n20882 & ~n43589 ;
  assign n43591 = ~n43587 & n43590 ;
  assign n43592 = ~n43581 & ~n43591 ;
  assign n43593 = ~n43580 & n43592 ;
  assign n43594 = \pi0626  & ~n23423 ;
  assign n43595 = ~n43589 & ~n43594 ;
  assign n43596 = ~n43172 & ~n43595 ;
  assign n43597 = n43169 & n43596 ;
  assign n43598 = n20881 & ~n43584 ;
  assign n43599 = ~n43597 & n43598 ;
  assign n43600 = ~n23856 & ~n43599 ;
  assign n43601 = n43593 & n43600 ;
  assign n43602 = ~n26803 & ~n43601 ;
  assign n43603 = ~n21067 & ~n43602 ;
  assign n43604 = ~n43574 & n43603 ;
  assign n43605 = ~n43214 & ~n43604 ;
  assign n43606 = ~n43195 & ~n43605 ;
  assign n43607 = ~\pi0630  & ~n42973 ;
  assign n43608 = \pi0630  & ~n42944 ;
  assign n43609 = ~n42941 & n43608 ;
  assign n43610 = \pi0792  & n43608 ;
  assign n43611 = ~n42962 & n43610 ;
  assign n43612 = ~n43609 & ~n43611 ;
  assign n43613 = ~n20846 & ~n43210 ;
  assign n43614 = ~n43208 & n43613 ;
  assign n43615 = ~n20846 & ~n20910 ;
  assign n43616 = ~n20910 & ~n42912 ;
  assign n43617 = ~n42916 & n43616 ;
  assign n43618 = ~n43615 & ~n43617 ;
  assign n43619 = ~n43614 & ~n43618 ;
  assign n43620 = ~n24761 & ~n43619 ;
  assign n43621 = n43612 & n43620 ;
  assign n43622 = ~n43607 & n43621 ;
  assign n43623 = ~n29722 & ~n43622 ;
  assign n43624 = ~n43195 & n43623 ;
  assign n43625 = n9948 & ~n43624 ;
  assign n43626 = ~n43606 & n43625 ;
  assign n43627 = ~n42652 & ~n43626 ;
  assign n43628 = \pi0199  & ~n9948 ;
  assign n43629 = \pi0199  & n21768 ;
  assign n43630 = \pi0199  & n21770 ;
  assign n43631 = ~n21734 & n43630 ;
  assign n43632 = ~n43629 & ~n43631 ;
  assign n43633 = ~n23380 & n43632 ;
  assign n43634 = ~\pi0199  & ~n21757 ;
  assign n43635 = n25669 & ~n43634 ;
  assign n43636 = n6861 & n43635 ;
  assign n43637 = ~\pi0199  & ~\pi0299  ;
  assign n43638 = ~n22078 & n43637 ;
  assign n43639 = ~n22085 & n43638 ;
  assign n43640 = ~n22075 & n43639 ;
  assign n43641 = ~\pi0199  & \pi0299  ;
  assign n43642 = ~n22051 & n43641 ;
  assign n43643 = ~n22061 & n43642 ;
  assign n43644 = ~n22048 & n43643 ;
  assign n43645 = \pi0039  & ~n43644 ;
  assign n43646 = ~n43640 & n43645 ;
  assign n43647 = ~n22099 & n43641 ;
  assign n43648 = ~n22686 & n43637 ;
  assign n43649 = ~n43647 & ~n43648 ;
  assign n43650 = \pi0199  & ~n21998 ;
  assign n43651 = ~n22004 & n43650 ;
  assign n43652 = n27217 & n43651 ;
  assign n43653 = n13558 & ~n22013 ;
  assign n43654 = n22011 & n43653 ;
  assign n43655 = ~\pi0039  & ~n43654 ;
  assign n43656 = ~n43652 & n43655 ;
  assign n43657 = n43649 & n43656 ;
  assign n43658 = ~n43646 & ~n43657 ;
  assign n43659 = \pi0199  & ~n21993 ;
  assign n43660 = ~n43657 & n43659 ;
  assign n43661 = ~n43658 & ~n43660 ;
  assign n43662 = n21764 & n43661 ;
  assign n43663 = ~n43636 & ~n43662 ;
  assign n43664 = \pi0199  & ~\pi0637  ;
  assign n43665 = n21768 & n43664 ;
  assign n43666 = n21770 & n43664 ;
  assign n43667 = ~n21734 & n43666 ;
  assign n43668 = ~n43665 & ~n43667 ;
  assign n43669 = \pi0199  & ~n6861 ;
  assign n43670 = n43668 & ~n43669 ;
  assign n43671 = n43663 & n43670 ;
  assign n43672 = ~\pi0637  & n43668 ;
  assign n43673 = ~\pi0778  & ~n43672 ;
  assign n43674 = ~n43671 & n43673 ;
  assign n43675 = n23380 & ~n43674 ;
  assign n43676 = ~n43633 & ~n43675 ;
  assign n43677 = \pi0625  & n43672 ;
  assign n43678 = \pi0625  & n43670 ;
  assign n43679 = n43663 & n43678 ;
  assign n43680 = ~n43677 & ~n43679 ;
  assign n43681 = ~\pi0625  & n43632 ;
  assign n43682 = \pi1153  & ~n43681 ;
  assign n43683 = n43680 & n43682 ;
  assign n43684 = ~\pi0625  & n43672 ;
  assign n43685 = ~\pi0625  & n43670 ;
  assign n43686 = n43663 & n43685 ;
  assign n43687 = ~n43684 & ~n43686 ;
  assign n43688 = \pi0625  & n43632 ;
  assign n43689 = ~\pi1153  & ~n43688 ;
  assign n43690 = n43687 & n43689 ;
  assign n43691 = ~n43683 & ~n43690 ;
  assign n43692 = \pi0778  & ~n43633 ;
  assign n43693 = ~n43691 & n43692 ;
  assign n43694 = ~n43676 & ~n43693 ;
  assign n43695 = n22162 & n43694 ;
  assign n43696 = ~n22162 & n43632 ;
  assign n43697 = ~\pi0792  & ~n43696 ;
  assign n43698 = ~n43695 & n43697 ;
  assign n43699 = ~\pi0647  & ~n43698 ;
  assign n43700 = \pi0647  & n43632 ;
  assign n43701 = n20897 & ~n43700 ;
  assign n43702 = ~n43699 & n43701 ;
  assign n43703 = \pi0628  & n43696 ;
  assign n43704 = n30310 & n43694 ;
  assign n43705 = ~n43703 & ~n43704 ;
  assign n43706 = ~\pi0628  & n43632 ;
  assign n43707 = \pi1156  & ~n43706 ;
  assign n43708 = n43705 & n43707 ;
  assign n43709 = ~\pi0628  & n43696 ;
  assign n43710 = n30317 & n43694 ;
  assign n43711 = ~n43709 & ~n43710 ;
  assign n43712 = \pi0628  & n43632 ;
  assign n43713 = ~\pi1156  & ~n43712 ;
  assign n43714 = n43711 & n43713 ;
  assign n43715 = ~n43708 & ~n43714 ;
  assign n43716 = \pi0792  & n43701 ;
  assign n43717 = ~n43715 & n43716 ;
  assign n43718 = ~n43702 & ~n43717 ;
  assign n43719 = \pi0647  & ~n43698 ;
  assign n43720 = ~\pi0647  & n43632 ;
  assign n43721 = n20849 & ~n43720 ;
  assign n43722 = ~n43719 & n43721 ;
  assign n43723 = \pi0792  & n43721 ;
  assign n43724 = ~n43715 & n43723 ;
  assign n43725 = ~n43722 & ~n43724 ;
  assign n43726 = \pi0199  & ~n20811 ;
  assign n43727 = n21768 & n43726 ;
  assign n43728 = n21770 & n43726 ;
  assign n43729 = ~n21734 & n43728 ;
  assign n43730 = ~n43727 & ~n43729 ;
  assign n43731 = n21776 & n43632 ;
  assign n43732 = n20811 & ~n43731 ;
  assign n43733 = n43730 & ~n43732 ;
  assign n43734 = n6861 & ~n25033 ;
  assign n43735 = ~n25028 & n43734 ;
  assign n43736 = \pi0199  & \pi0617  ;
  assign n43737 = ~n43735 & n43736 ;
  assign n43738 = \pi0199  & ~\pi0617  ;
  assign n43739 = n21768 & n43738 ;
  assign n43740 = n21770 & n43738 ;
  assign n43741 = ~n21734 & n43740 ;
  assign n43742 = ~n43739 & ~n43741 ;
  assign n43743 = ~\pi0199  & \pi0617  ;
  assign n43744 = \pi0603  & \pi0617  ;
  assign n43745 = ~n20783 & n43744 ;
  assign n43746 = n25039 & n43745 ;
  assign n43747 = ~n43743 & ~n43746 ;
  assign n43748 = n25040 & ~n43747 ;
  assign n43749 = ~\pi0038  & ~n43747 ;
  assign n43750 = n25023 & n43749 ;
  assign n43751 = ~n43748 & ~n43750 ;
  assign n43752 = n6861 & ~n43751 ;
  assign n43753 = n43742 & ~n43752 ;
  assign n43754 = ~n43737 & n43753 ;
  assign n43755 = ~n20985 & ~n43754 ;
  assign n43756 = n20985 & ~n43632 ;
  assign n43757 = ~n25588 & ~n43756 ;
  assign n43758 = n43730 & n43757 ;
  assign n43759 = ~n43755 & n43758 ;
  assign n43760 = ~n43733 & ~n43759 ;
  assign n43761 = n23424 & n43760 ;
  assign n43762 = ~n43755 & n43757 ;
  assign n43763 = ~\pi0781  & ~n43731 ;
  assign n43764 = ~n23423 & n43763 ;
  assign n43765 = ~n43762 & n43764 ;
  assign n43766 = n23423 & ~n43632 ;
  assign n43767 = n30376 & ~n43766 ;
  assign n43768 = ~n43765 & n43767 ;
  assign n43769 = ~n43761 & n43768 ;
  assign n43770 = ~n30376 & n43632 ;
  assign n43771 = ~n20910 & ~n43770 ;
  assign n43772 = ~n43769 & n43771 ;
  assign n43773 = n43725 & ~n43772 ;
  assign n43774 = n43718 & n43773 ;
  assign n43775 = \pi0787  & ~n43774 ;
  assign n43776 = \pi0629  & n43713 ;
  assign n43777 = n43711 & n43776 ;
  assign n43778 = n39058 & ~n43706 ;
  assign n43779 = n43705 & n43778 ;
  assign n43780 = n23880 & n24691 ;
  assign n43781 = ~n43632 & n43780 ;
  assign n43782 = ~n43765 & ~n43766 ;
  assign n43783 = ~n43761 & n43782 ;
  assign n43784 = ~n23880 & n24691 ;
  assign n43785 = ~n43783 & n43784 ;
  assign n43786 = ~n43781 & ~n43785 ;
  assign n43787 = ~n43779 & n43786 ;
  assign n43788 = ~n43777 & n43787 ;
  assign n43789 = \pi0792  & ~n43788 ;
  assign n43790 = n22160 & ~n43632 ;
  assign n43791 = ~\pi0641  & n43790 ;
  assign n43792 = n22160 & n43632 ;
  assign n43793 = ~\pi0641  & ~n43792 ;
  assign n43794 = ~n43694 & n43793 ;
  assign n43795 = ~n43791 & ~n43794 ;
  assign n43796 = \pi0199  & \pi0641  ;
  assign n43797 = n21768 & n43796 ;
  assign n43798 = n21770 & n43796 ;
  assign n43799 = ~n21734 & n43798 ;
  assign n43800 = ~n43797 & ~n43799 ;
  assign n43801 = n20777 & n43800 ;
  assign n43802 = n43795 & n43801 ;
  assign n43803 = n30606 & ~n43766 ;
  assign n43804 = ~n43765 & n43803 ;
  assign n43805 = ~n43761 & n43804 ;
  assign n43806 = \pi0199  & ~\pi0641  ;
  assign n43807 = n21768 & n43806 ;
  assign n43808 = n21770 & n43806 ;
  assign n43809 = ~n21734 & n43808 ;
  assign n43810 = ~n43807 & ~n43809 ;
  assign n43811 = n20776 & n43810 ;
  assign n43812 = ~n43805 & ~n43811 ;
  assign n43813 = \pi0641  & ~n43805 ;
  assign n43814 = ~n43812 & ~n43813 ;
  assign n43815 = ~n43694 & ~n43792 ;
  assign n43816 = ~n43790 & ~n43812 ;
  assign n43817 = ~n43815 & n43816 ;
  assign n43818 = ~n43814 & ~n43817 ;
  assign n43819 = ~n43802 & n43818 ;
  assign n43820 = \pi0788  & ~n43819 ;
  assign n43821 = ~n26119 & ~n43691 ;
  assign n43822 = \pi0609  & ~n43756 ;
  assign n43823 = ~n43755 & n43822 ;
  assign n43824 = ~\pi0609  & n43632 ;
  assign n43825 = n20864 & ~n43824 ;
  assign n43826 = ~n43823 & n43825 ;
  assign n43827 = ~\pi0609  & ~n43756 ;
  assign n43828 = ~n43755 & n43827 ;
  assign n43829 = \pi0609  & n43632 ;
  assign n43830 = n20865 & ~n43829 ;
  assign n43831 = ~n43828 & n43830 ;
  assign n43832 = n26125 & ~n43672 ;
  assign n43833 = ~n43671 & n43832 ;
  assign n43834 = ~n43831 & ~n43833 ;
  assign n43835 = ~n43826 & n43834 ;
  assign n43836 = ~n43821 & n43835 ;
  assign n43837 = \pi0785  & ~n43836 ;
  assign n43838 = n21022 & n43837 ;
  assign n43839 = ~\pi0199  & ~n6861 ;
  assign n43840 = ~\pi0199  & ~n25217 ;
  assign n43841 = ~n43839 & ~n43840 ;
  assign n43842 = n31753 & ~n43839 ;
  assign n43843 = n23572 & n43842 ;
  assign n43844 = ~n43841 & ~n43843 ;
  assign n43845 = ~\pi0038  & \pi0199  ;
  assign n43846 = ~n23567 & n43845 ;
  assign n43847 = n23565 & n43846 ;
  assign n43848 = ~\pi0617  & ~n25209 ;
  assign n43849 = ~n43847 & n43848 ;
  assign n43850 = n6861 & ~n43849 ;
  assign n43851 = ~n43844 & ~n43850 ;
  assign n43852 = n6861 & ~n25195 ;
  assign n43853 = \pi0038  & n43852 ;
  assign n43854 = ~n23558 & n43852 ;
  assign n43855 = n23557 & n43854 ;
  assign n43856 = ~n43853 & ~n43855 ;
  assign n43857 = ~\pi0199  & n43856 ;
  assign n43858 = \pi0199  & n23548 ;
  assign n43859 = ~n25191 & n43858 ;
  assign n43860 = ~n25190 & n43859 ;
  assign n43861 = \pi0617  & ~n43860 ;
  assign n43862 = ~n43857 & n43861 ;
  assign n43863 = ~n43851 & ~n43862 ;
  assign n43864 = \pi0625  & \pi0637  ;
  assign n43865 = n43863 & n43864 ;
  assign n43866 = ~n43737 & n43742 ;
  assign n43867 = \pi0625  & ~n43752 ;
  assign n43868 = ~\pi0637  & n43867 ;
  assign n43869 = n43866 & n43868 ;
  assign n43870 = ~\pi0625  & ~n43752 ;
  assign n43871 = n43866 & n43870 ;
  assign n43872 = \pi1153  & ~n43871 ;
  assign n43873 = ~n43869 & n43872 ;
  assign n43874 = ~n43865 & n43873 ;
  assign n43875 = \pi0608  & ~n43690 ;
  assign n43876 = ~n43874 & n43875 ;
  assign n43877 = ~\pi0625  & \pi0637  ;
  assign n43878 = n43863 & n43877 ;
  assign n43879 = ~\pi0625  & ~\pi0637  ;
  assign n43880 = n43754 & n43879 ;
  assign n43881 = n43866 & n43867 ;
  assign n43882 = ~\pi1153  & ~n43881 ;
  assign n43883 = ~n43880 & n43882 ;
  assign n43884 = ~n43878 & n43883 ;
  assign n43885 = ~\pi0608  & ~n43683 ;
  assign n43886 = ~n43884 & n43885 ;
  assign n43887 = ~n43876 & ~n43886 ;
  assign n43888 = \pi0778  & ~n43887 ;
  assign n43889 = \pi0637  & ~\pi0778  ;
  assign n43890 = n43863 & n43889 ;
  assign n43891 = ~\pi0637  & ~\pi0778  ;
  assign n43892 = n43754 & n43891 ;
  assign n43893 = ~n23808 & ~n43892 ;
  assign n43894 = ~n43890 & n43893 ;
  assign n43895 = n21022 & n43894 ;
  assign n43896 = ~n43888 & n43895 ;
  assign n43897 = ~n43838 & ~n43896 ;
  assign n43898 = ~n22147 & ~n43674 ;
  assign n43899 = \pi0781  & n23846 ;
  assign n43900 = n24348 & ~n43632 ;
  assign n43901 = ~n43899 & ~n43900 ;
  assign n43902 = ~n43898 & ~n43901 ;
  assign n43903 = \pi0778  & ~n43901 ;
  assign n43904 = ~n43691 & n43903 ;
  assign n43905 = ~n43902 & ~n43904 ;
  assign n43906 = n22155 & n43760 ;
  assign n43907 = \pi0789  & ~n21030 ;
  assign n43908 = \pi0789  & ~n21032 ;
  assign n43909 = ~n43632 & n43908 ;
  assign n43910 = ~n43907 & ~n43909 ;
  assign n43911 = ~n21038 & n43910 ;
  assign n43912 = ~n43906 & n43911 ;
  assign n43913 = n43905 & n43912 ;
  assign n43914 = n43897 & n43913 ;
  assign n43915 = n23683 & n43760 ;
  assign n43916 = n21032 & n43763 ;
  assign n43917 = ~n43762 & n43916 ;
  assign n43918 = ~n21032 & ~n43632 ;
  assign n43919 = ~n20876 & ~n43918 ;
  assign n43920 = \pi0789  & n43919 ;
  assign n43921 = ~n43917 & n43920 ;
  assign n43922 = ~n43915 & n43921 ;
  assign n43923 = ~n21038 & n43922 ;
  assign n43924 = ~n21038 & ~n31283 ;
  assign n43925 = n43694 & n43924 ;
  assign n43926 = ~n43923 & ~n43925 ;
  assign n43927 = ~n23856 & n43926 ;
  assign n43928 = ~n43914 & n43927 ;
  assign n43929 = ~n43820 & n43928 ;
  assign n43930 = ~n43789 & ~n43929 ;
  assign n43931 = ~n21067 & ~n43930 ;
  assign n43932 = ~n24761 & ~n43931 ;
  assign n43933 = ~n43775 & n43932 ;
  assign n43934 = ~\pi1157  & ~n43700 ;
  assign n43935 = ~n43699 & n43934 ;
  assign n43936 = \pi0792  & n43934 ;
  assign n43937 = ~n43715 & n43936 ;
  assign n43938 = ~n43935 & ~n43937 ;
  assign n43939 = \pi1157  & ~n43720 ;
  assign n43940 = ~n43719 & n43939 ;
  assign n43941 = \pi0792  & n43939 ;
  assign n43942 = ~n43715 & n43941 ;
  assign n43943 = ~n43940 & ~n43942 ;
  assign n43944 = n43938 & n43943 ;
  assign n43945 = n23415 & ~n43770 ;
  assign n43946 = ~n43769 & n43945 ;
  assign n43947 = ~n23415 & ~n43632 ;
  assign n43948 = ~n23414 & ~n43947 ;
  assign n43949 = ~n43946 & n43948 ;
  assign n43950 = \pi0787  & ~n43949 ;
  assign n43951 = ~n43944 & n43950 ;
  assign n43952 = \pi0790  & n43949 ;
  assign n43953 = ~\pi0787  & n43698 ;
  assign n43954 = n33084 & ~n43715 ;
  assign n43955 = ~n43953 & ~n43954 ;
  assign n43956 = \pi0790  & n23518 ;
  assign n43957 = n43955 & n43956 ;
  assign n43958 = ~n43952 & ~n43957 ;
  assign n43959 = ~n43951 & ~n43958 ;
  assign n43960 = n9948 & ~n43959 ;
  assign n43961 = ~n43933 & n43960 ;
  assign n43962 = ~n43628 & ~n43961 ;
  assign n43963 = \pi0200  & ~n9948 ;
  assign n43964 = \pi0200  & n21768 ;
  assign n43965 = \pi0200  & n21770 ;
  assign n43966 = ~n21734 & n43965 ;
  assign n43967 = ~n43964 & ~n43966 ;
  assign n43968 = ~n20811 & ~n43967 ;
  assign n43969 = n21776 & n43967 ;
  assign n43970 = n20811 & ~n43969 ;
  assign n43971 = ~n43968 & ~n43970 ;
  assign n43972 = \pi0200  & \pi0606  ;
  assign n43973 = n1289 & n43972 ;
  assign n43974 = n1287 & n43973 ;
  assign n43975 = ~n25040 & n43974 ;
  assign n43976 = ~n25033 & n43975 ;
  assign n43977 = ~n25028 & n43976 ;
  assign n43978 = \pi0606  & n1289 ;
  assign n43979 = n1287 & n43978 ;
  assign n43980 = ~n43972 & ~n43979 ;
  assign n43981 = ~\pi0200  & ~n25040 ;
  assign n43982 = ~n25024 & n43981 ;
  assign n43983 = ~n43980 & ~n43982 ;
  assign n43984 = ~n43977 & n43983 ;
  assign n43985 = ~n43967 & ~n43977 ;
  assign n43986 = ~n43984 & ~n43985 ;
  assign n43987 = ~n20985 & ~n43986 ;
  assign n43988 = n20985 & ~n43967 ;
  assign n43989 = ~n25588 & ~n43988 ;
  assign n43990 = ~n43968 & n43989 ;
  assign n43991 = ~n43987 & n43990 ;
  assign n43992 = ~n43971 & ~n43991 ;
  assign n43993 = \pi0781  & n43992 ;
  assign n43994 = ~n43987 & n43989 ;
  assign n43995 = ~\pi0781  & ~n43969 ;
  assign n43996 = ~n43994 & n43995 ;
  assign n43997 = n43203 & ~n43996 ;
  assign n43998 = ~n43993 & n43997 ;
  assign n43999 = ~n43203 & n43967 ;
  assign n44000 = n24691 & ~n43999 ;
  assign n44001 = ~n43998 & n44000 ;
  assign n44002 = ~\pi0625  & n43967 ;
  assign n44003 = \pi1153  & ~n44002 ;
  assign n44004 = ~\pi0200  & \pi0643  ;
  assign n44005 = ~n6861 & n44004 ;
  assign n44006 = \pi0200  & ~n21988 ;
  assign n44007 = ~n21987 & n44006 ;
  assign n44008 = \pi0200  & ~\pi0223  ;
  assign n44009 = ~n21928 & n44008 ;
  assign n44010 = n21902 & n44009 ;
  assign n44011 = ~n44007 & ~n44010 ;
  assign n44012 = ~\pi0200  & ~n22085 ;
  assign n44013 = ~n22078 & n44012 ;
  assign n44014 = ~n22075 & n44013 ;
  assign n44015 = ~\pi0299  & ~n44014 ;
  assign n44016 = n44011 & n44015 ;
  assign n44017 = n9627 & n44016 ;
  assign n44018 = ~n21969 & ~n21981 ;
  assign n44019 = ~\pi0215  & ~n21947 ;
  assign n44020 = n21937 & n44019 ;
  assign n44021 = ~n44018 & ~n44020 ;
  assign n44022 = \pi0200  & ~n44021 ;
  assign n44023 = ~\pi0200  & ~n22061 ;
  assign n44024 = ~n22051 & n44023 ;
  assign n44025 = ~n22048 & n44024 ;
  assign n44026 = \pi0299  & ~n44025 ;
  assign n44027 = n9627 & n44026 ;
  assign n44028 = ~n44022 & n44027 ;
  assign n44029 = ~n44017 & ~n44028 ;
  assign n44030 = ~\pi0200  & \pi0299  ;
  assign n44031 = ~n22099 & n44030 ;
  assign n44032 = ~\pi0200  & ~\pi0299  ;
  assign n44033 = ~n22686 & n44032 ;
  assign n44034 = ~n44031 & ~n44033 ;
  assign n44035 = \pi0200  & ~\pi0299  ;
  assign n44036 = ~n22013 & n44035 ;
  assign n44037 = n22011 & n44036 ;
  assign n44038 = ~\pi0039  & ~n44037 ;
  assign n44039 = \pi0200  & ~n21998 ;
  assign n44040 = ~n22004 & n44039 ;
  assign n44041 = n27217 & n44040 ;
  assign n44042 = ~\pi0038  & ~n44041 ;
  assign n44043 = n44038 & n44042 ;
  assign n44044 = n44034 & n44043 ;
  assign n44045 = \pi0643  & n1289 ;
  assign n44046 = n1287 & n44045 ;
  assign n44047 = ~n44004 & ~n44046 ;
  assign n44048 = ~\pi0200  & ~n21757 ;
  assign n44049 = n25669 & ~n44048 ;
  assign n44050 = ~n44047 & ~n44049 ;
  assign n44051 = ~n44044 & n44050 ;
  assign n44052 = n44029 & n44051 ;
  assign n44053 = ~n44005 & ~n44052 ;
  assign n44054 = ~\pi0643  & n43967 ;
  assign n44055 = n44053 & ~n44054 ;
  assign n44056 = \pi0625  & ~n44055 ;
  assign n44057 = n44003 & ~n44056 ;
  assign n44058 = \pi0625  & n43967 ;
  assign n44059 = ~\pi1153  & ~n44058 ;
  assign n44060 = ~\pi0625  & ~n44055 ;
  assign n44061 = n44059 & ~n44060 ;
  assign n44062 = ~n44057 & ~n44061 ;
  assign n44063 = n26065 & ~n44062 ;
  assign n44064 = ~\pi0778  & ~n44005 ;
  assign n44065 = ~n44052 & n44064 ;
  assign n44066 = ~n44054 & n44065 ;
  assign n44067 = n23885 & n44066 ;
  assign n44068 = ~n23885 & ~n43967 ;
  assign n44069 = ~\pi0628  & ~n44068 ;
  assign n44070 = ~n44067 & n44069 ;
  assign n44071 = ~n44063 & n44070 ;
  assign n44072 = \pi0628  & n43967 ;
  assign n44073 = ~\pi1156  & ~n44072 ;
  assign n44074 = \pi0629  & n44073 ;
  assign n44075 = ~n44071 & n44074 ;
  assign n44076 = \pi0628  & ~n44068 ;
  assign n44077 = ~n44067 & n44076 ;
  assign n44078 = ~n44063 & n44077 ;
  assign n44079 = ~\pi0628  & n43967 ;
  assign n44080 = \pi1156  & ~n44079 ;
  assign n44081 = ~\pi0629  & n44080 ;
  assign n44082 = ~n44078 & n44081 ;
  assign n44083 = ~n44075 & ~n44082 ;
  assign n44084 = ~n44001 & n44083 ;
  assign n44085 = n24724 & ~n44084 ;
  assign n44086 = \pi0200  & \pi0626  ;
  assign n44087 = n21768 & n44086 ;
  assign n44088 = n21770 & n44086 ;
  assign n44089 = ~n21734 & n44088 ;
  assign n44090 = ~n44087 & ~n44089 ;
  assign n44091 = n20882 & n44090 ;
  assign n44092 = \pi0200  & ~\pi0626  ;
  assign n44093 = n21768 & n44092 ;
  assign n44094 = n21770 & n44092 ;
  assign n44095 = ~n21734 & n44094 ;
  assign n44096 = ~n44093 & ~n44095 ;
  assign n44097 = ~\pi0626  & n20881 ;
  assign n44098 = n44096 & n44097 ;
  assign n44099 = ~n44091 & ~n44098 ;
  assign n44100 = n23424 & n43992 ;
  assign n44101 = ~n23423 & n43995 ;
  assign n44102 = ~n43994 & n44101 ;
  assign n44103 = n23423 & ~n43967 ;
  assign n44104 = ~n44102 & ~n44103 ;
  assign n44105 = ~n44100 & n44104 ;
  assign n44106 = ~\pi0626  & ~n44098 ;
  assign n44107 = ~n44105 & n44106 ;
  assign n44108 = ~n44099 & ~n44107 ;
  assign n44109 = n20881 & n44096 ;
  assign n44110 = ~n44103 & n44109 ;
  assign n44111 = ~n44102 & n44110 ;
  assign n44112 = ~n44100 & n44111 ;
  assign n44113 = n30780 & ~n44062 ;
  assign n44114 = n23380 & n44066 ;
  assign n44115 = ~n23380 & ~n43967 ;
  assign n44116 = n22160 & ~n43967 ;
  assign n44117 = n20951 & ~n44116 ;
  assign n44118 = ~n44115 & n44117 ;
  assign n44119 = ~n44114 & n44118 ;
  assign n44120 = ~n44113 & n44119 ;
  assign n44121 = n31306 & n43967 ;
  assign n44122 = ~n23856 & ~n44121 ;
  assign n44123 = ~n44120 & n44122 ;
  assign n44124 = ~n44112 & n44123 ;
  assign n44125 = ~n44108 & n44124 ;
  assign n44126 = ~n26803 & ~n44125 ;
  assign n44127 = ~n21067 & ~n44126 ;
  assign n44128 = ~n44085 & ~n44127 ;
  assign n44129 = n22155 & n43992 ;
  assign n44130 = ~n21034 & n44129 ;
  assign n44131 = \pi0778  & ~n44062 ;
  assign n44132 = ~n22147 & ~n44066 ;
  assign n44133 = ~n44131 & n44132 ;
  assign n44134 = n24348 & ~n43967 ;
  assign n44135 = ~n43899 & ~n44134 ;
  assign n44136 = ~n21034 & ~n44135 ;
  assign n44137 = ~n44133 & n44136 ;
  assign n44138 = ~n44130 & ~n44137 ;
  assign n44139 = ~n22117 & ~n22232 ;
  assign n44140 = n44049 & ~n44139 ;
  assign n44141 = \pi0200  & ~n23567 ;
  assign n44142 = n23565 & n44141 ;
  assign n44143 = ~n44140 & n44142 ;
  assign n44144 = n23572 & n31753 ;
  assign n44145 = ~\pi0038  & \pi0200  ;
  assign n44146 = ~n44140 & ~n44145 ;
  assign n44147 = ~n44144 & n44146 ;
  assign n44148 = ~n44143 & ~n44147 ;
  assign n44149 = ~\pi0606  & \pi0643  ;
  assign n44150 = n1289 & n44149 ;
  assign n44151 = n1287 & n44150 ;
  assign n44152 = n44148 & n44151 ;
  assign n44153 = ~\pi0643  & ~n43986 ;
  assign n44154 = \pi0200  & n23548 ;
  assign n44155 = ~n21484 & ~n44034 ;
  assign n44156 = ~n44154 & ~n44155 ;
  assign n44157 = ~\pi0039  & ~n44155 ;
  assign n44158 = ~n22683 & n44157 ;
  assign n44159 = ~n44156 & ~n44158 ;
  assign n44160 = ~\pi0038  & ~\pi0200  ;
  assign n44161 = ~n43150 & ~n44160 ;
  assign n44162 = n44159 & ~n44161 ;
  assign n44163 = ~\pi0200  & n43979 ;
  assign n44164 = ~n25195 & n44163 ;
  assign n44165 = n23555 & n44164 ;
  assign n44166 = ~n23556 & n44165 ;
  assign n44167 = \pi0200  & ~n6861 ;
  assign n44168 = \pi0200  & n43979 ;
  assign n44169 = ~n25188 & n44168 ;
  assign n44170 = ~n44167 & ~n44169 ;
  assign n44171 = ~n44166 & n44170 ;
  assign n44172 = \pi0643  & ~n44171 ;
  assign n44173 = ~n44162 & n44172 ;
  assign n44174 = ~n44153 & ~n44173 ;
  assign n44175 = ~n44152 & n44174 ;
  assign n44176 = ~\pi0625  & n20790 ;
  assign n44177 = \pi0778  & ~n44176 ;
  assign n44178 = ~n44175 & ~n44177 ;
  assign n44179 = ~n20985 & ~n25587 ;
  assign n44180 = ~n43986 & n44179 ;
  assign n44181 = n20985 & ~n25587 ;
  assign n44182 = ~n43967 & n44181 ;
  assign n44183 = n23808 & ~n44182 ;
  assign n44184 = ~n44180 & n44183 ;
  assign n44185 = n44178 & ~n44184 ;
  assign n44186 = n22740 & n43986 ;
  assign n44187 = ~n23781 & ~n44186 ;
  assign n44188 = \pi0608  & \pi0625  ;
  assign n44189 = ~n44152 & n44188 ;
  assign n44190 = n44174 & n44189 ;
  assign n44191 = n44187 & ~n44190 ;
  assign n44192 = ~n44061 & ~n44191 ;
  assign n44193 = n20858 & ~n43986 ;
  assign n44194 = ~\pi0608  & ~n44193 ;
  assign n44195 = ~n44057 & n44194 ;
  assign n44196 = \pi0778  & ~n44195 ;
  assign n44197 = ~n44184 & n44196 ;
  assign n44198 = ~n44192 & n44197 ;
  assign n44199 = ~n44185 & ~n44198 ;
  assign n44200 = \pi0609  & ~n43988 ;
  assign n44201 = ~n43987 & n44200 ;
  assign n44202 = ~\pi0609  & n43967 ;
  assign n44203 = n20864 & ~n44202 ;
  assign n44204 = ~n44201 & n44203 ;
  assign n44205 = ~n26119 & ~n44062 ;
  assign n44206 = ~n26124 & n44066 ;
  assign n44207 = ~\pi0609  & ~n43988 ;
  assign n44208 = ~n43987 & n44207 ;
  assign n44209 = \pi0609  & n43967 ;
  assign n44210 = n20865 & ~n44209 ;
  assign n44211 = ~n44208 & n44210 ;
  assign n44212 = ~n44206 & ~n44211 ;
  assign n44213 = ~n44205 & n44212 ;
  assign n44214 = ~n44204 & n44213 ;
  assign n44215 = \pi0785  & ~n44214 ;
  assign n44216 = n44199 & ~n44215 ;
  assign n44217 = n26700 & ~n44216 ;
  assign n44218 = n44138 & ~n44217 ;
  assign n44219 = ~n44114 & ~n44115 ;
  assign n44220 = ~n44113 & n44219 ;
  assign n44221 = n21050 & ~n44220 ;
  assign n44222 = ~\pi0619  & ~n43996 ;
  assign n44223 = ~n43993 & n44222 ;
  assign n44224 = \pi0619  & n43967 ;
  assign n44225 = n20874 & ~n44224 ;
  assign n44226 = ~n44223 & n44225 ;
  assign n44227 = ~n44221 & ~n44226 ;
  assign n44228 = \pi0619  & ~n43996 ;
  assign n44229 = ~n43993 & n44228 ;
  assign n44230 = ~\pi0619  & n43967 ;
  assign n44231 = n20875 & ~n44230 ;
  assign n44232 = ~n44229 & n44231 ;
  assign n44233 = ~n21038 & ~n44232 ;
  assign n44234 = n44227 & n44233 ;
  assign n44235 = ~n23177 & ~n44234 ;
  assign n44236 = ~n44085 & ~n44235 ;
  assign n44237 = n44218 & n44236 ;
  assign n44238 = ~n44128 & ~n44237 ;
  assign n44239 = ~n24761 & n44238 ;
  assign n44240 = ~n44067 & ~n44068 ;
  assign n44241 = ~n44063 & n44240 ;
  assign n44242 = ~\pi0792  & ~n44241 ;
  assign n44243 = \pi0647  & ~n44242 ;
  assign n44244 = ~\pi0647  & n43967 ;
  assign n44245 = \pi1157  & ~n44244 ;
  assign n44246 = ~n44243 & n44245 ;
  assign n44247 = ~n44078 & n44080 ;
  assign n44248 = ~n44071 & n44073 ;
  assign n44249 = ~n44247 & ~n44248 ;
  assign n44250 = \pi0792  & n44245 ;
  assign n44251 = ~n44249 & n44250 ;
  assign n44252 = ~n44246 & ~n44251 ;
  assign n44253 = n20846 & n43967 ;
  assign n44254 = ~n20910 & ~n44253 ;
  assign n44255 = n20846 & n44254 ;
  assign n44256 = ~n43999 & n44254 ;
  assign n44257 = ~n43998 & n44256 ;
  assign n44258 = ~n44255 & ~n44257 ;
  assign n44259 = ~\pi0630  & n44258 ;
  assign n44260 = n44252 & n44259 ;
  assign n44261 = ~\pi0647  & ~n44242 ;
  assign n44262 = \pi0647  & n43967 ;
  assign n44263 = ~\pi1157  & ~n44262 ;
  assign n44264 = ~n44261 & n44263 ;
  assign n44265 = \pi0792  & n44263 ;
  assign n44266 = ~n44249 & n44265 ;
  assign n44267 = ~n44264 & ~n44266 ;
  assign n44268 = \pi0630  & n44258 ;
  assign n44269 = n44267 & n44268 ;
  assign n44270 = ~n44260 & ~n44269 ;
  assign n44271 = n32298 & n44270 ;
  assign n44272 = \pi0787  & n44267 ;
  assign n44273 = ~n31367 & ~n43967 ;
  assign n44274 = ~\pi0644  & ~n44273 ;
  assign n44275 = \pi0644  & n43967 ;
  assign n44276 = n23413 & ~n44275 ;
  assign n44277 = ~n44274 & n44276 ;
  assign n44278 = n31367 & n44276 ;
  assign n44279 = ~n44105 & n44278 ;
  assign n44280 = ~n44277 & ~n44279 ;
  assign n44281 = \pi0644  & ~n44273 ;
  assign n44282 = ~\pi0644  & n43967 ;
  assign n44283 = n23412 & ~n44282 ;
  assign n44284 = ~n44281 & n44283 ;
  assign n44285 = n31367 & n44283 ;
  assign n44286 = ~n44105 & n44285 ;
  assign n44287 = ~n44284 & ~n44286 ;
  assign n44288 = n44280 & n44287 ;
  assign n44289 = n44252 & n44288 ;
  assign n44290 = n44272 & n44289 ;
  assign n44291 = ~\pi0787  & ~n44242 ;
  assign n44292 = n23518 & ~n44291 ;
  assign n44293 = n37542 & ~n44249 ;
  assign n44294 = ~n44292 & ~n44293 ;
  assign n44295 = n44288 & n44294 ;
  assign n44296 = \pi0790  & ~n44295 ;
  assign n44297 = ~n44290 & n44296 ;
  assign n44298 = ~n44271 & ~n44297 ;
  assign n44299 = ~n44239 & n44298 ;
  assign n44300 = n27408 & ~n44299 ;
  assign n44301 = ~n43963 & ~n44300 ;
  assign n44302 = ~\pi0332  & \pi0468  ;
  assign n44303 = ~n6712 & n44302 ;
  assign n44304 = ~\pi0032  & \pi0070  ;
  assign n44305 = ~\pi0332  & ~n44304 ;
  assign n44306 = \pi0096  & \pi0210  ;
  assign n44307 = ~\pi0332  & n44306 ;
  assign n44308 = ~n44305 & ~n44307 ;
  assign n44309 = ~\pi0070  & ~\pi0841  ;
  assign n44310 = n7147 & n44309 ;
  assign n44311 = ~n6712 & ~n44310 ;
  assign n44312 = ~n44308 & n44311 ;
  assign n44313 = ~n44303 & ~n44312 ;
  assign n44314 = \pi0947  & ~n6712 ;
  assign n44315 = ~n44308 & ~n44310 ;
  assign n44316 = \pi0332  & n44306 ;
  assign n44317 = \pi0947  & ~n44316 ;
  assign n44318 = ~n44315 & n44317 ;
  assign n44319 = ~n44314 & ~n44318 ;
  assign n44320 = n44313 & ~n44319 ;
  assign n44321 = ~\pi0332  & ~n6712 ;
  assign n44322 = ~\pi0947  & ~n44321 ;
  assign n44323 = ~n6706 & ~n44316 ;
  assign n44324 = n6712 & ~n44323 ;
  assign n44325 = n6712 & ~n44310 ;
  assign n44326 = ~n44308 & n44325 ;
  assign n44327 = ~n44324 & ~n44326 ;
  assign n44328 = n44322 & n44327 ;
  assign n44329 = ~n1292 & ~n44328 ;
  assign n44330 = ~n44320 & n44329 ;
  assign n44331 = ~\pi0059  & ~n44330 ;
  assign n44332 = ~\pi0095  & n1329 ;
  assign n44333 = n1261 & n44332 ;
  assign n44334 = n1354 & n44333 ;
  assign n44335 = n1358 & n44334 ;
  assign n44336 = ~\pi0070  & ~n44335 ;
  assign n44337 = \pi0210  & n1714 ;
  assign n44338 = ~n44336 & n44337 ;
  assign n44339 = \pi0210  & ~\pi0332  ;
  assign n44340 = \pi0032  & ~n44309 ;
  assign n44341 = ~\pi0040  & ~\pi0095  ;
  assign n44342 = n1262 & n44341 ;
  assign n44343 = ~n44340 & n44342 ;
  assign n44344 = n1261 & n44343 ;
  assign n44345 = n1354 & n44344 ;
  assign n44346 = n1358 & n44345 ;
  assign n44347 = \pi0032  & n44309 ;
  assign n44348 = n44305 & ~n44347 ;
  assign n44349 = ~n44346 & n44348 ;
  assign n44350 = ~n44339 & ~n44349 ;
  assign n44351 = ~n44338 & ~n44350 ;
  assign n44352 = ~\pi0468  & ~n44351 ;
  assign n44353 = \pi0332  & \pi0468  ;
  assign n44354 = ~n6712 & ~n44353 ;
  assign n44355 = ~n44352 & n44354 ;
  assign n44356 = n44317 & ~n44351 ;
  assign n44357 = ~n44314 & ~n44356 ;
  assign n44358 = ~n44355 & ~n44357 ;
  assign n44359 = ~n6712 & n44322 ;
  assign n44360 = n44322 & n44323 ;
  assign n44361 = ~n44351 & n44360 ;
  assign n44362 = ~n44359 & ~n44361 ;
  assign n44363 = n1291 & n44362 ;
  assign n44364 = ~n44358 & n44363 ;
  assign n44365 = ~n1291 & ~n44328 ;
  assign n44366 = ~n44320 & n44365 ;
  assign n44367 = \pi0055  & ~n44366 ;
  assign n44368 = ~n44364 & n44367 ;
  assign n44369 = n1292 & ~n44368 ;
  assign n44370 = n44331 & ~n44369 ;
  assign n44371 = \pi0070  & n44337 ;
  assign n44372 = n6967 & n44332 ;
  assign n44373 = n1351 & n44372 ;
  assign n44374 = n44337 & n44373 ;
  assign n44375 = ~n1350 & n44374 ;
  assign n44376 = ~n44371 & ~n44375 ;
  assign n44377 = ~\pi0468  & ~n44376 ;
  assign n44378 = n6967 & n44343 ;
  assign n44379 = n1351 & n44378 ;
  assign n44380 = ~n1350 & n44379 ;
  assign n44381 = n44348 & ~n44380 ;
  assign n44382 = ~\pi0468  & ~n44339 ;
  assign n44383 = ~n44381 & n44382 ;
  assign n44384 = ~n44377 & ~n44383 ;
  assign n44385 = \pi0947  & n44354 ;
  assign n44386 = n44384 & n44385 ;
  assign n44387 = \pi0332  & ~n6712 ;
  assign n44388 = ~n44314 & ~n44387 ;
  assign n44389 = \pi0468  & n6712 ;
  assign n44390 = ~\pi0332  & ~\pi0947  ;
  assign n44391 = ~n44389 & n44390 ;
  assign n44392 = ~n44316 & ~n44391 ;
  assign n44393 = ~n44376 & n44392 ;
  assign n44394 = ~n44339 & n44392 ;
  assign n44395 = ~n44381 & n44394 ;
  assign n44396 = ~n44393 & ~n44395 ;
  assign n44397 = n44388 & n44396 ;
  assign n44398 = ~n44386 & ~n44397 ;
  assign n44399 = n2403 & ~n44398 ;
  assign n44400 = n2342 & n8322 ;
  assign n44401 = n44362 & n44400 ;
  assign n44402 = ~n44358 & n44401 ;
  assign n44403 = \pi0299  & ~n44402 ;
  assign n44404 = ~n44399 & n44403 ;
  assign n44405 = \pi0198  & n1714 ;
  assign n44406 = ~n44336 & n44405 ;
  assign n44407 = \pi0198  & ~\pi0332  ;
  assign n44408 = ~n44349 & ~n44407 ;
  assign n44409 = ~n44406 & ~n44408 ;
  assign n44410 = ~\pi0468  & ~n44409 ;
  assign n44411 = \pi0587  & n44354 ;
  assign n44412 = n44400 & n44411 ;
  assign n44413 = ~n44410 & n44412 ;
  assign n44414 = \pi0070  & n44405 ;
  assign n44415 = n44373 & n44405 ;
  assign n44416 = ~n1350 & n44415 ;
  assign n44417 = ~n44414 & ~n44416 ;
  assign n44418 = ~\pi0468  & ~n44417 ;
  assign n44419 = ~\pi0468  & ~n44407 ;
  assign n44420 = ~n44381 & n44419 ;
  assign n44421 = ~n44418 & ~n44420 ;
  assign n44422 = \pi0587  & ~n44353 ;
  assign n44423 = ~n6712 & n44422 ;
  assign n44424 = n2403 & n44423 ;
  assign n44425 = n44421 & n44424 ;
  assign n44426 = ~n44413 & ~n44425 ;
  assign n44427 = ~\pi0332  & ~\pi0587  ;
  assign n44428 = ~n44389 & n44427 ;
  assign n44429 = \pi0096  & \pi0198  ;
  assign n44430 = \pi0332  & n44429 ;
  assign n44431 = ~n44428 & ~n44430 ;
  assign n44432 = ~n44417 & n44431 ;
  assign n44433 = ~n44407 & n44431 ;
  assign n44434 = ~n44381 & n44433 ;
  assign n44435 = ~n44432 & ~n44434 ;
  assign n44436 = \pi0587  & ~n6712 ;
  assign n44437 = ~n44387 & ~n44436 ;
  assign n44438 = n2403 & n44437 ;
  assign n44439 = n44435 & n44438 ;
  assign n44440 = n44400 & n44437 ;
  assign n44441 = ~\pi0299  & ~n44440 ;
  assign n44442 = ~\pi0299  & n44431 ;
  assign n44443 = ~n44409 & n44442 ;
  assign n44444 = ~n44441 & ~n44443 ;
  assign n44445 = ~n44439 & ~n44444 ;
  assign n44446 = n44426 & n44445 ;
  assign n44447 = ~\pi0074  & ~n44446 ;
  assign n44448 = ~n44404 & n44447 ;
  assign n44449 = ~\pi0074  & n2364 ;
  assign n44450 = n2342 & n44449 ;
  assign n44451 = ~\pi0096  & n44304 ;
  assign n44452 = ~\pi0332  & ~n44451 ;
  assign n44453 = ~\pi0198  & n44304 ;
  assign n44454 = n6971 & n44309 ;
  assign n44455 = ~n44453 & ~n44454 ;
  assign n44456 = n44452 & n44455 ;
  assign n44457 = n7343 & ~n44456 ;
  assign n44458 = n44321 & ~n44457 ;
  assign n44459 = ~\pi0299  & ~n7342 ;
  assign n44460 = ~n6712 & n44459 ;
  assign n44461 = ~n44430 & n44459 ;
  assign n44462 = ~n44456 & n44461 ;
  assign n44463 = ~n44460 & ~n44462 ;
  assign n44464 = ~n44458 & ~n44463 ;
  assign n44465 = ~n44450 & ~n44464 ;
  assign n44466 = ~\pi0055  & ~n44465 ;
  assign n44467 = ~\pi0055  & \pi0299  ;
  assign n44468 = n44328 & n44467 ;
  assign n44469 = n44313 & n44467 ;
  assign n44470 = ~n44319 & n44469 ;
  assign n44471 = ~n44468 & ~n44470 ;
  assign n44472 = ~n44466 & n44471 ;
  assign n44473 = n44331 & ~n44472 ;
  assign n44474 = ~n44448 & n44473 ;
  assign n44475 = ~n44370 & ~n44474 ;
  assign n44476 = \pi0057  & n44328 ;
  assign n44477 = \pi0057  & n44313 ;
  assign n44478 = ~n44319 & n44477 ;
  assign n44479 = ~n44476 & ~n44478 ;
  assign n44480 = n1291 & n1293 ;
  assign n44481 = n44362 & n44480 ;
  assign n44482 = ~n44358 & n44481 ;
  assign n44483 = ~n1291 & n1293 ;
  assign n44484 = ~n44328 & n44483 ;
  assign n44485 = ~n44320 & n44484 ;
  assign n44486 = ~n1293 & ~n44328 ;
  assign n44487 = ~n44320 & n44486 ;
  assign n44488 = \pi0059  & ~n44487 ;
  assign n44489 = ~n44485 & n44488 ;
  assign n44490 = ~n44482 & n44489 ;
  assign n44491 = n44479 & ~n44490 ;
  assign n44492 = n44475 & n44491 ;
  assign n44493 = \pi0057  & ~n44328 ;
  assign n44494 = ~n44320 & n44493 ;
  assign n44495 = \pi0233  & \pi0237  ;
  assign n44496 = ~\pi0201  & n44495 ;
  assign n44497 = ~n44494 & n44496 ;
  assign n44498 = ~n44492 & n44497 ;
  assign n44499 = n2511 & ~n7280 ;
  assign n44500 = ~n6735 & n44499 ;
  assign n44501 = n1259 & n44500 ;
  assign n44502 = n1249 & n44501 ;
  assign n44503 = n8410 & n44502 ;
  assign n44504 = \pi0055  & ~\pi0332  ;
  assign n44505 = ~n44503 & n44504 ;
  assign n44506 = n1292 & ~n44505 ;
  assign n44507 = \pi0332  & ~n1292 ;
  assign n44508 = \pi0057  & \pi0332  ;
  assign n44509 = ~\pi0059  & ~n44508 ;
  assign n44510 = ~n44507 & n44509 ;
  assign n44511 = ~n44506 & n44510 ;
  assign n44512 = \pi0332  & ~n13415 ;
  assign n44513 = ~n7315 & n44400 ;
  assign n44514 = n1281 & n44513 ;
  assign n44515 = n1260 & n44514 ;
  assign n44516 = ~n44512 & ~n44515 ;
  assign n44517 = ~\pi0074  & ~n44516 ;
  assign n44518 = ~\pi0468  & ~n7306 ;
  assign n44519 = ~n44389 & ~n44518 ;
  assign n44520 = n1714 & ~n44519 ;
  assign n44521 = n44373 & n44520 ;
  assign n44522 = ~n1350 & n44521 ;
  assign n44523 = ~\pi0332  & ~n44522 ;
  assign n44524 = ~\pi0074  & n2403 ;
  assign n44525 = ~n44523 & n44524 ;
  assign n44526 = ~n44517 & ~n44525 ;
  assign n44527 = \pi0074  & \pi0332  ;
  assign n44528 = ~\pi0055  & ~n44527 ;
  assign n44529 = n44510 & n44528 ;
  assign n44530 = n44526 & n44529 ;
  assign n44531 = ~n44511 & ~n44530 ;
  assign n44532 = \pi0059  & ~\pi0332  ;
  assign n44533 = ~n1292 & n44532 ;
  assign n44534 = \pi0055  & n44532 ;
  assign n44535 = ~n44533 & ~n44534 ;
  assign n44536 = ~\pi0057  & n44535 ;
  assign n44537 = ~n44508 & ~n44536 ;
  assign n44538 = ~n44508 & n44532 ;
  assign n44539 = ~n44503 & n44538 ;
  assign n44540 = ~n44537 & ~n44539 ;
  assign n44541 = ~\pi0201  & ~n44495 ;
  assign n44542 = n44540 & n44541 ;
  assign n44543 = n44531 & n44542 ;
  assign n44544 = n7284 & ~n20516 ;
  assign n44545 = n7343 & n20516 ;
  assign n44546 = ~n44544 & ~n44545 ;
  assign n44547 = ~n20516 & ~n44306 ;
  assign n44548 = n20515 & ~n44429 ;
  assign n44549 = n6848 & n44548 ;
  assign n44550 = n44495 & ~n44549 ;
  assign n44551 = ~n44547 & n44550 ;
  assign n44552 = ~n44546 & n44551 ;
  assign n44553 = \pi0201  & ~n44552 ;
  assign n44554 = ~n44543 & ~n44553 ;
  assign n44555 = ~n44498 & n44554 ;
  assign n44556 = ~\pi0233  & \pi0237  ;
  assign n44557 = ~\pi0202  & n44556 ;
  assign n44558 = ~n44494 & n44557 ;
  assign n44559 = ~n44492 & n44558 ;
  assign n44560 = ~\pi0202  & ~n44556 ;
  assign n44561 = n44540 & n44560 ;
  assign n44562 = n44531 & n44561 ;
  assign n44563 = ~n44547 & ~n44549 ;
  assign n44564 = ~n20516 & n44556 ;
  assign n44565 = n7284 & n44564 ;
  assign n44566 = n20516 & n44556 ;
  assign n44567 = n7343 & n44566 ;
  assign n44568 = ~n44565 & ~n44567 ;
  assign n44569 = n44563 & ~n44568 ;
  assign n44570 = \pi0202  & ~n44569 ;
  assign n44571 = ~n44562 & ~n44570 ;
  assign n44572 = ~n44559 & n44571 ;
  assign n44573 = ~\pi0233  & ~\pi0237  ;
  assign n44574 = ~\pi0203  & n44573 ;
  assign n44575 = ~n44494 & n44574 ;
  assign n44576 = ~n44492 & n44575 ;
  assign n44577 = ~\pi0203  & ~n44573 ;
  assign n44578 = n44540 & n44577 ;
  assign n44579 = n44531 & n44578 ;
  assign n44580 = ~n20516 & n44573 ;
  assign n44581 = n7284 & n44580 ;
  assign n44582 = n20516 & n44573 ;
  assign n44583 = n7343 & n44582 ;
  assign n44584 = ~n44581 & ~n44583 ;
  assign n44585 = n44563 & ~n44584 ;
  assign n44586 = \pi0203  & ~n44585 ;
  assign n44587 = ~n44579 & ~n44586 ;
  assign n44588 = ~n44576 & n44587 ;
  assign n44589 = ~n6860 & ~n20516 ;
  assign n44590 = ~n44547 & ~n44589 ;
  assign n44591 = ~n6888 & n44429 ;
  assign n44592 = ~n6851 & n44591 ;
  assign n44593 = n20516 & ~n44592 ;
  assign n44594 = \pi0204  & n44495 ;
  assign n44595 = ~n44593 & n44594 ;
  assign n44596 = n44590 & n44595 ;
  assign n44597 = ~n6709 & ~n44353 ;
  assign n44598 = ~n44352 & n44597 ;
  assign n44599 = \pi0907  & ~n6709 ;
  assign n44600 = \pi0907  & ~n44316 ;
  assign n44601 = ~n44351 & n44600 ;
  assign n44602 = ~n44599 & ~n44601 ;
  assign n44603 = ~n44598 & ~n44602 ;
  assign n44604 = ~\pi0332  & ~n6709 ;
  assign n44605 = ~\pi0907  & ~n44604 ;
  assign n44606 = ~\pi0662  & \pi0680  ;
  assign n44607 = n6708 & n44606 ;
  assign n44608 = ~\pi0332  & \pi0680  ;
  assign n44609 = ~n44607 & ~n44608 ;
  assign n44610 = n44605 & n44609 ;
  assign n44611 = n44323 & n44605 ;
  assign n44612 = ~n44351 & n44611 ;
  assign n44613 = ~n44610 & ~n44612 ;
  assign n44614 = n44400 & n44613 ;
  assign n44615 = ~n44603 & n44614 ;
  assign n44616 = \pi0299  & ~n44615 ;
  assign n44617 = \pi0332  & ~\pi0907  ;
  assign n44618 = ~n6709 & ~n44617 ;
  assign n44619 = ~\pi0907  & n44618 ;
  assign n44620 = ~n44353 & n44618 ;
  assign n44621 = n44384 & n44620 ;
  assign n44622 = ~n44619 & ~n44621 ;
  assign n44623 = n1287 & n2402 ;
  assign n44624 = ~n44622 & n44623 ;
  assign n44625 = ~n44430 & ~n44456 ;
  assign n44626 = ~\pi0468  & \pi0602  ;
  assign n44627 = \pi0468  & n6709 ;
  assign n44628 = ~n44626 & ~n44627 ;
  assign n44629 = ~\pi0299  & ~n44628 ;
  assign n44630 = n44625 & n44629 ;
  assign n44631 = n6709 & n44429 ;
  assign n44632 = ~\pi0299  & \pi0332  ;
  assign n44633 = ~n44631 & n44632 ;
  assign n44634 = ~n44450 & ~n44633 ;
  assign n44635 = ~n44630 & n44634 ;
  assign n44636 = ~\pi0055  & ~n44635 ;
  assign n44637 = n6709 & ~n44323 ;
  assign n44638 = n6709 & ~n44310 ;
  assign n44639 = ~n44308 & n44638 ;
  assign n44640 = ~n44637 & ~n44639 ;
  assign n44641 = n44605 & n44640 ;
  assign n44642 = n44467 & n44641 ;
  assign n44643 = ~n44315 & n44600 ;
  assign n44644 = ~n44599 & ~n44643 ;
  assign n44645 = ~n6709 & n44302 ;
  assign n44646 = ~n6709 & ~n44310 ;
  assign n44647 = ~n44308 & n44646 ;
  assign n44648 = ~n44645 & ~n44647 ;
  assign n44649 = n44467 & n44648 ;
  assign n44650 = ~n44644 & n44649 ;
  assign n44651 = ~n44642 & ~n44650 ;
  assign n44652 = ~n44636 & n44651 ;
  assign n44653 = ~n6852 & ~n44316 ;
  assign n44654 = ~n44376 & n44653 ;
  assign n44655 = ~n44339 & n44653 ;
  assign n44656 = ~n44381 & n44655 ;
  assign n44657 = ~n44654 & ~n44656 ;
  assign n44658 = ~n6709 & ~n6852 ;
  assign n44659 = n2403 & ~n44658 ;
  assign n44660 = n44657 & n44659 ;
  assign n44661 = ~n44652 & ~n44660 ;
  assign n44662 = ~n44624 & n44661 ;
  assign n44663 = n44616 & n44662 ;
  assign n44664 = n44480 & n44613 ;
  assign n44665 = ~n44603 & n44664 ;
  assign n44666 = ~n44644 & n44648 ;
  assign n44667 = n44483 & ~n44641 ;
  assign n44668 = ~n44666 & n44667 ;
  assign n44669 = ~n1293 & ~n44641 ;
  assign n44670 = ~n44666 & n44669 ;
  assign n44671 = \pi0059  & ~n44670 ;
  assign n44672 = ~n44668 & n44671 ;
  assign n44673 = ~n44665 & n44672 ;
  assign n44674 = n1291 & n44613 ;
  assign n44675 = ~n44603 & n44674 ;
  assign n44676 = ~n1291 & ~n44641 ;
  assign n44677 = ~n44666 & n44676 ;
  assign n44678 = \pi0055  & ~n44677 ;
  assign n44679 = ~n44675 & n44678 ;
  assign n44680 = ~n44673 & ~n44679 ;
  assign n44681 = \pi0074  & ~n44652 ;
  assign n44682 = ~n6888 & ~n44430 ;
  assign n44683 = ~n6851 & n44682 ;
  assign n44684 = ~n44409 & n44683 ;
  assign n44685 = \pi0332  & ~n44631 ;
  assign n44686 = n44400 & ~n44685 ;
  assign n44687 = ~n44684 & n44686 ;
  assign n44688 = ~\pi0299  & ~n44687 ;
  assign n44689 = ~n44417 & n44683 ;
  assign n44690 = ~n44407 & n44683 ;
  assign n44691 = ~n44381 & n44690 ;
  assign n44692 = ~n44689 & ~n44691 ;
  assign n44693 = n2403 & ~n44685 ;
  assign n44694 = n44692 & n44693 ;
  assign n44695 = ~n44652 & ~n44694 ;
  assign n44696 = n44688 & n44695 ;
  assign n44697 = ~n44681 & ~n44696 ;
  assign n44698 = n1292 & n44697 ;
  assign n44699 = n44680 & n44698 ;
  assign n44700 = ~n44663 & n44699 ;
  assign n44701 = ~n1292 & ~n44641 ;
  assign n44702 = ~n44666 & n44701 ;
  assign n44703 = ~\pi0059  & ~n44702 ;
  assign n44704 = ~n44673 & ~n44703 ;
  assign n44705 = ~\pi0057  & n44495 ;
  assign n44706 = ~n44704 & n44705 ;
  assign n44707 = ~n44700 & n44706 ;
  assign n44708 = \pi0057  & n44641 ;
  assign n44709 = \pi0057  & n44648 ;
  assign n44710 = ~n44644 & n44709 ;
  assign n44711 = ~n44708 & ~n44710 ;
  assign n44712 = n44495 & ~n44711 ;
  assign n44713 = n44495 & ~n44593 ;
  assign n44714 = n44590 & n44713 ;
  assign n44715 = \pi0204  & ~n44714 ;
  assign n44716 = n2511 & ~n6852 ;
  assign n44717 = ~n6851 & n44716 ;
  assign n44718 = n1259 & n44717 ;
  assign n44719 = n1249 & n44718 ;
  assign n44720 = n8410 & n44719 ;
  assign n44721 = n44504 & ~n44720 ;
  assign n44722 = n1292 & ~n44721 ;
  assign n44723 = n44510 & ~n44722 ;
  assign n44724 = ~\pi0299  & n44626 ;
  assign n44725 = ~\pi0299  & \pi0468  ;
  assign n44726 = n6709 & n44725 ;
  assign n44727 = ~n44724 & ~n44726 ;
  assign n44728 = \pi0299  & ~n6852 ;
  assign n44729 = ~n6851 & n44728 ;
  assign n44730 = n44727 & ~n44729 ;
  assign n44731 = n1281 & ~n44730 ;
  assign n44732 = n1260 & n44731 ;
  assign n44733 = ~\pi0332  & ~n44732 ;
  assign n44734 = ~\pi0332  & ~n44400 ;
  assign n44735 = ~n44733 & ~n44734 ;
  assign n44736 = \pi0299  & ~\pi0907  ;
  assign n44737 = ~\pi0299  & ~\pi0602  ;
  assign n44738 = ~\pi0468  & ~n44737 ;
  assign n44739 = ~n44736 & n44738 ;
  assign n44740 = ~n44627 & ~n44739 ;
  assign n44741 = n1714 & ~n44740 ;
  assign n44742 = n44373 & n44741 ;
  assign n44743 = ~n1350 & n44742 ;
  assign n44744 = ~n44735 & ~n44743 ;
  assign n44745 = ~n2403 & ~n44400 ;
  assign n44746 = ~\pi0332  & ~n2403 ;
  assign n44747 = ~n44732 & n44746 ;
  assign n44748 = ~n44745 & ~n44747 ;
  assign n44749 = ~\pi0074  & n44748 ;
  assign n44750 = ~n44744 & n44749 ;
  assign n44751 = \pi0332  & ~n44450 ;
  assign n44752 = ~\pi0055  & ~n44751 ;
  assign n44753 = n44510 & n44752 ;
  assign n44754 = ~n44750 & n44753 ;
  assign n44755 = ~n44723 & ~n44754 ;
  assign n44756 = n44538 & ~n44720 ;
  assign n44757 = ~n44537 & ~n44756 ;
  assign n44758 = ~n44495 & n44757 ;
  assign n44759 = n44755 & n44758 ;
  assign n44760 = ~n44715 & ~n44759 ;
  assign n44761 = ~n44712 & n44760 ;
  assign n44762 = ~n44707 & n44761 ;
  assign n44763 = ~n44596 & ~n44762 ;
  assign n44764 = n20516 & n44592 ;
  assign n44765 = ~n20516 & n44306 ;
  assign n44766 = n6860 & n44765 ;
  assign n44767 = ~n44764 & ~n44766 ;
  assign n44768 = \pi0205  & n44556 ;
  assign n44769 = ~n44767 & n44768 ;
  assign n44770 = ~\pi0057  & n44556 ;
  assign n44771 = ~n44704 & n44770 ;
  assign n44772 = ~n44700 & n44771 ;
  assign n44773 = n44556 & ~n44711 ;
  assign n44774 = n44556 & ~n44767 ;
  assign n44775 = \pi0205  & ~n44774 ;
  assign n44776 = ~n44556 & n44757 ;
  assign n44777 = n44755 & n44776 ;
  assign n44778 = ~n44775 & ~n44777 ;
  assign n44779 = ~n44773 & n44778 ;
  assign n44780 = ~n44772 & n44779 ;
  assign n44781 = ~n44769 & ~n44780 ;
  assign n44782 = \pi0233  & ~\pi0237  ;
  assign n44783 = \pi0206  & n44782 ;
  assign n44784 = ~n44767 & n44783 ;
  assign n44785 = ~\pi0057  & n44782 ;
  assign n44786 = ~n44704 & n44785 ;
  assign n44787 = ~n44700 & n44786 ;
  assign n44788 = ~n44711 & n44782 ;
  assign n44789 = ~n44767 & n44782 ;
  assign n44790 = \pi0206  & ~n44789 ;
  assign n44791 = n44757 & ~n44782 ;
  assign n44792 = n44755 & n44791 ;
  assign n44793 = ~n44790 & ~n44792 ;
  assign n44794 = ~n44788 & n44793 ;
  assign n44795 = ~n44787 & n44794 ;
  assign n44796 = ~n44784 & ~n44795 ;
  assign n44797 = n6861 & ~n20811 ;
  assign n44798 = ~n22124 & n44797 ;
  assign n44799 = ~n28084 & n44798 ;
  assign n44800 = n21777 & ~n43735 ;
  assign n44801 = n21768 & ~n21777 ;
  assign n44802 = n21770 & ~n21777 ;
  assign n44803 = ~n21734 & n44802 ;
  assign n44804 = ~n44801 & ~n44803 ;
  assign n44805 = n20811 & n44804 ;
  assign n44806 = ~n44800 & n44805 ;
  assign n44807 = ~n44799 & ~n44806 ;
  assign n44808 = n23424 & ~n44807 ;
  assign n44809 = ~\pi0781  & ~n23423 ;
  assign n44810 = n44804 & n44809 ;
  assign n44811 = ~n44800 & n44810 ;
  assign n44812 = n6861 & ~n21032 ;
  assign n44813 = \pi0789  & n44812 ;
  assign n44814 = ~n22124 & n44813 ;
  assign n44815 = ~n28084 & n44814 ;
  assign n44816 = ~n44811 & ~n44815 ;
  assign n44817 = n30376 & n44816 ;
  assign n44818 = ~n44808 & n44817 ;
  assign n44819 = n21768 & ~n30376 ;
  assign n44820 = n21770 & ~n30376 ;
  assign n44821 = ~n21734 & n44820 ;
  assign n44822 = ~n44819 & ~n44821 ;
  assign n44823 = ~\pi0207  & ~\pi0623  ;
  assign n44824 = n21768 & n44823 ;
  assign n44825 = n21770 & n44823 ;
  assign n44826 = ~n21734 & n44825 ;
  assign n44827 = ~n44824 & ~n44826 ;
  assign n44828 = ~\pi0207  & n44827 ;
  assign n44829 = n44822 & n44828 ;
  assign n44830 = ~n44818 & n44829 ;
  assign n44831 = ~\pi0207  & \pi0623  ;
  assign n44832 = n6861 & ~n20846 ;
  assign n44833 = n25040 & n44832 ;
  assign n44834 = ~\pi0038  & n44832 ;
  assign n44835 = n25023 & n44834 ;
  assign n44836 = ~n44833 & ~n44835 ;
  assign n44837 = n23832 & ~n23880 ;
  assign n44838 = \pi0623  & n44837 ;
  assign n44839 = ~n44836 & n44838 ;
  assign n44840 = ~n44831 & ~n44839 ;
  assign n44841 = n44827 & n44840 ;
  assign n44842 = n23419 & ~n44841 ;
  assign n44843 = ~n44830 & n44842 ;
  assign n44844 = ~\pi0207  & n21768 ;
  assign n44845 = ~\pi0207  & n21770 ;
  assign n44846 = ~n21734 & n44845 ;
  assign n44847 = ~n44844 & ~n44846 ;
  assign n44848 = n23416 & ~n44847 ;
  assign n44849 = \pi0790  & ~n44848 ;
  assign n44850 = ~n44843 & n44849 ;
  assign n44851 = n23074 & n23316 ;
  assign n44852 = n23021 & n23315 ;
  assign n44853 = ~n44851 & ~n44852 ;
  assign n44854 = ~\pi0625  & n21768 ;
  assign n44855 = ~\pi0625  & n21770 ;
  assign n44856 = ~n21734 & n44855 ;
  assign n44857 = ~n44854 & ~n44856 ;
  assign n44858 = \pi1153  & ~n44857 ;
  assign n44859 = n6861 & ~n25669 ;
  assign n44860 = ~n31625 & n44859 ;
  assign n44861 = n24550 & ~n44860 ;
  assign n44862 = ~n44858 & ~n44861 ;
  assign n44863 = \pi0625  & n21768 ;
  assign n44864 = \pi0625  & n21770 ;
  assign n44865 = ~n21734 & n44864 ;
  assign n44866 = ~n44863 & ~n44865 ;
  assign n44867 = ~\pi1153  & ~n44866 ;
  assign n44868 = n24561 & ~n44860 ;
  assign n44869 = ~n44867 & ~n44868 ;
  assign n44870 = n44862 & n44869 ;
  assign n44871 = n22148 & ~n44870 ;
  assign n44872 = n22151 & ~n44860 ;
  assign n44873 = n21768 & n22147 ;
  assign n44874 = n21770 & n22147 ;
  assign n44875 = ~n21734 & n44874 ;
  assign n44876 = ~n44873 & ~n44875 ;
  assign n44877 = n22849 & n44876 ;
  assign n44878 = ~n44872 & n44877 ;
  assign n44879 = ~n44871 & n44878 ;
  assign n44880 = ~n21768 & ~n22849 ;
  assign n44881 = ~n28084 & n44880 ;
  assign n44882 = n33294 & ~n44881 ;
  assign n44883 = ~n44879 & n44882 ;
  assign n44884 = n21768 & ~n33294 ;
  assign n44885 = n21770 & ~n33294 ;
  assign n44886 = ~n21734 & n44885 ;
  assign n44887 = ~n44884 & ~n44886 ;
  assign n44888 = ~\pi0207  & \pi0710  ;
  assign n44889 = n44887 & n44888 ;
  assign n44890 = ~n44883 & n44889 ;
  assign n44891 = ~n20861 & n23380 ;
  assign n44892 = n6861 & n44891 ;
  assign n44893 = ~n22117 & n44892 ;
  assign n44894 = ~n22160 & n33294 ;
  assign n44895 = n44893 & n44894 ;
  assign n44896 = ~n22109 & n44895 ;
  assign n44897 = \pi0207  & \pi0710  ;
  assign n44898 = ~n44896 & n44897 ;
  assign n44899 = ~\pi0710  & n44847 ;
  assign n44900 = n23518 & ~n44899 ;
  assign n44901 = ~n44898 & n44900 ;
  assign n44902 = ~n44890 & n44901 ;
  assign n44903 = n44853 & ~n44902 ;
  assign n44904 = n44850 & n44903 ;
  assign n44905 = ~\pi0647  & ~n44899 ;
  assign n44906 = ~n44898 & n44905 ;
  assign n44907 = ~n44890 & n44906 ;
  assign n44908 = ~\pi0207  & \pi0647  ;
  assign n44909 = n21768 & n44908 ;
  assign n44910 = n21770 & n44908 ;
  assign n44911 = ~n21734 & n44910 ;
  assign n44912 = ~n44909 & ~n44911 ;
  assign n44913 = ~\pi1157  & n44912 ;
  assign n44914 = ~n44907 & n44913 ;
  assign n44915 = \pi0647  & ~n44899 ;
  assign n44916 = ~n44898 & n44915 ;
  assign n44917 = ~n44890 & n44916 ;
  assign n44918 = ~\pi0207  & ~\pi0647  ;
  assign n44919 = n21768 & n44918 ;
  assign n44920 = n21770 & n44918 ;
  assign n44921 = ~n21734 & n44920 ;
  assign n44922 = ~n44919 & ~n44921 ;
  assign n44923 = \pi1157  & n44922 ;
  assign n44924 = ~n44917 & n44923 ;
  assign n44925 = ~n44914 & ~n44924 ;
  assign n44926 = \pi0787  & n44850 ;
  assign n44927 = ~n44925 & n44926 ;
  assign n44928 = ~n44904 & ~n44927 ;
  assign n44929 = ~n23318 & ~n44928 ;
  assign n44930 = ~\pi0710  & ~n44841 ;
  assign n44931 = ~n44830 & n44930 ;
  assign n44932 = ~n21067 & ~n44931 ;
  assign n44933 = \pi0630  & n44913 ;
  assign n44934 = ~n44907 & n44933 ;
  assign n44935 = ~\pi0630  & n44923 ;
  assign n44936 = ~n44917 & n44935 ;
  assign n44937 = ~n44830 & ~n44841 ;
  assign n44938 = ~n20910 & ~n44937 ;
  assign n44939 = ~n44936 & ~n44938 ;
  assign n44940 = ~n44934 & n44939 ;
  assign n44941 = \pi0787  & ~n44940 ;
  assign n44942 = ~n44932 & ~n44941 ;
  assign n44943 = ~n44929 & n44942 ;
  assign n44944 = \pi0626  & ~\pi1158  ;
  assign n44945 = ~\pi0641  & \pi0788  ;
  assign n44946 = n44944 & n44945 ;
  assign n44947 = \pi0641  & \pi0788  ;
  assign n44948 = n20776 & n44947 ;
  assign n44949 = ~n44946 & ~n44948 ;
  assign n44950 = ~n22160 & ~n44949 ;
  assign n44951 = n44893 & n44950 ;
  assign n44952 = ~n22109 & n44951 ;
  assign n44953 = ~n23856 & n44952 ;
  assign n44954 = ~n21038 & ~n23856 ;
  assign n44955 = ~\pi0625  & \pi0778  ;
  assign n44956 = ~n20790 & n44955 ;
  assign n44957 = \pi0625  & \pi0778  ;
  assign n44958 = ~n20788 & n44957 ;
  assign n44959 = ~n44956 & ~n44958 ;
  assign n44960 = n6861 & n44959 ;
  assign n44961 = n25217 & n44960 ;
  assign n44962 = n31753 & n44960 ;
  assign n44963 = n23572 & n44962 ;
  assign n44964 = ~n44961 & ~n44963 ;
  assign n44965 = ~n20858 & ~n30491 ;
  assign n44966 = n20789 & n44965 ;
  assign n44967 = n31631 & n44966 ;
  assign n44968 = ~n22109 & n44967 ;
  assign n44969 = ~n21776 & ~n44968 ;
  assign n44970 = n44964 & n44969 ;
  assign n44971 = ~n20861 & n20866 ;
  assign n44972 = ~n22109 & n44971 ;
  assign n44973 = n31631 & n44972 ;
  assign n44974 = ~n44970 & n44973 ;
  assign n44975 = n44964 & ~n44968 ;
  assign n44976 = ~n23808 & ~n44975 ;
  assign n44977 = ~n44974 & ~n44976 ;
  assign n44978 = n26700 & ~n44977 ;
  assign n44979 = ~n20861 & ~n22147 ;
  assign n44980 = \pi0618  & \pi0781  ;
  assign n44981 = n20869 & n44980 ;
  assign n44982 = ~\pi0618  & \pi0781  ;
  assign n44983 = n20870 & n44982 ;
  assign n44984 = ~n44981 & ~n44983 ;
  assign n44985 = n44979 & ~n44984 ;
  assign n44986 = n31631 & n44985 ;
  assign n44987 = ~n22109 & n44986 ;
  assign n44988 = ~n21034 & n44987 ;
  assign n44989 = ~\pi0648  & \pi0789  ;
  assign n44990 = n21031 & n44989 ;
  assign n44991 = \pi0648  & \pi1159  ;
  assign n44992 = ~\pi0619  & \pi0789  ;
  assign n44993 = n44991 & n44992 ;
  assign n44994 = ~n44990 & ~n44993 ;
  assign n44995 = n44893 & ~n44994 ;
  assign n44996 = ~n22109 & n44995 ;
  assign n44997 = ~n44988 & ~n44996 ;
  assign n44998 = ~n44978 & n44997 ;
  assign n44999 = n44954 & ~n44998 ;
  assign n45000 = ~n44953 & ~n44999 ;
  assign n45001 = n20944 & n22932 ;
  assign n45002 = ~\pi0628  & \pi0792  ;
  assign n45003 = n20844 & n45002 ;
  assign n45004 = ~n45001 & ~n45003 ;
  assign n45005 = n22162 & ~n45004 ;
  assign n45006 = n44893 & n45005 ;
  assign n45007 = ~n22109 & n45006 ;
  assign n45008 = \pi0207  & ~n45007 ;
  assign n45009 = n45000 & n45008 ;
  assign n45010 = ~\pi0623  & ~n45009 ;
  assign n45011 = \pi0710  & ~n44941 ;
  assign n45012 = ~n44929 & n45011 ;
  assign n45013 = n45010 & n45012 ;
  assign n45014 = n21768 & n22155 ;
  assign n45015 = n21770 & n22155 ;
  assign n45016 = ~n21734 & n45015 ;
  assign n45017 = ~n45014 & ~n45016 ;
  assign n45018 = n44876 & n45017 ;
  assign n45019 = ~n44872 & n45018 ;
  assign n45020 = ~n44871 & n45019 ;
  assign n45021 = ~n21768 & n22155 ;
  assign n45022 = ~n28084 & n45021 ;
  assign n45023 = n22162 & ~n45022 ;
  assign n45024 = ~n45020 & n45023 ;
  assign n45025 = n21768 & n22160 ;
  assign n45026 = n21770 & n22160 ;
  assign n45027 = ~n21734 & n45026 ;
  assign n45028 = ~n45025 & ~n45027 ;
  assign n45029 = n21768 & n22161 ;
  assign n45030 = n21770 & n22161 ;
  assign n45031 = ~n21734 & n45030 ;
  assign n45032 = ~n45029 & ~n45031 ;
  assign n45033 = n45028 & n45032 ;
  assign n45034 = ~n45024 & n45033 ;
  assign n45035 = ~n23880 & ~n44816 ;
  assign n45036 = n23424 & ~n23880 ;
  assign n45037 = ~n44807 & n45036 ;
  assign n45038 = ~n45035 & ~n45037 ;
  assign n45039 = n6861 & n23880 ;
  assign n45040 = ~n22124 & n45039 ;
  assign n45041 = ~n28084 & n45040 ;
  assign n45042 = n24691 & ~n45041 ;
  assign n45043 = n45038 & n45042 ;
  assign n45044 = ~\pi0628  & ~n45043 ;
  assign n45045 = n45034 & n45044 ;
  assign n45046 = \pi0628  & n1289 ;
  assign n45047 = n1287 & n45046 ;
  assign n45048 = ~n22124 & n45047 ;
  assign n45049 = ~n28084 & n45048 ;
  assign n45050 = n20844 & ~n45049 ;
  assign n45051 = ~n45043 & ~n45050 ;
  assign n45052 = \pi0792  & ~n45051 ;
  assign n45053 = ~n45045 & n45052 ;
  assign n45054 = ~\pi0628  & n21768 ;
  assign n45055 = ~\pi0628  & n21770 ;
  assign n45056 = ~n21734 & n45055 ;
  assign n45057 = ~n45054 & ~n45056 ;
  assign n45058 = ~\pi0629  & ~n45057 ;
  assign n45059 = n20944 & n45058 ;
  assign n45060 = n45001 & ~n45034 ;
  assign n45061 = ~n45059 & ~n45060 ;
  assign n45062 = ~n45053 & n45061 ;
  assign n45063 = ~\pi0207  & n45062 ;
  assign n45064 = n31631 & n44979 ;
  assign n45065 = ~n22109 & n45064 ;
  assign n45066 = \pi0618  & n20869 ;
  assign n45067 = ~n45065 & n45066 ;
  assign n45068 = n6861 & n25040 ;
  assign n45069 = n21764 & n25023 ;
  assign n45070 = ~n45068 & ~n45069 ;
  assign n45071 = \pi0618  & n21777 ;
  assign n45072 = ~n45070 & n45071 ;
  assign n45073 = n30730 & ~n45072 ;
  assign n45074 = ~n45067 & ~n45073 ;
  assign n45075 = ~n23830 & n25040 ;
  assign n45076 = ~\pi0038  & ~n23830 ;
  assign n45077 = n25023 & n45076 ;
  assign n45078 = ~n45075 & ~n45077 ;
  assign n45079 = \pi0619  & n6861 ;
  assign n45080 = n21777 & n45079 ;
  assign n45081 = ~n45078 & n45080 ;
  assign n45082 = n20875 & n45081 ;
  assign n45083 = ~\pi1159  & n21028 ;
  assign n45084 = n6861 & n45083 ;
  assign n45085 = n21777 & n45084 ;
  assign n45086 = ~n45078 & n45085 ;
  assign n45087 = \pi1159  & n21028 ;
  assign n45088 = n44893 & n45087 ;
  assign n45089 = ~n22109 & n45088 ;
  assign n45090 = ~\pi1159  & n21029 ;
  assign n45091 = n44893 & n45090 ;
  assign n45092 = ~n22109 & n45091 ;
  assign n45093 = ~n45089 & ~n45092 ;
  assign n45094 = ~n45086 & n45093 ;
  assign n45095 = ~n45082 & n45094 ;
  assign n45096 = \pi0789  & ~n45095 ;
  assign n45097 = \pi0781  & ~n45096 ;
  assign n45098 = ~n45074 & n45097 ;
  assign n45099 = ~n25195 & n44960 ;
  assign n45100 = \pi0038  & n45099 ;
  assign n45101 = ~n23558 & n45099 ;
  assign n45102 = n23557 & n45101 ;
  assign n45103 = ~n45100 & ~n45102 ;
  assign n45104 = \pi0609  & n45103 ;
  assign n45105 = ~n20861 & n31631 ;
  assign n45106 = ~n22109 & n45105 ;
  assign n45107 = ~\pi0609  & ~n45106 ;
  assign n45108 = \pi1155  & ~n45107 ;
  assign n45109 = ~n45104 & n45108 ;
  assign n45110 = n22755 & n31631 ;
  assign n45111 = ~n22109 & n45110 ;
  assign n45112 = \pi1153  & ~n45111 ;
  assign n45113 = n1289 & n22740 ;
  assign n45114 = n1287 & n45113 ;
  assign n45115 = n25040 & n45114 ;
  assign n45116 = ~\pi0038  & n45114 ;
  assign n45117 = n25023 & n45116 ;
  assign n45118 = ~n45115 & ~n45117 ;
  assign n45119 = n45112 & n45118 ;
  assign n45120 = \pi0778  & ~n45119 ;
  assign n45121 = n22740 & n31631 ;
  assign n45122 = ~n22109 & n45121 ;
  assign n45123 = ~\pi1153  & ~n45122 ;
  assign n45124 = n1289 & n22755 ;
  assign n45125 = n1287 & n45124 ;
  assign n45126 = n25040 & n45125 ;
  assign n45127 = ~\pi0038  & n45125 ;
  assign n45128 = n25023 & n45127 ;
  assign n45129 = ~n45126 & ~n45128 ;
  assign n45130 = n45123 & n45129 ;
  assign n45131 = n45108 & ~n45130 ;
  assign n45132 = n45120 & n45131 ;
  assign n45133 = ~n45109 & ~n45132 ;
  assign n45134 = n1289 & n20999 ;
  assign n45135 = n1287 & n45134 ;
  assign n45136 = ~n20985 & n45135 ;
  assign n45137 = n25040 & n45136 ;
  assign n45138 = ~\pi0038  & n45136 ;
  assign n45139 = n25023 & n45138 ;
  assign n45140 = ~n45137 & ~n45139 ;
  assign n45141 = \pi0660  & n45140 ;
  assign n45142 = n45133 & n45141 ;
  assign n45143 = n22816 & n45142 ;
  assign n45144 = ~\pi0609  & n45103 ;
  assign n45145 = \pi0609  & ~n45106 ;
  assign n45146 = ~n45144 & ~n45145 ;
  assign n45147 = ~n45130 & ~n45145 ;
  assign n45148 = n45120 & n45147 ;
  assign n45149 = ~n45146 & ~n45148 ;
  assign n45150 = ~\pi1155  & ~n45149 ;
  assign n45151 = n1289 & n21774 ;
  assign n45152 = n1287 & n45151 ;
  assign n45153 = ~n20985 & n45152 ;
  assign n45154 = n25040 & n45153 ;
  assign n45155 = ~\pi0038  & n45153 ;
  assign n45156 = n25023 & n45155 ;
  assign n45157 = ~n45154 & ~n45156 ;
  assign n45158 = ~\pi0660  & n45157 ;
  assign n45159 = n22816 & n45158 ;
  assign n45160 = ~n45150 & n45159 ;
  assign n45161 = ~n45143 & ~n45160 ;
  assign n45162 = n45120 & ~n45130 ;
  assign n45163 = ~\pi0785  & n45103 ;
  assign n45164 = \pi0618  & n45163 ;
  assign n45165 = ~n45162 & n45164 ;
  assign n45166 = ~\pi0618  & ~n45065 ;
  assign n45167 = \pi1154  & ~n45166 ;
  assign n45168 = ~n45165 & n45167 ;
  assign n45169 = n45161 & n45168 ;
  assign n45170 = n21777 & n25612 ;
  assign n45171 = ~n45070 & n45170 ;
  assign n45172 = \pi0627  & ~n45171 ;
  assign n45173 = n45097 & n45172 ;
  assign n45174 = ~n45169 & n45173 ;
  assign n45175 = ~n45098 & ~n45174 ;
  assign n45176 = \pi0785  & ~n33630 ;
  assign n45177 = n45142 & n45176 ;
  assign n45178 = n45158 & n45176 ;
  assign n45179 = ~n45150 & n45178 ;
  assign n45180 = ~n45177 & ~n45179 ;
  assign n45181 = ~n33630 & n45163 ;
  assign n45182 = ~n45162 & n45181 ;
  assign n45183 = ~n21034 & ~n45182 ;
  assign n45184 = n45180 & n45183 ;
  assign n45185 = ~n45096 & ~n45184 ;
  assign n45186 = n44954 & ~n45185 ;
  assign n45187 = n45175 & n45186 ;
  assign n45188 = n23832 & n25040 ;
  assign n45189 = ~\pi0038  & n23832 ;
  assign n45190 = n25023 & n45189 ;
  assign n45191 = ~n45188 & ~n45190 ;
  assign n45192 = n1289 & n20948 ;
  assign n45193 = n1287 & n45192 ;
  assign n45194 = ~n45191 & n45193 ;
  assign n45195 = n20949 & ~n22160 ;
  assign n45196 = n44893 & n45195 ;
  assign n45197 = ~n22109 & n45196 ;
  assign n45198 = ~\pi1158  & ~n45197 ;
  assign n45199 = ~n45194 & n45198 ;
  assign n45200 = \pi0788  & ~n45199 ;
  assign n45201 = n1289 & n20949 ;
  assign n45202 = n1287 & n45201 ;
  assign n45203 = ~n45191 & n45202 ;
  assign n45204 = n20948 & ~n22160 ;
  assign n45205 = n44893 & n45204 ;
  assign n45206 = ~n22109 & n45205 ;
  assign n45207 = \pi1158  & ~n45206 ;
  assign n45208 = ~n45203 & n45207 ;
  assign n45209 = ~n23856 & ~n45208 ;
  assign n45210 = n45200 & n45209 ;
  assign n45211 = ~n22160 & n22932 ;
  assign n45212 = n44893 & n45211 ;
  assign n45213 = ~n22109 & n45212 ;
  assign n45214 = ~n22161 & n45213 ;
  assign n45215 = n6861 & n22166 ;
  assign n45216 = ~n23880 & n45215 ;
  assign n45217 = n23832 & n45216 ;
  assign n45218 = n25040 & n45217 ;
  assign n45219 = ~\pi0038  & n45217 ;
  assign n45220 = n25023 & n45219 ;
  assign n45221 = ~n45218 & ~n45220 ;
  assign n45222 = \pi1156  & n45221 ;
  assign n45223 = ~n45214 & n45222 ;
  assign n45224 = ~n22160 & n22166 ;
  assign n45225 = n44893 & n45224 ;
  assign n45226 = ~n22109 & n45225 ;
  assign n45227 = ~n22161 & n45226 ;
  assign n45228 = n6861 & n22932 ;
  assign n45229 = ~n23880 & n45228 ;
  assign n45230 = n23832 & n45229 ;
  assign n45231 = n25040 & n45230 ;
  assign n45232 = ~\pi0038  & n45230 ;
  assign n45233 = n25023 & n45232 ;
  assign n45234 = ~n45231 & ~n45233 ;
  assign n45235 = ~\pi1156  & n45234 ;
  assign n45236 = ~n45227 & n45235 ;
  assign n45237 = ~n45223 & ~n45236 ;
  assign n45238 = \pi0792  & n45237 ;
  assign n45239 = \pi0207  & ~n45238 ;
  assign n45240 = ~n45210 & n45239 ;
  assign n45241 = ~n45187 & n45240 ;
  assign n45242 = ~n45063 & ~n45241 ;
  assign n45243 = ~n31283 & ~n45022 ;
  assign n45244 = ~n45020 & n45243 ;
  assign n45245 = ~n22124 & n44812 ;
  assign n45246 = ~n28084 & n45245 ;
  assign n45247 = ~n20876 & ~n45246 ;
  assign n45248 = ~n23683 & n45247 ;
  assign n45249 = ~n44799 & n45247 ;
  assign n45250 = ~n44806 & n45249 ;
  assign n45251 = ~n45248 & ~n45250 ;
  assign n45252 = ~\pi0781  & n21032 ;
  assign n45253 = n44804 & n45252 ;
  assign n45254 = ~n44800 & n45253 ;
  assign n45255 = \pi0789  & ~n45254 ;
  assign n45256 = ~n45251 & n45255 ;
  assign n45257 = ~n21038 & ~n45256 ;
  assign n45258 = ~n45244 & n45257 ;
  assign n45259 = ~\pi0641  & ~n44881 ;
  assign n45260 = ~n44879 & n45259 ;
  assign n45261 = \pi0641  & n21768 ;
  assign n45262 = \pi0641  & n21770 ;
  assign n45263 = ~n21734 & n45262 ;
  assign n45264 = ~n45261 & ~n45263 ;
  assign n45265 = n44944 & n45264 ;
  assign n45266 = ~n45260 & n45265 ;
  assign n45267 = \pi0788  & n45266 ;
  assign n45268 = ~n44879 & ~n44881 ;
  assign n45269 = n30606 & ~n44816 ;
  assign n45270 = n23424 & n30606 ;
  assign n45271 = ~n44807 & n45270 ;
  assign n45272 = ~n45269 & ~n45271 ;
  assign n45273 = \pi0641  & n45272 ;
  assign n45274 = n45268 & n45273 ;
  assign n45275 = ~\pi0641  & n21768 ;
  assign n45276 = ~\pi0641  & n21770 ;
  assign n45277 = ~n21734 & n45276 ;
  assign n45278 = ~n45275 & ~n45277 ;
  assign n45279 = n20776 & n45278 ;
  assign n45280 = n45272 & ~n45279 ;
  assign n45281 = \pi0788  & ~n45280 ;
  assign n45282 = ~n45274 & n45281 ;
  assign n45283 = ~n45267 & ~n45282 ;
  assign n45284 = ~n45258 & n45283 ;
  assign n45285 = ~n44872 & n44876 ;
  assign n45286 = n20871 & ~n44799 ;
  assign n45287 = ~n44806 & n45286 ;
  assign n45288 = n45285 & ~n45287 ;
  assign n45289 = ~n44871 & n45288 ;
  assign n45290 = ~n23667 & ~n45287 ;
  assign n45291 = \pi0781  & ~n45290 ;
  assign n45292 = ~n45289 & n45291 ;
  assign n45293 = n6861 & ~n25191 ;
  assign n45294 = n23548 & n45293 ;
  assign n45295 = ~n25190 & n45294 ;
  assign n45296 = ~\pi0778  & ~n45295 ;
  assign n45297 = ~\pi0785  & ~n45296 ;
  assign n45298 = n21022 & ~n45297 ;
  assign n45299 = n22727 & ~n25191 ;
  assign n45300 = n23548 & n45299 ;
  assign n45301 = ~n25190 & n45300 ;
  assign n45302 = n22734 & ~n25033 ;
  assign n45303 = ~n25028 & n45302 ;
  assign n45304 = ~n45301 & ~n45303 ;
  assign n45305 = \pi1153  & n45304 ;
  assign n45306 = \pi0608  & ~n45305 ;
  assign n45307 = n44869 & n45306 ;
  assign n45308 = \pi0778  & ~n45307 ;
  assign n45309 = n22734 & ~n25191 ;
  assign n45310 = n23548 & n45309 ;
  assign n45311 = ~n25190 & n45310 ;
  assign n45312 = n22727 & ~n25033 ;
  assign n45313 = ~n25028 & n45312 ;
  assign n45314 = ~n45311 & ~n45313 ;
  assign n45315 = ~\pi1153  & n45314 ;
  assign n45316 = ~\pi0608  & ~n45315 ;
  assign n45317 = n44862 & n45316 ;
  assign n45318 = n21022 & ~n45317 ;
  assign n45319 = n45308 & n45318 ;
  assign n45320 = ~n45298 & ~n45319 ;
  assign n45321 = ~n45292 & n45320 ;
  assign n45322 = \pi0609  & n45296 ;
  assign n45323 = \pi0609  & ~n45317 ;
  assign n45324 = n45308 & n45323 ;
  assign n45325 = ~n45322 & ~n45324 ;
  assign n45326 = n23613 & ~n44870 ;
  assign n45327 = ~\pi0609  & ~\pi0778  ;
  assign n45328 = ~n44860 & n45327 ;
  assign n45329 = n31812 & ~n43735 ;
  assign n45330 = n21768 & ~n32768 ;
  assign n45331 = n21770 & ~n32768 ;
  assign n45332 = ~n21734 & n45331 ;
  assign n45333 = ~n45330 & ~n45332 ;
  assign n45334 = \pi0660  & n45333 ;
  assign n45335 = ~n45329 & n45334 ;
  assign n45336 = ~n45328 & n45335 ;
  assign n45337 = ~n45326 & n45336 ;
  assign n45338 = n45325 & n45337 ;
  assign n45339 = n22767 & ~n43735 ;
  assign n45340 = n20865 & n45333 ;
  assign n45341 = ~n45339 & n45340 ;
  assign n45342 = \pi1155  & n22788 ;
  assign n45343 = ~n43735 & n45342 ;
  assign n45344 = n21768 & ~n32759 ;
  assign n45345 = n21770 & ~n32759 ;
  assign n45346 = ~n21734 & n45345 ;
  assign n45347 = ~n45344 & ~n45346 ;
  assign n45348 = ~\pi0660  & n45347 ;
  assign n45349 = ~n45343 & n45348 ;
  assign n45350 = ~n45341 & ~n45349 ;
  assign n45351 = ~n45338 & n45350 ;
  assign n45352 = ~\pi1155  & n21768 ;
  assign n45353 = ~\pi1155  & n21770 ;
  assign n45354 = ~n21734 & n45353 ;
  assign n45355 = ~n45352 & ~n45354 ;
  assign n45356 = ~n22767 & ~n45355 ;
  assign n45357 = ~n45329 & ~n45356 ;
  assign n45358 = n31121 & n45357 ;
  assign n45359 = ~\pi0609  & ~n45317 ;
  assign n45360 = n45308 & n45359 ;
  assign n45361 = ~n45295 & n45327 ;
  assign n45362 = n23638 & ~n44870 ;
  assign n45363 = \pi0609  & ~\pi0778  ;
  assign n45364 = ~n44860 & n45363 ;
  assign n45365 = \pi0785  & ~n45364 ;
  assign n45366 = ~n45362 & n45365 ;
  assign n45367 = ~n45361 & n45366 ;
  assign n45368 = ~n45360 & n45367 ;
  assign n45369 = ~n45358 & ~n45368 ;
  assign n45370 = ~n45292 & ~n45369 ;
  assign n45371 = ~n45351 & n45370 ;
  assign n45372 = ~n45321 & ~n45371 ;
  assign n45373 = ~n21034 & n45283 ;
  assign n45374 = n45372 & n45373 ;
  assign n45375 = ~n45284 & ~n45374 ;
  assign n45376 = ~n23856 & ~n45241 ;
  assign n45377 = ~n45375 & n45376 ;
  assign n45378 = ~n45242 & ~n45377 ;
  assign n45379 = \pi0623  & n45012 ;
  assign n45380 = ~n45378 & n45379 ;
  assign n45381 = ~n45013 & ~n45380 ;
  assign n45382 = ~n44943 & n45381 ;
  assign n45383 = ~\pi0628  & n45032 ;
  assign n45384 = n45028 & n45383 ;
  assign n45385 = ~n45024 & n45384 ;
  assign n45386 = ~n20844 & ~n20887 ;
  assign n45387 = ~n45049 & ~n45386 ;
  assign n45388 = \pi0792  & n45387 ;
  assign n45389 = ~n45385 & n45388 ;
  assign n45390 = n45033 & n45057 ;
  assign n45391 = ~n45024 & n45390 ;
  assign n45392 = ~n22932 & n45057 ;
  assign n45393 = n20944 & ~n45392 ;
  assign n45394 = ~n45391 & n45393 ;
  assign n45395 = ~n45389 & ~n45394 ;
  assign n45396 = ~\pi0625  & ~n25209 ;
  assign n45397 = ~n25204 & n45396 ;
  assign n45398 = ~\pi0625  & ~n6861 ;
  assign n45399 = n44866 & ~n45398 ;
  assign n45400 = ~n45397 & n45399 ;
  assign n45401 = ~\pi1153  & ~n45400 ;
  assign n45402 = ~\pi0608  & n44862 ;
  assign n45403 = ~n45401 & n45402 ;
  assign n45404 = \pi0778  & ~n45403 ;
  assign n45405 = \pi0625  & ~n25209 ;
  assign n45406 = ~n25204 & n45405 ;
  assign n45407 = \pi0625  & ~n6861 ;
  assign n45408 = n44857 & ~n45407 ;
  assign n45409 = ~n45406 & n45408 ;
  assign n45410 = \pi1153  & ~n45409 ;
  assign n45411 = \pi0608  & n44869 ;
  assign n45412 = ~n45410 & n45411 ;
  assign n45413 = n45404 & ~n45412 ;
  assign n45414 = ~\pi0778  & ~n6861 ;
  assign n45415 = ~\pi0778  & ~n25209 ;
  assign n45416 = ~n25204 & n45415 ;
  assign n45417 = ~n45414 & ~n45416 ;
  assign n45418 = ~\pi0785  & n45417 ;
  assign n45419 = ~n45413 & n45418 ;
  assign n45420 = ~\pi0785  & ~n45419 ;
  assign n45421 = ~\pi0609  & ~n45417 ;
  assign n45422 = ~\pi0609  & ~n45412 ;
  assign n45423 = n45404 & n45422 ;
  assign n45424 = ~n45421 & ~n45423 ;
  assign n45425 = \pi1155  & n21768 ;
  assign n45426 = \pi1155  & n21770 ;
  assign n45427 = ~n21734 & n45426 ;
  assign n45428 = ~n45425 & ~n45427 ;
  assign n45429 = ~\pi0660  & n45428 ;
  assign n45430 = ~n45362 & ~n45364 ;
  assign n45431 = n45429 & n45430 ;
  assign n45432 = n45424 & n45431 ;
  assign n45433 = n20864 & ~n21768 ;
  assign n45434 = ~n28084 & n45433 ;
  assign n45435 = n20865 & ~n21768 ;
  assign n45436 = ~n28084 & n45435 ;
  assign n45437 = ~n45434 & ~n45436 ;
  assign n45438 = ~n45432 & n45437 ;
  assign n45439 = \pi0609  & ~n45417 ;
  assign n45440 = \pi0609  & ~n45412 ;
  assign n45441 = n45404 & n45440 ;
  assign n45442 = ~n45439 & ~n45441 ;
  assign n45443 = ~n45326 & ~n45328 ;
  assign n45444 = \pi0660  & n45355 ;
  assign n45445 = n45443 & n45444 ;
  assign n45446 = n45442 & n45445 ;
  assign n45447 = ~n45419 & ~n45446 ;
  assign n45448 = n45438 & n45447 ;
  assign n45449 = ~n45420 & ~n45448 ;
  assign n45450 = n20869 & ~n45449 ;
  assign n45451 = ~\pi0618  & ~n20870 ;
  assign n45452 = ~\pi0618  & n44876 ;
  assign n45453 = ~n44872 & n45452 ;
  assign n45454 = ~n44871 & n45453 ;
  assign n45455 = ~n45451 & ~n45454 ;
  assign n45456 = ~n45450 & ~n45455 ;
  assign n45457 = n20870 & ~n45419 ;
  assign n45458 = ~\pi0785  & n45457 ;
  assign n45459 = ~n45446 & n45457 ;
  assign n45460 = n45438 & n45459 ;
  assign n45461 = ~n45458 & ~n45460 ;
  assign n45462 = \pi0618  & ~n20869 ;
  assign n45463 = \pi0618  & n44876 ;
  assign n45464 = ~n44872 & n45463 ;
  assign n45465 = ~n44871 & n45464 ;
  assign n45466 = ~n45462 & ~n45465 ;
  assign n45467 = n45461 & ~n45466 ;
  assign n45468 = \pi0781  & ~n45467 ;
  assign n45469 = ~n45456 & n45468 ;
  assign n45470 = ~\pi0781  & ~n45449 ;
  assign n45471 = \pi0619  & n45017 ;
  assign n45472 = ~n45470 & n45471 ;
  assign n45473 = ~n45469 & n45472 ;
  assign n45474 = ~n45020 & ~n45022 ;
  assign n45475 = ~\pi0619  & ~n45474 ;
  assign n45476 = n44991 & ~n45475 ;
  assign n45477 = ~n45473 & n45476 ;
  assign n45478 = ~n20876 & n21768 ;
  assign n45479 = ~n20876 & n21770 ;
  assign n45480 = ~n21734 & n45479 ;
  assign n45481 = ~n45478 & ~n45480 ;
  assign n45482 = \pi0789  & n45481 ;
  assign n45483 = ~n45477 & n45482 ;
  assign n45484 = ~\pi0619  & n45017 ;
  assign n45485 = ~n45470 & n45484 ;
  assign n45486 = ~n45469 & n45485 ;
  assign n45487 = ~\pi0648  & ~\pi1159  ;
  assign n45488 = \pi0619  & ~n45474 ;
  assign n45489 = n45487 & ~n45488 ;
  assign n45490 = ~n45486 & n45489 ;
  assign n45491 = ~\pi0788  & ~n45490 ;
  assign n45492 = n45483 & n45491 ;
  assign n45493 = ~\pi0789  & n45017 ;
  assign n45494 = ~n45470 & n45493 ;
  assign n45495 = ~\pi0788  & n45494 ;
  assign n45496 = ~n45469 & n45495 ;
  assign n45497 = ~n23856 & ~n45496 ;
  assign n45498 = ~n45492 & n45497 ;
  assign n45499 = n45395 & ~n45498 ;
  assign n45500 = ~\pi1158  & n45264 ;
  assign n45501 = ~\pi0626  & ~n45490 ;
  assign n45502 = n45483 & n45501 ;
  assign n45503 = ~\pi0626  & n45494 ;
  assign n45504 = ~n45469 & n45503 ;
  assign n45505 = ~n23719 & ~n45260 ;
  assign n45506 = ~n45504 & ~n45505 ;
  assign n45507 = ~n45502 & n45506 ;
  assign n45508 = n45500 & ~n45507 ;
  assign n45509 = \pi1158  & n45278 ;
  assign n45510 = \pi0626  & ~n45490 ;
  assign n45511 = n45483 & n45510 ;
  assign n45512 = \pi0626  & n45494 ;
  assign n45513 = ~n45469 & n45512 ;
  assign n45514 = \pi0641  & ~n44881 ;
  assign n45515 = ~n44879 & n45514 ;
  assign n45516 = ~n23733 & ~n45515 ;
  assign n45517 = ~n45513 & ~n45516 ;
  assign n45518 = ~n45511 & n45517 ;
  assign n45519 = n45509 & ~n45518 ;
  assign n45520 = ~n45508 & ~n45519 ;
  assign n45521 = \pi0788  & n45395 ;
  assign n45522 = ~n45520 & n45521 ;
  assign n45523 = ~n45499 & ~n45522 ;
  assign n45524 = \pi0623  & ~n45378 ;
  assign n45525 = ~\pi0207  & ~n45524 ;
  assign n45526 = ~n44943 & n45525 ;
  assign n45527 = ~n45523 & n45526 ;
  assign n45528 = ~n45382 & ~n45527 ;
  assign n45529 = \pi0790  & n44928 ;
  assign n45530 = n27408 & ~n45529 ;
  assign n45531 = ~n45528 & n45530 ;
  assign n45532 = \pi0207  & ~n27408 ;
  assign n45533 = ~n45531 & ~n45532 ;
  assign n45534 = ~\pi0208  & ~\pi0607  ;
  assign n45535 = n21768 & n45534 ;
  assign n45536 = n21770 & n45534 ;
  assign n45537 = ~n21734 & n45536 ;
  assign n45538 = ~n45535 & ~n45537 ;
  assign n45539 = ~\pi0208  & n45538 ;
  assign n45540 = n44822 & n45539 ;
  assign n45541 = ~n44818 & n45540 ;
  assign n45542 = ~\pi0208  & \pi0607  ;
  assign n45543 = \pi0607  & n44837 ;
  assign n45544 = ~n44836 & n45543 ;
  assign n45545 = ~n45542 & ~n45544 ;
  assign n45546 = n45538 & n45545 ;
  assign n45547 = n23419 & ~n45546 ;
  assign n45548 = ~n45541 & n45547 ;
  assign n45549 = ~\pi0208  & n21768 ;
  assign n45550 = ~\pi0208  & n21770 ;
  assign n45551 = ~n21734 & n45550 ;
  assign n45552 = ~n45549 & ~n45551 ;
  assign n45553 = n23416 & ~n45552 ;
  assign n45554 = \pi0790  & ~n45553 ;
  assign n45555 = ~n45548 & n45554 ;
  assign n45556 = ~\pi0208  & \pi0638  ;
  assign n45557 = n44887 & n45556 ;
  assign n45558 = ~n44883 & n45557 ;
  assign n45559 = \pi0208  & \pi0638  ;
  assign n45560 = ~n44896 & n45559 ;
  assign n45561 = ~\pi0638  & n45552 ;
  assign n45562 = n23518 & ~n45561 ;
  assign n45563 = ~n45560 & n45562 ;
  assign n45564 = ~n45558 & n45563 ;
  assign n45565 = n44853 & ~n45564 ;
  assign n45566 = n45555 & n45565 ;
  assign n45567 = ~\pi0647  & ~n45560 ;
  assign n45568 = ~n45561 & n45567 ;
  assign n45569 = ~n45558 & n45568 ;
  assign n45570 = ~\pi0208  & \pi0647  ;
  assign n45571 = n21768 & n45570 ;
  assign n45572 = n21770 & n45570 ;
  assign n45573 = ~n21734 & n45572 ;
  assign n45574 = ~n45571 & ~n45573 ;
  assign n45575 = ~\pi1157  & n45574 ;
  assign n45576 = ~n45569 & n45575 ;
  assign n45577 = \pi0647  & ~n45560 ;
  assign n45578 = ~n45561 & n45577 ;
  assign n45579 = ~n45558 & n45578 ;
  assign n45580 = ~\pi0208  & ~\pi0647  ;
  assign n45581 = n21768 & n45580 ;
  assign n45582 = n21770 & n45580 ;
  assign n45583 = ~n21734 & n45582 ;
  assign n45584 = ~n45581 & ~n45583 ;
  assign n45585 = \pi1157  & n45584 ;
  assign n45586 = ~n45579 & n45585 ;
  assign n45587 = ~n45576 & ~n45586 ;
  assign n45588 = \pi0787  & n45555 ;
  assign n45589 = ~n45587 & n45588 ;
  assign n45590 = ~n45566 & ~n45589 ;
  assign n45591 = ~n23318 & ~n45590 ;
  assign n45592 = n20897 & n45574 ;
  assign n45593 = ~n45569 & n45592 ;
  assign n45594 = n20849 & n45584 ;
  assign n45595 = ~n45579 & n45594 ;
  assign n45596 = ~n45541 & ~n45546 ;
  assign n45597 = ~n20910 & ~n45596 ;
  assign n45598 = ~n45595 & ~n45597 ;
  assign n45599 = ~n45593 & n45598 ;
  assign n45600 = \pi0787  & ~n45599 ;
  assign n45601 = ~n45591 & ~n45600 ;
  assign n45602 = \pi0790  & n45590 ;
  assign n45603 = ~n45601 & ~n45602 ;
  assign n45604 = ~n23856 & ~n45375 ;
  assign n45605 = ~\pi0208  & n45062 ;
  assign n45606 = ~n45604 & n45605 ;
  assign n45607 = \pi0208  & ~n45238 ;
  assign n45608 = ~n45210 & n45607 ;
  assign n45609 = ~n45187 & n45608 ;
  assign n45610 = \pi0607  & ~n45609 ;
  assign n45611 = ~n45606 & n45610 ;
  assign n45612 = ~\pi0208  & ~n45611 ;
  assign n45613 = ~n45523 & n45612 ;
  assign n45614 = \pi0208  & ~n45007 ;
  assign n45615 = n45000 & n45614 ;
  assign n45616 = ~\pi0607  & ~n45615 ;
  assign n45617 = ~n45610 & ~n45616 ;
  assign n45618 = n45605 & ~n45616 ;
  assign n45619 = ~n45604 & n45618 ;
  assign n45620 = ~n45617 & ~n45619 ;
  assign n45621 = \pi0638  & n45620 ;
  assign n45622 = ~n45613 & n45621 ;
  assign n45623 = ~\pi0638  & ~n45546 ;
  assign n45624 = ~n45541 & n45623 ;
  assign n45625 = ~n21067 & ~n45624 ;
  assign n45626 = ~n45602 & n45625 ;
  assign n45627 = ~n45622 & n45626 ;
  assign n45628 = ~n45603 & ~n45627 ;
  assign n45629 = n27408 & ~n45628 ;
  assign n45630 = \pi0208  & ~n27408 ;
  assign n45631 = ~n45629 & ~n45630 ;
  assign n45632 = ~n21067 & n23318 ;
  assign n45633 = ~n45062 & n45632 ;
  assign n45634 = ~n23856 & n45632 ;
  assign n45635 = ~n45375 & n45634 ;
  assign n45636 = ~n45633 & ~n45635 ;
  assign n45637 = ~n44883 & n44887 ;
  assign n45638 = ~\pi0647  & n20910 ;
  assign n45639 = ~\pi0647  & n44822 ;
  assign n45640 = ~n44818 & n45639 ;
  assign n45641 = ~n45638 & ~n45640 ;
  assign n45642 = n45637 & ~n45641 ;
  assign n45643 = \pi0647  & n1289 ;
  assign n45644 = n1287 & n45643 ;
  assign n45645 = ~n22124 & n45644 ;
  assign n45646 = ~n28084 & n45645 ;
  assign n45647 = n20897 & ~n45646 ;
  assign n45648 = n20910 & ~n45647 ;
  assign n45649 = n44822 & ~n45647 ;
  assign n45650 = ~n44818 & n45649 ;
  assign n45651 = ~n45648 & ~n45650 ;
  assign n45652 = \pi0787  & n45651 ;
  assign n45653 = ~n45642 & n45652 ;
  assign n45654 = ~\pi0647  & n21768 ;
  assign n45655 = ~\pi0647  & n21770 ;
  assign n45656 = ~n21734 & n45655 ;
  assign n45657 = ~n45654 & ~n45656 ;
  assign n45658 = ~\pi0630  & ~n45657 ;
  assign n45659 = ~n20908 & ~n45658 ;
  assign n45660 = n44887 & ~n45658 ;
  assign n45661 = ~n44883 & n45660 ;
  assign n45662 = ~n45659 & ~n45661 ;
  assign n45663 = n24994 & n45662 ;
  assign n45664 = ~n45653 & ~n45663 ;
  assign n45665 = n23318 & ~n45664 ;
  assign n45666 = ~n21088 & ~n43173 ;
  assign n45667 = ~n21768 & ~n28084 ;
  assign n45668 = ~n45666 & ~n45667 ;
  assign n45669 = ~n45666 & ~n45668 ;
  assign n45670 = n44822 & ~n45668 ;
  assign n45671 = ~n44818 & n45670 ;
  assign n45672 = ~n45669 & ~n45671 ;
  assign n45673 = n23317 & n45672 ;
  assign n45674 = n21768 & n23942 ;
  assign n45675 = n21770 & n23942 ;
  assign n45676 = ~n21734 & n45675 ;
  assign n45677 = ~n45674 & ~n45676 ;
  assign n45678 = n23518 & ~n45677 ;
  assign n45679 = ~n45673 & ~n45678 ;
  assign n45680 = n26068 & ~n45637 ;
  assign n45681 = n45679 & ~n45680 ;
  assign n45682 = ~n45665 & n45681 ;
  assign n45683 = n45636 & n45682 ;
  assign n45684 = \pi0790  & ~n45683 ;
  assign n45685 = ~\pi0790  & ~n21067 ;
  assign n45686 = ~n45062 & n45685 ;
  assign n45687 = ~n23856 & n45685 ;
  assign n45688 = ~n45375 & n45687 ;
  assign n45689 = ~n45686 & ~n45688 ;
  assign n45690 = ~\pi0790  & ~n45664 ;
  assign n45691 = n9948 & ~n45690 ;
  assign n45692 = n45689 & n45691 ;
  assign n45693 = \pi0639  & n45692 ;
  assign n45694 = ~n45684 & n45693 ;
  assign n45695 = \pi0790  & n45672 ;
  assign n45696 = ~\pi0790  & ~n21088 ;
  assign n45697 = n21088 & n21768 ;
  assign n45698 = n21088 & n21770 ;
  assign n45699 = ~n21734 & n45698 ;
  assign n45700 = ~n45697 & ~n45699 ;
  assign n45701 = ~\pi0790  & ~n45700 ;
  assign n45702 = n9948 & ~n45701 ;
  assign n45703 = ~n45696 & n45702 ;
  assign n45704 = n44822 & n45702 ;
  assign n45705 = ~n44818 & n45704 ;
  assign n45706 = ~n45703 & ~n45705 ;
  assign n45707 = ~\pi0639  & ~n45706 ;
  assign n45708 = ~n45695 & n45707 ;
  assign n45709 = ~\pi0209  & \pi0622  ;
  assign n45710 = ~n45708 & n45709 ;
  assign n45711 = ~n45694 & n45710 ;
  assign n45712 = ~\pi0639  & n1289 ;
  assign n45713 = n1287 & n45712 ;
  assign n45714 = n9948 & n45713 ;
  assign n45715 = ~n22124 & n45714 ;
  assign n45716 = ~n28084 & n45715 ;
  assign n45717 = ~\pi0209  & ~\pi0622  ;
  assign n45718 = ~n45716 & n45717 ;
  assign n45719 = ~n45711 & ~n45718 ;
  assign n45720 = ~\pi0647  & n44887 ;
  assign n45721 = ~n44883 & n45720 ;
  assign n45722 = ~n20897 & ~n21064 ;
  assign n45723 = ~n45646 & ~n45722 ;
  assign n45724 = \pi0787  & n45723 ;
  assign n45725 = ~n45721 & n45724 ;
  assign n45726 = n44887 & n45657 ;
  assign n45727 = ~n44883 & n45726 ;
  assign n45728 = ~n20908 & n45657 ;
  assign n45729 = n24994 & ~n45728 ;
  assign n45730 = ~n45727 & n45729 ;
  assign n45731 = ~n45725 & ~n45730 ;
  assign n45732 = n23315 & n45731 ;
  assign n45733 = n23316 & n45677 ;
  assign n45734 = n23942 & n45733 ;
  assign n45735 = n44887 & n45733 ;
  assign n45736 = ~n44883 & n45735 ;
  assign n45737 = ~n45734 & ~n45736 ;
  assign n45738 = ~n45732 & n45737 ;
  assign n45739 = ~n21067 & n45737 ;
  assign n45740 = n45523 & n45739 ;
  assign n45741 = ~n45738 & ~n45740 ;
  assign n45742 = n6861 & n23317 ;
  assign n45743 = ~n22124 & n45742 ;
  assign n45744 = ~n28084 & n45743 ;
  assign n45745 = \pi0790  & ~n45744 ;
  assign n45746 = \pi0644  & n45745 ;
  assign n45747 = ~n45741 & n45746 ;
  assign n45748 = n23316 & n45731 ;
  assign n45749 = n23315 & n45677 ;
  assign n45750 = n23942 & n45749 ;
  assign n45751 = n44887 & n45749 ;
  assign n45752 = ~n44883 & n45751 ;
  assign n45753 = ~n45750 & ~n45752 ;
  assign n45754 = ~n45748 & n45753 ;
  assign n45755 = ~n21067 & n45753 ;
  assign n45756 = n45523 & n45755 ;
  assign n45757 = ~n45754 & ~n45756 ;
  assign n45758 = ~\pi0644  & n45745 ;
  assign n45759 = ~n45757 & n45758 ;
  assign n45760 = ~n45747 & ~n45759 ;
  assign n45761 = n45523 & n45685 ;
  assign n45762 = ~\pi0790  & ~n45731 ;
  assign n45763 = n9948 & ~n45762 ;
  assign n45764 = \pi0639  & n45763 ;
  assign n45765 = ~n45761 & n45764 ;
  assign n45766 = ~n45711 & n45765 ;
  assign n45767 = n45760 & n45766 ;
  assign n45768 = ~n45719 & ~n45767 ;
  assign n45769 = n20906 & n44837 ;
  assign n45770 = ~n44836 & n45769 ;
  assign n45771 = n20908 & n44894 ;
  assign n45772 = n44893 & n45771 ;
  assign n45773 = ~n22109 & n45772 ;
  assign n45774 = \pi1157  & ~n45773 ;
  assign n45775 = ~n45770 & n45774 ;
  assign n45776 = n20908 & n44837 ;
  assign n45777 = ~n44836 & n45776 ;
  assign n45778 = n20906 & n44894 ;
  assign n45779 = n44893 & n45778 ;
  assign n45780 = ~n22109 & n45779 ;
  assign n45781 = ~\pi1157  & ~n45780 ;
  assign n45782 = ~n45777 & n45781 ;
  assign n45783 = ~n45775 & ~n45782 ;
  assign n45784 = \pi0787  & n45783 ;
  assign n45785 = ~n45238 & ~n45784 ;
  assign n45786 = ~n45210 & n45785 ;
  assign n45787 = ~n45187 & n45786 ;
  assign n45788 = \pi0787  & ~n21066 ;
  assign n45789 = ~n45783 & n45788 ;
  assign n45790 = n9948 & ~n24761 ;
  assign n45791 = ~n45789 & n45790 ;
  assign n45792 = ~n45787 & n45791 ;
  assign n45793 = \pi0622  & \pi0639  ;
  assign n45794 = ~\pi1160  & ~n23942 ;
  assign n45795 = n44894 & n45794 ;
  assign n45796 = n44893 & n45795 ;
  assign n45797 = ~n22109 & n45796 ;
  assign n45798 = n30987 & n44837 ;
  assign n45799 = ~n44836 & n45798 ;
  assign n45800 = ~n45797 & ~n45799 ;
  assign n45801 = n23312 & ~n45800 ;
  assign n45802 = \pi1160  & ~n23942 ;
  assign n45803 = n44894 & n45802 ;
  assign n45804 = n44893 & n45803 ;
  assign n45805 = ~n22109 & n45804 ;
  assign n45806 = n31010 & n44837 ;
  assign n45807 = ~n44836 & n45806 ;
  assign n45808 = ~n45805 & ~n45807 ;
  assign n45809 = n23313 & ~n45808 ;
  assign n45810 = ~n45801 & ~n45809 ;
  assign n45811 = \pi0790  & n9948 ;
  assign n45812 = ~n45810 & n45811 ;
  assign n45813 = n45793 & ~n45812 ;
  assign n45814 = ~n45792 & n45813 ;
  assign n45815 = \pi0790  & n44894 ;
  assign n45816 = n44893 & n45815 ;
  assign n45817 = ~n22109 & n45816 ;
  assign n45818 = n26068 & n45817 ;
  assign n45819 = ~\pi0057  & \pi0639  ;
  assign n45820 = n6848 & n45819 ;
  assign n45821 = n45818 & n45820 ;
  assign n45822 = n30823 & n44952 ;
  assign n45823 = ~n21038 & n30823 ;
  assign n45824 = ~n44998 & n45823 ;
  assign n45825 = ~n45822 & ~n45824 ;
  assign n45826 = ~n21067 & n45007 ;
  assign n45827 = \pi0787  & ~\pi1157  ;
  assign n45828 = n20906 & n45827 ;
  assign n45829 = ~\pi0630  & \pi0787  ;
  assign n45830 = n20925 & n45829 ;
  assign n45831 = ~n45828 & ~n45830 ;
  assign n45832 = n44894 & ~n45831 ;
  assign n45833 = n44893 & n45832 ;
  assign n45834 = ~n22109 & n45833 ;
  assign n45835 = ~n45826 & ~n45834 ;
  assign n45836 = n45825 & n45835 ;
  assign n45837 = ~n24761 & n45820 ;
  assign n45838 = ~n45836 & n45837 ;
  assign n45839 = ~n45821 & ~n45838 ;
  assign n45840 = n6861 & n23832 ;
  assign n45841 = \pi0790  & n43173 ;
  assign n45842 = ~n23880 & ~n45841 ;
  assign n45843 = n21092 & n45842 ;
  assign n45844 = n9948 & n45843 ;
  assign n45845 = n45840 & n45844 ;
  assign n45846 = n25040 & n45845 ;
  assign n45847 = ~\pi0038  & n45845 ;
  assign n45848 = n25023 & n45847 ;
  assign n45849 = ~n45846 & ~n45848 ;
  assign n45850 = \pi0622  & ~n45849 ;
  assign n45851 = ~n45793 & ~n45850 ;
  assign n45852 = n45839 & n45851 ;
  assign n45853 = \pi0209  & ~n45852 ;
  assign n45854 = ~n45814 & n45853 ;
  assign n45855 = ~n45768 & ~n45854 ;
  assign n45856 = \pi0634  & n26930 ;
  assign n45857 = \pi0633  & \pi0947  ;
  assign n45858 = ~n45856 & ~n45857 ;
  assign n45859 = ~n21740 & ~n45858 ;
  assign n45860 = ~n21738 & n45859 ;
  assign n45861 = ~\pi0210  & ~\pi0299  ;
  assign n45862 = ~n27218 & ~n45861 ;
  assign n45863 = n21737 & ~n45861 ;
  assign n45864 = n21232 & n45863 ;
  assign n45865 = ~n45862 & ~n45864 ;
  assign n45866 = ~n45860 & n45865 ;
  assign n45867 = ~n21205 & ~n45858 ;
  assign n45868 = \pi0299  & ~n45867 ;
  assign n45869 = ~n21238 & n45868 ;
  assign n45870 = ~\pi0039  & ~n45869 ;
  assign n45871 = ~n45866 & n45870 ;
  assign n45872 = \pi0210  & n21334 ;
  assign n45873 = ~n21330 & n45872 ;
  assign n45874 = ~\pi0634  & ~n6709 ;
  assign n45875 = n6735 & n45874 ;
  assign n45876 = \pi0907  & ~n45875 ;
  assign n45877 = ~n21285 & n45876 ;
  assign n45878 = ~\pi0210  & ~n6709 ;
  assign n45879 = n6735 & n45878 ;
  assign n45880 = \pi0907  & ~n45879 ;
  assign n45881 = n21285 & n45880 ;
  assign n45882 = ~n45877 & ~n45881 ;
  assign n45883 = \pi0210  & ~n21306 ;
  assign n45884 = ~n21903 & n45883 ;
  assign n45885 = \pi0634  & ~n21290 ;
  assign n45886 = ~n21325 & n45885 ;
  assign n45887 = \pi0634  & n21291 ;
  assign n45888 = ~n21305 & n45887 ;
  assign n45889 = ~n6736 & ~n45888 ;
  assign n45890 = ~n45886 & n45889 ;
  assign n45891 = ~n45884 & n45890 ;
  assign n45892 = ~n45882 & ~n45891 ;
  assign n45893 = ~n21694 & ~n45892 ;
  assign n45894 = ~n45873 & n45893 ;
  assign n45895 = n2352 & ~n45857 ;
  assign n45896 = ~n45856 & n45895 ;
  assign n45897 = ~\pi0215  & ~n45896 ;
  assign n45898 = ~n21285 & n45897 ;
  assign n45899 = ~\pi0210  & n2352 ;
  assign n45900 = ~\pi0215  & ~n45899 ;
  assign n45901 = n21285 & n45900 ;
  assign n45902 = ~n45898 & ~n45901 ;
  assign n45903 = ~\pi0947  & ~n45902 ;
  assign n45904 = n45892 & n45903 ;
  assign n45905 = \pi0210  & n6713 ;
  assign n45906 = n21285 & n45905 ;
  assign n45907 = \pi0210  & ~n6713 ;
  assign n45908 = ~n45906 & ~n45907 ;
  assign n45909 = n21694 & n45908 ;
  assign n45910 = n21355 & ~n45906 ;
  assign n45911 = ~n21290 & ~n45906 ;
  assign n45912 = ~n21325 & n45911 ;
  assign n45913 = ~n45910 & ~n45912 ;
  assign n45914 = ~n21352 & n21694 ;
  assign n45915 = ~n45913 & n45914 ;
  assign n45916 = ~n45909 & ~n45915 ;
  assign n45917 = ~\pi0907  & n45903 ;
  assign n45918 = n45916 & n45917 ;
  assign n45919 = ~n45904 & ~n45918 ;
  assign n45920 = ~n45894 & ~n45919 ;
  assign n45921 = \pi0633  & ~n21290 ;
  assign n45922 = ~n21325 & n45921 ;
  assign n45923 = \pi0633  & n21291 ;
  assign n45924 = ~n21305 & n45923 ;
  assign n45925 = ~n2352 & ~n6736 ;
  assign n45926 = ~n45924 & n45925 ;
  assign n45927 = ~n45922 & n45926 ;
  assign n45928 = ~n45884 & n45927 ;
  assign n45929 = ~\pi0633  & ~n6709 ;
  assign n45930 = n6735 & n45929 ;
  assign n45931 = \pi0947  & ~n45930 ;
  assign n45932 = ~n21285 & n45931 ;
  assign n45933 = \pi0947  & ~n45879 ;
  assign n45934 = n21285 & n45933 ;
  assign n45935 = ~n45932 & ~n45934 ;
  assign n45936 = ~n2352 & n45935 ;
  assign n45937 = ~n45902 & ~n45936 ;
  assign n45938 = ~n45928 & n45937 ;
  assign n45939 = ~n6706 & n45907 ;
  assign n45940 = n21403 & n45939 ;
  assign n45941 = ~n21399 & n45940 ;
  assign n45942 = n6706 & n45907 ;
  assign n45943 = n21285 & n45942 ;
  assign n45944 = n21694 & ~n45906 ;
  assign n45945 = ~n45943 & n45944 ;
  assign n45946 = ~n45941 & n45945 ;
  assign n45947 = ~\pi0907  & n21694 ;
  assign n45948 = ~\pi0120  & ~n6709 ;
  assign n45949 = n6735 & n45948 ;
  assign n45950 = n21277 & n45949 ;
  assign n45951 = n1281 & n45950 ;
  assign n45952 = n1260 & n45951 ;
  assign n45953 = \pi0120  & ~n6709 ;
  assign n45954 = n6735 & n45953 ;
  assign n45955 = n1281 & n45954 ;
  assign n45956 = n1260 & n45955 ;
  assign n45957 = ~n45952 & ~n45956 ;
  assign n45958 = n1689 & ~n45957 ;
  assign n45959 = \pi0210  & ~n45958 ;
  assign n45960 = ~\pi0907  & n45959 ;
  assign n45961 = n22183 & n45960 ;
  assign n45962 = ~n45947 & ~n45961 ;
  assign n45963 = ~n45946 & ~n45962 ;
  assign n45964 = ~\pi0633  & ~n6736 ;
  assign n45965 = ~n21403 & n45964 ;
  assign n45966 = ~n21393 & n45964 ;
  assign n45967 = n21398 & n45966 ;
  assign n45968 = ~n45965 & ~n45967 ;
  assign n45969 = ~\pi0210  & ~n6736 ;
  assign n45970 = n21403 & n45969 ;
  assign n45971 = ~n21399 & n45970 ;
  assign n45972 = ~n45935 & ~n45971 ;
  assign n45973 = n45968 & n45972 ;
  assign n45974 = ~\pi0634  & ~n6736 ;
  assign n45975 = ~n21403 & n45974 ;
  assign n45976 = ~n21393 & n45974 ;
  assign n45977 = n21398 & n45976 ;
  assign n45978 = ~n45975 & ~n45977 ;
  assign n45979 = ~n45971 & n45978 ;
  assign n45980 = ~n45882 & n45979 ;
  assign n45981 = ~n45973 & ~n45980 ;
  assign n45982 = ~n45963 & n45981 ;
  assign n45983 = \pi0215  & ~\pi0947  ;
  assign n45984 = \pi0215  & n45968 ;
  assign n45985 = n45972 & n45984 ;
  assign n45986 = ~n45983 & ~n45985 ;
  assign n45987 = ~n45982 & ~n45986 ;
  assign n45988 = \pi0299  & ~n45987 ;
  assign n45989 = ~n45938 & n45988 ;
  assign n45990 = ~n45920 & n45989 ;
  assign n45991 = \pi0039  & ~n45990 ;
  assign n45992 = ~\pi0038  & ~n45991 ;
  assign n45993 = n2165 & ~n45857 ;
  assign n45994 = ~n45856 & n45993 ;
  assign n45995 = ~\pi0223  & ~n45994 ;
  assign n45996 = ~n21285 & n45995 ;
  assign n45997 = ~\pi0210  & n2165 ;
  assign n45998 = ~\pi0223  & ~n45997 ;
  assign n45999 = n21285 & n45998 ;
  assign n46000 = ~n45996 & ~n45999 ;
  assign n46001 = \pi0634  & ~n6714 ;
  assign n46002 = \pi0907  & ~n46001 ;
  assign n46003 = ~n21285 & n46002 ;
  assign n46004 = \pi0210  & ~n6714 ;
  assign n46005 = \pi0907  & ~n46004 ;
  assign n46006 = n21285 & n46005 ;
  assign n46007 = ~n46003 & ~n46006 ;
  assign n46008 = ~n6713 & n42734 ;
  assign n46009 = ~n21403 & n46008 ;
  assign n46010 = ~n21393 & n46008 ;
  assign n46011 = n21398 & n46010 ;
  assign n46012 = ~n46009 & ~n46011 ;
  assign n46013 = \pi0210  & ~n6706 ;
  assign n46014 = ~n6713 & n46013 ;
  assign n46015 = n21403 & n46014 ;
  assign n46016 = ~n21399 & n46015 ;
  assign n46017 = n46012 & ~n46016 ;
  assign n46018 = ~n46007 & n46017 ;
  assign n46019 = ~\pi0907  & ~n45906 ;
  assign n46020 = ~n45943 & n46019 ;
  assign n46021 = ~n45941 & n46020 ;
  assign n46022 = ~\pi0947  & ~n46021 ;
  assign n46023 = ~n46018 & n46022 ;
  assign n46024 = ~\pi0633  & n6713 ;
  assign n46025 = \pi0947  & ~n46024 ;
  assign n46026 = ~n21285 & n46025 ;
  assign n46027 = ~\pi0210  & n6713 ;
  assign n46028 = \pi0947  & ~n46027 ;
  assign n46029 = n21285 & n46028 ;
  assign n46030 = ~n46026 & ~n46029 ;
  assign n46031 = n6761 & n46030 ;
  assign n46032 = ~n21403 & n43044 ;
  assign n46033 = ~n21393 & n43044 ;
  assign n46034 = n21398 & n46033 ;
  assign n46035 = ~n46032 & ~n46034 ;
  assign n46036 = n21403 & n46013 ;
  assign n46037 = ~n21399 & n46036 ;
  assign n46038 = ~\pi0633  & ~n6713 ;
  assign n46039 = ~n6714 & ~n46038 ;
  assign n46040 = ~n21285 & n46039 ;
  assign n46041 = ~\pi0210  & ~n6713 ;
  assign n46042 = ~n6714 & ~n46041 ;
  assign n46043 = n21285 & n46042 ;
  assign n46044 = ~n46040 & ~n46043 ;
  assign n46045 = n6761 & n46044 ;
  assign n46046 = ~n46037 & n46045 ;
  assign n46047 = n46035 & n46046 ;
  assign n46048 = ~n46031 & ~n46047 ;
  assign n46049 = ~n46023 & ~n46048 ;
  assign n46050 = ~n6761 & ~n45973 ;
  assign n46051 = ~\pi0947  & n45959 ;
  assign n46052 = n22183 & n46051 ;
  assign n46053 = ~\pi0947  & ~n45882 ;
  assign n46054 = n45979 & n46053 ;
  assign n46055 = ~n46052 & ~n46054 ;
  assign n46056 = n46050 & n46055 ;
  assign n46057 = \pi0223  & ~n46056 ;
  assign n46058 = ~n46049 & n46057 ;
  assign n46059 = n46000 & ~n46058 ;
  assign n46060 = ~n6761 & n45935 ;
  assign n46061 = n17234 & ~n45924 ;
  assign n46062 = ~n45922 & n46061 ;
  assign n46063 = ~n45884 & n46062 ;
  assign n46064 = ~n46060 & ~n46063 ;
  assign n46065 = \pi0947  & ~n46064 ;
  assign n46066 = \pi0210  & ~\pi0907  ;
  assign n46067 = n21334 & n46066 ;
  assign n46068 = ~n21330 & n46067 ;
  assign n46069 = ~n45892 & ~n46064 ;
  assign n46070 = ~n46068 & n46069 ;
  assign n46071 = ~n46065 & ~n46070 ;
  assign n46072 = ~\pi0907  & n45908 ;
  assign n46073 = ~\pi0907  & ~n21352 ;
  assign n46074 = ~n45913 & n46073 ;
  assign n46075 = ~n46072 & ~n46074 ;
  assign n46076 = ~\pi0947  & n46007 ;
  assign n46077 = ~n45886 & ~n45888 ;
  assign n46078 = ~n45884 & n46077 ;
  assign n46079 = ~\pi0947  & ~n6706 ;
  assign n46080 = ~n6713 & n46079 ;
  assign n46081 = ~n46078 & n46080 ;
  assign n46082 = ~n46076 & ~n46081 ;
  assign n46083 = n46075 & ~n46082 ;
  assign n46084 = ~n45922 & ~n45924 ;
  assign n46085 = ~n45884 & n46084 ;
  assign n46086 = ~n6706 & ~n46030 ;
  assign n46087 = ~n46085 & n46086 ;
  assign n46088 = ~n46030 & ~n46044 ;
  assign n46089 = n6761 & ~n46088 ;
  assign n46090 = ~n46087 & n46089 ;
  assign n46091 = ~n46083 & n46090 ;
  assign n46092 = n46071 & ~n46091 ;
  assign n46093 = ~n2165 & ~n46058 ;
  assign n46094 = ~n46092 & n46093 ;
  assign n46095 = ~n46059 & ~n46094 ;
  assign n46096 = ~\pi0038  & ~\pi0299  ;
  assign n46097 = ~n46095 & n46096 ;
  assign n46098 = ~n45992 & ~n46097 ;
  assign n46099 = ~n45871 & ~n46098 ;
  assign n46100 = ~\pi0210  & ~n11834 ;
  assign n46101 = \pi0210  & ~n21757 ;
  assign n46102 = n1689 & ~n45858 ;
  assign n46103 = n8413 & n46102 ;
  assign n46104 = n1354 & n46103 ;
  assign n46105 = n1358 & n46104 ;
  assign n46106 = \pi0038  & ~n46105 ;
  assign n46107 = ~n46101 & n46106 ;
  assign n46108 = ~n46100 & ~n46107 ;
  assign n46109 = ~n46099 & n46108 ;
  assign n46110 = n6861 & n9948 ;
  assign n46111 = \pi0210  & ~n46110 ;
  assign n46112 = ~n46109 & ~n46111 ;
  assign n46113 = \pi0606  & \pi0643  ;
  assign n46114 = ~n27107 & n43150 ;
  assign n46115 = ~n28108 & n46114 ;
  assign n46116 = n1281 & n6861 ;
  assign n46117 = n28115 & n46116 ;
  assign n46118 = \pi0643  & ~n46117 ;
  assign n46119 = ~n46115 & n46118 ;
  assign n46120 = ~n46113 & ~n46119 ;
  assign n46121 = \pi0211  & ~n43979 ;
  assign n46122 = \pi0211  & ~n28105 ;
  assign n46123 = n28102 & n46122 ;
  assign n46124 = ~n46121 & ~n46123 ;
  assign n46125 = ~n46120 & ~n46124 ;
  assign n46126 = n9948 & n43979 ;
  assign n46127 = ~n27269 & n46126 ;
  assign n46128 = ~\pi0606  & n1289 ;
  assign n46129 = n1287 & n46128 ;
  assign n46130 = ~\pi0038  & n46129 ;
  assign n46131 = n21765 & n46129 ;
  assign n46132 = n1638 & n46131 ;
  assign n46133 = ~n46130 & ~n46132 ;
  assign n46134 = ~\pi0643  & n46133 ;
  assign n46135 = ~\pi0643  & n21770 ;
  assign n46136 = ~n21734 & n46135 ;
  assign n46137 = ~n46134 & ~n46136 ;
  assign n46138 = n9948 & n46137 ;
  assign n46139 = \pi0211  & ~n46138 ;
  assign n46140 = ~n46127 & n46139 ;
  assign n46141 = ~\pi0057  & ~\pi0211  ;
  assign n46142 = n6848 & n46141 ;
  assign n46143 = ~n27308 & ~n27310 ;
  assign n46144 = \pi0606  & ~\pi0643  ;
  assign n46145 = n1289 & n46144 ;
  assign n46146 = n1287 & n46145 ;
  assign n46147 = ~n46143 & n46146 ;
  assign n46148 = n46142 & n46147 ;
  assign n46149 = ~n28061 & n46129 ;
  assign n46150 = ~n28052 & n43979 ;
  assign n46151 = ~n46149 & ~n46150 ;
  assign n46152 = \pi0643  & n46142 ;
  assign n46153 = ~n46151 & n46152 ;
  assign n46154 = ~n46148 & ~n46153 ;
  assign n46155 = ~n46140 & n46154 ;
  assign n46156 = ~n46125 & n46155 ;
  assign n46157 = ~\pi0607  & n1289 ;
  assign n46158 = n1287 & n46157 ;
  assign n46159 = ~n22124 & n46158 ;
  assign n46160 = ~n28084 & n46159 ;
  assign n46161 = ~\pi0638  & ~n46160 ;
  assign n46162 = n27408 & ~n46161 ;
  assign n46163 = \pi0607  & n1289 ;
  assign n46164 = n1287 & n46163 ;
  assign n46165 = n27408 & n46164 ;
  assign n46166 = ~n27269 & n46165 ;
  assign n46167 = ~n46162 & ~n46166 ;
  assign n46168 = ~\pi0212  & n46167 ;
  assign n46169 = \pi0607  & \pi0638  ;
  assign n46170 = \pi0638  & ~n46117 ;
  assign n46171 = ~n46115 & n46170 ;
  assign n46172 = ~n46169 & ~n46171 ;
  assign n46173 = ~\pi0212  & ~n46164 ;
  assign n46174 = ~\pi0212  & ~n28105 ;
  assign n46175 = n28102 & n46174 ;
  assign n46176 = ~n46173 & ~n46175 ;
  assign n46177 = ~n46172 & ~n46176 ;
  assign n46178 = ~n46168 & ~n46177 ;
  assign n46179 = ~\pi0607  & ~n6861 ;
  assign n46180 = ~\pi0607  & ~n28057 ;
  assign n46181 = ~n28060 & n46180 ;
  assign n46182 = ~n46179 & ~n46181 ;
  assign n46183 = ~\pi0607  & \pi0638  ;
  assign n46184 = \pi0638  & n1289 ;
  assign n46185 = n1287 & n46184 ;
  assign n46186 = ~n46183 & ~n46185 ;
  assign n46187 = ~n28048 & ~n46183 ;
  assign n46188 = ~n28051 & n46187 ;
  assign n46189 = ~n46186 & ~n46188 ;
  assign n46190 = n46182 & n46189 ;
  assign n46191 = \pi0607  & ~\pi0638  ;
  assign n46192 = n6861 & n46191 ;
  assign n46193 = ~n46143 & n46192 ;
  assign n46194 = ~n46190 & ~n46193 ;
  assign n46195 = ~\pi0057  & \pi0212  ;
  assign n46196 = n6848 & n46195 ;
  assign n46197 = ~n46194 & n46196 ;
  assign n46198 = n46178 & ~n46197 ;
  assign n46199 = ~\pi0622  & n45713 ;
  assign n46200 = ~n22124 & n46199 ;
  assign n46201 = ~n28084 & n46200 ;
  assign n46202 = ~n46115 & ~n46117 ;
  assign n46203 = ~\pi0622  & \pi0639  ;
  assign n46204 = ~n46202 & n46203 ;
  assign n46205 = ~n46201 & ~n46204 ;
  assign n46206 = ~\pi0057  & ~\pi0213  ;
  assign n46207 = n6848 & n46206 ;
  assign n46208 = ~n46205 & n46207 ;
  assign n46209 = \pi0639  & ~n6861 ;
  assign n46210 = \pi0639  & ~n28105 ;
  assign n46211 = n28102 & n46210 ;
  assign n46212 = ~n46209 & ~n46211 ;
  assign n46213 = ~\pi0639  & ~n27232 ;
  assign n46214 = ~n27268 & n46213 ;
  assign n46215 = ~\pi0639  & ~n6861 ;
  assign n46216 = \pi0622  & ~n46215 ;
  assign n46217 = ~n46214 & n46216 ;
  assign n46218 = n46207 & n46217 ;
  assign n46219 = n46212 & n46218 ;
  assign n46220 = ~n46208 & ~n46219 ;
  assign n46221 = ~\pi0622  & ~n6861 ;
  assign n46222 = ~\pi0622  & ~n28057 ;
  assign n46223 = ~n28060 & n46222 ;
  assign n46224 = ~n46221 & ~n46223 ;
  assign n46225 = \pi0639  & n1289 ;
  assign n46226 = n1287 & n46225 ;
  assign n46227 = ~n46203 & ~n46226 ;
  assign n46228 = ~n28048 & ~n46203 ;
  assign n46229 = ~n28051 & n46228 ;
  assign n46230 = ~n46227 & ~n46229 ;
  assign n46231 = n46224 & n46230 ;
  assign n46232 = \pi0622  & ~\pi0639  ;
  assign n46233 = n6861 & n46232 ;
  assign n46234 = ~n46143 & n46233 ;
  assign n46235 = \pi0213  & ~n46234 ;
  assign n46236 = ~n46231 & n46235 ;
  assign n46237 = \pi0213  & ~n27408 ;
  assign n46238 = ~n46236 & ~n46237 ;
  assign n46239 = n46220 & n46238 ;
  assign n46240 = ~\pi0623  & n1289 ;
  assign n46241 = n1287 & n46240 ;
  assign n46242 = ~n22124 & n46241 ;
  assign n46243 = ~n28084 & n46242 ;
  assign n46244 = ~\pi0710  & ~n46243 ;
  assign n46245 = n27408 & ~n46244 ;
  assign n46246 = \pi0623  & n1289 ;
  assign n46247 = n1287 & n46246 ;
  assign n46248 = n27408 & n46247 ;
  assign n46249 = ~n27269 & n46248 ;
  assign n46250 = ~n46245 & ~n46249 ;
  assign n46251 = ~\pi0214  & n46250 ;
  assign n46252 = \pi0623  & \pi0710  ;
  assign n46253 = \pi0710  & ~n46117 ;
  assign n46254 = ~n46115 & n46253 ;
  assign n46255 = ~n46252 & ~n46254 ;
  assign n46256 = ~\pi0214  & ~n46247 ;
  assign n46257 = ~\pi0214  & ~n28105 ;
  assign n46258 = n28102 & n46257 ;
  assign n46259 = ~n46256 & ~n46258 ;
  assign n46260 = ~n46255 & ~n46259 ;
  assign n46261 = ~n46251 & ~n46260 ;
  assign n46262 = ~\pi0623  & ~n6861 ;
  assign n46263 = ~\pi0623  & ~n28057 ;
  assign n46264 = ~n28060 & n46263 ;
  assign n46265 = ~n46262 & ~n46264 ;
  assign n46266 = ~\pi0623  & \pi0710  ;
  assign n46267 = \pi0710  & n1289 ;
  assign n46268 = n1287 & n46267 ;
  assign n46269 = ~n46266 & ~n46268 ;
  assign n46270 = ~n28048 & ~n46266 ;
  assign n46271 = ~n28051 & n46270 ;
  assign n46272 = ~n46269 & ~n46271 ;
  assign n46273 = n46265 & n46272 ;
  assign n46274 = \pi0623  & ~\pi0710  ;
  assign n46275 = n6861 & n46274 ;
  assign n46276 = ~n46143 & n46275 ;
  assign n46277 = ~n46273 & ~n46276 ;
  assign n46278 = ~\pi0057  & \pi0214  ;
  assign n46279 = n6848 & n46278 ;
  assign n46280 = ~n46277 & n46279 ;
  assign n46281 = n46261 & ~n46280 ;
  assign n46282 = \pi0681  & \pi0907  ;
  assign n46283 = ~\pi0947  & ~n46282 ;
  assign n46284 = ~n29026 & n46283 ;
  assign n46285 = \pi0642  & n6761 ;
  assign n46286 = n6761 & ~n21407 ;
  assign n46287 = ~n46285 & ~n46286 ;
  assign n46288 = ~\pi0616  & ~n21632 ;
  assign n46289 = ~n21631 & n46288 ;
  assign n46290 = ~n6709 & ~n21570 ;
  assign n46291 = ~n46285 & n46290 ;
  assign n46292 = ~n46289 & n46291 ;
  assign n46293 = ~n46287 & ~n46292 ;
  assign n46294 = n6707 & n6708 ;
  assign n46295 = n21403 & n46294 ;
  assign n46296 = ~n21399 & n46295 ;
  assign n46297 = ~\pi0642  & ~n46296 ;
  assign n46298 = ~n21615 & n46297 ;
  assign n46299 = ~n21645 & n46298 ;
  assign n46300 = ~\pi0642  & n6709 ;
  assign n46301 = ~n46296 & n46300 ;
  assign n46302 = ~n6761 & ~n46301 ;
  assign n46303 = ~n46299 & n46302 ;
  assign n46304 = \pi0947  & ~n46303 ;
  assign n46305 = ~n46293 & n46304 ;
  assign n46306 = ~\pi0947  & n46282 ;
  assign n46307 = \pi0223  & ~n46306 ;
  assign n46308 = n46305 & n46307 ;
  assign n46309 = n21651 & n46307 ;
  assign n46310 = ~n27183 & n46309 ;
  assign n46311 = ~n46308 & ~n46310 ;
  assign n46312 = ~n21285 & n21370 ;
  assign n46313 = n21363 & n21370 ;
  assign n46314 = ~n46312 & ~n46313 ;
  assign n46315 = n21355 & ~n46314 ;
  assign n46316 = ~n21290 & ~n46314 ;
  assign n46317 = ~n21325 & n46316 ;
  assign n46318 = ~n46315 & ~n46317 ;
  assign n46319 = ~\pi0603  & n21370 ;
  assign n46320 = ~n21285 & n46319 ;
  assign n46321 = ~\pi0642  & ~n6711 ;
  assign n46322 = ~n21285 & n46321 ;
  assign n46323 = ~n6709 & ~n46322 ;
  assign n46324 = ~n46320 & n46323 ;
  assign n46325 = n46318 & n46324 ;
  assign n46326 = ~\pi0642  & ~n21352 ;
  assign n46327 = n21355 & n46326 ;
  assign n46328 = ~n21290 & n46326 ;
  assign n46329 = ~n21325 & n46328 ;
  assign n46330 = ~n46327 & ~n46329 ;
  assign n46331 = n6709 & n46330 ;
  assign n46332 = ~n46325 & ~n46331 ;
  assign n46333 = n6761 & n46332 ;
  assign n46334 = ~\pi0642  & ~n6761 ;
  assign n46335 = ~n21334 & n46334 ;
  assign n46336 = n6713 & n46334 ;
  assign n46337 = ~n21329 & n46336 ;
  assign n46338 = ~n46335 & ~n46337 ;
  assign n46339 = ~n46333 & n46338 ;
  assign n46340 = \pi0947  & ~n46339 ;
  assign n46341 = ~n2165 & ~n46340 ;
  assign n46342 = n46311 & n46341 ;
  assign n46343 = ~n46284 & n46342 ;
  assign n46344 = \pi0642  & \pi0947  ;
  assign n46345 = ~n46306 & ~n46344 ;
  assign n46346 = n2165 & ~n46345 ;
  assign n46347 = ~n21285 & n46346 ;
  assign n46348 = ~\pi0223  & ~n46347 ;
  assign n46349 = ~n21905 & n46282 ;
  assign n46350 = ~n22039 & n46349 ;
  assign n46351 = ~\pi0947  & ~n46350 ;
  assign n46352 = ~n6709 & ~n21286 ;
  assign n46353 = n21328 & n46352 ;
  assign n46354 = n6709 & ~n21306 ;
  assign n46355 = ~n21903 & n46354 ;
  assign n46356 = \pi0642  & ~\pi0662  ;
  assign n46357 = n6708 & n46356 ;
  assign n46358 = ~n46355 & n46357 ;
  assign n46359 = ~n46353 & n46358 ;
  assign n46360 = ~\pi0642  & \pi0947  ;
  assign n46361 = ~\pi0662  & \pi0947  ;
  assign n46362 = n6708 & n46361 ;
  assign n46363 = ~n46360 & ~n46362 ;
  assign n46364 = \pi0947  & ~n21286 ;
  assign n46365 = n21328 & n46364 ;
  assign n46366 = n46363 & ~n46365 ;
  assign n46367 = ~n46359 & ~n46366 ;
  assign n46368 = ~n46351 & ~n46367 ;
  assign n46369 = ~n6761 & ~n46368 ;
  assign n46370 = ~n2165 & ~n46369 ;
  assign n46371 = \pi0616  & n46306 ;
  assign n46372 = ~n21577 & n46306 ;
  assign n46373 = ~n21576 & n46372 ;
  assign n46374 = ~n46371 & ~n46373 ;
  assign n46375 = ~n21570 & ~n46374 ;
  assign n46376 = ~\pi0947  & n6761 ;
  assign n46377 = ~n21285 & n46357 ;
  assign n46378 = n21882 & n46357 ;
  assign n46379 = ~n46377 & ~n46378 ;
  assign n46380 = n21355 & ~n46379 ;
  assign n46381 = ~n21290 & ~n46379 ;
  assign n46382 = ~n21325 & n46381 ;
  assign n46383 = ~n46380 & ~n46382 ;
  assign n46384 = ~\pi0680  & n46357 ;
  assign n46385 = ~n21285 & n46384 ;
  assign n46386 = \pi0642  & ~n21586 ;
  assign n46387 = ~n21285 & n46386 ;
  assign n46388 = n6761 & ~n46387 ;
  assign n46389 = ~n46385 & n46388 ;
  assign n46390 = n46383 & n46389 ;
  assign n46391 = ~n46376 & ~n46390 ;
  assign n46392 = ~n46375 & ~n46391 ;
  assign n46393 = n46370 & ~n46392 ;
  assign n46394 = n46348 & ~n46393 ;
  assign n46395 = ~\pi0215  & ~\pi0299  ;
  assign n46396 = n2352 & ~n46345 ;
  assign n46397 = ~\pi0215  & n46396 ;
  assign n46398 = ~n21285 & n46397 ;
  assign n46399 = ~n46395 & ~n46398 ;
  assign n46400 = ~n21582 & n46357 ;
  assign n46401 = ~\pi0680  & n46400 ;
  assign n46402 = ~n21352 & n46400 ;
  assign n46403 = ~n21405 & n46402 ;
  assign n46404 = ~n46401 & ~n46403 ;
  assign n46405 = \pi0947  & ~n46387 ;
  assign n46406 = n46404 & n46405 ;
  assign n46407 = \pi0223  & n46406 ;
  assign n46408 = ~n21615 & ~n21645 ;
  assign n46409 = ~n22079 & ~n27180 ;
  assign n46410 = \pi0223  & ~n46409 ;
  assign n46411 = ~n46408 & n46410 ;
  assign n46412 = ~n46407 & ~n46411 ;
  assign n46413 = ~\pi0616  & n6761 ;
  assign n46414 = ~n21632 & n46413 ;
  assign n46415 = ~n21631 & n46414 ;
  assign n46416 = \pi0616  & n6761 ;
  assign n46417 = n21285 & n46416 ;
  assign n46418 = n46282 & ~n46417 ;
  assign n46419 = ~n46415 & n46418 ;
  assign n46420 = \pi0223  & ~\pi0947  ;
  assign n46421 = ~n46419 & n46420 ;
  assign n46422 = n46412 & ~n46421 ;
  assign n46423 = ~n46399 & n46422 ;
  assign n46424 = n24388 & n46422 ;
  assign n46425 = n46368 & n46424 ;
  assign n46426 = ~n46423 & ~n46425 ;
  assign n46427 = ~n46394 & ~n46426 ;
  assign n46428 = \pi0299  & ~n46399 ;
  assign n46429 = n27078 & n46368 ;
  assign n46430 = ~n46428 & ~n46429 ;
  assign n46431 = \pi0039  & n46430 ;
  assign n46432 = ~\pi0223  & ~n46344 ;
  assign n46433 = ~n46306 & n46432 ;
  assign n46434 = ~n22316 & ~n46433 ;
  assign n46435 = ~\pi0222  & ~\pi0224  ;
  assign n46436 = n21285 & n46435 ;
  assign n46437 = ~n46434 & ~n46436 ;
  assign n46438 = n46311 & ~n46437 ;
  assign n46439 = ~\pi0299  & ~n46438 ;
  assign n46440 = n46431 & n46439 ;
  assign n46441 = ~n46427 & n46440 ;
  assign n46442 = ~n46343 & n46441 ;
  assign n46443 = ~\pi0947  & ~n27082 ;
  assign n46444 = ~n21724 & n46443 ;
  assign n46445 = \pi0299  & ~n46306 ;
  assign n46446 = \pi0947  & ~n46301 ;
  assign n46447 = ~n46299 & n46446 ;
  assign n46448 = n46445 & ~n46447 ;
  assign n46449 = ~n46444 & n46448 ;
  assign n46450 = \pi0215  & ~n46449 ;
  assign n46451 = n46431 & ~n46450 ;
  assign n46452 = ~n46427 & n46451 ;
  assign n46453 = ~n21205 & n46345 ;
  assign n46454 = ~n21238 & n46453 ;
  assign n46455 = ~n2259 & ~n26957 ;
  assign n46456 = ~n2259 & n21237 ;
  assign n46457 = n21232 & n46456 ;
  assign n46458 = ~n46455 & ~n46457 ;
  assign n46459 = ~n46454 & n46458 ;
  assign n46460 = ~n21740 & n46345 ;
  assign n46461 = ~n21738 & n46460 ;
  assign n46462 = \pi0215  & ~\pi0299  ;
  assign n46463 = ~n27218 & ~n46462 ;
  assign n46464 = n21737 & ~n46462 ;
  assign n46465 = n21232 & n46464 ;
  assign n46466 = ~n46463 & ~n46465 ;
  assign n46467 = ~n46461 & n46466 ;
  assign n46468 = ~n46459 & ~n46467 ;
  assign n46469 = ~\pi0039  & n46468 ;
  assign n46470 = ~\pi0038  & ~n46469 ;
  assign n46471 = ~n46452 & n46470 ;
  assign n46472 = ~n46442 & n46471 ;
  assign n46473 = n46110 & n46472 ;
  assign n46474 = ~\pi0215  & ~n21757 ;
  assign n46475 = n1689 & ~n46344 ;
  assign n46476 = ~n46306 & n46475 ;
  assign n46477 = n8413 & n46476 ;
  assign n46478 = n1354 & n46477 ;
  assign n46479 = n1358 & n46478 ;
  assign n46480 = n11835 & ~n46479 ;
  assign n46481 = ~n46474 & n46480 ;
  assign n46482 = \pi0215  & ~n46110 ;
  assign n46483 = ~n46481 & ~n46482 ;
  assign n46484 = ~n46473 & n46483 ;
  assign n46485 = \pi0662  & \pi0907  ;
  assign n46486 = ~\pi0947  & n46485 ;
  assign n46487 = \pi0614  & \pi0947  ;
  assign n46488 = ~n46486 & ~n46487 ;
  assign n46489 = ~n6761 & n46488 ;
  assign n46490 = ~n21334 & n46489 ;
  assign n46491 = n6713 & n46489 ;
  assign n46492 = ~n21329 & n46491 ;
  assign n46493 = ~n46490 & ~n46492 ;
  assign n46494 = ~n46435 & n46493 ;
  assign n46495 = \pi0947  & ~n21602 ;
  assign n46496 = ~n21599 & n46495 ;
  assign n46497 = n6761 & n46496 ;
  assign n46498 = n21593 & ~n46485 ;
  assign n46499 = ~n21602 & ~n46485 ;
  assign n46500 = ~n21599 & n46499 ;
  assign n46501 = ~n46498 & ~n46500 ;
  assign n46502 = ~\pi0947  & ~n46501 ;
  assign n46503 = n6761 & ~n21581 ;
  assign n46504 = n46502 & n46503 ;
  assign n46505 = ~n46497 & ~n46504 ;
  assign n46506 = n46494 & n46505 ;
  assign n46507 = n2165 & n21285 ;
  assign n46508 = \pi0216  & ~n46507 ;
  assign n46509 = ~\pi0223  & ~n46487 ;
  assign n46510 = ~n46486 & n46509 ;
  assign n46511 = ~n22316 & ~n46510 ;
  assign n46512 = n46508 & ~n46511 ;
  assign n46513 = ~n46506 & n46512 ;
  assign n46514 = \pi0223  & ~n46486 ;
  assign n46515 = \pi0614  & n6761 ;
  assign n46516 = \pi0616  & ~n6709 ;
  assign n46517 = ~n21285 & n46516 ;
  assign n46518 = ~n6709 & ~n21285 ;
  assign n46519 = ~\pi0616  & n6710 ;
  assign n46520 = ~n6709 & n46519 ;
  assign n46521 = ~n46518 & ~n46520 ;
  assign n46522 = ~n21622 & ~n46521 ;
  assign n46523 = ~n21619 & n46522 ;
  assign n46524 = ~n46517 & ~n46523 ;
  assign n46525 = n46286 & n46524 ;
  assign n46526 = n21429 & n42695 ;
  assign n46527 = n21429 & n21908 ;
  assign n46528 = n21520 & n46527 ;
  assign n46529 = ~n46526 & ~n46528 ;
  assign n46530 = \pi0947  & n6761 ;
  assign n46531 = ~\pi0614  & \pi0947  ;
  assign n46532 = ~n46296 & n46531 ;
  assign n46533 = ~n46530 & ~n46532 ;
  assign n46534 = n46529 & ~n46533 ;
  assign n46535 = ~n46525 & n46534 ;
  assign n46536 = ~n46515 & n46535 ;
  assign n46537 = \pi0216  & n46536 ;
  assign n46538 = \pi0216  & n21651 ;
  assign n46539 = ~n27183 & n46538 ;
  assign n46540 = ~n46537 & ~n46539 ;
  assign n46541 = n46514 & ~n46540 ;
  assign n46542 = \pi0616  & n46486 ;
  assign n46543 = ~n21577 & n46486 ;
  assign n46544 = ~n21576 & n46543 ;
  assign n46545 = ~n46542 & ~n46544 ;
  assign n46546 = ~n21570 & ~n46545 ;
  assign n46547 = n2165 & ~n46488 ;
  assign n46548 = ~n21285 & n46547 ;
  assign n46549 = n6761 & ~n21588 ;
  assign n46550 = ~n21585 & n46549 ;
  assign n46551 = \pi0680  & n46549 ;
  assign n46552 = n21359 & n46551 ;
  assign n46553 = ~n46550 & ~n46552 ;
  assign n46554 = ~n46376 & n46553 ;
  assign n46555 = ~n46548 & ~n46554 ;
  assign n46556 = ~n46546 & n46555 ;
  assign n46557 = n46435 & ~n46488 ;
  assign n46558 = ~n21285 & n46557 ;
  assign n46559 = n2165 & ~n46558 ;
  assign n46560 = ~n46355 & n46487 ;
  assign n46561 = ~n46353 & n46560 ;
  assign n46562 = ~n21905 & n46486 ;
  assign n46563 = ~n22039 & n46562 ;
  assign n46564 = ~n46561 & ~n46563 ;
  assign n46565 = ~n6761 & ~n46558 ;
  assign n46566 = n46564 & n46565 ;
  assign n46567 = ~n46559 & ~n46566 ;
  assign n46568 = ~\pi0223  & n46567 ;
  assign n46569 = ~n46556 & n46568 ;
  assign n46570 = \pi0223  & n21587 ;
  assign n46571 = ~n21285 & n46570 ;
  assign n46572 = ~n46420 & ~n46571 ;
  assign n46573 = \pi0223  & n6708 ;
  assign n46574 = n21583 & n46573 ;
  assign n46575 = ~n21582 & n46574 ;
  assign n46576 = ~\pi0680  & n46575 ;
  assign n46577 = ~n21352 & n46575 ;
  assign n46578 = ~n21405 & n46577 ;
  assign n46579 = ~n46576 & ~n46578 ;
  assign n46580 = n46572 & n46579 ;
  assign n46581 = ~\pi0216  & n46580 ;
  assign n46582 = ~\pi0216  & ~n46409 ;
  assign n46583 = ~n46408 & n46582 ;
  assign n46584 = ~n46581 & ~n46583 ;
  assign n46585 = ~\pi0216  & ~\pi0947  ;
  assign n46586 = ~n46417 & n46485 ;
  assign n46587 = ~n46415 & n46586 ;
  assign n46588 = n46585 & ~n46587 ;
  assign n46589 = n46584 & ~n46588 ;
  assign n46590 = ~n46569 & ~n46589 ;
  assign n46591 = ~n46541 & ~n46590 ;
  assign n46592 = ~n46513 & n46591 ;
  assign n46593 = ~n21740 & ~n46488 ;
  assign n46594 = ~n21738 & n46593 ;
  assign n46595 = \pi0216  & n21740 ;
  assign n46596 = \pi0216  & n21737 ;
  assign n46597 = n21232 & n46596 ;
  assign n46598 = ~n46595 & ~n46597 ;
  assign n46599 = ~\pi0299  & n46598 ;
  assign n46600 = ~n46594 & n46599 ;
  assign n46601 = ~n21205 & ~n46488 ;
  assign n46602 = ~n21238 & n46601 ;
  assign n46603 = ~n13621 & ~n26957 ;
  assign n46604 = ~n13621 & n21237 ;
  assign n46605 = n21232 & n46604 ;
  assign n46606 = ~n46603 & ~n46605 ;
  assign n46607 = ~n46602 & n46606 ;
  assign n46608 = ~\pi0039  & ~n46607 ;
  assign n46609 = ~n46600 & n46608 ;
  assign n46610 = n46096 & ~n46609 ;
  assign n46611 = ~n46592 & n46610 ;
  assign n46612 = ~\pi0614  & ~n46296 ;
  assign n46613 = \pi0947  & ~n46612 ;
  assign n46614 = \pi0947  & ~n6709 ;
  assign n46615 = n42695 & n46614 ;
  assign n46616 = n21908 & n46614 ;
  assign n46617 = n21520 & n46616 ;
  assign n46618 = ~n46615 & ~n46617 ;
  assign n46619 = ~n46613 & n46618 ;
  assign n46620 = \pi0216  & \pi0299  ;
  assign n46621 = ~n46486 & n46620 ;
  assign n46622 = n46619 & n46621 ;
  assign n46623 = ~\pi0947  & ~n46486 ;
  assign n46624 = ~n21286 & ~n46486 ;
  assign n46625 = n21520 & n46624 ;
  assign n46626 = ~n46623 & ~n46625 ;
  assign n46627 = ~\pi0216  & ~n46626 ;
  assign n46628 = ~\pi0680  & n21585 ;
  assign n46629 = ~n21352 & n21585 ;
  assign n46630 = ~n21405 & n46629 ;
  assign n46631 = ~n46628 & ~n46630 ;
  assign n46632 = \pi0947  & ~n21588 ;
  assign n46633 = ~\pi0216  & n46632 ;
  assign n46634 = n46631 & n46633 ;
  assign n46635 = ~n46627 & ~n46634 ;
  assign n46636 = \pi0215  & n46635 ;
  assign n46637 = ~\pi0216  & ~n21286 ;
  assign n46638 = n21520 & n46637 ;
  assign n46639 = ~n46585 & ~n46638 ;
  assign n46640 = ~n46408 & ~n46639 ;
  assign n46641 = \pi0039  & ~n46640 ;
  assign n46642 = n46636 & n46641 ;
  assign n46643 = ~n27982 & ~n46642 ;
  assign n46644 = ~n46622 & ~n46643 ;
  assign n46645 = n46443 & ~n46643 ;
  assign n46646 = ~n21724 & n46645 ;
  assign n46647 = ~n46644 & ~n46646 ;
  assign n46648 = \pi0216  & n6730 ;
  assign n46649 = n21694 & n46648 ;
  assign n46650 = ~n21711 & n46649 ;
  assign n46651 = \pi0216  & ~n6732 ;
  assign n46652 = n21334 & n46651 ;
  assign n46653 = ~n21330 & n46652 ;
  assign n46654 = \pi0216  & n46487 ;
  assign n46655 = \pi0216  & ~\pi0947  ;
  assign n46656 = n46485 & n46655 ;
  assign n46657 = ~n46654 & ~n46656 ;
  assign n46658 = n2352 & ~n46488 ;
  assign n46659 = ~n21285 & n46658 ;
  assign n46660 = n46657 & ~n46659 ;
  assign n46661 = \pi0221  & ~n46564 ;
  assign n46662 = n46660 & ~n46661 ;
  assign n46663 = ~n46653 & n46662 ;
  assign n46664 = ~n46650 & n46663 ;
  assign n46665 = n43041 & ~n46664 ;
  assign n46666 = n46647 & ~n46665 ;
  assign n46667 = ~\pi0038  & ~n46609 ;
  assign n46668 = n46666 & n46667 ;
  assign n46669 = ~\pi0216  & ~n11834 ;
  assign n46670 = \pi0216  & ~n21757 ;
  assign n46671 = n1689 & ~n46488 ;
  assign n46672 = n8413 & n46671 ;
  assign n46673 = n26939 & n46672 ;
  assign n46674 = n10323 & n46673 ;
  assign n46675 = \pi0038  & ~n46674 ;
  assign n46676 = ~n46670 & n46675 ;
  assign n46677 = ~n46669 & ~n46676 ;
  assign n46678 = ~n46668 & n46677 ;
  assign n46679 = ~n46611 & n46678 ;
  assign n46680 = \pi0216  & ~n46110 ;
  assign n46681 = ~n46679 & ~n46680 ;
  assign n46682 = ~n21768 & n27408 ;
  assign n46683 = \pi0695  & ~n46682 ;
  assign n46684 = \pi0695  & n21770 ;
  assign n46685 = ~n21734 & n46684 ;
  assign n46686 = ~n46683 & ~n46685 ;
  assign n46687 = ~\pi0217  & n46686 ;
  assign n46688 = \pi0695  & n46687 ;
  assign n46689 = ~n45761 & n45763 ;
  assign n46690 = n46687 & n46689 ;
  assign n46691 = n45760 & n46690 ;
  assign n46692 = ~n46688 & ~n46691 ;
  assign n46693 = ~\pi0057  & ~\pi0695  ;
  assign n46694 = n6848 & n46693 ;
  assign n46695 = n45818 & n46694 ;
  assign n46696 = ~n24761 & n46694 ;
  assign n46697 = ~n45836 & n46696 ;
  assign n46698 = ~n46695 & ~n46697 ;
  assign n46699 = \pi0217  & n46698 ;
  assign n46700 = ~\pi0612  & ~n46699 ;
  assign n46701 = n46692 & n46700 ;
  assign n46702 = ~\pi0695  & ~n45692 ;
  assign n46703 = ~\pi0695  & \pi0790  ;
  assign n46704 = ~n45683 & n46703 ;
  assign n46705 = ~n46702 & ~n46704 ;
  assign n46706 = \pi0695  & n45706 ;
  assign n46707 = \pi0695  & \pi0790  ;
  assign n46708 = n45672 & n46707 ;
  assign n46709 = ~n46706 & ~n46708 ;
  assign n46710 = ~\pi0217  & n46709 ;
  assign n46711 = n46705 & n46710 ;
  assign n46712 = ~\pi0217  & \pi0612  ;
  assign n46713 = \pi0612  & \pi0695  ;
  assign n46714 = ~n45849 & n46713 ;
  assign n46715 = ~n46712 & ~n46714 ;
  assign n46716 = \pi0612  & ~\pi0695  ;
  assign n46717 = n46715 & ~n46716 ;
  assign n46718 = ~n45812 & n46715 ;
  assign n46719 = ~n45792 & n46718 ;
  assign n46720 = ~n46717 & ~n46719 ;
  assign n46721 = ~n46711 & n46720 ;
  assign n46722 = ~n46701 & ~n46721 ;
  assign n46723 = \pi0218  & n44573 ;
  assign n46724 = ~n44593 & n46723 ;
  assign n46725 = n44590 & n46724 ;
  assign n46726 = ~\pi0057  & n44573 ;
  assign n46727 = ~n44704 & n46726 ;
  assign n46728 = ~n44700 & n46727 ;
  assign n46729 = n44573 & ~n44711 ;
  assign n46730 = n44573 & ~n44593 ;
  assign n46731 = n44590 & n46730 ;
  assign n46732 = \pi0218  & ~n46731 ;
  assign n46733 = ~n44573 & n44757 ;
  assign n46734 = n44755 & n46733 ;
  assign n46735 = ~n46732 & ~n46734 ;
  assign n46736 = ~n46729 & n46735 ;
  assign n46737 = ~n46728 & n46736 ;
  assign n46738 = ~n46725 & ~n46737 ;
  assign n46739 = \pi0617  & \pi0637  ;
  assign n46740 = \pi0637  & ~n46117 ;
  assign n46741 = ~n46115 & n46740 ;
  assign n46742 = ~n46739 & ~n46741 ;
  assign n46743 = \pi0617  & n1289 ;
  assign n46744 = n1287 & n46743 ;
  assign n46745 = \pi0219  & ~n46744 ;
  assign n46746 = \pi0219  & ~n28105 ;
  assign n46747 = n28102 & n46746 ;
  assign n46748 = ~n46745 & ~n46747 ;
  assign n46749 = ~n46742 & ~n46748 ;
  assign n46750 = ~\pi0057  & ~\pi0219  ;
  assign n46751 = n6848 & n46750 ;
  assign n46752 = ~\pi0617  & ~n6861 ;
  assign n46753 = ~\pi0617  & ~n28057 ;
  assign n46754 = ~n28060 & n46753 ;
  assign n46755 = ~n46752 & ~n46754 ;
  assign n46756 = ~\pi0617  & \pi0637  ;
  assign n46757 = \pi0637  & n1289 ;
  assign n46758 = n1287 & n46757 ;
  assign n46759 = ~n46756 & ~n46758 ;
  assign n46760 = ~n28048 & ~n46756 ;
  assign n46761 = ~n28051 & n46760 ;
  assign n46762 = ~n46759 & ~n46761 ;
  assign n46763 = n46755 & n46762 ;
  assign n46764 = \pi0617  & ~\pi0637  ;
  assign n46765 = n6861 & n46764 ;
  assign n46766 = ~n46143 & n46765 ;
  assign n46767 = ~n46763 & ~n46766 ;
  assign n46768 = n46751 & ~n46767 ;
  assign n46769 = \pi0617  & ~n27232 ;
  assign n46770 = ~n27268 & n46769 ;
  assign n46771 = ~\pi0617  & n21768 ;
  assign n46772 = ~\pi0617  & n21770 ;
  assign n46773 = ~n21734 & n46772 ;
  assign n46774 = ~n46771 & ~n46773 ;
  assign n46775 = \pi0617  & ~n6861 ;
  assign n46776 = n27408 & ~n46775 ;
  assign n46777 = n46774 & n46776 ;
  assign n46778 = ~n46770 & n46777 ;
  assign n46779 = ~\pi0057  & \pi0637  ;
  assign n46780 = n6848 & n46779 ;
  assign n46781 = \pi0219  & ~n46780 ;
  assign n46782 = ~n46778 & n46781 ;
  assign n46783 = ~n46768 & ~n46782 ;
  assign n46784 = ~n46749 & n46783 ;
  assign n46785 = ~\pi0220  & n44782 ;
  assign n46786 = ~n44494 & n46785 ;
  assign n46787 = ~n44492 & n46786 ;
  assign n46788 = ~\pi0220  & ~n44782 ;
  assign n46789 = n44540 & n46788 ;
  assign n46790 = n44531 & n46789 ;
  assign n46791 = ~n44549 & n44782 ;
  assign n46792 = ~n44547 & n46791 ;
  assign n46793 = ~n44546 & n46792 ;
  assign n46794 = \pi0220  & ~n46793 ;
  assign n46795 = ~n46790 & ~n46794 ;
  assign n46796 = ~n46787 & n46795 ;
  assign n46797 = \pi0661  & \pi0907  ;
  assign n46798 = ~n27077 & ~n46797 ;
  assign n46799 = n6730 & ~n46797 ;
  assign n46800 = ~n21696 & n46799 ;
  assign n46801 = ~n46798 & ~n46800 ;
  assign n46802 = n21694 & ~n46798 ;
  assign n46803 = ~n21711 & n46802 ;
  assign n46804 = ~n46801 & ~n46803 ;
  assign n46805 = \pi0616  & \pi0947  ;
  assign n46806 = ~\pi0216  & n46805 ;
  assign n46807 = n46585 & n46797 ;
  assign n46808 = ~n46806 & ~n46807 ;
  assign n46809 = ~\pi0215  & ~n46808 ;
  assign n46810 = ~n21285 & n46809 ;
  assign n46811 = ~n6936 & ~n46810 ;
  assign n46812 = ~\pi0947  & ~n46811 ;
  assign n46813 = ~n46355 & n46805 ;
  assign n46814 = ~n46353 & n46813 ;
  assign n46815 = ~\pi0947  & n46797 ;
  assign n46816 = ~n21905 & n46815 ;
  assign n46817 = ~n22039 & n46816 ;
  assign n46818 = ~n46814 & ~n46817 ;
  assign n46819 = ~\pi0215  & \pi0216  ;
  assign n46820 = ~\pi0947  & n46819 ;
  assign n46821 = ~n46818 & n46820 ;
  assign n46822 = ~n46812 & ~n46821 ;
  assign n46823 = ~n46804 & ~n46822 ;
  assign n46824 = ~n21328 & n21660 ;
  assign n46825 = ~\pi0614  & ~n21574 ;
  assign n46826 = ~n21573 & n46825 ;
  assign n46827 = ~n6706 & ~n21577 ;
  assign n46828 = n21660 & n46827 ;
  assign n46829 = ~n46826 & n46828 ;
  assign n46830 = ~n46824 & ~n46829 ;
  assign n46831 = ~\pi0642  & n21674 ;
  assign n46832 = ~n21334 & n46831 ;
  assign n46833 = n6713 & n46831 ;
  assign n46834 = ~n21329 & n46833 ;
  assign n46835 = ~n46832 & ~n46834 ;
  assign n46836 = n21674 & n46357 ;
  assign n46837 = ~n46355 & n46836 ;
  assign n46838 = ~n46353 & n46837 ;
  assign n46839 = \pi0947  & ~n46838 ;
  assign n46840 = n46835 & n46839 ;
  assign n46841 = n46830 & n46840 ;
  assign n46842 = \pi0221  & ~n46841 ;
  assign n46843 = ~n46818 & n46819 ;
  assign n46844 = n46811 & ~n46843 ;
  assign n46845 = ~n46842 & ~n46844 ;
  assign n46846 = ~\pi0947  & ~n46815 ;
  assign n46847 = ~n21681 & ~n46815 ;
  assign n46848 = n21668 & n46847 ;
  assign n46849 = ~n46846 & ~n46848 ;
  assign n46850 = ~\pi0221  & ~n46849 ;
  assign n46851 = ~\pi0221  & ~\pi0947  ;
  assign n46852 = ~\pi0221  & ~n21286 ;
  assign n46853 = n21520 & n46852 ;
  assign n46854 = ~n46851 & ~n46853 ;
  assign n46855 = ~n46408 & ~n46854 ;
  assign n46856 = \pi0215  & ~n46855 ;
  assign n46857 = ~n46850 & n46856 ;
  assign n46858 = \pi0221  & ~\pi0947  ;
  assign n46859 = ~n46797 & n46858 ;
  assign n46860 = n21600 & ~n21624 ;
  assign n46861 = n21520 & n46352 ;
  assign n46862 = \pi0221  & ~n46815 ;
  assign n46863 = ~\pi0616  & n46862 ;
  assign n46864 = ~n46296 & n46863 ;
  assign n46865 = ~n46861 & n46864 ;
  assign n46866 = ~n46860 & n46865 ;
  assign n46867 = ~n46859 & ~n46866 ;
  assign n46868 = n46857 & n46867 ;
  assign n46869 = n46443 & n46857 ;
  assign n46870 = ~n21724 & n46869 ;
  assign n46871 = ~n46868 & ~n46870 ;
  assign n46872 = \pi0299  & n46871 ;
  assign n46873 = ~n46845 & n46872 ;
  assign n46874 = ~n46823 & n46873 ;
  assign n46875 = \pi0039  & ~n46874 ;
  assign n46876 = ~\pi0947  & ~n46797 ;
  assign n46877 = ~n29026 & n46876 ;
  assign n46878 = ~n6761 & ~n46838 ;
  assign n46879 = n46835 & n46878 ;
  assign n46880 = n46830 & n46879 ;
  assign n46881 = ~n46435 & n46880 ;
  assign n46882 = \pi0680  & n21359 ;
  assign n46883 = n21585 & ~n46882 ;
  assign n46884 = n21674 & n46883 ;
  assign n46885 = ~n21602 & n21674 ;
  assign n46886 = ~n21599 & n46885 ;
  assign n46887 = ~n46884 & ~n46886 ;
  assign n46888 = \pi0947  & ~n46887 ;
  assign n46889 = ~n21577 & n21660 ;
  assign n46890 = ~n46826 & n46889 ;
  assign n46891 = n6758 & n6759 ;
  assign n46892 = n6757 & n46891 ;
  assign n46893 = ~n46890 & n46892 ;
  assign n46894 = \pi0947  & ~n46893 ;
  assign n46895 = ~n46435 & ~n46894 ;
  assign n46896 = ~n46888 & n46895 ;
  assign n46897 = ~n46881 & ~n46896 ;
  assign n46898 = ~n46877 & ~n46897 ;
  assign n46899 = \pi0616  & n46815 ;
  assign n46900 = ~n21577 & n46815 ;
  assign n46901 = ~n21576 & n46900 ;
  assign n46902 = ~n46899 & ~n46901 ;
  assign n46903 = ~n21570 & ~n46902 ;
  assign n46904 = ~n46805 & ~n46815 ;
  assign n46905 = n2165 & ~n46904 ;
  assign n46906 = ~n21285 & n46905 ;
  assign n46907 = ~\pi0223  & ~n46906 ;
  assign n46908 = n6761 & ~n21681 ;
  assign n46909 = ~n21664 & n46908 ;
  assign n46910 = \pi0680  & n46908 ;
  assign n46911 = n21359 & n46910 ;
  assign n46912 = ~n46909 & ~n46911 ;
  assign n46913 = ~n46376 & n46912 ;
  assign n46914 = n46907 & ~n46913 ;
  assign n46915 = ~n46903 & n46914 ;
  assign n46916 = n46435 & n46907 ;
  assign n46917 = ~n6761 & n46907 ;
  assign n46918 = n46818 & n46917 ;
  assign n46919 = ~n46916 & ~n46918 ;
  assign n46920 = ~n46415 & ~n46417 ;
  assign n46921 = n21668 & ~n21681 ;
  assign n46922 = \pi0947  & ~n46921 ;
  assign n46923 = ~n46920 & ~n46922 ;
  assign n46924 = ~n46408 & ~n46409 ;
  assign n46925 = n46849 & ~n46924 ;
  assign n46926 = ~n46923 & n46925 ;
  assign n46927 = \pi0223  & ~n46926 ;
  assign n46928 = ~\pi0221  & ~n46927 ;
  assign n46929 = n46919 & n46928 ;
  assign n46930 = ~n46915 & n46929 ;
  assign n46931 = ~\pi0299  & ~n46930 ;
  assign n46932 = ~\pi0223  & ~n46805 ;
  assign n46933 = ~n46815 & n46932 ;
  assign n46934 = ~n21285 & n46933 ;
  assign n46935 = ~n22316 & ~n46934 ;
  assign n46936 = n46931 & ~n46935 ;
  assign n46937 = ~n46898 & n46936 ;
  assign n46938 = n1689 & ~n46904 ;
  assign n46939 = n8413 & n46938 ;
  assign n46940 = n26939 & n46939 ;
  assign n46941 = n10323 & n46940 ;
  assign n46942 = \pi0038  & ~n46941 ;
  assign n46943 = \pi0221  & ~n21757 ;
  assign n46944 = n46942 & ~n46943 ;
  assign n46945 = \pi0947  & ~n21678 ;
  assign n46946 = ~n21672 & n46945 ;
  assign n46947 = \pi0947  & n21660 ;
  assign n46948 = ~n21659 & n46947 ;
  assign n46949 = n6761 & ~n46948 ;
  assign n46950 = ~n46946 & n46949 ;
  assign n46951 = \pi0223  & ~n46815 ;
  assign n46952 = ~n46950 & n46951 ;
  assign n46953 = ~\pi0947  & ~n21654 ;
  assign n46954 = ~n21657 & n46953 ;
  assign n46955 = n46951 & n46954 ;
  assign n46956 = ~n21684 & n46955 ;
  assign n46957 = ~n46952 & ~n46956 ;
  assign n46958 = \pi0221  & n46957 ;
  assign n46959 = ~\pi0616  & ~n46296 ;
  assign n46960 = ~n46861 & n46959 ;
  assign n46961 = ~n46860 & n46960 ;
  assign n46962 = \pi0947  & ~n46961 ;
  assign n46963 = \pi0947  & ~n46962 ;
  assign n46964 = n21627 & ~n46962 ;
  assign n46965 = ~n21726 & n46964 ;
  assign n46966 = ~n46963 & ~n46965 ;
  assign n46967 = \pi0221  & ~n6761 ;
  assign n46968 = n46966 & n46967 ;
  assign n46969 = ~n46958 & ~n46968 ;
  assign n46970 = ~\pi0299  & n46969 ;
  assign n46971 = ~n46930 & n46970 ;
  assign n46972 = ~n46944 & ~n46971 ;
  assign n46973 = ~n46937 & n46972 ;
  assign n46974 = n46875 & n46973 ;
  assign n46975 = \pi0038  & ~n46944 ;
  assign n46976 = ~n21205 & n46904 ;
  assign n46977 = ~n21238 & n46976 ;
  assign n46978 = \pi0221  & \pi0299  ;
  assign n46979 = ~n26957 & ~n46978 ;
  assign n46980 = n21237 & ~n46978 ;
  assign n46981 = n21232 & n46980 ;
  assign n46982 = ~n46979 & ~n46981 ;
  assign n46983 = ~n46977 & n46982 ;
  assign n46984 = ~n21740 & n46904 ;
  assign n46985 = ~n21738 & n46984 ;
  assign n46986 = \pi0221  & ~\pi0299  ;
  assign n46987 = ~n27218 & ~n46986 ;
  assign n46988 = n21737 & ~n46986 ;
  assign n46989 = n21232 & n46988 ;
  assign n46990 = ~n46987 & ~n46989 ;
  assign n46991 = ~n46985 & n46990 ;
  assign n46992 = ~n46983 & ~n46991 ;
  assign n46993 = ~\pi0039  & ~n46944 ;
  assign n46994 = ~n46992 & n46993 ;
  assign n46995 = ~n46975 & ~n46994 ;
  assign n46996 = n11834 & n46995 ;
  assign n46997 = ~n46974 & n46996 ;
  assign n46998 = ~\pi0221  & ~n46110 ;
  assign n46999 = ~n46997 & ~n46998 ;
  assign n47000 = \pi0222  & n21768 ;
  assign n47001 = n20985 & n47000 ;
  assign n47002 = ~\pi0223  & n21612 ;
  assign n47003 = ~n21606 & n47002 ;
  assign n47004 = \pi0039  & n21688 ;
  assign n47005 = ~n47003 & n47004 ;
  assign n47006 = ~n2297 & ~n47005 ;
  assign n47007 = n25541 & ~n47006 ;
  assign n47008 = ~\pi0038  & \pi0222  ;
  assign n47009 = n21743 & n47008 ;
  assign n47010 = n20985 & n47009 ;
  assign n47011 = ~n47007 & n47010 ;
  assign n47012 = ~n47001 & ~n47011 ;
  assign n47013 = ~n25588 & n47012 ;
  assign n47014 = ~n47007 & n47009 ;
  assign n47015 = n21776 & ~n47000 ;
  assign n47016 = ~n47014 & n47015 ;
  assign n47017 = ~\pi0781  & ~n47016 ;
  assign n47018 = ~n47013 & n47017 ;
  assign n47019 = \pi0222  & n21272 ;
  assign n47020 = \pi0299  & ~\pi0616  ;
  assign n47021 = n21474 & n47020 ;
  assign n47022 = ~n21472 & n47021 ;
  assign n47023 = ~\pi0299  & ~\pi0616  ;
  assign n47024 = n21481 & n47023 ;
  assign n47025 = n21477 & n47023 ;
  assign n47026 = ~n21263 & n47025 ;
  assign n47027 = ~n47024 & ~n47026 ;
  assign n47028 = ~n47022 & n47027 ;
  assign n47029 = ~\pi0222  & \pi0299  ;
  assign n47030 = ~n21475 & n47029 ;
  assign n47031 = ~\pi0222  & ~\pi0299  ;
  assign n47032 = ~n21481 & n47031 ;
  assign n47033 = ~n21478 & n47032 ;
  assign n47034 = ~\pi0039  & ~n47033 ;
  assign n47035 = ~n47030 & n47034 ;
  assign n47036 = n47028 & n47035 ;
  assign n47037 = ~n47019 & n47036 ;
  assign n47038 = ~\pi0038  & ~n47037 ;
  assign n47039 = \pi0222  & ~n21757 ;
  assign n47040 = \pi0603  & \pi0616  ;
  assign n47041 = ~n20783 & n47040 ;
  assign n47042 = n1689 & n47041 ;
  assign n47043 = n8413 & n47042 ;
  assign n47044 = n1354 & n47043 ;
  assign n47045 = n1358 & n47044 ;
  assign n47046 = \pi0038  & ~n47045 ;
  assign n47047 = ~n47039 & n47046 ;
  assign n47048 = n6861 & ~n47047 ;
  assign n47049 = ~n47038 & n47048 ;
  assign n47050 = \pi0222  & ~n6861 ;
  assign n47051 = \pi0616  & ~n1689 ;
  assign n47052 = ~n47041 & ~n47051 ;
  assign n47053 = ~n21639 & n47052 ;
  assign n47054 = ~n21615 & n47053 ;
  assign n47055 = ~n21645 & n47054 ;
  assign n47056 = n6707 & n47052 ;
  assign n47057 = ~n22183 & n47056 ;
  assign n47058 = n6708 & ~n47057 ;
  assign n47059 = ~n47055 & n47058 ;
  assign n47060 = ~n21615 & n47052 ;
  assign n47061 = ~n21645 & n47060 ;
  assign n47062 = ~n6708 & ~n47061 ;
  assign n47063 = ~n6761 & ~n47062 ;
  assign n47064 = ~n47059 & n47063 ;
  assign n47065 = ~n6707 & ~n20784 ;
  assign n47066 = ~n21285 & n47065 ;
  assign n47067 = ~n21633 & ~n47066 ;
  assign n47068 = ~n46289 & ~n47067 ;
  assign n47069 = n6707 & ~n47041 ;
  assign n47070 = ~n21352 & n47069 ;
  assign n47071 = ~n21405 & n47070 ;
  assign n47072 = n6708 & ~n47071 ;
  assign n47073 = ~n47068 & n47072 ;
  assign n47074 = ~\pi0616  & ~n6708 ;
  assign n47075 = ~n21632 & n47074 ;
  assign n47076 = ~n21631 & n47075 ;
  assign n47077 = ~n20784 & ~n21285 ;
  assign n47078 = \pi0616  & ~n6708 ;
  assign n47079 = ~n47077 & n47078 ;
  assign n47080 = n6761 & ~n47079 ;
  assign n47081 = ~n47076 & n47080 ;
  assign n47082 = ~n47073 & n47081 ;
  assign n47083 = \pi0222  & ~n47082 ;
  assign n47084 = ~n47064 & n47083 ;
  assign n47085 = ~n6706 & n6708 ;
  assign n47086 = n6707 & n47085 ;
  assign n47087 = n21403 & n47086 ;
  assign n47088 = ~n21399 & n47087 ;
  assign n47089 = ~\pi0222  & \pi0616  ;
  assign n47090 = n20784 & n47089 ;
  assign n47091 = ~n21285 & n47090 ;
  assign n47092 = ~n47088 & n47091 ;
  assign n47093 = ~n22079 & n47092 ;
  assign n47094 = \pi0223  & ~n47093 ;
  assign n47095 = ~\pi0299  & n47094 ;
  assign n47096 = ~n47084 & n47095 ;
  assign n47097 = \pi0039  & ~n47096 ;
  assign n47098 = ~n21346 & n47069 ;
  assign n47099 = n6707 & n20783 ;
  assign n47100 = ~n21290 & n47099 ;
  assign n47101 = ~n21325 & n47100 ;
  assign n47102 = n6708 & ~n47101 ;
  assign n47103 = ~n47098 & n47102 ;
  assign n47104 = n6707 & n47103 ;
  assign n47105 = ~\pi0616  & ~n21328 ;
  assign n47106 = ~\pi0616  & n46827 ;
  assign n47107 = ~n46826 & n47106 ;
  assign n47108 = ~n47105 & ~n47107 ;
  assign n47109 = \pi0616  & ~n20784 ;
  assign n47110 = ~n21339 & n47109 ;
  assign n47111 = ~n21337 & n47110 ;
  assign n47112 = n47103 & ~n47111 ;
  assign n47113 = n47108 & n47112 ;
  assign n47114 = ~n47104 & ~n47113 ;
  assign n47115 = ~n6708 & ~n47111 ;
  assign n47116 = n47108 & n47115 ;
  assign n47117 = ~n6761 & ~n47116 ;
  assign n47118 = n47114 & n47117 ;
  assign n47119 = ~n21359 & n47069 ;
  assign n47120 = n6708 & ~n47119 ;
  assign n47121 = \pi0616  & ~n47077 ;
  assign n47122 = \pi0616  & ~n47121 ;
  assign n47123 = ~n21577 & ~n47121 ;
  assign n47124 = ~n21576 & n47123 ;
  assign n47125 = ~n47122 & ~n47124 ;
  assign n47126 = ~n6707 & ~n47125 ;
  assign n47127 = n47120 & ~n47126 ;
  assign n47128 = ~n6708 & n47125 ;
  assign n47129 = n6761 & ~n47128 ;
  assign n47130 = ~n47127 & n47129 ;
  assign n47131 = \pi0222  & ~n47130 ;
  assign n47132 = ~n47118 & n47131 ;
  assign n47133 = ~n6707 & n47041 ;
  assign n47134 = ~n21329 & n47133 ;
  assign n47135 = n44606 & n47040 ;
  assign n47136 = ~n21346 & n47135 ;
  assign n47137 = n6708 & ~n47136 ;
  assign n47138 = ~n47134 & n47137 ;
  assign n47139 = ~n6708 & ~n21286 ;
  assign n47140 = n21328 & n47139 ;
  assign n47141 = ~n6708 & ~n47041 ;
  assign n47142 = ~n6761 & ~n47141 ;
  assign n47143 = ~n47140 & n47142 ;
  assign n47144 = ~n47138 & n47143 ;
  assign n47145 = ~n6709 & ~n21516 ;
  assign n47146 = n46416 & ~n47145 ;
  assign n47147 = ~n21487 & n47146 ;
  assign n47148 = \pi0224  & ~n47147 ;
  assign n47149 = ~n47144 & n47148 ;
  assign n47150 = ~n21285 & n47041 ;
  assign n47151 = ~\pi0224  & ~n47150 ;
  assign n47152 = ~\pi0222  & ~n47151 ;
  assign n47153 = ~n47149 & n47152 ;
  assign n47154 = n43384 & ~n47153 ;
  assign n47155 = ~n47132 & n47154 ;
  assign n47156 = \pi0616  & n6709 ;
  assign n47157 = \pi0616  & n20784 ;
  assign n47158 = ~n21285 & n47157 ;
  assign n47159 = ~n47156 & ~n47158 ;
  assign n47160 = ~n6709 & ~n47159 ;
  assign n47161 = n20784 & ~n47159 ;
  assign n47162 = ~n21359 & n47161 ;
  assign n47163 = ~n47160 & ~n47162 ;
  assign n47164 = n6732 & n47163 ;
  assign n47165 = ~\pi0222  & n6732 ;
  assign n47166 = ~n47140 & ~n47141 ;
  assign n47167 = ~\pi0222  & n47166 ;
  assign n47168 = ~n47138 & n47167 ;
  assign n47169 = ~n47165 & ~n47168 ;
  assign n47170 = ~n47164 & ~n47169 ;
  assign n47171 = ~n6732 & ~n47062 ;
  assign n47172 = ~n47059 & n47171 ;
  assign n47173 = ~n47076 & ~n47079 ;
  assign n47174 = n6732 & n47173 ;
  assign n47175 = ~n47073 & n47174 ;
  assign n47176 = \pi0215  & \pi0222  ;
  assign n47177 = ~n47175 & n47176 ;
  assign n47178 = ~n47172 & n47177 ;
  assign n47179 = \pi0215  & n47091 ;
  assign n47180 = ~n47088 & n47179 ;
  assign n47181 = ~n22055 & n47180 ;
  assign n47182 = \pi0299  & ~n47181 ;
  assign n47183 = ~n47178 & n47182 ;
  assign n47184 = ~\pi0216  & ~\pi0221  ;
  assign n47185 = n47183 & ~n47184 ;
  assign n47186 = ~n47170 & n47185 ;
  assign n47187 = \pi0222  & n21285 ;
  assign n47188 = n2352 & ~n47187 ;
  assign n47189 = ~n47150 & n47188 ;
  assign n47190 = ~\pi0215  & ~n47189 ;
  assign n47191 = n47182 & ~n47190 ;
  assign n47192 = ~n47178 & n47191 ;
  assign n47193 = n47048 & ~n47192 ;
  assign n47194 = ~n47186 & n47193 ;
  assign n47195 = n6732 & ~n47128 ;
  assign n47196 = ~n47127 & n47195 ;
  assign n47197 = \pi0222  & ~n47196 ;
  assign n47198 = ~n6732 & ~n47116 ;
  assign n47199 = n47114 & n47198 ;
  assign n47200 = n47193 & ~n47199 ;
  assign n47201 = n47197 & n47200 ;
  assign n47202 = ~n47194 & ~n47201 ;
  assign n47203 = ~n47155 & ~n47202 ;
  assign n47204 = n47097 & n47203 ;
  assign n47205 = ~n47050 & ~n47204 ;
  assign n47206 = ~n47049 & n47205 ;
  assign n47207 = ~n20985 & n47017 ;
  assign n47208 = ~n47206 & n47207 ;
  assign n47209 = ~n47018 & ~n47208 ;
  assign n47210 = ~\pi0619  & n47209 ;
  assign n47211 = \pi0619  & ~n47000 ;
  assign n47212 = ~n47014 & n47211 ;
  assign n47213 = ~\pi1159  & ~n47212 ;
  assign n47214 = ~n47210 & n47213 ;
  assign n47215 = ~n47000 & ~n47014 ;
  assign n47216 = \pi0618  & ~\pi1154  ;
  assign n47217 = ~n47215 & n47216 ;
  assign n47218 = \pi0618  & ~n47000 ;
  assign n47219 = ~n47014 & n47218 ;
  assign n47220 = ~\pi1154  & ~n47219 ;
  assign n47221 = ~n47016 & n47220 ;
  assign n47222 = ~n47217 & ~n47221 ;
  assign n47223 = ~n20985 & ~n47206 ;
  assign n47224 = n47013 & ~n47217 ;
  assign n47225 = ~n47223 & n47224 ;
  assign n47226 = ~n47222 & ~n47225 ;
  assign n47227 = ~\pi0618  & \pi1154  ;
  assign n47228 = ~n47215 & n47227 ;
  assign n47229 = ~\pi0618  & ~n47000 ;
  assign n47230 = ~n47014 & n47229 ;
  assign n47231 = \pi1154  & ~n47230 ;
  assign n47232 = ~n47016 & n47231 ;
  assign n47233 = ~n47228 & ~n47232 ;
  assign n47234 = n47013 & ~n47228 ;
  assign n47235 = ~n47223 & n47234 ;
  assign n47236 = ~n47233 & ~n47235 ;
  assign n47237 = ~n47226 & ~n47236 ;
  assign n47238 = \pi0781  & n47213 ;
  assign n47239 = ~n47237 & n47238 ;
  assign n47240 = ~n47214 & ~n47239 ;
  assign n47241 = \pi0619  & n47209 ;
  assign n47242 = ~\pi0619  & ~n47000 ;
  assign n47243 = ~n47014 & n47242 ;
  assign n47244 = \pi1159  & ~n47243 ;
  assign n47245 = ~n47241 & n47244 ;
  assign n47246 = \pi0781  & n47244 ;
  assign n47247 = ~n47237 & n47246 ;
  assign n47248 = ~n47245 & ~n47247 ;
  assign n47249 = n47240 & n47248 ;
  assign n47250 = n39235 & ~n47249 ;
  assign n47251 = ~\pi0789  & ~n47209 ;
  assign n47252 = ~n23880 & n47251 ;
  assign n47253 = n39241 & ~n47237 ;
  assign n47254 = ~n47252 & ~n47253 ;
  assign n47255 = \pi0661  & n1689 ;
  assign n47256 = n20855 & n47255 ;
  assign n47257 = n8413 & n47256 ;
  assign n47258 = n1354 & n47257 ;
  assign n47259 = n1358 & n47258 ;
  assign n47260 = \pi0038  & ~n47259 ;
  assign n47261 = ~n47039 & n47260 ;
  assign n47262 = n6861 & ~n47261 ;
  assign n47263 = ~\pi0222  & \pi0625  ;
  assign n47264 = ~n22727 & ~n47263 ;
  assign n47265 = ~n47262 & ~n47264 ;
  assign n47266 = ~\pi0661  & \pi0681  ;
  assign n47267 = n21580 & n47266 ;
  assign n47268 = n21359 & n44606 ;
  assign n47269 = \pi0616  & ~n47268 ;
  assign n47270 = ~n21577 & ~n47268 ;
  assign n47271 = ~n21576 & n47270 ;
  assign n47272 = ~n47269 & ~n47271 ;
  assign n47273 = ~n21570 & ~n47272 ;
  assign n47274 = ~n21359 & n44606 ;
  assign n47275 = n6708 & ~n47274 ;
  assign n47276 = ~n47273 & n47275 ;
  assign n47277 = ~n47267 & ~n47276 ;
  assign n47278 = ~n21889 & n21892 ;
  assign n47279 = \pi0661  & n47278 ;
  assign n47280 = \pi0616  & ~n21570 ;
  assign n47281 = ~n21570 & ~n21577 ;
  assign n47282 = ~n21576 & n47281 ;
  assign n47283 = ~n47280 & ~n47282 ;
  assign n47284 = \pi0661  & ~\pi0680  ;
  assign n47285 = n47283 & n47284 ;
  assign n47286 = ~n47279 & ~n47285 ;
  assign n47287 = n6761 & n47286 ;
  assign n47288 = n47277 & n47287 ;
  assign n47289 = \pi0661  & ~n21972 ;
  assign n47290 = ~n21970 & n47289 ;
  assign n47291 = ~n21672 & n47290 ;
  assign n47292 = n6761 & n47291 ;
  assign n47293 = ~\pi0661  & ~n21654 ;
  assign n47294 = ~n21657 & n47293 ;
  assign n47295 = n6761 & n47294 ;
  assign n47296 = ~n21684 & n47295 ;
  assign n47297 = ~n47292 & ~n47296 ;
  assign n47298 = n21954 & ~n21961 ;
  assign n47299 = \pi0661  & ~n47298 ;
  assign n47300 = ~n6706 & ~n21639 ;
  assign n47301 = ~n21637 & n47300 ;
  assign n47302 = ~n21635 & n47301 ;
  assign n47303 = n6708 & n21520 ;
  assign n47304 = ~n47302 & n47303 ;
  assign n47305 = n21615 & n47266 ;
  assign n47306 = n6711 & n47266 ;
  assign n47307 = ~n21624 & n47306 ;
  assign n47308 = ~n47305 & ~n47307 ;
  assign n47309 = ~n6761 & n47308 ;
  assign n47310 = ~n47304 & n47309 ;
  assign n47311 = ~n47299 & n47310 ;
  assign n47312 = \pi0222  & ~n47311 ;
  assign n47313 = n47297 & n47312 ;
  assign n47314 = ~\pi0222  & \pi0661  ;
  assign n47315 = ~n22079 & n47314 ;
  assign n47316 = n22054 & n47315 ;
  assign n47317 = \pi0223  & ~n47316 ;
  assign n47318 = ~n47313 & n47317 ;
  assign n47319 = \pi0680  & ~n21917 ;
  assign n47320 = ~n21914 & n47319 ;
  assign n47321 = \pi0661  & ~n6761 ;
  assign n47322 = ~n47320 & n47321 ;
  assign n47323 = n22274 & n47322 ;
  assign n47324 = ~\pi0661  & ~n6761 ;
  assign n47325 = ~n21334 & n47324 ;
  assign n47326 = n6713 & n47324 ;
  assign n47327 = ~n21329 & n47326 ;
  assign n47328 = ~n47325 & ~n47327 ;
  assign n47329 = ~n47323 & n47328 ;
  assign n47330 = \pi0222  & n47329 ;
  assign n47331 = ~n47318 & n47330 ;
  assign n47332 = ~n47288 & n47331 ;
  assign n47333 = \pi0661  & \pi0680  ;
  assign n47334 = ~n20854 & n47333 ;
  assign n47335 = ~n21285 & n47334 ;
  assign n47336 = ~\pi0224  & ~n47335 ;
  assign n47337 = ~\pi0222  & ~n47336 ;
  assign n47338 = ~\pi0223  & ~n47337 ;
  assign n47339 = \pi0661  & n20855 ;
  assign n47340 = ~n21905 & n47339 ;
  assign n47341 = ~n22039 & n47340 ;
  assign n47342 = ~n6761 & n47341 ;
  assign n47343 = \pi0224  & ~n47342 ;
  assign n47344 = n6761 & n47333 ;
  assign n47345 = n22030 & n47344 ;
  assign n47346 = ~n22025 & n47344 ;
  assign n47347 = n22033 & n47346 ;
  assign n47348 = ~n47345 & ~n47347 ;
  assign n47349 = ~\pi0223  & n47348 ;
  assign n47350 = n47343 & n47349 ;
  assign n47351 = ~n47338 & ~n47350 ;
  assign n47352 = ~n47318 & n47351 ;
  assign n47353 = ~\pi0299  & ~n47352 ;
  assign n47354 = ~n47332 & n47353 ;
  assign n47355 = \pi0039  & ~n47354 ;
  assign n47356 = n47188 & ~n47335 ;
  assign n47357 = ~\pi0215  & ~n47356 ;
  assign n47358 = n22030 & n47333 ;
  assign n47359 = ~n22025 & n47333 ;
  assign n47360 = n22033 & n47359 ;
  assign n47361 = ~n47358 & ~n47360 ;
  assign n47362 = n6732 & n47361 ;
  assign n47363 = ~n6732 & ~n47341 ;
  assign n47364 = ~\pi0222  & ~n47363 ;
  assign n47365 = ~n47362 & n47364 ;
  assign n47366 = ~n2352 & ~n47365 ;
  assign n47367 = n47357 & ~n47366 ;
  assign n47368 = n6732 & n47286 ;
  assign n47369 = n47277 & n47368 ;
  assign n47370 = ~\pi0661  & ~n6732 ;
  assign n47371 = ~n21334 & n47370 ;
  assign n47372 = n6713 & n47370 ;
  assign n47373 = ~n21329 & n47372 ;
  assign n47374 = ~n47371 & ~n47373 ;
  assign n47375 = \pi0661  & ~n6732 ;
  assign n47376 = ~n47320 & n47375 ;
  assign n47377 = n22274 & n47376 ;
  assign n47378 = \pi0222  & ~n47377 ;
  assign n47379 = n47374 & n47378 ;
  assign n47380 = n47357 & n47379 ;
  assign n47381 = ~n47369 & n47380 ;
  assign n47382 = ~n47367 & ~n47381 ;
  assign n47383 = n6732 & n47291 ;
  assign n47384 = n6732 & n47294 ;
  assign n47385 = ~n21684 & n47384 ;
  assign n47386 = ~n47383 & ~n47385 ;
  assign n47387 = ~n6732 & n47308 ;
  assign n47388 = ~n47304 & n47387 ;
  assign n47389 = ~n47299 & n47388 ;
  assign n47390 = \pi0222  & ~n47389 ;
  assign n47391 = n47386 & n47390 ;
  assign n47392 = ~n22055 & n47314 ;
  assign n47393 = n22054 & n47392 ;
  assign n47394 = \pi0299  & ~n47393 ;
  assign n47395 = ~n47391 & n47394 ;
  assign n47396 = ~n21948 & ~n47395 ;
  assign n47397 = n47382 & ~n47396 ;
  assign n47398 = n47355 & ~n47397 ;
  assign n47399 = ~n22102 & ~n47333 ;
  assign n47400 = ~n22101 & n47399 ;
  assign n47401 = \pi0198  & n22002 ;
  assign n47402 = ~\pi0198  & ~n21996 ;
  assign n47403 = \pi0222  & ~n47402 ;
  assign n47404 = ~n47401 & n47403 ;
  assign n47405 = ~n47400 & ~n47404 ;
  assign n47406 = ~\pi0198  & ~\pi0222  ;
  assign n47407 = n21203 & n47406 ;
  assign n47408 = ~n22096 & n47407 ;
  assign n47409 = \pi0198  & ~\pi0222  ;
  assign n47410 = n21236 & n47409 ;
  assign n47411 = n22094 & n47410 ;
  assign n47412 = ~n47408 & ~n47411 ;
  assign n47413 = ~\pi0299  & n47412 ;
  assign n47414 = n47405 & n47413 ;
  assign n47415 = ~\pi0039  & n47414 ;
  assign n47416 = ~n22097 & ~n47333 ;
  assign n47417 = ~n22095 & n47416 ;
  assign n47418 = \pi0210  & n22002 ;
  assign n47419 = ~\pi0210  & ~n21996 ;
  assign n47420 = \pi0222  & ~n47419 ;
  assign n47421 = ~n47418 & n47420 ;
  assign n47422 = ~n47417 & ~n47421 ;
  assign n47423 = \pi0299  & n47422 ;
  assign n47424 = ~n22095 & ~n22097 ;
  assign n47425 = ~\pi0222  & ~n47424 ;
  assign n47426 = ~\pi0039  & ~n47425 ;
  assign n47427 = n47423 & n47426 ;
  assign n47428 = ~n47415 & ~n47427 ;
  assign n47429 = ~\pi0038  & n47428 ;
  assign n47430 = ~n47264 & n47429 ;
  assign n47431 = ~n47398 & n47430 ;
  assign n47432 = ~n47265 & ~n47431 ;
  assign n47433 = ~\pi0625  & ~n47000 ;
  assign n47434 = ~n47014 & n47433 ;
  assign n47435 = \pi1153  & ~n47434 ;
  assign n47436 = n47432 & n47435 ;
  assign n47437 = ~\pi0222  & ~\pi0625  ;
  assign n47438 = ~n22734 & ~n47437 ;
  assign n47439 = ~n47262 & ~n47438 ;
  assign n47440 = n47429 & ~n47438 ;
  assign n47441 = ~n47398 & n47440 ;
  assign n47442 = ~n47439 & ~n47441 ;
  assign n47443 = \pi0625  & ~n47000 ;
  assign n47444 = ~n47014 & n47443 ;
  assign n47445 = ~\pi1153  & ~n47444 ;
  assign n47446 = n47442 & n47445 ;
  assign n47447 = ~n47436 & ~n47446 ;
  assign n47448 = n26065 & ~n47447 ;
  assign n47449 = ~n47050 & ~n47262 ;
  assign n47450 = ~n47050 & n47429 ;
  assign n47451 = ~n47398 & n47450 ;
  assign n47452 = ~n47449 & ~n47451 ;
  assign n47453 = n26739 & n47452 ;
  assign n47454 = ~n23885 & n47000 ;
  assign n47455 = ~n23885 & n47009 ;
  assign n47456 = ~n47007 & n47455 ;
  assign n47457 = ~n47454 & ~n47456 ;
  assign n47458 = ~\pi0628  & n47457 ;
  assign n47459 = ~n47453 & n47458 ;
  assign n47460 = ~n47448 & n47459 ;
  assign n47461 = \pi0628  & ~n47000 ;
  assign n47462 = ~n47014 & n47461 ;
  assign n47463 = n20844 & ~n47462 ;
  assign n47464 = ~n47460 & n47463 ;
  assign n47465 = \pi0628  & n47457 ;
  assign n47466 = ~n47453 & n47465 ;
  assign n47467 = ~n47448 & n47466 ;
  assign n47468 = ~\pi0628  & ~n47000 ;
  assign n47469 = ~n47014 & n47468 ;
  assign n47470 = n20843 & ~n47469 ;
  assign n47471 = ~n47467 & n47470 ;
  assign n47472 = ~n47464 & ~n47471 ;
  assign n47473 = n23880 & n47000 ;
  assign n47474 = n23880 & n47009 ;
  assign n47475 = ~n47007 & n47474 ;
  assign n47476 = ~n47473 & ~n47475 ;
  assign n47477 = n47472 & n47476 ;
  assign n47478 = n47254 & n47477 ;
  assign n47479 = ~n47250 & n47478 ;
  assign n47480 = ~n24691 & n47472 ;
  assign n47481 = n24724 & ~n47480 ;
  assign n47482 = ~n47479 & n47481 ;
  assign n47483 = ~\pi0609  & n47012 ;
  assign n47484 = \pi0609  & ~n47000 ;
  assign n47485 = ~n47014 & n47484 ;
  assign n47486 = n20865 & ~n47485 ;
  assign n47487 = ~n47483 & n47486 ;
  assign n47488 = ~n20985 & n47486 ;
  assign n47489 = ~n47206 & n47488 ;
  assign n47490 = ~n47487 & ~n47489 ;
  assign n47491 = ~n26119 & ~n47447 ;
  assign n47492 = n26125 & n47452 ;
  assign n47493 = \pi0609  & n47012 ;
  assign n47494 = ~\pi0609  & ~n47000 ;
  assign n47495 = ~n47014 & n47494 ;
  assign n47496 = n20864 & ~n47495 ;
  assign n47497 = ~n47493 & n47496 ;
  assign n47498 = ~n20985 & n47496 ;
  assign n47499 = ~n47206 & n47498 ;
  assign n47500 = ~n47497 & ~n47499 ;
  assign n47501 = ~n47492 & n47500 ;
  assign n47502 = ~n47491 & n47501 ;
  assign n47503 = n47490 & n47502 ;
  assign n47504 = \pi0785  & ~n21021 ;
  assign n47505 = ~n21018 & n47504 ;
  assign n47506 = ~n47503 & n47505 ;
  assign n47507 = \pi0222  & ~n6761 ;
  assign n47508 = n47125 & n47266 ;
  assign n47509 = ~n47127 & ~n47508 ;
  assign n47510 = ~\pi0680  & ~n47125 ;
  assign n47511 = ~\pi0616  & \pi0680  ;
  assign n47512 = \pi0680  & n22276 ;
  assign n47513 = ~n21285 & n47512 ;
  assign n47514 = ~n47511 & ~n47513 ;
  assign n47515 = ~n22265 & ~n47514 ;
  assign n47516 = ~n22262 & n47515 ;
  assign n47517 = \pi0661  & ~n47516 ;
  assign n47518 = ~n47510 & n47517 ;
  assign n47519 = \pi0222  & ~n47518 ;
  assign n47520 = n47509 & n47519 ;
  assign n47521 = ~n47507 & ~n47520 ;
  assign n47522 = ~n47041 & n47266 ;
  assign n47523 = ~n21286 & n47266 ;
  assign n47524 = n21328 & n47523 ;
  assign n47525 = ~n47522 & ~n47524 ;
  assign n47526 = \pi0616  & ~n21286 ;
  assign n47527 = n21328 & n47526 ;
  assign n47528 = ~n22023 & n47109 ;
  assign n47529 = ~n21306 & n47528 ;
  assign n47530 = ~n22022 & n47529 ;
  assign n47531 = \pi0680  & ~n47530 ;
  assign n47532 = ~n47527 & n47531 ;
  assign n47533 = n47525 & n47532 ;
  assign n47534 = ~n47138 & n47533 ;
  assign n47535 = ~n22308 & n47534 ;
  assign n47536 = ~\pi0680  & n47041 ;
  assign n47537 = ~n21329 & n47536 ;
  assign n47538 = \pi0661  & ~n47537 ;
  assign n47539 = ~n47138 & ~n47538 ;
  assign n47540 = n47525 & n47539 ;
  assign n47541 = ~n21285 & n22218 ;
  assign n47542 = ~\pi0616  & n47333 ;
  assign n47543 = ~n47541 & n47542 ;
  assign n47544 = ~n21285 & ~n22276 ;
  assign n47545 = \pi0616  & n47333 ;
  assign n47546 = ~n47544 & n47545 ;
  assign n47547 = ~n47543 & ~n47546 ;
  assign n47548 = ~n47150 & ~n47333 ;
  assign n47549 = ~\pi0224  & ~n47548 ;
  assign n47550 = n47547 & n47549 ;
  assign n47551 = ~\pi0222  & ~n47550 ;
  assign n47552 = ~n6761 & n47551 ;
  assign n47553 = ~n47540 & n47552 ;
  assign n47554 = ~n47535 & n47553 ;
  assign n47555 = \pi0616  & ~\pi0681  ;
  assign n47556 = n6707 & n47555 ;
  assign n47557 = n20784 & n47556 ;
  assign n47558 = ~n21352 & n47557 ;
  assign n47559 = ~n6706 & ~n21306 ;
  assign n47560 = ~n21903 & n47559 ;
  assign n47561 = n47558 & ~n47560 ;
  assign n47562 = ~\pi0661  & ~n47150 ;
  assign n47563 = ~n6709 & ~n47562 ;
  assign n47564 = n6761 & ~n47563 ;
  assign n47565 = ~n47561 & n47564 ;
  assign n47566 = \pi0224  & ~n47565 ;
  assign n47567 = n47551 & ~n47566 ;
  assign n47568 = \pi0616  & ~n47544 ;
  assign n47569 = \pi0680  & ~n47568 ;
  assign n47570 = ~n22341 & n47569 ;
  assign n47571 = ~\pi0680  & ~n20783 ;
  assign n47572 = n47040 & n47571 ;
  assign n47573 = ~n21285 & n47572 ;
  assign n47574 = \pi0661  & n6761 ;
  assign n47575 = ~n47573 & n47574 ;
  assign n47576 = n47551 & n47575 ;
  assign n47577 = ~n47570 & n47576 ;
  assign n47578 = ~n47567 & ~n47577 ;
  assign n47579 = ~\pi0223  & n47578 ;
  assign n47580 = ~n47554 & n47579 ;
  assign n47581 = n47521 & n47580 ;
  assign n47582 = ~n47111 & n47266 ;
  assign n47583 = n47108 & n47582 ;
  assign n47584 = n47114 & ~n47583 ;
  assign n47585 = ~n20783 & n43424 ;
  assign n47586 = ~n21329 & n47585 ;
  assign n47587 = ~\pi0603  & ~n20854 ;
  assign n47588 = ~n21327 & n21336 ;
  assign n47589 = ~n47587 & ~n47588 ;
  assign n47590 = ~\pi0642  & ~n22242 ;
  assign n47591 = \pi0603  & ~n21306 ;
  assign n47592 = ~n21903 & n47591 ;
  assign n47593 = n47590 & ~n47592 ;
  assign n47594 = n47589 & n47593 ;
  assign n47595 = ~n21286 & ~n21327 ;
  assign n47596 = \pi0642  & n20854 ;
  assign n47597 = ~n47595 & n47596 ;
  assign n47598 = n6711 & ~n47597 ;
  assign n47599 = ~n47594 & n47598 ;
  assign n47600 = ~n47586 & n47599 ;
  assign n47601 = ~n21327 & n47526 ;
  assign n47602 = \pi0616  & ~n22276 ;
  assign n47603 = \pi0680  & ~n47602 ;
  assign n47604 = ~n47601 & n47603 ;
  assign n47605 = n20784 & ~n21329 ;
  assign n47606 = \pi0614  & ~\pi0616  ;
  assign n47607 = ~n20854 & n47606 ;
  assign n47608 = ~n21286 & n47606 ;
  assign n47609 = ~n21327 & n47608 ;
  assign n47610 = ~n47607 & ~n47609 ;
  assign n47611 = ~n47605 & ~n47610 ;
  assign n47612 = n47604 & ~n47611 ;
  assign n47613 = ~n47600 & n47612 ;
  assign n47614 = \pi0661  & ~n47111 ;
  assign n47615 = n47108 & n47614 ;
  assign n47616 = ~n47333 & ~n47615 ;
  assign n47617 = ~n47613 & ~n47616 ;
  assign n47618 = n47584 & ~n47617 ;
  assign n47619 = ~n47540 & n47551 ;
  assign n47620 = ~n47535 & n47619 ;
  assign n47621 = ~n6761 & n47579 ;
  assign n47622 = ~n47620 & n47621 ;
  assign n47623 = ~n47618 & n47622 ;
  assign n47624 = \pi0614  & ~n22219 ;
  assign n47625 = ~n47514 & ~n47624 ;
  assign n47626 = ~n22221 & n47625 ;
  assign n47627 = ~n22217 & n47626 ;
  assign n47628 = ~\pi0616  & ~\pi0680  ;
  assign n47629 = ~\pi0680  & ~n20784 ;
  assign n47630 = ~n21285 & n47629 ;
  assign n47631 = ~n47628 & ~n47630 ;
  assign n47632 = ~n46289 & ~n47631 ;
  assign n47633 = \pi0616  & \pi0680  ;
  assign n47634 = n22276 & n47633 ;
  assign n47635 = ~n21285 & n47634 ;
  assign n47636 = \pi0661  & ~n47635 ;
  assign n47637 = ~n47632 & n47636 ;
  assign n47638 = ~n47627 & n47637 ;
  assign n47639 = ~\pi0616  & n47266 ;
  assign n47640 = ~n21632 & n47639 ;
  assign n47641 = ~n21631 & n47640 ;
  assign n47642 = \pi0616  & n47266 ;
  assign n47643 = ~n47077 & n47642 ;
  assign n47644 = ~n47641 & ~n47643 ;
  assign n47645 = ~n47073 & n47644 ;
  assign n47646 = ~n47638 & n47645 ;
  assign n47647 = \pi0222  & ~n47646 ;
  assign n47648 = ~\pi0222  & n22352 ;
  assign n47649 = ~\pi0222  & n22349 ;
  assign n47650 = n21392 & n47649 ;
  assign n47651 = ~n47648 & ~n47650 ;
  assign n47652 = n47333 & ~n47651 ;
  assign n47653 = n6761 & ~n47092 ;
  assign n47654 = ~n47652 & n47653 ;
  assign n47655 = ~n47647 & n47654 ;
  assign n47656 = ~n22192 & n22197 ;
  assign n47657 = ~n22188 & n47512 ;
  assign n47658 = ~n47511 & ~n47657 ;
  assign n47659 = ~n47656 & ~n47658 ;
  assign n47660 = ~n22191 & n47659 ;
  assign n47661 = ~\pi0680  & n47052 ;
  assign n47662 = ~n21615 & n47661 ;
  assign n47663 = ~n21645 & n47662 ;
  assign n47664 = \pi0661  & ~n47663 ;
  assign n47665 = ~n47660 & n47664 ;
  assign n47666 = ~n47061 & n47266 ;
  assign n47667 = ~n47059 & ~n47666 ;
  assign n47668 = ~n47665 & n47667 ;
  assign n47669 = \pi0222  & ~n47668 ;
  assign n47670 = ~n21516 & ~n47333 ;
  assign n47671 = ~n20784 & n20854 ;
  assign n47672 = ~n21285 & ~n47671 ;
  assign n47673 = ~n47670 & n47672 ;
  assign n47674 = \pi0616  & n47673 ;
  assign n47675 = ~n21615 & n47674 ;
  assign n47676 = n21369 & ~n22356 ;
  assign n47677 = n22241 & n47542 ;
  assign n47678 = n22331 & n47542 ;
  assign n47679 = ~n21285 & n47678 ;
  assign n47680 = ~n47677 & ~n47679 ;
  assign n47681 = n21419 & ~n47680 ;
  assign n47682 = n6706 & ~n47680 ;
  assign n47683 = ~n21425 & n47682 ;
  assign n47684 = ~n47681 & ~n47683 ;
  assign n47685 = ~n47676 & ~n47684 ;
  assign n47686 = ~n47675 & ~n47685 ;
  assign n47687 = n6709 & ~n47150 ;
  assign n47688 = n6709 & n21403 ;
  assign n47689 = ~n21399 & n47688 ;
  assign n47690 = ~n47687 & ~n47689 ;
  assign n47691 = ~\pi0222  & n47690 ;
  assign n47692 = ~n47686 & n47691 ;
  assign n47693 = ~n6761 & ~n47692 ;
  assign n47694 = ~n47669 & n47693 ;
  assign n47695 = \pi0223  & ~n47694 ;
  assign n47696 = ~n47655 & n47695 ;
  assign n47697 = ~\pi0299  & ~n47696 ;
  assign n47698 = ~n47623 & n47697 ;
  assign n47699 = ~n47581 & n47698 ;
  assign n47700 = \pi0039  & ~n47699 ;
  assign n47701 = \pi0222  & ~n2352 ;
  assign n47702 = ~n47518 & n47701 ;
  assign n47703 = n47509 & n47702 ;
  assign n47704 = ~\pi0222  & ~n47563 ;
  assign n47705 = ~n47561 & n47704 ;
  assign n47706 = n6732 & ~n47705 ;
  assign n47707 = ~n2352 & ~n47706 ;
  assign n47708 = n47314 & ~n47573 ;
  assign n47709 = ~n2352 & n47708 ;
  assign n47710 = ~n47570 & n47709 ;
  assign n47711 = ~n47707 & ~n47710 ;
  assign n47712 = ~n47041 & ~n47333 ;
  assign n47713 = ~\pi0616  & n22218 ;
  assign n47714 = ~n47712 & n47713 ;
  assign n47715 = ~n21285 & n47714 ;
  assign n47716 = ~n47041 & ~n47545 ;
  assign n47717 = ~n22276 & ~n47716 ;
  assign n47718 = ~n21285 & n47717 ;
  assign n47719 = ~n47715 & ~n47718 ;
  assign n47720 = n47188 & n47719 ;
  assign n47721 = ~\pi0215  & ~n47720 ;
  assign n47722 = n47711 & n47721 ;
  assign n47723 = ~n47703 & n47722 ;
  assign n47724 = \pi0222  & ~n47583 ;
  assign n47725 = n47114 & n47724 ;
  assign n47726 = ~n47617 & n47725 ;
  assign n47727 = ~\pi0222  & ~n47540 ;
  assign n47728 = ~n47535 & n47727 ;
  assign n47729 = ~n6732 & n47721 ;
  assign n47730 = ~n47728 & n47729 ;
  assign n47731 = ~n47726 & n47730 ;
  assign n47732 = ~n47723 & ~n47731 ;
  assign n47733 = n6732 & ~n47092 ;
  assign n47734 = ~n47652 & n47733 ;
  assign n47735 = ~n47647 & n47734 ;
  assign n47736 = ~n6732 & ~n47691 ;
  assign n47737 = ~n6732 & ~n47675 ;
  assign n47738 = ~n47685 & n47737 ;
  assign n47739 = ~n47736 & ~n47738 ;
  assign n47740 = \pi0215  & n47739 ;
  assign n47741 = n47176 & ~n47668 ;
  assign n47742 = ~n47740 & ~n47741 ;
  assign n47743 = ~n47735 & ~n47742 ;
  assign n47744 = \pi0299  & ~n47743 ;
  assign n47745 = n47732 & n47744 ;
  assign n47746 = n47700 & ~n47745 ;
  assign n47747 = ~\pi0603  & n47402 ;
  assign n47748 = n21258 & n22002 ;
  assign n47749 = ~n47747 & ~n47748 ;
  assign n47750 = ~n22241 & n47749 ;
  assign n47751 = n22669 & n47750 ;
  assign n47752 = ~\pi0616  & n21481 ;
  assign n47753 = ~\pi0616  & n21477 ;
  assign n47754 = ~n21263 & n47753 ;
  assign n47755 = ~n47752 & ~n47754 ;
  assign n47756 = ~\pi0299  & n47755 ;
  assign n47757 = ~n22330 & ~n47333 ;
  assign n47758 = ~n22673 & n47757 ;
  assign n47759 = ~n22671 & n47758 ;
  assign n47760 = n22669 & n47759 ;
  assign n47761 = n47756 & ~n47760 ;
  assign n47762 = ~n47751 & n47761 ;
  assign n47763 = \pi0603  & ~\pi0616  ;
  assign n47764 = ~n21473 & n47763 ;
  assign n47765 = ~n21472 & n47764 ;
  assign n47766 = \pi0299  & ~n47765 ;
  assign n47767 = ~n21243 & n47757 ;
  assign n47768 = ~n21249 & n47767 ;
  assign n47769 = n22661 & n47768 ;
  assign n47770 = ~\pi0603  & n47419 ;
  assign n47771 = \pi0210  & ~\pi0603  ;
  assign n47772 = n22002 & n47771 ;
  assign n47773 = ~n47770 & ~n47772 ;
  assign n47774 = ~n21243 & ~n22241 ;
  assign n47775 = ~n21249 & n47774 ;
  assign n47776 = n47773 & n47775 ;
  assign n47777 = ~n47769 & ~n47776 ;
  assign n47778 = n47766 & n47777 ;
  assign n47779 = \pi0222  & ~n47778 ;
  assign n47780 = ~n47762 & n47779 ;
  assign n47781 = ~\pi0039  & \pi0222  ;
  assign n47782 = \pi0661  & n22676 ;
  assign n47783 = \pi0616  & n21481 ;
  assign n47784 = \pi0616  & n21477 ;
  assign n47785 = ~n21263 & n47784 ;
  assign n47786 = ~n47783 & ~n47785 ;
  assign n47787 = ~\pi0299  & n47786 ;
  assign n47788 = ~n47782 & n47787 ;
  assign n47789 = \pi0661  & ~n22657 ;
  assign n47790 = ~n22660 & n47789 ;
  assign n47791 = n22664 & n47790 ;
  assign n47792 = ~n21473 & n47040 ;
  assign n47793 = ~n21472 & n47792 ;
  assign n47794 = \pi0299  & ~n47793 ;
  assign n47795 = ~n47791 & n47794 ;
  assign n47796 = ~\pi0039  & ~n47795 ;
  assign n47797 = ~n47788 & n47796 ;
  assign n47798 = ~n47781 & ~n47797 ;
  assign n47799 = ~n47780 & ~n47798 ;
  assign n47800 = ~\pi0038  & ~n47799 ;
  assign n47801 = ~n47746 & n47800 ;
  assign n47802 = ~\pi0616  & ~n22232 ;
  assign n47803 = ~n47712 & ~n47802 ;
  assign n47804 = n21756 & n47803 ;
  assign n47805 = n1358 & n47804 ;
  assign n47806 = \pi0038  & ~n47805 ;
  assign n47807 = ~n47039 & n47806 ;
  assign n47808 = n1689 & n22276 ;
  assign n47809 = ~\pi0222  & ~\pi0616  ;
  assign n47810 = ~\pi0039  & \pi0616  ;
  assign n47811 = n47333 & n47810 ;
  assign n47812 = ~n47809 & ~n47811 ;
  assign n47813 = n47808 & ~n47812 ;
  assign n47814 = n1281 & n47813 ;
  assign n47815 = n1260 & n47814 ;
  assign n47816 = \pi0038  & n47815 ;
  assign n47817 = n6861 & ~n47816 ;
  assign n47818 = ~n47807 & n47817 ;
  assign n47819 = ~n47801 & n47818 ;
  assign n47820 = ~n47438 & ~n47819 ;
  assign n47821 = ~n47204 & ~n47264 ;
  assign n47822 = ~n47049 & n47821 ;
  assign n47823 = ~\pi1153  & ~n47822 ;
  assign n47824 = ~n47820 & n47823 ;
  assign n47825 = ~\pi0608  & ~n47436 ;
  assign n47826 = ~n47824 & n47825 ;
  assign n47827 = ~n47264 & ~n47819 ;
  assign n47828 = ~n47204 & ~n47438 ;
  assign n47829 = ~n47049 & n47828 ;
  assign n47830 = \pi1153  & ~n47829 ;
  assign n47831 = ~n47827 & n47830 ;
  assign n47832 = \pi0608  & ~n47446 ;
  assign n47833 = ~n47831 & n47832 ;
  assign n47834 = ~n47826 & ~n47833 ;
  assign n47835 = \pi0778  & ~n47834 ;
  assign n47836 = ~\pi0222  & ~\pi0778  ;
  assign n47837 = ~n23622 & ~n47836 ;
  assign n47838 = ~n23808 & n47837 ;
  assign n47839 = ~n23808 & n47818 ;
  assign n47840 = ~n47801 & n47839 ;
  assign n47841 = ~n47838 & ~n47840 ;
  assign n47842 = n21022 & ~n47841 ;
  assign n47843 = ~n47835 & n47842 ;
  assign n47844 = ~n47506 & ~n47843 ;
  assign n47845 = ~\pi0778  & n47452 ;
  assign n47846 = ~n22147 & ~n47845 ;
  assign n47847 = n22147 & ~n47000 ;
  assign n47848 = ~n47014 & n47847 ;
  assign n47849 = ~n47846 & ~n47848 ;
  assign n47850 = \pi0778  & ~n47848 ;
  assign n47851 = ~n47447 & n47850 ;
  assign n47852 = ~n47849 & ~n47851 ;
  assign n47853 = n23667 & ~n47852 ;
  assign n47854 = \pi0627  & n47226 ;
  assign n47855 = ~\pi0627  & n47236 ;
  assign n47856 = ~n47854 & ~n47855 ;
  assign n47857 = ~n47853 & n47856 ;
  assign n47858 = \pi0781  & ~n47857 ;
  assign n47859 = n47844 & ~n47858 ;
  assign n47860 = n29803 & ~n47859 ;
  assign n47861 = ~\pi0648  & ~n47248 ;
  assign n47862 = n23380 & ~n47845 ;
  assign n47863 = ~n23380 & ~n47000 ;
  assign n47864 = ~n47014 & n47863 ;
  assign n47865 = n21050 & ~n47864 ;
  assign n47866 = ~n47862 & n47865 ;
  assign n47867 = \pi0778  & n47865 ;
  assign n47868 = ~n47447 & n47867 ;
  assign n47869 = ~n47866 & ~n47868 ;
  assign n47870 = n20874 & ~n47212 ;
  assign n47871 = ~n47210 & n47870 ;
  assign n47872 = \pi0781  & n47870 ;
  assign n47873 = ~n47237 & n47872 ;
  assign n47874 = ~n47871 & ~n47873 ;
  assign n47875 = n47869 & n47874 ;
  assign n47876 = ~n47861 & n47875 ;
  assign n47877 = n36155 & ~n47876 ;
  assign n47878 = ~n47860 & ~n47877 ;
  assign n47879 = n30823 & ~n47878 ;
  assign n47880 = \pi0778  & ~n47447 ;
  assign n47881 = ~n22160 & n47862 ;
  assign n47882 = ~n47880 & n47881 ;
  assign n47883 = ~n26186 & ~n47000 ;
  assign n47884 = ~n47014 & n47883 ;
  assign n47885 = n20951 & ~n47884 ;
  assign n47886 = ~n47882 & n47885 ;
  assign n47887 = n21806 & ~n47237 ;
  assign n47888 = \pi0626  & ~n47251 ;
  assign n47889 = ~n47887 & n47888 ;
  assign n47890 = ~\pi0626  & ~n47000 ;
  assign n47891 = ~n47014 & n47890 ;
  assign n47892 = n20881 & ~n47891 ;
  assign n47893 = ~n47889 & n47892 ;
  assign n47894 = \pi0789  & n47892 ;
  assign n47895 = ~n47249 & n47894 ;
  assign n47896 = ~n47893 & ~n47895 ;
  assign n47897 = ~n47886 & n47896 ;
  assign n47898 = \pi0789  & ~n47249 ;
  assign n47899 = ~n47251 & ~n47887 ;
  assign n47900 = ~\pi0626  & n47899 ;
  assign n47901 = ~n47898 & n47900 ;
  assign n47902 = \pi0626  & ~n47000 ;
  assign n47903 = ~n47014 & n47902 ;
  assign n47904 = n20882 & ~n47903 ;
  assign n47905 = ~n47901 & n47904 ;
  assign n47906 = n47897 & ~n47905 ;
  assign n47907 = \pi0788  & n30823 ;
  assign n47908 = ~n47906 & n47907 ;
  assign n47909 = ~n47879 & ~n47908 ;
  assign n47910 = ~n47482 & n47909 ;
  assign n47911 = n23412 & n47000 ;
  assign n47912 = n23412 & n47009 ;
  assign n47913 = ~n47007 & n47912 ;
  assign n47914 = ~n47911 & ~n47913 ;
  assign n47915 = ~\pi0644  & ~n47914 ;
  assign n47916 = ~\pi0644  & n23413 ;
  assign n47917 = n21092 & n47916 ;
  assign n47918 = ~n47254 & n47917 ;
  assign n47919 = n39235 & n47917 ;
  assign n47920 = ~n47249 & n47919 ;
  assign n47921 = ~n47918 & ~n47920 ;
  assign n47922 = ~n47915 & n47921 ;
  assign n47923 = n21092 & n23412 ;
  assign n47924 = \pi0644  & ~n47254 ;
  assign n47925 = \pi0644  & n39235 ;
  assign n47926 = ~n47249 & n47925 ;
  assign n47927 = ~n47924 & ~n47926 ;
  assign n47928 = n47923 & ~n47927 ;
  assign n47929 = n23413 & n47000 ;
  assign n47930 = n23413 & n47009 ;
  assign n47931 = ~n47007 & n47930 ;
  assign n47932 = ~n47929 & ~n47931 ;
  assign n47933 = \pi0644  & ~n47932 ;
  assign n47934 = ~n23907 & n47457 ;
  assign n47935 = ~n47453 & n47934 ;
  assign n47936 = ~n47448 & n47935 ;
  assign n47937 = n23907 & ~n47000 ;
  assign n47938 = ~n47014 & n47937 ;
  assign n47939 = n23518 & ~n47938 ;
  assign n47940 = ~n47936 & n47939 ;
  assign n47941 = ~n23414 & ~n31367 ;
  assign n47942 = n47000 & n47941 ;
  assign n47943 = n47009 & n47941 ;
  assign n47944 = ~n47007 & n47943 ;
  assign n47945 = ~n47942 & ~n47944 ;
  assign n47946 = n44853 & n47945 ;
  assign n47947 = ~n47940 & n47946 ;
  assign n47948 = ~\pi0647  & ~n47000 ;
  assign n47949 = ~n47014 & n47948 ;
  assign n47950 = \pi1157  & ~n47949 ;
  assign n47951 = ~n47938 & n47950 ;
  assign n47952 = ~n47936 & n47951 ;
  assign n47953 = n20923 & ~n47215 ;
  assign n47954 = \pi0787  & ~n47953 ;
  assign n47955 = ~n47952 & n47954 ;
  assign n47956 = \pi0647  & ~n47000 ;
  assign n47957 = ~n47014 & n47956 ;
  assign n47958 = ~\pi1157  & ~n47957 ;
  assign n47959 = ~n47938 & n47958 ;
  assign n47960 = ~n47936 & n47959 ;
  assign n47961 = n21064 & ~n47215 ;
  assign n47962 = n47945 & ~n47961 ;
  assign n47963 = ~n47960 & n47962 ;
  assign n47964 = n47955 & n47963 ;
  assign n47965 = ~n47947 & ~n47964 ;
  assign n47966 = ~n47933 & ~n47965 ;
  assign n47967 = ~n47928 & n47966 ;
  assign n47968 = n47922 & n47967 ;
  assign n47969 = \pi0790  & ~n47968 ;
  assign n47970 = ~\pi0630  & n47953 ;
  assign n47971 = ~\pi0630  & n47951 ;
  assign n47972 = ~n47936 & n47971 ;
  assign n47973 = ~n47970 & ~n47972 ;
  assign n47974 = \pi0630  & n47961 ;
  assign n47975 = \pi0630  & n47959 ;
  assign n47976 = ~n47936 & n47975 ;
  assign n47977 = ~n47974 & ~n47976 ;
  assign n47978 = n47973 & n47977 ;
  assign n47979 = \pi0787  & ~n47978 ;
  assign n47980 = ~n20846 & n47476 ;
  assign n47981 = n47254 & n47980 ;
  assign n47982 = ~n47250 & n47981 ;
  assign n47983 = n20846 & ~n47000 ;
  assign n47984 = ~n47014 & n47983 ;
  assign n47985 = ~n24996 & ~n47984 ;
  assign n47986 = ~n47982 & n47985 ;
  assign n47987 = ~n47979 & ~n47986 ;
  assign n47988 = ~n47969 & n47987 ;
  assign n47989 = n47910 & n47988 ;
  assign n47990 = n24761 & n47922 ;
  assign n47991 = n47967 & n47990 ;
  assign n47992 = n9948 & ~n47991 ;
  assign n47993 = ~n47989 & n47992 ;
  assign n47994 = \pi0222  & ~n27408 ;
  assign n47995 = ~n47993 & ~n47994 ;
  assign n47996 = \pi0223  & ~n27408 ;
  assign n47997 = ~n9948 & ~n47996 ;
  assign n47998 = \pi0223  & ~\pi0778  ;
  assign n47999 = ~n6861 & n47998 ;
  assign n48000 = \pi0680  & \pi0681  ;
  assign n48001 = n2165 & ~n20854 ;
  assign n48002 = n48000 & n48001 ;
  assign n48003 = ~n21285 & n48002 ;
  assign n48004 = ~\pi0223  & ~n48003 ;
  assign n48005 = \pi0681  & n20855 ;
  assign n48006 = ~n21905 & n48005 ;
  assign n48007 = ~n22039 & n48006 ;
  assign n48008 = ~n6761 & n48007 ;
  assign n48009 = ~n2165 & n48008 ;
  assign n48010 = \pi0680  & n22030 ;
  assign n48011 = \pi0680  & ~n22025 ;
  assign n48012 = n22033 & n48011 ;
  assign n48013 = ~n48010 & ~n48012 ;
  assign n48014 = \pi0681  & n6761 ;
  assign n48015 = ~n2165 & n48014 ;
  assign n48016 = ~n48013 & n48015 ;
  assign n48017 = ~n48009 & ~n48016 ;
  assign n48018 = n48004 & n48017 ;
  assign n48019 = \pi0681  & ~n47298 ;
  assign n48020 = ~n21726 & ~n48019 ;
  assign n48021 = ~n6761 & ~n48020 ;
  assign n48022 = n6761 & n21668 ;
  assign n48023 = ~n21661 & n48022 ;
  assign n48024 = n21683 & n48023 ;
  assign n48025 = ~n21970 & ~n21972 ;
  assign n48026 = ~n21672 & n48025 ;
  assign n48027 = n48014 & ~n48026 ;
  assign n48028 = \pi0223  & ~n48027 ;
  assign n48029 = ~n48024 & n48028 ;
  assign n48030 = ~n48021 & n48029 ;
  assign n48031 = n27982 & ~n48030 ;
  assign n48032 = ~n48018 & n48031 ;
  assign n48033 = n6732 & n21593 ;
  assign n48034 = n6732 & ~n21602 ;
  assign n48035 = ~n21599 & n48034 ;
  assign n48036 = ~n48033 & ~n48035 ;
  assign n48037 = n22274 & ~n47320 ;
  assign n48038 = \pi0681  & ~n48037 ;
  assign n48039 = ~\pi0661  & n6707 ;
  assign n48040 = ~n21905 & ~n48039 ;
  assign n48041 = ~n22039 & n48040 ;
  assign n48042 = n21306 & n48039 ;
  assign n48043 = ~n21290 & n48039 ;
  assign n48044 = ~n21325 & n48043 ;
  assign n48045 = ~n48042 & ~n48044 ;
  assign n48046 = ~\pi0681  & n48045 ;
  assign n48047 = ~n48041 & n48046 ;
  assign n48048 = ~n6732 & ~n48047 ;
  assign n48049 = ~n48038 & n48048 ;
  assign n48050 = \pi0223  & ~n48049 ;
  assign n48051 = n48036 & n48050 ;
  assign n48052 = ~\pi0680  & n47283 ;
  assign n48053 = ~n47278 & ~n48052 ;
  assign n48054 = \pi0223  & \pi0681  ;
  assign n48055 = ~n48049 & n48054 ;
  assign n48056 = ~n48053 & n48055 ;
  assign n48057 = n22030 & n48000 ;
  assign n48058 = ~n22025 & n48000 ;
  assign n48059 = n22033 & n48058 ;
  assign n48060 = ~n48057 & ~n48059 ;
  assign n48061 = n6732 & n48060 ;
  assign n48062 = ~n6732 & ~n48007 ;
  assign n48063 = ~\pi0223  & ~n48062 ;
  assign n48064 = ~n48061 & n48063 ;
  assign n48065 = ~\pi0215  & ~n47184 ;
  assign n48066 = ~n48064 & n48065 ;
  assign n48067 = ~n48056 & n48066 ;
  assign n48068 = ~n48051 & n48067 ;
  assign n48069 = \pi0223  & n21285 ;
  assign n48070 = n2352 & ~n48069 ;
  assign n48071 = ~n20854 & n48000 ;
  assign n48072 = ~n21285 & n48071 ;
  assign n48073 = ~\pi0215  & ~n48072 ;
  assign n48074 = n48070 & n48073 ;
  assign n48075 = ~n6732 & n48020 ;
  assign n48076 = \pi0681  & ~n48026 ;
  assign n48077 = n6732 & ~n48076 ;
  assign n48078 = ~n21684 & n48077 ;
  assign n48079 = \pi0223  & ~n48078 ;
  assign n48080 = ~n48075 & n48079 ;
  assign n48081 = ~\pi0223  & \pi0681  ;
  assign n48082 = ~n22055 & n48081 ;
  assign n48083 = n22054 & n48082 ;
  assign n48084 = \pi0215  & ~n48083 ;
  assign n48085 = ~n48080 & n48084 ;
  assign n48086 = \pi0039  & \pi0299  ;
  assign n48087 = ~n48085 & n48086 ;
  assign n48088 = ~n48074 & n48087 ;
  assign n48089 = ~n48068 & n48088 ;
  assign n48090 = ~n48032 & ~n48089 ;
  assign n48091 = n21737 & n22094 ;
  assign n48092 = ~n22102 & ~n48091 ;
  assign n48093 = ~\pi0223  & ~n48092 ;
  assign n48094 = \pi0223  & ~n47402 ;
  assign n48095 = ~\pi0299  & ~n48094 ;
  assign n48096 = n21268 & n22002 ;
  assign n48097 = ~n48095 & ~n48096 ;
  assign n48098 = ~n22102 & ~n48000 ;
  assign n48099 = ~n22101 & n48098 ;
  assign n48100 = ~n48097 & ~n48099 ;
  assign n48101 = ~n48093 & n48100 ;
  assign n48102 = ~\pi0223  & ~n47424 ;
  assign n48103 = ~n22097 & ~n48000 ;
  assign n48104 = ~n22095 & n48103 ;
  assign n48105 = \pi0223  & ~n47419 ;
  assign n48106 = \pi0299  & ~n48105 ;
  assign n48107 = \pi0210  & \pi0299  ;
  assign n48108 = n22002 & n48107 ;
  assign n48109 = ~n48106 & ~n48108 ;
  assign n48110 = ~n48104 & ~n48109 ;
  assign n48111 = ~n48102 & n48110 ;
  assign n48112 = ~n48101 & ~n48111 ;
  assign n48113 = ~\pi0039  & ~n48112 ;
  assign n48114 = ~\pi0038  & ~n48113 ;
  assign n48115 = n48090 & n48114 ;
  assign n48116 = \pi0223  & ~n21757 ;
  assign n48117 = \pi0681  & n1689 ;
  assign n48118 = n20855 & n48117 ;
  assign n48119 = n8413 & n48118 ;
  assign n48120 = n1354 & n48119 ;
  assign n48121 = n1358 & n48120 ;
  assign n48122 = \pi0038  & ~n48121 ;
  assign n48123 = ~n48116 & n48122 ;
  assign n48124 = n25171 & ~n48123 ;
  assign n48125 = ~n48115 & n48124 ;
  assign n48126 = ~n47999 & ~n48125 ;
  assign n48127 = n23885 & ~n23907 ;
  assign n48128 = ~n48126 & n48127 ;
  assign n48129 = n6861 & ~n48123 ;
  assign n48130 = ~n48115 & n48129 ;
  assign n48131 = ~\pi0223  & \pi0625  ;
  assign n48132 = ~n22727 & ~n48131 ;
  assign n48133 = ~n48130 & ~n48132 ;
  assign n48134 = ~n21768 & ~n21770 ;
  assign n48135 = n2297 & ~n21768 ;
  assign n48136 = \pi0039  & ~n6761 ;
  assign n48137 = \pi0039  & n21658 ;
  assign n48138 = ~n21684 & n48137 ;
  assign n48139 = ~n48136 & ~n48138 ;
  assign n48140 = n21651 & ~n21768 ;
  assign n48141 = ~n48139 & n48140 ;
  assign n48142 = ~n48135 & ~n48141 ;
  assign n48143 = ~n21731 & ~n48142 ;
  assign n48144 = n21714 & n48143 ;
  assign n48145 = ~n48134 & ~n48144 ;
  assign n48146 = \pi0223  & \pi1153  ;
  assign n48147 = n48145 & n48146 ;
  assign n48148 = ~n24550 & ~n48147 ;
  assign n48149 = ~n48133 & ~n48148 ;
  assign n48150 = ~\pi0223  & ~\pi0625  ;
  assign n48151 = ~n22734 & ~n48150 ;
  assign n48152 = ~n48130 & ~n48151 ;
  assign n48153 = \pi0223  & ~\pi1153  ;
  assign n48154 = n48145 & n48153 ;
  assign n48155 = ~n24561 & ~n48154 ;
  assign n48156 = ~n48152 & ~n48155 ;
  assign n48157 = ~n48149 & ~n48156 ;
  assign n48158 = \pi0778  & n48127 ;
  assign n48159 = ~n48157 & n48158 ;
  assign n48160 = ~n48128 & ~n48159 ;
  assign n48161 = \pi0223  & ~n48127 ;
  assign n48162 = n48145 & n48161 ;
  assign n48163 = \pi0647  & ~n48162 ;
  assign n48164 = n48160 & n48163 ;
  assign n48165 = \pi0223  & \pi1157  ;
  assign n48166 = n48145 & n48165 ;
  assign n48167 = ~n20925 & ~n48166 ;
  assign n48168 = ~n48164 & ~n48167 ;
  assign n48169 = ~\pi0647  & ~n48162 ;
  assign n48170 = n48160 & n48169 ;
  assign n48171 = \pi0223  & ~\pi1157  ;
  assign n48172 = n48145 & n48171 ;
  assign n48173 = ~n22945 & ~n48172 ;
  assign n48174 = ~n48170 & ~n48173 ;
  assign n48175 = ~n48168 & ~n48174 ;
  assign n48176 = \pi0223  & n48145 ;
  assign n48177 = n23314 & n23317 ;
  assign n48178 = ~n47941 & ~n48177 ;
  assign n48179 = ~n48176 & ~n48178 ;
  assign n48180 = n23419 & n30376 ;
  assign n48181 = ~n48179 & ~n48180 ;
  assign n48182 = ~\pi0781  & n21776 ;
  assign n48183 = ~n48176 & n48182 ;
  assign n48184 = n20985 & ~n48176 ;
  assign n48185 = ~\pi0781  & ~n25588 ;
  assign n48186 = n48184 & n48185 ;
  assign n48187 = ~\pi0223  & \pi0642  ;
  assign n48188 = n21481 & n48187 ;
  assign n48189 = n21477 & n48187 ;
  assign n48190 = ~n21263 & n48189 ;
  assign n48191 = ~n48188 & ~n48190 ;
  assign n48192 = ~\pi0299  & n48191 ;
  assign n48193 = \pi0223  & n21266 ;
  assign n48194 = \pi0198  & \pi0223  ;
  assign n48195 = n21247 & n48194 ;
  assign n48196 = ~n48193 & ~n48195 ;
  assign n48197 = ~\pi0642  & n21481 ;
  assign n48198 = ~\pi0642  & n21477 ;
  assign n48199 = ~n21263 & n48198 ;
  assign n48200 = ~n48197 & ~n48199 ;
  assign n48201 = n21265 & n48200 ;
  assign n48202 = ~n48196 & n48201 ;
  assign n48203 = n48192 & ~n48202 ;
  assign n48204 = \pi0603  & n48187 ;
  assign n48205 = ~n21473 & n48204 ;
  assign n48206 = ~\pi0039  & n48205 ;
  assign n48207 = ~n21472 & n48206 ;
  assign n48208 = ~n21479 & ~n48207 ;
  assign n48209 = n6710 & ~n21473 ;
  assign n48210 = ~n21472 & n48209 ;
  assign n48211 = ~\pi0039  & \pi0223  ;
  assign n48212 = ~n48210 & n48211 ;
  assign n48213 = ~n21251 & n48212 ;
  assign n48214 = n48208 & ~n48213 ;
  assign n48215 = ~n48203 & ~n48214 ;
  assign n48216 = n47585 & ~n48039 ;
  assign n48217 = ~n21329 & n48216 ;
  assign n48218 = \pi0642  & ~\pi0661  ;
  assign n48219 = n44606 & n48218 ;
  assign n48220 = \pi0603  & n48219 ;
  assign n48221 = ~\pi0681  & ~n48220 ;
  assign n48222 = ~\pi0681  & ~n21306 ;
  assign n48223 = ~n21345 & n48222 ;
  assign n48224 = ~n48221 & ~n48223 ;
  assign n48225 = ~n48217 & ~n48224 ;
  assign n48226 = \pi0681  & ~n21286 ;
  assign n48227 = n21328 & n48226 ;
  assign n48228 = \pi0681  & ~n47585 ;
  assign n48229 = ~n48227 & ~n48228 ;
  assign n48230 = ~n6761 & n48229 ;
  assign n48231 = ~n48225 & n48230 ;
  assign n48232 = ~n20783 & n48220 ;
  assign n48233 = ~n21352 & n48232 ;
  assign n48234 = n21355 & n48233 ;
  assign n48235 = ~n21290 & n48233 ;
  assign n48236 = ~n21325 & n48235 ;
  assign n48237 = ~n48234 & ~n48236 ;
  assign n48238 = \pi0642  & ~n48039 ;
  assign n48239 = n20784 & n48238 ;
  assign n48240 = ~n21285 & n48239 ;
  assign n48241 = ~\pi0681  & ~n48240 ;
  assign n48242 = n48237 & n48241 ;
  assign n48243 = ~\pi0681  & n6761 ;
  assign n48244 = n6761 & n47585 ;
  assign n48245 = ~n21285 & n48244 ;
  assign n48246 = ~n48243 & ~n48245 ;
  assign n48247 = ~n48242 & ~n48246 ;
  assign n48248 = ~n46435 & ~n48247 ;
  assign n48249 = ~n48231 & n48248 ;
  assign n48250 = ~\pi0223  & ~n46435 ;
  assign n48251 = ~\pi0223  & n47585 ;
  assign n48252 = ~n21285 & n48251 ;
  assign n48253 = ~n48250 & ~n48252 ;
  assign n48254 = ~n48249 & ~n48253 ;
  assign n48255 = n1689 & ~n47585 ;
  assign n48256 = n1281 & n48255 ;
  assign n48257 = n1260 & n48256 ;
  assign n48258 = n48039 & n48257 ;
  assign n48259 = ~n21352 & n48258 ;
  assign n48260 = ~n21405 & n48259 ;
  assign n48261 = ~\pi0681  & n48039 ;
  assign n48262 = ~n48260 & n48261 ;
  assign n48263 = \pi0642  & ~n47077 ;
  assign n48264 = ~n47121 & ~n48263 ;
  assign n48265 = ~n46289 & n48264 ;
  assign n48266 = ~n6711 & ~n47585 ;
  assign n48267 = ~n21285 & n48266 ;
  assign n48268 = ~\pi0681  & ~n48267 ;
  assign n48269 = ~n48260 & n48268 ;
  assign n48270 = ~n48265 & n48269 ;
  assign n48271 = ~n48262 & ~n48270 ;
  assign n48272 = \pi0681  & ~n48267 ;
  assign n48273 = ~n48265 & n48272 ;
  assign n48274 = n6761 & ~n48273 ;
  assign n48275 = n48271 & n48274 ;
  assign n48276 = n21370 & ~n21624 ;
  assign n48277 = \pi0642  & ~n1689 ;
  assign n48278 = ~n47585 & ~n48277 ;
  assign n48279 = ~n6706 & n48278 ;
  assign n48280 = ~n21285 & n48279 ;
  assign n48281 = ~n48039 & n48280 ;
  assign n48282 = ~n48039 & n48278 ;
  assign n48283 = ~n21520 & n48282 ;
  assign n48284 = ~n48281 & ~n48283 ;
  assign n48285 = ~n48276 & ~n48284 ;
  assign n48286 = n48039 & n48278 ;
  assign n48287 = ~n21403 & n48286 ;
  assign n48288 = ~n21393 & n48286 ;
  assign n48289 = n21398 & n48288 ;
  assign n48290 = ~n48287 & ~n48289 ;
  assign n48291 = ~\pi0681  & n48290 ;
  assign n48292 = ~n48285 & n48291 ;
  assign n48293 = ~n21520 & n48278 ;
  assign n48294 = ~n48280 & ~n48293 ;
  assign n48295 = ~n48276 & ~n48294 ;
  assign n48296 = \pi0681  & ~n48295 ;
  assign n48297 = ~n6761 & ~n48296 ;
  assign n48298 = ~n48292 & n48297 ;
  assign n48299 = \pi0223  & ~n48298 ;
  assign n48300 = ~n48275 & n48299 ;
  assign n48301 = ~\pi0299  & ~n48300 ;
  assign n48302 = ~n48254 & n48301 ;
  assign n48303 = \pi0039  & ~n48302 ;
  assign n48304 = ~\pi0038  & ~n48303 ;
  assign n48305 = ~n20784 & n48238 ;
  assign n48306 = ~n21339 & n48305 ;
  assign n48307 = ~n21337 & n48306 ;
  assign n48308 = ~\pi0642  & ~n48039 ;
  assign n48309 = ~n21905 & n48308 ;
  assign n48310 = ~n22039 & n48309 ;
  assign n48311 = ~n48307 & ~n48310 ;
  assign n48312 = ~n47585 & ~n48045 ;
  assign n48313 = ~\pi0681  & ~n48312 ;
  assign n48314 = n48311 & n48313 ;
  assign n48315 = \pi0642  & \pi0681  ;
  assign n48316 = ~n21341 & n48315 ;
  assign n48317 = \pi0681  & n21905 ;
  assign n48318 = \pi0681  & n21908 ;
  assign n48319 = n21328 & n48318 ;
  assign n48320 = ~n48317 & ~n48319 ;
  assign n48321 = ~\pi0642  & ~n48320 ;
  assign n48322 = ~n48316 & ~n48321 ;
  assign n48323 = ~n6732 & n48322 ;
  assign n48324 = ~n48314 & n48323 ;
  assign n48325 = ~n21359 & ~n21371 ;
  assign n48326 = ~\pi0603  & ~n21285 ;
  assign n48327 = ~\pi0642  & ~n48267 ;
  assign n48328 = ~n48326 & n48327 ;
  assign n48329 = ~n48325 & n48328 ;
  assign n48330 = n6711 & ~n20784 ;
  assign n48331 = ~n21285 & n48330 ;
  assign n48332 = ~n43050 & ~n48331 ;
  assign n48333 = ~n48267 & n48332 ;
  assign n48334 = ~n48329 & ~n48333 ;
  assign n48335 = \pi0681  & ~n48334 ;
  assign n48336 = ~\pi0681  & n46330 ;
  assign n48337 = ~\pi0681  & ~n48039 ;
  assign n48338 = n6732 & ~n48337 ;
  assign n48339 = ~n48336 & n48338 ;
  assign n48340 = ~n21359 & n48338 ;
  assign n48341 = n21365 & n48340 ;
  assign n48342 = ~n48339 & ~n48341 ;
  assign n48343 = n6732 & ~n48039 ;
  assign n48344 = ~n48333 & n48343 ;
  assign n48345 = ~n48329 & n48344 ;
  assign n48346 = n48342 & ~n48345 ;
  assign n48347 = ~n48335 & ~n48346 ;
  assign n48348 = \pi0223  & ~n48347 ;
  assign n48349 = ~n48324 & n48348 ;
  assign n48350 = ~\pi0907  & n6729 ;
  assign n48351 = n6728 & n48350 ;
  assign n48352 = n48229 & ~n48351 ;
  assign n48353 = ~n48225 & n48352 ;
  assign n48354 = ~n21285 & n47585 ;
  assign n48355 = \pi0681  & ~n48354 ;
  assign n48356 = n48351 & ~n48355 ;
  assign n48357 = ~n48242 & n48356 ;
  assign n48358 = ~\pi0947  & ~n48357 ;
  assign n48359 = ~n48353 & n48358 ;
  assign n48360 = ~\pi0223  & ~\pi0947  ;
  assign n48361 = ~\pi0223  & n48229 ;
  assign n48362 = ~n48225 & n48361 ;
  assign n48363 = ~n48360 & ~n48362 ;
  assign n48364 = ~n48359 & ~n48363 ;
  assign n48365 = ~n47184 & ~n48364 ;
  assign n48366 = ~n48349 & n48365 ;
  assign n48367 = n2352 & ~n47585 ;
  assign n48368 = ~n21285 & n48367 ;
  assign n48369 = ~\pi0223  & n2352 ;
  assign n48370 = n21285 & n48369 ;
  assign n48371 = ~n48368 & ~n48370 ;
  assign n48372 = ~\pi0215  & n48371 ;
  assign n48373 = ~n48366 & n48372 ;
  assign n48374 = n6732 & ~n48273 ;
  assign n48375 = n48271 & n48374 ;
  assign n48376 = ~n6732 & ~n48296 ;
  assign n48377 = ~n48292 & n48376 ;
  assign n48378 = \pi0215  & \pi0223  ;
  assign n48379 = ~n48377 & n48378 ;
  assign n48380 = ~n48375 & n48379 ;
  assign n48381 = n21516 & n48219 ;
  assign n48382 = ~n21405 & n48381 ;
  assign n48383 = n48241 & ~n48382 ;
  assign n48384 = n21615 & n48291 ;
  assign n48385 = ~n48383 & ~n48384 ;
  assign n48386 = \pi0642  & n21515 ;
  assign n48387 = \pi0642  & n21516 ;
  assign n48388 = ~n21520 & n48387 ;
  assign n48389 = ~n48386 & ~n48388 ;
  assign n48390 = \pi0681  & n48389 ;
  assign n48391 = n48385 & ~n48390 ;
  assign n48392 = \pi0947  & ~n48391 ;
  assign n48393 = ~\pi0223  & ~n48392 ;
  assign n48394 = n6732 & n47585 ;
  assign n48395 = ~n21285 & n48394 ;
  assign n48396 = ~\pi0947  & ~n48395 ;
  assign n48397 = ~\pi0947  & n48241 ;
  assign n48398 = ~n48382 & n48397 ;
  assign n48399 = ~n48396 & ~n48398 ;
  assign n48400 = \pi0215  & n48399 ;
  assign n48401 = \pi0215  & ~n48351 ;
  assign n48402 = n48391 & n48401 ;
  assign n48403 = ~n48400 & ~n48402 ;
  assign n48404 = n48393 & ~n48403 ;
  assign n48405 = ~\pi0038  & \pi0299  ;
  assign n48406 = ~n48404 & n48405 ;
  assign n48407 = ~n48380 & n48406 ;
  assign n48408 = ~n48373 & n48407 ;
  assign n48409 = ~n48304 & ~n48408 ;
  assign n48410 = ~n48215 & ~n48409 ;
  assign n48411 = \pi0038  & ~n43121 ;
  assign n48412 = ~\pi0223  & ~n21289 ;
  assign n48413 = ~\pi0039  & ~n48257 ;
  assign n48414 = ~n48412 & n48413 ;
  assign n48415 = n48411 & ~n48414 ;
  assign n48416 = n6861 & ~n48415 ;
  assign n48417 = ~n48410 & n48416 ;
  assign n48418 = \pi0223  & ~n6861 ;
  assign n48419 = ~n20985 & ~n48418 ;
  assign n48420 = n48185 & n48419 ;
  assign n48421 = ~n48417 & n48420 ;
  assign n48422 = ~n48186 & ~n48421 ;
  assign n48423 = ~n48183 & n48422 ;
  assign n48424 = ~n23423 & ~n48423 ;
  assign n48425 = n20811 & ~n25588 ;
  assign n48426 = n48184 & n48425 ;
  assign n48427 = n48419 & n48425 ;
  assign n48428 = ~n48417 & n48427 ;
  assign n48429 = ~n48426 & ~n48428 ;
  assign n48430 = n20811 & n21776 ;
  assign n48431 = ~n48176 & n48430 ;
  assign n48432 = ~n20811 & ~n48176 ;
  assign n48433 = ~n48431 & ~n48432 ;
  assign n48434 = n48429 & n48433 ;
  assign n48435 = n23424 & ~n48434 ;
  assign n48436 = ~n48424 & ~n48435 ;
  assign n48437 = n23423 & ~n48176 ;
  assign n48438 = ~n48179 & ~n48437 ;
  assign n48439 = n48436 & n48438 ;
  assign n48440 = ~n48181 & ~n48439 ;
  assign n48441 = \pi0787  & ~n48440 ;
  assign n48442 = ~n48175 & n48441 ;
  assign n48443 = \pi0790  & ~n48442 ;
  assign n48444 = \pi0787  & n23518 ;
  assign n48445 = n23518 & ~n48162 ;
  assign n48446 = n48160 & n48445 ;
  assign n48447 = ~n48444 & ~n48446 ;
  assign n48448 = n48436 & ~n48437 ;
  assign n48449 = n48180 & ~n48448 ;
  assign n48450 = n48447 & ~n48449 ;
  assign n48451 = ~n48179 & n48450 ;
  assign n48452 = ~n47996 & ~n48451 ;
  assign n48453 = n48443 & n48452 ;
  assign n48454 = ~n47997 & ~n48453 ;
  assign n48455 = \pi0223  & n24691 ;
  assign n48456 = n48145 & n48455 ;
  assign n48457 = ~n43784 & ~n48456 ;
  assign n48458 = n23880 & ~n48457 ;
  assign n48459 = ~n48437 & ~n48457 ;
  assign n48460 = n48436 & n48459 ;
  assign n48461 = ~n48458 & ~n48460 ;
  assign n48462 = \pi0778  & ~n48157 ;
  assign n48463 = n23885 & n48126 ;
  assign n48464 = ~n48462 & n48463 ;
  assign n48465 = ~n23885 & ~n48176 ;
  assign n48466 = ~\pi0628  & n20844 ;
  assign n48467 = \pi0223  & n20844 ;
  assign n48468 = n48145 & n48467 ;
  assign n48469 = ~n48466 & ~n48468 ;
  assign n48470 = ~n48465 & ~n48469 ;
  assign n48471 = ~n48464 & n48470 ;
  assign n48472 = \pi0628  & n20843 ;
  assign n48473 = \pi0223  & n20843 ;
  assign n48474 = n48145 & n48473 ;
  assign n48475 = ~n48472 & ~n48474 ;
  assign n48476 = ~n48465 & ~n48475 ;
  assign n48477 = ~n48464 & n48476 ;
  assign n48478 = \pi0223  & ~\pi0628  ;
  assign n48479 = n20843 & n48478 ;
  assign n48480 = n48145 & n48479 ;
  assign n48481 = \pi0223  & \pi0628  ;
  assign n48482 = n20844 & n48481 ;
  assign n48483 = n48145 & n48482 ;
  assign n48484 = ~n48480 & ~n48483 ;
  assign n48485 = ~n48477 & n48484 ;
  assign n48486 = ~n48471 & n48485 ;
  assign n48487 = n48461 & n48486 ;
  assign n48488 = \pi0792  & ~n48487 ;
  assign n48489 = n22155 & ~n48431 ;
  assign n48490 = ~n48432 & n48489 ;
  assign n48491 = n48429 & n48490 ;
  assign n48492 = ~n21034 & n48491 ;
  assign n48493 = ~n22147 & n48126 ;
  assign n48494 = ~n48462 & n48493 ;
  assign n48495 = ~n22147 & n23667 ;
  assign n48496 = \pi0223  & n23667 ;
  assign n48497 = n48145 & n48496 ;
  assign n48498 = ~n48495 & ~n48497 ;
  assign n48499 = \pi0781  & ~n48498 ;
  assign n48500 = ~n21034 & n48499 ;
  assign n48501 = ~n48494 & n48500 ;
  assign n48502 = ~n48492 & ~n48501 ;
  assign n48503 = n1689 & ~n22218 ;
  assign n48504 = n1259 & n48503 ;
  assign n48505 = n1249 & n48504 ;
  assign n48506 = \pi0642  & ~n22276 ;
  assign n48507 = n48000 & ~n48506 ;
  assign n48508 = n1281 & n48507 ;
  assign n48509 = n48505 & n48508 ;
  assign n48510 = ~n48000 & n48255 ;
  assign n48511 = n1281 & n48510 ;
  assign n48512 = n1260 & n48511 ;
  assign n48513 = \pi0223  & ~n48512 ;
  assign n48514 = ~n48509 & n48513 ;
  assign n48515 = n1281 & n47808 ;
  assign n48516 = n1260 & n48515 ;
  assign n48517 = ~\pi0642  & n20854 ;
  assign n48518 = ~n20783 & n21572 ;
  assign n48519 = ~n48517 & ~n48518 ;
  assign n48520 = n48000 & n48519 ;
  assign n48521 = ~n48516 & n48520 ;
  assign n48522 = n47585 & ~n48000 ;
  assign n48523 = n48411 & ~n48522 ;
  assign n48524 = ~n48521 & n48523 ;
  assign n48525 = ~n48514 & n48524 ;
  assign n48526 = ~\pi0223  & n48411 ;
  assign n48527 = ~n21289 & n48526 ;
  assign n48528 = \pi0039  & n48411 ;
  assign n48529 = ~n48527 & ~n48528 ;
  assign n48530 = n6861 & n48529 ;
  assign n48531 = ~n48525 & n48530 ;
  assign n48532 = ~n48418 & ~n48531 ;
  assign n48533 = \pi0223  & ~n48210 ;
  assign n48534 = ~n22330 & ~n48000 ;
  assign n48535 = ~n21243 & n48534 ;
  assign n48536 = ~n21249 & n48535 ;
  assign n48537 = n22661 & n48536 ;
  assign n48538 = ~n47776 & ~n48537 ;
  assign n48539 = n48533 & n48538 ;
  assign n48540 = ~n21472 & n48205 ;
  assign n48541 = \pi0299  & ~n48540 ;
  assign n48542 = ~n22657 & n48081 ;
  assign n48543 = ~n22660 & n48542 ;
  assign n48544 = n22664 & n48543 ;
  assign n48545 = n48541 & ~n48544 ;
  assign n48546 = ~n48539 & n48545 ;
  assign n48547 = ~\pi0039  & n48546 ;
  assign n48548 = \pi0223  & n48200 ;
  assign n48549 = ~n22673 & n48534 ;
  assign n48550 = ~n22671 & n48549 ;
  assign n48551 = n22669 & n48550 ;
  assign n48552 = n48548 & ~n48551 ;
  assign n48553 = ~n47751 & n48552 ;
  assign n48554 = n22676 & n48081 ;
  assign n48555 = n48192 & ~n48554 ;
  assign n48556 = ~\pi0039  & n48555 ;
  assign n48557 = ~n48553 & n48556 ;
  assign n48558 = ~n48547 & ~n48557 ;
  assign n48559 = ~\pi0038  & ~\pi0223  ;
  assign n48560 = ~n43150 & ~n48559 ;
  assign n48561 = ~n48558 & ~n48560 ;
  assign n48562 = ~n48521 & ~n48522 ;
  assign n48563 = ~\pi0223  & ~n21285 ;
  assign n48564 = ~n48562 & n48563 ;
  assign n48565 = ~n48514 & ~n48564 ;
  assign n48566 = n48070 & n48565 ;
  assign n48567 = ~\pi0215  & n48566 ;
  assign n48568 = ~n6732 & ~n48314 ;
  assign n48569 = ~n48000 & n48322 ;
  assign n48570 = n20854 & ~n47595 ;
  assign n48571 = n46321 & ~n48570 ;
  assign n48572 = ~n47605 & n48571 ;
  assign n48573 = ~n22242 & ~n47592 ;
  assign n48574 = n47589 & n48573 ;
  assign n48575 = n21370 & ~n48574 ;
  assign n48576 = \pi0680  & ~n48506 ;
  assign n48577 = \pi0642  & ~n21286 ;
  assign n48578 = ~n21327 & n48577 ;
  assign n48579 = n48576 & ~n48578 ;
  assign n48580 = ~n48575 & n48579 ;
  assign n48581 = ~n48572 & n48580 ;
  assign n48582 = ~n48569 & ~n48581 ;
  assign n48583 = n48568 & ~n48582 ;
  assign n48584 = ~\pi0680  & ~n48333 ;
  assign n48585 = ~n48329 & n48584 ;
  assign n48586 = \pi0681  & ~n48585 ;
  assign n48587 = n1281 & ~n48506 ;
  assign n48588 = n48505 & n48587 ;
  assign n48589 = ~n6711 & ~n48588 ;
  assign n48590 = ~\pi0120  & ~n6711 ;
  assign n48591 = ~n21301 & n48590 ;
  assign n48592 = ~n48589 & ~n48591 ;
  assign n48593 = \pi0680  & n48592 ;
  assign n48594 = ~\pi0642  & ~n22218 ;
  assign n48595 = ~n22218 & n22276 ;
  assign n48596 = ~n21285 & n48595 ;
  assign n48597 = ~n48594 & ~n48596 ;
  assign n48598 = ~n21371 & ~n48597 ;
  assign n48599 = ~n21359 & n48598 ;
  assign n48600 = n22256 & ~n48597 ;
  assign n48601 = ~n48599 & ~n48600 ;
  assign n48602 = \pi0642  & n22276 ;
  assign n48603 = ~n21285 & n48602 ;
  assign n48604 = n6711 & ~n48603 ;
  assign n48605 = n48601 & n48604 ;
  assign n48606 = n48593 & ~n48605 ;
  assign n48607 = n48586 & ~n48606 ;
  assign n48608 = ~n48346 & ~n48607 ;
  assign n48609 = \pi0223  & ~n48608 ;
  assign n48610 = ~n48583 & n48609 ;
  assign n48611 = ~n2352 & ~n48610 ;
  assign n48612 = n21370 & ~n22302 ;
  assign n48613 = n21328 & n48577 ;
  assign n48614 = \pi0642  & ~n20784 ;
  assign n48615 = ~n22023 & n48614 ;
  assign n48616 = ~n21306 & n48615 ;
  assign n48617 = ~n22022 & n48616 ;
  assign n48618 = \pi0680  & ~n48617 ;
  assign n48619 = ~n48613 & n48618 ;
  assign n48620 = ~n22496 & n48619 ;
  assign n48621 = ~n48612 & n48620 ;
  assign n48622 = ~n22311 & n46321 ;
  assign n48623 = ~n48225 & ~n48622 ;
  assign n48624 = n48621 & n48623 ;
  assign n48625 = ~n48000 & n48229 ;
  assign n48626 = ~n48225 & n48625 ;
  assign n48627 = ~n6732 & ~n48626 ;
  assign n48628 = ~n48624 & n48627 ;
  assign n48629 = n6711 & ~n22276 ;
  assign n48630 = ~n21285 & n48629 ;
  assign n48631 = ~n43050 & ~n48630 ;
  assign n48632 = ~n22333 & ~n48631 ;
  assign n48633 = ~n21362 & n48632 ;
  assign n48634 = ~n21364 & n48633 ;
  assign n48635 = \pi0642  & n6711 ;
  assign n48636 = ~n22276 & n48635 ;
  assign n48637 = ~n21285 & n48636 ;
  assign n48638 = ~n6711 & ~n21285 ;
  assign n48639 = \pi0680  & ~n48638 ;
  assign n48640 = \pi0681  & n48639 ;
  assign n48641 = n48000 & ~n48597 ;
  assign n48642 = ~n48640 & ~n48641 ;
  assign n48643 = ~n48637 & ~n48642 ;
  assign n48644 = ~n48634 & n48643 ;
  assign n48645 = ~\pi0680  & \pi0681  ;
  assign n48646 = ~n48354 & n48645 ;
  assign n48647 = ~n48242 & ~n48646 ;
  assign n48648 = ~n48644 & n48647 ;
  assign n48649 = n6732 & ~n48648 ;
  assign n48650 = ~\pi0223  & ~n48649 ;
  assign n48651 = ~n48628 & n48650 ;
  assign n48652 = ~\pi0215  & ~n48651 ;
  assign n48653 = n48611 & n48652 ;
  assign n48654 = ~n48567 & ~n48653 ;
  assign n48655 = n6732 & ~n48383 ;
  assign n48656 = n21392 & n48632 ;
  assign n48657 = n48643 & ~n48656 ;
  assign n48658 = ~\pi0223  & ~n48646 ;
  assign n48659 = ~n48657 & n48658 ;
  assign n48660 = n48655 & n48659 ;
  assign n48661 = ~\pi0223  & ~n6732 ;
  assign n48662 = n48385 & n48661 ;
  assign n48663 = \pi0215  & ~n48662 ;
  assign n48664 = \pi0680  & ~n46321 ;
  assign n48665 = \pi0680  & n21419 ;
  assign n48666 = ~n21425 & n21877 ;
  assign n48667 = ~n48665 & ~n48666 ;
  assign n48668 = ~n22333 & ~n48667 ;
  assign n48669 = ~n48664 & ~n48668 ;
  assign n48670 = n21370 & ~n22356 ;
  assign n48671 = n21370 & ~n22454 ;
  assign n48672 = ~n22455 & n48671 ;
  assign n48673 = ~n48670 & ~n48672 ;
  assign n48674 = ~n21516 & ~n22023 ;
  assign n48675 = ~n21615 & ~n48674 ;
  assign n48676 = \pi0642  & ~n48675 ;
  assign n48677 = n48673 & ~n48676 ;
  assign n48678 = ~n48669 & n48677 ;
  assign n48679 = \pi0642  & ~\pi0680  ;
  assign n48680 = n21515 & n48679 ;
  assign n48681 = n21516 & n48679 ;
  assign n48682 = ~n21520 & n48681 ;
  assign n48683 = ~n48680 & ~n48682 ;
  assign n48684 = \pi0681  & n48683 ;
  assign n48685 = \pi0215  & n48684 ;
  assign n48686 = ~n48678 & n48685 ;
  assign n48687 = ~n48663 & ~n48686 ;
  assign n48688 = ~n48660 & ~n48687 ;
  assign n48689 = \pi0299  & ~n48688 ;
  assign n48690 = ~n48000 & ~n48273 ;
  assign n48691 = \pi0616  & n48593 ;
  assign n48692 = n22214 & n22216 ;
  assign n48693 = ~n21285 & n22276 ;
  assign n48694 = \pi0642  & ~n48693 ;
  assign n48695 = n48593 & ~n48694 ;
  assign n48696 = ~n48692 & n48695 ;
  assign n48697 = ~n48691 & ~n48696 ;
  assign n48698 = ~n48690 & n48697 ;
  assign n48699 = n6732 & ~n48262 ;
  assign n48700 = ~n48270 & n48699 ;
  assign n48701 = ~n48698 & n48700 ;
  assign n48702 = \pi0680  & ~n22197 ;
  assign n48703 = \pi0680  & n21516 ;
  assign n48704 = ~n22183 & n48703 ;
  assign n48705 = ~n48702 & ~n48704 ;
  assign n48706 = ~n6711 & n22188 ;
  assign n48707 = ~n21515 & n48706 ;
  assign n48708 = ~n21521 & n48707 ;
  assign n48709 = ~n22188 & n22276 ;
  assign n48710 = \pi0642  & ~n48709 ;
  assign n48711 = ~n48708 & ~n48710 ;
  assign n48712 = ~n48705 & n48711 ;
  assign n48713 = ~\pi0680  & n48280 ;
  assign n48714 = ~\pi0680  & n48278 ;
  assign n48715 = ~n21520 & n48714 ;
  assign n48716 = ~n48713 & ~n48715 ;
  assign n48717 = ~n48276 & ~n48716 ;
  assign n48718 = \pi0681  & ~n48717 ;
  assign n48719 = ~n48712 & n48718 ;
  assign n48720 = ~n6732 & ~n48292 ;
  assign n48721 = ~n48719 & n48720 ;
  assign n48722 = \pi0223  & \pi0299  ;
  assign n48723 = ~n48721 & n48722 ;
  assign n48724 = ~n48701 & n48723 ;
  assign n48725 = ~n48689 & ~n48724 ;
  assign n48726 = n48654 & ~n48725 ;
  assign n48727 = n2165 & ~n48522 ;
  assign n48728 = ~n48521 & n48727 ;
  assign n48729 = ~n46507 & ~n48728 ;
  assign n48730 = n43384 & n48729 ;
  assign n48731 = n6761 & n48271 ;
  assign n48732 = ~n48698 & n48731 ;
  assign n48733 = ~n6761 & ~n48292 ;
  assign n48734 = ~n48719 & n48733 ;
  assign n48735 = n43374 & ~n48734 ;
  assign n48736 = ~n48732 & n48735 ;
  assign n48737 = \pi0039  & ~n48736 ;
  assign n48738 = ~n48730 & n48737 ;
  assign n48739 = ~n6761 & n48626 ;
  assign n48740 = ~n6761 & n48621 ;
  assign n48741 = n48623 & n48740 ;
  assign n48742 = ~n48739 & ~n48741 ;
  assign n48743 = n6761 & ~n48646 ;
  assign n48744 = ~n48242 & n48743 ;
  assign n48745 = ~n48644 & n48744 ;
  assign n48746 = ~n2165 & ~n48745 ;
  assign n48747 = n48737 & n48746 ;
  assign n48748 = n48742 & n48747 ;
  assign n48749 = ~n48738 & ~n48748 ;
  assign n48750 = ~n48560 & ~n48749 ;
  assign n48751 = ~n48726 & n48750 ;
  assign n48752 = ~n48561 & ~n48751 ;
  assign n48753 = ~n48532 & n48752 ;
  assign n48754 = \pi0625  & ~n48753 ;
  assign n48755 = \pi1153  & n48151 ;
  assign n48756 = \pi1153  & n48416 ;
  assign n48757 = ~n48410 & n48756 ;
  assign n48758 = ~n48755 & ~n48757 ;
  assign n48759 = ~n48754 & ~n48758 ;
  assign n48760 = ~n44177 & ~n48532 ;
  assign n48761 = n48752 & n48760 ;
  assign n48762 = \pi0608  & n48155 ;
  assign n48763 = \pi0608  & ~n48151 ;
  assign n48764 = ~n48130 & n48763 ;
  assign n48765 = ~n48762 & ~n48764 ;
  assign n48766 = ~n48761 & ~n48765 ;
  assign n48767 = ~n48759 & n48766 ;
  assign n48768 = \pi0778  & ~n48148 ;
  assign n48769 = ~n48133 & n48768 ;
  assign n48770 = n20858 & n48416 ;
  assign n48771 = ~n48410 & n48770 ;
  assign n48772 = \pi0223  & n20858 ;
  assign n48773 = ~n6861 & n48772 ;
  assign n48774 = ~\pi0608  & ~n48773 ;
  assign n48775 = ~n48771 & n48774 ;
  assign n48776 = \pi0778  & ~n48775 ;
  assign n48777 = ~n48769 & ~n48776 ;
  assign n48778 = ~n48761 & n48777 ;
  assign n48779 = ~n23808 & ~n48778 ;
  assign n48780 = ~n48767 & n48779 ;
  assign n48781 = n26700 & n48780 ;
  assign n48782 = ~\pi0609  & n48184 ;
  assign n48783 = ~\pi0609  & n48419 ;
  assign n48784 = ~n48417 & n48783 ;
  assign n48785 = ~n48782 & ~n48784 ;
  assign n48786 = ~\pi0609  & n20865 ;
  assign n48787 = \pi0223  & n20865 ;
  assign n48788 = n48145 & n48787 ;
  assign n48789 = ~n48786 & ~n48788 ;
  assign n48790 = n48785 & ~n48789 ;
  assign n48791 = ~n26119 & ~n48157 ;
  assign n48792 = ~n26124 & n47999 ;
  assign n48793 = ~n26124 & n48124 ;
  assign n48794 = ~n48115 & n48793 ;
  assign n48795 = ~n48792 & ~n48794 ;
  assign n48796 = \pi0609  & n48184 ;
  assign n48797 = \pi0609  & n48419 ;
  assign n48798 = ~n48417 & n48797 ;
  assign n48799 = ~n48796 & ~n48798 ;
  assign n48800 = \pi0609  & n20864 ;
  assign n48801 = \pi0223  & n20864 ;
  assign n48802 = n48145 & n48801 ;
  assign n48803 = ~n48800 & ~n48802 ;
  assign n48804 = n48799 & ~n48803 ;
  assign n48805 = n48795 & ~n48804 ;
  assign n48806 = ~n48791 & n48805 ;
  assign n48807 = ~n48790 & n48806 ;
  assign n48808 = n43534 & ~n48807 ;
  assign n48809 = ~n48781 & ~n48808 ;
  assign n48810 = n48502 & n48809 ;
  assign n48811 = n23683 & ~n48434 ;
  assign n48812 = \pi0223  & ~n20876 ;
  assign n48813 = n48145 & n48812 ;
  assign n48814 = ~n24969 & ~n48813 ;
  assign n48815 = ~n21032 & ~n48814 ;
  assign n48816 = ~n48183 & ~n48814 ;
  assign n48817 = n48422 & n48816 ;
  assign n48818 = ~n48815 & ~n48817 ;
  assign n48819 = ~n48811 & ~n48818 ;
  assign n48820 = \pi0789  & n48819 ;
  assign n48821 = n30780 & ~n48157 ;
  assign n48822 = \pi0223  & ~n23380 ;
  assign n48823 = n48145 & n48822 ;
  assign n48824 = n23380 & n47999 ;
  assign n48825 = n23380 & n48124 ;
  assign n48826 = ~n48115 & n48825 ;
  assign n48827 = ~n48824 & ~n48826 ;
  assign n48828 = ~n48823 & n48827 ;
  assign n48829 = ~n48821 & n48828 ;
  assign n48830 = n23701 & ~n48829 ;
  assign n48831 = ~n48820 & ~n48830 ;
  assign n48832 = ~n21038 & n48831 ;
  assign n48833 = n48810 & n48832 ;
  assign n48834 = \pi0223  & n22160 ;
  assign n48835 = n48145 & n48834 ;
  assign n48836 = n20951 & ~n48835 ;
  assign n48837 = ~n22160 & ~n48829 ;
  assign n48838 = n48836 & ~n48837 ;
  assign n48839 = \pi0223  & ~\pi0626  ;
  assign n48840 = n48145 & n48839 ;
  assign n48841 = ~n43582 & ~n48840 ;
  assign n48842 = n48436 & ~n48841 ;
  assign n48843 = \pi0223  & \pi0626  ;
  assign n48844 = n48145 & n48843 ;
  assign n48845 = n20882 & ~n48844 ;
  assign n48846 = ~n48842 & n48845 ;
  assign n48847 = ~n48838 & ~n48846 ;
  assign n48848 = ~n43594 & ~n48844 ;
  assign n48849 = n48436 & ~n48848 ;
  assign n48850 = n20881 & ~n48840 ;
  assign n48851 = ~n48849 & n48850 ;
  assign n48852 = ~n23856 & ~n48851 ;
  assign n48853 = n48847 & n48852 ;
  assign n48854 = ~n26803 & ~n48853 ;
  assign n48855 = ~n48833 & ~n48854 ;
  assign n48856 = ~n48488 & ~n48855 ;
  assign n48857 = ~n21067 & ~n48856 ;
  assign n48858 = ~\pi0630  & ~n48167 ;
  assign n48859 = ~n48164 & n48858 ;
  assign n48860 = \pi0630  & ~n48173 ;
  assign n48861 = ~n48170 & n48860 ;
  assign n48862 = ~n48859 & ~n48861 ;
  assign n48863 = ~n20846 & n23880 ;
  assign n48864 = ~n48176 & n48863 ;
  assign n48865 = \pi0223  & ~n20910 ;
  assign n48866 = n48145 & n48865 ;
  assign n48867 = ~n43615 & ~n48866 ;
  assign n48868 = ~n48864 & ~n48867 ;
  assign n48869 = ~n30376 & n48868 ;
  assign n48870 = ~n48437 & n48868 ;
  assign n48871 = n48436 & n48870 ;
  assign n48872 = ~n48869 & ~n48871 ;
  assign n48873 = ~n24761 & n48872 ;
  assign n48874 = n48862 & n48873 ;
  assign n48875 = ~n29722 & ~n48874 ;
  assign n48876 = ~n47996 & ~n48875 ;
  assign n48877 = ~n48857 & n48876 ;
  assign n48878 = n48454 & ~n48877 ;
  assign n48879 = \pi0224  & n21768 ;
  assign n48880 = \pi0626  & n48879 ;
  assign n48881 = ~\pi0038  & \pi0224  ;
  assign n48882 = n21743 & n48881 ;
  assign n48883 = \pi0626  & n48882 ;
  assign n48884 = ~n47007 & n48883 ;
  assign n48885 = ~n48880 & ~n48884 ;
  assign n48886 = n20882 & n48885 ;
  assign n48887 = \pi0626  & n48886 ;
  assign n48888 = ~n47007 & n48882 ;
  assign n48889 = ~n48879 & ~n48888 ;
  assign n48890 = n20828 & ~n48889 ;
  assign n48891 = n23830 & ~n48879 ;
  assign n48892 = ~n48888 & n48891 ;
  assign n48893 = \pi0781  & n20811 ;
  assign n48894 = ~n48892 & ~n48893 ;
  assign n48895 = \pi0603  & \pi0614  ;
  assign n48896 = ~n20783 & n48895 ;
  assign n48897 = ~n21285 & ~n48896 ;
  assign n48898 = ~n6712 & ~n48897 ;
  assign n48899 = ~\pi0680  & ~n48898 ;
  assign n48900 = n21355 & ~n48896 ;
  assign n48901 = ~n21290 & ~n48896 ;
  assign n48902 = ~n21325 & n48901 ;
  assign n48903 = ~n48900 & ~n48902 ;
  assign n48904 = ~n21352 & ~n48898 ;
  assign n48905 = ~n48903 & n48904 ;
  assign n48906 = ~n48899 & ~n48905 ;
  assign n48907 = \pi0680  & ~n21352 ;
  assign n48908 = ~n48903 & n48907 ;
  assign n48909 = n21586 & ~n48908 ;
  assign n48910 = n48906 & n48909 ;
  assign n48911 = ~n21576 & ~n21577 ;
  assign n48912 = ~\pi0616  & n48909 ;
  assign n48913 = ~n48911 & n48912 ;
  assign n48914 = ~n48910 & ~n48913 ;
  assign n48915 = \pi0616  & ~n48898 ;
  assign n48916 = ~n21577 & ~n48898 ;
  assign n48917 = ~n21576 & n48916 ;
  assign n48918 = ~n48915 & ~n48917 ;
  assign n48919 = ~n21586 & n48918 ;
  assign n48920 = n48914 & ~n48919 ;
  assign n48921 = n6761 & n48920 ;
  assign n48922 = \pi0224  & ~n48921 ;
  assign n48923 = ~n21352 & ~n48896 ;
  assign n48924 = ~n21405 & n48923 ;
  assign n48925 = \pi0680  & ~n48924 ;
  assign n48926 = n21586 & n48925 ;
  assign n48927 = ~n46289 & ~n48898 ;
  assign n48928 = ~\pi0680  & n21586 ;
  assign n48929 = ~n48927 & n48928 ;
  assign n48930 = ~n48926 & ~n48929 ;
  assign n48931 = n6761 & n21586 ;
  assign n48932 = n6761 & ~n48898 ;
  assign n48933 = ~n46289 & n48932 ;
  assign n48934 = ~n48931 & ~n48933 ;
  assign n48935 = n48930 & ~n48934 ;
  assign n48936 = \pi0680  & n21403 ;
  assign n48937 = ~n21399 & n48936 ;
  assign n48938 = \pi0614  & \pi0680  ;
  assign n48939 = ~n21417 & n48938 ;
  assign n48940 = ~n48937 & ~n48939 ;
  assign n48941 = n21586 & ~n48940 ;
  assign n48942 = n6706 & ~n21425 ;
  assign n48943 = \pi0614  & ~n21419 ;
  assign n48944 = ~n48942 & n48943 ;
  assign n48945 = n42695 & ~n47606 ;
  assign n48946 = n21908 & ~n47606 ;
  assign n48947 = n21520 & n48946 ;
  assign n48948 = ~n48945 & ~n48947 ;
  assign n48949 = ~n48944 & n48948 ;
  assign n48950 = n48928 & ~n48949 ;
  assign n48951 = ~n48941 & ~n48950 ;
  assign n48952 = ~n21586 & ~n48949 ;
  assign n48953 = ~n6761 & ~n48952 ;
  assign n48954 = n48951 & n48953 ;
  assign n48955 = ~n48935 & ~n48954 ;
  assign n48956 = \pi0224  & n48955 ;
  assign n48957 = ~\pi0224  & ~n20783 ;
  assign n48958 = n48895 & n48957 ;
  assign n48959 = ~n21285 & n48958 ;
  assign n48960 = ~n47088 & n48959 ;
  assign n48961 = ~n22079 & n48960 ;
  assign n48962 = \pi0223  & ~n48961 ;
  assign n48963 = ~n48956 & n48962 ;
  assign n48964 = ~n6706 & ~n21570 ;
  assign n48965 = ~\pi0614  & ~n48964 ;
  assign n48966 = n21328 & n48965 ;
  assign n48967 = n21328 & n46825 ;
  assign n48968 = ~n21573 & n48967 ;
  assign n48969 = ~\pi0616  & n48968 ;
  assign n48970 = ~n48966 & ~n48969 ;
  assign n48971 = \pi0680  & n48896 ;
  assign n48972 = ~n21306 & ~n21903 ;
  assign n48973 = \pi0680  & ~n48895 ;
  assign n48974 = \pi0680  & ~n21306 ;
  assign n48975 = ~n21345 & n48974 ;
  assign n48976 = ~n48973 & ~n48975 ;
  assign n48977 = n48972 & ~n48976 ;
  assign n48978 = ~n48971 & ~n48977 ;
  assign n48979 = \pi0614  & ~n21341 ;
  assign n48980 = n48978 & ~n48979 ;
  assign n48981 = n48970 & n48980 ;
  assign n48982 = \pi0680  & ~n48896 ;
  assign n48983 = ~n48977 & n48982 ;
  assign n48984 = n21586 & ~n48983 ;
  assign n48985 = ~n48981 & n48984 ;
  assign n48986 = ~n6761 & n21586 ;
  assign n48987 = ~n6761 & ~n48979 ;
  assign n48988 = n48970 & n48987 ;
  assign n48989 = ~n48986 & ~n48988 ;
  assign n48990 = ~n48985 & ~n48989 ;
  assign n48991 = ~n48963 & ~n48990 ;
  assign n48992 = n48922 & n48991 ;
  assign n48993 = ~\pi0299  & n48963 ;
  assign n48994 = ~n21586 & ~n48896 ;
  assign n48995 = ~n21286 & ~n21586 ;
  assign n48996 = n21328 & n48995 ;
  assign n48997 = ~n48994 & ~n48996 ;
  assign n48998 = ~n6761 & ~n48997 ;
  assign n48999 = ~\pi0680  & ~n48896 ;
  assign n49000 = ~\pi0680  & ~n21286 ;
  assign n49001 = n21328 & n49000 ;
  assign n49002 = ~n48999 & ~n49001 ;
  assign n49003 = n48976 & n49002 ;
  assign n49004 = n48986 & ~n49003 ;
  assign n49005 = ~n48998 & ~n49004 ;
  assign n49006 = \pi0614  & n6709 ;
  assign n49007 = \pi0614  & n20784 ;
  assign n49008 = ~n21285 & n49007 ;
  assign n49009 = ~n49006 & ~n49008 ;
  assign n49010 = ~n6709 & ~n49009 ;
  assign n49011 = n20784 & ~n49009 ;
  assign n49012 = ~n21359 & n49011 ;
  assign n49013 = ~n49010 & ~n49012 ;
  assign n49014 = n6761 & n49013 ;
  assign n49015 = n6148 & ~n49014 ;
  assign n49016 = n49005 & n49015 ;
  assign n49017 = ~\pi0224  & \pi0614  ;
  assign n49018 = ~\pi0222  & \pi0603  ;
  assign n49019 = ~n20783 & n49018 ;
  assign n49020 = n49017 & n49019 ;
  assign n49021 = ~n21285 & n49020 ;
  assign n49022 = ~\pi0223  & ~n49021 ;
  assign n49023 = ~\pi0299  & n49022 ;
  assign n49024 = ~n49016 & n49023 ;
  assign n49025 = ~n48993 & ~n49024 ;
  assign n49026 = ~n48992 & ~n49025 ;
  assign n49027 = n9627 & n49026 ;
  assign n49028 = ~n21285 & n48896 ;
  assign n49029 = \pi0224  & n21285 ;
  assign n49030 = n2352 & ~n49029 ;
  assign n49031 = ~n49028 & n49030 ;
  assign n49032 = ~\pi0215  & ~n49031 ;
  assign n49033 = ~n6732 & ~n48997 ;
  assign n49034 = ~n6732 & n21586 ;
  assign n49035 = ~n49003 & n49034 ;
  assign n49036 = ~n49033 & ~n49035 ;
  assign n49037 = n6732 & n49013 ;
  assign n49038 = ~\pi0224  & ~n49037 ;
  assign n49039 = n49036 & n49038 ;
  assign n49040 = ~n2352 & ~n49039 ;
  assign n49041 = n49032 & ~n49040 ;
  assign n49042 = n6732 & n48920 ;
  assign n49043 = \pi0224  & ~n49042 ;
  assign n49044 = ~n6732 & ~n48979 ;
  assign n49045 = n48970 & n49044 ;
  assign n49046 = ~n49034 & ~n49045 ;
  assign n49047 = ~n48985 & ~n49046 ;
  assign n49048 = n49032 & ~n49047 ;
  assign n49049 = n49043 & n49048 ;
  assign n49050 = ~n49041 & ~n49049 ;
  assign n49051 = ~n22055 & n48960 ;
  assign n49052 = \pi0299  & ~n49051 ;
  assign n49053 = ~n21948 & ~n49052 ;
  assign n49054 = ~n6732 & ~n48952 ;
  assign n49055 = n48951 & n49054 ;
  assign n49056 = \pi0224  & ~n49055 ;
  assign n49057 = n6732 & n21586 ;
  assign n49058 = n6732 & ~n48898 ;
  assign n49059 = ~n46289 & n49058 ;
  assign n49060 = ~n49057 & ~n49059 ;
  assign n49061 = n48930 & ~n49060 ;
  assign n49062 = ~n21948 & ~n49061 ;
  assign n49063 = n49056 & n49062 ;
  assign n49064 = ~n49053 & ~n49063 ;
  assign n49065 = n9627 & n49064 ;
  assign n49066 = n49050 & n49065 ;
  assign n49067 = ~n49027 & ~n49066 ;
  assign n49068 = n21481 & n49017 ;
  assign n49069 = n21477 & n49017 ;
  assign n49070 = ~n21263 & n49069 ;
  assign n49071 = ~n49068 & ~n49070 ;
  assign n49072 = ~\pi0299  & ~n49071 ;
  assign n49073 = ~\pi0614  & n21481 ;
  assign n49074 = ~\pi0614  & n21477 ;
  assign n49075 = ~n21263 & n49074 ;
  assign n49076 = ~n49073 & ~n49075 ;
  assign n49077 = n21265 & n49076 ;
  assign n49078 = \pi0224  & n21266 ;
  assign n49079 = \pi0198  & \pi0224  ;
  assign n49080 = n21247 & n49079 ;
  assign n49081 = ~n49078 & ~n49080 ;
  assign n49082 = ~\pi0299  & ~n49081 ;
  assign n49083 = n49077 & n49082 ;
  assign n49084 = ~n49072 & ~n49083 ;
  assign n49085 = ~n21473 & n48895 ;
  assign n49086 = ~n21472 & n49085 ;
  assign n49087 = \pi0224  & ~n43275 ;
  assign n49088 = \pi0299  & ~n49087 ;
  assign n49089 = n21247 & n48107 ;
  assign n49090 = ~n49088 & ~n49089 ;
  assign n49091 = n49086 & ~n49090 ;
  assign n49092 = \pi0224  & n21205 ;
  assign n49093 = \pi0224  & n21237 ;
  assign n49094 = n21232 & n49093 ;
  assign n49095 = ~n49092 & ~n49094 ;
  assign n49096 = \pi0299  & ~n49095 ;
  assign n49097 = ~\pi0039  & ~n49096 ;
  assign n49098 = ~n49091 & n49097 ;
  assign n49099 = ~\pi0038  & n49098 ;
  assign n49100 = n49084 & n49099 ;
  assign n49101 = \pi0224  & ~n21757 ;
  assign n49102 = n1689 & n48896 ;
  assign n49103 = n8413 & n49102 ;
  assign n49104 = n1354 & n49103 ;
  assign n49105 = n1358 & n49104 ;
  assign n49106 = \pi0038  & ~n49105 ;
  assign n49107 = ~n49101 & n49106 ;
  assign n49108 = n26645 & ~n49107 ;
  assign n49109 = ~n49100 & n49108 ;
  assign n49110 = n49067 & n49109 ;
  assign n49111 = n20985 & n48879 ;
  assign n49112 = n20985 & n48882 ;
  assign n49113 = ~n47007 & n49112 ;
  assign n49114 = ~n49111 & ~n49113 ;
  assign n49115 = \pi0224  & ~n6861 ;
  assign n49116 = ~n20985 & n49115 ;
  assign n49117 = ~n25588 & ~n49116 ;
  assign n49118 = n49114 & n49117 ;
  assign n49119 = ~n49110 & n49118 ;
  assign n49120 = n21776 & ~n48879 ;
  assign n49121 = ~n48888 & n49120 ;
  assign n49122 = ~n48892 & ~n49121 ;
  assign n49123 = ~n49119 & n49122 ;
  assign n49124 = ~n48894 & ~n49123 ;
  assign n49125 = ~\pi0619  & ~n48879 ;
  assign n49126 = ~n48888 & n49125 ;
  assign n49127 = \pi1159  & ~n49126 ;
  assign n49128 = \pi0781  & n49127 ;
  assign n49129 = ~n49121 & n49127 ;
  assign n49130 = ~n49119 & n49129 ;
  assign n49131 = ~n49128 & ~n49130 ;
  assign n49132 = ~n49124 & ~n49131 ;
  assign n49133 = ~n48890 & ~n49132 ;
  assign n49134 = \pi0789  & ~n49133 ;
  assign n49135 = \pi0619  & n48879 ;
  assign n49136 = \pi0619  & n48882 ;
  assign n49137 = ~n47007 & n49136 ;
  assign n49138 = ~n49135 & ~n49137 ;
  assign n49139 = \pi0619  & ~n48879 ;
  assign n49140 = ~n48888 & n49139 ;
  assign n49141 = \pi0781  & ~n49140 ;
  assign n49142 = ~n49121 & ~n49140 ;
  assign n49143 = ~n49119 & n49142 ;
  assign n49144 = ~n49141 & ~n49143 ;
  assign n49145 = ~n49124 & ~n49144 ;
  assign n49146 = n49138 & ~n49145 ;
  assign n49147 = n31279 & ~n49146 ;
  assign n49148 = ~n49134 & ~n49147 ;
  assign n49149 = ~\pi0789  & ~n49121 ;
  assign n49150 = ~n49119 & n49149 ;
  assign n49151 = ~n21806 & ~n49150 ;
  assign n49152 = ~n49124 & ~n49151 ;
  assign n49153 = n48886 & ~n49152 ;
  assign n49154 = n49148 & n49153 ;
  assign n49155 = ~n48887 & ~n49154 ;
  assign n49156 = ~\pi0626  & n48879 ;
  assign n49157 = ~\pi0626  & n48882 ;
  assign n49158 = ~n47007 & n49157 ;
  assign n49159 = ~n49156 & ~n49158 ;
  assign n49160 = n20881 & n49159 ;
  assign n49161 = ~\pi0626  & n49160 ;
  assign n49162 = ~n49152 & n49160 ;
  assign n49163 = n49148 & n49162 ;
  assign n49164 = ~n49161 & ~n49163 ;
  assign n49165 = n31306 & ~n48879 ;
  assign n49166 = ~n48888 & n49165 ;
  assign n49167 = \pi0662  & n1689 ;
  assign n49168 = n20855 & n49167 ;
  assign n49169 = n8413 & n49168 ;
  assign n49170 = n1354 & n49169 ;
  assign n49171 = n1358 & n49170 ;
  assign n49172 = \pi0038  & ~n49171 ;
  assign n49173 = ~n49101 & n49172 ;
  assign n49174 = n6861 & ~n49173 ;
  assign n49175 = \pi0038  & n49174 ;
  assign n49176 = ~\pi0662  & ~n26996 ;
  assign n49177 = ~\pi0662  & ~n6732 ;
  assign n49178 = ~n6732 & ~n21961 ;
  assign n49179 = n21954 & n49178 ;
  assign n49180 = ~n49177 & ~n49179 ;
  assign n49181 = ~n49176 & ~n49180 ;
  assign n49182 = \pi0662  & ~n21972 ;
  assign n49183 = ~n21970 & n49182 ;
  assign n49184 = ~n21672 & n49183 ;
  assign n49185 = n6732 & n49184 ;
  assign n49186 = ~\pi0662  & ~n21654 ;
  assign n49187 = ~n21657 & n49186 ;
  assign n49188 = n6732 & n49187 ;
  assign n49189 = ~n21684 & n49188 ;
  assign n49190 = ~n49185 & ~n49189 ;
  assign n49191 = \pi0224  & n49190 ;
  assign n49192 = ~n49181 & n49191 ;
  assign n49193 = ~\pi0224  & \pi0662  ;
  assign n49194 = ~n22055 & n49193 ;
  assign n49195 = n22054 & n49194 ;
  assign n49196 = \pi0215  & ~n49195 ;
  assign n49197 = ~n49192 & n49196 ;
  assign n49198 = \pi0299  & ~n49197 ;
  assign n49199 = \pi0662  & n47278 ;
  assign n49200 = \pi0662  & ~\pi0680  ;
  assign n49201 = n47283 & n49200 ;
  assign n49202 = ~n49199 & ~n49201 ;
  assign n49203 = ~\pi0662  & ~n21593 ;
  assign n49204 = ~n21709 & n49203 ;
  assign n49205 = ~\pi0662  & \pi0681  ;
  assign n49206 = n47283 & n49205 ;
  assign n49207 = ~n49204 & ~n49206 ;
  assign n49208 = n49202 & n49207 ;
  assign n49209 = \pi0662  & \pi0680  ;
  assign n49210 = n22030 & n49209 ;
  assign n49211 = ~n22025 & n49209 ;
  assign n49212 = n22033 & n49211 ;
  assign n49213 = ~n49210 & ~n49212 ;
  assign n49214 = n6732 & n49213 ;
  assign n49215 = \pi0662  & n20855 ;
  assign n49216 = ~n21905 & n49215 ;
  assign n49217 = ~n22039 & n49216 ;
  assign n49218 = ~n6732 & ~n49217 ;
  assign n49219 = ~\pi0224  & ~n49218 ;
  assign n49220 = ~n49214 & n49219 ;
  assign n49221 = n21446 & ~n49220 ;
  assign n49222 = n49208 & n49221 ;
  assign n49223 = ~n6732 & ~n21334 ;
  assign n49224 = n6713 & ~n6732 ;
  assign n49225 = ~n21329 & n49224 ;
  assign n49226 = ~n49223 & ~n49225 ;
  assign n49227 = \pi0224  & n49226 ;
  assign n49228 = \pi0224  & ~n6707 ;
  assign n49229 = ~n48037 & n49228 ;
  assign n49230 = ~n49227 & ~n49229 ;
  assign n49231 = ~n47184 & ~n49220 ;
  assign n49232 = n49230 & n49231 ;
  assign n49233 = ~n20854 & n49209 ;
  assign n49234 = ~n21285 & n49233 ;
  assign n49235 = n49030 & ~n49234 ;
  assign n49236 = ~n49232 & ~n49235 ;
  assign n49237 = ~n49222 & n49236 ;
  assign n49238 = ~\pi0215  & ~n49237 ;
  assign n49239 = n49198 & ~n49238 ;
  assign n49240 = n6761 & n49213 ;
  assign n49241 = ~n6761 & ~n49217 ;
  assign n49242 = n6148 & ~n49241 ;
  assign n49243 = ~n49240 & n49242 ;
  assign n49244 = n48001 & n49209 ;
  assign n49245 = ~n21285 & n49244 ;
  assign n49246 = ~\pi0223  & ~n49245 ;
  assign n49247 = n6761 & n49246 ;
  assign n49248 = ~n49243 & n49247 ;
  assign n49249 = n49208 & n49248 ;
  assign n49250 = ~n49243 & n49246 ;
  assign n49251 = ~n6707 & ~n48037 ;
  assign n49252 = ~n6761 & ~n21335 ;
  assign n49253 = ~n49251 & n49252 ;
  assign n49254 = \pi0224  & ~n49253 ;
  assign n49255 = n49250 & ~n49254 ;
  assign n49256 = ~n49249 & ~n49255 ;
  assign n49257 = ~\pi0662  & ~n6761 ;
  assign n49258 = ~n6761 & ~n21961 ;
  assign n49259 = n21954 & n49258 ;
  assign n49260 = ~n49257 & ~n49259 ;
  assign n49261 = ~n49176 & ~n49260 ;
  assign n49262 = n6761 & n49184 ;
  assign n49263 = n6761 & n49187 ;
  assign n49264 = ~n21684 & n49263 ;
  assign n49265 = ~n49262 & ~n49264 ;
  assign n49266 = \pi0224  & n49265 ;
  assign n49267 = ~n49261 & n49266 ;
  assign n49268 = ~n22079 & n49193 ;
  assign n49269 = n22054 & n49268 ;
  assign n49270 = \pi0223  & ~n49269 ;
  assign n49271 = ~n49267 & n49270 ;
  assign n49272 = ~\pi0299  & ~n49271 ;
  assign n49273 = n49256 & n49272 ;
  assign n49274 = \pi0039  & ~n49273 ;
  assign n49275 = ~n49239 & n49274 ;
  assign n49276 = ~\pi0224  & ~n47424 ;
  assign n49277 = ~n22097 & ~n49209 ;
  assign n49278 = ~n22095 & n49277 ;
  assign n49279 = \pi0224  & ~n47419 ;
  assign n49280 = \pi0299  & ~n49279 ;
  assign n49281 = ~n48108 & ~n49280 ;
  assign n49282 = ~n49278 & ~n49281 ;
  assign n49283 = ~n49276 & n49282 ;
  assign n49284 = ~\pi0224  & ~n48092 ;
  assign n49285 = ~n22102 & ~n49209 ;
  assign n49286 = ~n48091 & n49285 ;
  assign n49287 = \pi0224  & ~n47402 ;
  assign n49288 = ~\pi0299  & ~n49287 ;
  assign n49289 = ~n48096 & ~n49288 ;
  assign n49290 = ~n49286 & ~n49289 ;
  assign n49291 = ~n49284 & n49290 ;
  assign n49292 = ~n49283 & ~n49291 ;
  assign n49293 = ~\pi0039  & n49292 ;
  assign n49294 = n49174 & ~n49293 ;
  assign n49295 = ~n49275 & n49294 ;
  assign n49296 = ~n49175 & ~n49295 ;
  assign n49297 = ~\pi0224  & \pi0625  ;
  assign n49298 = ~n22727 & ~n49297 ;
  assign n49299 = n49296 & ~n49298 ;
  assign n49300 = ~\pi0625  & ~n48879 ;
  assign n49301 = ~n48888 & n49300 ;
  assign n49302 = \pi1153  & ~n49301 ;
  assign n49303 = ~n49299 & n49302 ;
  assign n49304 = ~\pi0224  & ~\pi0625  ;
  assign n49305 = ~n22734 & ~n49304 ;
  assign n49306 = n49296 & ~n49305 ;
  assign n49307 = \pi0625  & ~n48879 ;
  assign n49308 = ~n48888 & n49307 ;
  assign n49309 = ~\pi1153  & ~n49308 ;
  assign n49310 = ~n49306 & n49309 ;
  assign n49311 = ~n49303 & ~n49310 ;
  assign n49312 = n30780 & ~n49311 ;
  assign n49313 = ~n49115 & n49296 ;
  assign n49314 = n31274 & ~n49313 ;
  assign n49315 = n22160 & n48879 ;
  assign n49316 = n22160 & n48882 ;
  assign n49317 = ~n47007 & n49316 ;
  assign n49318 = ~n49315 & ~n49317 ;
  assign n49319 = n20951 & n49318 ;
  assign n49320 = ~n23380 & n48879 ;
  assign n49321 = ~n23380 & n48882 ;
  assign n49322 = ~n47007 & n49321 ;
  assign n49323 = ~n49320 & ~n49322 ;
  assign n49324 = n49319 & n49323 ;
  assign n49325 = ~n49314 & n49324 ;
  assign n49326 = ~n49312 & n49325 ;
  assign n49327 = ~n49166 & ~n49326 ;
  assign n49328 = n49164 & n49327 ;
  assign n49329 = n49155 & n49328 ;
  assign n49330 = \pi0788  & ~n49329 ;
  assign n49331 = ~\pi0680  & n48949 ;
  assign n49332 = ~n22191 & ~n47656 ;
  assign n49333 = \pi0614  & ~n48709 ;
  assign n49334 = \pi0680  & ~n49333 ;
  assign n49335 = n49332 & n49334 ;
  assign n49336 = ~n49331 & ~n49335 ;
  assign n49337 = \pi0662  & n49336 ;
  assign n49338 = ~\pi0662  & ~n6708 ;
  assign n49339 = ~n48948 & n49338 ;
  assign n49340 = \pi0614  & n49338 ;
  assign n49341 = ~n21419 & n49340 ;
  assign n49342 = ~n48942 & n49341 ;
  assign n49343 = \pi0224  & ~n49342 ;
  assign n49344 = ~n49339 & n49343 ;
  assign n49345 = n48951 & n49344 ;
  assign n49346 = ~n49337 & n49345 ;
  assign n49347 = \pi0614  & n21515 ;
  assign n49348 = \pi0614  & n21516 ;
  assign n49349 = ~n21520 & n49348 ;
  assign n49350 = ~n49347 & ~n49349 ;
  assign n49351 = n22454 & n48938 ;
  assign n49352 = n22023 & n48938 ;
  assign n49353 = ~n21520 & n49352 ;
  assign n49354 = ~n49351 & ~n49353 ;
  assign n49355 = n49350 & n49354 ;
  assign n49356 = \pi0662  & ~n49355 ;
  assign n49357 = ~\pi0614  & ~n22333 ;
  assign n49358 = ~n48667 & n49357 ;
  assign n49359 = ~\pi0616  & ~\pi0642  ;
  assign n49360 = ~n22356 & n49359 ;
  assign n49361 = \pi0662  & ~n49360 ;
  assign n49362 = n49358 & n49361 ;
  assign n49363 = ~n49356 & ~n49362 ;
  assign n49364 = ~\pi0662  & ~n20783 ;
  assign n49365 = n48895 & n49364 ;
  assign n49366 = ~n21285 & n49365 ;
  assign n49367 = ~n47088 & n49366 ;
  assign n49368 = ~n21615 & n49367 ;
  assign n49369 = ~\pi0224  & ~n49368 ;
  assign n49370 = n49363 & n49369 ;
  assign n49371 = ~n6761 & ~n49370 ;
  assign n49372 = ~n49346 & n49371 ;
  assign n49373 = \pi0223  & ~n49372 ;
  assign n49374 = ~n48927 & n49200 ;
  assign n49375 = \pi0614  & ~n48516 ;
  assign n49376 = n1281 & n48505 ;
  assign n49377 = ~\pi0614  & ~n49376 ;
  assign n49378 = ~n22532 & ~n49377 ;
  assign n49379 = ~n49375 & n49378 ;
  assign n49380 = \pi0616  & ~n49379 ;
  assign n49381 = \pi0614  & ~n48693 ;
  assign n49382 = ~n22221 & ~n49381 ;
  assign n49383 = ~n49380 & n49382 ;
  assign n49384 = ~n22217 & n49383 ;
  assign n49385 = \pi0616  & ~n49375 ;
  assign n49386 = n49378 & n49385 ;
  assign n49387 = n49209 & ~n49386 ;
  assign n49388 = ~n49384 & n49387 ;
  assign n49389 = ~n49374 & ~n49388 ;
  assign n49390 = ~\pi0662  & n47074 ;
  assign n49391 = ~n21632 & n49390 ;
  assign n49392 = ~n21631 & n49391 ;
  assign n49393 = ~n6712 & n49338 ;
  assign n49394 = ~n48897 & n49393 ;
  assign n49395 = \pi0224  & ~n49394 ;
  assign n49396 = ~n49392 & n49395 ;
  assign n49397 = n48930 & n49396 ;
  assign n49398 = n49389 & n49397 ;
  assign n49399 = ~\pi0614  & \pi0616  ;
  assign n49400 = ~n47541 & n49399 ;
  assign n49401 = ~n47568 & ~n49400 ;
  assign n49402 = \pi0680  & ~n49401 ;
  assign n49403 = \pi0662  & ~n49402 ;
  assign n49404 = ~\pi0224  & ~n49367 ;
  assign n49405 = ~n49403 & n49404 ;
  assign n49406 = \pi0680  & ~n22354 ;
  assign n49407 = ~n49028 & n49404 ;
  assign n49408 = ~n49406 & n49407 ;
  assign n49409 = ~n49405 & ~n49408 ;
  assign n49410 = n6761 & n49409 ;
  assign n49411 = ~n49398 & n49410 ;
  assign n49412 = ~\pi0299  & ~n49411 ;
  assign n49413 = n49373 & n49412 ;
  assign n49414 = n21586 & ~n49003 ;
  assign n49415 = ~n48896 & n49338 ;
  assign n49416 = ~n21286 & n49338 ;
  assign n49417 = n21328 & n49416 ;
  assign n49418 = ~n49415 & ~n49417 ;
  assign n49419 = ~n49414 & n49418 ;
  assign n49420 = ~\pi0224  & ~n49419 ;
  assign n49421 = ~n20784 & n22025 ;
  assign n49422 = ~n21329 & ~n49421 ;
  assign n49423 = \pi0614  & n49422 ;
  assign n49424 = \pi0680  & ~n49423 ;
  assign n49425 = n49002 & ~n49424 ;
  assign n49426 = ~\pi0614  & ~n22025 ;
  assign n49427 = n21341 & n49426 ;
  assign n49428 = ~n6711 & ~n49427 ;
  assign n49429 = n49002 & ~n49428 ;
  assign n49430 = ~n22308 & n49429 ;
  assign n49431 = ~n49425 & ~n49430 ;
  assign n49432 = n49193 & n49431 ;
  assign n49433 = ~n49420 & ~n49432 ;
  assign n49434 = \pi0224  & ~n49338 ;
  assign n49435 = \pi0224  & ~n48979 ;
  assign n49436 = n48970 & n49435 ;
  assign n49437 = ~n49434 & ~n49436 ;
  assign n49438 = ~n48985 & ~n49437 ;
  assign n49439 = ~\pi0680  & ~n48979 ;
  assign n49440 = n48970 & n49439 ;
  assign n49441 = ~n48570 & n49399 ;
  assign n49442 = ~n47605 & n49441 ;
  assign n49443 = \pi0614  & ~n22276 ;
  assign n49444 = \pi0614  & ~n21286 ;
  assign n49445 = ~n21327 & n49444 ;
  assign n49446 = ~n49443 & ~n49445 ;
  assign n49447 = \pi0680  & n49446 ;
  assign n49448 = ~n49442 & n49447 ;
  assign n49449 = ~n47600 & n49448 ;
  assign n49450 = \pi0662  & ~n49449 ;
  assign n49451 = ~n49440 & n49450 ;
  assign n49452 = n49438 & ~n49451 ;
  assign n49453 = n21275 & ~n49452 ;
  assign n49454 = n49433 & n49453 ;
  assign n49455 = ~\pi0680  & ~n48918 ;
  assign n49456 = n47606 & ~n48693 ;
  assign n49457 = \pi0680  & ~n49375 ;
  assign n49458 = n49378 & n49457 ;
  assign n49459 = ~n47511 & ~n49458 ;
  assign n49460 = ~n49456 & ~n49459 ;
  assign n49461 = ~n22262 & n49460 ;
  assign n49462 = \pi0662  & ~n49461 ;
  assign n49463 = ~n49455 & n49462 ;
  assign n49464 = n48918 & n49338 ;
  assign n49465 = \pi0224  & ~n49464 ;
  assign n49466 = n48914 & n49465 ;
  assign n49467 = ~n49463 & n49466 ;
  assign n49468 = n22340 & ~n49028 ;
  assign n49469 = ~n22336 & n49468 ;
  assign n49470 = ~\pi0680  & ~n49028 ;
  assign n49471 = n49403 & ~n49470 ;
  assign n49472 = ~n49469 & n49471 ;
  assign n49473 = n6709 & n21583 ;
  assign n49474 = n20784 & n21583 ;
  assign n49475 = ~n21285 & n49474 ;
  assign n49476 = ~n49473 & ~n49475 ;
  assign n49477 = ~n6709 & ~n49476 ;
  assign n49478 = n20784 & ~n49476 ;
  assign n49479 = ~n21359 & n49478 ;
  assign n49480 = ~n49477 & ~n49479 ;
  assign n49481 = ~\pi0224  & n49480 ;
  assign n49482 = ~n49472 & n49481 ;
  assign n49483 = n21368 & ~n49482 ;
  assign n49484 = ~n49467 & n49483 ;
  assign n49485 = ~n20784 & n49233 ;
  assign n49486 = ~n21285 & n49485 ;
  assign n49487 = ~n49028 & ~n49486 ;
  assign n49488 = n46435 & ~n49487 ;
  assign n49489 = n43384 & ~n49488 ;
  assign n49490 = ~n49484 & n49489 ;
  assign n49491 = ~n49454 & n49490 ;
  assign n49492 = ~n49413 & ~n49491 ;
  assign n49493 = ~n49398 & n49409 ;
  assign n49494 = \pi0299  & n6732 ;
  assign n49495 = ~n49493 & n49494 ;
  assign n49496 = ~n6732 & n49344 ;
  assign n49497 = n48951 & n49496 ;
  assign n49498 = ~n49337 & n49497 ;
  assign n49499 = ~n6732 & n49369 ;
  assign n49500 = n49363 & n49499 ;
  assign n49501 = \pi0215  & ~n49500 ;
  assign n49502 = ~n49498 & n49501 ;
  assign n49503 = \pi0299  & ~n49502 ;
  assign n49504 = \pi0039  & ~n49503 ;
  assign n49505 = ~n49495 & n49504 ;
  assign n49506 = ~n6732 & ~n49452 ;
  assign n49507 = n49433 & n49506 ;
  assign n49508 = n6732 & ~n49482 ;
  assign n49509 = ~n47184 & ~n49508 ;
  assign n49510 = ~n47184 & ~n49463 ;
  assign n49511 = n49466 & n49510 ;
  assign n49512 = ~n49509 & ~n49511 ;
  assign n49513 = ~n49507 & ~n49512 ;
  assign n49514 = ~\pi0224  & ~n49487 ;
  assign n49515 = ~\pi0614  & n49209 ;
  assign n49516 = n49376 & n49515 ;
  assign n49517 = \pi0614  & n49209 ;
  assign n49518 = n48516 & n49517 ;
  assign n49519 = ~n49516 & ~n49518 ;
  assign n49520 = n1689 & ~n48896 ;
  assign n49521 = ~n49209 & n49520 ;
  assign n49522 = n1281 & n49521 ;
  assign n49523 = n1260 & n49522 ;
  assign n49524 = \pi0224  & ~n49523 ;
  assign n49525 = n49519 & n49524 ;
  assign n49526 = n49030 & ~n49525 ;
  assign n49527 = ~n49514 & n49526 ;
  assign n49528 = n43041 & ~n49527 ;
  assign n49529 = ~n49513 & n49528 ;
  assign n49530 = ~n49505 & ~n49529 ;
  assign n49531 = n49492 & ~n49530 ;
  assign n49532 = \pi0614  & n21481 ;
  assign n49533 = \pi0614  & n21477 ;
  assign n49534 = ~n21263 & n49533 ;
  assign n49535 = ~n49532 & ~n49534 ;
  assign n49536 = ~\pi0224  & ~n49535 ;
  assign n49537 = ~n22330 & n49209 ;
  assign n49538 = n22669 & n49537 ;
  assign n49539 = ~n22671 & ~n22673 ;
  assign n49540 = ~\pi0224  & n49539 ;
  assign n49541 = n49538 & n49540 ;
  assign n49542 = ~n49536 & ~n49541 ;
  assign n49543 = ~\pi0299  & ~n49542 ;
  assign n49544 = ~n22330 & ~n49209 ;
  assign n49545 = n22669 & n49544 ;
  assign n49546 = n49539 & n49545 ;
  assign n49547 = ~n47751 & ~n49546 ;
  assign n49548 = \pi0224  & n49076 ;
  assign n49549 = ~\pi0299  & n49548 ;
  assign n49550 = n49547 & n49549 ;
  assign n49551 = ~n49543 & ~n49550 ;
  assign n49552 = ~\pi0039  & ~n49551 ;
  assign n49553 = \pi0210  & n21247 ;
  assign n49554 = n49087 & ~n49553 ;
  assign n49555 = n49086 & ~n49554 ;
  assign n49556 = n49095 & ~n49209 ;
  assign n49557 = ~n49555 & n49556 ;
  assign n49558 = ~n49209 & ~n49557 ;
  assign n49559 = \pi0603  & ~\pi0614  ;
  assign n49560 = \pi0224  & n49559 ;
  assign n49561 = ~n21473 & n49560 ;
  assign n49562 = ~n21472 & n49561 ;
  assign n49563 = \pi0224  & n47773 ;
  assign n49564 = n47775 & n49563 ;
  assign n49565 = ~n49562 & ~n49564 ;
  assign n49566 = ~n21243 & ~n22330 ;
  assign n49567 = ~n21249 & n49566 ;
  assign n49568 = n22661 & n49567 ;
  assign n49569 = ~\pi0224  & ~n49086 ;
  assign n49570 = ~n49568 & n49569 ;
  assign n49571 = ~n49557 & ~n49570 ;
  assign n49572 = n49565 & n49571 ;
  assign n49573 = ~n49558 & ~n49572 ;
  assign n49574 = ~\pi0039  & \pi0299  ;
  assign n49575 = ~n49573 & n49574 ;
  assign n49576 = ~n49552 & ~n49575 ;
  assign n49577 = ~\pi0038  & n49576 ;
  assign n49578 = ~n49531 & n49577 ;
  assign n49579 = n21754 & n49485 ;
  assign n49580 = n1266 & n49579 ;
  assign n49581 = n1354 & n49580 ;
  assign n49582 = n1358 & n49581 ;
  assign n49583 = n49107 & ~n49582 ;
  assign n49584 = n6861 & ~n49583 ;
  assign n49585 = ~n49578 & n49584 ;
  assign n49586 = ~n49305 & ~n49585 ;
  assign n49587 = n6861 & ~n49107 ;
  assign n49588 = ~n49100 & n49587 ;
  assign n49589 = n49067 & n49588 ;
  assign n49590 = ~n49298 & ~n49589 ;
  assign n49591 = ~\pi1153  & ~n49590 ;
  assign n49592 = ~n49586 & n49591 ;
  assign n49593 = ~\pi0608  & ~n49302 ;
  assign n49594 = ~\pi0608  & ~n49298 ;
  assign n49595 = n49296 & n49594 ;
  assign n49596 = ~n49593 & ~n49595 ;
  assign n49597 = ~n49592 & ~n49596 ;
  assign n49598 = ~n49298 & ~n49585 ;
  assign n49599 = ~n49305 & ~n49589 ;
  assign n49600 = \pi1153  & ~n49599 ;
  assign n49601 = ~n49598 & n49600 ;
  assign n49602 = \pi0608  & ~n49309 ;
  assign n49603 = \pi0608  & ~n49305 ;
  assign n49604 = n49296 & n49603 ;
  assign n49605 = ~n49602 & ~n49604 ;
  assign n49606 = ~n49601 & ~n49605 ;
  assign n49607 = ~n49597 & ~n49606 ;
  assign n49608 = \pi0778  & ~n49607 ;
  assign n49609 = ~\pi0224  & ~\pi0778  ;
  assign n49610 = ~n23622 & ~n49609 ;
  assign n49611 = ~n23808 & n49610 ;
  assign n49612 = ~n23808 & n49584 ;
  assign n49613 = ~n49578 & n49612 ;
  assign n49614 = ~n49611 & ~n49613 ;
  assign n49615 = n21022 & ~n49614 ;
  assign n49616 = ~n49608 & n49615 ;
  assign n49617 = ~n20811 & ~n48879 ;
  assign n49618 = ~n48888 & n49617 ;
  assign n49619 = ~n20811 & ~n49618 ;
  assign n49620 = ~n49121 & ~n49618 ;
  assign n49621 = ~n49119 & n49620 ;
  assign n49622 = ~n49619 & ~n49621 ;
  assign n49623 = n20871 & ~n49622 ;
  assign n49624 = \pi0781  & n49623 ;
  assign n49625 = ~n22147 & ~n49115 ;
  assign n49626 = n49296 & n49625 ;
  assign n49627 = ~n22148 & ~n49626 ;
  assign n49628 = n22147 & ~n48879 ;
  assign n49629 = ~n48888 & n49628 ;
  assign n49630 = n49627 & ~n49629 ;
  assign n49631 = \pi0778  & ~n49629 ;
  assign n49632 = ~n49311 & n49631 ;
  assign n49633 = ~n49630 & ~n49632 ;
  assign n49634 = n24348 & ~n49633 ;
  assign n49635 = ~n49624 & ~n49634 ;
  assign n49636 = ~n26119 & ~n49311 ;
  assign n49637 = n26125 & ~n49313 ;
  assign n49638 = ~\pi0609  & ~n49116 ;
  assign n49639 = n49114 & n49638 ;
  assign n49640 = ~n49110 & n49639 ;
  assign n49641 = \pi0609  & ~n48879 ;
  assign n49642 = ~n48888 & n49641 ;
  assign n49643 = n20865 & ~n49642 ;
  assign n49644 = ~n49640 & n49643 ;
  assign n49645 = \pi0609  & ~n49116 ;
  assign n49646 = n49114 & n49645 ;
  assign n49647 = ~n49110 & n49646 ;
  assign n49648 = ~\pi0609  & ~n48879 ;
  assign n49649 = ~n48888 & n49648 ;
  assign n49650 = n20864 & ~n49649 ;
  assign n49651 = ~n49647 & n49650 ;
  assign n49652 = ~n49644 & ~n49651 ;
  assign n49653 = ~n49637 & n49652 ;
  assign n49654 = ~n49636 & n49653 ;
  assign n49655 = n47505 & ~n49654 ;
  assign n49656 = ~n21038 & ~n49655 ;
  assign n49657 = n49635 & n49656 ;
  assign n49658 = ~n49616 & n49657 ;
  assign n49659 = ~n23856 & ~n30434 ;
  assign n49660 = ~n49658 & n49659 ;
  assign n49661 = ~n49314 & n49323 ;
  assign n49662 = ~n49312 & n49661 ;
  assign n49663 = n21050 & ~n49662 ;
  assign n49664 = ~\pi0648  & ~n49133 ;
  assign n49665 = n20874 & ~n49146 ;
  assign n49666 = ~n49664 & ~n49665 ;
  assign n49667 = ~n49663 & n49666 ;
  assign n49668 = \pi0789  & ~n23856 ;
  assign n49669 = ~n49667 & n49668 ;
  assign n49670 = ~n49660 & ~n49669 ;
  assign n49671 = ~n21067 & ~n49670 ;
  assign n49672 = ~n49330 & n49671 ;
  assign n49673 = ~n23880 & ~n49152 ;
  assign n49674 = n49148 & n49673 ;
  assign n49675 = n23880 & ~n48879 ;
  assign n49676 = ~n48888 & n49675 ;
  assign n49677 = n20846 & ~n48879 ;
  assign n49678 = ~n48888 & n49677 ;
  assign n49679 = ~n20910 & ~n49678 ;
  assign n49680 = ~n49676 & n49679 ;
  assign n49681 = ~n49674 & n49680 ;
  assign n49682 = n20923 & ~n48889 ;
  assign n49683 = ~\pi0630  & n49682 ;
  assign n49684 = n26065 & ~n49311 ;
  assign n49685 = n26739 & ~n49313 ;
  assign n49686 = ~n23885 & n48879 ;
  assign n49687 = ~n23885 & n48882 ;
  assign n49688 = ~n47007 & n49687 ;
  assign n49689 = ~n49686 & ~n49688 ;
  assign n49690 = ~n23907 & n49689 ;
  assign n49691 = ~n49685 & n49690 ;
  assign n49692 = ~n49684 & n49691 ;
  assign n49693 = n23907 & ~n48879 ;
  assign n49694 = ~n48888 & n49693 ;
  assign n49695 = ~\pi0647  & ~n48879 ;
  assign n49696 = ~n48888 & n49695 ;
  assign n49697 = \pi1157  & ~n49696 ;
  assign n49698 = ~n49694 & n49697 ;
  assign n49699 = ~\pi0630  & n49698 ;
  assign n49700 = ~n49692 & n49699 ;
  assign n49701 = ~n49683 & ~n49700 ;
  assign n49702 = ~n24761 & n49701 ;
  assign n49703 = n20846 & ~n20910 ;
  assign n49704 = ~n48889 & n49703 ;
  assign n49705 = n21064 & ~n48889 ;
  assign n49706 = \pi0630  & n49705 ;
  assign n49707 = \pi0647  & ~n48879 ;
  assign n49708 = ~n48888 & n49707 ;
  assign n49709 = ~\pi1157  & ~n49708 ;
  assign n49710 = ~n49694 & n49709 ;
  assign n49711 = \pi0630  & n49710 ;
  assign n49712 = ~n49692 & n49711 ;
  assign n49713 = ~n49706 & ~n49712 ;
  assign n49714 = ~n49704 & n49713 ;
  assign n49715 = n49702 & n49714 ;
  assign n49716 = ~n49681 & n49715 ;
  assign n49717 = ~n29722 & ~n49716 ;
  assign n49718 = ~\pi0628  & n49689 ;
  assign n49719 = ~n49685 & n49718 ;
  assign n49720 = ~n49684 & n49719 ;
  assign n49721 = \pi0628  & ~n48879 ;
  assign n49722 = ~n48888 & n49721 ;
  assign n49723 = n20844 & ~n49722 ;
  assign n49724 = ~n49720 & n49723 ;
  assign n49725 = \pi0628  & n49689 ;
  assign n49726 = ~n49685 & n49725 ;
  assign n49727 = ~n49684 & n49726 ;
  assign n49728 = ~\pi0628  & ~n48879 ;
  assign n49729 = ~n48888 & n49728 ;
  assign n49730 = n20843 & ~n49729 ;
  assign n49731 = ~n49727 & n49730 ;
  assign n49732 = ~n49724 & ~n49731 ;
  assign n49733 = ~n21067 & ~n49732 ;
  assign n49734 = n24691 & ~n49676 ;
  assign n49735 = ~n21067 & n49734 ;
  assign n49736 = ~n49674 & n49735 ;
  assign n49737 = ~n49733 & ~n49736 ;
  assign n49738 = \pi0792  & ~n49737 ;
  assign n49739 = n27408 & ~n49738 ;
  assign n49740 = ~n49717 & n49739 ;
  assign n49741 = ~n49672 & n49740 ;
  assign n49742 = n48180 & ~n49152 ;
  assign n49743 = n49148 & n49742 ;
  assign n49744 = ~n48178 & ~n48879 ;
  assign n49745 = ~n48888 & n49744 ;
  assign n49746 = ~n23518 & ~n49745 ;
  assign n49747 = ~\pi0787  & ~n49694 ;
  assign n49748 = ~n49745 & n49747 ;
  assign n49749 = ~n49692 & n49748 ;
  assign n49750 = ~n49746 & ~n49749 ;
  assign n49751 = ~n49743 & ~n49750 ;
  assign n49752 = ~n49692 & n49698 ;
  assign n49753 = ~n49682 & ~n49752 ;
  assign n49754 = ~n49692 & n49710 ;
  assign n49755 = ~n49705 & ~n49754 ;
  assign n49756 = n49753 & n49755 ;
  assign n49757 = \pi0787  & ~n49745 ;
  assign n49758 = ~n49743 & n49757 ;
  assign n49759 = ~n49756 & n49758 ;
  assign n49760 = ~n49751 & ~n49759 ;
  assign n49761 = n45811 & n49760 ;
  assign n49762 = ~\pi0224  & ~n27408 ;
  assign n49763 = ~n49761 & ~n49762 ;
  assign n49764 = ~n49741 & n49763 ;
  assign n49765 = \pi0056  & n2404 ;
  assign n49766 = \pi0137  & n49765 ;
  assign n49767 = n2403 & n49766 ;
  assign n49768 = n1281 & n49767 ;
  assign n49769 = n1260 & n49768 ;
  assign n49770 = ~\pi0062  & n2467 ;
  assign n49771 = n2327 & n20521 ;
  assign n49772 = n1281 & n49771 ;
  assign n49773 = ~\pi0054  & ~\pi0092  ;
  assign n49774 = n1286 & n49773 ;
  assign n49775 = ~n6621 & n49774 ;
  assign n49776 = n1259 & n49775 ;
  assign n49777 = n1249 & n49776 ;
  assign n49778 = n49772 & n49777 ;
  assign n49779 = ~\pi0062  & n10015 ;
  assign n49780 = n49778 & n49779 ;
  assign n49781 = ~n49770 & ~n49780 ;
  assign n49782 = n49769 & ~n49781 ;
  assign n49783 = \pi0087  & n1259 ;
  assign n49784 = n1249 & n49783 ;
  assign n49785 = n49772 & n49784 ;
  assign n49786 = ~\pi0075  & ~n49785 ;
  assign n49787 = \pi0087  & n49786 ;
  assign n49788 = \pi0038  & ~\pi0137  ;
  assign n49789 = ~n6693 & ~n49788 ;
  assign n49790 = \pi0039  & \pi0137  ;
  assign n49791 = n1281 & n49790 ;
  assign n49792 = n1260 & n49791 ;
  assign n49793 = ~\pi0038  & ~n49792 ;
  assign n49794 = n49789 & ~n49793 ;
  assign n49795 = ~n1639 & ~n1667 ;
  assign n49796 = ~n2088 & n49795 ;
  assign n49797 = ~n1744 & n49796 ;
  assign n49798 = ~\pi0137  & ~n1694 ;
  assign n49799 = ~n2088 & n49798 ;
  assign n49800 = ~\pi0332  & ~n49799 ;
  assign n49801 = ~n49797 & n49800 ;
  assign n49802 = n1963 & ~n13614 ;
  assign n49803 = n1626 & n49802 ;
  assign n49804 = ~n1616 & n49803 ;
  assign n49805 = ~n1614 & n49804 ;
  assign n49806 = ~n1639 & ~n1655 ;
  assign n49807 = ~n1631 & n49806 ;
  assign n49808 = ~n49805 & n49807 ;
  assign n49809 = \pi0095  & n1638 ;
  assign n49810 = \pi0137  & \pi0332  ;
  assign n49811 = ~n49809 & n49810 ;
  assign n49812 = ~n49808 & n49811 ;
  assign n49813 = \pi0332  & n1694 ;
  assign n49814 = n1329 & n13614 ;
  assign n49815 = ~\pi0032  & ~n49814 ;
  assign n49816 = \pi0332  & n49815 ;
  assign n49817 = ~n1368 & n49816 ;
  assign n49818 = ~n49813 & ~n49817 ;
  assign n49819 = ~\pi0137  & ~n49818 ;
  assign n49820 = n2070 & ~n49819 ;
  assign n49821 = ~n49812 & n49820 ;
  assign n49822 = ~n49801 & n49821 ;
  assign n49823 = ~n1694 & n8675 ;
  assign n49824 = ~\pi0032  & ~n1329 ;
  assign n49825 = ~\pi0032  & \pi0096  ;
  assign n49826 = ~n8552 & n49825 ;
  assign n49827 = ~n49824 & ~n49826 ;
  assign n49828 = n49823 & n49827 ;
  assign n49829 = ~n1715 & n49828 ;
  assign n49830 = ~n1694 & ~n8675 ;
  assign n49831 = ~\pi1093  & ~n49830 ;
  assign n49832 = ~\pi0032  & ~\pi1093  ;
  assign n49833 = ~n1368 & n49832 ;
  assign n49834 = ~n49831 & ~n49833 ;
  assign n49835 = ~n49829 & ~n49834 ;
  assign n49836 = n13767 & n49835 ;
  assign n49837 = n13767 & ~n49830 ;
  assign n49838 = ~\pi0032  & n13767 ;
  assign n49839 = ~n1368 & n49838 ;
  assign n49840 = ~n49837 & ~n49839 ;
  assign n49841 = n1329 & ~n8582 ;
  assign n49842 = n49823 & n49841 ;
  assign n49843 = ~n1772 & n49842 ;
  assign n49844 = ~n1771 & n49843 ;
  assign n49845 = \pi0032  & n8675 ;
  assign n49846 = n1665 & n49845 ;
  assign n49847 = \pi1093  & ~n49846 ;
  assign n49848 = ~n49844 & n49847 ;
  assign n49849 = ~n49840 & n49848 ;
  assign n49850 = ~n49836 & ~n49849 ;
  assign n49851 = ~\pi0137  & ~n8799 ;
  assign n49852 = \pi1093  & n1694 ;
  assign n49853 = ~\pi0032  & \pi1093  ;
  assign n49854 = ~n1368 & n49853 ;
  assign n49855 = ~n49852 & ~n49854 ;
  assign n49856 = ~n49835 & n49855 ;
  assign n49857 = n49851 & ~n49856 ;
  assign n49858 = n49850 & ~n49857 ;
  assign n49859 = ~n1639 & n49858 ;
  assign n49860 = ~n1744 & n49859 ;
  assign n49861 = ~\pi0137  & n49858 ;
  assign n49862 = ~\pi0332  & ~n49861 ;
  assign n49863 = ~n49860 & n49862 ;
  assign n49864 = \pi1093  & n49815 ;
  assign n49865 = ~n1368 & n49864 ;
  assign n49866 = ~n49852 & ~n49865 ;
  assign n49867 = n49851 & ~n49866 ;
  assign n49868 = ~n1368 & n49815 ;
  assign n49869 = n49830 & ~n49868 ;
  assign n49870 = ~n49829 & ~n49869 ;
  assign n49871 = \pi0070  & n1261 ;
  assign n49872 = n1354 & n49871 ;
  assign n49873 = n1358 & n49872 ;
  assign n49874 = n8675 & n49873 ;
  assign n49875 = ~n1694 & n49874 ;
  assign n49876 = n49841 & n49875 ;
  assign n49877 = ~\pi1093  & ~n49876 ;
  assign n49878 = n49851 & n49877 ;
  assign n49879 = n49870 & n49878 ;
  assign n49880 = ~n49867 & ~n49879 ;
  assign n49881 = \pi0332  & ~n49880 ;
  assign n49882 = ~n49869 & ~n49876 ;
  assign n49883 = \pi0332  & n49882 ;
  assign n49884 = ~n49850 & n49883 ;
  assign n49885 = ~n49881 & ~n49884 ;
  assign n49886 = ~n2070 & n49885 ;
  assign n49887 = ~n49812 & n49886 ;
  assign n49888 = ~n49863 & n49887 ;
  assign n49889 = ~n49822 & ~n49888 ;
  assign n49890 = ~\pi0210  & n49889 ;
  assign n49891 = n1336 & ~n1639 ;
  assign n49892 = ~n2088 & n49891 ;
  assign n49893 = ~n1762 & n49892 ;
  assign n49894 = ~\pi0137  & n1751 ;
  assign n49895 = ~n2088 & n49894 ;
  assign n49896 = n44339 & ~n49895 ;
  assign n49897 = ~n49893 & n49896 ;
  assign n49898 = ~n1632 & n2054 ;
  assign n49899 = ~n1631 & n49898 ;
  assign n49900 = ~n49805 & n49899 ;
  assign n49901 = ~\pi0095  & ~\pi0137  ;
  assign n49902 = ~n1632 & n49901 ;
  assign n49903 = ~n49868 & n49902 ;
  assign n49904 = \pi0095  & \pi0137  ;
  assign n49905 = n1638 & n49904 ;
  assign n49906 = \pi0332  & ~n49905 ;
  assign n49907 = ~n49903 & n49906 ;
  assign n49908 = \pi0210  & n49907 ;
  assign n49909 = ~n49900 & n49908 ;
  assign n49910 = \pi0299  & ~n49909 ;
  assign n49911 = ~n49897 & n49910 ;
  assign n49912 = ~n49890 & n49911 ;
  assign n49913 = ~n49812 & ~n49819 ;
  assign n49914 = n7234 & n49913 ;
  assign n49915 = ~n49801 & n49914 ;
  assign n49916 = ~\pi0198  & ~n49915 ;
  assign n49917 = ~n49812 & n49885 ;
  assign n49918 = ~n7234 & n49917 ;
  assign n49919 = ~n49863 & n49918 ;
  assign n49920 = n49916 & ~n49919 ;
  assign n49921 = n44407 & ~n49895 ;
  assign n49922 = ~n49893 & n49921 ;
  assign n49923 = \pi0198  & n49907 ;
  assign n49924 = ~n49900 & n49923 ;
  assign n49925 = ~\pi0299  & ~n49924 ;
  assign n49926 = ~n49922 & n49925 ;
  assign n49927 = ~n49920 & n49926 ;
  assign n49928 = ~n49912 & ~n49927 ;
  assign n49929 = ~\pi0039  & n49789 ;
  assign n49930 = ~n49928 & n49929 ;
  assign n49931 = ~n49794 & ~n49930 ;
  assign n49932 = ~n6684 & n6795 ;
  assign n49933 = ~\pi0137  & ~n49932 ;
  assign n49934 = n6787 & ~n49933 ;
  assign n49935 = n1359 & n49934 ;
  assign n49936 = n49786 & ~n49935 ;
  assign n49937 = n49931 & n49936 ;
  assign n49938 = ~n49787 & ~n49937 ;
  assign n49939 = n2363 & n6784 ;
  assign n49940 = n1266 & n49939 ;
  assign n49941 = ~n49933 & n49940 ;
  assign n49942 = n1359 & n49941 ;
  assign n49943 = \pi0075  & ~n49942 ;
  assign n49944 = ~\pi0074  & ~\pi0092  ;
  assign n49945 = n1286 & n49944 ;
  assign n49946 = n1259 & n49945 ;
  assign n49947 = n1249 & n49946 ;
  assign n49948 = n49772 & n49947 ;
  assign n49949 = ~n2511 & ~n49948 ;
  assign n49950 = ~\pi0092  & ~n49949 ;
  assign n49951 = ~n49943 & n49950 ;
  assign n49952 = n49938 & n49951 ;
  assign n49953 = \pi0092  & n1286 ;
  assign n49954 = ~\pi0100  & \pi0137  ;
  assign n49955 = n1288 & n49954 ;
  assign n49956 = n49953 & n49955 ;
  assign n49957 = n1259 & n49956 ;
  assign n49958 = n1281 & n49957 ;
  assign n49959 = n1249 & n49958 ;
  assign n49960 = ~\pi0054  & ~n49959 ;
  assign n49961 = ~n49949 & ~n49960 ;
  assign n49962 = n1259 & n2324 ;
  assign n49963 = n1249 & n49962 ;
  assign n49964 = n49772 & n49963 ;
  assign n49965 = n2375 & n49964 ;
  assign n49966 = ~\pi0055  & ~n49965 ;
  assign n49967 = ~n49961 & n49966 ;
  assign n49968 = ~n49952 & n49967 ;
  assign n49969 = ~n8436 & ~n49781 ;
  assign n49970 = ~n49968 & n49969 ;
  assign n49971 = ~n49782 & ~n49970 ;
  assign n49972 = n10015 & n49778 ;
  assign n49973 = ~n2467 & ~n49972 ;
  assign n49974 = n2404 & n13466 ;
  assign n49975 = n49774 & n49974 ;
  assign n49976 = n1259 & n49975 ;
  assign n49977 = n1249 & n49976 ;
  assign n49978 = n49772 & n49977 ;
  assign n49979 = n2467 & ~n49978 ;
  assign n49980 = ~n49973 & ~n49979 ;
  assign n49981 = n49971 & ~n49980 ;
  assign n49982 = \pi0228  & \pi0231  ;
  assign n49983 = \pi0054  & ~n49982 ;
  assign n49984 = ~\pi0074  & ~n49983 ;
  assign n49985 = ~\pi0062  & ~n49982 ;
  assign n49986 = ~n8513 & n49985 ;
  assign n49987 = ~n1292 & ~n49986 ;
  assign n49988 = \pi0074  & n49982 ;
  assign n49989 = n2364 & n2375 ;
  assign n49990 = ~n49988 & ~n49989 ;
  assign n49991 = n1259 & ~n49990 ;
  assign n49992 = n1249 & n49991 ;
  assign n49993 = n6858 & n49992 ;
  assign n49994 = n2362 & n49993 ;
  assign n49995 = ~\pi0055  & ~n49988 ;
  assign n49996 = ~n49994 & n49995 ;
  assign n49997 = ~n49987 & n49996 ;
  assign n49998 = ~n49984 & n49997 ;
  assign n49999 = n1259 & n16777 ;
  assign n50000 = n1249 & n49999 ;
  assign n50001 = n6858 & n50000 ;
  assign n50002 = \pi0075  & n49982 ;
  assign n50003 = ~\pi0092  & ~n50002 ;
  assign n50004 = ~n50001 & n50003 ;
  assign n50005 = \pi0092  & ~n49982 ;
  assign n50006 = ~n8495 & n50005 ;
  assign n50007 = ~n50004 & ~n50006 ;
  assign n50008 = n1281 & n9627 ;
  assign n50009 = n1260 & n50008 ;
  assign n50010 = n8453 & n50009 ;
  assign n50011 = ~\pi0038  & n1281 ;
  assign n50012 = n1260 & n50011 ;
  assign n50013 = ~n1288 & ~n50012 ;
  assign n50014 = \pi0095  & ~n50013 ;
  assign n50015 = n1626 & ~n1630 ;
  assign n50016 = \pi0051  & ~n1868 ;
  assign n50017 = \pi0035  & n1354 ;
  assign n50018 = n1358 & n50017 ;
  assign n50019 = ~n1832 & ~n50018 ;
  assign n50020 = ~\pi0093  & ~n50018 ;
  assign n50021 = ~n1860 & n50020 ;
  assign n50022 = ~n50019 & ~n50021 ;
  assign n50023 = ~\pi0070  & ~n1868 ;
  assign n50024 = n50022 & n50023 ;
  assign n50025 = ~n50016 & ~n50024 ;
  assign n50026 = n1626 & n1963 ;
  assign n50027 = n50025 & n50026 ;
  assign n50028 = ~n50015 & ~n50027 ;
  assign n50029 = \pi0032  & ~n6688 ;
  assign n50030 = ~n6685 & n50029 ;
  assign n50031 = ~n50013 & ~n50030 ;
  assign n50032 = n50028 & n50031 ;
  assign n50033 = ~n50014 & ~n50032 ;
  assign n50034 = n1640 & n8453 ;
  assign n50035 = ~n50033 & n50034 ;
  assign n50036 = ~n50010 & ~n50035 ;
  assign n50037 = ~\pi0100  & n49982 ;
  assign n50038 = ~\pi0087  & ~n49982 ;
  assign n50039 = ~n6859 & n50038 ;
  assign n50040 = ~n2362 & ~n50039 ;
  assign n50041 = ~n50037 & ~n50040 ;
  assign n50042 = n50036 & n50041 ;
  assign n50043 = \pi0087  & ~n49982 ;
  assign n50044 = ~n8484 & n50043 ;
  assign n50045 = ~\pi0075  & ~n50044 ;
  assign n50046 = ~n50006 & n50045 ;
  assign n50047 = ~n50042 & n50046 ;
  assign n50048 = ~n50007 & ~n50047 ;
  assign n50049 = ~\pi0054  & n49997 ;
  assign n50050 = n50048 & n50049 ;
  assign n50051 = ~n49998 & ~n50050 ;
  assign n50052 = \pi0055  & ~n49982 ;
  assign n50053 = ~\pi0056  & ~n50052 ;
  assign n50054 = n1292 & ~n50053 ;
  assign n50055 = n49985 & ~n50053 ;
  assign n50056 = ~n8513 & n50055 ;
  assign n50057 = ~n50054 & ~n50056 ;
  assign n50058 = \pi0062  & ~n49982 ;
  assign n50059 = ~n8522 & n50058 ;
  assign n50060 = n50057 & ~n50059 ;
  assign n50061 = n50051 & n50060 ;
  assign n50062 = n2467 & ~n50061 ;
  assign n50063 = ~n2467 & ~n49982 ;
  assign n50064 = ~n50062 & ~n50063 ;
  assign n50065 = ~n6809 & n13028 ;
  assign n50066 = ~n6809 & n13030 ;
  assign n50067 = n1542 & n50066 ;
  assign n50068 = ~n50065 & ~n50067 ;
  assign n50069 = n1389 & ~n50068 ;
  assign n50070 = ~n13027 & n50069 ;
  assign n50071 = ~\pi0091  & ~n1391 ;
  assign n50072 = n7114 & n13053 ;
  assign n50073 = n1315 & n50072 ;
  assign n50074 = ~n13059 & n50073 ;
  assign n50075 = ~n13052 & n50074 ;
  assign n50076 = n50071 & ~n50075 ;
  assign n50077 = ~n50070 & n50076 ;
  assign n50078 = ~\pi0058  & n1323 ;
  assign n50079 = n1322 & n50078 ;
  assign n50080 = ~n7069 & n50079 ;
  assign n50081 = ~n50077 & n50080 ;
  assign n50082 = \pi0829  & ~\pi1093  ;
  assign n50083 = ~n6699 & ~n50082 ;
  assign n50084 = ~n50081 & ~n50083 ;
  assign n50085 = ~\pi0829  & ~\pi1093  ;
  assign n50086 = ~\pi0091  & \pi0824  ;
  assign n50087 = n6809 & n50086 ;
  assign n50088 = ~n1391 & n50087 ;
  assign n50089 = n50085 & n50088 ;
  assign n50090 = ~n15408 & ~n50082 ;
  assign n50091 = ~\pi0058  & n1325 ;
  assign n50092 = n1398 & n50091 ;
  assign n50093 = n1319 & n50092 ;
  assign n50094 = ~n11815 & ~n50082 ;
  assign n50095 = ~n50093 & n50094 ;
  assign n50096 = ~n50090 & ~n50095 ;
  assign n50097 = ~n6931 & n50088 ;
  assign n50098 = ~n50096 & n50097 ;
  assign n50099 = ~n50089 & ~n50098 ;
  assign n50100 = ~n50084 & n50099 ;
  assign n50101 = \pi0072  & ~n1628 ;
  assign n50102 = n2575 & ~n50101 ;
  assign n50103 = ~n6931 & ~n50096 ;
  assign n50104 = ~n6704 & ~n50085 ;
  assign n50105 = ~n50103 & n50104 ;
  assign n50106 = n1389 & ~n13052 ;
  assign n50107 = ~n13027 & n50106 ;
  assign n50108 = n50071 & ~n50107 ;
  assign n50109 = n50080 & ~n50108 ;
  assign n50110 = ~n50105 & ~n50109 ;
  assign n50111 = n50102 & ~n50110 ;
  assign n50112 = n50100 & n50111 ;
  assign n50113 = \pi0072  & n2575 ;
  assign n50114 = n1628 & n50113 ;
  assign n50115 = ~\pi0039  & ~n50114 ;
  assign n50116 = ~n50112 & n50115 ;
  assign n50117 = ~n13699 & ~n50116 ;
  assign n50118 = ~n6703 & ~n10050 ;
  assign n50119 = n1329 & n15411 ;
  assign n50120 = ~n50118 & n50119 ;
  assign n50121 = ~\pi0096  & n50120 ;
  assign n50122 = n1721 & n50120 ;
  assign n50123 = n1319 & n50122 ;
  assign n50124 = ~n50121 & ~n50123 ;
  assign n50125 = n13386 & ~n50124 ;
  assign n50126 = ~n13731 & n50125 ;
  assign n50127 = \pi1091  & ~n13630 ;
  assign n50128 = n6921 & n50127 ;
  assign n50129 = \pi0039  & ~n13627 ;
  assign n50130 = \pi0039  & ~\pi0223  ;
  assign n50131 = n2165 & n50130 ;
  assign n50132 = ~n8387 & n50131 ;
  assign n50133 = ~n50129 & ~n50132 ;
  assign n50134 = n13386 & ~n50133 ;
  assign n50135 = n50128 & n50134 ;
  assign n50136 = ~n9635 & ~n50135 ;
  assign n50137 = ~n50126 & n50136 ;
  assign n50138 = n4520 & n46110 ;
  assign n50139 = n1638 & n50138 ;
  assign n50140 = n9948 & n43150 ;
  assign n50141 = ~n50139 & ~n50140 ;
  assign n50142 = ~\pi0038  & ~\pi0039  ;
  assign n50143 = ~\pi0120  & ~n21277 ;
  assign n50144 = n6705 & n6722 ;
  assign n50145 = \pi0120  & n50144 ;
  assign n50146 = ~n50143 & ~n50145 ;
  assign n50147 = n2280 & n50146 ;
  assign n50148 = ~n6714 & ~n50143 ;
  assign n50149 = n2280 & n50148 ;
  assign n50150 = n21686 & ~n50149 ;
  assign n50151 = ~n50147 & n50150 ;
  assign n50152 = n45957 & ~n50147 ;
  assign n50153 = \pi0223  & ~n6761 ;
  assign n50154 = n50152 & n50153 ;
  assign n50155 = ~\pi0299  & ~n50154 ;
  assign n50156 = ~n50151 & n50155 ;
  assign n50157 = ~n50147 & ~n50149 ;
  assign n50158 = n22426 & n50157 ;
  assign n50159 = \pi0299  & ~n50158 ;
  assign n50160 = n22526 & n50152 ;
  assign n50161 = ~\pi0215  & n21509 ;
  assign n50162 = ~n50160 & ~n50161 ;
  assign n50163 = n50159 & n50162 ;
  assign n50164 = ~n50156 & ~n50163 ;
  assign n50165 = n1281 & ~n6736 ;
  assign n50166 = n1260 & n50165 ;
  assign n50167 = ~n17053 & ~n50166 ;
  assign n50168 = ~n6761 & n45957 ;
  assign n50169 = n50167 & n50168 ;
  assign n50170 = ~n6810 & n8648 ;
  assign n50171 = \pi1091  & ~n50170 ;
  assign n50172 = ~n21301 & n50171 ;
  assign n50173 = n1281 & ~n21295 ;
  assign n50174 = n1260 & n50173 ;
  assign n50175 = \pi1091  & n50170 ;
  assign n50176 = ~n50174 & n50175 ;
  assign n50177 = ~n50172 & ~n50176 ;
  assign n50178 = ~\pi1091  & ~n6922 ;
  assign n50179 = ~n21301 & n50178 ;
  assign n50180 = ~\pi1091  & n6922 ;
  assign n50181 = ~n50174 & n50180 ;
  assign n50182 = ~n50179 & ~n50181 ;
  assign n50183 = n50177 & n50182 ;
  assign n50184 = ~\pi0120  & n50168 ;
  assign n50185 = ~n50183 & n50184 ;
  assign n50186 = ~n50169 & ~n50185 ;
  assign n50187 = ~n2165 & n50186 ;
  assign n50188 = ~\pi0120  & ~n50183 ;
  assign n50189 = \pi0120  & ~n2280 ;
  assign n50190 = n6714 & ~n50189 ;
  assign n50191 = ~n50188 & n50190 ;
  assign n50192 = n6761 & ~n50149 ;
  assign n50193 = ~n50191 & n50192 ;
  assign n50194 = n50187 & ~n50193 ;
  assign n50195 = ~\pi0223  & n21560 ;
  assign n50196 = ~n50163 & n50195 ;
  assign n50197 = ~n50194 & n50196 ;
  assign n50198 = ~n50164 & ~n50197 ;
  assign n50199 = n50159 & ~n50160 ;
  assign n50200 = ~n6732 & n45957 ;
  assign n50201 = n50167 & n50200 ;
  assign n50202 = ~\pi0120  & n50200 ;
  assign n50203 = ~n50183 & n50202 ;
  assign n50204 = ~n50201 & ~n50203 ;
  assign n50205 = ~n2352 & n50204 ;
  assign n50206 = n6732 & ~n50149 ;
  assign n50207 = ~n50191 & n50206 ;
  assign n50208 = n50205 & ~n50207 ;
  assign n50209 = n50199 & n50208 ;
  assign n50210 = ~\pi0038  & ~n50209 ;
  assign n50211 = ~n50198 & n50210 ;
  assign n50212 = ~n50142 & ~n50211 ;
  assign n50213 = ~n50141 & n50212 ;
  assign n50214 = \pi0829  & \pi1091  ;
  assign n50215 = ~\pi0095  & n50214 ;
  assign n50216 = n13053 & n50215 ;
  assign n50217 = ~n21212 & n50216 ;
  assign n50218 = n21223 & n50217 ;
  assign n50219 = ~n6924 & n50218 ;
  assign n50220 = ~n6924 & n21215 ;
  assign n50221 = ~n21211 & n50220 ;
  assign n50222 = ~n50219 & ~n50221 ;
  assign n50223 = n1264 & n6924 ;
  assign n50224 = ~\pi0824  & ~n50214 ;
  assign n50225 = n6809 & ~n50224 ;
  assign n50226 = n1264 & ~n50225 ;
  assign n50227 = ~n50223 & ~n50226 ;
  assign n50228 = ~n21187 & ~n50227 ;
  assign n50229 = ~n21180 & n50228 ;
  assign n50230 = \pi1093  & n6684 ;
  assign n50231 = ~n50229 & n50230 ;
  assign n50232 = n50222 & n50231 ;
  assign n50233 = n1264 & ~n9012 ;
  assign n50234 = ~n21187 & n50233 ;
  assign n50235 = ~n21180 & n50234 ;
  assign n50236 = ~n6924 & n21134 ;
  assign n50237 = ~n2585 & n50236 ;
  assign n50238 = ~n21150 & n50237 ;
  assign n50239 = n21167 & n50237 ;
  assign n50240 = n21166 & n50239 ;
  assign n50241 = ~n50238 & ~n50240 ;
  assign n50242 = ~n6684 & n50241 ;
  assign n50243 = ~n21187 & n50223 ;
  assign n50244 = ~n21180 & n50243 ;
  assign n50245 = \pi1093  & ~n50244 ;
  assign n50246 = n50242 & n50245 ;
  assign n50247 = ~n50235 & n50246 ;
  assign n50248 = n1264 & ~n6811 ;
  assign n50249 = ~n21187 & n50248 ;
  assign n50250 = ~n21180 & n50249 ;
  assign n50251 = ~\pi0252  & n21186 ;
  assign n50252 = ~\pi0035  & n1320 ;
  assign n50253 = n1618 & n50252 ;
  assign n50254 = n1326 & n50253 ;
  assign n50255 = ~n1392 & n50254 ;
  assign n50256 = ~\pi0040  & ~n50255 ;
  assign n50257 = n21181 & ~n50256 ;
  assign n50258 = ~\pi0040  & ~\pi0047  ;
  assign n50259 = ~n21174 & n50258 ;
  assign n50260 = \pi0252  & ~n50259 ;
  assign n50261 = n50257 & n50260 ;
  assign n50262 = ~n50251 & ~n50261 ;
  assign n50263 = n6811 & ~n50262 ;
  assign n50264 = ~\pi1093  & ~n50263 ;
  assign n50265 = ~n50250 & n50264 ;
  assign n50266 = ~\pi0039  & ~n50141 ;
  assign n50267 = ~n50265 & n50266 ;
  assign n50268 = ~n50247 & n50267 ;
  assign n50269 = ~n50232 & n50268 ;
  assign n50270 = ~n50213 & ~n50269 ;
  assign n50271 = ~n1325 & n1858 ;
  assign n50272 = ~n1596 & n1597 ;
  assign n50273 = ~n1571 & ~n1581 ;
  assign n50274 = ~\pi0102  & ~n1529 ;
  assign n50275 = n1557 & ~n50274 ;
  assign n50276 = ~\pi0081  & n1557 ;
  assign n50277 = ~n1522 & n50276 ;
  assign n50278 = ~n50275 & ~n50277 ;
  assign n50279 = ~\pi0088  & ~\pi0098  ;
  assign n50280 = ~n50278 & n50279 ;
  assign n50281 = ~n1551 & n1557 ;
  assign n50282 = n7056 & ~n50281 ;
  assign n50283 = ~n50280 & n50282 ;
  assign n50284 = n1249 & n7059 ;
  assign n50285 = \pi0053  & n1340 ;
  assign n50286 = n1249 & n50285 ;
  assign n50287 = ~n50284 & ~n50286 ;
  assign n50288 = ~\pi0086  & n50287 ;
  assign n50289 = ~n50283 & n50288 ;
  assign n50290 = ~n1571 & ~n1574 ;
  assign n50291 = ~n50289 & n50290 ;
  assign n50292 = ~n50273 & ~n50291 ;
  assign n50293 = ~\pi0108  & n1597 ;
  assign n50294 = n50292 & n50293 ;
  assign n50295 = ~n50272 & ~n50294 ;
  assign n50296 = ~n1599 & n1858 ;
  assign n50297 = n50295 & n50296 ;
  assign n50298 = ~n50271 & ~n50297 ;
  assign n50299 = n1397 & ~n50298 ;
  assign n50300 = ~n1401 & n1858 ;
  assign n50301 = ~\pi0035  & ~\pi0093  ;
  assign n50302 = ~n50300 & n50301 ;
  assign n50303 = ~n50299 & n50302 ;
  assign n50304 = ~\pi0070  & n50303 ;
  assign n50305 = ~\pi0070  & ~n19328 ;
  assign n50306 = ~n1864 & ~n1868 ;
  assign n50307 = ~n50305 & n50306 ;
  assign n50308 = ~n50304 & n50307 ;
  assign n50309 = ~\pi1082  & n1621 ;
  assign n50310 = ~\pi0032  & ~n50309 ;
  assign n50311 = \pi0051  & n1867 ;
  assign n50312 = n1963 & ~n50311 ;
  assign n50313 = n50310 & n50312 ;
  assign n50314 = ~n50308 & n50313 ;
  assign n50315 = ~n1630 & n50310 ;
  assign n50316 = ~n1639 & ~n2589 ;
  assign n50317 = ~n50315 & n50316 ;
  assign n50318 = ~n50314 & n50317 ;
  assign n50319 = n1288 & ~n49809 ;
  assign n50320 = ~n50318 & n50319 ;
  assign n50321 = \pi0039  & ~n2280 ;
  assign n50322 = n8381 & n8387 ;
  assign n50323 = n6716 & n6917 ;
  assign n50324 = ~n6702 & n50323 ;
  assign n50325 = ~n6704 & n6809 ;
  assign n50326 = n50324 & n50325 ;
  assign n50327 = ~n50322 & n50326 ;
  assign n50328 = \pi0039  & n11859 ;
  assign n50329 = n6716 & n6718 ;
  assign n50330 = n50328 & n50329 ;
  assign n50331 = ~n50327 & n50330 ;
  assign n50332 = ~n50321 & ~n50331 ;
  assign n50333 = ~\pi0038  & ~n50332 ;
  assign n50334 = n1638 & n6629 ;
  assign n50335 = \pi0087  & ~n50334 ;
  assign n50336 = ~n6693 & ~n50335 ;
  assign n50337 = ~n50333 & n50336 ;
  assign n50338 = ~n50320 & n50337 ;
  assign n50339 = ~\pi0087  & n6789 ;
  assign n50340 = \pi0087  & n6629 ;
  assign n50341 = n1638 & n50340 ;
  assign n50342 = ~n50339 & ~n50341 ;
  assign n50343 = n7265 & n50342 ;
  assign n50344 = ~n50338 & n50343 ;
  assign n50345 = ~\pi0054  & ~n8421 ;
  assign n50346 = ~n8412 & n19402 ;
  assign n50347 = ~n50345 & n50346 ;
  assign n50348 = ~n50344 & n50347 ;
  assign n50349 = \pi0055  & ~\pi0074  ;
  assign n50350 = n6630 & n50349 ;
  assign n50351 = n1638 & n50350 ;
  assign n50352 = ~\pi0055  & \pi0074  ;
  assign n50353 = n6630 & n50352 ;
  assign n50354 = n1638 & n50353 ;
  assign n50355 = ~n50351 & ~n50354 ;
  assign n50356 = n1292 & n2467 ;
  assign n50357 = n50355 & n50356 ;
  assign n50358 = ~n50348 & n50357 ;
  assign n50359 = n2467 & ~n19403 ;
  assign n50360 = ~n8441 & ~n50359 ;
  assign n50361 = ~n50358 & n50360 ;
  assign n50362 = ~\pi0230  & ~\pi0233  ;
  assign n50363 = \pi0199  & ~\pi1153  ;
  assign n50364 = n44032 & ~n50363 ;
  assign n50365 = ~\pi0199  & ~\pi1155  ;
  assign n50366 = \pi0207  & ~\pi1154  ;
  assign n50367 = ~n50365 & n50366 ;
  assign n50368 = n50364 & n50367 ;
  assign n50369 = \pi0208  & n50368 ;
  assign n50370 = \pi0199  & \pi0200  ;
  assign n50371 = ~n12691 & ~n50370 ;
  assign n50372 = ~\pi0299  & ~n50363 ;
  assign n50373 = n50371 & n50372 ;
  assign n50374 = \pi1155  & ~n13558 ;
  assign n50375 = ~\pi0299  & ~n50374 ;
  assign n50376 = ~n50373 & n50375 ;
  assign n50377 = \pi0207  & \pi1154  ;
  assign n50378 = \pi0208  & n50377 ;
  assign n50379 = ~n50376 & n50378 ;
  assign n50380 = ~n50369 & ~n50379 ;
  assign n50381 = ~\pi0207  & \pi0208  ;
  assign n50382 = \pi1155  & n13645 ;
  assign n50383 = \pi0199  & ~\pi0200  ;
  assign n50384 = ~\pi0299  & ~n50383 ;
  assign n50385 = ~n50382 & n50384 ;
  assign n50386 = \pi1154  & ~n50385 ;
  assign n50387 = ~\pi0199  & \pi1155  ;
  assign n50388 = n44035 & n50387 ;
  assign n50389 = ~\pi1154  & ~n50388 ;
  assign n50390 = ~\pi0299  & ~n12691 ;
  assign n50391 = \pi0200  & ~n50387 ;
  assign n50392 = n50390 & ~n50391 ;
  assign n50393 = ~n50389 & n50392 ;
  assign n50394 = \pi0200  & ~\pi1155  ;
  assign n50395 = \pi1156  & n13550 ;
  assign n50396 = ~n50394 & n50395 ;
  assign n50397 = ~n50393 & ~n50396 ;
  assign n50398 = ~n50386 & n50397 ;
  assign n50399 = n50381 & ~n50398 ;
  assign n50400 = n50380 & ~n50399 ;
  assign n50401 = ~\pi0299  & ~\pi1156  ;
  assign n50402 = ~\pi0200  & \pi1155  ;
  assign n50403 = n13558 & ~n50402 ;
  assign n50404 = ~n50401 & ~n50403 ;
  assign n50405 = \pi0199  & ~\pi1155  ;
  assign n50406 = ~\pi0200  & ~\pi1156  ;
  assign n50407 = ~n50405 & n50406 ;
  assign n50408 = \pi0207  & ~n50407 ;
  assign n50409 = ~n50404 & n50408 ;
  assign n50410 = ~\pi0207  & ~\pi0299  ;
  assign n50411 = ~\pi0208  & ~n50410 ;
  assign n50412 = \pi0299  & ~\pi1154  ;
  assign n50413 = \pi1157  & ~n50412 ;
  assign n50414 = n50411 & n50413 ;
  assign n50415 = ~n50409 & n50414 ;
  assign n50416 = \pi0299  & \pi1154  ;
  assign n50417 = ~\pi0208  & n50416 ;
  assign n50418 = \pi0207  & ~\pi0208  ;
  assign n50419 = ~\pi0299  & \pi1155  ;
  assign n50420 = n50383 & n50419 ;
  assign n50421 = ~\pi1156  & ~n50420 ;
  assign n50422 = ~\pi0299  & ~n50405 ;
  assign n50423 = n50371 & n50422 ;
  assign n50424 = ~n50421 & n50423 ;
  assign n50425 = n50418 & n50424 ;
  assign n50426 = ~n50417 & ~n50425 ;
  assign n50427 = ~\pi1157  & ~n50426 ;
  assign n50428 = ~n50415 & ~n50427 ;
  assign n50429 = n50400 & n50428 ;
  assign n50430 = \pi0211  & \pi0214  ;
  assign n50431 = ~n50429 & n50430 ;
  assign n50432 = ~\pi0299  & ~n50371 ;
  assign n50433 = ~\pi1155  & ~n13550 ;
  assign n50434 = ~n50432 & ~n50433 ;
  assign n50435 = \pi0299  & \pi1155  ;
  assign n50436 = ~\pi0207  & ~n50435 ;
  assign n50437 = ~\pi0208  & ~n50436 ;
  assign n50438 = \pi1155  & n50383 ;
  assign n50439 = n50401 & ~n50438 ;
  assign n50440 = n50437 & ~n50439 ;
  assign n50441 = n50434 & n50440 ;
  assign n50442 = ~\pi0211  & ~\pi0214  ;
  assign n50443 = ~n50430 & ~n50442 ;
  assign n50444 = n50441 & n50443 ;
  assign n50445 = \pi0207  & ~n50395 ;
  assign n50446 = ~n50436 & ~n50445 ;
  assign n50447 = ~n50383 & n50401 ;
  assign n50448 = ~\pi1155  & ~n50447 ;
  assign n50449 = ~n44035 & ~n50436 ;
  assign n50450 = ~n50448 & n50449 ;
  assign n50451 = ~n50446 & ~n50450 ;
  assign n50452 = ~\pi0208  & \pi1157  ;
  assign n50453 = n50443 & n50452 ;
  assign n50454 = ~n50451 & n50453 ;
  assign n50455 = ~n50444 & ~n50454 ;
  assign n50456 = ~n50373 & ~n50374 ;
  assign n50457 = \pi1154  & ~n50456 ;
  assign n50458 = ~\pi0299  & ~\pi1155  ;
  assign n50459 = n50383 & n50458 ;
  assign n50460 = \pi1153  & ~\pi1154  ;
  assign n50461 = n50459 & n50460 ;
  assign n50462 = ~\pi1153  & n13558 ;
  assign n50463 = ~\pi1154  & \pi1155  ;
  assign n50464 = ~n44035 & n50463 ;
  assign n50465 = ~n50462 & n50464 ;
  assign n50466 = ~n50461 & ~n50465 ;
  assign n50467 = \pi0207  & n50466 ;
  assign n50468 = ~n50457 & n50467 ;
  assign n50469 = ~n50396 & n50436 ;
  assign n50470 = ~n50393 & n50469 ;
  assign n50471 = \pi0208  & n50443 ;
  assign n50472 = ~n50470 & n50471 ;
  assign n50473 = ~n50468 & n50472 ;
  assign n50474 = n50455 & ~n50473 ;
  assign n50475 = ~\pi0299  & \pi1156  ;
  assign n50476 = ~n13645 & n50475 ;
  assign n50477 = ~n50438 & n50476 ;
  assign n50478 = n50418 & ~n50421 ;
  assign n50479 = ~n50477 & n50478 ;
  assign n50480 = ~\pi0208  & \pi0299  ;
  assign n50481 = ~n50421 & n50480 ;
  assign n50482 = ~n50479 & ~n50481 ;
  assign n50483 = \pi0299  & \pi1156  ;
  assign n50484 = n50452 & n50483 ;
  assign n50485 = ~n50370 & ~n50405 ;
  assign n50486 = n50475 & n50485 ;
  assign n50487 = ~\pi0200  & ~n50405 ;
  assign n50488 = n50401 & n50487 ;
  assign n50489 = ~n50486 & ~n50488 ;
  assign n50490 = \pi0207  & n50452 ;
  assign n50491 = ~n50489 & n50490 ;
  assign n50492 = ~n50484 & ~n50491 ;
  assign n50493 = n50482 & n50492 ;
  assign n50494 = ~\pi0199  & \pi1156  ;
  assign n50495 = ~n50394 & n50494 ;
  assign n50496 = ~n50483 & ~n50495 ;
  assign n50497 = ~\pi0207  & n50496 ;
  assign n50498 = ~n50393 & n50497 ;
  assign n50499 = \pi0207  & ~n50483 ;
  assign n50500 = \pi0208  & ~n50499 ;
  assign n50501 = ~n50498 & n50500 ;
  assign n50502 = ~\pi1153  & ~n13550 ;
  assign n50503 = \pi1154  & n50371 ;
  assign n50504 = ~n50502 & n50503 ;
  assign n50505 = ~\pi1154  & ~n50365 ;
  assign n50506 = n50364 & n50505 ;
  assign n50507 = n13550 & n50402 ;
  assign n50508 = ~n50506 & ~n50507 ;
  assign n50509 = ~n50504 & n50508 ;
  assign n50510 = ~\pi1153  & \pi1154  ;
  assign n50511 = ~\pi0299  & \pi1154  ;
  assign n50512 = ~n50370 & n50511 ;
  assign n50513 = ~n50510 & ~n50512 ;
  assign n50514 = ~n50506 & n50513 ;
  assign n50515 = n12409 & ~n50514 ;
  assign n50516 = ~n50509 & n50515 ;
  assign n50517 = ~n50501 & ~n50516 ;
  assign n50518 = n50493 & n50517 ;
  assign n50519 = n50442 & ~n50518 ;
  assign n50520 = n50474 & ~n50519 ;
  assign n50521 = ~n50431 & n50520 ;
  assign n50522 = \pi0212  & ~n50521 ;
  assign n50523 = \pi0207  & ~n50514 ;
  assign n50524 = ~n50509 & n50523 ;
  assign n50525 = \pi0208  & ~n50396 ;
  assign n50526 = ~n50393 & n50525 ;
  assign n50527 = ~n12409 & ~n50526 ;
  assign n50528 = ~\pi1157  & ~n50527 ;
  assign n50529 = ~n50524 & n50528 ;
  assign n50530 = \pi0207  & n50424 ;
  assign n50531 = ~\pi0208  & ~\pi1157  ;
  assign n50532 = ~n50530 & n50531 ;
  assign n50533 = ~n50529 & ~n50532 ;
  assign n50534 = \pi1157  & ~n50411 ;
  assign n50535 = \pi0207  & \pi1157  ;
  assign n50536 = ~n50407 & n50535 ;
  assign n50537 = ~n50404 & n50536 ;
  assign n50538 = ~n50534 & ~n50537 ;
  assign n50539 = ~\pi0299  & ~n50382 ;
  assign n50540 = n50496 & n50539 ;
  assign n50541 = ~n50386 & n50540 ;
  assign n50542 = ~\pi0207  & n50541 ;
  assign n50543 = \pi1153  & ~n50384 ;
  assign n50544 = \pi0207  & ~\pi0299  ;
  assign n50545 = ~n50507 & n50544 ;
  assign n50546 = ~n50543 & n50545 ;
  assign n50547 = ~n50504 & n50546 ;
  assign n50548 = \pi0208  & ~n50547 ;
  assign n50549 = ~n50542 & n50548 ;
  assign n50550 = ~n50538 & ~n50549 ;
  assign n50551 = ~\pi0211  & ~n50550 ;
  assign n50552 = n50533 & n50551 ;
  assign n50553 = \pi0211  & ~n50518 ;
  assign n50554 = \pi0214  & ~n50553 ;
  assign n50555 = ~n50552 & n50554 ;
  assign n50556 = ~\pi0212  & \pi0214  ;
  assign n50557 = ~\pi1157  & ~n50532 ;
  assign n50558 = ~n50524 & ~n50527 ;
  assign n50559 = \pi0207  & ~n50489 ;
  assign n50560 = ~\pi0208  & ~n50559 ;
  assign n50561 = ~n50532 & ~n50560 ;
  assign n50562 = ~n50558 & n50561 ;
  assign n50563 = ~n50557 & ~n50562 ;
  assign n50564 = ~\pi0212  & ~n50529 ;
  assign n50565 = ~n50563 & n50564 ;
  assign n50566 = ~n50556 & ~n50565 ;
  assign n50567 = ~n50555 & ~n50566 ;
  assign n50568 = ~n50522 & ~n50567 ;
  assign n50569 = n46751 & ~n50568 ;
  assign n50570 = ~\pi0212  & ~\pi0214  ;
  assign n50571 = ~\pi0211  & ~n50570 ;
  assign n50572 = \pi0219  & n50571 ;
  assign n50573 = \pi0219  & ~n50529 ;
  assign n50574 = ~n50563 & n50573 ;
  assign n50575 = ~n50572 & ~n50574 ;
  assign n50576 = \pi0211  & n9948 ;
  assign n50577 = \pi0208  & ~n50470 ;
  assign n50578 = ~n50468 & n50577 ;
  assign n50579 = ~n50451 & n50452 ;
  assign n50580 = ~n50441 & n50556 ;
  assign n50581 = ~n50579 & n50580 ;
  assign n50582 = ~n50578 & n50581 ;
  assign n50583 = ~n50507 & ~n50543 ;
  assign n50584 = ~n50504 & n50583 ;
  assign n50585 = \pi0207  & ~n50584 ;
  assign n50586 = \pi0299  & ~\pi1153  ;
  assign n50587 = ~\pi0207  & ~n50586 ;
  assign n50588 = ~n50541 & n50587 ;
  assign n50589 = ~n50585 & ~n50588 ;
  assign n50590 = \pi0208  & ~n50589 ;
  assign n50591 = ~n50421 & ~n50477 ;
  assign n50592 = n50418 & n50591 ;
  assign n50593 = ~\pi1157  & ~n50480 ;
  assign n50594 = ~n50592 & n50593 ;
  assign n50595 = n50538 & ~n50586 ;
  assign n50596 = ~n50594 & n50595 ;
  assign n50597 = n12255 & ~n50596 ;
  assign n50598 = ~n50590 & n50597 ;
  assign n50599 = ~n50582 & ~n50598 ;
  assign n50600 = \pi0212  & ~\pi0214  ;
  assign n50601 = ~n50415 & n50600 ;
  assign n50602 = ~n50427 & n50601 ;
  assign n50603 = n50400 & n50602 ;
  assign n50604 = n9948 & ~n50603 ;
  assign n50605 = n50599 & n50604 ;
  assign n50606 = ~n50576 & ~n50605 ;
  assign n50607 = ~n50575 & ~n50606 ;
  assign n50608 = ~\pi0211  & \pi1155  ;
  assign n50609 = \pi0211  & \pi1154  ;
  assign n50610 = ~n50608 & ~n50609 ;
  assign n50611 = n12255 & ~n50610 ;
  assign n50612 = ~\pi0211  & \pi1156  ;
  assign n50613 = \pi0211  & \pi1155  ;
  assign n50614 = ~n50612 & ~n50613 ;
  assign n50615 = n50600 & ~n50614 ;
  assign n50616 = ~n50611 & ~n50615 ;
  assign n50617 = ~\pi0211  & \pi1157  ;
  assign n50618 = \pi0211  & \pi1156  ;
  assign n50619 = ~n50617 & ~n50618 ;
  assign n50620 = n50556 & ~n50619 ;
  assign n50621 = ~\pi0219  & ~n50620 ;
  assign n50622 = n50616 & n50621 ;
  assign n50623 = \pi0214  & n50608 ;
  assign n50624 = ~\pi0212  & ~n50623 ;
  assign n50625 = ~\pi0211  & \pi1153  ;
  assign n50626 = n12255 & ~n50625 ;
  assign n50627 = ~\pi0211  & \pi1154  ;
  assign n50628 = ~\pi0214  & ~n50627 ;
  assign n50629 = ~n50626 & ~n50628 ;
  assign n50630 = ~n50624 & n50629 ;
  assign n50631 = \pi0219  & ~n50630 ;
  assign n50632 = ~n27408 & ~n50631 ;
  assign n50633 = ~n50622 & n50632 ;
  assign n50634 = ~\pi0213  & ~n50633 ;
  assign n50635 = \pi0199  & \pi1142  ;
  assign n50636 = ~\pi0200  & ~n50635 ;
  assign n50637 = ~\pi0199  & \pi1143  ;
  assign n50638 = n50636 & ~n50637 ;
  assign n50639 = ~\pi0199  & \pi1142  ;
  assign n50640 = \pi0200  & ~n50639 ;
  assign n50641 = \pi0208  & n50544 ;
  assign n50642 = ~n50640 & n50641 ;
  assign n50643 = ~n50638 & n50642 ;
  assign n50644 = ~\pi0199  & \pi1144  ;
  assign n50645 = ~\pi0299  & ~n50644 ;
  assign n50646 = n50636 & n50645 ;
  assign n50647 = n44035 & ~n50637 ;
  assign n50648 = n50381 & ~n50647 ;
  assign n50649 = ~n50646 & n50648 ;
  assign n50650 = ~n50643 & ~n50649 ;
  assign n50651 = n50636 & ~n50644 ;
  assign n50652 = \pi0200  & ~n50637 ;
  assign n50653 = n50418 & ~n50652 ;
  assign n50654 = ~n50651 & n50653 ;
  assign n50655 = n50650 & ~n50654 ;
  assign n50656 = n20516 & ~n50655 ;
  assign n50657 = \pi0211  & \pi1143  ;
  assign n50658 = ~\pi0211  & \pi1144  ;
  assign n50659 = ~n50657 & ~n50658 ;
  assign n50660 = ~n12255 & ~n50659 ;
  assign n50661 = ~\pi0211  & \pi1143  ;
  assign n50662 = n12255 & n50661 ;
  assign n50663 = \pi0211  & \pi1142  ;
  assign n50664 = n12255 & n50663 ;
  assign n50665 = ~n50662 & ~n50664 ;
  assign n50666 = ~n50660 & n50665 ;
  assign n50667 = ~\pi0219  & n50666 ;
  assign n50668 = ~\pi0211  & \pi1142  ;
  assign n50669 = \pi0219  & ~n50668 ;
  assign n50670 = ~\pi0057  & \pi0299  ;
  assign n50671 = ~n50570 & n50670 ;
  assign n50672 = n6848 & n50671 ;
  assign n50673 = ~n50669 & n50672 ;
  assign n50674 = ~n50667 & n50673 ;
  assign n50675 = ~n50656 & ~n50674 ;
  assign n50676 = \pi0219  & ~n50571 ;
  assign n50677 = ~n9948 & ~n50676 ;
  assign n50678 = \pi0213  & ~n50677 ;
  assign n50679 = ~n12255 & ~n50570 ;
  assign n50680 = ~n50659 & n50679 ;
  assign n50681 = ~n50662 & ~n50680 ;
  assign n50682 = ~\pi0219  & ~n50681 ;
  assign n50683 = \pi0219  & \pi1142  ;
  assign n50684 = ~n50664 & ~n50683 ;
  assign n50685 = \pi0213  & n50684 ;
  assign n50686 = ~n50682 & n50685 ;
  assign n50687 = ~n50678 & ~n50686 ;
  assign n50688 = n50675 & ~n50687 ;
  assign n50689 = ~\pi0211  & \pi0219  ;
  assign n50690 = n50435 & n50556 ;
  assign n50691 = n50689 & n50690 ;
  assign n50692 = ~\pi0214  & n50416 ;
  assign n50693 = \pi0214  & \pi0299  ;
  assign n50694 = \pi1153  & n50693 ;
  assign n50695 = ~n50692 & ~n50694 ;
  assign n50696 = \pi0212  & n50689 ;
  assign n50697 = ~n50695 & n50696 ;
  assign n50698 = ~n50691 & ~n50697 ;
  assign n50699 = n27408 & ~n50698 ;
  assign n50700 = n50616 & ~n50620 ;
  assign n50701 = ~\pi0219  & \pi0299  ;
  assign n50702 = n27408 & n50701 ;
  assign n50703 = ~n50700 & n50702 ;
  assign n50704 = ~n50699 & ~n50703 ;
  assign n50705 = ~n50656 & n50704 ;
  assign n50706 = n50634 & n50705 ;
  assign n50707 = ~n50688 & ~n50706 ;
  assign n50708 = \pi0209  & n50707 ;
  assign n50709 = n50634 & ~n50708 ;
  assign n50710 = ~n50607 & n50709 ;
  assign n50711 = ~n50569 & n50710 ;
  assign n50712 = ~n50529 & ~n50563 ;
  assign n50713 = \pi0211  & \pi0219  ;
  assign n50714 = ~n50570 & ~n50713 ;
  assign n50715 = ~n50712 & ~n50714 ;
  assign n50716 = n50538 & ~n50594 ;
  assign n50717 = \pi0299  & ~\pi1142  ;
  assign n50718 = n50716 & ~n50717 ;
  assign n50719 = n50466 & n50544 ;
  assign n50720 = ~n50457 & n50719 ;
  assign n50721 = ~n50386 & n50496 ;
  assign n50722 = ~n50382 & n50410 ;
  assign n50723 = ~\pi1154  & ~\pi1156  ;
  assign n50724 = ~\pi0207  & ~n50723 ;
  assign n50725 = ~n50722 & ~n50724 ;
  assign n50726 = n50721 & ~n50725 ;
  assign n50727 = ~n50720 & ~n50726 ;
  assign n50728 = \pi0208  & ~n50717 ;
  assign n50729 = n50727 & n50728 ;
  assign n50730 = ~n50718 & ~n50729 ;
  assign n50731 = ~n12257 & n50714 ;
  assign n50732 = n50730 & n50731 ;
  assign n50733 = n27408 & ~n50732 ;
  assign n50734 = ~n50715 & n50733 ;
  assign n50735 = \pi1154  & ~n50459 ;
  assign n50736 = \pi0299  & ~\pi1143  ;
  assign n50737 = ~n50458 & ~n50736 ;
  assign n50738 = ~n50432 & n50737 ;
  assign n50739 = n50735 & ~n50738 ;
  assign n50740 = \pi0299  & \pi1143  ;
  assign n50741 = ~\pi1154  & ~n50740 ;
  assign n50742 = ~n50388 & n50741 ;
  assign n50743 = ~\pi1156  & ~n50742 ;
  assign n50744 = ~n50739 & n50743 ;
  assign n50745 = \pi0200  & \pi1154  ;
  assign n50746 = ~n50387 & n50745 ;
  assign n50747 = ~n50416 & ~n50746 ;
  assign n50748 = ~n50740 & ~n50747 ;
  assign n50749 = n43637 & ~n50394 ;
  assign n50750 = n50741 & ~n50749 ;
  assign n50751 = \pi1156  & ~n50750 ;
  assign n50752 = ~n50748 & n50751 ;
  assign n50753 = ~\pi0207  & ~n50752 ;
  assign n50754 = ~n50744 & n50753 ;
  assign n50755 = \pi0207  & ~n50740 ;
  assign n50756 = \pi0208  & ~n50755 ;
  assign n50757 = \pi0208  & ~n50514 ;
  assign n50758 = ~n50509 & n50757 ;
  assign n50759 = ~n50756 & ~n50758 ;
  assign n50760 = ~n50754 & ~n50759 ;
  assign n50761 = n50480 & ~n50736 ;
  assign n50762 = n50418 & ~n50736 ;
  assign n50763 = n50591 & n50762 ;
  assign n50764 = ~n50761 & ~n50763 ;
  assign n50765 = ~\pi1157  & ~n50764 ;
  assign n50766 = ~\pi0299  & ~n50487 ;
  assign n50767 = ~n50486 & n50766 ;
  assign n50768 = \pi0207  & ~n50736 ;
  assign n50769 = n50452 & n50768 ;
  assign n50770 = ~n50767 & n50769 ;
  assign n50771 = n50452 & n50740 ;
  assign n50772 = ~\pi0211  & n12255 ;
  assign n50773 = \pi0211  & n50679 ;
  assign n50774 = ~n50772 & ~n50773 ;
  assign n50775 = ~n50771 & ~n50774 ;
  assign n50776 = ~n50770 & n50775 ;
  assign n50777 = ~n50765 & n50776 ;
  assign n50778 = ~n50760 & n50777 ;
  assign n50779 = \pi0299  & ~\pi1144  ;
  assign n50780 = ~n50458 & ~n50779 ;
  assign n50781 = ~n50432 & n50780 ;
  assign n50782 = n50735 & ~n50781 ;
  assign n50783 = \pi0299  & \pi1144  ;
  assign n50784 = ~\pi1154  & ~n50783 ;
  assign n50785 = ~n50388 & n50784 ;
  assign n50786 = ~\pi1156  & ~n50785 ;
  assign n50787 = ~n50782 & n50786 ;
  assign n50788 = ~n50747 & ~n50783 ;
  assign n50789 = ~n50749 & n50784 ;
  assign n50790 = \pi1156  & ~n50789 ;
  assign n50791 = ~n50788 & n50790 ;
  assign n50792 = ~\pi0207  & ~n50791 ;
  assign n50793 = ~n50787 & n50792 ;
  assign n50794 = \pi0207  & ~n50783 ;
  assign n50795 = \pi0208  & ~n50794 ;
  assign n50796 = ~n50758 & ~n50795 ;
  assign n50797 = ~n50793 & ~n50796 ;
  assign n50798 = n50480 & ~n50779 ;
  assign n50799 = n50418 & ~n50779 ;
  assign n50800 = n50591 & n50799 ;
  assign n50801 = ~n50798 & ~n50800 ;
  assign n50802 = ~\pi1157  & ~n50801 ;
  assign n50803 = n50490 & ~n50779 ;
  assign n50804 = ~n50767 & n50803 ;
  assign n50805 = ~\pi0211  & n50679 ;
  assign n50806 = n50452 & n50783 ;
  assign n50807 = n50805 & ~n50806 ;
  assign n50808 = ~n50804 & n50807 ;
  assign n50809 = ~n50802 & n50808 ;
  assign n50810 = ~n50797 & n50809 ;
  assign n50811 = ~n50778 & ~n50810 ;
  assign n50812 = ~\pi0219  & ~n50811 ;
  assign n50813 = ~\pi0209  & ~n50812 ;
  assign n50814 = n50734 & n50813 ;
  assign n50815 = ~\pi0209  & ~n50678 ;
  assign n50816 = ~n50686 & n50815 ;
  assign n50817 = ~n50708 & ~n50816 ;
  assign n50818 = ~n50814 & n50817 ;
  assign n50819 = \pi0230  & ~n50818 ;
  assign n50820 = ~n50711 & n50819 ;
  assign n50821 = ~n50362 & ~n50820 ;
  assign n50822 = ~\pi0230  & ~\pi0234  ;
  assign n50823 = ~\pi1154  & ~n50507 ;
  assign n50824 = ~\pi0299  & ~n50370 ;
  assign n50825 = ~\pi1155  & n12691 ;
  assign n50826 = n50824 & ~n50825 ;
  assign n50827 = ~n50823 & n50826 ;
  assign n50828 = \pi0207  & ~n50435 ;
  assign n50829 = ~n50827 & n50828 ;
  assign n50830 = ~\pi0211  & ~n50829 ;
  assign n50831 = n50577 & n50830 ;
  assign n50832 = ~n50396 & ~n50435 ;
  assign n50833 = ~n50393 & n50832 ;
  assign n50834 = ~\pi0211  & n50437 ;
  assign n50835 = ~n50833 & n50834 ;
  assign n50836 = \pi0214  & ~n50835 ;
  assign n50837 = ~n50831 & n50836 ;
  assign n50838 = ~\pi0207  & ~n50386 ;
  assign n50839 = n50397 & n50838 ;
  assign n50840 = ~\pi0299  & n50370 ;
  assign n50841 = n12691 & n50458 ;
  assign n50842 = ~n50840 & ~n50841 ;
  assign n50843 = ~n50823 & n50842 ;
  assign n50844 = \pi0207  & ~n50843 ;
  assign n50845 = \pi0208  & \pi0211  ;
  assign n50846 = ~n50844 & n50845 ;
  assign n50847 = ~n50839 & n50846 ;
  assign n50848 = ~\pi0207  & n50416 ;
  assign n50849 = ~n50386 & ~n50848 ;
  assign n50850 = n50397 & n50849 ;
  assign n50851 = ~\pi0207  & ~n50416 ;
  assign n50852 = ~\pi0208  & \pi0211  ;
  assign n50853 = ~n50851 & n50852 ;
  assign n50854 = ~n50850 & n50853 ;
  assign n50855 = ~n50847 & ~n50854 ;
  assign n50856 = n50837 & n50855 ;
  assign n50857 = \pi0212  & ~n50856 ;
  assign n50858 = n50437 & ~n50833 ;
  assign n50859 = \pi0211  & n50858 ;
  assign n50860 = \pi0211  & ~n50829 ;
  assign n50861 = n50577 & n50860 ;
  assign n50862 = ~n50859 & ~n50861 ;
  assign n50863 = \pi0211  & ~\pi0214  ;
  assign n50864 = n12409 & n50827 ;
  assign n50865 = ~n50501 & ~n50864 ;
  assign n50866 = ~n50393 & n50496 ;
  assign n50867 = ~\pi0207  & ~n50483 ;
  assign n50868 = ~\pi0208  & ~n50867 ;
  assign n50869 = ~n50866 & n50868 ;
  assign n50870 = ~\pi0214  & ~n50869 ;
  assign n50871 = n50865 & n50870 ;
  assign n50872 = ~n50863 & ~n50871 ;
  assign n50873 = n50862 & ~n50872 ;
  assign n50874 = n50857 & ~n50873 ;
  assign n50875 = \pi0207  & n50827 ;
  assign n50876 = ~\pi0207  & ~\pi0208  ;
  assign n50877 = ~n12409 & ~n50876 ;
  assign n50878 = ~\pi0214  & ~n50877 ;
  assign n50879 = ~n50875 & n50878 ;
  assign n50880 = ~\pi0214  & ~n12409 ;
  assign n50881 = ~n50396 & n50880 ;
  assign n50882 = ~n50393 & n50881 ;
  assign n50883 = ~\pi0212  & ~n50882 ;
  assign n50884 = ~n50879 & n50883 ;
  assign n50885 = n50865 & ~n50869 ;
  assign n50886 = ~\pi0211  & ~n50885 ;
  assign n50887 = \pi0214  & n50862 ;
  assign n50888 = ~n50886 & n50887 ;
  assign n50889 = n50884 & ~n50888 ;
  assign n50890 = ~n50874 & ~n50889 ;
  assign n50891 = ~\pi0219  & n50890 ;
  assign n50892 = ~\pi0057  & \pi0213  ;
  assign n50893 = n6848 & n50892 ;
  assign n50894 = ~n50875 & ~n50877 ;
  assign n50895 = ~n12409 & ~n50396 ;
  assign n50896 = ~n50393 & n50895 ;
  assign n50897 = ~n50571 & ~n50896 ;
  assign n50898 = ~n50894 & n50897 ;
  assign n50899 = \pi0219  & ~n50898 ;
  assign n50900 = n50893 & ~n50899 ;
  assign n50901 = \pi0208  & ~\pi0211  ;
  assign n50902 = ~n50844 & n50901 ;
  assign n50903 = ~n50839 & n50902 ;
  assign n50904 = ~\pi0208  & ~\pi0211  ;
  assign n50905 = ~n50851 & n50904 ;
  assign n50906 = ~n50850 & n50905 ;
  assign n50907 = ~n50903 & ~n50906 ;
  assign n50908 = ~n50570 & n50892 ;
  assign n50909 = n6848 & n50908 ;
  assign n50910 = ~n50907 & n50909 ;
  assign n50911 = ~n50900 & ~n50910 ;
  assign n50912 = ~n50891 & ~n50911 ;
  assign n50913 = ~\pi0214  & ~n50907 ;
  assign n50914 = \pi0207  & n50541 ;
  assign n50915 = n50411 & ~n50914 ;
  assign n50916 = n50544 & ~n50843 ;
  assign n50917 = \pi0208  & ~n50916 ;
  assign n50918 = ~n50542 & n50917 ;
  assign n50919 = ~n50915 & ~n50918 ;
  assign n50920 = \pi0211  & ~n50586 ;
  assign n50921 = ~\pi0214  & n50920 ;
  assign n50922 = ~n50919 & n50921 ;
  assign n50923 = ~n50913 & ~n50922 ;
  assign n50924 = \pi0211  & ~n50877 ;
  assign n50925 = ~n50875 & n50924 ;
  assign n50926 = \pi0211  & ~n12409 ;
  assign n50927 = ~n50396 & n50926 ;
  assign n50928 = ~n50393 & n50927 ;
  assign n50929 = \pi0214  & ~n50928 ;
  assign n50930 = ~n50925 & n50929 ;
  assign n50931 = \pi0211  & n50930 ;
  assign n50932 = ~n50586 & n50930 ;
  assign n50933 = ~n50919 & n50932 ;
  assign n50934 = ~n50931 & ~n50933 ;
  assign n50935 = n50923 & n50934 ;
  assign n50936 = \pi0219  & ~n50877 ;
  assign n50937 = ~n50875 & n50936 ;
  assign n50938 = \pi0219  & ~n12409 ;
  assign n50939 = ~n50396 & n50938 ;
  assign n50940 = ~n50393 & n50939 ;
  assign n50941 = \pi0212  & n9948 ;
  assign n50942 = ~n50940 & n50941 ;
  assign n50943 = ~n50937 & n50942 ;
  assign n50944 = ~n50935 & n50943 ;
  assign n50945 = \pi0211  & \pi1153  ;
  assign n50946 = ~n50627 & ~n50945 ;
  assign n50947 = ~n12255 & n50946 ;
  assign n50948 = ~\pi0219  & ~n50570 ;
  assign n50949 = ~n50626 & n50948 ;
  assign n50950 = ~n50947 & n50949 ;
  assign n50951 = ~n27408 & n50950 ;
  assign n50952 = ~\pi1152  & ~n50951 ;
  assign n50953 = ~n50919 & n50920 ;
  assign n50954 = \pi0214  & ~\pi0219  ;
  assign n50955 = n50907 & n50954 ;
  assign n50956 = ~n50953 & n50955 ;
  assign n50957 = n9948 & ~n50940 ;
  assign n50958 = ~n50937 & n50957 ;
  assign n50959 = ~\pi0219  & ~n50884 ;
  assign n50960 = n50958 & ~n50959 ;
  assign n50961 = ~n50956 & n50960 ;
  assign n50962 = n50952 & ~n50961 ;
  assign n50963 = ~n50944 & n50962 ;
  assign n50964 = ~\pi0213  & ~n50963 ;
  assign n50965 = \pi0212  & \pi1153  ;
  assign n50966 = ~n50442 & n50965 ;
  assign n50967 = ~\pi0211  & \pi0214  ;
  assign n50968 = \pi0212  & ~n50967 ;
  assign n50969 = ~n50628 & n50968 ;
  assign n50970 = ~n50966 & ~n50969 ;
  assign n50971 = n50556 & ~n50946 ;
  assign n50972 = ~\pi0219  & ~n50971 ;
  assign n50973 = n50970 & n50972 ;
  assign n50974 = n50677 & ~n50973 ;
  assign n50975 = \pi1152  & ~n50974 ;
  assign n50976 = ~n50956 & ~n50959 ;
  assign n50977 = ~\pi0211  & n50586 ;
  assign n50978 = \pi0214  & ~n50977 ;
  assign n50979 = \pi0212  & n50978 ;
  assign n50980 = ~n50919 & n50979 ;
  assign n50981 = n50600 & ~n50907 ;
  assign n50982 = n50600 & n50920 ;
  assign n50983 = ~n50919 & n50982 ;
  assign n50984 = ~n50981 & ~n50983 ;
  assign n50985 = ~n50980 & n50984 ;
  assign n50986 = ~n50976 & n50985 ;
  assign n50987 = n9948 & ~n50899 ;
  assign n50988 = n9948 & n50571 ;
  assign n50989 = ~n50919 & n50988 ;
  assign n50990 = ~n50987 & ~n50989 ;
  assign n50991 = ~n50986 & ~n50990 ;
  assign n50992 = n50975 & ~n50991 ;
  assign n50993 = n50964 & ~n50992 ;
  assign n50994 = ~n50912 & ~n50993 ;
  assign n50995 = \pi0209  & ~n50994 ;
  assign n50996 = ~\pi0230  & \pi0234  ;
  assign n50997 = ~\pi0057  & \pi1152  ;
  assign n50998 = n6848 & n50997 ;
  assign n50999 = ~\pi1153  & ~n15351 ;
  assign n51000 = ~n50513 & ~n50999 ;
  assign n51001 = ~\pi0199  & ~\pi1153  ;
  assign n51002 = ~\pi0299  & ~n51001 ;
  assign n51003 = n50371 & n51002 ;
  assign n51004 = ~n12409 & ~n51003 ;
  assign n51005 = ~n51000 & n51004 ;
  assign n51006 = ~n50571 & ~n50876 ;
  assign n51007 = ~\pi1153  & n12691 ;
  assign n51008 = n50824 & ~n51007 ;
  assign n51009 = n12409 & ~n51008 ;
  assign n51010 = n51006 & ~n51009 ;
  assign n51011 = ~n51005 & n51010 ;
  assign n51012 = ~n50571 & ~n51011 ;
  assign n51013 = ~\pi0200  & ~\pi1153  ;
  assign n51014 = ~\pi0199  & ~n51013 ;
  assign n51015 = n50384 & ~n51014 ;
  assign n51016 = \pi0207  & ~n50412 ;
  assign n51017 = \pi0208  & n51016 ;
  assign n51018 = ~n51015 & n51017 ;
  assign n51019 = \pi1154  & ~n50390 ;
  assign n51020 = ~n51003 & ~n51019 ;
  assign n51021 = ~n51000 & n51020 ;
  assign n51022 = n50381 & ~n51021 ;
  assign n51023 = ~n51018 & ~n51022 ;
  assign n51024 = ~n50416 & ~n51003 ;
  assign n51025 = ~n51000 & n51024 ;
  assign n51026 = ~\pi0208  & ~n50851 ;
  assign n51027 = ~n51025 & n51026 ;
  assign n51028 = ~n51011 & ~n51027 ;
  assign n51029 = n51023 & n51028 ;
  assign n51030 = ~n51012 & ~n51029 ;
  assign n51031 = \pi0219  & n51030 ;
  assign n51032 = n50998 & n51031 ;
  assign n51033 = ~\pi0299  & \pi1153  ;
  assign n51034 = n13645 & n51033 ;
  assign n51035 = ~\pi1154  & ~n51034 ;
  assign n51036 = ~\pi0199  & \pi1153  ;
  assign n51037 = \pi1154  & n44035 ;
  assign n51038 = ~n51036 & n51037 ;
  assign n51039 = ~n51035 & ~n51038 ;
  assign n51040 = ~n50383 & n50410 ;
  assign n51041 = ~n51039 & n51040 ;
  assign n51042 = ~n50383 & n50544 ;
  assign n51043 = ~n51014 & n51042 ;
  assign n51044 = \pi0208  & ~n51043 ;
  assign n51045 = ~n51041 & n51044 ;
  assign n51046 = n50384 & ~n51039 ;
  assign n51047 = n50437 & ~n51046 ;
  assign n51048 = ~n51045 & ~n51047 ;
  assign n51049 = ~\pi1154  & n12691 ;
  assign n51050 = n50410 & n51049 ;
  assign n51051 = \pi0299  & ~\pi1155  ;
  assign n51052 = \pi0211  & ~n51051 ;
  assign n51053 = ~n51050 & n51052 ;
  assign n51054 = ~n51048 & n51053 ;
  assign n51055 = ~n50483 & ~n51003 ;
  assign n51056 = ~n51000 & n51055 ;
  assign n51057 = ~\pi0207  & ~n51056 ;
  assign n51058 = \pi0299  & ~\pi1156  ;
  assign n51059 = \pi0207  & ~n51058 ;
  assign n51060 = ~n51015 & n51059 ;
  assign n51061 = \pi0208  & ~n51060 ;
  assign n51062 = ~n51057 & n51061 ;
  assign n51063 = ~\pi0208  & ~n50483 ;
  assign n51064 = ~n51003 & n51063 ;
  assign n51065 = ~n51000 & n51064 ;
  assign n51066 = ~n50483 & n50876 ;
  assign n51067 = ~\pi0211  & ~n51066 ;
  assign n51068 = ~n51065 & n51067 ;
  assign n51069 = ~n51062 & n51068 ;
  assign n51070 = ~n51054 & ~n51069 ;
  assign n51071 = n50679 & n51070 ;
  assign n51072 = ~n50876 & ~n51009 ;
  assign n51073 = ~n51005 & n51072 ;
  assign n51074 = n50570 & ~n51073 ;
  assign n51075 = ~\pi0219  & ~n51074 ;
  assign n51076 = ~n51071 & n51075 ;
  assign n51077 = n51023 & ~n51027 ;
  assign n51078 = \pi0211  & ~n51077 ;
  assign n51079 = ~\pi0211  & ~n51051 ;
  assign n51080 = ~n51050 & n51079 ;
  assign n51081 = ~n51048 & n51080 ;
  assign n51082 = n12255 & ~n51081 ;
  assign n51083 = ~n51078 & n51082 ;
  assign n51084 = n50998 & ~n51083 ;
  assign n51085 = n51076 & n51084 ;
  assign n51086 = ~n51032 & ~n51085 ;
  assign n51087 = ~\pi0057  & ~\pi1152  ;
  assign n51088 = n6848 & n51087 ;
  assign n51089 = \pi0207  & n51034 ;
  assign n51090 = ~\pi1153  & n44035 ;
  assign n51091 = ~n13558 & n50377 ;
  assign n51092 = ~n51090 & n51091 ;
  assign n51093 = ~n51089 & ~n51092 ;
  assign n51094 = ~n50848 & n51093 ;
  assign n51095 = ~\pi0208  & ~n51094 ;
  assign n51096 = \pi1154  & ~n13558 ;
  assign n51097 = ~n51090 & n51096 ;
  assign n51098 = ~\pi0207  & ~n51034 ;
  assign n51099 = ~n51097 & n51098 ;
  assign n51100 = ~\pi0299  & ~\pi1153  ;
  assign n51101 = ~n50412 & ~n51100 ;
  assign n51102 = ~n50390 & n51101 ;
  assign n51103 = \pi0207  & ~n51102 ;
  assign n51104 = \pi0208  & ~n51103 ;
  assign n51105 = ~n51099 & n51104 ;
  assign n51106 = ~\pi0211  & ~n51105 ;
  assign n51107 = ~n51095 & n51106 ;
  assign n51108 = \pi0219  & ~n50570 ;
  assign n51109 = \pi0200  & ~\pi1153  ;
  assign n51110 = n13550 & ~n51109 ;
  assign n51111 = \pi1154  & ~n51110 ;
  assign n51112 = ~n51035 & ~n51111 ;
  assign n51113 = n50877 & n51112 ;
  assign n51114 = n12691 & n50544 ;
  assign n51115 = \pi0208  & \pi1153  ;
  assign n51116 = n51114 & n51115 ;
  assign n51117 = \pi0211  & ~n51116 ;
  assign n51118 = ~n51113 & n51117 ;
  assign n51119 = n51108 & ~n51118 ;
  assign n51120 = ~n51107 & n51119 ;
  assign n51121 = n50570 & n50877 ;
  assign n51122 = n51112 & n51121 ;
  assign n51123 = n50570 & n51115 ;
  assign n51124 = n51114 & n51123 ;
  assign n51125 = ~n51122 & ~n51124 ;
  assign n51126 = ~n51120 & n51125 ;
  assign n51127 = n51088 & ~n51126 ;
  assign n51128 = ~\pi0211  & ~n50483 ;
  assign n51129 = ~n51116 & n51128 ;
  assign n51130 = ~n51113 & n51129 ;
  assign n51131 = n50679 & ~n51130 ;
  assign n51132 = ~n50772 & ~n51131 ;
  assign n51133 = n13645 & n50460 ;
  assign n51134 = ~n50412 & ~n51133 ;
  assign n51135 = ~n51051 & ~n51134 ;
  assign n51136 = ~n13558 & ~n51090 ;
  assign n51137 = \pi1154  & ~n50433 ;
  assign n51138 = n51136 & n51137 ;
  assign n51139 = ~n51135 & ~n51138 ;
  assign n51140 = \pi0207  & n51139 ;
  assign n51141 = n50437 & ~n51140 ;
  assign n51142 = ~\pi0207  & n51139 ;
  assign n51143 = ~n51051 & ~n51100 ;
  assign n51144 = ~n50390 & n51143 ;
  assign n51145 = \pi0207  & ~n51144 ;
  assign n51146 = \pi0208  & ~n51145 ;
  assign n51147 = ~n51142 & n51146 ;
  assign n51148 = ~n51141 & ~n51147 ;
  assign n51149 = ~n51132 & ~n51148 ;
  assign n51150 = n50805 & ~n51130 ;
  assign n51151 = ~n51095 & ~n51105 ;
  assign n51152 = n12256 & ~n51151 ;
  assign n51153 = ~n51150 & ~n51152 ;
  assign n51154 = ~n51149 & n51153 ;
  assign n51155 = ~\pi0219  & n51088 ;
  assign n51156 = ~n51154 & n51155 ;
  assign n51157 = ~n51127 & ~n51156 ;
  assign n51158 = \pi0213  & n51157 ;
  assign n51159 = n51086 & n51158 ;
  assign n51160 = ~\pi0209  & ~n51159 ;
  assign n51161 = n50556 & ~n50614 ;
  assign n51162 = ~\pi0219  & ~n51161 ;
  assign n51163 = n50616 & n51162 ;
  assign n51164 = \pi0219  & ~n50627 ;
  assign n51165 = \pi0213  & ~n51164 ;
  assign n51166 = n50677 & n51165 ;
  assign n51167 = ~n51163 & n51166 ;
  assign n51168 = ~n51160 & ~n51167 ;
  assign n51169 = ~n12256 & n50948 ;
  assign n51170 = ~n51116 & ~n51169 ;
  assign n51171 = ~n51113 & n51170 ;
  assign n51172 = n27408 & ~n51171 ;
  assign n51173 = n50952 & ~n51172 ;
  assign n51174 = ~\pi0219  & ~\pi1152  ;
  assign n51175 = ~n50951 & n51174 ;
  assign n51176 = ~\pi1153  & ~n44032 ;
  assign n51177 = n51096 & ~n51176 ;
  assign n51178 = ~\pi0299  & ~n13645 ;
  assign n51179 = n50460 & ~n51178 ;
  assign n51180 = ~n51177 & ~n51179 ;
  assign n51181 = ~\pi0207  & ~n51180 ;
  assign n51182 = \pi0207  & \pi1153  ;
  assign n51183 = ~n50390 & n51182 ;
  assign n51184 = \pi0208  & ~n51183 ;
  assign n51185 = ~n51181 & n51184 ;
  assign n51186 = \pi0207  & ~n51180 ;
  assign n51187 = \pi0299  & \pi1153  ;
  assign n51188 = ~\pi0207  & n51187 ;
  assign n51189 = ~\pi0208  & ~n51188 ;
  assign n51190 = ~n51186 & n51189 ;
  assign n51191 = ~n51185 & ~n51190 ;
  assign n51192 = ~n50774 & ~n51191 ;
  assign n51193 = n50679 & ~n51095 ;
  assign n51194 = n51106 & n51193 ;
  assign n51195 = ~n51192 & ~n51194 ;
  assign n51196 = n51175 & ~n51195 ;
  assign n51197 = ~n51173 & ~n51196 ;
  assign n51198 = \pi0211  & ~n50876 ;
  assign n51199 = ~n50570 & n51198 ;
  assign n51200 = ~n51009 & n51199 ;
  assign n51201 = ~n51005 & n51200 ;
  assign n51202 = n50411 & ~n51046 ;
  assign n51203 = ~n51045 & ~n51202 ;
  assign n51204 = n50571 & ~n51203 ;
  assign n51205 = ~n51201 & ~n51204 ;
  assign n51206 = \pi0219  & ~n51073 ;
  assign n51207 = ~n51108 & ~n51206 ;
  assign n51208 = n51205 & ~n51207 ;
  assign n51209 = n9948 & ~n51208 ;
  assign n51210 = n50975 & ~n51209 ;
  assign n51211 = ~\pi0211  & ~n51077 ;
  assign n51212 = ~\pi0207  & \pi1154  ;
  assign n51213 = ~n13558 & n51212 ;
  assign n51214 = ~n51176 & n51213 ;
  assign n51215 = ~\pi1153  & ~n13558 ;
  assign n51216 = ~\pi0207  & ~n51215 ;
  assign n51217 = ~n50432 & n51216 ;
  assign n51218 = ~n51214 & ~n51217 ;
  assign n51219 = ~\pi1153  & ~n50390 ;
  assign n51220 = \pi0207  & ~n50840 ;
  assign n51221 = ~n51219 & n51220 ;
  assign n51222 = n51218 & ~n51221 ;
  assign n51223 = n50845 & ~n51222 ;
  assign n51224 = \pi0207  & ~n51215 ;
  assign n51225 = ~n50432 & n51224 ;
  assign n51226 = n51091 & ~n51176 ;
  assign n51227 = ~n51188 & ~n51226 ;
  assign n51228 = ~n51225 & n51227 ;
  assign n51229 = n50852 & ~n51228 ;
  assign n51230 = ~\pi0214  & ~n51229 ;
  assign n51231 = ~n51223 & n51230 ;
  assign n51232 = ~n51211 & n51231 ;
  assign n51233 = \pi0211  & ~n51203 ;
  assign n51234 = n50904 & ~n51228 ;
  assign n51235 = \pi0214  & ~n50901 ;
  assign n51236 = \pi0214  & ~n51221 ;
  assign n51237 = n51218 & n51236 ;
  assign n51238 = ~n51235 & ~n51237 ;
  assign n51239 = ~n51234 & ~n51238 ;
  assign n51240 = ~n51233 & n51239 ;
  assign n51241 = \pi0212  & ~n51240 ;
  assign n51242 = ~n51232 & n51241 ;
  assign n51243 = ~\pi0214  & ~n51073 ;
  assign n51244 = ~\pi0212  & ~n51243 ;
  assign n51245 = \pi0214  & ~n51229 ;
  assign n51246 = ~n51223 & n51245 ;
  assign n51247 = ~n51211 & n51246 ;
  assign n51248 = n51244 & ~n51247 ;
  assign n51249 = ~n51242 & ~n51248 ;
  assign n51250 = ~\pi0219  & n50975 ;
  assign n51251 = n51249 & n51250 ;
  assign n51252 = ~n51210 & ~n51251 ;
  assign n51253 = n51197 & n51252 ;
  assign n51254 = ~\pi0213  & ~n51253 ;
  assign n51255 = ~n51168 & ~n51254 ;
  assign n51256 = ~n50996 & ~n51255 ;
  assign n51257 = ~n50995 & n51256 ;
  assign n51258 = ~n50822 & ~n51257 ;
  assign n51259 = ~\pi0230  & ~\pi0235  ;
  assign n51260 = ~n50480 & ~n50592 ;
  assign n51261 = ~\pi1157  & ~n50421 ;
  assign n51262 = ~n51260 & n51261 ;
  assign n51263 = ~\pi1156  & n50388 ;
  assign n51264 = n50496 & ~n51263 ;
  assign n51265 = n12409 & ~n51264 ;
  assign n51266 = n50381 & n50591 ;
  assign n51267 = ~n51265 & ~n51266 ;
  assign n51268 = ~\pi1157  & ~n51267 ;
  assign n51269 = \pi0208  & \pi1157  ;
  assign n51270 = \pi0207  & n51269 ;
  assign n51271 = ~n51264 & n51270 ;
  assign n51272 = \pi1156  & ~n50403 ;
  assign n51273 = ~n50488 & ~n51272 ;
  assign n51274 = ~\pi0207  & n51269 ;
  assign n51275 = ~n51273 & n51274 ;
  assign n51276 = ~n51271 & ~n51275 ;
  assign n51277 = n50492 & n51276 ;
  assign n51278 = ~n51268 & n51277 ;
  assign n51279 = ~n51262 & n51278 ;
  assign n51280 = \pi0211  & ~n51279 ;
  assign n51281 = ~n50409 & n50411 ;
  assign n51282 = n50617 & n51281 ;
  assign n51283 = ~n50382 & n50544 ;
  assign n51284 = n50496 & n51283 ;
  assign n51285 = \pi0208  & ~n51284 ;
  assign n51286 = ~\pi0207  & ~n50407 ;
  assign n51287 = ~n50404 & n51286 ;
  assign n51288 = n50617 & ~n51287 ;
  assign n51289 = n51285 & n51288 ;
  assign n51290 = ~n51282 & ~n51289 ;
  assign n51291 = ~\pi0208  & ~n50530 ;
  assign n51292 = ~\pi0207  & ~n50424 ;
  assign n51293 = \pi0207  & ~n51263 ;
  assign n51294 = n50525 & n51293 ;
  assign n51295 = ~n51292 & ~n51294 ;
  assign n51296 = ~n51291 & n51295 ;
  assign n51297 = ~\pi0211  & ~\pi1157  ;
  assign n51298 = n51296 & n51297 ;
  assign n51299 = n51290 & ~n51298 ;
  assign n51300 = n50679 & n51299 ;
  assign n51301 = ~n51280 & n51300 ;
  assign n51302 = n50772 & ~n51262 ;
  assign n51303 = n51278 & n51302 ;
  assign n51304 = ~\pi1157  & ~n50433 ;
  assign n51305 = ~n50432 & n51304 ;
  assign n51306 = n50440 & n51305 ;
  assign n51307 = \pi1155  & ~n51178 ;
  assign n51308 = ~n50396 & ~n51307 ;
  assign n51309 = \pi0207  & ~n51308 ;
  assign n51310 = ~\pi0207  & ~n50401 ;
  assign n51311 = ~\pi0207  & \pi1155  ;
  assign n51312 = n50383 & n51311 ;
  assign n51313 = ~n51310 & ~n51312 ;
  assign n51314 = n50434 & ~n51313 ;
  assign n51315 = ~n51309 & ~n51314 ;
  assign n51316 = \pi0208  & ~\pi1157  ;
  assign n51317 = ~n51315 & n51316 ;
  assign n51318 = ~n51306 & ~n51317 ;
  assign n51319 = ~\pi0207  & n50395 ;
  assign n51320 = ~\pi0207  & ~n44035 ;
  assign n51321 = ~n50448 & n51320 ;
  assign n51322 = ~n51319 & ~n51321 ;
  assign n51323 = ~n51309 & n51322 ;
  assign n51324 = n51269 & ~n51323 ;
  assign n51325 = n12256 & ~n50579 ;
  assign n51326 = ~n51324 & n51325 ;
  assign n51327 = n51318 & n51326 ;
  assign n51328 = ~n51303 & ~n51327 ;
  assign n51329 = ~\pi0207  & n50489 ;
  assign n51330 = ~n51294 & ~n51329 ;
  assign n51331 = ~n50560 & n51330 ;
  assign n51332 = \pi1157  & n50570 ;
  assign n51333 = ~n51331 & n51332 ;
  assign n51334 = ~\pi1157  & n50570 ;
  assign n51335 = ~n51296 & n51334 ;
  assign n51336 = ~n51333 & ~n51335 ;
  assign n51337 = n51328 & n51336 ;
  assign n51338 = ~n51301 & n51337 ;
  assign n51339 = ~\pi0219  & ~n51338 ;
  assign n51340 = ~\pi1157  & ~n50679 ;
  assign n51341 = n51296 & n51340 ;
  assign n51342 = \pi1157  & ~n50679 ;
  assign n51343 = n51331 & n51342 ;
  assign n51344 = \pi0219  & ~n51343 ;
  assign n51345 = ~n51341 & n51344 ;
  assign n51346 = \pi0209  & ~n51345 ;
  assign n51347 = \pi0211  & ~\pi1157  ;
  assign n51348 = ~n51296 & n51347 ;
  assign n51349 = \pi0211  & \pi1157  ;
  assign n51350 = ~n51331 & n51349 ;
  assign n51351 = n50679 & ~n51350 ;
  assign n51352 = ~n51348 & n51351 ;
  assign n51353 = ~\pi0211  & ~n50579 ;
  assign n51354 = ~n51324 & n51353 ;
  assign n51355 = n51318 & n51354 ;
  assign n51356 = \pi0209  & ~n51355 ;
  assign n51357 = n51352 & n51356 ;
  assign n51358 = ~n51346 & ~n51357 ;
  assign n51359 = n27408 & ~n51358 ;
  assign n51360 = ~n51339 & n51359 ;
  assign n51361 = \pi1154  & n12409 ;
  assign n51362 = ~n51110 & n51361 ;
  assign n51363 = ~\pi1154  & n12409 ;
  assign n51364 = ~n51034 & n51363 ;
  assign n51365 = ~n51362 & ~n51364 ;
  assign n51366 = ~n50876 & n51365 ;
  assign n51367 = n51128 & ~n51366 ;
  assign n51368 = ~n50509 & ~n50514 ;
  assign n51369 = ~n12409 & n51128 ;
  assign n51370 = ~n51368 & n51369 ;
  assign n51371 = ~n51367 & ~n51370 ;
  assign n51372 = n12255 & ~n51371 ;
  assign n51373 = ~\pi0207  & n50466 ;
  assign n51374 = ~n50457 & n51373 ;
  assign n51375 = \pi0208  & ~n51140 ;
  assign n51376 = ~n51374 & n51375 ;
  assign n51377 = n50437 & ~n50466 ;
  assign n51378 = \pi1154  & n50437 ;
  assign n51379 = ~n50456 & n51378 ;
  assign n51380 = ~n51377 & ~n51379 ;
  assign n51381 = \pi0211  & n51380 ;
  assign n51382 = n12255 & n51381 ;
  assign n51383 = ~n51376 & n51382 ;
  assign n51384 = ~n51372 & ~n51383 ;
  assign n51385 = \pi0299  & n50618 ;
  assign n51386 = ~n51366 & ~n51385 ;
  assign n51387 = ~n12409 & ~n51385 ;
  assign n51388 = ~n51368 & n51387 ;
  assign n51389 = ~n51386 & ~n51388 ;
  assign n51390 = ~n12255 & ~n50617 ;
  assign n51391 = ~n51389 & n51390 ;
  assign n51392 = n50411 & ~n50547 ;
  assign n51393 = ~n50570 & n50617 ;
  assign n51394 = ~n51392 & n51393 ;
  assign n51395 = n50410 & ~n50507 ;
  assign n51396 = ~n50543 & n51395 ;
  assign n51397 = ~n50504 & n51396 ;
  assign n51398 = n51016 & ~n51133 ;
  assign n51399 = ~n51097 & n51398 ;
  assign n51400 = \pi0208  & ~n51399 ;
  assign n51401 = ~n51397 & n51400 ;
  assign n51402 = ~n12255 & ~n51401 ;
  assign n51403 = n51394 & n51402 ;
  assign n51404 = n50570 & ~n51366 ;
  assign n51405 = ~n12409 & n50570 ;
  assign n51406 = ~n51368 & n51405 ;
  assign n51407 = ~n51404 & ~n51406 ;
  assign n51408 = ~n51403 & n51407 ;
  assign n51409 = ~n51391 & n51408 ;
  assign n51410 = n51384 & n51409 ;
  assign n51411 = ~\pi0219  & ~n51410 ;
  assign n51412 = ~n12409 & ~n51368 ;
  assign n51413 = ~n50679 & n51366 ;
  assign n51414 = ~n51412 & n51413 ;
  assign n51415 = \pi0219  & ~n51414 ;
  assign n51416 = ~\pi0209  & ~n51415 ;
  assign n51417 = \pi0211  & ~n51366 ;
  assign n51418 = n50926 & ~n51368 ;
  assign n51419 = ~n51417 & ~n51418 ;
  assign n51420 = n50679 & n51419 ;
  assign n51421 = ~\pi0211  & n51380 ;
  assign n51422 = ~\pi0209  & ~n51421 ;
  assign n51423 = ~\pi0209  & ~n51374 ;
  assign n51424 = n51375 & n51423 ;
  assign n51425 = ~n51422 & ~n51424 ;
  assign n51426 = n51420 & ~n51425 ;
  assign n51427 = ~n51416 & ~n51426 ;
  assign n51428 = n9948 & ~n51427 ;
  assign n51429 = ~n51411 & n51428 ;
  assign n51430 = n12255 & ~n50614 ;
  assign n51431 = n50600 & ~n50619 ;
  assign n51432 = ~n51430 & ~n51431 ;
  assign n51433 = n50621 & n51432 ;
  assign n51434 = n50608 & n50679 ;
  assign n51435 = \pi0219  & ~n51434 ;
  assign n51436 = ~n9948 & ~n51435 ;
  assign n51437 = ~n51433 & n51436 ;
  assign n51438 = \pi0213  & ~n51437 ;
  assign n51439 = ~n51429 & n51438 ;
  assign n51440 = ~n51360 & n51439 ;
  assign n51441 = ~\pi0299  & ~\pi1157  ;
  assign n51442 = n50482 & n51441 ;
  assign n51443 = n51267 & n51442 ;
  assign n51444 = n51285 & ~n51287 ;
  assign n51445 = \pi1157  & ~n51281 ;
  assign n51446 = ~n51444 & n51445 ;
  assign n51447 = n50920 & ~n51446 ;
  assign n51448 = ~n51443 & n51447 ;
  assign n51449 = \pi0207  & \pi0208  ;
  assign n51450 = ~n50388 & ~n50416 ;
  assign n51451 = ~n50396 & n51450 ;
  assign n51452 = n51449 & ~n51451 ;
  assign n51453 = \pi1154  & ~n50477 ;
  assign n51454 = ~n50423 & ~n51453 ;
  assign n51455 = \pi0208  & ~n51313 ;
  assign n51456 = ~n51454 & n51455 ;
  assign n51457 = ~n51452 & ~n51456 ;
  assign n51458 = n50426 & n51457 ;
  assign n51459 = n51297 & ~n51458 ;
  assign n51460 = n50413 & n51281 ;
  assign n51461 = n50413 & ~n51287 ;
  assign n51462 = n51285 & n51461 ;
  assign n51463 = ~n51460 & ~n51462 ;
  assign n51464 = ~\pi0211  & ~n51463 ;
  assign n51465 = n12255 & ~n51464 ;
  assign n51466 = ~n51459 & n51465 ;
  assign n51467 = ~n51448 & n51466 ;
  assign n51468 = ~\pi0219  & n51467 ;
  assign n51469 = ~\pi1157  & ~n51458 ;
  assign n51470 = \pi0211  & n51463 ;
  assign n51471 = ~n51469 & n51470 ;
  assign n51472 = n51336 & ~n51355 ;
  assign n51473 = ~n51471 & n51472 ;
  assign n51474 = ~n50679 & n51336 ;
  assign n51475 = ~\pi0219  & ~n51474 ;
  assign n51476 = ~n51473 & n51475 ;
  assign n51477 = ~n51468 & ~n51476 ;
  assign n51478 = \pi0209  & ~n51348 ;
  assign n51479 = n51351 & n51478 ;
  assign n51480 = ~n50586 & ~n51446 ;
  assign n51481 = ~n51443 & n51480 ;
  assign n51482 = ~\pi0211  & ~n51481 ;
  assign n51483 = n51479 & ~n51482 ;
  assign n51484 = ~n51346 & ~n51483 ;
  assign n51485 = n27408 & ~n51484 ;
  assign n51486 = n51477 & n51485 ;
  assign n51487 = ~\pi0208  & n51188 ;
  assign n51488 = n50418 & ~n50584 ;
  assign n51489 = ~n51487 & ~n51488 ;
  assign n51490 = n50381 & ~n50584 ;
  assign n51491 = ~n51180 & n51449 ;
  assign n51492 = ~\pi0211  & ~n51491 ;
  assign n51493 = ~n51490 & n51492 ;
  assign n51494 = n51489 & n51493 ;
  assign n51495 = ~\pi0209  & ~n51494 ;
  assign n51496 = n51420 & n51495 ;
  assign n51497 = ~n51416 & ~n51496 ;
  assign n51498 = \pi0219  & n9948 ;
  assign n51499 = n50679 & n51421 ;
  assign n51500 = ~n51376 & n51499 ;
  assign n51501 = ~n50376 & n51212 ;
  assign n51502 = ~\pi0207  & ~\pi1154  ;
  assign n51503 = ~n50365 & n51502 ;
  assign n51504 = n50364 & n51503 ;
  assign n51505 = n51093 & ~n51504 ;
  assign n51506 = ~n51501 & n51505 ;
  assign n51507 = \pi0208  & ~n51506 ;
  assign n51508 = \pi0208  & n50772 ;
  assign n51509 = n50679 & n50845 ;
  assign n51510 = ~n51508 & ~n51509 ;
  assign n51511 = ~n50376 & n50377 ;
  assign n51512 = ~n50368 & ~n50848 ;
  assign n51513 = ~n50774 & n51512 ;
  assign n51514 = ~n51511 & n51513 ;
  assign n51515 = n51510 & ~n51514 ;
  assign n51516 = ~n51507 & ~n51515 ;
  assign n51517 = ~n51500 & ~n51516 ;
  assign n51518 = n12256 & ~n51491 ;
  assign n51519 = ~n51490 & n51518 ;
  assign n51520 = n51489 & n51519 ;
  assign n51521 = n51407 & ~n51520 ;
  assign n51522 = n9948 & n51521 ;
  assign n51523 = n51517 & n51522 ;
  assign n51524 = ~n51498 & ~n51523 ;
  assign n51525 = ~n51497 & ~n51524 ;
  assign n51526 = \pi0219  & ~n50625 ;
  assign n51527 = ~n9948 & ~n51526 ;
  assign n51528 = ~\pi0219  & n12255 ;
  assign n51529 = ~n50946 & n51528 ;
  assign n51530 = ~n50610 & n50679 ;
  assign n51531 = \pi0219  & n50679 ;
  assign n51532 = ~n51530 & ~n51531 ;
  assign n51533 = ~n51529 & n51532 ;
  assign n51534 = n51527 & ~n51533 ;
  assign n51535 = ~\pi0213  & ~n51534 ;
  assign n51536 = ~n51525 & n51535 ;
  assign n51537 = ~n51486 & n51536 ;
  assign n51538 = ~n51440 & ~n51537 ;
  assign n51539 = \pi0230  & ~n51538 ;
  assign n51540 = ~n51259 & ~n51539 ;
  assign n51541 = \pi0075  & ~\pi0092  ;
  assign n51542 = ~n8416 & n51541 ;
  assign n51543 = ~\pi0054  & ~n8420 ;
  assign n51544 = ~n6837 & n51543 ;
  assign n51545 = ~n51542 & n51544 ;
  assign n51546 = n1292 & ~n50354 ;
  assign n51547 = ~n51545 & n51546 ;
  assign n51548 = ~\pi0100  & n6629 ;
  assign n51549 = n1638 & n51548 ;
  assign n51550 = ~n16448 & ~n51549 ;
  assign n51551 = n50009 & ~n51550 ;
  assign n51552 = n1640 & ~n51550 ;
  assign n51553 = ~n50033 & n51552 ;
  assign n51554 = ~n51551 & ~n51553 ;
  assign n51555 = n2364 & n50342 ;
  assign n51556 = n51546 & n51555 ;
  assign n51557 = n51554 & n51556 ;
  assign n51558 = ~n51547 & ~n51557 ;
  assign n51559 = \pi0056  & ~\pi0062  ;
  assign n51560 = ~n6833 & n51559 ;
  assign n51561 = n2467 & ~n51560 ;
  assign n51562 = ~n16284 & n51561 ;
  assign n51563 = n51558 & n51562 ;
  assign n51564 = ~\pi0230  & \pi0237  ;
  assign n51565 = \pi0207  & n50752 ;
  assign n51566 = \pi0207  & n50743 ;
  assign n51567 = ~n50739 & n51566 ;
  assign n51568 = ~n51565 & ~n51567 ;
  assign n51569 = ~\pi0207  & ~n50736 ;
  assign n51570 = \pi0208  & ~n51569 ;
  assign n51571 = ~n50438 & n51178 ;
  assign n51572 = ~n50439 & ~n51571 ;
  assign n51573 = ~\pi0200  & \pi1157  ;
  assign n51574 = ~\pi0199  & n51573 ;
  assign n51575 = \pi0208  & ~n51574 ;
  assign n51576 = ~n51572 & n51575 ;
  assign n51577 = ~n51570 & ~n51576 ;
  assign n51578 = n51568 & ~n51577 ;
  assign n51579 = ~\pi0208  & ~n50740 ;
  assign n51580 = \pi0211  & ~n51579 ;
  assign n51581 = ~\pi0200  & ~\pi1158  ;
  assign n51582 = ~\pi0199  & ~n51581 ;
  assign n51583 = \pi1156  & ~n50840 ;
  assign n51584 = ~n51582 & ~n51583 ;
  assign n51585 = ~\pi0299  & n50371 ;
  assign n51586 = \pi0199  & ~\pi1158  ;
  assign n51587 = ~n51581 & ~n51586 ;
  assign n51588 = ~n51585 & ~n51587 ;
  assign n51589 = ~n51584 & ~n51588 ;
  assign n51590 = n50544 & n51589 ;
  assign n51591 = ~\pi0299  & \pi1158  ;
  assign n51592 = n12691 & n51591 ;
  assign n51593 = \pi0199  & \pi1156  ;
  assign n51594 = \pi1156  & \pi1158  ;
  assign n51595 = ~n51593 & ~n51594 ;
  assign n51596 = ~n51592 & n51595 ;
  assign n51597 = ~\pi0200  & \pi0207  ;
  assign n51598 = ~\pi0208  & n51597 ;
  assign n51599 = ~n51596 & n51598 ;
  assign n51600 = ~n50452 & ~n51599 ;
  assign n51601 = \pi0211  & ~n51600 ;
  assign n51602 = n51590 & n51601 ;
  assign n51603 = ~n51580 & ~n51602 ;
  assign n51604 = ~n51578 & ~n51603 ;
  assign n51605 = \pi0207  & n50791 ;
  assign n51606 = \pi0207  & n50786 ;
  assign n51607 = ~n50782 & n51606 ;
  assign n51608 = ~n51605 & ~n51607 ;
  assign n51609 = ~\pi0207  & ~n50779 ;
  assign n51610 = \pi0208  & ~n51609 ;
  assign n51611 = ~n51576 & ~n51610 ;
  assign n51612 = n51608 & ~n51611 ;
  assign n51613 = ~\pi0208  & ~n50783 ;
  assign n51614 = ~\pi0211  & ~n51613 ;
  assign n51615 = ~\pi0211  & ~n51600 ;
  assign n51616 = n51590 & n51615 ;
  assign n51617 = ~n51614 & ~n51616 ;
  assign n51618 = ~n51612 & ~n51617 ;
  assign n51619 = ~n51604 & ~n51618 ;
  assign n51620 = \pi0214  & n51619 ;
  assign n51621 = ~\pi0200  & ~n51593 ;
  assign n51622 = n50824 & ~n51621 ;
  assign n51623 = \pi1157  & ~n51592 ;
  assign n51624 = ~n51622 & n51623 ;
  assign n51625 = \pi0207  & ~n51624 ;
  assign n51626 = n44032 & n51593 ;
  assign n51627 = ~\pi1157  & ~n51626 ;
  assign n51628 = ~n51592 & n51627 ;
  assign n51629 = n51625 & ~n51628 ;
  assign n51630 = \pi0299  & \pi1145  ;
  assign n51631 = ~\pi0208  & ~n51630 ;
  assign n51632 = ~\pi0211  & n51631 ;
  assign n51633 = ~n51629 & n51632 ;
  assign n51634 = ~n50747 & ~n51630 ;
  assign n51635 = ~\pi1154  & ~n51630 ;
  assign n51636 = ~n50749 & n51635 ;
  assign n51637 = \pi1156  & ~n51636 ;
  assign n51638 = ~n51634 & n51637 ;
  assign n51639 = \pi0207  & n51638 ;
  assign n51640 = \pi0299  & ~\pi1145  ;
  assign n51641 = ~n50385 & ~n51640 ;
  assign n51642 = \pi1154  & ~n51641 ;
  assign n51643 = ~n50388 & n51635 ;
  assign n51644 = ~\pi1156  & ~n51643 ;
  assign n51645 = \pi0207  & n51644 ;
  assign n51646 = ~n51642 & n51645 ;
  assign n51647 = ~n51639 & ~n51646 ;
  assign n51648 = ~\pi0207  & ~n51640 ;
  assign n51649 = \pi0208  & ~n51648 ;
  assign n51650 = ~n51576 & ~n51649 ;
  assign n51651 = ~\pi0211  & ~n51650 ;
  assign n51652 = n51647 & n51651 ;
  assign n51653 = ~n51633 & ~n51652 ;
  assign n51654 = ~\pi0214  & ~n51653 ;
  assign n51655 = n51590 & ~n51600 ;
  assign n51656 = n51613 & ~n51655 ;
  assign n51657 = ~n51612 & ~n51656 ;
  assign n51658 = n50863 & ~n51657 ;
  assign n51659 = ~n51654 & ~n51658 ;
  assign n51660 = \pi0212  & n51659 ;
  assign n51661 = ~n51620 & n51660 ;
  assign n51662 = \pi0219  & ~n50661 ;
  assign n51663 = n50677 & ~n51662 ;
  assign n51664 = \pi0213  & ~n51663 ;
  assign n51665 = ~\pi0211  & \pi1145  ;
  assign n51666 = \pi0211  & \pi1144  ;
  assign n51667 = ~n51665 & ~n51666 ;
  assign n51668 = ~n12255 & n51667 ;
  assign n51669 = n12255 & n50659 ;
  assign n51670 = ~n50570 & ~n51669 ;
  assign n51671 = ~n51668 & n51670 ;
  assign n51672 = \pi0213  & ~\pi0219  ;
  assign n51673 = ~n51671 & n51672 ;
  assign n51674 = ~n51664 & ~n51673 ;
  assign n51675 = \pi0207  & ~n50396 ;
  assign n51676 = ~n50393 & n51675 ;
  assign n51677 = ~n51292 & ~n51676 ;
  assign n51678 = n51316 & n51677 ;
  assign n51679 = n44032 & n50418 ;
  assign n51680 = ~\pi1157  & n51679 ;
  assign n51681 = ~n51596 & n51680 ;
  assign n51682 = \pi1156  & n50383 ;
  assign n51683 = ~n51582 & ~n51682 ;
  assign n51684 = ~\pi0208  & n50544 ;
  assign n51685 = \pi1157  & n51684 ;
  assign n51686 = ~n51683 & n51685 ;
  assign n51687 = ~n51681 & ~n51686 ;
  assign n51688 = ~n51678 & n51687 ;
  assign n51689 = ~n51329 & ~n51676 ;
  assign n51690 = n51269 & n51689 ;
  assign n51691 = ~\pi0214  & ~n51690 ;
  assign n51692 = n51688 & n51691 ;
  assign n51693 = ~\pi0212  & ~n51692 ;
  assign n51694 = ~\pi0219  & ~n51693 ;
  assign n51695 = n50954 & ~n51653 ;
  assign n51696 = \pi0211  & n50954 ;
  assign n51697 = ~n51657 & n51696 ;
  assign n51698 = ~n51695 & ~n51697 ;
  assign n51699 = ~n51694 & n51698 ;
  assign n51700 = ~n51674 & ~n51699 ;
  assign n51701 = ~n51661 & n51700 ;
  assign n51702 = ~n50571 & ~n51690 ;
  assign n51703 = n51688 & n51702 ;
  assign n51704 = n50571 & ~n51577 ;
  assign n51705 = n51568 & n51704 ;
  assign n51706 = n50571 & n51579 ;
  assign n51707 = ~n51655 & n51706 ;
  assign n51708 = ~n51705 & ~n51707 ;
  assign n51709 = ~n51703 & n51708 ;
  assign n51710 = \pi0219  & ~n51709 ;
  assign n51711 = n27408 & ~n51710 ;
  assign n51712 = ~n51674 & ~n51711 ;
  assign n51713 = ~\pi0209  & ~n51712 ;
  assign n51714 = ~n51701 & n51713 ;
  assign n51715 = ~\pi0230  & ~\pi0237  ;
  assign n51716 = \pi0199  & \pi1143  ;
  assign n51717 = ~\pi0200  & ~n51716 ;
  assign n51718 = ~n50644 & n51717 ;
  assign n51719 = n50641 & ~n50652 ;
  assign n51720 = ~n51718 & n51719 ;
  assign n51721 = ~\pi0199  & \pi1145  ;
  assign n51722 = n51717 & ~n51721 ;
  assign n51723 = \pi0200  & ~n50644 ;
  assign n51724 = n50877 & ~n51723 ;
  assign n51725 = ~n51722 & n51724 ;
  assign n51726 = ~n51720 & ~n51725 ;
  assign n51727 = ~\pi0299  & ~n51726 ;
  assign n51728 = n50701 & ~n51668 ;
  assign n51729 = n51670 & n51728 ;
  assign n51730 = ~n50570 & n50689 ;
  assign n51731 = n50740 & n51730 ;
  assign n51732 = ~n51729 & ~n51731 ;
  assign n51733 = ~n51727 & n51732 ;
  assign n51734 = n9948 & ~n51733 ;
  assign n51735 = ~n51674 & ~n51734 ;
  assign n51736 = ~n51715 & n51735 ;
  assign n51737 = ~\pi0211  & \pi1158  ;
  assign n51738 = ~n51349 & ~n51737 ;
  assign n51739 = n50556 & ~n51738 ;
  assign n51740 = ~\pi0219  & ~n51739 ;
  assign n51741 = n51432 & n51740 ;
  assign n51742 = n50701 & ~n51741 ;
  assign n51743 = n50483 & n50689 ;
  assign n51744 = n50556 & n51743 ;
  assign n51745 = ~\pi0214  & n50435 ;
  assign n51746 = \pi1154  & n50693 ;
  assign n51747 = ~n51745 & ~n51746 ;
  assign n51748 = n50696 & ~n51747 ;
  assign n51749 = ~n51744 & ~n51748 ;
  assign n51750 = ~n51727 & n51749 ;
  assign n51751 = ~n51742 & n51750 ;
  assign n51752 = ~\pi0057  & \pi0209  ;
  assign n51753 = n6848 & n51752 ;
  assign n51754 = ~n51751 & n51753 ;
  assign n51755 = \pi0214  & n50627 ;
  assign n51756 = \pi1155  & n50442 ;
  assign n51757 = ~n51755 & ~n51756 ;
  assign n51758 = ~n9948 & ~n51757 ;
  assign n51759 = \pi0212  & n51758 ;
  assign n51760 = ~\pi0212  & \pi1156  ;
  assign n51761 = n50967 & n51760 ;
  assign n51762 = \pi0219  & ~n51761 ;
  assign n51763 = ~n9948 & ~n51762 ;
  assign n51764 = ~\pi0213  & ~n51763 ;
  assign n51765 = ~n51759 & n51764 ;
  assign n51766 = ~\pi0213  & ~\pi0219  ;
  assign n51767 = ~n51739 & n51766 ;
  assign n51768 = n51432 & n51767 ;
  assign n51769 = \pi0209  & ~n51768 ;
  assign n51770 = ~n51765 & n51769 ;
  assign n51771 = ~n51715 & ~n51770 ;
  assign n51772 = ~n51754 & n51771 ;
  assign n51773 = ~n51736 & ~n51772 ;
  assign n51774 = ~n51714 & ~n51773 ;
  assign n51775 = \pi1158  & n50541 ;
  assign n51776 = ~\pi1158  & ~n50396 ;
  assign n51777 = ~n50393 & n51776 ;
  assign n51778 = \pi0207  & ~n51777 ;
  assign n51779 = ~n51775 & n51778 ;
  assign n51780 = \pi0299  & ~\pi1158  ;
  assign n51781 = ~\pi0207  & ~n51780 ;
  assign n51782 = n51572 & n51781 ;
  assign n51783 = \pi0208  & ~n51782 ;
  assign n51784 = ~n51779 & n51783 ;
  assign n51785 = \pi0299  & \pi1158  ;
  assign n51786 = \pi0207  & \pi1158  ;
  assign n51787 = n12691 & n51786 ;
  assign n51788 = ~n51785 & ~n51787 ;
  assign n51789 = \pi0207  & n51626 ;
  assign n51790 = n51788 & ~n51789 ;
  assign n51791 = ~\pi0208  & n51790 ;
  assign n51792 = ~\pi1157  & ~n51791 ;
  assign n51793 = ~n51784 & n51792 ;
  assign n51794 = n50490 & ~n51624 ;
  assign n51795 = n50452 & ~n51788 ;
  assign n51796 = ~\pi0211  & ~n51795 ;
  assign n51797 = ~n51794 & n51796 ;
  assign n51798 = ~n51793 & n51797 ;
  assign n51799 = \pi0214  & ~n51269 ;
  assign n51800 = ~n50404 & ~n50407 ;
  assign n51801 = n51781 & ~n51800 ;
  assign n51802 = \pi0214  & ~n51801 ;
  assign n51803 = ~n51779 & n51802 ;
  assign n51804 = ~n51799 & ~n51803 ;
  assign n51805 = n51798 & ~n51804 ;
  assign n51806 = \pi0211  & ~n51681 ;
  assign n51807 = ~n51678 & n51806 ;
  assign n51808 = ~\pi0299  & n51683 ;
  assign n51809 = n50411 & ~n51808 ;
  assign n51810 = \pi1157  & n51809 ;
  assign n51811 = \pi0208  & ~n51287 ;
  assign n51812 = \pi1157  & n51811 ;
  assign n51813 = ~n50914 & n51812 ;
  assign n51814 = ~n51810 & ~n51813 ;
  assign n51815 = \pi0214  & n51814 ;
  assign n51816 = n51807 & n51815 ;
  assign n51817 = n51693 & ~n51816 ;
  assign n51818 = ~n51805 & n51817 ;
  assign n51819 = ~\pi0212  & ~\pi0219  ;
  assign n51820 = ~n51678 & ~n51681 ;
  assign n51821 = n51814 & n51820 ;
  assign n51822 = n50442 & ~n51821 ;
  assign n51823 = ~\pi0207  & n50591 ;
  assign n51824 = \pi0208  & n50496 ;
  assign n51825 = ~n50393 & n51824 ;
  assign n51826 = ~n50381 & ~n51825 ;
  assign n51827 = ~n51823 & ~n51826 ;
  assign n51828 = n51063 & n51596 ;
  assign n51829 = n51063 & ~n51597 ;
  assign n51830 = ~\pi1157  & ~n51829 ;
  assign n51831 = ~n51828 & n51830 ;
  assign n51832 = ~n51827 & n51831 ;
  assign n51833 = n50452 & n50544 ;
  assign n51834 = ~n51683 & n51833 ;
  assign n51835 = ~n50484 & ~n51834 ;
  assign n51836 = ~\pi0207  & n51273 ;
  assign n51837 = ~n50495 & n50499 ;
  assign n51838 = ~n50393 & n51837 ;
  assign n51839 = ~n51836 & ~n51838 ;
  assign n51840 = n51269 & n51839 ;
  assign n51841 = n51835 & ~n51840 ;
  assign n51842 = ~n51832 & n51841 ;
  assign n51843 = n50443 & ~n51842 ;
  assign n51844 = ~n51822 & ~n51843 ;
  assign n51845 = n51269 & ~n51322 ;
  assign n51846 = ~n50833 & n51270 ;
  assign n51847 = ~n51845 & ~n51846 ;
  assign n51848 = n50435 & n50452 ;
  assign n51849 = n51589 & n51833 ;
  assign n51850 = ~n51848 & ~n51849 ;
  assign n51851 = n51847 & n51850 ;
  assign n51852 = n50430 & ~n51851 ;
  assign n51853 = n12409 & ~n50833 ;
  assign n51854 = n50434 & n51455 ;
  assign n51855 = ~n51596 & n51679 ;
  assign n51856 = ~\pi0208  & n50435 ;
  assign n51857 = ~n51855 & ~n51856 ;
  assign n51858 = ~n51854 & n51857 ;
  assign n51859 = ~n51853 & n51858 ;
  assign n51860 = ~\pi1157  & n50430 ;
  assign n51861 = ~n51859 & n51860 ;
  assign n51862 = ~\pi0219  & ~n51861 ;
  assign n51863 = ~n51852 & n51862 ;
  assign n51864 = n51844 & n51863 ;
  assign n51865 = ~n51819 & ~n51864 ;
  assign n51866 = ~n51818 & ~n51865 ;
  assign n51867 = ~\pi0214  & ~n51851 ;
  assign n51868 = ~\pi0214  & ~\pi1157  ;
  assign n51869 = ~n51859 & n51868 ;
  assign n51870 = ~n51867 & ~n51869 ;
  assign n51871 = \pi0214  & \pi1157  ;
  assign n51872 = \pi0214  & n51679 ;
  assign n51873 = ~n51596 & n51872 ;
  assign n51874 = ~n51871 & ~n51873 ;
  assign n51875 = n51590 & ~n51874 ;
  assign n51876 = ~\pi0208  & \pi0212  ;
  assign n51877 = ~n50416 & n51876 ;
  assign n51878 = ~n50600 & ~n51877 ;
  assign n51879 = ~n51875 & ~n51878 ;
  assign n51880 = ~\pi0207  & ~n50412 ;
  assign n51881 = \pi1157  & ~n51880 ;
  assign n51882 = \pi1157  & ~n50407 ;
  assign n51883 = ~n50404 & n51882 ;
  assign n51884 = ~n51881 & ~n51883 ;
  assign n51885 = ~\pi1157  & ~n51855 ;
  assign n51886 = ~n51313 & ~n51454 ;
  assign n51887 = n51885 & ~n51886 ;
  assign n51888 = n51884 & ~n51887 ;
  assign n51889 = \pi0208  & ~n50386 ;
  assign n51890 = n50397 & n51889 ;
  assign n51891 = ~n50381 & ~n51890 ;
  assign n51892 = \pi0212  & ~n51891 ;
  assign n51893 = ~n51888 & n51892 ;
  assign n51894 = ~n51879 & ~n51893 ;
  assign n51895 = n51870 & ~n51894 ;
  assign n51896 = ~n50484 & n50556 ;
  assign n51897 = ~n51834 & n51896 ;
  assign n51898 = ~n51840 & n51897 ;
  assign n51899 = ~n51832 & n51898 ;
  assign n51900 = ~n51703 & ~n51899 ;
  assign n51901 = ~n51895 & n51900 ;
  assign n51902 = \pi0211  & ~n51703 ;
  assign n51903 = \pi0219  & ~n51902 ;
  assign n51904 = ~n51901 & n51903 ;
  assign n51905 = n27408 & ~n51904 ;
  assign n51906 = ~n51866 & n51905 ;
  assign n51907 = ~n51765 & ~n51768 ;
  assign n51908 = ~n51773 & ~n51907 ;
  assign n51909 = ~n51906 & n51908 ;
  assign n51910 = ~n51774 & ~n51909 ;
  assign n51911 = ~n51564 & n51910 ;
  assign n51912 = ~\pi0230  & \pi0238  ;
  assign n51913 = ~\pi0211  & n51187 ;
  assign n51914 = n51108 & n51913 ;
  assign n51915 = \pi0200  & \pi0207  ;
  assign n51916 = \pi0208  & n51915 ;
  assign n51917 = n43637 & ~n50876 ;
  assign n51918 = ~n51916 & n51917 ;
  assign n51919 = ~n12409 & n51013 ;
  assign n51920 = ~n50948 & ~n51919 ;
  assign n51921 = n51918 & n51920 ;
  assign n51922 = ~n51914 & ~n51921 ;
  assign n51923 = \pi0219  & n51922 ;
  assign n51924 = ~\pi0299  & ~n51014 ;
  assign n51925 = ~\pi0211  & ~n50412 ;
  assign n51926 = n50411 & n51925 ;
  assign n51927 = ~n51924 & n51926 ;
  assign n51928 = n12255 & n51927 ;
  assign n51929 = \pi0207  & ~n50390 ;
  assign n51930 = ~\pi0207  & \pi0299  ;
  assign n51931 = ~\pi0199  & ~\pi0207  ;
  assign n51932 = ~n51013 & n51931 ;
  assign n51933 = ~n51930 & ~n51932 ;
  assign n51934 = ~n51929 & n51933 ;
  assign n51935 = ~n50412 & n50901 ;
  assign n51936 = n12255 & n51935 ;
  assign n51937 = ~n51934 & n51936 ;
  assign n51938 = ~n51928 & ~n51937 ;
  assign n51939 = n50876 & n51187 ;
  assign n51940 = \pi1153  & ~n13558 ;
  assign n51941 = ~n13646 & ~n51940 ;
  assign n51942 = n50418 & ~n51941 ;
  assign n51943 = ~n51939 & ~n51942 ;
  assign n51944 = \pi0208  & \pi0299  ;
  assign n51945 = ~\pi0199  & \pi0208  ;
  assign n51946 = ~n51915 & n51945 ;
  assign n51947 = ~n51944 & ~n51946 ;
  assign n51948 = ~\pi0200  & ~\pi0207  ;
  assign n51949 = n51001 & n51948 ;
  assign n51950 = ~n50586 & ~n51949 ;
  assign n51951 = ~n51947 & n51950 ;
  assign n51952 = n51943 & ~n51951 ;
  assign n51953 = n12256 & ~n51952 ;
  assign n51954 = n51938 & ~n51953 ;
  assign n51955 = n50411 & n50679 ;
  assign n51956 = ~n51924 & n51955 ;
  assign n51957 = \pi0208  & n50679 ;
  assign n51958 = ~n51934 & n51957 ;
  assign n51959 = ~n51956 & ~n51958 ;
  assign n51960 = \pi0299  & n50610 ;
  assign n51961 = ~n51959 & ~n51960 ;
  assign n51962 = n51922 & ~n51961 ;
  assign n51963 = n51954 & n51962 ;
  assign n51964 = ~n51923 & ~n51963 ;
  assign n51965 = ~\pi0057  & ~\pi1151  ;
  assign n51966 = n6848 & n51965 ;
  assign n51967 = n51964 & n51966 ;
  assign n51968 = ~n51934 & n51935 ;
  assign n51969 = ~n51927 & ~n51968 ;
  assign n51970 = n50371 & n50544 ;
  assign n51971 = ~\pi0207  & n12691 ;
  assign n51972 = \pi0208  & ~\pi0299  ;
  assign n51973 = ~n50370 & n51972 ;
  assign n51974 = ~n51971 & n51973 ;
  assign n51975 = ~n51970 & ~n51974 ;
  assign n51976 = \pi0299  & n50945 ;
  assign n51977 = n12691 & n50945 ;
  assign n51978 = n50877 & n51977 ;
  assign n51979 = ~n51976 & ~n51978 ;
  assign n51980 = n51975 & n51979 ;
  assign n51981 = n51969 & n51980 ;
  assign n51982 = n12255 & ~n51981 ;
  assign n51983 = n12691 & n51033 ;
  assign n51984 = n50877 & n51983 ;
  assign n51985 = ~\pi0219  & ~n51984 ;
  assign n51986 = n51975 & n51985 ;
  assign n51987 = ~n50948 & ~n51986 ;
  assign n51988 = n51015 & ~n51220 ;
  assign n51989 = \pi0208  & ~n51988 ;
  assign n51990 = n50411 & ~n51043 ;
  assign n51991 = ~n51989 & ~n51990 ;
  assign n51992 = n50679 & ~n51960 ;
  assign n51993 = ~n51991 & n51992 ;
  assign n51994 = ~n51987 & ~n51993 ;
  assign n51995 = ~n51982 & n51994 ;
  assign n51996 = ~\pi0057  & \pi1151  ;
  assign n51997 = n6848 & n51996 ;
  assign n51998 = \pi0219  & n51975 ;
  assign n51999 = n51997 & ~n51998 ;
  assign n52000 = ~\pi0211  & \pi0299  ;
  assign n52001 = \pi0211  & \pi0299  ;
  assign n52002 = n12691 & ~n52001 ;
  assign n52003 = n50877 & n52002 ;
  assign n52004 = ~n52000 & ~n52003 ;
  assign n52005 = n15351 & n50877 ;
  assign n52006 = n50570 & ~n52005 ;
  assign n52007 = ~n52004 & ~n52006 ;
  assign n52008 = \pi1153  & n51996 ;
  assign n52009 = n6848 & n52008 ;
  assign n52010 = n52007 & n52009 ;
  assign n52011 = ~n51999 & ~n52010 ;
  assign n52012 = ~n51995 & ~n52011 ;
  assign n52013 = \pi1152  & ~n52012 ;
  assign n52014 = ~n51967 & n52013 ;
  assign n52015 = \pi1153  & n51966 ;
  assign n52016 = n52007 & n52015 ;
  assign n52017 = n50948 & n51966 ;
  assign n52018 = ~\pi1152  & ~n52017 ;
  assign n52019 = ~n52016 & n52018 ;
  assign n52020 = ~n50416 & ~n51984 ;
  assign n52021 = ~\pi0211  & ~n52020 ;
  assign n52022 = n12255 & n51979 ;
  assign n52023 = ~n52021 & n52022 ;
  assign n52024 = \pi0299  & ~n50610 ;
  assign n52025 = ~n51984 & ~n52024 ;
  assign n52026 = n50679 & n52025 ;
  assign n52027 = ~n52023 & ~n52026 ;
  assign n52028 = n51174 & ~n52027 ;
  assign n52029 = ~n52019 & ~n52028 ;
  assign n52030 = ~\pi0209  & n52029 ;
  assign n52031 = n44032 & n50877 ;
  assign n52032 = n50371 & n50641 ;
  assign n52033 = ~n52031 & ~n52032 ;
  assign n52034 = ~\pi0212  & ~n51007 ;
  assign n52035 = ~n52033 & n52034 ;
  assign n52036 = ~n50556 & ~n52035 ;
  assign n52037 = ~\pi1153  & n43637 ;
  assign n52038 = \pi1155  & ~n44035 ;
  assign n52039 = ~n52037 & n52038 ;
  assign n52040 = n44032 & ~n51001 ;
  assign n52041 = ~n52032 & ~n52040 ;
  assign n52042 = ~n52039 & n52041 ;
  assign n52043 = ~n50371 & n50641 ;
  assign n52044 = ~n50435 & n50876 ;
  assign n52045 = ~n50641 & n52044 ;
  assign n52046 = ~n52043 & ~n52045 ;
  assign n52047 = ~\pi0299  & n52046 ;
  assign n52048 = ~n52042 & n52047 ;
  assign n52049 = \pi0214  & ~n52024 ;
  assign n52050 = ~n52048 & n52049 ;
  assign n52051 = ~n52036 & ~n52050 ;
  assign n52052 = n50442 & ~n52046 ;
  assign n52053 = n50442 & ~n52039 ;
  assign n52054 = n52041 & n52053 ;
  assign n52055 = ~n52052 & ~n52054 ;
  assign n52056 = ~\pi1153  & n50430 ;
  assign n52057 = ~n50390 & n52056 ;
  assign n52058 = ~n50371 & n50544 ;
  assign n52059 = \pi0200  & n50410 ;
  assign n52060 = \pi0208  & ~n52059 ;
  assign n52061 = ~n52058 & n52060 ;
  assign n52062 = ~\pi0299  & ~n51597 ;
  assign n52063 = ~\pi0208  & ~n52062 ;
  assign n52064 = n50430 & ~n52063 ;
  assign n52065 = ~n52061 & n52064 ;
  assign n52066 = ~n52057 & ~n52065 ;
  assign n52067 = ~n50416 & n50443 ;
  assign n52068 = \pi0212  & ~n52067 ;
  assign n52069 = \pi0212  & ~n51007 ;
  assign n52070 = ~n52033 & n52069 ;
  assign n52071 = ~n52068 & ~n52070 ;
  assign n52072 = n52066 & ~n52071 ;
  assign n52073 = n52055 & n52072 ;
  assign n52074 = ~n52051 & ~n52073 ;
  assign n52075 = ~\pi0219  & n52074 ;
  assign n52076 = ~\pi0219  & n51996 ;
  assign n52077 = n6848 & n52076 ;
  assign n52078 = \pi0211  & n52033 ;
  assign n52079 = ~\pi0211  & ~n52063 ;
  assign n52080 = ~n52061 & n52079 ;
  assign n52081 = ~n52078 & ~n52080 ;
  assign n52082 = ~n51219 & n52081 ;
  assign n52083 = ~n50570 & n51997 ;
  assign n52084 = ~n51007 & n51997 ;
  assign n52085 = ~n52033 & n52084 ;
  assign n52086 = ~n52083 & ~n52085 ;
  assign n52087 = n52082 & ~n52086 ;
  assign n52088 = ~n52077 & ~n52087 ;
  assign n52089 = ~\pi0209  & ~n52088 ;
  assign n52090 = ~n52075 & n52089 ;
  assign n52091 = ~n52030 & ~n52090 ;
  assign n52092 = ~n52014 & ~n52091 ;
  assign n52093 = n12255 & ~n50946 ;
  assign n52094 = ~\pi0219  & ~n51530 ;
  assign n52095 = ~n52093 & n52094 ;
  assign n52096 = ~\pi1153  & n50689 ;
  assign n52097 = n50677 & ~n52096 ;
  assign n52098 = ~n52095 & n52097 ;
  assign n52099 = ~n52092 & ~n52098 ;
  assign n52100 = \pi0211  & n50556 ;
  assign n52101 = n50556 & n51380 ;
  assign n52102 = ~n52100 & ~n52101 ;
  assign n52103 = \pi0207  & ~n50824 ;
  assign n52104 = ~n51144 & n52103 ;
  assign n52105 = \pi0208  & ~n52104 ;
  assign n52106 = ~n51374 & n52105 ;
  assign n52107 = ~\pi1154  & ~n51100 ;
  assign n52108 = \pi0207  & ~n52107 ;
  assign n52109 = ~n52058 & ~n52108 ;
  assign n52110 = ~n51019 & ~n52109 ;
  assign n52111 = ~n51000 & n52110 ;
  assign n52112 = ~n52100 & ~n52111 ;
  assign n52113 = n52106 & n52112 ;
  assign n52114 = ~n52102 & ~n52113 ;
  assign n52115 = ~n51501 & ~n51504 ;
  assign n52116 = ~\pi0299  & n50460 ;
  assign n52117 = n50371 & n52116 ;
  assign n52118 = ~n51019 & ~n52117 ;
  assign n52119 = ~n51000 & n52118 ;
  assign n52120 = \pi0207  & ~n52119 ;
  assign n52121 = n52115 & ~n52120 ;
  assign n52122 = n50845 & ~n52121 ;
  assign n52123 = ~n51511 & n51512 ;
  assign n52124 = n50852 & ~n52123 ;
  assign n52125 = ~\pi0219  & ~n52124 ;
  assign n52126 = ~n52122 & n52125 ;
  assign n52127 = n52114 & n52126 ;
  assign n52128 = \pi1153  & ~n50432 ;
  assign n52129 = ~n51000 & ~n52128 ;
  assign n52130 = n12409 & ~n52129 ;
  assign n52131 = ~n51490 & ~n52130 ;
  assign n52132 = n51489 & n52131 ;
  assign n52133 = n50430 & ~n52132 ;
  assign n52134 = \pi0212  & ~n52133 ;
  assign n52135 = n50442 & ~n51380 ;
  assign n52136 = n50442 & ~n52111 ;
  assign n52137 = n52106 & n52136 ;
  assign n52138 = ~n52135 & ~n52137 ;
  assign n52139 = n50471 & ~n52121 ;
  assign n52140 = ~\pi0208  & n50443 ;
  assign n52141 = ~n52123 & n52140 ;
  assign n52142 = ~\pi0219  & ~n52141 ;
  assign n52143 = ~n52139 & n52142 ;
  assign n52144 = n52138 & n52143 ;
  assign n52145 = n52134 & n52144 ;
  assign n52146 = ~n52127 & ~n52145 ;
  assign n52147 = n12409 & ~n52117 ;
  assign n52148 = ~n51000 & n52147 ;
  assign n52149 = ~n50876 & ~n52148 ;
  assign n52150 = ~n50570 & n50713 ;
  assign n52151 = ~n52149 & n52150 ;
  assign n52152 = ~n12409 & n52150 ;
  assign n52153 = ~n51368 & n52152 ;
  assign n52154 = ~n52151 & ~n52153 ;
  assign n52155 = n51730 & n52132 ;
  assign n52156 = n50570 & ~n52149 ;
  assign n52157 = ~n51406 & ~n52156 ;
  assign n52158 = n51753 & n52157 ;
  assign n52159 = ~n52155 & n52158 ;
  assign n52160 = n52154 & n52159 ;
  assign n52161 = n52146 & n52160 ;
  assign n52162 = n52099 & ~n52161 ;
  assign n52163 = \pi0213  & ~n52162 ;
  assign n52164 = n50625 & n50679 ;
  assign n52165 = n12257 & ~n52164 ;
  assign n52166 = n50677 & ~n52165 ;
  assign n52167 = \pi1151  & ~n52166 ;
  assign n52168 = \pi0208  & ~n51397 ;
  assign n52169 = ~n52111 & n52168 ;
  assign n52170 = n50571 & ~n51392 ;
  assign n52171 = ~n52169 & n52170 ;
  assign n52172 = \pi0211  & ~n50570 ;
  assign n52173 = ~n52149 & n52172 ;
  assign n52174 = ~n12409 & n52172 ;
  assign n52175 = ~n51368 & n52174 ;
  assign n52176 = ~n52173 & ~n52175 ;
  assign n52177 = ~n52171 & n52176 ;
  assign n52178 = n27408 & n52157 ;
  assign n52179 = n52177 & n52178 ;
  assign n52180 = ~n46751 & ~n52179 ;
  assign n52181 = n52167 & n52180 ;
  assign n52182 = n50967 & n52132 ;
  assign n52183 = ~\pi0214  & ~n52149 ;
  assign n52184 = n50880 & ~n51368 ;
  assign n52185 = ~n52183 & ~n52184 ;
  assign n52186 = n50430 & ~n52149 ;
  assign n52187 = ~n12409 & n50430 ;
  assign n52188 = ~n51368 & n52187 ;
  assign n52189 = ~n52186 & ~n52188 ;
  assign n52190 = n52185 & n52189 ;
  assign n52191 = ~n52182 & n52190 ;
  assign n52192 = ~\pi0212  & ~n52191 ;
  assign n52193 = n50442 & ~n52132 ;
  assign n52194 = n50863 & n52149 ;
  assign n52195 = ~n51412 & n52194 ;
  assign n52196 = \pi0212  & ~n52195 ;
  assign n52197 = ~n52193 & n52196 ;
  assign n52198 = n50967 & n52149 ;
  assign n52199 = ~n51412 & n52198 ;
  assign n52200 = ~n51392 & ~n52169 ;
  assign n52201 = n50430 & ~n52200 ;
  assign n52202 = ~n52199 & ~n52201 ;
  assign n52203 = n52197 & n52202 ;
  assign n52204 = ~n52192 & ~n52203 ;
  assign n52205 = ~\pi0219  & n52167 ;
  assign n52206 = ~n52204 & n52205 ;
  assign n52207 = ~n52181 & ~n52206 ;
  assign n52208 = ~\pi0219  & n50625 ;
  assign n52209 = n50679 & n52208 ;
  assign n52210 = ~n9948 & n52209 ;
  assign n52211 = ~\pi1151  & ~n52210 ;
  assign n52212 = ~\pi0219  & n50679 ;
  assign n52213 = ~\pi0211  & n52212 ;
  assign n52214 = n52132 & n52213 ;
  assign n52215 = \pi0211  & ~n52149 ;
  assign n52216 = ~n51418 & ~n52215 ;
  assign n52217 = n52212 & ~n52216 ;
  assign n52218 = ~n52214 & ~n52217 ;
  assign n52219 = ~n52149 & ~n52212 ;
  assign n52220 = ~n12409 & ~n52212 ;
  assign n52221 = ~n51368 & n52220 ;
  assign n52222 = ~n52219 & ~n52221 ;
  assign n52223 = n27408 & n52222 ;
  assign n52224 = n52218 & n52223 ;
  assign n52225 = n52211 & ~n52224 ;
  assign n52226 = ~\pi1152  & ~n52225 ;
  assign n52227 = n52207 & n52226 ;
  assign n52228 = \pi0209  & ~n52227 ;
  assign n52229 = ~n9948 & n51169 ;
  assign n52230 = ~\pi0211  & ~\pi1153  ;
  assign n52231 = ~n12255 & n52230 ;
  assign n52232 = n52229 & ~n52231 ;
  assign n52233 = ~n12257 & n50677 ;
  assign n52234 = \pi1151  & ~n52233 ;
  assign n52235 = ~n52232 & n52234 ;
  assign n52236 = n50430 & ~n51392 ;
  assign n52237 = ~n52169 & n52236 ;
  assign n52238 = ~n52182 & ~n52237 ;
  assign n52239 = ~\pi0212  & n52185 ;
  assign n52240 = n52238 & n52239 ;
  assign n52241 = \pi0212  & ~n50442 ;
  assign n52242 = ~n52200 & n52241 ;
  assign n52243 = \pi0212  & n50442 ;
  assign n52244 = ~n52132 & n52243 ;
  assign n52245 = ~n52242 & ~n52244 ;
  assign n52246 = ~\pi0219  & n52245 ;
  assign n52247 = ~n52240 & n52246 ;
  assign n52248 = ~n52180 & ~n52247 ;
  assign n52249 = n52235 & ~n52248 ;
  assign n52250 = \pi1151  & \pi1152  ;
  assign n52251 = \pi1152  & ~n52231 ;
  assign n52252 = n52229 & n52251 ;
  assign n52253 = ~n52250 & ~n52252 ;
  assign n52254 = ~\pi0219  & ~n52240 ;
  assign n52255 = n50863 & ~n52200 ;
  assign n52256 = ~n52193 & ~n52255 ;
  assign n52257 = n50967 & ~n52200 ;
  assign n52258 = n50430 & n52149 ;
  assign n52259 = ~n51412 & n52258 ;
  assign n52260 = ~n52257 & ~n52259 ;
  assign n52261 = n52256 & n52260 ;
  assign n52262 = \pi0212  & ~n52261 ;
  assign n52263 = n52254 & ~n52262 ;
  assign n52264 = \pi0219  & ~n52149 ;
  assign n52265 = n50938 & ~n51368 ;
  assign n52266 = ~n52264 & ~n52265 ;
  assign n52267 = n50998 & n52266 ;
  assign n52268 = ~n52263 & n52267 ;
  assign n52269 = n52253 & ~n52268 ;
  assign n52270 = ~n52249 & ~n52269 ;
  assign n52271 = n52228 & ~n52270 ;
  assign n52272 = ~n52163 & n52271 ;
  assign n52273 = ~\pi0214  & \pi1153  ;
  assign n52274 = ~\pi0214  & ~\pi0299  ;
  assign n52275 = ~n12691 & n52274 ;
  assign n52276 = ~n52273 & ~n52275 ;
  assign n52277 = n52081 & ~n52276 ;
  assign n52278 = \pi0214  & ~n51007 ;
  assign n52279 = ~n52033 & n52278 ;
  assign n52280 = \pi0212  & ~n52001 ;
  assign n52281 = ~n51984 & n52280 ;
  assign n52282 = ~n50600 & ~n52281 ;
  assign n52283 = ~n52279 & ~n52282 ;
  assign n52284 = ~\pi0219  & n52283 ;
  assign n52285 = ~n52277 & n52284 ;
  assign n52286 = ~n51007 & ~n52033 ;
  assign n52287 = n50570 & ~n52286 ;
  assign n52288 = n52082 & ~n52287 ;
  assign n52289 = n51819 & ~n52288 ;
  assign n52290 = ~n52285 & ~n52289 ;
  assign n52291 = ~n51984 & ~n52001 ;
  assign n52292 = ~\pi0214  & ~n52005 ;
  assign n52293 = \pi0212  & ~n52292 ;
  assign n52294 = ~n52291 & n52293 ;
  assign n52295 = ~\pi0219  & ~n52005 ;
  assign n52296 = ~\pi0212  & n50967 ;
  assign n52297 = n51187 & n52296 ;
  assign n52298 = n52295 & ~n52297 ;
  assign n52299 = ~n52294 & n52298 ;
  assign n52300 = \pi1153  & n52292 ;
  assign n52301 = n52007 & n52300 ;
  assign n52302 = n52211 & ~n52301 ;
  assign n52303 = n52299 & n52302 ;
  assign n52304 = \pi0219  & ~n52005 ;
  assign n52305 = ~\pi0057  & \pi1153  ;
  assign n52306 = n6848 & n52305 ;
  assign n52307 = ~n52304 & n52306 ;
  assign n52308 = n52007 & n52307 ;
  assign n52309 = n52211 & ~n52308 ;
  assign n52310 = ~n51984 & ~n52000 ;
  assign n52311 = ~n50570 & ~n52310 ;
  assign n52312 = ~n52286 & ~n52311 ;
  assign n52313 = \pi0219  & n52312 ;
  assign n52314 = ~n52309 & ~n52313 ;
  assign n52315 = ~n52303 & n52314 ;
  assign n52316 = n27408 & n52315 ;
  assign n52317 = n52290 & n52316 ;
  assign n52318 = ~n52167 & ~n52309 ;
  assign n52319 = ~n52303 & n52318 ;
  assign n52320 = ~\pi0209  & ~\pi1152  ;
  assign n52321 = ~n52319 & n52320 ;
  assign n52322 = ~n52317 & n52321 ;
  assign n52323 = \pi0211  & n51990 ;
  assign n52324 = n50845 & ~n51988 ;
  assign n52325 = ~n52323 & ~n52324 ;
  assign n52326 = \pi1153  & n12691 ;
  assign n52327 = n50877 & n52326 ;
  assign n52328 = ~n51187 & ~n52327 ;
  assign n52329 = ~\pi0214  & n51975 ;
  assign n52330 = n52328 & n52329 ;
  assign n52331 = n52325 & n52330 ;
  assign n52332 = \pi0214  & ~n51990 ;
  assign n52333 = ~n51989 & n52332 ;
  assign n52334 = \pi0212  & ~n52333 ;
  assign n52335 = ~n52331 & n52334 ;
  assign n52336 = ~\pi0219  & ~n52335 ;
  assign n52337 = \pi0214  & n52328 ;
  assign n52338 = n51975 & n52337 ;
  assign n52339 = n52325 & n52338 ;
  assign n52340 = ~\pi0214  & ~n51984 ;
  assign n52341 = n51975 & n52340 ;
  assign n52342 = ~\pi0212  & ~n52341 ;
  assign n52343 = ~n52339 & n52342 ;
  assign n52344 = n52235 & ~n52343 ;
  assign n52345 = n52336 & n52344 ;
  assign n52346 = ~\pi1151  & ~n52232 ;
  assign n52347 = n51918 & ~n51919 ;
  assign n52348 = \pi0219  & ~n52347 ;
  assign n52349 = n9948 & ~n52348 ;
  assign n52350 = n52346 & ~n52349 ;
  assign n52351 = ~\pi0211  & ~n51951 ;
  assign n52352 = n51943 & n52351 ;
  assign n52353 = ~n51959 & ~n52352 ;
  assign n52354 = ~n50679 & ~n51919 ;
  assign n52355 = n51918 & n52354 ;
  assign n52356 = n12255 & n52000 ;
  assign n52357 = ~\pi0219  & ~n52356 ;
  assign n52358 = ~n52355 & n52357 ;
  assign n52359 = n52346 & n52358 ;
  assign n52360 = ~n52353 & n52359 ;
  assign n52361 = ~n52350 & ~n52360 ;
  assign n52362 = n50571 & n51990 ;
  assign n52363 = \pi0208  & n50571 ;
  assign n52364 = ~n51988 & n52363 ;
  assign n52365 = ~n52362 & ~n52364 ;
  assign n52366 = \pi0219  & ~n51984 ;
  assign n52367 = n51975 & n52366 ;
  assign n52368 = n52365 & n52367 ;
  assign n52369 = n9948 & ~n52368 ;
  assign n52370 = n52235 & ~n52369 ;
  assign n52371 = n52361 & ~n52370 ;
  assign n52372 = ~n52345 & n52371 ;
  assign n52373 = ~\pi0209  & \pi1152  ;
  assign n52374 = ~n52372 & n52373 ;
  assign n52375 = ~\pi0213  & ~n52374 ;
  assign n52376 = ~n52322 & n52375 ;
  assign n52377 = ~n52163 & ~n52376 ;
  assign n52378 = \pi0230  & ~n52377 ;
  assign n52379 = ~n52272 & n52378 ;
  assign n52380 = ~n51912 & ~n52379 ;
  assign n52381 = ~\pi0230  & ~\pi0239  ;
  assign n52382 = ~\pi0214  & n50418 ;
  assign n52383 = ~n50397 & n52382 ;
  assign n52384 = n51819 & ~n52383 ;
  assign n52385 = ~n50868 & n51128 ;
  assign n52386 = n50496 & n51128 ;
  assign n52387 = ~n50393 & n52386 ;
  assign n52388 = ~n52385 & ~n52387 ;
  assign n52389 = \pi0211  & ~n50435 ;
  assign n52390 = \pi0214  & ~n52389 ;
  assign n52391 = \pi0214  & n50437 ;
  assign n52392 = ~n50833 & n52391 ;
  assign n52393 = ~n52390 & ~n52392 ;
  assign n52394 = n52388 & ~n52393 ;
  assign n52395 = n52384 & ~n52394 ;
  assign n52396 = ~\pi0212  & \pi0219  ;
  assign n52397 = ~n52383 & n52396 ;
  assign n52398 = ~n50386 & ~n50416 ;
  assign n52399 = n50397 & n52398 ;
  assign n52400 = \pi0211  & ~n50396 ;
  assign n52401 = ~n50393 & n52400 ;
  assign n52402 = \pi0211  & ~n50418 ;
  assign n52403 = \pi0214  & ~n52402 ;
  assign n52404 = ~n50416 & ~n50418 ;
  assign n52405 = n52403 & ~n52404 ;
  assign n52406 = ~n52401 & n52405 ;
  assign n52407 = ~n52399 & n52406 ;
  assign n52408 = n52397 & ~n52407 ;
  assign n52409 = \pi0212  & ~n50418 ;
  assign n52410 = \pi0212  & ~n50396 ;
  assign n52411 = ~n50393 & n52410 ;
  assign n52412 = ~n52409 & ~n52411 ;
  assign n52413 = n9948 & n52412 ;
  assign n52414 = ~n52408 & n52413 ;
  assign n52415 = ~n52395 & n52414 ;
  assign n52416 = ~n9948 & ~n51164 ;
  assign n52417 = \pi0219  & n50556 ;
  assign n52418 = ~n51161 & ~n52417 ;
  assign n52419 = n52416 & ~n52418 ;
  assign n52420 = ~\pi0209  & ~\pi0213  ;
  assign n52421 = ~n52419 & n52420 ;
  assign n52422 = ~n52415 & n52421 ;
  assign n52423 = ~n51683 & n51684 ;
  assign n52424 = ~\pi0214  & \pi1157  ;
  assign n52425 = ~\pi0214  & n51679 ;
  assign n52426 = ~n51596 & n52425 ;
  assign n52427 = ~n52424 & ~n52426 ;
  assign n52428 = n52423 & ~n52427 ;
  assign n52429 = n52396 & ~n52428 ;
  assign n52430 = ~\pi0211  & ~n50416 ;
  assign n52431 = ~n51655 & n52430 ;
  assign n52432 = ~n51874 & n52423 ;
  assign n52433 = ~n50967 & ~n52432 ;
  assign n52434 = ~n52431 & ~n52433 ;
  assign n52435 = n52429 & ~n52434 ;
  assign n52436 = \pi0212  & ~n52423 ;
  assign n52437 = \pi0212  & ~\pi1157  ;
  assign n52438 = ~n51855 & n52437 ;
  assign n52439 = ~n52436 & ~n52438 ;
  assign n52440 = n9948 & n52439 ;
  assign n52441 = n51819 & ~n52428 ;
  assign n52442 = n52440 & ~n52441 ;
  assign n52443 = ~n51655 & n52389 ;
  assign n52444 = n51128 & ~n52423 ;
  assign n52445 = ~\pi1157  & n51128 ;
  assign n52446 = ~n51855 & n52445 ;
  assign n52447 = ~n52444 & ~n52446 ;
  assign n52448 = \pi0214  & n52447 ;
  assign n52449 = n52440 & n52448 ;
  assign n52450 = ~n52443 & n52449 ;
  assign n52451 = ~n52442 & ~n52450 ;
  assign n52452 = ~n52435 & ~n52451 ;
  assign n52453 = ~\pi0213  & ~n52419 ;
  assign n52454 = \pi0209  & n52453 ;
  assign n52455 = ~n52452 & n52454 ;
  assign n52456 = ~n52422 & ~n52455 ;
  assign n52457 = ~n50418 & n51785 ;
  assign n52458 = n50418 & ~n51777 ;
  assign n52459 = ~n51775 & n52458 ;
  assign n52460 = ~n52457 & ~n52459 ;
  assign n52461 = n50967 & ~n52460 ;
  assign n52462 = \pi1157  & ~n51944 ;
  assign n52463 = ~n50411 & n52462 ;
  assign n52464 = \pi0207  & n52462 ;
  assign n52465 = n50541 & n52464 ;
  assign n52466 = ~n52463 & ~n52465 ;
  assign n52467 = ~\pi1157  & ~n50418 ;
  assign n52468 = ~\pi1157  & ~n50396 ;
  assign n52469 = ~n50393 & n52468 ;
  assign n52470 = ~n52467 & ~n52469 ;
  assign n52471 = n50430 & n52470 ;
  assign n52472 = n52466 & n52471 ;
  assign n52473 = n52384 & ~n52472 ;
  assign n52474 = ~n52461 & n52473 ;
  assign n52475 = ~\pi0057  & ~\pi0209  ;
  assign n52476 = n6848 & n52475 ;
  assign n52477 = n52412 & n52476 ;
  assign n52478 = ~n52397 & n52477 ;
  assign n52479 = ~n52401 & n52403 ;
  assign n52480 = n52388 & n52479 ;
  assign n52481 = n52477 & n52480 ;
  assign n52482 = ~n52478 & ~n52481 ;
  assign n52483 = ~n52474 & ~n52482 ;
  assign n52484 = \pi0208  & ~n51785 ;
  assign n52485 = ~n50452 & ~n52484 ;
  assign n52486 = ~n51791 & n52485 ;
  assign n52487 = n51797 & ~n52486 ;
  assign n52488 = ~\pi0299  & n52462 ;
  assign n52489 = n51683 & n52488 ;
  assign n52490 = ~n52463 & ~n52489 ;
  assign n52491 = ~n51885 & n52490 ;
  assign n52492 = \pi0211  & ~n52491 ;
  assign n52493 = \pi0214  & ~n52492 ;
  assign n52494 = ~n52487 & n52493 ;
  assign n52495 = n52441 & ~n52494 ;
  assign n52496 = \pi0209  & n9948 ;
  assign n52497 = n52439 & n52496 ;
  assign n52498 = \pi0211  & ~n52423 ;
  assign n52499 = n51347 & ~n51855 ;
  assign n52500 = ~n52498 & ~n52499 ;
  assign n52501 = n52448 & n52500 ;
  assign n52502 = n52429 & ~n52501 ;
  assign n52503 = n52497 & ~n52502 ;
  assign n52504 = ~n52495 & n52503 ;
  assign n52505 = ~n51740 & n51763 ;
  assign n52506 = \pi0213  & ~n52505 ;
  assign n52507 = ~n52504 & n52506 ;
  assign n52508 = ~n52483 & n52507 ;
  assign n52509 = n52456 & ~n52508 ;
  assign n52510 = \pi0230  & ~n52509 ;
  assign n52511 = ~n52381 & ~n52510 ;
  assign n52512 = n12257 & ~n50805 ;
  assign n52513 = n50677 & ~n52512 ;
  assign n52514 = \pi1147  & n52513 ;
  assign n52515 = ~\pi0199  & \pi1146  ;
  assign n52516 = \pi0199  & \pi1145  ;
  assign n52517 = ~\pi0200  & ~n52516 ;
  assign n52518 = ~n52515 & n52517 ;
  assign n52519 = \pi0200  & ~n51721 ;
  assign n52520 = n50544 & ~n52519 ;
  assign n52521 = ~n52518 & n52520 ;
  assign n52522 = ~n50877 & ~n52521 ;
  assign n52523 = \pi0200  & ~n52515 ;
  assign n52524 = ~\pi0299  & ~n52523 ;
  assign n52525 = n50383 & ~n52516 ;
  assign n52526 = n52524 & ~n52525 ;
  assign n52527 = ~n12409 & ~n52526 ;
  assign n52528 = ~n52522 & ~n52527 ;
  assign n52529 = ~n50571 & n52528 ;
  assign n52530 = \pi0219  & ~n52529 ;
  assign n52531 = n50418 & ~n52525 ;
  assign n52532 = n52524 & n52531 ;
  assign n52533 = ~\pi0208  & ~n52532 ;
  assign n52534 = ~\pi0299  & n52533 ;
  assign n52535 = \pi0299  & \pi1146  ;
  assign n52536 = ~n52521 & ~n52535 ;
  assign n52537 = ~n51449 & ~n52525 ;
  assign n52538 = n52524 & n52537 ;
  assign n52539 = ~\pi0299  & ~n52538 ;
  assign n52540 = n52536 & n52539 ;
  assign n52541 = ~n52534 & ~n52540 ;
  assign n52542 = n50571 & n52541 ;
  assign n52543 = n52530 & ~n52542 ;
  assign n52544 = n9948 & ~n52543 ;
  assign n52545 = ~\pi0219  & ~n52528 ;
  assign n52546 = \pi0212  & ~n50443 ;
  assign n52547 = ~n52296 & ~n52546 ;
  assign n52548 = n52541 & ~n52547 ;
  assign n52549 = n52545 & ~n52548 ;
  assign n52550 = \pi1147  & ~n52549 ;
  assign n52551 = n52544 & n52550 ;
  assign n52552 = ~n52514 & ~n52551 ;
  assign n52553 = n44032 & n52516 ;
  assign n52554 = n44035 & n52515 ;
  assign n52555 = ~n52553 & ~n52554 ;
  assign n52556 = ~n12409 & n52555 ;
  assign n52557 = ~\pi0057  & ~\pi1147  ;
  assign n52558 = n6848 & n52557 ;
  assign n52559 = ~n52556 & n52558 ;
  assign n52560 = ~n52522 & n52559 ;
  assign n52561 = ~\pi0211  & ~\pi1147  ;
  assign n52562 = ~\pi0219  & n52561 ;
  assign n52563 = n50679 & n52562 ;
  assign n52564 = ~n52560 & ~n52563 ;
  assign n52565 = ~\pi0207  & ~n52525 ;
  assign n52566 = n52524 & n52565 ;
  assign n52567 = n52536 & ~n52566 ;
  assign n52568 = n52517 & n52566 ;
  assign n52569 = \pi0208  & ~n52568 ;
  assign n52570 = ~n52567 & n52569 ;
  assign n52571 = n50418 & ~n52555 ;
  assign n52572 = n12577 & n50679 ;
  assign n52573 = n20516 & n52572 ;
  assign n52574 = ~n52571 & n52573 ;
  assign n52575 = ~n52570 & n52574 ;
  assign n52576 = ~n52564 & ~n52575 ;
  assign n52577 = \pi1149  & ~n52576 ;
  assign n52578 = n52552 & n52577 ;
  assign n52579 = ~\pi1148  & ~n52578 ;
  assign n52580 = \pi0211  & n52541 ;
  assign n52581 = \pi0212  & n52580 ;
  assign n52582 = ~\pi0299  & ~n52571 ;
  assign n52583 = ~n52570 & n52582 ;
  assign n52584 = n12255 & ~n52583 ;
  assign n52585 = ~n52581 & ~n52584 ;
  assign n52586 = n50430 & n52541 ;
  assign n52587 = n52545 & ~n52586 ;
  assign n52588 = n52585 & n52587 ;
  assign n52589 = n52544 & ~n52549 ;
  assign n52590 = ~n52588 & n52589 ;
  assign n52591 = ~\pi1149  & ~n52233 ;
  assign n52592 = ~n52560 & n52591 ;
  assign n52593 = ~n52590 & n52592 ;
  assign n52594 = ~\pi1147  & ~\pi1149  ;
  assign n52595 = ~n52560 & n52594 ;
  assign n52596 = ~\pi0209  & ~n52595 ;
  assign n52597 = ~n52593 & n52596 ;
  assign n52598 = n52579 & n52597 ;
  assign n52599 = ~\pi0211  & n52541 ;
  assign n52600 = \pi0212  & n50954 ;
  assign n52601 = ~n52528 & n52600 ;
  assign n52602 = ~n52599 & n52601 ;
  assign n52603 = ~\pi0299  & ~n50570 ;
  assign n52604 = ~n52571 & n52603 ;
  assign n52605 = ~\pi0219  & n52604 ;
  assign n52606 = ~n52570 & n52605 ;
  assign n52607 = ~n50948 & n52556 ;
  assign n52608 = ~n50877 & ~n50948 ;
  assign n52609 = ~n52521 & n52608 ;
  assign n52610 = ~n52607 & ~n52609 ;
  assign n52611 = n9948 & n52610 ;
  assign n52612 = ~n52606 & n52611 ;
  assign n52613 = ~n52602 & n52612 ;
  assign n52614 = ~\pi1147  & ~n52229 ;
  assign n52615 = ~n52613 & n52614 ;
  assign n52616 = \pi0299  & ~n50570 ;
  assign n52617 = ~\pi0219  & ~n52616 ;
  assign n52618 = ~n52528 & n52617 ;
  assign n52619 = n9948 & ~n52618 ;
  assign n52620 = ~n52543 & n52619 ;
  assign n52621 = ~n9948 & n50714 ;
  assign n52622 = \pi1147  & ~n52621 ;
  assign n52623 = ~n52620 & n52622 ;
  assign n52624 = ~n52615 & ~n52623 ;
  assign n52625 = \pi1149  & n52624 ;
  assign n52626 = ~\pi0209  & \pi1148  ;
  assign n52627 = n52625 & n52626 ;
  assign n52628 = ~\pi0219  & ~n9948 ;
  assign n52629 = \pi0212  & n50443 ;
  assign n52630 = ~n52100 & ~n52629 ;
  assign n52631 = n52628 & ~n52630 ;
  assign n52632 = ~\pi1147  & ~n52631 ;
  assign n52633 = n50570 & ~n52556 ;
  assign n52634 = ~n52522 & n52633 ;
  assign n52635 = n52587 & ~n52634 ;
  assign n52636 = n52585 & n52635 ;
  assign n52637 = n52613 & ~n52636 ;
  assign n52638 = n52632 & ~n52637 ;
  assign n52639 = ~\pi0219  & ~n52241 ;
  assign n52640 = ~n52100 & n52639 ;
  assign n52641 = n50677 & ~n52640 ;
  assign n52642 = \pi1147  & ~n52641 ;
  assign n52643 = n52587 & n52642 ;
  assign n52644 = n52585 & n52643 ;
  assign n52645 = ~\pi1149  & ~n52642 ;
  assign n52646 = ~\pi1149  & n9948 ;
  assign n52647 = ~n52543 & n52646 ;
  assign n52648 = ~n52645 & ~n52647 ;
  assign n52649 = ~n52644 & ~n52648 ;
  assign n52650 = n52626 & n52649 ;
  assign n52651 = ~n52638 & n52650 ;
  assign n52652 = ~n52627 & ~n52651 ;
  assign n52653 = ~n52598 & n52652 ;
  assign n52654 = ~n52061 & ~n52063 ;
  assign n52655 = \pi0211  & ~n52654 ;
  assign n52656 = ~\pi0211  & ~n52033 ;
  assign n52657 = \pi0214  & ~n52656 ;
  assign n52658 = ~n52655 & n52657 ;
  assign n52659 = n12255 & ~n52658 ;
  assign n52660 = \pi0212  & ~\pi0219  ;
  assign n52661 = ~\pi0214  & ~\pi0219  ;
  assign n52662 = n52033 & n52661 ;
  assign n52663 = ~n52660 & ~n52662 ;
  assign n52664 = n50954 & ~n52081 ;
  assign n52665 = n52663 & ~n52664 ;
  assign n52666 = \pi0212  & n52081 ;
  assign n52667 = ~n52658 & n52666 ;
  assign n52668 = ~n52665 & ~n52667 ;
  assign n52669 = ~n52659 & n52668 ;
  assign n52670 = ~\pi0214  & n52033 ;
  assign n52671 = ~\pi0212  & ~n52670 ;
  assign n52672 = \pi0214  & ~n52081 ;
  assign n52673 = n52671 & ~n52672 ;
  assign n52674 = \pi0219  & ~n52666 ;
  assign n52675 = ~n52673 & n52674 ;
  assign n52676 = n9948 & ~n52675 ;
  assign n52677 = ~n52669 & n52676 ;
  assign n52678 = \pi1147  & ~n52513 ;
  assign n52679 = ~n52677 & n52678 ;
  assign n52680 = n12691 & n50877 ;
  assign n52681 = n20516 & n52680 ;
  assign n52682 = ~n20516 & n52572 ;
  assign n52683 = ~n52681 & ~n52682 ;
  assign n52684 = ~\pi1147  & n52683 ;
  assign n52685 = ~\pi1148  & \pi1149  ;
  assign n52686 = ~n52684 & n52685 ;
  assign n52687 = ~n52679 & n52686 ;
  assign n52688 = \pi1147  & ~\pi1149  ;
  assign n52689 = ~n12257 & n52688 ;
  assign n52690 = n50677 & n52689 ;
  assign n52691 = ~\pi1148  & n52690 ;
  assign n52692 = ~\pi0211  & n50693 ;
  assign n52693 = ~\pi0219  & ~n52692 ;
  assign n52694 = n51975 & n52693 ;
  assign n52695 = ~n52660 & ~n52694 ;
  assign n52696 = ~\pi0214  & ~n52000 ;
  assign n52697 = n51975 & n52696 ;
  assign n52698 = \pi0212  & ~n52697 ;
  assign n52699 = \pi0214  & ~n52001 ;
  assign n52700 = n51975 & n52699 ;
  assign n52701 = n52698 & ~n52700 ;
  assign n52702 = ~n52695 & ~n52701 ;
  assign n52703 = ~\pi0199  & ~\pi0208  ;
  assign n52704 = ~\pi0199  & ~n51915 ;
  assign n52705 = n50384 & n52704 ;
  assign n52706 = ~n52703 & ~n52705 ;
  assign n52707 = ~n51975 & n52706 ;
  assign n52708 = ~\pi0299  & ~n52707 ;
  assign n52709 = n9948 & ~n51975 ;
  assign n52710 = n9948 & ~n50676 ;
  assign n52711 = \pi0219  & ~n52000 ;
  assign n52712 = n52710 & ~n52711 ;
  assign n52713 = ~n52709 & ~n52712 ;
  assign n52714 = ~n52708 & ~n52713 ;
  assign n52715 = ~n52702 & n52714 ;
  assign n52716 = \pi0299  & n50430 ;
  assign n52717 = ~\pi0212  & ~n52716 ;
  assign n52718 = n51975 & n52717 ;
  assign n52719 = ~\pi0214  & n52001 ;
  assign n52720 = \pi0212  & ~n52719 ;
  assign n52721 = ~n52692 & n52720 ;
  assign n52722 = n51975 & n52721 ;
  assign n52723 = ~n52718 & ~n52722 ;
  assign n52724 = n12577 & ~n52723 ;
  assign n52725 = ~\pi0219  & ~\pi0299  ;
  assign n52726 = ~\pi0211  & n52725 ;
  assign n52727 = ~n52707 & n52726 ;
  assign n52728 = n52688 & ~n52727 ;
  assign n52729 = ~n52724 & n52728 ;
  assign n52730 = ~\pi1148  & n52729 ;
  assign n52731 = n52715 & n52730 ;
  assign n52732 = ~n52691 & ~n52731 ;
  assign n52733 = n52616 & n52710 ;
  assign n52734 = ~n52640 & n52733 ;
  assign n52735 = ~n52709 & ~n52734 ;
  assign n52736 = n52642 & n52735 ;
  assign n52737 = ~n50877 & ~n51929 ;
  assign n52738 = ~\pi0299  & ~n51971 ;
  assign n52739 = ~n12409 & n51178 ;
  assign n52740 = n52738 & ~n52739 ;
  assign n52741 = ~n52737 & n52740 ;
  assign n52742 = \pi0219  & ~n52741 ;
  assign n52743 = n9948 & ~n52742 ;
  assign n52744 = n52632 & ~n52743 ;
  assign n52745 = ~n52736 & ~n52744 ;
  assign n52746 = ~\pi1149  & ~n52745 ;
  assign n52747 = ~\pi0299  & n52739 ;
  assign n52748 = ~\pi0299  & ~n50877 ;
  assign n52749 = ~n51929 & n52748 ;
  assign n52750 = ~n52747 & ~n52749 ;
  assign n52751 = ~\pi0207  & \pi0211  ;
  assign n52752 = n12691 & n52751 ;
  assign n52753 = ~n52001 & ~n52752 ;
  assign n52754 = \pi0214  & ~n52753 ;
  assign n52755 = n52750 & ~n52754 ;
  assign n52756 = \pi0212  & ~n52755 ;
  assign n52757 = n50570 & ~n52741 ;
  assign n52758 = n50556 & ~n52750 ;
  assign n52759 = ~n52757 & ~n52758 ;
  assign n52760 = ~n52756 & n52759 ;
  assign n52761 = \pi0214  & n52750 ;
  assign n52762 = ~n52001 & ~n52741 ;
  assign n52763 = ~n52761 & n52762 ;
  assign n52764 = \pi0212  & ~n52763 ;
  assign n52765 = n52760 & n52764 ;
  assign n52766 = ~\pi0219  & ~n52716 ;
  assign n52767 = ~n52741 & n52766 ;
  assign n52768 = ~n52660 & ~n52767 ;
  assign n52769 = n52632 & ~n52768 ;
  assign n52770 = ~\pi1149  & n52769 ;
  assign n52771 = ~n52765 & n52770 ;
  assign n52772 = ~n52746 & ~n52771 ;
  assign n52773 = ~\pi0214  & ~n51918 ;
  assign n52774 = ~\pi0212  & ~n52773 ;
  assign n52775 = n13550 & n50418 ;
  assign n52776 = \pi0214  & ~\pi0299  ;
  assign n52777 = ~n52775 & n52776 ;
  assign n52778 = n51947 & n52777 ;
  assign n52779 = n52774 & ~n52778 ;
  assign n52780 = ~\pi0219  & ~n52779 ;
  assign n52781 = ~\pi0299  & ~n52775 ;
  assign n52782 = n51947 & n52781 ;
  assign n52783 = \pi0212  & ~n52782 ;
  assign n52784 = ~\pi0211  & ~n52782 ;
  assign n52785 = \pi0211  & n51918 ;
  assign n52786 = \pi0214  & ~n52785 ;
  assign n52787 = ~n52784 & n52786 ;
  assign n52788 = n52783 & ~n52787 ;
  assign n52789 = n52780 & ~n52788 ;
  assign n52790 = n9948 & n51918 ;
  assign n52791 = ~\pi1147  & n52790 ;
  assign n52792 = ~\pi1147  & n9948 ;
  assign n52793 = ~n52304 & n52792 ;
  assign n52794 = ~n52791 & ~n52793 ;
  assign n52795 = ~n52789 & ~n52794 ;
  assign n52796 = ~\pi1147  & n52229 ;
  assign n52797 = ~\pi1147  & \pi1149  ;
  assign n52798 = n50824 & ~n50876 ;
  assign n52799 = n9948 & n52798 ;
  assign n52800 = ~n52733 & ~n52799 ;
  assign n52801 = \pi1149  & ~n52621 ;
  assign n52802 = n52800 & n52801 ;
  assign n52803 = ~n52797 & ~n52802 ;
  assign n52804 = ~n52796 & ~n52803 ;
  assign n52805 = ~n52795 & n52804 ;
  assign n52806 = \pi1148  & ~n52805 ;
  assign n52807 = n52772 & n52806 ;
  assign n52808 = n52732 & ~n52807 ;
  assign n52809 = ~n52687 & n52808 ;
  assign n52810 = \pi0209  & ~n52809 ;
  assign n52811 = \pi0213  & \pi0230  ;
  assign n52812 = ~n52810 & n52811 ;
  assign n52813 = n52653 & n52812 ;
  assign n52814 = \pi0211  & \pi1146  ;
  assign n52815 = n50600 & n52814 ;
  assign n52816 = ~\pi0211  & \pi1146  ;
  assign n52817 = \pi0211  & \pi1145  ;
  assign n52818 = ~n52816 & ~n52817 ;
  assign n52819 = n12255 & ~n52818 ;
  assign n52820 = ~n52815 & ~n52819 ;
  assign n52821 = n50556 & n52814 ;
  assign n52822 = ~n51108 & ~n52821 ;
  assign n52823 = n52820 & n52822 ;
  assign n52824 = \pi0219  & ~n51665 ;
  assign n52825 = ~n27408 & ~n52824 ;
  assign n52826 = ~n52823 & n52825 ;
  assign n52827 = ~n9948 & n52572 ;
  assign n52828 = \pi1147  & ~n52827 ;
  assign n52829 = ~n52826 & n52828 ;
  assign n52830 = n50571 & ~n51640 ;
  assign n52831 = n52541 & n52830 ;
  assign n52832 = n52530 & ~n52831 ;
  assign n52833 = n27408 & ~n52832 ;
  assign n52834 = n52829 & ~n52833 ;
  assign n52835 = \pi0211  & ~n51640 ;
  assign n52836 = n52541 & n52835 ;
  assign n52837 = \pi0299  & ~n52818 ;
  assign n52838 = \pi0214  & ~n52837 ;
  assign n52839 = n52533 & n52838 ;
  assign n52840 = ~n52538 & n52838 ;
  assign n52841 = n52536 & n52840 ;
  assign n52842 = ~n52839 & ~n52841 ;
  assign n52843 = ~n52586 & n52842 ;
  assign n52844 = ~n52836 & ~n52843 ;
  assign n52845 = \pi0211  & ~\pi1146  ;
  assign n52846 = \pi0299  & ~n52845 ;
  assign n52847 = ~\pi0214  & ~n52846 ;
  assign n52848 = n52533 & n52847 ;
  assign n52849 = ~n52538 & n52847 ;
  assign n52850 = n52536 & n52849 ;
  assign n52851 = ~n52848 & ~n52850 ;
  assign n52852 = \pi0212  & n52851 ;
  assign n52853 = ~n52844 & n52852 ;
  assign n52854 = \pi0211  & n52535 ;
  assign n52855 = n52556 & ~n52854 ;
  assign n52856 = ~n50877 & ~n52854 ;
  assign n52857 = ~n52521 & n52856 ;
  assign n52858 = ~n52855 & ~n52857 ;
  assign n52859 = n50878 & ~n52521 ;
  assign n52860 = n50880 & n52555 ;
  assign n52861 = ~\pi0212  & ~n52860 ;
  assign n52862 = ~n52859 & n52861 ;
  assign n52863 = n52858 & n52862 ;
  assign n52864 = ~\pi0219  & ~n52863 ;
  assign n52865 = ~\pi0214  & ~n52528 ;
  assign n52866 = ~\pi0212  & ~n52865 ;
  assign n52867 = n52829 & ~n52866 ;
  assign n52868 = ~n52528 & n52829 ;
  assign n52869 = ~n52599 & n52868 ;
  assign n52870 = ~n52867 & ~n52869 ;
  assign n52871 = n52864 & ~n52870 ;
  assign n52872 = ~n52853 & n52871 ;
  assign n52873 = ~n52834 & ~n52872 ;
  assign n52874 = ~\pi1147  & ~n52825 ;
  assign n52875 = ~\pi1147  & n52822 ;
  assign n52876 = n52820 & n52875 ;
  assign n52877 = ~n52874 & ~n52876 ;
  assign n52878 = ~\pi0209  & n52877 ;
  assign n52879 = \pi0219  & ~n52634 ;
  assign n52880 = ~\pi0211  & ~n51630 ;
  assign n52881 = ~n52571 & n52880 ;
  assign n52882 = ~n52570 & n52881 ;
  assign n52883 = ~\pi1145  & n52000 ;
  assign n52884 = \pi0211  & n52556 ;
  assign n52885 = n50924 & ~n52521 ;
  assign n52886 = ~n52884 & ~n52885 ;
  assign n52887 = ~n50570 & n52886 ;
  assign n52888 = ~n52883 & n52887 ;
  assign n52889 = ~n52882 & n52888 ;
  assign n52890 = n52879 & ~n52889 ;
  assign n52891 = n9948 & ~n52890 ;
  assign n52892 = ~n52571 & n52838 ;
  assign n52893 = ~n52570 & n52892 ;
  assign n52894 = ~\pi0214  & ~n52858 ;
  assign n52895 = n50693 & n52818 ;
  assign n52896 = \pi0212  & ~n52895 ;
  assign n52897 = ~n52894 & n52896 ;
  assign n52898 = ~n52893 & n52897 ;
  assign n52899 = n52864 & ~n52898 ;
  assign n52900 = ~\pi0209  & ~n52899 ;
  assign n52901 = n52891 & n52900 ;
  assign n52902 = ~n52878 & ~n52901 ;
  assign n52903 = n52873 & ~n52902 ;
  assign n52904 = n50689 & n51630 ;
  assign n52905 = n52710 & n52904 ;
  assign n52906 = ~n52815 & ~n52821 ;
  assign n52907 = ~n52819 & n52906 ;
  assign n52908 = \pi0299  & n46750 ;
  assign n52909 = n6848 & n52908 ;
  assign n52910 = ~n52907 & n52909 ;
  assign n52911 = ~n52905 & ~n52910 ;
  assign n52912 = ~n52877 & n52911 ;
  assign n52913 = ~\pi1149  & ~n52912 ;
  assign n52914 = ~\pi1148  & ~n52829 ;
  assign n52915 = n51975 & ~n52837 ;
  assign n52916 = n12255 & ~n52915 ;
  assign n52917 = ~\pi1146  & n52001 ;
  assign n52918 = n50679 & ~n52917 ;
  assign n52919 = ~n52916 & ~n52918 ;
  assign n52920 = ~\pi0211  & n51630 ;
  assign n52921 = n51108 & n52920 ;
  assign n52922 = ~n50948 & n52707 ;
  assign n52923 = ~n52921 & ~n52922 ;
  assign n52924 = n52919 & n52923 ;
  assign n52925 = ~n50701 & ~n52921 ;
  assign n52926 = ~n52707 & n52925 ;
  assign n52927 = n9948 & ~n52926 ;
  assign n52928 = ~\pi1148  & n52927 ;
  assign n52929 = ~n52924 & n52928 ;
  assign n52930 = ~n52914 & ~n52929 ;
  assign n52931 = n52913 & ~n52930 ;
  assign n52932 = \pi1148  & ~n52829 ;
  assign n52933 = n51975 & ~n52846 ;
  assign n52934 = n50679 & ~n52933 ;
  assign n52935 = n50570 & ~n51975 ;
  assign n52936 = ~\pi0219  & ~n52935 ;
  assign n52937 = ~n52916 & n52936 ;
  assign n52938 = ~n52934 & n52937 ;
  assign n52939 = \pi0219  & ~n52920 ;
  assign n52940 = n52710 & ~n52939 ;
  assign n52941 = ~n52709 & ~n52940 ;
  assign n52942 = \pi1148  & ~n52941 ;
  assign n52943 = ~n52938 & n52942 ;
  assign n52944 = ~n52932 & ~n52943 ;
  assign n52945 = n9948 & n52741 ;
  assign n52946 = n52912 & ~n52945 ;
  assign n52947 = ~\pi1149  & ~n52946 ;
  assign n52948 = ~n52944 & n52947 ;
  assign n52949 = ~n52931 & ~n52948 ;
  assign n52950 = \pi0209  & ~n52949 ;
  assign n52951 = n51972 & ~n52059 ;
  assign n52952 = ~n52058 & n52951 ;
  assign n52953 = ~n51679 & ~n52535 ;
  assign n52954 = n50430 & n52953 ;
  assign n52955 = ~n52952 & n52954 ;
  assign n52956 = n50967 & ~n52063 ;
  assign n52957 = ~n52061 & n52956 ;
  assign n52958 = ~n52955 & ~n52957 ;
  assign n52959 = n52671 & n52958 ;
  assign n52960 = ~\pi0219  & ~n52959 ;
  assign n52961 = \pi0214  & ~n51679 ;
  assign n52962 = ~n52837 & n52961 ;
  assign n52963 = ~n52952 & n52962 ;
  assign n52964 = \pi0212  & ~n52963 ;
  assign n52965 = n50863 & n52953 ;
  assign n52966 = ~n52952 & n52965 ;
  assign n52967 = n50442 & ~n52063 ;
  assign n52968 = ~n52061 & n52967 ;
  assign n52969 = ~n52966 & ~n52968 ;
  assign n52970 = n52964 & n52969 ;
  assign n52971 = n52829 & ~n52970 ;
  assign n52972 = n52960 & n52971 ;
  assign n52973 = ~n52681 & n52912 ;
  assign n52974 = \pi0219  & n52033 ;
  assign n52975 = n9948 & ~n52974 ;
  assign n52976 = n52828 & ~n52940 ;
  assign n52977 = ~n52826 & n52976 ;
  assign n52978 = ~n52975 & n52977 ;
  assign n52979 = ~n52973 & ~n52978 ;
  assign n52980 = ~n52972 & n52979 ;
  assign n52981 = ~\pi1148  & ~n52980 ;
  assign n52982 = n50571 & ~n52782 ;
  assign n52983 = ~n50571 & n51918 ;
  assign n52984 = \pi0219  & ~n52983 ;
  assign n52985 = ~n52982 & n52984 ;
  assign n52986 = ~\pi0057  & n13550 ;
  assign n52987 = n6848 & n52986 ;
  assign n52988 = ~n52985 & n52987 ;
  assign n52989 = ~n52940 & ~n52988 ;
  assign n52990 = ~\pi0214  & n52814 ;
  assign n52991 = \pi0214  & ~n52818 ;
  assign n52992 = ~n51918 & ~n52991 ;
  assign n52993 = ~n52990 & n52992 ;
  assign n52994 = n52783 & ~n52993 ;
  assign n52995 = ~\pi0212  & n51918 ;
  assign n52996 = n50556 & n52854 ;
  assign n52997 = ~\pi0219  & ~n52996 ;
  assign n52998 = ~n52995 & n52997 ;
  assign n52999 = ~n52994 & n52998 ;
  assign n53000 = ~n52989 & ~n52999 ;
  assign n53001 = \pi1148  & ~n52877 ;
  assign n53002 = ~n53000 & n53001 ;
  assign n53003 = \pi0219  & ~n52798 ;
  assign n53004 = n9948 & ~n53003 ;
  assign n53005 = ~\pi0299  & n50876 ;
  assign n53006 = ~n50840 & ~n53005 ;
  assign n53007 = \pi0212  & \pi0299  ;
  assign n53008 = ~n50442 & n53007 ;
  assign n53009 = \pi0212  & ~n53008 ;
  assign n53010 = n53006 & n53009 ;
  assign n53011 = ~\pi0212  & ~n50876 ;
  assign n53012 = n50824 & n53011 ;
  assign n53013 = ~\pi0211  & ~\pi0212  ;
  assign n53014 = n50693 & n53013 ;
  assign n53015 = ~\pi0219  & ~n53014 ;
  assign n53016 = ~n53012 & n53015 ;
  assign n53017 = ~n53010 & n53016 ;
  assign n53018 = n53004 & ~n53017 ;
  assign n53019 = \pi1148  & ~n53018 ;
  assign n53020 = n52829 & n53019 ;
  assign n53021 = n52911 & n53020 ;
  assign n53022 = \pi0209  & \pi1149  ;
  assign n53023 = ~n53021 & n53022 ;
  assign n53024 = ~n53002 & n53023 ;
  assign n53025 = ~n52981 & n53024 ;
  assign n53026 = ~\pi0213  & ~n53025 ;
  assign n53027 = ~n52950 & n53026 ;
  assign n53028 = ~n52903 & n53027 ;
  assign n53029 = \pi0230  & n53028 ;
  assign n53030 = ~\pi0230  & ~\pi0240  ;
  assign n53031 = ~n53029 & ~n53030 ;
  assign n53032 = ~n52813 & n53031 ;
  assign n53033 = \pi0219  & ~n52007 ;
  assign n53034 = n9948 & ~n53033 ;
  assign n53035 = n52167 & ~n53034 ;
  assign n53036 = n52167 & ~n52301 ;
  assign n53037 = n52299 & n53036 ;
  assign n53038 = ~n53035 & ~n53037 ;
  assign n53039 = n12577 & n51187 ;
  assign n53040 = n50679 & n53039 ;
  assign n53041 = ~\pi1151  & ~n53040 ;
  assign n53042 = ~n52210 & n53041 ;
  assign n53043 = ~\pi1152  & ~n53042 ;
  assign n53044 = ~\pi1150  & n53043 ;
  assign n53045 = n53038 & n53044 ;
  assign n53046 = ~\pi1149  & n53045 ;
  assign n53047 = n52299 & ~n52301 ;
  assign n53048 = n53034 & ~n53047 ;
  assign n53049 = ~\pi0212  & \pi0299  ;
  assign n53050 = ~\pi0212  & n12691 ;
  assign n53051 = n50877 & n53050 ;
  assign n53052 = ~n53049 & ~n53051 ;
  assign n53053 = ~n52292 & ~n53052 ;
  assign n53054 = ~n52000 & n53053 ;
  assign n53055 = n50442 & ~n52005 ;
  assign n53056 = \pi0212  & n12691 ;
  assign n53057 = n50877 & n53056 ;
  assign n53058 = ~n53007 & ~n53057 ;
  assign n53059 = ~n53055 & ~n53058 ;
  assign n53060 = ~\pi0219  & ~n53059 ;
  assign n53061 = ~n53054 & n53060 ;
  assign n53062 = n53034 & ~n53061 ;
  assign n53063 = n52235 & ~n53062 ;
  assign n53064 = ~n53048 & n53063 ;
  assign n53065 = ~n50570 & n50701 ;
  assign n53066 = ~n12256 & n53065 ;
  assign n53067 = ~n52231 & n53066 ;
  assign n53068 = ~\pi1151  & ~n53067 ;
  assign n53069 = ~n52232 & n53068 ;
  assign n53070 = ~\pi1150  & \pi1152  ;
  assign n53071 = ~n53069 & n53070 ;
  assign n53072 = ~\pi1149  & n53071 ;
  assign n53073 = ~n53064 & n53072 ;
  assign n53074 = ~n53046 & ~n53073 ;
  assign n53075 = n52346 & ~n52743 ;
  assign n53076 = ~\pi0214  & n52741 ;
  assign n53077 = ~\pi0212  & ~n53076 ;
  assign n53078 = n50978 & n52750 ;
  assign n53079 = n53077 & ~n53078 ;
  assign n53080 = \pi0214  & n52753 ;
  assign n53081 = n52750 & n53080 ;
  assign n53082 = \pi0212  & ~n53081 ;
  assign n53083 = ~\pi0214  & ~n50977 ;
  assign n53084 = n52750 & n53083 ;
  assign n53085 = n53082 & ~n53084 ;
  assign n53086 = ~n53079 & ~n53085 ;
  assign n53087 = ~\pi0219  & n52346 ;
  assign n53088 = ~n53086 & n53087 ;
  assign n53089 = ~n53075 & ~n53088 ;
  assign n53090 = n9948 & ~n52985 ;
  assign n53091 = \pi0211  & ~n52782 ;
  assign n53092 = ~\pi0211  & ~n50586 ;
  assign n53093 = ~n13558 & n50411 ;
  assign n53094 = n51947 & ~n53093 ;
  assign n53095 = n53092 & ~n53094 ;
  assign n53096 = ~n53091 & ~n53095 ;
  assign n53097 = ~\pi0214  & n53096 ;
  assign n53098 = n52783 & ~n53097 ;
  assign n53099 = ~n51918 & n52661 ;
  assign n53100 = ~n52660 & ~n53099 ;
  assign n53101 = n50954 & n53096 ;
  assign n53102 = n53100 & ~n53101 ;
  assign n53103 = ~n53098 & ~n53102 ;
  assign n53104 = n53090 & ~n53103 ;
  assign n53105 = n52235 & ~n53104 ;
  assign n53106 = n53089 & ~n53105 ;
  assign n53107 = \pi1152  & ~n53106 ;
  assign n53108 = \pi0212  & n51918 ;
  assign n53109 = n52546 & ~n52782 ;
  assign n53110 = ~n53108 & ~n53109 ;
  assign n53111 = ~n53096 & ~n53110 ;
  assign n53112 = ~\pi0219  & ~n52785 ;
  assign n53113 = ~n53095 & n53112 ;
  assign n53114 = n53100 & ~n53113 ;
  assign n53115 = ~n53111 & ~n53114 ;
  assign n53116 = n53090 & ~n53115 ;
  assign n53117 = \pi1151  & ~\pi1152  ;
  assign n53118 = ~n52166 & n53117 ;
  assign n53119 = ~n53116 & n53118 ;
  assign n53120 = ~\pi1151  & ~n9948 ;
  assign n53121 = ~n52210 & n53120 ;
  assign n53122 = ~\pi1152  & n53121 ;
  assign n53123 = n52212 & n52753 ;
  assign n53124 = ~n50977 & n53123 ;
  assign n53125 = n52750 & n53124 ;
  assign n53126 = ~n52212 & n52741 ;
  assign n53127 = ~n53125 & ~n53126 ;
  assign n53128 = ~\pi1152  & n52211 ;
  assign n53129 = n53127 & n53128 ;
  assign n53130 = ~n53122 & ~n53129 ;
  assign n53131 = ~\pi1149  & n53130 ;
  assign n53132 = ~n53119 & n53131 ;
  assign n53133 = \pi1150  & n53132 ;
  assign n53134 = ~n53107 & n53133 ;
  assign n53135 = n53074 & ~n53134 ;
  assign n53136 = n52167 & ~n52676 ;
  assign n53137 = ~\pi0219  & \pi1151  ;
  assign n53138 = ~n52166 & n53137 ;
  assign n53139 = \pi0212  & ~n52658 ;
  assign n53140 = ~n52671 & ~n53139 ;
  assign n53141 = \pi0211  & ~n52033 ;
  assign n53142 = ~n52654 & n53092 ;
  assign n53143 = ~n53141 & ~n53142 ;
  assign n53144 = ~n52659 & n53143 ;
  assign n53145 = ~n53140 & ~n53144 ;
  assign n53146 = n53138 & ~n53145 ;
  assign n53147 = ~n53136 & ~n53146 ;
  assign n53148 = ~\pi1152  & ~n52211 ;
  assign n53149 = ~\pi0211  & n50701 ;
  assign n53150 = n50679 & n53149 ;
  assign n53151 = ~n52707 & ~n53150 ;
  assign n53152 = n9948 & ~n50977 ;
  assign n53153 = ~\pi1152  & n53152 ;
  assign n53154 = ~n53151 & n53153 ;
  assign n53155 = ~n53148 & ~n53154 ;
  assign n53156 = n53147 & ~n53155 ;
  assign n53157 = \pi1152  & ~n52346 ;
  assign n53158 = ~n12256 & ~n52231 ;
  assign n53159 = ~\pi0219  & ~n51585 ;
  assign n53160 = ~n53158 & n53159 ;
  assign n53161 = n52707 & ~n53160 ;
  assign n53162 = ~\pi0219  & n52616 ;
  assign n53163 = ~n53160 & n53162 ;
  assign n53164 = ~n53161 & ~n53163 ;
  assign n53165 = \pi1152  & n27408 ;
  assign n53166 = ~n53164 & n53165 ;
  assign n53167 = ~n53157 & ~n53166 ;
  assign n53168 = ~\pi1150  & n53167 ;
  assign n53169 = n50430 & ~n52654 ;
  assign n53170 = ~n50430 & ~n52033 ;
  assign n53171 = ~n53169 & ~n53170 ;
  assign n53172 = ~\pi0219  & ~n53008 ;
  assign n53173 = n53171 & n53172 ;
  assign n53174 = ~n52288 & n53173 ;
  assign n53175 = n52676 & ~n53174 ;
  assign n53176 = ~\pi1150  & n52235 ;
  assign n53177 = ~n53175 & n53176 ;
  assign n53178 = ~n53168 & ~n53177 ;
  assign n53179 = ~n53156 & ~n53178 ;
  assign n53180 = ~\pi0219  & ~\pi1153  ;
  assign n53181 = ~n53008 & n53180 ;
  assign n53182 = ~n52798 & n53181 ;
  assign n53183 = n50430 & n53007 ;
  assign n53184 = ~\pi0219  & ~n53183 ;
  assign n53185 = ~n52711 & ~n53184 ;
  assign n53186 = n52710 & n53185 ;
  assign n53187 = ~n53018 & ~n53186 ;
  assign n53188 = ~n53182 & ~n53187 ;
  assign n53189 = \pi1150  & \pi1151  ;
  assign n53190 = ~n52166 & n53189 ;
  assign n53191 = ~n53188 & n53190 ;
  assign n53192 = ~\pi1152  & n9948 ;
  assign n53193 = ~n51975 & n53192 ;
  assign n53194 = ~n53117 & ~n53193 ;
  assign n53195 = \pi1150  & ~n53043 ;
  assign n53196 = n53194 & n53195 ;
  assign n53197 = \pi1149  & ~n53196 ;
  assign n53198 = ~n53191 & n53197 ;
  assign n53199 = n12577 & ~n53008 ;
  assign n53200 = ~n52798 & n53199 ;
  assign n53201 = ~n52800 & ~n53200 ;
  assign n53202 = n52235 & ~n53201 ;
  assign n53203 = ~n53188 & n53202 ;
  assign n53204 = \pi1152  & ~n53203 ;
  assign n53205 = n51975 & ~n52000 ;
  assign n53206 = n12255 & ~n53205 ;
  assign n53207 = n52936 & ~n53206 ;
  assign n53208 = ~\pi0299  & n51975 ;
  assign n53209 = n50679 & ~n50977 ;
  assign n53210 = ~n53208 & n53209 ;
  assign n53211 = n52346 & ~n53210 ;
  assign n53212 = n53207 & n53211 ;
  assign n53213 = n9948 & ~n51998 ;
  assign n53214 = n52346 & ~n53213 ;
  assign n53215 = \pi1149  & ~n53214 ;
  assign n53216 = ~n53212 & n53215 ;
  assign n53217 = n53204 & n53216 ;
  assign n53218 = ~n53198 & ~n53217 ;
  assign n53219 = ~n53179 & ~n53218 ;
  assign n53220 = n53135 & ~n53219 ;
  assign n53221 = ~\pi0209  & ~n53220 ;
  assign n53222 = ~n52317 & ~n52319 ;
  assign n53223 = \pi0209  & ~\pi1152  ;
  assign n53224 = ~n53222 & n53223 ;
  assign n53225 = \pi0209  & \pi1152  ;
  assign n53226 = n52372 & n53225 ;
  assign n53227 = n52811 & ~n53226 ;
  assign n53228 = ~n53224 & n53227 ;
  assign n53229 = ~n53221 & n53228 ;
  assign n53230 = \pi1151  & ~n52229 ;
  assign n53231 = ~n50430 & n51990 ;
  assign n53232 = \pi0208  & ~n50430 ;
  assign n53233 = ~n51988 & n53232 ;
  assign n53234 = ~n53231 & ~n53233 ;
  assign n53235 = n51975 & ~n51984 ;
  assign n53236 = \pi0214  & ~n53235 ;
  assign n53237 = n53234 & ~n53236 ;
  assign n53238 = \pi0212  & ~n53237 ;
  assign n53239 = ~n52333 & n52342 ;
  assign n53240 = ~\pi0219  & \pi1152  ;
  assign n53241 = ~n53239 & n53240 ;
  assign n53242 = ~n53238 & n53241 ;
  assign n53243 = n27408 & ~n52367 ;
  assign n53244 = ~n53242 & n53243 ;
  assign n53245 = \pi0219  & ~\pi1152  ;
  assign n53246 = n52033 & n53245 ;
  assign n53247 = ~\pi0299  & n51219 ;
  assign n53248 = ~\pi0299  & ~n52063 ;
  assign n53249 = ~n52061 & n53248 ;
  assign n53250 = ~n53247 & ~n53249 ;
  assign n53251 = ~\pi0214  & ~n52063 ;
  assign n53252 = ~n52061 & n53251 ;
  assign n53253 = \pi0212  & ~n53252 ;
  assign n53254 = n53250 & n53253 ;
  assign n53255 = ~n52672 & n53254 ;
  assign n53256 = ~n52036 & n53250 ;
  assign n53257 = n51174 & ~n53256 ;
  assign n53258 = ~n53255 & n53257 ;
  assign n53259 = ~n53246 & ~n53258 ;
  assign n53260 = n53244 & n53259 ;
  assign n53261 = n53230 & ~n53260 ;
  assign n53262 = ~n51984 & n52725 ;
  assign n53263 = ~n52294 & n53262 ;
  assign n53264 = ~n52347 & n53263 ;
  assign n53265 = ~\pi0219  & ~n53054 ;
  assign n53266 = \pi0214  & ~n52000 ;
  assign n53267 = ~n52003 & n53266 ;
  assign n53268 = n53059 & ~n53267 ;
  assign n53269 = ~n52347 & ~n53268 ;
  assign n53270 = n53265 & n53269 ;
  assign n53271 = ~n53264 & ~n53270 ;
  assign n53272 = \pi1152  & n9948 ;
  assign n53273 = ~n52348 & n53272 ;
  assign n53274 = n53271 & n53273 ;
  assign n53275 = ~\pi1151  & ~n52631 ;
  assign n53276 = n53265 & ~n53268 ;
  assign n53277 = n9948 & ~n52366 ;
  assign n53278 = ~\pi1152  & n53277 ;
  assign n53279 = ~n53263 & n53278 ;
  assign n53280 = ~n53276 & n53279 ;
  assign n53281 = n53275 & ~n53280 ;
  assign n53282 = ~n53274 & n53281 ;
  assign n53283 = ~\pi1149  & ~n53282 ;
  assign n53284 = ~n53261 & n53283 ;
  assign n53285 = ~\pi1151  & ~n52641 ;
  assign n53286 = ~n52712 & ~n53277 ;
  assign n53287 = ~n52349 & n53286 ;
  assign n53288 = \pi1152  & n53287 ;
  assign n53289 = \pi0208  & ~n51934 ;
  assign n53290 = n12255 & ~n50411 ;
  assign n53291 = ~\pi0299  & n12255 ;
  assign n53292 = ~n51014 & n53291 ;
  assign n53293 = ~n53290 & ~n53292 ;
  assign n53294 = ~n53289 & ~n53293 ;
  assign n53295 = ~n52006 & ~n52291 ;
  assign n53296 = ~n12255 & ~n52347 ;
  assign n53297 = ~n53295 & n53296 ;
  assign n53298 = ~n53294 & ~n53297 ;
  assign n53299 = n53240 & ~n53298 ;
  assign n53300 = ~n53288 & ~n53299 ;
  assign n53301 = ~n53263 & n53277 ;
  assign n53302 = ~n53276 & n53301 ;
  assign n53303 = n51985 & ~n52294 ;
  assign n53304 = ~n53286 & ~n53303 ;
  assign n53305 = ~\pi1152  & ~n53304 ;
  assign n53306 = ~n53302 & n53305 ;
  assign n53307 = n53300 & ~n53306 ;
  assign n53308 = n53285 & ~n53307 ;
  assign n53309 = n50998 & ~n52368 ;
  assign n53310 = \pi0208  & \pi0212  ;
  assign n53311 = ~n51988 & n53310 ;
  assign n53312 = \pi0212  & n50411 ;
  assign n53313 = ~n51043 & n53312 ;
  assign n53314 = ~\pi0219  & ~n53313 ;
  assign n53315 = ~n53311 & n53314 ;
  assign n53316 = ~n53239 & n53315 ;
  assign n53317 = n53309 & ~n53316 ;
  assign n53318 = \pi1151  & ~n52621 ;
  assign n53319 = n51088 & ~n52313 ;
  assign n53320 = ~n52287 & n53250 ;
  assign n53321 = ~\pi0219  & ~n53320 ;
  assign n53322 = n53319 & ~n53321 ;
  assign n53323 = n53318 & ~n53322 ;
  assign n53324 = ~n53317 & n53323 ;
  assign n53325 = \pi1149  & ~n53324 ;
  assign n53326 = ~n53308 & n53325 ;
  assign n53327 = \pi1150  & ~n53326 ;
  assign n53328 = ~n53284 & n53327 ;
  assign n53329 = n51819 & n52312 ;
  assign n53330 = ~\pi0214  & ~n52310 ;
  assign n53331 = ~\pi0214  & ~n51007 ;
  assign n53332 = ~n52033 & n53331 ;
  assign n53333 = ~n53330 & ~n53332 ;
  assign n53334 = ~\pi0219  & n53333 ;
  assign n53335 = n52283 & n53334 ;
  assign n53336 = ~n53329 & ~n53335 ;
  assign n53337 = n53319 & n53336 ;
  assign n53338 = \pi1151  & ~n52513 ;
  assign n53339 = ~n51991 & ~n52547 ;
  assign n53340 = n51986 & ~n53339 ;
  assign n53341 = n53309 & ~n53340 ;
  assign n53342 = n53338 & ~n53341 ;
  assign n53343 = ~n53337 & n53342 ;
  assign n53344 = ~\pi1151  & ~n52233 ;
  assign n53345 = \pi1152  & ~n52347 ;
  assign n53346 = ~\pi0219  & n53345 ;
  assign n53347 = ~n52294 & n53346 ;
  assign n53348 = ~n53287 & ~n53347 ;
  assign n53349 = n53344 & ~n53348 ;
  assign n53350 = ~\pi1151  & ~\pi1152  ;
  assign n53351 = ~n52233 & n53350 ;
  assign n53352 = ~n53304 & n53351 ;
  assign n53353 = ~n53349 & ~n53352 ;
  assign n53354 = \pi1149  & n53353 ;
  assign n53355 = ~n53343 & n53354 ;
  assign n53356 = \pi1149  & ~\pi1150  ;
  assign n53357 = n51990 & n52572 ;
  assign n53358 = \pi0208  & n52572 ;
  assign n53359 = ~n51988 & n53358 ;
  assign n53360 = ~n53357 & ~n53359 ;
  assign n53361 = n53235 & n53360 ;
  assign n53362 = ~n9948 & ~n52572 ;
  assign n53363 = n52250 & ~n53362 ;
  assign n53364 = ~n53361 & n53363 ;
  assign n53365 = \pi1151  & ~n53362 ;
  assign n53366 = ~\pi1152  & ~n51007 ;
  assign n53367 = ~n52033 & n53366 ;
  assign n53368 = ~\pi0211  & ~\pi1152  ;
  assign n53369 = n50701 & n53368 ;
  assign n53370 = n50679 & n53369 ;
  assign n53371 = n9948 & ~n53370 ;
  assign n53372 = ~n53367 & n53371 ;
  assign n53373 = n53365 & ~n53372 ;
  assign n53374 = ~\pi1152  & n51984 ;
  assign n53375 = \pi1152  & ~n51919 ;
  assign n53376 = n51918 & n53375 ;
  assign n53377 = ~n53374 & ~n53376 ;
  assign n53378 = n51966 & ~n53377 ;
  assign n53379 = ~\pi1150  & ~n53378 ;
  assign n53380 = ~n53373 & n53379 ;
  assign n53381 = ~n53364 & n53380 ;
  assign n53382 = ~n53356 & ~n53381 ;
  assign n53383 = ~n53355 & ~n53382 ;
  assign n53384 = \pi0209  & ~n53383 ;
  assign n53385 = ~n53328 & n53384 ;
  assign n53386 = ~n52743 & n53275 ;
  assign n53387 = ~n52768 & n53275 ;
  assign n53388 = ~n52765 & n53387 ;
  assign n53389 = ~n53386 & ~n53388 ;
  assign n53390 = \pi1150  & ~n53230 ;
  assign n53391 = n9948 & ~n52304 ;
  assign n53392 = ~n52790 & ~n53391 ;
  assign n53393 = \pi1150  & ~n53392 ;
  assign n53394 = ~n52789 & n53393 ;
  assign n53395 = ~n53390 & ~n53394 ;
  assign n53396 = n53389 & ~n53395 ;
  assign n53397 = ~\pi1150  & \pi1151  ;
  assign n53398 = ~n52683 & n53397 ;
  assign n53399 = ~\pi1149  & ~n53398 ;
  assign n53400 = ~n53396 & n53399 ;
  assign n53401 = ~n52734 & n53285 ;
  assign n53402 = ~n52709 & n53401 ;
  assign n53403 = n52800 & n53318 ;
  assign n53404 = \pi1150  & ~n53403 ;
  assign n53405 = ~n53402 & n53404 ;
  assign n53406 = \pi1149  & ~n53405 ;
  assign n53407 = n53338 & n53406 ;
  assign n53408 = ~n52677 & n53407 ;
  assign n53409 = ~\pi1150  & ~n52727 ;
  assign n53410 = ~n52724 & n53409 ;
  assign n53411 = n52715 & n53410 ;
  assign n53412 = ~\pi1150  & ~n12257 ;
  assign n53413 = n50677 & n53412 ;
  assign n53414 = ~n53397 & ~n53413 ;
  assign n53415 = \pi1149  & n53414 ;
  assign n53416 = ~n53405 & n53415 ;
  assign n53417 = ~n53411 & n53416 ;
  assign n53418 = ~\pi0209  & ~n53417 ;
  assign n53419 = ~n53408 & n53418 ;
  assign n53420 = ~n53400 & n53419 ;
  assign n53421 = ~\pi0213  & \pi0230  ;
  assign n53422 = ~n53420 & n53421 ;
  assign n53423 = ~n53385 & n53422 ;
  assign n53424 = ~\pi0230  & ~\pi0241  ;
  assign n53425 = ~n53423 & ~n53424 ;
  assign n53426 = ~n53229 & n53425 ;
  assign n53427 = \pi0199  & \pi1144  ;
  assign n53428 = ~\pi0200  & ~n53427 ;
  assign n53429 = ~n51721 & n53428 ;
  assign n53430 = ~\pi0299  & n12409 ;
  assign n53431 = ~n51723 & n53430 ;
  assign n53432 = ~n53429 & n53431 ;
  assign n53433 = ~n52515 & n53428 ;
  assign n53434 = ~\pi0299  & n50381 ;
  assign n53435 = ~n52519 & n53434 ;
  assign n53436 = ~n53433 & n53435 ;
  assign n53437 = ~n53432 & ~n53436 ;
  assign n53438 = ~\pi0299  & n50418 ;
  assign n53439 = ~n52519 & n53438 ;
  assign n53440 = ~n53433 & n53439 ;
  assign n53441 = \pi0211  & ~n51630 ;
  assign n53442 = ~n53440 & n53441 ;
  assign n53443 = n53437 & n53442 ;
  assign n53444 = ~\pi0211  & ~n52535 ;
  assign n53445 = ~n53440 & n53444 ;
  assign n53446 = n53437 & n53445 ;
  assign n53447 = ~n53443 & ~n53446 ;
  assign n53448 = ~\pi0214  & ~n53447 ;
  assign n53449 = ~n51630 & ~n53440 ;
  assign n53450 = n53437 & n53449 ;
  assign n53451 = n50967 & n53450 ;
  assign n53452 = ~n50783 & ~n53440 ;
  assign n53453 = n53437 & n53452 ;
  assign n53454 = n50430 & n53453 ;
  assign n53455 = ~n53451 & ~n53454 ;
  assign n53456 = ~n53448 & n53455 ;
  assign n53457 = \pi0212  & n53456 ;
  assign n53458 = n50600 & ~n52818 ;
  assign n53459 = n12255 & ~n51667 ;
  assign n53460 = ~n53458 & ~n53459 ;
  assign n53461 = n50556 & ~n52818 ;
  assign n53462 = ~\pi0219  & ~n53461 ;
  assign n53463 = n53460 & n53462 ;
  assign n53464 = \pi0219  & ~n50658 ;
  assign n53465 = n50677 & ~n53464 ;
  assign n53466 = ~n53463 & n53465 ;
  assign n53467 = \pi0213  & ~n53466 ;
  assign n53468 = ~\pi0299  & ~n52519 ;
  assign n53469 = ~n53433 & n53468 ;
  assign n53470 = n50877 & n53469 ;
  assign n53471 = ~\pi0214  & ~n53470 ;
  assign n53472 = ~\pi0219  & n53437 ;
  assign n53473 = n53471 & n53472 ;
  assign n53474 = ~n52660 & ~n53473 ;
  assign n53475 = n50954 & ~n53447 ;
  assign n53476 = n53474 & ~n53475 ;
  assign n53477 = n53467 & ~n53476 ;
  assign n53478 = ~n53457 & n53477 ;
  assign n53479 = n50571 & ~n53453 ;
  assign n53480 = n9948 & n53479 ;
  assign n53481 = \pi0219  & ~n53470 ;
  assign n53482 = n53437 & n53481 ;
  assign n53483 = n9948 & ~n51730 ;
  assign n53484 = ~n53482 & n53483 ;
  assign n53485 = ~n53480 & ~n53484 ;
  assign n53486 = n53467 & n53485 ;
  assign n53487 = \pi0299  & ~n50666 ;
  assign n53488 = n50948 & ~n53440 ;
  assign n53489 = ~n53487 & n53488 ;
  assign n53490 = n50570 & ~n53470 ;
  assign n53491 = ~n53489 & ~n53490 ;
  assign n53492 = \pi0299  & \pi1142  ;
  assign n53493 = n51730 & ~n53492 ;
  assign n53494 = ~n53440 & n53493 ;
  assign n53495 = n50713 & ~n53470 ;
  assign n53496 = ~n53494 & ~n53495 ;
  assign n53497 = n53491 & n53496 ;
  assign n53498 = ~\pi0213  & ~n50677 ;
  assign n53499 = ~\pi0213  & \pi0219  ;
  assign n53500 = ~\pi0213  & ~n50662 ;
  assign n53501 = ~n50680 & n53500 ;
  assign n53502 = ~n53499 & ~n53501 ;
  assign n53503 = n50684 & ~n53502 ;
  assign n53504 = ~n53498 & ~n53503 ;
  assign n53505 = n53437 & ~n53504 ;
  assign n53506 = ~n53497 & n53505 ;
  assign n53507 = ~n9948 & n53498 ;
  assign n53508 = ~n9948 & n50684 ;
  assign n53509 = ~n53502 & n53508 ;
  assign n53510 = ~n53507 & ~n53509 ;
  assign n53511 = \pi0209  & \pi0230  ;
  assign n53512 = n53510 & n53511 ;
  assign n53513 = ~n53506 & n53512 ;
  assign n53514 = ~n53486 & n53513 ;
  assign n53515 = ~n53478 & n53514 ;
  assign n53516 = ~n50570 & n50658 ;
  assign n53517 = \pi0219  & ~n53516 ;
  assign n53518 = \pi0299  & ~n53517 ;
  assign n53519 = n9948 & n53518 ;
  assign n53520 = ~n53463 & n53519 ;
  assign n53521 = n53467 & ~n53520 ;
  assign n53522 = ~n50656 & n53521 ;
  assign n53523 = ~\pi0209  & ~n53522 ;
  assign n53524 = ~\pi0213  & n50684 ;
  assign n53525 = ~n50682 & n53524 ;
  assign n53526 = ~n53498 & ~n53525 ;
  assign n53527 = n50675 & ~n53526 ;
  assign n53528 = \pi0230  & ~n53527 ;
  assign n53529 = n53523 & n53528 ;
  assign n53530 = ~\pi0230  & \pi0242  ;
  assign n53531 = ~n53529 & ~n53530 ;
  assign n53532 = ~n53515 & n53531 ;
  assign n53533 = ~\pi0083  & ~\pi0085  ;
  assign n53534 = ~\pi0081  & n53533 ;
  assign n53535 = \pi0314  & \pi0802  ;
  assign n53536 = \pi0276  & ~\pi1091  ;
  assign n53537 = n53535 & n53536 ;
  assign n53538 = ~n53534 & n53537 ;
  assign n53539 = \pi0276  & n53535 ;
  assign n53540 = ~n53534 & n53539 ;
  assign n53541 = \pi0271  & ~\pi1091  ;
  assign n53542 = \pi0273  & n53541 ;
  assign n53543 = n53540 & n53542 ;
  assign n53544 = ~\pi0199  & n53543 ;
  assign n53545 = ~n53533 & n53535 ;
  assign n53546 = ~\pi1091  & ~n53545 ;
  assign n53547 = ~\pi0276  & ~\pi1091  ;
  assign n53548 = ~\pi0271  & ~\pi1091  ;
  assign n53549 = ~n53547 & ~n53548 ;
  assign n53550 = \pi0273  & n53549 ;
  assign n53551 = ~n53546 & n53550 ;
  assign n53552 = ~\pi1091  & ~n53551 ;
  assign n53553 = ~n53544 & n53552 ;
  assign n53554 = n53538 & ~n53553 ;
  assign n53555 = ~n53543 & ~n53551 ;
  assign n53556 = ~\pi1091  & n53555 ;
  assign n53557 = ~\pi0199  & ~n53556 ;
  assign n53558 = \pi0276  & n53545 ;
  assign n53559 = ~\pi1091  & ~n53558 ;
  assign n53560 = ~\pi0273  & ~\pi1091  ;
  assign n53561 = ~n53548 & ~n53560 ;
  assign n53562 = ~\pi0200  & n53561 ;
  assign n53563 = ~n53559 & n53562 ;
  assign n53564 = ~\pi0299  & ~n53563 ;
  assign n53565 = ~n53557 & n53564 ;
  assign n53566 = ~n53554 & n53565 ;
  assign n53567 = ~n53559 & n53561 ;
  assign n53568 = \pi0299  & ~n53543 ;
  assign n53569 = ~n53567 & n53568 ;
  assign n53570 = \pi1155  & ~n53569 ;
  assign n53571 = ~n53566 & n53570 ;
  assign n53572 = \pi0199  & n53561 ;
  assign n53573 = ~n53559 & n53572 ;
  assign n53574 = n53564 & ~n53573 ;
  assign n53575 = ~n53554 & n53574 ;
  assign n53576 = \pi0299  & n53542 ;
  assign n53577 = n53540 & n53576 ;
  assign n53578 = ~\pi0200  & ~n53538 ;
  assign n53579 = ~n53568 & ~n53578 ;
  assign n53580 = ~n53553 & n53579 ;
  assign n53581 = ~n53577 & ~n53580 ;
  assign n53582 = ~\pi0243  & ~n53581 ;
  assign n53583 = ~n53575 & n53582 ;
  assign n53584 = n53571 & ~n53583 ;
  assign n53585 = ~n53553 & ~n53578 ;
  assign n53586 = ~\pi0299  & ~n53573 ;
  assign n53587 = ~n53585 & n53586 ;
  assign n53588 = \pi0273  & \pi0276  ;
  assign n53589 = n53541 & n53588 ;
  assign n53590 = n53545 & n53589 ;
  assign n53591 = \pi0299  & ~n53590 ;
  assign n53592 = ~n53587 & ~n53591 ;
  assign n53593 = ~n53566 & n53592 ;
  assign n53594 = \pi0299  & ~n53561 ;
  assign n53595 = \pi0299  & ~\pi1091  ;
  assign n53596 = ~n53558 & n53595 ;
  assign n53597 = ~n53594 & ~n53596 ;
  assign n53598 = ~n53564 & n53597 ;
  assign n53599 = n53538 & n53597 ;
  assign n53600 = ~n53553 & n53599 ;
  assign n53601 = ~n53598 & ~n53600 ;
  assign n53602 = \pi0243  & n53601 ;
  assign n53603 = ~n53593 & n53602 ;
  assign n53604 = \pi1155  & ~n53583 ;
  assign n53605 = ~n53603 & n53604 ;
  assign n53606 = ~n53584 & ~n53605 ;
  assign n53607 = ~\pi0243  & ~\pi1155  ;
  assign n53608 = ~\pi0299  & ~\pi1091  ;
  assign n53609 = n53555 & n53608 ;
  assign n53610 = ~n13558 & ~n53609 ;
  assign n53611 = ~n53585 & ~n53610 ;
  assign n53612 = ~n53575 & ~n53611 ;
  assign n53613 = ~n53569 & n53612 ;
  assign n53614 = n53607 & ~n53613 ;
  assign n53615 = \pi0243  & ~\pi1091  ;
  assign n53616 = ~n53568 & ~n53575 ;
  assign n53617 = ~n53615 & ~n53616 ;
  assign n53618 = ~n53568 & ~n53586 ;
  assign n53619 = ~n53580 & ~n53618 ;
  assign n53620 = \pi0243  & ~\pi1155  ;
  assign n53621 = ~n53619 & n53620 ;
  assign n53622 = ~n53566 & n53621 ;
  assign n53623 = ~n53617 & ~n53622 ;
  assign n53624 = ~n53614 & n53623 ;
  assign n53625 = n53606 & n53624 ;
  assign n53626 = \pi1156  & ~n53625 ;
  assign n53627 = \pi0243  & ~\pi0299  ;
  assign n53628 = \pi0243  & n53542 ;
  assign n53629 = n53540 & n53628 ;
  assign n53630 = ~n53627 & ~n53629 ;
  assign n53631 = ~n53564 & ~n53630 ;
  assign n53632 = n53538 & ~n53630 ;
  assign n53633 = ~n53553 & n53632 ;
  assign n53634 = ~n53631 & ~n53633 ;
  assign n53635 = ~\pi1156  & ~n53586 ;
  assign n53636 = ~\pi1156  & n53538 ;
  assign n53637 = ~n53553 & n53636 ;
  assign n53638 = ~n53635 & ~n53637 ;
  assign n53639 = ~n53634 & ~n53638 ;
  assign n53640 = ~\pi1155  & n53597 ;
  assign n53641 = ~n53611 & n53640 ;
  assign n53642 = ~n53620 & ~n53641 ;
  assign n53643 = \pi1155  & ~\pi1156  ;
  assign n53644 = n53538 & ~n53568 ;
  assign n53645 = ~n53553 & n53644 ;
  assign n53646 = ~\pi1156  & ~n53577 ;
  assign n53647 = ~n53645 & n53646 ;
  assign n53648 = ~n53643 & ~n53647 ;
  assign n53649 = n53642 & ~n53648 ;
  assign n53650 = ~n53639 & ~n53649 ;
  assign n53651 = ~\pi0243  & n53569 ;
  assign n53652 = ~\pi0243  & ~\pi0299  ;
  assign n53653 = ~n53585 & n53652 ;
  assign n53654 = ~n53651 & ~n53653 ;
  assign n53655 = \pi1155  & n53634 ;
  assign n53656 = n53654 & n53655 ;
  assign n53657 = ~n53650 & ~n53656 ;
  assign n53658 = \pi1157  & ~n53657 ;
  assign n53659 = ~n53626 & n53658 ;
  assign n53660 = ~n53577 & ~n53645 ;
  assign n53661 = n53538 & ~n53591 ;
  assign n53662 = ~n53553 & n53661 ;
  assign n53663 = ~\pi0243  & ~\pi1091  ;
  assign n53664 = \pi0299  & n53590 ;
  assign n53665 = n53663 & ~n53664 ;
  assign n53666 = ~n53662 & n53665 ;
  assign n53667 = ~\pi1155  & ~n53666 ;
  assign n53668 = n53660 & n53667 ;
  assign n53669 = ~\pi1156  & ~n53607 ;
  assign n53670 = ~n53647 & ~n53669 ;
  assign n53671 = ~n53668 & ~n53670 ;
  assign n53672 = \pi1155  & ~n53615 ;
  assign n53673 = n53572 & n53672 ;
  assign n53674 = ~n53559 & n53673 ;
  assign n53675 = ~n53656 & ~n53674 ;
  assign n53676 = n53671 & n53675 ;
  assign n53677 = ~n53554 & ~n53610 ;
  assign n53678 = ~n53569 & ~n53677 ;
  assign n53679 = \pi0243  & ~n53678 ;
  assign n53680 = ~\pi0243  & n53542 ;
  assign n53681 = n53540 & n53680 ;
  assign n53682 = ~n53652 & ~n53681 ;
  assign n53683 = ~n53586 & ~n53682 ;
  assign n53684 = n53538 & ~n53682 ;
  assign n53685 = ~n53553 & n53684 ;
  assign n53686 = ~n53683 & ~n53685 ;
  assign n53687 = ~\pi1155  & ~n53538 ;
  assign n53688 = ~n53568 & n53687 ;
  assign n53689 = \pi1156  & ~n53688 ;
  assign n53690 = \pi1156  & n53564 ;
  assign n53691 = ~n53554 & n53690 ;
  assign n53692 = ~n53689 & ~n53691 ;
  assign n53693 = n53686 & ~n53692 ;
  assign n53694 = ~n53679 & n53693 ;
  assign n53695 = ~\pi1157  & ~n53694 ;
  assign n53696 = ~n53676 & n53695 ;
  assign n53697 = \pi0211  & ~n53696 ;
  assign n53698 = ~n53659 & n53697 ;
  assign n53699 = ~n53679 & n53686 ;
  assign n53700 = ~\pi0243  & ~n53577 ;
  assign n53701 = ~n53580 & n53700 ;
  assign n53702 = ~n53554 & n53564 ;
  assign n53703 = \pi0243  & ~n53569 ;
  assign n53704 = ~n53702 & n53703 ;
  assign n53705 = ~n53701 & ~n53704 ;
  assign n53706 = n53699 & ~n53705 ;
  assign n53707 = \pi1155  & ~n53706 ;
  assign n53708 = ~\pi0211  & ~n53670 ;
  assign n53709 = ~n53668 & n53708 ;
  assign n53710 = ~n53707 & n53709 ;
  assign n53711 = \pi0211  & ~\pi0219  ;
  assign n53712 = ~\pi1155  & ~n53569 ;
  assign n53713 = ~n53702 & n53712 ;
  assign n53714 = n53581 & n53713 ;
  assign n53715 = ~n53692 & ~n53714 ;
  assign n53716 = n53699 & n53715 ;
  assign n53717 = ~\pi0219  & ~\pi1157  ;
  assign n53718 = ~n53716 & n53717 ;
  assign n53719 = ~n53711 & ~n53718 ;
  assign n53720 = ~n53710 & ~n53719 ;
  assign n53721 = ~n53614 & ~n53622 ;
  assign n53722 = n53606 & n53721 ;
  assign n53723 = \pi1156  & ~n53722 ;
  assign n53724 = \pi1157  & n53705 ;
  assign n53725 = \pi1157  & ~n53639 ;
  assign n53726 = ~n53649 & n53725 ;
  assign n53727 = ~n53724 & ~n53726 ;
  assign n53728 = ~\pi0219  & ~n53727 ;
  assign n53729 = ~n53723 & n53728 ;
  assign n53730 = ~n53720 & ~n53729 ;
  assign n53731 = ~n53698 & ~n53730 ;
  assign n53732 = \pi0253  & \pi0254  ;
  assign n53733 = ~\pi0263  & \pi0267  ;
  assign n53734 = n53732 & n53733 ;
  assign n53735 = ~\pi0219  & n53734 ;
  assign n53736 = \pi0243  & ~n53591 ;
  assign n53737 = n53538 & n53736 ;
  assign n53738 = ~n53553 & n53737 ;
  assign n53739 = ~n53564 & n53736 ;
  assign n53740 = ~n53738 & ~n53739 ;
  assign n53741 = n53654 & n53740 ;
  assign n53742 = \pi1155  & ~n53741 ;
  assign n53743 = ~n53564 & ~n53591 ;
  assign n53744 = ~n53662 & ~n53743 ;
  assign n53745 = \pi0243  & n53538 ;
  assign n53746 = ~n53553 & n53745 ;
  assign n53747 = \pi0243  & ~n53586 ;
  assign n53748 = ~n53746 & ~n53747 ;
  assign n53749 = ~n53744 & ~n53748 ;
  assign n53750 = n53597 & ~n53611 ;
  assign n53751 = ~\pi0243  & ~n53750 ;
  assign n53752 = ~n53749 & ~n53751 ;
  assign n53753 = ~n53742 & n53752 ;
  assign n53754 = ~\pi1156  & ~n53753 ;
  assign n53755 = \pi0211  & ~n53754 ;
  assign n53756 = ~n53575 & n53597 ;
  assign n53757 = ~\pi0243  & ~n53756 ;
  assign n53758 = ~n53587 & n53736 ;
  assign n53759 = ~n53566 & n53758 ;
  assign n53760 = ~n53757 & ~n53759 ;
  assign n53761 = \pi1156  & ~n53760 ;
  assign n53762 = \pi1155  & n53654 ;
  assign n53763 = ~n53566 & n53736 ;
  assign n53764 = n53762 & ~n53763 ;
  assign n53765 = \pi1156  & n53642 ;
  assign n53766 = ~n53764 & n53765 ;
  assign n53767 = ~n53761 & ~n53766 ;
  assign n53768 = \pi1157  & n53767 ;
  assign n53769 = n53755 & n53768 ;
  assign n53770 = ~n53591 & ~n53677 ;
  assign n53771 = n50458 & ~n53585 ;
  assign n53772 = \pi0243  & ~n53771 ;
  assign n53773 = n53770 & n53772 ;
  assign n53774 = n53688 & ~n53702 ;
  assign n53775 = ~n53586 & n53597 ;
  assign n53776 = ~n53600 & ~n53775 ;
  assign n53777 = ~\pi0243  & n53776 ;
  assign n53778 = ~n53774 & n53777 ;
  assign n53779 = ~n53773 & ~n53778 ;
  assign n53780 = \pi1156  & ~n53779 ;
  assign n53781 = ~n53677 & ~n53740 ;
  assign n53782 = \pi0243  & \pi1155  ;
  assign n53783 = \pi1155  & n53597 ;
  assign n53784 = ~n53782 & ~n53783 ;
  assign n53785 = n53586 & ~n53782 ;
  assign n53786 = ~n53585 & n53785 ;
  assign n53787 = ~n53784 & ~n53786 ;
  assign n53788 = ~n53781 & n53787 ;
  assign n53789 = ~\pi1155  & ~n53663 ;
  assign n53790 = ~n53664 & n53789 ;
  assign n53791 = ~n53662 & n53790 ;
  assign n53792 = ~\pi1156  & ~n53664 ;
  assign n53793 = ~n53662 & n53792 ;
  assign n53794 = ~n53669 & ~n53793 ;
  assign n53795 = ~n53791 & ~n53794 ;
  assign n53796 = ~n53788 & n53795 ;
  assign n53797 = ~\pi1157  & ~n53796 ;
  assign n53798 = ~n53780 & n53797 ;
  assign n53799 = ~n53769 & ~n53798 ;
  assign n53800 = ~\pi0243  & n53597 ;
  assign n53801 = ~n53575 & n53800 ;
  assign n53802 = ~n53578 & ~n53591 ;
  assign n53803 = ~n53553 & n53802 ;
  assign n53804 = ~n53664 & ~n53803 ;
  assign n53805 = n53801 & ~n53804 ;
  assign n53806 = \pi1155  & \pi1156  ;
  assign n53807 = ~n53805 & n53806 ;
  assign n53808 = ~n53603 & n53807 ;
  assign n53809 = ~n53617 & ~n53751 ;
  assign n53810 = n53760 & n53809 ;
  assign n53811 = ~\pi1155  & \pi1156  ;
  assign n53812 = ~n53810 & n53811 ;
  assign n53813 = ~n53808 & ~n53812 ;
  assign n53814 = ~n53591 & ~n53611 ;
  assign n53815 = ~\pi0243  & ~n53814 ;
  assign n53816 = ~\pi1155  & n53748 ;
  assign n53817 = ~n53815 & n53816 ;
  assign n53818 = ~\pi0243  & \pi1155  ;
  assign n53819 = ~n53804 & n53818 ;
  assign n53820 = ~n53602 & ~n53819 ;
  assign n53821 = ~\pi1156  & n53820 ;
  assign n53822 = ~n53817 & n53821 ;
  assign n53823 = n50617 & ~n53822 ;
  assign n53824 = n53813 & n53823 ;
  assign n53825 = n53734 & ~n53824 ;
  assign n53826 = n53799 & n53825 ;
  assign n53827 = ~n53735 & ~n53826 ;
  assign n53828 = ~n53731 & ~n53827 ;
  assign n53829 = ~\pi0299  & \pi1091  ;
  assign n53830 = ~n50370 & n53829 ;
  assign n53831 = ~n50825 & n53830 ;
  assign n53832 = ~n53663 & ~n53831 ;
  assign n53833 = \pi1156  & ~n53832 ;
  assign n53834 = \pi1091  & ~n15351 ;
  assign n53835 = n51583 & n53834 ;
  assign n53836 = ~n53833 & ~n53835 ;
  assign n53837 = n50383 & n53829 ;
  assign n53838 = ~n53663 & ~n53837 ;
  assign n53839 = \pi1091  & \pi1155  ;
  assign n53840 = ~n53663 & ~n53839 ;
  assign n53841 = n44032 & ~n53840 ;
  assign n53842 = n53838 & ~n53841 ;
  assign n53843 = ~\pi1156  & ~n53842 ;
  assign n53844 = \pi1157  & ~n53843 ;
  assign n53845 = n53836 & n53844 ;
  assign n53846 = \pi0199  & \pi1091  ;
  assign n53847 = ~\pi0299  & n53846 ;
  assign n53848 = n53672 & ~n53847 ;
  assign n53849 = \pi1156  & ~n53848 ;
  assign n53850 = ~\pi1155  & ~n53615 ;
  assign n53851 = ~n13645 & n53829 ;
  assign n53852 = n53850 & ~n53851 ;
  assign n53853 = ~\pi1157  & ~n53852 ;
  assign n53854 = n53849 & n53853 ;
  assign n53855 = ~\pi1156  & n53840 ;
  assign n53856 = \pi1091  & ~\pi1156  ;
  assign n53857 = ~n15351 & n53856 ;
  assign n53858 = ~n53855 & ~n53857 ;
  assign n53859 = ~\pi1157  & ~n53858 ;
  assign n53860 = \pi0211  & ~n53859 ;
  assign n53861 = ~n53854 & n53860 ;
  assign n53862 = ~n53845 & n53861 ;
  assign n53863 = n53832 & n53849 ;
  assign n53864 = ~\pi1155  & ~n53838 ;
  assign n53865 = \pi0200  & \pi1091  ;
  assign n53866 = ~\pi0299  & n53865 ;
  assign n53867 = n53672 & ~n53866 ;
  assign n53868 = ~\pi1156  & ~n53867 ;
  assign n53869 = ~n53864 & n53868 ;
  assign n53870 = ~n53863 & ~n53869 ;
  assign n53871 = \pi1157  & ~n53870 ;
  assign n53872 = \pi0200  & ~\pi1156  ;
  assign n53873 = n53829 & n53872 ;
  assign n53874 = n53848 & ~n53873 ;
  assign n53875 = \pi1091  & ~n13646 ;
  assign n53876 = n53850 & ~n53873 ;
  assign n53877 = ~n53875 & n53876 ;
  assign n53878 = ~n53874 & ~n53877 ;
  assign n53879 = ~\pi1157  & n53878 ;
  assign n53880 = ~\pi0211  & ~n53879 ;
  assign n53881 = ~n53871 & n53880 ;
  assign n53882 = ~n53862 & ~n53881 ;
  assign n53883 = ~\pi0219  & ~n53882 ;
  assign n53884 = ~n50383 & n53829 ;
  assign n53885 = n53850 & ~n53884 ;
  assign n53886 = ~n53867 & ~n53885 ;
  assign n53887 = ~\pi1156  & ~n53886 ;
  assign n53888 = n50617 & ~n53887 ;
  assign n53889 = n53836 & n53888 ;
  assign n53890 = ~\pi1156  & n51349 ;
  assign n53891 = n51349 & ~n53663 ;
  assign n53892 = ~n53831 & n53891 ;
  assign n53893 = ~n53890 & ~n53892 ;
  assign n53894 = ~n53843 & ~n53893 ;
  assign n53895 = \pi0219  & ~n53894 ;
  assign n53896 = \pi0299  & \pi1091  ;
  assign n53897 = ~n53878 & ~n53896 ;
  assign n53898 = ~\pi1157  & ~n53897 ;
  assign n53899 = n53895 & ~n53898 ;
  assign n53900 = ~n53889 & n53899 ;
  assign n53901 = n27408 & ~n53900 ;
  assign n53902 = ~n53883 & n53901 ;
  assign n53903 = \pi0272  & \pi0283  ;
  assign n53904 = \pi0268  & \pi0275  ;
  assign n53905 = n53903 & n53904 ;
  assign n53906 = \pi1091  & \pi1157  ;
  assign n53907 = n50689 & n53906 ;
  assign n53908 = ~n50608 & ~n50618 ;
  assign n53909 = ~\pi0219  & \pi1091  ;
  assign n53910 = ~n53908 & n53909 ;
  assign n53911 = ~n53907 & ~n53910 ;
  assign n53912 = ~n27408 & ~n53663 ;
  assign n53913 = n53911 & n53912 ;
  assign n53914 = ~n53905 & ~n53913 ;
  assign n53915 = ~n53902 & n53914 ;
  assign n53916 = ~n53734 & n53900 ;
  assign n53917 = ~\pi0219  & ~n53734 ;
  assign n53918 = ~n53882 & n53917 ;
  assign n53919 = ~n53916 & ~n53918 ;
  assign n53920 = ~\pi0230  & n27408 ;
  assign n53921 = n53919 & n53920 ;
  assign n53922 = ~n53915 & n53921 ;
  assign n53923 = ~n53828 & n53922 ;
  assign n53924 = ~n53543 & n53615 ;
  assign n53925 = ~n53551 & n53924 ;
  assign n53926 = \pi1091  & n53908 ;
  assign n53927 = ~n53681 & ~n53926 ;
  assign n53928 = ~n53925 & n53927 ;
  assign n53929 = ~\pi0219  & ~n53928 ;
  assign n53930 = ~\pi0243  & ~n53561 ;
  assign n53931 = ~n53558 & n53663 ;
  assign n53932 = ~n53930 & ~n53931 ;
  assign n53933 = \pi0276  & n53541 ;
  assign n53934 = n53545 & n53933 ;
  assign n53935 = \pi0243  & \pi0273  ;
  assign n53936 = n53934 & n53935 ;
  assign n53937 = n53536 & n53545 ;
  assign n53938 = n50617 & ~n53615 ;
  assign n53939 = ~n53937 & n53938 ;
  assign n53940 = ~n53936 & ~n53939 ;
  assign n53941 = \pi0219  & n53940 ;
  assign n53942 = n53932 & n53941 ;
  assign n53943 = n53734 & ~n53942 ;
  assign n53944 = ~n53929 & n53943 ;
  assign n53945 = ~n9948 & n53734 ;
  assign n53946 = ~n53913 & ~n53945 ;
  assign n53947 = ~n53944 & ~n53946 ;
  assign n53948 = n53905 & ~n53947 ;
  assign n53949 = ~\pi0230  & ~n53948 ;
  assign n53950 = ~n53915 & n53949 ;
  assign n53951 = ~\pi0219  & ~n53908 ;
  assign n53952 = \pi1157  & n50689 ;
  assign n53953 = \pi0230  & ~n53952 ;
  assign n53954 = ~n20516 & n53953 ;
  assign n53955 = ~n53951 & n53954 ;
  assign n53956 = \pi0199  & ~n51573 ;
  assign n53957 = ~n50825 & ~n53956 ;
  assign n53958 = ~n53872 & n53957 ;
  assign n53959 = \pi0230  & n20515 ;
  assign n53960 = n6848 & n53959 ;
  assign n53961 = ~n53958 & n53960 ;
  assign n53962 = ~n53955 & ~n53961 ;
  assign n53963 = ~n53950 & n53962 ;
  assign n53964 = ~n53923 & n53963 ;
  assign n53965 = ~\pi0230  & \pi0244  ;
  assign n53966 = n52891 & ~n52899 ;
  assign n53967 = ~n52877 & ~n53966 ;
  assign n53968 = n52873 & ~n53967 ;
  assign n53969 = \pi0209  & \pi0213  ;
  assign n53970 = ~n53968 & n53969 ;
  assign n53971 = ~\pi0213  & ~n51663 ;
  assign n53972 = ~n51671 & n51766 ;
  assign n53973 = ~n53971 & ~n53972 ;
  assign n53974 = \pi0219  & \pi0299  ;
  assign n53975 = ~n50661 & n53974 ;
  assign n53976 = \pi1147  & ~n53975 ;
  assign n53977 = n9948 & n53976 ;
  assign n53978 = ~n52543 & n53977 ;
  assign n53979 = ~n53973 & ~n53978 ;
  assign n53980 = ~n52528 & n52661 ;
  assign n53981 = ~n52660 & ~n53980 ;
  assign n53982 = ~\pi0211  & n51640 ;
  assign n53983 = ~\pi1144  & n52001 ;
  assign n53984 = ~n53982 & ~n53983 ;
  assign n53985 = n52541 & n53984 ;
  assign n53986 = n50954 & ~n53985 ;
  assign n53987 = n53981 & ~n53986 ;
  assign n53988 = n50659 & n50693 ;
  assign n53989 = \pi0212  & ~n53988 ;
  assign n53990 = n53984 & n53989 ;
  assign n53991 = n52541 & n53990 ;
  assign n53992 = \pi0214  & n53989 ;
  assign n53993 = n52541 & n53992 ;
  assign n53994 = ~n53991 & ~n53993 ;
  assign n53995 = ~n53973 & n53994 ;
  assign n53996 = ~n53987 & n53995 ;
  assign n53997 = ~n53979 & ~n53996 ;
  assign n53998 = ~\pi0214  & ~n53985 ;
  assign n53999 = ~n52583 & n53989 ;
  assign n54000 = ~n53998 & n53999 ;
  assign n54001 = n52862 & n53984 ;
  assign n54002 = n52541 & n54001 ;
  assign n54003 = ~n52583 & n54002 ;
  assign n54004 = n52633 & ~n52859 ;
  assign n54005 = ~\pi0219  & ~n54004 ;
  assign n54006 = ~n54003 & n54005 ;
  assign n54007 = ~n54000 & n54006 ;
  assign n54008 = n52558 & ~n52879 ;
  assign n54009 = ~\pi0211  & ~n50740 ;
  assign n54010 = ~n52571 & n54009 ;
  assign n54011 = ~n52570 & n54010 ;
  assign n54012 = ~\pi1143  & n52000 ;
  assign n54013 = ~n50570 & ~n54012 ;
  assign n54014 = n52558 & n54013 ;
  assign n54015 = n52886 & n54014 ;
  assign n54016 = ~n54011 & n54015 ;
  assign n54017 = ~n54008 & ~n54016 ;
  assign n54018 = ~n54007 & ~n54017 ;
  assign n54019 = \pi0209  & ~n54018 ;
  assign n54020 = ~n53997 & n54019 ;
  assign n54021 = ~\pi0230  & ~\pi0244  ;
  assign n54022 = n46207 & ~n51733 ;
  assign n54023 = ~\pi0219  & ~n51671 ;
  assign n54024 = ~\pi0213  & n51663 ;
  assign n54025 = ~n54023 & n54024 ;
  assign n54026 = ~\pi0209  & ~n54025 ;
  assign n54027 = ~n54022 & n54026 ;
  assign n54028 = ~n54021 & ~n54027 ;
  assign n54029 = \pi0299  & ~n52907 ;
  assign n54030 = ~n52877 & ~n54029 ;
  assign n54031 = n12255 & ~n52837 ;
  assign n54032 = ~n12255 & ~n52846 ;
  assign n54033 = n9948 & ~n54032 ;
  assign n54034 = ~n54031 & n54033 ;
  assign n54035 = n50948 & n54034 ;
  assign n54036 = ~n54030 & n54035 ;
  assign n54037 = ~\pi1147  & n52909 ;
  assign n54038 = ~n52907 & n54037 ;
  assign n54039 = \pi1147  & n12577 ;
  assign n54040 = n50679 & n54039 ;
  assign n54041 = ~n9948 & n54040 ;
  assign n54042 = ~n54038 & ~n54041 ;
  assign n54043 = ~n52826 & n54042 ;
  assign n54044 = ~\pi0299  & n9948 ;
  assign n54045 = ~n51726 & n54044 ;
  assign n54046 = n9948 & n52921 ;
  assign n54047 = ~n54045 & ~n54046 ;
  assign n54048 = n54043 & n54047 ;
  assign n54049 = ~n54036 & n54048 ;
  assign n54050 = \pi0213  & ~n54021 ;
  assign n54051 = ~n54049 & n54050 ;
  assign n54052 = ~n54028 & ~n54051 ;
  assign n54053 = ~n54020 & ~n54052 ;
  assign n54054 = ~n53970 & n54053 ;
  assign n54055 = ~n53965 & ~n54054 ;
  assign n54056 = ~\pi0230  & \pi0245  ;
  assign n54057 = ~n52535 & ~n53440 ;
  assign n54058 = n53437 & n54057 ;
  assign n54059 = n50571 & ~n54058 ;
  assign n54060 = n9948 & n54059 ;
  assign n54061 = ~n53484 & ~n54060 ;
  assign n54062 = \pi1147  & n52229 ;
  assign n54063 = \pi0219  & \pi1146  ;
  assign n54064 = n12255 & n52814 ;
  assign n54065 = ~n54063 & ~n54064 ;
  assign n54066 = n50677 & ~n54065 ;
  assign n54067 = n50805 & n52229 ;
  assign n54068 = ~n54066 & ~n54067 ;
  assign n54069 = ~n54062 & n54068 ;
  assign n54070 = n54061 & n54069 ;
  assign n54071 = \pi1148  & ~n54070 ;
  assign n54072 = ~\pi0299  & ~n53440 ;
  assign n54073 = n53437 & n54072 ;
  assign n54074 = n50967 & ~n54073 ;
  assign n54075 = n50430 & ~n54058 ;
  assign n54076 = ~n54074 & ~n54075 ;
  assign n54077 = ~\pi0214  & ~n54073 ;
  assign n54078 = n54076 & ~n54077 ;
  assign n54079 = \pi0212  & ~n54078 ;
  assign n54080 = \pi1147  & ~n52229 ;
  assign n54081 = ~n54066 & n54080 ;
  assign n54082 = n53437 & n53471 ;
  assign n54083 = ~\pi0212  & ~n54073 ;
  assign n54084 = ~n54082 & n54083 ;
  assign n54085 = n54081 & ~n54084 ;
  assign n54086 = ~n54079 & n54085 ;
  assign n54087 = ~\pi0219  & n54086 ;
  assign n54088 = ~\pi0212  & ~n54082 ;
  assign n54089 = \pi0211  & \pi0212  ;
  assign n54090 = n52535 & n54089 ;
  assign n54091 = ~n50600 & ~n54090 ;
  assign n54092 = \pi0212  & ~\pi0299  ;
  assign n54093 = n53447 & n54092 ;
  assign n54094 = n54091 & ~n54093 ;
  assign n54095 = ~n54088 & n54094 ;
  assign n54096 = \pi0214  & ~n54091 ;
  assign n54097 = \pi0214  & n54092 ;
  assign n54098 = n53447 & n54097 ;
  assign n54099 = ~n54096 & ~n54098 ;
  assign n54100 = ~\pi0211  & ~n54073 ;
  assign n54101 = n53437 & ~n53470 ;
  assign n54102 = ~n54100 & n54101 ;
  assign n54103 = n54099 & n54102 ;
  assign n54104 = ~n54095 & ~n54103 ;
  assign n54105 = ~\pi1147  & ~n54066 ;
  assign n54106 = ~n54067 & n54105 ;
  assign n54107 = ~\pi0219  & n54106 ;
  assign n54108 = ~n54104 & n54107 ;
  assign n54109 = ~n54087 & ~n54108 ;
  assign n54110 = n54071 & n54109 ;
  assign n54111 = ~n52642 & ~n54081 ;
  assign n54112 = n54061 & ~n54111 ;
  assign n54113 = ~n52001 & ~n53470 ;
  assign n54114 = n53437 & n54113 ;
  assign n54115 = ~\pi0214  & ~n54114 ;
  assign n54116 = n54076 & ~n54115 ;
  assign n54117 = \pi0212  & ~n54116 ;
  assign n54118 = n54088 & ~n54114 ;
  assign n54119 = ~\pi0219  & ~n54111 ;
  assign n54120 = ~n54118 & n54119 ;
  assign n54121 = ~n54117 & n54120 ;
  assign n54122 = ~n54112 & ~n54121 ;
  assign n54123 = ~n54082 & ~n54094 ;
  assign n54124 = ~\pi0219  & ~n53470 ;
  assign n54125 = n53437 & n54124 ;
  assign n54126 = ~n52660 & ~n54125 ;
  assign n54127 = n54105 & ~n54126 ;
  assign n54128 = ~n54123 & n54127 ;
  assign n54129 = n54061 & n54105 ;
  assign n54130 = ~\pi1148  & ~n54129 ;
  assign n54131 = ~n54128 & n54130 ;
  assign n54132 = n54122 & n54131 ;
  assign n54133 = ~\pi0209  & \pi0213  ;
  assign n54134 = ~n54132 & n54133 ;
  assign n54135 = ~n54110 & n54134 ;
  assign n54136 = \pi0199  & \pi1146  ;
  assign n54137 = ~\pi0200  & ~n54136 ;
  assign n54138 = n50824 & ~n54137 ;
  assign n54139 = ~n12409 & ~n54138 ;
  assign n54140 = ~n52001 & n54139 ;
  assign n54141 = n50383 & ~n54136 ;
  assign n54142 = \pi0207  & ~n54141 ;
  assign n54143 = n52524 & n54142 ;
  assign n54144 = ~n50877 & ~n52001 ;
  assign n54145 = ~n54143 & n54144 ;
  assign n54146 = ~n54140 & ~n54145 ;
  assign n54147 = \pi0214  & n54146 ;
  assign n54148 = ~n50877 & ~n54143 ;
  assign n54149 = ~\pi0214  & ~n54139 ;
  assign n54150 = ~n54148 & n54149 ;
  assign n54151 = ~\pi0212  & ~n54150 ;
  assign n54152 = ~n54147 & n54151 ;
  assign n54153 = ~\pi0299  & n54137 ;
  assign n54154 = ~\pi0299  & ~n50418 ;
  assign n54155 = ~n50840 & ~n54154 ;
  assign n54156 = ~n54153 & n54155 ;
  assign n54157 = \pi0214  & n54156 ;
  assign n54158 = ~n50370 & n50410 ;
  assign n54159 = ~n54137 & n54158 ;
  assign n54160 = ~n52535 & ~n54159 ;
  assign n54161 = ~n54143 & n54160 ;
  assign n54162 = \pi0208  & \pi0214  ;
  assign n54163 = ~n54161 & n54162 ;
  assign n54164 = ~n54157 & ~n54163 ;
  assign n54165 = n50824 & ~n54141 ;
  assign n54166 = ~n12409 & ~n54165 ;
  assign n54167 = ~n54148 & ~n54166 ;
  assign n54168 = \pi0199  & ~\pi1146  ;
  assign n54169 = \pi0208  & ~\pi1146  ;
  assign n54170 = n51915 & n54169 ;
  assign n54171 = ~n54168 & ~n54170 ;
  assign n54172 = n52798 & n54171 ;
  assign n54173 = ~\pi0299  & ~n54172 ;
  assign n54174 = ~\pi0211  & ~n54173 ;
  assign n54175 = ~n54167 & ~n54174 ;
  assign n54176 = ~n54164 & ~n54175 ;
  assign n54177 = ~\pi0214  & n54146 ;
  assign n54178 = \pi0212  & ~n54177 ;
  assign n54179 = ~n54176 & n54178 ;
  assign n54180 = ~n54152 & ~n54179 ;
  assign n54181 = ~\pi0219  & ~\pi1146  ;
  assign n54182 = ~n50443 & n54181 ;
  assign n54183 = ~n53172 & ~n54182 ;
  assign n54184 = ~n54180 & ~n54183 ;
  assign n54185 = n50570 & ~n54139 ;
  assign n54186 = ~n54148 & n54185 ;
  assign n54187 = \pi0219  & ~n54186 ;
  assign n54188 = \pi0211  & n54139 ;
  assign n54189 = n50924 & ~n54143 ;
  assign n54190 = ~n54188 & ~n54189 ;
  assign n54191 = ~n50570 & n54190 ;
  assign n54192 = \pi0208  & ~n54161 ;
  assign n54193 = ~\pi0208  & n52535 ;
  assign n54194 = n50418 & n54138 ;
  assign n54195 = ~n54193 & ~n54194 ;
  assign n54196 = ~n54192 & n54195 ;
  assign n54197 = n54191 & ~n54196 ;
  assign n54198 = n54187 & ~n54197 ;
  assign n54199 = n27408 & ~n54198 ;
  assign n54200 = ~n54184 & n54199 ;
  assign n54201 = ~n54111 & ~n54200 ;
  assign n54202 = ~\pi1148  & ~n54105 ;
  assign n54203 = n44032 & n54136 ;
  assign n54204 = ~n52554 & ~n54203 ;
  assign n54205 = n12409 & ~n54204 ;
  assign n54206 = \pi0208  & \pi1146  ;
  assign n54207 = ~n50384 & n54206 ;
  assign n54208 = ~n54205 & ~n54207 ;
  assign n54209 = \pi0200  & ~\pi0207  ;
  assign n54210 = ~n52515 & n54209 ;
  assign n54211 = ~n51930 & ~n54210 ;
  assign n54212 = n52031 & ~n54141 ;
  assign n54213 = n54211 & n54212 ;
  assign n54214 = n54208 & ~n54213 ;
  assign n54215 = \pi1146  & ~n50384 ;
  assign n54216 = \pi0207  & ~n54204 ;
  assign n54217 = ~n54215 & ~n54216 ;
  assign n54218 = ~\pi0299  & ~n54217 ;
  assign n54219 = ~n54214 & n54218 ;
  assign n54220 = n53183 & n54215 ;
  assign n54221 = \pi0207  & n53183 ;
  assign n54222 = ~n54204 & n54221 ;
  assign n54223 = ~n54220 & ~n54222 ;
  assign n54224 = ~\pi0219  & n54223 ;
  assign n54225 = ~n54219 & n54224 ;
  assign n54226 = n9948 & ~n54225 ;
  assign n54227 = n44032 & ~n50876 ;
  assign n54228 = ~n12409 & ~n54227 ;
  assign n54229 = ~n54204 & ~n54228 ;
  assign n54230 = \pi0219  & ~n54229 ;
  assign n54231 = ~n51108 & ~n54230 ;
  assign n54232 = ~n54193 & ~n54207 ;
  assign n54233 = ~n54205 & n54232 ;
  assign n54234 = ~n54213 & n54233 ;
  assign n54235 = \pi0211  & ~n54229 ;
  assign n54236 = n44032 & ~n54136 ;
  assign n54237 = n44035 & ~n52515 ;
  assign n54238 = ~n54236 & ~n54237 ;
  assign n54239 = ~n50570 & n54238 ;
  assign n54240 = ~n54235 & n54239 ;
  assign n54241 = ~n54234 & n54240 ;
  assign n54242 = ~n54231 & ~n54241 ;
  assign n54243 = ~\pi1148  & ~n54242 ;
  assign n54244 = n54226 & n54243 ;
  assign n54245 = ~n54202 & ~n54244 ;
  assign n54246 = ~n54201 & ~n54245 ;
  assign n54247 = ~\pi0212  & ~\pi0299  ;
  assign n54248 = ~n54214 & n54247 ;
  assign n54249 = ~n50556 & ~n54248 ;
  assign n54250 = ~\pi0299  & ~n54214 ;
  assign n54251 = n54235 & ~n54250 ;
  assign n54252 = ~\pi0211  & ~\pi0299  ;
  assign n54253 = n54214 & n54252 ;
  assign n54254 = ~n54251 & ~n54253 ;
  assign n54255 = ~n54249 & n54254 ;
  assign n54256 = ~\pi0219  & ~n54255 ;
  assign n54257 = ~\pi0214  & n54253 ;
  assign n54258 = ~\pi0214  & n54235 ;
  assign n54259 = ~n54250 & n54258 ;
  assign n54260 = ~n54257 & ~n54259 ;
  assign n54261 = \pi0214  & ~n52854 ;
  assign n54262 = \pi0212  & ~n54261 ;
  assign n54263 = n54092 & ~n54214 ;
  assign n54264 = ~n54262 & ~n54263 ;
  assign n54265 = n54260 & ~n54264 ;
  assign n54266 = n54256 & ~n54265 ;
  assign n54267 = n50880 & ~n54165 ;
  assign n54268 = n50878 & ~n54143 ;
  assign n54269 = ~n54267 & ~n54268 ;
  assign n54270 = ~\pi0212  & ~n54173 ;
  assign n54271 = n54269 & n54270 ;
  assign n54272 = ~\pi0219  & ~n54271 ;
  assign n54273 = \pi0212  & ~n54173 ;
  assign n54274 = n50430 & ~n52535 ;
  assign n54275 = ~n54172 & n54274 ;
  assign n54276 = n54273 & ~n54275 ;
  assign n54277 = n54272 & ~n54276 ;
  assign n54278 = ~n50571 & ~n54166 ;
  assign n54279 = ~n54148 & n54278 ;
  assign n54280 = \pi0219  & ~n54279 ;
  assign n54281 = ~n52535 & ~n54172 ;
  assign n54282 = n50571 & ~n54281 ;
  assign n54283 = n54280 & ~n54282 ;
  assign n54284 = n27408 & ~n54283 ;
  assign n54285 = ~n54277 & n54284 ;
  assign n54286 = n54081 & ~n54285 ;
  assign n54287 = ~\pi0299  & ~n50571 ;
  assign n54288 = ~n54214 & n54287 ;
  assign n54289 = \pi0219  & ~n54288 ;
  assign n54290 = n50571 & ~n54234 ;
  assign n54291 = n54289 & ~n54290 ;
  assign n54292 = \pi1148  & n27408 ;
  assign n54293 = ~n54291 & n54292 ;
  assign n54294 = ~n54286 & n54293 ;
  assign n54295 = ~n54266 & n54294 ;
  assign n54296 = \pi1148  & ~n54106 ;
  assign n54297 = ~n54286 & n54296 ;
  assign n54298 = n53969 & ~n54297 ;
  assign n54299 = ~n54295 & n54298 ;
  assign n54300 = ~n54246 & n54299 ;
  assign n54301 = ~n54135 & ~n54300 ;
  assign n54302 = ~\pi0230  & ~\pi0245  ;
  assign n54303 = ~n52837 & ~n54250 ;
  assign n54304 = ~n54249 & ~n54303 ;
  assign n54305 = ~\pi0214  & \pi0299  ;
  assign n54306 = ~n52818 & n54305 ;
  assign n54307 = n50693 & ~n51667 ;
  assign n54308 = ~n54306 & ~n54307 ;
  assign n54309 = \pi0212  & ~n54308 ;
  assign n54310 = ~n54263 & ~n54309 ;
  assign n54311 = ~\pi0219  & n54310 ;
  assign n54312 = ~n54304 & n54311 ;
  assign n54313 = ~\pi0299  & ~n54207 ;
  assign n54314 = ~n54205 & n54313 ;
  assign n54315 = ~n54213 & n54314 ;
  assign n54316 = n50571 & ~n50779 ;
  assign n54317 = ~n54315 & n54316 ;
  assign n54318 = n54289 & ~n54317 ;
  assign n54319 = n52558 & ~n54318 ;
  assign n54320 = ~n54312 & n54319 ;
  assign n54321 = ~\pi0057  & \pi1147  ;
  assign n54322 = n6848 & n54321 ;
  assign n54323 = ~n54172 & n54308 ;
  assign n54324 = \pi0212  & ~n54323 ;
  assign n54325 = ~\pi0219  & ~n54324 ;
  assign n54326 = n52838 & ~n54172 ;
  assign n54327 = ~\pi0212  & ~n54326 ;
  assign n54328 = n54269 & n54327 ;
  assign n54329 = n54325 & ~n54328 ;
  assign n54330 = ~n50783 & ~n54172 ;
  assign n54331 = n50571 & ~n54330 ;
  assign n54332 = n54280 & ~n54331 ;
  assign n54333 = ~n54329 & ~n54332 ;
  assign n54334 = n54322 & n54333 ;
  assign n54335 = \pi1148  & ~n54334 ;
  assign n54336 = ~n54320 & n54335 ;
  assign n54337 = \pi0209  & ~n54336 ;
  assign n54338 = ~\pi0213  & ~n53466 ;
  assign n54339 = ~\pi0209  & ~n53485 ;
  assign n54340 = n54338 & ~n54339 ;
  assign n54341 = ~n53476 & n54338 ;
  assign n54342 = ~n53457 & n54341 ;
  assign n54343 = ~n54340 & ~n54342 ;
  assign n54344 = ~n54337 & ~n54343 ;
  assign n54345 = n50570 & n54229 ;
  assign n54346 = \pi0299  & ~n52818 ;
  assign n54347 = ~\pi0299  & ~n54204 ;
  assign n54348 = ~n54214 & n54347 ;
  assign n54349 = ~n54346 & ~n54348 ;
  assign n54350 = n50556 & ~n54349 ;
  assign n54351 = ~n54345 & ~n54350 ;
  assign n54352 = n54238 & ~n54310 ;
  assign n54353 = ~\pi0219  & ~n54352 ;
  assign n54354 = n54351 & n54353 ;
  assign n54355 = n54238 & ~n54315 ;
  assign n54356 = ~n50570 & ~n50779 ;
  assign n54357 = ~n54235 & n54356 ;
  assign n54358 = n54355 & n54357 ;
  assign n54359 = ~n51730 & ~n54230 ;
  assign n54360 = ~n54358 & ~n54359 ;
  assign n54361 = n52558 & ~n54360 ;
  assign n54362 = ~n54354 & n54361 ;
  assign n54363 = ~\pi0212  & n54150 ;
  assign n54364 = ~n52837 & ~n54172 ;
  assign n54365 = ~\pi0212  & ~n54364 ;
  assign n54366 = ~n54164 & n54365 ;
  assign n54367 = ~n54363 & ~n54366 ;
  assign n54368 = ~\pi0219  & ~n54156 ;
  assign n54369 = ~n54192 & n54368 ;
  assign n54370 = ~n54325 & ~n54369 ;
  assign n54371 = n54367 & ~n54370 ;
  assign n54372 = n6848 & ~n54187 ;
  assign n54373 = ~\pi0211  & n54330 ;
  assign n54374 = ~\pi0211  & ~n54156 ;
  assign n54375 = ~n54192 & n54374 ;
  assign n54376 = ~n54373 & ~n54375 ;
  assign n54377 = n6848 & n54191 ;
  assign n54378 = n54376 & n54377 ;
  assign n54379 = ~n54372 & ~n54378 ;
  assign n54380 = n54321 & ~n54379 ;
  assign n54381 = ~n54371 & n54380 ;
  assign n54382 = ~n54362 & ~n54381 ;
  assign n54383 = ~\pi1148  & ~n54343 ;
  assign n54384 = n54382 & n54383 ;
  assign n54385 = ~n54344 & ~n54384 ;
  assign n54386 = ~n54302 & n54385 ;
  assign n54387 = n54301 & n54386 ;
  assign n54388 = ~n54056 & ~n54387 ;
  assign n54389 = n50693 & n52814 ;
  assign n54390 = ~n52741 & ~n54389 ;
  assign n54391 = ~n52768 & n54390 ;
  assign n54392 = ~n52765 & n54391 ;
  assign n54393 = n52710 & n52750 ;
  assign n54394 = ~n52743 & ~n54393 ;
  assign n54395 = \pi0219  & ~\pi1146  ;
  assign n54396 = ~n52741 & n54395 ;
  assign n54397 = ~\pi1150  & ~n54396 ;
  assign n54398 = ~n54394 & n54397 ;
  assign n54399 = ~n54392 & n54398 ;
  assign n54400 = \pi0219  & ~n52535 ;
  assign n54401 = n52710 & ~n54400 ;
  assign n54402 = ~n52988 & ~n54401 ;
  assign n54403 = \pi0212  & ~n52787 ;
  assign n54404 = n52773 & ~n53091 ;
  assign n54405 = n54403 & ~n54404 ;
  assign n54406 = n50430 & ~n52782 ;
  assign n54407 = ~\pi0219  & ~n51918 ;
  assign n54408 = ~n54406 & n54407 ;
  assign n54409 = ~n54405 & n54408 ;
  assign n54410 = ~n54402 & ~n54409 ;
  assign n54411 = n51972 & n52704 ;
  assign n54412 = ~\pi0219  & ~n52535 ;
  assign n54413 = ~n52775 & n54412 ;
  assign n54414 = ~n54411 & n54413 ;
  assign n54415 = ~\pi0212  & n50430 ;
  assign n54416 = ~n52782 & n54415 ;
  assign n54417 = ~n52995 & ~n54416 ;
  assign n54418 = n54414 & n54417 ;
  assign n54419 = ~n54405 & n54418 ;
  assign n54420 = \pi1150  & ~n54419 ;
  assign n54421 = n54410 & n54420 ;
  assign n54422 = ~n54111 & ~n54421 ;
  assign n54423 = ~n54399 & n54422 ;
  assign n54424 = n52774 & ~n52787 ;
  assign n54425 = ~\pi0219  & n53110 ;
  assign n54426 = ~n54424 & n54425 ;
  assign n54427 = \pi1150  & n9948 ;
  assign n54428 = ~n52985 & n54427 ;
  assign n54429 = ~n54426 & n54428 ;
  assign n54430 = ~n54419 & n54429 ;
  assign n54431 = n54410 & n54430 ;
  assign n54432 = ~\pi0219  & ~n53052 ;
  assign n54433 = ~n52767 & ~n54432 ;
  assign n54434 = ~\pi1146  & ~n52741 ;
  assign n54435 = ~\pi1150  & ~n54434 ;
  assign n54436 = n54433 & n54435 ;
  assign n54437 = ~n54394 & n54436 ;
  assign n54438 = n52790 & n54428 ;
  assign n54439 = ~n54426 & n54438 ;
  assign n54440 = n54105 & ~n54439 ;
  assign n54441 = ~n54437 & n54440 ;
  assign n54442 = ~n54431 & n54441 ;
  assign n54443 = ~\pi1148  & ~n54442 ;
  assign n54444 = ~n54423 & n54443 ;
  assign n54445 = ~n52709 & ~n54401 ;
  assign n54446 = n51975 & n54261 ;
  assign n54447 = n52698 & ~n54446 ;
  assign n54448 = ~n52695 & ~n54447 ;
  assign n54449 = ~n54445 & ~n54448 ;
  assign n54450 = ~n52700 & ~n53205 ;
  assign n54451 = n52698 & n54450 ;
  assign n54452 = ~n52723 & ~n54451 ;
  assign n54453 = ~n54106 & ~n54445 ;
  assign n54454 = ~n54452 & n54453 ;
  assign n54455 = ~n54449 & ~n54454 ;
  assign n54456 = ~\pi0219  & ~n52814 ;
  assign n54457 = ~n54400 & ~n54456 ;
  assign n54458 = ~n53184 & n54457 ;
  assign n54459 = n52710 & n54458 ;
  assign n54460 = ~n53018 & ~n54459 ;
  assign n54461 = n54106 & n54460 ;
  assign n54462 = ~n52798 & ~n53066 ;
  assign n54463 = n9948 & ~n54462 ;
  assign n54464 = \pi1146  & n52616 ;
  assign n54465 = n52710 & n54464 ;
  assign n54466 = ~n54463 & ~n54465 ;
  assign n54467 = n54081 & n54466 ;
  assign n54468 = \pi1150  & ~n54467 ;
  assign n54469 = ~n54461 & n54468 ;
  assign n54470 = n54069 & ~n54469 ;
  assign n54471 = n54455 & n54470 ;
  assign n54472 = \pi1148  & ~\pi1150  ;
  assign n54473 = \pi1148  & ~n54467 ;
  assign n54474 = ~n54461 & n54473 ;
  assign n54475 = ~n54472 & ~n54474 ;
  assign n54476 = ~n54471 & ~n54475 ;
  assign n54477 = \pi1149  & ~n54476 ;
  assign n54478 = ~n54444 & n54477 ;
  assign n54479 = ~n52975 & ~n54401 ;
  assign n54480 = n54081 & n54479 ;
  assign n54481 = \pi1150  & n54480 ;
  assign n54482 = n52958 & n53253 ;
  assign n54483 = ~\pi0212  & ~n52033 ;
  assign n54484 = ~\pi0219  & ~n54483 ;
  assign n54485 = ~n53053 & n54484 ;
  assign n54486 = ~n54482 & n54485 ;
  assign n54487 = \pi1150  & n54081 ;
  assign n54488 = n54486 & n54487 ;
  assign n54489 = ~n54481 & ~n54488 ;
  assign n54490 = n52665 & ~n54479 ;
  assign n54491 = ~\pi0214  & ~n52081 ;
  assign n54492 = \pi0212  & ~n54491 ;
  assign n54493 = ~n52952 & n52953 ;
  assign n54494 = \pi0211  & ~n54493 ;
  assign n54495 = n52657 & ~n54494 ;
  assign n54496 = ~n54479 & ~n54495 ;
  assign n54497 = n54492 & n54496 ;
  assign n54498 = ~n54490 & ~n54497 ;
  assign n54499 = \pi1150  & n54106 ;
  assign n54500 = n54498 & n54499 ;
  assign n54501 = n54489 & ~n54500 ;
  assign n54502 = ~n52707 & n52725 ;
  assign n54503 = ~n52702 & ~n54502 ;
  assign n54504 = ~\pi1150  & ~n54062 ;
  assign n54505 = n54068 & n54504 ;
  assign n54506 = n54106 & n54505 ;
  assign n54507 = ~n54503 & n54506 ;
  assign n54508 = n52706 & n52709 ;
  assign n54509 = ~n54401 & ~n54508 ;
  assign n54510 = n52617 & ~n52707 ;
  assign n54511 = n52001 & n54181 ;
  assign n54512 = ~n50679 & n54511 ;
  assign n54513 = ~n54510 & ~n54512 ;
  assign n54514 = ~n54509 & n54513 ;
  assign n54515 = ~\pi1150  & n54069 ;
  assign n54516 = ~n54514 & n54515 ;
  assign n54517 = \pi1148  & ~n54516 ;
  assign n54518 = ~n54507 & n54517 ;
  assign n54519 = n54501 & n54518 ;
  assign n54520 = \pi1150  & n12691 ;
  assign n54521 = n50877 & n54520 ;
  assign n54522 = n20516 & n54521 ;
  assign n54523 = n54105 & ~n54459 ;
  assign n54524 = ~n54522 & n54523 ;
  assign n54525 = ~n54401 & ~n54522 ;
  assign n54526 = ~n54111 & n54525 ;
  assign n54527 = ~n54524 & ~n54526 ;
  assign n54528 = ~\pi1146  & ~n50443 ;
  assign n54529 = n53008 & ~n54528 ;
  assign n54530 = ~\pi0299  & \pi1150  ;
  assign n54531 = n12691 & n54530 ;
  assign n54532 = n50877 & n54531 ;
  assign n54533 = n50556 & n52001 ;
  assign n54534 = ~\pi0219  & ~n54533 ;
  assign n54535 = ~n54532 & n54534 ;
  assign n54536 = ~n54529 & n54535 ;
  assign n54537 = ~n54111 & n54536 ;
  assign n54538 = ~\pi1148  & ~n54537 ;
  assign n54539 = n54527 & n54538 ;
  assign n54540 = ~\pi1149  & ~n54539 ;
  assign n54541 = ~n54519 & n54540 ;
  assign n54542 = ~\pi0213  & ~n54541 ;
  assign n54543 = ~n54478 & n54542 ;
  assign n54544 = ~n52420 & ~n54543 ;
  assign n54545 = ~\pi0209  & ~n54297 ;
  assign n54546 = ~n54295 & n54545 ;
  assign n54547 = ~n54246 & n54546 ;
  assign n54548 = \pi0230  & ~n54547 ;
  assign n54549 = ~n54544 & n54548 ;
  assign n54550 = ~\pi0230  & \pi0246  ;
  assign n54551 = ~\pi0219  & ~n54273 ;
  assign n54552 = ~n54271 & n54551 ;
  assign n54553 = n50571 & ~n54173 ;
  assign n54554 = n54280 & ~n54553 ;
  assign n54555 = n6848 & ~n54554 ;
  assign n54556 = ~n54552 & n54555 ;
  assign n54557 = n54321 & ~n54556 ;
  assign n54558 = n6848 & ~n50948 ;
  assign n54559 = n54287 & n54558 ;
  assign n54560 = ~n54214 & n54559 ;
  assign n54561 = n50714 & ~n54315 ;
  assign n54562 = n52557 & ~n54561 ;
  assign n54563 = ~n54560 & n54562 ;
  assign n54564 = ~\pi0057  & ~n54563 ;
  assign n54565 = ~n54557 & n54564 ;
  assign n54566 = ~n50714 & ~n54565 ;
  assign n54567 = n54322 & n54552 ;
  assign n54568 = n54322 & n54554 ;
  assign n54569 = ~n54567 & ~n54568 ;
  assign n54570 = n6848 & ~n54560 ;
  assign n54571 = n54562 & n54570 ;
  assign n54572 = \pi1150  & ~n54571 ;
  assign n54573 = n54569 & n54572 ;
  assign n54574 = ~n54566 & n54573 ;
  assign n54575 = \pi0219  & ~\pi0299  ;
  assign n54576 = ~n54207 & n54575 ;
  assign n54577 = ~n54205 & n54576 ;
  assign n54578 = ~n54213 & n54577 ;
  assign n54579 = ~n50571 & n53974 ;
  assign n54580 = ~\pi1150  & ~n54579 ;
  assign n54581 = n52558 & n54580 ;
  assign n54582 = ~n54578 & n54581 ;
  assign n54583 = \pi0214  & n54238 ;
  assign n54584 = ~n54315 & n54583 ;
  assign n54585 = ~n52001 & ~n54229 ;
  assign n54586 = ~n54584 & n54585 ;
  assign n54587 = \pi0212  & ~n54586 ;
  assign n54588 = ~\pi0219  & ~n52001 ;
  assign n54589 = ~n54229 & n54588 ;
  assign n54590 = ~n52661 & ~n54589 ;
  assign n54591 = ~n54250 & ~n54590 ;
  assign n54592 = ~n54587 & n54591 ;
  assign n54593 = n54582 & ~n54592 ;
  assign n54594 = \pi1149  & \pi1150  ;
  assign n54595 = ~n53200 & n54321 ;
  assign n54596 = ~n54552 & n54595 ;
  assign n54597 = n54555 & n54596 ;
  assign n54598 = \pi1149  & ~n52641 ;
  assign n54599 = ~n54597 & n54598 ;
  assign n54600 = ~n54594 & ~n54599 ;
  assign n54601 = ~n54593 & ~n54600 ;
  assign n54602 = ~n54574 & n54601 ;
  assign n54603 = n52699 & ~n54229 ;
  assign n54604 = ~n54250 & n54603 ;
  assign n54605 = \pi0212  & ~n54604 ;
  assign n54606 = n54260 & n54605 ;
  assign n54607 = n54256 & ~n54606 ;
  assign n54608 = n52558 & ~n54579 ;
  assign n54609 = ~n54578 & n54608 ;
  assign n54610 = n54322 & ~n54554 ;
  assign n54611 = n52699 & ~n54172 ;
  assign n54612 = \pi0212  & ~n54611 ;
  assign n54613 = n54269 & n54612 ;
  assign n54614 = ~\pi0212  & ~n54166 ;
  assign n54615 = ~n54148 & n54614 ;
  assign n54616 = ~\pi0219  & ~n54615 ;
  assign n54617 = ~n54613 & n54616 ;
  assign n54618 = n54610 & ~n54617 ;
  assign n54619 = ~\pi1150  & ~n52233 ;
  assign n54620 = n53184 & ~n54250 ;
  assign n54621 = n54609 & ~n54620 ;
  assign n54622 = n54619 & ~n54621 ;
  assign n54623 = ~n54618 & n54622 ;
  assign n54624 = n54609 & ~n54623 ;
  assign n54625 = ~n54607 & n54624 ;
  assign n54626 = ~\pi1149  & n54623 ;
  assign n54627 = ~\pi0214  & n54175 ;
  assign n54628 = n54612 & ~n54627 ;
  assign n54629 = ~\pi0212  & n54269 ;
  assign n54630 = ~n54175 & n54629 ;
  assign n54631 = ~\pi0219  & ~n54630 ;
  assign n54632 = ~n54628 & n54631 ;
  assign n54633 = n54610 & ~n54632 ;
  assign n54634 = \pi1150  & ~n52513 ;
  assign n54635 = ~\pi1149  & n54634 ;
  assign n54636 = ~n54633 & n54635 ;
  assign n54637 = ~n54626 & ~n54636 ;
  assign n54638 = ~n54625 & ~n54637 ;
  assign n54639 = \pi1148  & ~n54638 ;
  assign n54640 = ~n54602 & n54639 ;
  assign n54641 = \pi1150  & ~n52229 ;
  assign n54642 = ~\pi0219  & \pi1147  ;
  assign n54643 = n50936 & ~n54143 ;
  assign n54644 = \pi0219  & n54139 ;
  assign n54645 = ~n54643 & ~n54644 ;
  assign n54646 = \pi1147  & ~n54645 ;
  assign n54647 = n9948 & ~n54646 ;
  assign n54648 = ~n54642 & n54647 ;
  assign n54649 = \pi0212  & ~n54156 ;
  assign n54650 = ~n54192 & n54649 ;
  assign n54651 = n12255 & n54175 ;
  assign n54652 = ~n54650 & ~n54651 ;
  assign n54653 = n54151 & n54164 ;
  assign n54654 = n54647 & ~n54653 ;
  assign n54655 = n54652 & n54654 ;
  assign n54656 = ~n54648 & ~n54655 ;
  assign n54657 = n54641 & n54656 ;
  assign n54658 = \pi0219  & n54229 ;
  assign n54659 = ~\pi0214  & n54229 ;
  assign n54660 = ~\pi0212  & ~n54659 ;
  assign n54661 = ~n54584 & n54660 ;
  assign n54662 = ~n54230 & ~n54661 ;
  assign n54663 = ~n54658 & ~n54662 ;
  assign n54664 = ~\pi0211  & ~n54355 ;
  assign n54665 = \pi0214  & ~n54235 ;
  assign n54666 = ~n54664 & n54665 ;
  assign n54667 = ~\pi0214  & n54238 ;
  assign n54668 = ~n54315 & n54667 ;
  assign n54669 = \pi0212  & ~n54668 ;
  assign n54670 = ~n54658 & n54669 ;
  assign n54671 = ~n54666 & n54670 ;
  assign n54672 = ~n54663 & ~n54671 ;
  assign n54673 = ~\pi1147  & n54641 ;
  assign n54674 = ~n54672 & n54673 ;
  assign n54675 = ~n54657 & ~n54674 ;
  assign n54676 = \pi1147  & n54139 ;
  assign n54677 = \pi1147  & ~n50877 ;
  assign n54678 = ~n54143 & n54677 ;
  assign n54679 = ~n54676 & ~n54678 ;
  assign n54680 = ~\pi0211  & \pi1150  ;
  assign n54681 = ~\pi0219  & n54680 ;
  assign n54682 = n50679 & n54681 ;
  assign n54683 = n27408 & ~n54682 ;
  assign n54684 = n54229 & n54683 ;
  assign n54685 = ~n54322 & ~n54684 ;
  assign n54686 = n54679 & ~n54685 ;
  assign n54687 = ~\pi1149  & ~n54686 ;
  assign n54688 = ~\pi1148  & ~n54687 ;
  assign n54689 = ~\pi1148  & n54682 ;
  assign n54690 = ~n20516 & n54689 ;
  assign n54691 = ~\pi1147  & n54238 ;
  assign n54692 = n54689 & n54691 ;
  assign n54693 = ~n54234 & n54692 ;
  assign n54694 = ~n54690 & ~n54693 ;
  assign n54695 = ~n54688 & n54694 ;
  assign n54696 = n52558 & ~n54230 ;
  assign n54697 = \pi0219  & n54696 ;
  assign n54698 = n52280 & ~n54229 ;
  assign n54699 = ~n12255 & ~n54698 ;
  assign n54700 = ~n54665 & ~n54699 ;
  assign n54701 = ~\pi0211  & ~n54699 ;
  assign n54702 = ~n54355 & n54701 ;
  assign n54703 = ~n54700 & ~n54702 ;
  assign n54704 = \pi0214  & n52001 ;
  assign n54705 = ~\pi0212  & ~n54704 ;
  assign n54706 = ~n54229 & n54705 ;
  assign n54707 = n54696 & ~n54706 ;
  assign n54708 = n54703 & n54707 ;
  assign n54709 = ~n54697 & ~n54708 ;
  assign n54710 = n54322 & n54645 ;
  assign n54711 = ~n54152 & n54710 ;
  assign n54712 = ~n54179 & n54711 ;
  assign n54713 = \pi0219  & n54322 ;
  assign n54714 = ~n54139 & n54713 ;
  assign n54715 = ~n54148 & n54714 ;
  assign n54716 = ~\pi1150  & ~n52631 ;
  assign n54717 = ~n54715 & n54716 ;
  assign n54718 = ~n54712 & n54717 ;
  assign n54719 = n54709 & n54718 ;
  assign n54720 = ~n54695 & ~n54719 ;
  assign n54721 = n54675 & n54720 ;
  assign n54722 = ~\pi1149  & ~n54694 ;
  assign n54723 = ~\pi1148  & ~\pi1149  ;
  assign n54724 = n54686 & n54723 ;
  assign n54725 = ~n54722 & ~n54724 ;
  assign n54726 = ~\pi0209  & n54725 ;
  assign n54727 = ~n54721 & n54726 ;
  assign n54728 = ~n54640 & n54727 ;
  assign n54729 = ~\pi1149  & \pi1150  ;
  assign n54730 = ~n52683 & n54729 ;
  assign n54731 = \pi1149  & ~n54641 ;
  assign n54732 = \pi1149  & ~n53392 ;
  assign n54733 = ~n52789 & n54732 ;
  assign n54734 = ~n54731 & ~n54733 ;
  assign n54735 = ~n54730 & n54734 ;
  assign n54736 = ~\pi1148  & n54735 ;
  assign n54737 = ~n52631 & ~n52743 ;
  assign n54738 = ~n52631 & ~n52768 ;
  assign n54739 = ~n52765 & n54738 ;
  assign n54740 = ~n54737 & ~n54739 ;
  assign n54741 = ~\pi1148  & ~\pi1150  ;
  assign n54742 = ~n54740 & n54741 ;
  assign n54743 = ~n54736 & ~n54742 ;
  assign n54744 = \pi0209  & ~n54743 ;
  assign n54745 = ~\pi1149  & ~n54619 ;
  assign n54746 = ~n52724 & ~n52727 ;
  assign n54747 = ~\pi1149  & n54746 ;
  assign n54748 = n52715 & n54747 ;
  assign n54749 = ~n54745 & ~n54748 ;
  assign n54750 = ~n52641 & ~n52709 ;
  assign n54751 = ~n52734 & n54750 ;
  assign n54752 = ~\pi1150  & n54751 ;
  assign n54753 = \pi1150  & ~n52621 ;
  assign n54754 = n52800 & n54753 ;
  assign n54755 = \pi1149  & ~n54754 ;
  assign n54756 = ~n54752 & n54755 ;
  assign n54757 = n54749 & ~n54756 ;
  assign n54758 = n54634 & ~n54756 ;
  assign n54759 = ~n52677 & n54758 ;
  assign n54760 = ~n54757 & ~n54759 ;
  assign n54761 = \pi0209  & \pi1148  ;
  assign n54762 = ~n54760 & n54761 ;
  assign n54763 = ~n54744 & ~n54762 ;
  assign n54764 = n52811 & n54763 ;
  assign n54765 = ~n54728 & n54764 ;
  assign n54766 = ~n54550 & ~n54765 ;
  assign n54767 = ~n54549 & n54766 ;
  assign n54768 = ~n52677 & n53338 ;
  assign n54769 = \pi1147  & ~n54768 ;
  assign n54770 = n53060 & n53171 ;
  assign n54771 = n9948 & ~n54770 ;
  assign n54772 = ~n52675 & n54771 ;
  assign n54773 = ~n52669 & n54772 ;
  assign n54774 = n53344 & ~n54773 ;
  assign n54775 = n54769 & ~n54774 ;
  assign n54776 = ~n52005 & n53184 ;
  assign n54777 = n9948 & ~n54776 ;
  assign n54778 = ~n53033 & n54777 ;
  assign n54779 = n53344 & ~n54778 ;
  assign n54780 = n9948 & ~n12255 ;
  assign n54781 = ~n52304 & n54780 ;
  assign n54782 = n52007 & n54781 ;
  assign n54783 = n53338 & ~n54782 ;
  assign n54784 = ~n54778 & n54783 ;
  assign n54785 = ~\pi1147  & ~n54784 ;
  assign n54786 = ~n54779 & n54785 ;
  assign n54787 = n54741 & ~n54786 ;
  assign n54788 = ~n54775 & n54787 ;
  assign n54789 = \pi0212  & ~n52654 ;
  assign n54790 = n54485 & ~n54789 ;
  assign n54791 = n9948 & ~n54790 ;
  assign n54792 = ~n52675 & n54791 ;
  assign n54793 = n53318 & ~n54792 ;
  assign n54794 = \pi1147  & ~n54793 ;
  assign n54795 = n53285 & ~n54772 ;
  assign n54796 = n54794 & ~n54795 ;
  assign n54797 = n52007 & n53391 ;
  assign n54798 = n53318 & ~n54797 ;
  assign n54799 = ~\pi1147  & ~n53285 ;
  assign n54800 = ~n54798 & n54799 ;
  assign n54801 = n52792 & ~n53033 ;
  assign n54802 = ~n53061 & n54801 ;
  assign n54803 = \pi1150  & ~n54802 ;
  assign n54804 = ~n54800 & n54803 ;
  assign n54805 = ~\pi1148  & n54804 ;
  assign n54806 = ~n54796 & n54805 ;
  assign n54807 = ~n53090 & n53285 ;
  assign n54808 = n53285 & n54408 ;
  assign n54809 = ~n54405 & n54808 ;
  assign n54810 = ~n54807 & ~n54809 ;
  assign n54811 = ~\pi0219  & ~n52783 ;
  assign n54812 = ~n52779 & n54811 ;
  assign n54813 = n53090 & ~n54812 ;
  assign n54814 = n53318 & ~n54813 ;
  assign n54815 = ~\pi1147  & ~n54814 ;
  assign n54816 = n54810 & n54815 ;
  assign n54817 = \pi1147  & ~n53403 ;
  assign n54818 = ~n53201 & n53285 ;
  assign n54819 = n54817 & ~n54818 ;
  assign n54820 = \pi1150  & ~n54819 ;
  assign n54821 = ~n54816 & n54820 ;
  assign n54822 = \pi1148  & n54821 ;
  assign n54823 = n53090 & ~n54426 ;
  assign n54824 = ~n54409 & n54823 ;
  assign n54825 = n53344 & ~n54824 ;
  assign n54826 = ~\pi1147  & ~n53338 ;
  assign n54827 = ~\pi1147  & n53090 ;
  assign n54828 = ~n54426 & n54827 ;
  assign n54829 = ~n54826 & ~n54828 ;
  assign n54830 = ~n54825 & ~n54829 ;
  assign n54831 = n53187 & n53338 ;
  assign n54832 = ~n52799 & ~n53186 ;
  assign n54833 = n53344 & n54832 ;
  assign n54834 = \pi1147  & ~n54833 ;
  assign n54835 = ~n54831 & n54834 ;
  assign n54836 = ~\pi1150  & ~n54835 ;
  assign n54837 = \pi1148  & n54836 ;
  assign n54838 = ~n54830 & n54837 ;
  assign n54839 = ~n54822 & ~n54838 ;
  assign n54840 = ~n54806 & n54839 ;
  assign n54841 = ~n54788 & n54840 ;
  assign n54842 = \pi1149  & n54841 ;
  assign n54843 = ~n50701 & ~n52707 ;
  assign n54844 = ~n50679 & ~n52692 ;
  assign n54845 = n51975 & n54844 ;
  assign n54846 = n9948 & ~n54845 ;
  assign n54847 = ~n54843 & n54846 ;
  assign n54848 = n53230 & ~n54847 ;
  assign n54849 = \pi1147  & ~n54848 ;
  assign n54850 = ~\pi0219  & ~n20516 ;
  assign n54851 = ~n52630 & n54850 ;
  assign n54852 = ~\pi1151  & ~n54851 ;
  assign n54853 = ~n20516 & n51169 ;
  assign n54854 = \pi1151  & ~n54853 ;
  assign n54855 = ~\pi1147  & ~n54854 ;
  assign n54856 = ~n54852 & n54855 ;
  assign n54857 = \pi1150  & ~n54856 ;
  assign n54858 = ~n54849 & n54857 ;
  assign n54859 = \pi0219  & ~n52707 ;
  assign n54860 = n9948 & ~n54859 ;
  assign n54861 = ~\pi0219  & ~n52723 ;
  assign n54862 = ~n54502 & ~n54861 ;
  assign n54863 = n54860 & n54862 ;
  assign n54864 = n53275 & n54857 ;
  assign n54865 = ~n54863 & n54864 ;
  assign n54866 = ~n54858 & ~n54865 ;
  assign n54867 = ~n52827 & ~n53150 ;
  assign n54868 = ~n52707 & n54867 ;
  assign n54869 = ~n53362 & ~n54868 ;
  assign n54870 = \pi1147  & \pi1151  ;
  assign n54871 = \pi1147  & n52706 ;
  assign n54872 = n52709 & n54871 ;
  assign n54873 = ~n54870 & ~n54872 ;
  assign n54874 = n54869 & ~n54873 ;
  assign n54875 = ~\pi1147  & \pi1151  ;
  assign n54876 = n12577 & n54875 ;
  assign n54877 = n50679 & n54876 ;
  assign n54878 = ~n20516 & n54877 ;
  assign n54879 = ~\pi1150  & ~n54878 ;
  assign n54880 = ~n54874 & n54879 ;
  assign n54881 = n54723 & ~n54880 ;
  assign n54882 = n54866 & n54881 ;
  assign n54883 = ~n53362 & n54875 ;
  assign n54884 = n52558 & ~n53362 ;
  assign n54885 = n52741 & n54884 ;
  assign n54886 = ~n54883 & ~n54885 ;
  assign n54887 = ~\pi1150  & n54886 ;
  assign n54888 = n9948 & ~n53126 ;
  assign n54889 = n52750 & n53123 ;
  assign n54890 = ~\pi1150  & ~n54889 ;
  assign n54891 = n54888 & n54890 ;
  assign n54892 = ~n54887 & ~n54891 ;
  assign n54893 = ~\pi1149  & n54892 ;
  assign n54894 = \pi1151  & ~n52827 ;
  assign n54895 = ~n53213 & n54894 ;
  assign n54896 = ~n52695 & n54894 ;
  assign n54897 = ~n54451 & n54896 ;
  assign n54898 = ~n54895 & ~n54897 ;
  assign n54899 = \pi1147  & n9948 ;
  assign n54900 = ~n51975 & n54899 ;
  assign n54901 = ~n54870 & ~n54900 ;
  assign n54902 = ~\pi1149  & ~n54901 ;
  assign n54903 = n54898 & n54902 ;
  assign n54904 = ~n54893 & ~n54903 ;
  assign n54905 = \pi1148  & ~n54904 ;
  assign n54906 = ~\pi1147  & ~n53230 ;
  assign n54907 = ~\pi1147  & n52743 ;
  assign n54908 = n52760 & n54907 ;
  assign n54909 = ~n54906 & ~n54908 ;
  assign n54910 = n53389 & ~n54909 ;
  assign n54911 = \pi1147  & ~n53275 ;
  assign n54912 = \pi1147  & n53213 ;
  assign n54913 = ~n54861 & n54912 ;
  assign n54914 = ~n54911 & ~n54913 ;
  assign n54915 = \pi1150  & n54914 ;
  assign n54916 = ~n52695 & ~n54451 ;
  assign n54917 = n53213 & ~n54916 ;
  assign n54918 = ~n53213 & n53230 ;
  assign n54919 = ~\pi0219  & n53230 ;
  assign n54920 = ~n52723 & n54919 ;
  assign n54921 = ~n54918 & ~n54920 ;
  assign n54922 = \pi1150  & ~n54921 ;
  assign n54923 = ~n54917 & n54922 ;
  assign n54924 = ~n54915 & ~n54923 ;
  assign n54925 = ~n54910 & ~n54924 ;
  assign n54926 = n54905 & ~n54925 ;
  assign n54927 = ~n54882 & ~n54926 ;
  assign n54928 = ~n54842 & n54927 ;
  assign n54929 = \pi0213  & ~n54928 ;
  assign n54930 = ~\pi0213  & ~n52809 ;
  assign n54931 = ~\pi0209  & ~n54930 ;
  assign n54932 = \pi0230  & n54931 ;
  assign n54933 = ~n54929 & n54932 ;
  assign n54934 = ~\pi0230  & ~\pi0247  ;
  assign n54935 = ~\pi1151  & ~n52827 ;
  assign n54936 = ~n52695 & n54935 ;
  assign n54937 = ~n54451 & n54936 ;
  assign n54938 = ~n53213 & n54935 ;
  assign n54939 = ~n53018 & n54894 ;
  assign n54940 = ~\pi1147  & ~n54939 ;
  assign n54941 = ~n54938 & n54940 ;
  assign n54942 = ~n54937 & n54941 ;
  assign n54943 = \pi1150  & n54942 ;
  assign n54944 = ~n52513 & n52713 ;
  assign n54945 = ~n52513 & ~n52695 ;
  assign n54946 = ~n52701 & n54945 ;
  assign n54947 = ~n54944 & ~n54946 ;
  assign n54948 = ~\pi1151  & ~n54947 ;
  assign n54949 = \pi1147  & ~n54831 ;
  assign n54950 = \pi1150  & n54949 ;
  assign n54951 = ~n54948 & n54950 ;
  assign n54952 = ~n54943 & ~n54951 ;
  assign n54953 = ~\pi1148  & \pi1150  ;
  assign n54954 = ~\pi1151  & ~n52513 ;
  assign n54955 = ~n52714 & n54954 ;
  assign n54956 = ~n52695 & n54954 ;
  assign n54957 = ~n52701 & n54956 ;
  assign n54958 = ~n54955 & ~n54957 ;
  assign n54959 = \pi1147  & n54958 ;
  assign n54960 = ~\pi1147  & ~n54935 ;
  assign n54961 = ~n54894 & n54960 ;
  assign n54962 = n52558 & ~n54894 ;
  assign n54963 = ~n53151 & n54962 ;
  assign n54964 = ~n54961 & ~n54963 ;
  assign n54965 = ~n54959 & n54964 ;
  assign n54966 = n53338 & n54964 ;
  assign n54967 = ~n52677 & n54966 ;
  assign n54968 = ~n54965 & ~n54967 ;
  assign n54969 = n52558 & ~n53151 ;
  assign n54970 = ~n54960 & ~n54969 ;
  assign n54971 = n52975 & ~n54970 ;
  assign n54972 = ~n52668 & n54971 ;
  assign n54973 = ~\pi1148  & ~n54972 ;
  assign n54974 = ~n54968 & n54973 ;
  assign n54975 = ~n54953 & ~n54974 ;
  assign n54976 = n54952 & ~n54975 ;
  assign n54977 = ~\pi1151  & ~n52229 ;
  assign n54978 = ~n53213 & n54977 ;
  assign n54979 = ~\pi0219  & n54977 ;
  assign n54980 = ~n52723 & n54979 ;
  assign n54981 = ~n54978 & ~n54980 ;
  assign n54982 = n53230 & ~n54463 ;
  assign n54983 = ~\pi1147  & \pi1150  ;
  assign n54984 = ~n54982 & n54983 ;
  assign n54985 = n54981 & n54984 ;
  assign n54986 = n53213 & n54984 ;
  assign n54987 = ~n54916 & n54986 ;
  assign n54988 = ~n54985 & ~n54987 ;
  assign n54989 = ~\pi1151  & ~n52709 ;
  assign n54990 = ~n52621 & ~n52733 ;
  assign n54991 = n54989 & n54990 ;
  assign n54992 = \pi1150  & ~n54991 ;
  assign n54993 = n54817 & n54992 ;
  assign n54994 = \pi1148  & ~n54993 ;
  assign n54995 = n54988 & n54994 ;
  assign n54996 = \pi1149  & ~n54995 ;
  assign n54997 = n52975 & ~n54485 ;
  assign n54998 = n52975 & n53253 ;
  assign n54999 = ~n52672 & n54998 ;
  assign n55000 = ~n54997 & ~n54999 ;
  assign n55001 = n53230 & n55000 ;
  assign n55002 = ~n54847 & n54977 ;
  assign n55003 = ~\pi1147  & ~n55002 ;
  assign n55004 = ~n55001 & n55003 ;
  assign n55005 = n53356 & n55004 ;
  assign n55006 = \pi1147  & n52714 ;
  assign n55007 = ~n52702 & n55006 ;
  assign n55008 = ~\pi1151  & ~n52621 ;
  assign n55009 = ~n54847 & n55008 ;
  assign n55010 = \pi1147  & ~n55009 ;
  assign n55011 = ~n55007 & ~n55010 ;
  assign n55012 = n53356 & ~n55011 ;
  assign n55013 = ~n54793 & n55012 ;
  assign n55014 = ~n55005 & ~n55013 ;
  assign n55015 = ~n54996 & n55014 ;
  assign n55016 = ~\pi0213  & ~n55015 ;
  assign n55017 = ~n54976 & n55016 ;
  assign n55018 = \pi1151  & ~n52641 ;
  assign n55019 = \pi1147  & ~n55018 ;
  assign n55020 = ~n52985 & n54899 ;
  assign n55021 = ~n55019 & ~n55020 ;
  assign n55022 = n54408 & ~n55019 ;
  assign n55023 = ~n54405 & n55022 ;
  assign n55024 = ~n55021 & ~n55023 ;
  assign n55025 = ~n52641 & ~n52768 ;
  assign n55026 = ~n52764 & n55025 ;
  assign n55027 = ~n52641 & ~n54393 ;
  assign n55028 = ~n52743 & n55027 ;
  assign n55029 = \pi1150  & ~n55028 ;
  assign n55030 = ~n55026 & n55029 ;
  assign n55031 = ~n53189 & ~n55030 ;
  assign n55032 = n55024 & ~n55031 ;
  assign n55033 = ~\pi1147  & n53389 ;
  assign n55034 = \pi1151  & ~n52631 ;
  assign n55035 = ~\pi0219  & n54417 ;
  assign n55036 = ~n54405 & n55035 ;
  assign n55037 = ~n53392 & ~n55036 ;
  assign n55038 = n55034 & ~n55037 ;
  assign n55039 = \pi1150  & ~n55038 ;
  assign n55040 = n55033 & n55039 ;
  assign n55041 = ~n55032 & ~n55040 ;
  assign n55042 = ~\pi1147  & ~n54852 ;
  assign n55043 = ~n53391 & n55034 ;
  assign n55044 = ~n53268 & n55034 ;
  assign n55045 = n53265 & n55044 ;
  assign n55046 = ~n55043 & ~n55045 ;
  assign n55047 = n55042 & n55046 ;
  assign n55048 = ~n53062 & n55018 ;
  assign n55049 = \pi1147  & ~n53401 ;
  assign n55050 = ~n55048 & n55049 ;
  assign n55051 = ~n55047 & ~n55050 ;
  assign n55052 = ~\pi1150  & ~n55051 ;
  assign n55053 = \pi1148  & ~n55052 ;
  assign n55054 = n55041 & n55053 ;
  assign n55055 = n52234 & ~n54824 ;
  assign n55056 = ~n52233 & ~n54433 ;
  assign n55057 = ~n52233 & ~n54393 ;
  assign n55058 = ~n52743 & n55057 ;
  assign n55059 = ~n55056 & ~n55058 ;
  assign n55060 = ~\pi1151  & ~n55059 ;
  assign n55061 = \pi1147  & ~n55060 ;
  assign n55062 = ~n55055 & n55061 ;
  assign n55063 = \pi1151  & ~n52790 ;
  assign n55064 = \pi1150  & n55063 ;
  assign n55065 = n52558 & n52741 ;
  assign n55066 = \pi1150  & ~n54875 ;
  assign n55067 = ~n55065 & n55066 ;
  assign n55068 = ~n55064 & ~n55067 ;
  assign n55069 = ~\pi1148  & ~n55068 ;
  assign n55070 = ~n55062 & n55069 ;
  assign n55071 = n52234 & ~n54778 ;
  assign n55072 = ~n53186 & n53344 ;
  assign n55073 = \pi1147  & ~n55072 ;
  assign n55074 = ~n55071 & n55073 ;
  assign n55075 = n12691 & n54875 ;
  assign n55076 = n50877 & n55075 ;
  assign n55077 = n20516 & n55076 ;
  assign n55078 = ~\pi1150  & ~n55077 ;
  assign n55079 = ~\pi1148  & n55078 ;
  assign n55080 = ~n55074 & n55079 ;
  assign n55081 = ~\pi1149  & ~n55080 ;
  assign n55082 = ~n55070 & n55081 ;
  assign n55083 = ~\pi0213  & n55082 ;
  assign n55084 = ~n55054 & n55083 ;
  assign n55085 = \pi0213  & ~n53417 ;
  assign n55086 = ~n53408 & n55085 ;
  assign n55087 = ~n53400 & n55086 ;
  assign n55088 = \pi0209  & ~n55087 ;
  assign n55089 = \pi0230  & n55088 ;
  assign n55090 = ~n55084 & n55089 ;
  assign n55091 = ~n55017 & n55090 ;
  assign n55092 = ~n54934 & ~n55091 ;
  assign n55093 = ~n54933 & n55092 ;
  assign n55094 = \pi1152  & ~n53403 ;
  assign n55095 = ~n54792 & n55008 ;
  assign n55096 = n55094 & ~n55095 ;
  assign n55097 = \pi1151  & ~n52709 ;
  assign n55098 = n54990 & n55097 ;
  assign n55099 = ~\pi1152  & ~n55098 ;
  assign n55100 = \pi1150  & ~n55099 ;
  assign n55101 = \pi1150  & n55009 ;
  assign n55102 = ~n52715 & n55101 ;
  assign n55103 = ~n55100 & ~n55102 ;
  assign n55104 = ~n55096 & ~n55103 ;
  assign n55105 = ~\pi1152  & ~n53401 ;
  assign n55106 = ~\pi1151  & n55105 ;
  assign n55107 = ~n55028 & n55105 ;
  assign n55108 = ~n55026 & n55107 ;
  assign n55109 = ~n55106 & ~n55108 ;
  assign n55110 = \pi1148  & \pi1149  ;
  assign n55111 = ~n55109 & n55110 ;
  assign n55112 = ~\pi1150  & ~n53090 ;
  assign n55113 = ~\pi1150  & n54408 ;
  assign n55114 = ~n54405 & n55113 ;
  assign n55115 = ~n55112 & ~n55114 ;
  assign n55116 = n55018 & ~n55115 ;
  assign n55117 = ~\pi1150  & ~\pi1152  ;
  assign n55118 = ~\pi1150  & n53285 ;
  assign n55119 = ~n53062 & n55118 ;
  assign n55120 = ~n55117 & ~n55119 ;
  assign n55121 = n55110 & n55120 ;
  assign n55122 = ~n55116 & n55121 ;
  assign n55123 = ~n55111 & ~n55122 ;
  assign n55124 = ~n55104 & ~n55123 ;
  assign n55125 = ~n52743 & n55034 ;
  assign n55126 = ~n52768 & n55034 ;
  assign n55127 = ~n52765 & n55126 ;
  assign n55128 = ~n55125 & ~n55127 ;
  assign n55129 = ~\pi1152  & ~n54852 ;
  assign n55130 = n55128 & n55129 ;
  assign n55131 = ~n53268 & n53275 ;
  assign n55132 = n53265 & n55131 ;
  assign n55133 = n53275 & ~n53391 ;
  assign n55134 = \pi1152  & ~n55133 ;
  assign n55135 = ~n55132 & n55134 ;
  assign n55136 = ~\pi1150  & ~n55135 ;
  assign n55137 = ~\pi1150  & n55034 ;
  assign n55138 = ~n55037 & n55137 ;
  assign n55139 = ~n55136 & ~n55138 ;
  assign n55140 = ~n55130 & ~n55139 ;
  assign n55141 = n53213 & ~n54861 ;
  assign n55142 = n53230 & ~n55141 ;
  assign n55143 = ~n54917 & n55142 ;
  assign n55144 = ~\pi1152  & ~n55002 ;
  assign n55145 = ~n55143 & n55144 ;
  assign n55146 = \pi1152  & ~n54982 ;
  assign n55147 = \pi1150  & ~n55146 ;
  assign n55148 = \pi1150  & n54977 ;
  assign n55149 = n55000 & n55148 ;
  assign n55150 = ~n55147 & ~n55149 ;
  assign n55151 = ~n55145 & ~n55150 ;
  assign n55152 = n52685 & ~n55151 ;
  assign n55153 = ~n55140 & n55152 ;
  assign n55154 = ~n55124 & ~n55153 ;
  assign n55155 = ~\pi0213  & ~n55154 ;
  assign n55156 = \pi1151  & ~n54947 ;
  assign n55157 = ~\pi1152  & n54958 ;
  assign n55158 = ~n55156 & n55157 ;
  assign n55159 = \pi1150  & n55158 ;
  assign n55160 = ~n52677 & n54954 ;
  assign n55161 = \pi1152  & ~n54831 ;
  assign n55162 = \pi1150  & n55161 ;
  assign n55163 = ~n55160 & n55162 ;
  assign n55164 = ~n55159 & ~n55163 ;
  assign n55165 = \pi1151  & ~n55059 ;
  assign n55166 = ~\pi1152  & ~n55072 ;
  assign n55167 = ~\pi1150  & n55166 ;
  assign n55168 = ~n55165 & n55167 ;
  assign n55169 = n53070 & ~n54779 ;
  assign n55170 = \pi1148  & ~n55169 ;
  assign n55171 = \pi1148  & n52234 ;
  assign n55172 = ~n54824 & n55171 ;
  assign n55173 = ~n55170 & ~n55172 ;
  assign n55174 = ~n55168 & ~n55173 ;
  assign n55175 = n55164 & n55174 ;
  assign n55176 = \pi1148  & ~\pi1149  ;
  assign n55177 = \pi1152  & ~n54935 ;
  assign n55178 = ~n54939 & n55177 ;
  assign n55179 = \pi1152  & n52975 ;
  assign n55180 = ~n54939 & n55179 ;
  assign n55181 = ~n52668 & n55180 ;
  assign n55182 = ~n55178 & ~n55181 ;
  assign n55183 = ~\pi1152  & ~n54935 ;
  assign n55184 = n51088 & ~n53151 ;
  assign n55185 = ~n55183 & ~n55184 ;
  assign n55186 = n54898 & ~n55185 ;
  assign n55187 = \pi1150  & ~n55186 ;
  assign n55188 = n55182 & n55187 ;
  assign n55189 = n9948 & n53117 ;
  assign n55190 = n52741 & n55189 ;
  assign n55191 = ~\pi0057  & n52250 ;
  assign n55192 = n6848 & n55191 ;
  assign n55193 = n51918 & n55192 ;
  assign n55194 = ~\pi1151  & \pi1152  ;
  assign n55195 = n12691 & n55194 ;
  assign n55196 = n50877 & n55195 ;
  assign n55197 = n20516 & n55196 ;
  assign n55198 = ~\pi1150  & ~n55197 ;
  assign n55199 = ~n55193 & n55198 ;
  assign n55200 = ~n55190 & n55199 ;
  assign n55201 = ~\pi1149  & ~n55200 ;
  assign n55202 = ~n55188 & n55201 ;
  assign n55203 = ~n55176 & ~n55202 ;
  assign n55204 = ~\pi0213  & ~n55203 ;
  assign n55205 = ~n55175 & n55204 ;
  assign n55206 = ~n55155 & ~n55205 ;
  assign n55207 = n55094 & ~n55160 ;
  assign n55208 = n52715 & n54746 ;
  assign n55209 = n53344 & ~n55208 ;
  assign n55210 = \pi1151  & n54751 ;
  assign n55211 = ~\pi1152  & ~n55210 ;
  assign n55212 = ~n55209 & n55211 ;
  assign n55213 = \pi1150  & ~n55212 ;
  assign n55214 = ~n55207 & n55213 ;
  assign n55215 = n53117 & n54740 ;
  assign n55216 = ~\pi1151  & ~n52682 ;
  assign n55217 = ~n52681 & n55216 ;
  assign n55218 = \pi1152  & ~n55217 ;
  assign n55219 = ~n53230 & n55218 ;
  assign n55220 = ~n53392 & n55218 ;
  assign n55221 = ~n52789 & n55220 ;
  assign n55222 = ~n55219 & ~n55221 ;
  assign n55223 = ~\pi1150  & n55222 ;
  assign n55224 = ~n55215 & n55223 ;
  assign n55225 = \pi0213  & ~n55224 ;
  assign n55226 = ~n55214 & n55225 ;
  assign n55227 = \pi0209  & ~n55226 ;
  assign n55228 = n55206 & n55227 ;
  assign n55229 = \pi0230  & n55228 ;
  assign n55230 = \pi1152  & ~n54793 ;
  assign n55231 = ~n55160 & n55230 ;
  assign n55232 = ~n54772 & n55018 ;
  assign n55233 = ~\pi1152  & ~n55232 ;
  assign n55234 = ~n54774 & n55233 ;
  assign n55235 = \pi1150  & ~n55234 ;
  assign n55236 = ~n55231 & n55235 ;
  assign n55237 = ~\pi1152  & n52706 ;
  assign n55238 = n52709 & n55237 ;
  assign n55239 = ~n53117 & ~n55238 ;
  assign n55240 = ~n55034 & ~n55239 ;
  assign n55241 = n54860 & ~n55239 ;
  assign n55242 = n54862 & n55241 ;
  assign n55243 = ~n55240 & ~n55242 ;
  assign n55244 = n50998 & ~n53151 ;
  assign n55245 = ~n55177 & ~n55244 ;
  assign n55246 = ~n54848 & ~n55245 ;
  assign n55247 = ~\pi1150  & ~n55246 ;
  assign n55248 = n55243 & n55247 ;
  assign n55249 = ~\pi1149  & ~n55248 ;
  assign n55250 = ~n55236 & n55249 ;
  assign n55251 = n53187 & n54954 ;
  assign n55252 = n55094 & ~n55251 ;
  assign n55253 = ~n53201 & n55018 ;
  assign n55254 = ~\pi1152  & ~n54833 ;
  assign n55255 = ~n55253 & n55254 ;
  assign n55256 = ~n55252 & ~n55255 ;
  assign n55257 = \pi1150  & n55256 ;
  assign n55258 = \pi1149  & ~n55257 ;
  assign n55259 = ~n54937 & ~n54938 ;
  assign n55260 = \pi1152  & n55259 ;
  assign n55261 = ~n55143 & n55260 ;
  assign n55262 = ~n53194 & n53213 ;
  assign n55263 = ~n54861 & n55262 ;
  assign n55264 = ~n53194 & ~n55034 ;
  assign n55265 = ~\pi1150  & ~n55264 ;
  assign n55266 = ~n55263 & n55265 ;
  assign n55267 = ~n55261 & n55266 ;
  assign n55268 = n55258 & ~n55267 ;
  assign n55269 = \pi1148  & ~n55268 ;
  assign n55270 = ~n55250 & n55269 ;
  assign n55271 = n52250 & n54853 ;
  assign n55272 = n52682 & n55194 ;
  assign n55273 = ~n55271 & ~n55272 ;
  assign n55274 = ~\pi0219  & n53117 ;
  assign n55275 = ~n20516 & n55274 ;
  assign n55276 = ~n52630 & n55275 ;
  assign n55277 = ~\pi1150  & ~n55276 ;
  assign n55278 = n55273 & n55277 ;
  assign n55279 = ~\pi1149  & ~n55278 ;
  assign n55280 = ~\pi1148  & ~n55279 ;
  assign n55281 = ~\pi1152  & ~n54779 ;
  assign n55282 = ~n55048 & n55281 ;
  assign n55283 = \pi1150  & ~n55282 ;
  assign n55284 = ~n53062 & n54798 ;
  assign n55285 = ~n54782 & n54954 ;
  assign n55286 = ~n54778 & n55285 ;
  assign n55287 = \pi1152  & ~n55286 ;
  assign n55288 = ~n55284 & n55287 ;
  assign n55289 = ~\pi1148  & ~n55288 ;
  assign n55290 = n55283 & n55289 ;
  assign n55291 = ~n55280 & ~n55290 ;
  assign n55292 = \pi0213  & n55291 ;
  assign n55293 = ~n53090 & n55018 ;
  assign n55294 = n54408 & n55018 ;
  assign n55295 = ~n54405 & n55294 ;
  assign n55296 = ~n55293 & ~n55295 ;
  assign n55297 = ~\pi1152  & n55296 ;
  assign n55298 = ~n54825 & n55297 ;
  assign n55299 = ~n54823 & n54954 ;
  assign n55300 = \pi1152  & ~n54814 ;
  assign n55301 = ~n55299 & n55300 ;
  assign n55302 = \pi1150  & ~n55301 ;
  assign n55303 = ~n55298 & n55302 ;
  assign n55304 = \pi1149  & ~n55303 ;
  assign n55305 = n52741 & n53192 ;
  assign n55306 = ~n53117 & ~n55305 ;
  assign n55307 = n55128 & ~n55306 ;
  assign n55308 = ~\pi1151  & ~n54889 ;
  assign n55309 = n54888 & n55308 ;
  assign n55310 = ~\pi1151  & n53362 ;
  assign n55311 = \pi1152  & ~n55310 ;
  assign n55312 = ~n55309 & n55311 ;
  assign n55313 = ~\pi1150  & ~n55312 ;
  assign n55314 = n52743 & n52760 ;
  assign n55315 = ~\pi1150  & n53230 ;
  assign n55316 = ~n55314 & n55315 ;
  assign n55317 = ~n55313 & ~n55316 ;
  assign n55318 = ~n55307 & ~n55317 ;
  assign n55319 = \pi0213  & ~n55318 ;
  assign n55320 = n55304 & n55319 ;
  assign n55321 = ~n55292 & ~n55320 ;
  assign n55322 = ~n55270 & ~n55321 ;
  assign n55323 = \pi1148  & ~n54760 ;
  assign n55324 = ~\pi0213  & n54743 ;
  assign n55325 = ~n55323 & n55324 ;
  assign n55326 = ~\pi0209  & ~n55325 ;
  assign n55327 = \pi0230  & n55326 ;
  assign n55328 = ~n55322 & n55327 ;
  assign n55329 = ~n55229 & ~n55328 ;
  assign n55330 = ~\pi0230  & ~\pi0248  ;
  assign n55331 = n55329 & ~n55330 ;
  assign n55332 = n50877 & n51088 ;
  assign n55333 = n51112 & n55332 ;
  assign n55334 = n51088 & n51116 ;
  assign n55335 = ~n53117 & ~n55334 ;
  assign n55336 = ~n55333 & n55335 ;
  assign n55337 = ~n55034 & ~n55336 ;
  assign n55338 = \pi0219  & ~n51116 ;
  assign n55339 = n9948 & ~n55338 ;
  assign n55340 = n9948 & n50877 ;
  assign n55341 = n51112 & n55340 ;
  assign n55342 = ~n55339 & ~n55341 ;
  assign n55343 = ~n55336 & ~n55342 ;
  assign n55344 = ~n55337 & ~n55343 ;
  assign n55345 = \pi0214  & n51117 ;
  assign n55346 = ~n51113 & n55345 ;
  assign n55347 = n50411 & ~n51399 ;
  assign n55348 = \pi0208  & ~n50544 ;
  assign n55349 = n12691 & n51115 ;
  assign n55350 = ~n55348 & ~n55349 ;
  assign n55351 = ~n51133 & n51880 ;
  assign n55352 = ~n51097 & n55351 ;
  assign n55353 = ~n55350 & ~n55352 ;
  assign n55354 = ~n55347 & ~n55353 ;
  assign n55355 = n50967 & n55354 ;
  assign n55356 = ~n55346 & ~n55355 ;
  assign n55357 = ~\pi0211  & n51115 ;
  assign n55358 = n51114 & n55357 ;
  assign n55359 = ~\pi0214  & ~n55358 ;
  assign n55360 = \pi0212  & ~n55359 ;
  assign n55361 = ~\pi0211  & n50877 ;
  assign n55362 = \pi0212  & n55361 ;
  assign n55363 = n51112 & n55362 ;
  assign n55364 = ~n55360 & ~n55363 ;
  assign n55365 = n54089 & ~n55354 ;
  assign n55366 = n55364 & ~n55365 ;
  assign n55367 = n55356 & ~n55366 ;
  assign n55368 = \pi1154  & ~n50430 ;
  assign n55369 = n51110 & n55368 ;
  assign n55370 = ~\pi1154  & ~n50430 ;
  assign n55371 = n51034 & n55370 ;
  assign n55372 = ~n55369 & ~n55371 ;
  assign n55373 = n50877 & ~n55372 ;
  assign n55374 = ~n50430 & n51115 ;
  assign n55375 = n51114 & n55374 ;
  assign n55376 = ~\pi0219  & ~n55375 ;
  assign n55377 = ~n55373 & n55376 ;
  assign n55378 = ~n52660 & ~n55377 ;
  assign n55379 = n50430 & ~n52660 ;
  assign n55380 = ~n55354 & n55379 ;
  assign n55381 = ~n55378 & ~n55380 ;
  assign n55382 = ~n55337 & n55381 ;
  assign n55383 = ~n55367 & n55382 ;
  assign n55384 = ~n55344 & ~n55383 ;
  assign n55385 = ~\pi1150  & n55384 ;
  assign n55386 = ~n51209 & n54954 ;
  assign n55387 = ~\pi0212  & n51243 ;
  assign n55388 = ~\pi0211  & ~n51203 ;
  assign n55389 = ~n51009 & n51198 ;
  assign n55390 = ~n51005 & n55389 ;
  assign n55391 = \pi0214  & ~n55390 ;
  assign n55392 = ~\pi0212  & n55391 ;
  assign n55393 = ~n55388 & n55392 ;
  assign n55394 = ~n55387 & ~n55393 ;
  assign n55395 = ~\pi0214  & n55390 ;
  assign n55396 = n50442 & ~n51203 ;
  assign n55397 = ~n55395 & ~n55396 ;
  assign n55398 = n50430 & ~n51203 ;
  assign n55399 = ~\pi0211  & ~n50876 ;
  assign n55400 = ~n51009 & n55399 ;
  assign n55401 = \pi0214  & ~n51005 ;
  assign n55402 = n55400 & n55401 ;
  assign n55403 = \pi0212  & ~n55402 ;
  assign n55404 = ~n55398 & n55403 ;
  assign n55405 = n55397 & n55404 ;
  assign n55406 = n55394 & ~n55405 ;
  assign n55407 = ~\pi0219  & n54954 ;
  assign n55408 = ~n55406 & n55407 ;
  assign n55409 = ~n55386 & ~n55408 ;
  assign n55410 = \pi1152  & ~n53318 ;
  assign n55411 = \pi0214  & n51203 ;
  assign n55412 = n51244 & ~n55411 ;
  assign n55413 = \pi0212  & ~n51203 ;
  assign n55414 = ~\pi0219  & ~n55413 ;
  assign n55415 = ~n55412 & n55414 ;
  assign n55416 = \pi1152  & ~n55415 ;
  assign n55417 = n51209 & n55416 ;
  assign n55418 = ~n55410 & ~n55417 ;
  assign n55419 = n55409 & ~n55418 ;
  assign n55420 = \pi1150  & n55419 ;
  assign n55421 = ~\pi0219  & ~n55412 ;
  assign n55422 = ~n55388 & n55391 ;
  assign n55423 = ~\pi0214  & n51203 ;
  assign n55424 = \pi0212  & ~n55423 ;
  assign n55425 = ~n55422 & n55424 ;
  assign n55426 = n55421 & ~n55425 ;
  assign n55427 = n9948 & ~n51206 ;
  assign n55428 = ~n55426 & n55427 ;
  assign n55429 = n53230 & ~n55428 ;
  assign n55430 = ~n51073 & ~n52212 ;
  assign n55431 = n53272 & ~n55430 ;
  assign n55432 = ~n55177 & ~n55431 ;
  assign n55433 = n52212 & ~n55390 ;
  assign n55434 = ~n55177 & n55433 ;
  assign n55435 = ~n55388 & n55434 ;
  assign n55436 = ~n55432 & ~n55435 ;
  assign n55437 = ~\pi1150  & n55436 ;
  assign n55438 = ~n55429 & n55437 ;
  assign n55439 = ~\pi1152  & ~n12257 ;
  assign n55440 = n50677 & n55439 ;
  assign n55441 = ~n53117 & ~n55440 ;
  assign n55442 = ~\pi0211  & n55354 ;
  assign n55443 = ~n50570 & ~n51118 ;
  assign n55444 = ~n55442 & n55443 ;
  assign n55445 = \pi0219  & n51125 ;
  assign n55446 = ~n55444 & n55445 ;
  assign n55447 = n9948 & ~n55446 ;
  assign n55448 = n50430 & ~n55354 ;
  assign n55449 = ~n55373 & ~n55375 ;
  assign n55450 = ~\pi0212  & n50877 ;
  assign n55451 = n51112 & n55450 ;
  assign n55452 = ~\pi0212  & n51115 ;
  assign n55453 = n51114 & n55452 ;
  assign n55454 = ~\pi0219  & ~n55453 ;
  assign n55455 = ~n55451 & n55454 ;
  assign n55456 = n55449 & n55455 ;
  assign n55457 = ~n55448 & n55456 ;
  assign n55458 = ~\pi0212  & n55454 ;
  assign n55459 = ~n55451 & n55458 ;
  assign n55460 = ~\pi1152  & ~n55459 ;
  assign n55461 = ~n55457 & n55460 ;
  assign n55462 = n55447 & n55461 ;
  assign n55463 = n55441 & ~n55462 ;
  assign n55464 = \pi0214  & n55354 ;
  assign n55465 = ~n55366 & ~n55464 ;
  assign n55466 = n55381 & ~n55465 ;
  assign n55467 = n55447 & ~n55466 ;
  assign n55468 = n55018 & ~n55467 ;
  assign n55469 = \pi1150  & ~n55468 ;
  assign n55470 = ~n55463 & n55469 ;
  assign n55471 = ~n55438 & ~n55470 ;
  assign n55472 = ~n55420 & n55471 ;
  assign n55473 = ~n55385 & n55472 ;
  assign n55474 = ~\pi0213  & ~n55473 ;
  assign n55475 = \pi0213  & n51197 ;
  assign n55476 = n51252 & n55475 ;
  assign n55477 = \pi0209  & ~n55476 ;
  assign n55478 = \pi0230  & n55477 ;
  assign n55479 = ~n55474 & n55478 ;
  assign n55480 = \pi0214  & n53096 ;
  assign n55481 = \pi0299  & ~n50946 ;
  assign n55482 = n52773 & ~n55481 ;
  assign n55483 = \pi0212  & ~n55482 ;
  assign n55484 = ~n55480 & n55483 ;
  assign n55485 = \pi0299  & n50946 ;
  assign n55486 = n53053 & ~n55485 ;
  assign n55487 = ~\pi0219  & ~n52995 ;
  assign n55488 = \pi1151  & n55487 ;
  assign n55489 = ~n55486 & n55488 ;
  assign n55490 = ~n55484 & n55489 ;
  assign n55491 = ~\pi1151  & ~n54778 ;
  assign n55492 = \pi1151  & ~n53090 ;
  assign n55493 = ~n55491 & ~n55492 ;
  assign n55494 = ~n55490 & n55493 ;
  assign n55495 = \pi0299  & ~n12255 ;
  assign n55496 = ~n50946 & n55495 ;
  assign n55497 = ~n51913 & ~n55496 ;
  assign n55498 = ~n50947 & n50948 ;
  assign n55499 = ~n55497 & n55498 ;
  assign n55500 = n51966 & n55499 ;
  assign n55501 = ~\pi1150  & ~n55500 ;
  assign n55502 = n50975 & n55501 ;
  assign n55503 = ~n55494 & n55502 ;
  assign n55504 = ~n51169 & ~n52741 ;
  assign n55505 = n51997 & ~n55504 ;
  assign n55506 = n50952 & ~n55505 ;
  assign n55507 = n55501 & n55506 ;
  assign n55508 = n52750 & ~n55485 ;
  assign n55509 = n50679 & ~n55508 ;
  assign n55510 = ~n50586 & n52750 ;
  assign n55511 = n50772 & ~n55510 ;
  assign n55512 = ~n55509 & ~n55511 ;
  assign n55513 = n51175 & n55501 ;
  assign n55514 = ~n55512 & n55513 ;
  assign n55515 = ~n55507 & ~n55514 ;
  assign n55516 = \pi0213  & n55515 ;
  assign n55517 = ~n55503 & n55516 ;
  assign n55518 = ~\pi0209  & ~n55517 ;
  assign n55519 = n6848 & ~n54859 ;
  assign n55520 = ~n6848 & n50950 ;
  assign n55521 = n51965 & ~n55520 ;
  assign n55522 = ~n55519 & n55521 ;
  assign n55523 = ~n52329 & ~n55485 ;
  assign n55524 = ~n52708 & n55523 ;
  assign n55525 = ~\pi0212  & ~n55524 ;
  assign n55526 = ~\pi0214  & ~n55485 ;
  assign n55527 = ~n52708 & n55526 ;
  assign n55528 = ~\pi0211  & \pi0212  ;
  assign n55529 = n50586 & n55528 ;
  assign n55530 = ~n50600 & ~n55529 ;
  assign n55531 = \pi0212  & ~n52000 ;
  assign n55532 = ~n52707 & n55531 ;
  assign n55533 = n55530 & ~n55532 ;
  assign n55534 = ~n55527 & ~n55533 ;
  assign n55535 = ~n55525 & ~n55534 ;
  assign n55536 = ~\pi0219  & n55521 ;
  assign n55537 = ~n55535 & n55536 ;
  assign n55538 = ~n55522 & ~n55537 ;
  assign n55539 = ~\pi1152  & ~n55538 ;
  assign n55540 = n51975 & n52274 ;
  assign n55541 = n50946 & n54305 ;
  assign n55542 = ~n55540 & ~n55541 ;
  assign n55543 = \pi0214  & ~n51913 ;
  assign n55544 = n51975 & n55543 ;
  assign n55545 = \pi0212  & ~n55544 ;
  assign n55546 = n55542 & n55545 ;
  assign n55547 = ~\pi0219  & ~n55546 ;
  assign n55548 = n50693 & n50946 ;
  assign n55549 = n51975 & n52776 ;
  assign n55550 = ~n55548 & ~n55549 ;
  assign n55551 = ~\pi0212  & ~n52329 ;
  assign n55552 = n55550 & n55551 ;
  assign n55553 = \pi1151  & ~n55552 ;
  assign n55554 = n55547 & n55553 ;
  assign n55555 = \pi1151  & ~n6848 ;
  assign n55556 = \pi0219  & \pi1151  ;
  assign n55557 = n51975 & n55556 ;
  assign n55558 = ~n55555 & ~n55557 ;
  assign n55559 = ~\pi0057  & n55558 ;
  assign n55560 = ~n55554 & n55559 ;
  assign n55561 = n50952 & ~n55560 ;
  assign n55562 = n50586 & n50967 ;
  assign n55563 = ~n55541 & ~n55562 ;
  assign n55564 = \pi0212  & n55563 ;
  assign n55565 = ~n52654 & n55564 ;
  assign n55566 = ~n55486 & ~n55565 ;
  assign n55567 = n54484 & n55566 ;
  assign n55568 = ~\pi1151  & n9948 ;
  assign n55569 = ~n55567 & n55568 ;
  assign n55570 = ~n52675 & n55569 ;
  assign n55571 = ~\pi0219  & ~n52798 ;
  assign n55572 = n50970 & ~n55496 ;
  assign n55573 = n52616 & ~n55572 ;
  assign n55574 = n55571 & ~n55573 ;
  assign n55575 = ~n52712 & ~n53004 ;
  assign n55576 = \pi1151  & ~n55575 ;
  assign n55577 = ~n55574 & n55576 ;
  assign n55578 = n50975 & ~n55577 ;
  assign n55579 = ~n55570 & n55578 ;
  assign n55580 = ~n55561 & ~n55579 ;
  assign n55581 = ~n55539 & n55580 ;
  assign n55582 = ~\pi0209  & \pi1150  ;
  assign n55583 = ~n55581 & n55582 ;
  assign n55584 = ~n55518 & ~n55583 ;
  assign n55585 = ~\pi0213  & ~n55224 ;
  assign n55586 = ~n55214 & n55585 ;
  assign n55587 = \pi0230  & ~n55586 ;
  assign n55588 = ~n55584 & n55587 ;
  assign n55589 = ~\pi0230  & ~\pi0249  ;
  assign n55590 = ~n55588 & ~n55589 ;
  assign n55591 = ~n55479 & n55590 ;
  assign n55592 = ~\pi0087  & ~\pi0250  ;
  assign n55593 = n10017 & n55592 ;
  assign n55594 = ~\pi0038  & n10094 ;
  assign n55595 = n6784 & n55594 ;
  assign n55596 = n1266 & n55595 ;
  assign n55597 = n1354 & n55596 ;
  assign n55598 = n1358 & n55597 ;
  assign n55599 = n55593 & n55598 ;
  assign n55600 = n1578 & n2402 ;
  assign n55601 = n13771 & n55600 ;
  assign n55602 = n13788 & n55601 ;
  assign n55603 = ~n6789 & ~n55602 ;
  assign n55604 = ~\pi0075  & n55593 ;
  assign n55605 = ~n55603 & n55604 ;
  assign n55606 = ~n55599 & ~n55605 ;
  assign n55607 = ~\pi0476  & n13645 ;
  assign n55608 = ~\pi0199  & ~\pi0200  ;
  assign n55609 = \pi0897  & n55608 ;
  assign n55610 = ~n55607 & ~n55609 ;
  assign n55611 = \pi0200  & \pi1039  ;
  assign n55612 = ~\pi0200  & \pi1053  ;
  assign n55613 = ~\pi0199  & ~n55612 ;
  assign n55614 = ~n55611 & n55613 ;
  assign n55615 = ~n55610 & ~n55614 ;
  assign n55616 = \pi0251  & n55610 ;
  assign n55617 = ~n55615 & ~n55616 ;
  assign n55618 = \pi0057  & n13815 ;
  assign n55619 = n10003 & ~n55618 ;
  assign n55620 = ~\pi0057  & \pi1092  ;
  assign n55621 = n55619 & ~n55620 ;
  assign n55622 = ~\pi0979  & ~\pi0984  ;
  assign n55623 = \pi1001  & n55622 ;
  assign n55624 = n6720 & n9627 ;
  assign n55625 = n55623 & n55624 ;
  assign n55626 = n27402 & n55625 ;
  assign n55627 = n6705 & n55626 ;
  assign n55628 = ~n50322 & n55627 ;
  assign n55629 = n12966 & n55628 ;
  assign n55630 = ~\pi0252  & n55619 ;
  assign n55631 = ~n55629 & n55630 ;
  assign n55632 = ~n55621 & ~n55631 ;
  assign n55633 = ~n12971 & n13816 ;
  assign n55634 = ~n10003 & ~n55633 ;
  assign n55635 = n55632 & ~n55634 ;
  assign n55636 = ~n6709 & n13816 ;
  assign n55637 = n6735 & n55636 ;
  assign n55638 = ~n6732 & n55637 ;
  assign n55639 = n6720 & ~n6810 ;
  assign n55640 = ~\pi0287  & \pi1001  ;
  assign n55641 = n55622 & n55640 ;
  assign n55642 = n55639 & n55641 ;
  assign n55643 = n1259 & n55642 ;
  assign n55644 = n1281 & n55643 ;
  assign n55645 = n1249 & n55644 ;
  assign n55646 = ~\pi0252  & ~n55645 ;
  assign n55647 = \pi1091  & n10049 ;
  assign n55648 = ~n13630 & n55647 ;
  assign n55649 = n6921 & n55648 ;
  assign n55650 = ~n55646 & n55649 ;
  assign n55651 = ~n6736 & ~n55650 ;
  assign n55652 = \pi0252  & n10049 ;
  assign n55653 = n1249 & n10049 ;
  assign n55654 = n55644 & n55653 ;
  assign n55655 = ~n55652 & ~n55654 ;
  assign n55656 = ~n6954 & n55655 ;
  assign n55657 = ~n6732 & ~n55656 ;
  assign n55658 = n55651 & n55657 ;
  assign n55659 = ~n55638 & ~n55658 ;
  assign n55660 = \pi0299  & ~n6732 ;
  assign n55661 = \pi0299  & ~n13816 ;
  assign n55662 = \pi0299  & ~n6706 ;
  assign n55663 = ~n6713 & n55662 ;
  assign n55664 = ~n55661 & ~n55663 ;
  assign n55665 = ~n55660 & n55664 ;
  assign n55666 = n6714 & ~n55650 ;
  assign n55667 = ~n55656 & ~n55660 ;
  assign n55668 = n55666 & n55667 ;
  assign n55669 = ~n55665 & ~n55668 ;
  assign n55670 = n55659 & n55669 ;
  assign n55671 = n12971 & ~n55670 ;
  assign n55672 = ~n6761 & n55637 ;
  assign n55673 = ~n6761 & ~n55656 ;
  assign n55674 = n55651 & n55673 ;
  assign n55675 = ~n55672 & ~n55674 ;
  assign n55676 = ~\pi0299  & ~n6761 ;
  assign n55677 = ~\pi0299  & ~n13816 ;
  assign n55678 = ~\pi0299  & ~n6706 ;
  assign n55679 = ~n6713 & n55678 ;
  assign n55680 = ~n55677 & ~n55679 ;
  assign n55681 = ~n55676 & n55680 ;
  assign n55682 = ~n55656 & ~n55676 ;
  assign n55683 = n55666 & n55682 ;
  assign n55684 = ~n55681 & ~n55683 ;
  assign n55685 = n55675 & n55684 ;
  assign n55686 = n55632 & ~n55685 ;
  assign n55687 = n55671 & n55686 ;
  assign n55688 = ~n55635 & ~n55687 ;
  assign n55689 = ~n50701 & ~n52001 ;
  assign n55690 = ~n50384 & n55689 ;
  assign n55691 = n9948 & n55690 ;
  assign n55692 = ~n9948 & n50689 ;
  assign n55693 = ~n55691 & ~n55692 ;
  assign n55694 = ~\pi1151  & \pi1153  ;
  assign n55695 = ~n55693 & n55694 ;
  assign n55696 = ~n44035 & ~n50462 ;
  assign n55697 = n12577 & ~n55696 ;
  assign n55698 = \pi0211  & ~n50364 ;
  assign n55699 = ~n55697 & ~n55698 ;
  assign n55700 = ~n44035 & ~n50502 ;
  assign n55701 = n50689 & ~n55700 ;
  assign n55702 = n51997 & ~n55701 ;
  assign n55703 = n55699 & n55702 ;
  assign n55704 = ~n55695 & ~n55703 ;
  assign n55705 = ~\pi1152  & ~n55704 ;
  assign n55706 = \pi1153  & n50689 ;
  assign n55707 = ~n50432 & n55706 ;
  assign n55708 = ~\pi1151  & ~n13648 ;
  assign n55709 = ~n50373 & n55708 ;
  assign n55710 = ~n55707 & n55709 ;
  assign n55711 = ~n44032 & ~n52000 ;
  assign n55712 = \pi1153  & ~n55711 ;
  assign n55713 = ~n13550 & ~n50701 ;
  assign n55714 = \pi1151  & n55713 ;
  assign n55715 = ~n55712 & n55714 ;
  assign n55716 = n50998 & ~n55715 ;
  assign n55717 = ~n55710 & n55716 ;
  assign n55718 = \pi0219  & ~\pi1153  ;
  assign n55719 = ~n50713 & ~n55718 ;
  assign n55720 = \pi1151  & ~n13647 ;
  assign n55721 = \pi1152  & ~n12577 ;
  assign n55722 = ~n55720 & ~n55721 ;
  assign n55723 = n55719 & ~n55722 ;
  assign n55724 = ~n9948 & n55723 ;
  assign n55725 = \pi0230  & ~n55724 ;
  assign n55726 = ~n55717 & n55725 ;
  assign n55727 = ~n55705 & n55726 ;
  assign n55728 = ~\pi0230  & ~\pi1152  ;
  assign n55729 = \pi1091  & n55698 ;
  assign n55730 = \pi1091  & n12577 ;
  assign n55731 = ~n55696 & n55730 ;
  assign n55732 = ~n55729 & ~n55731 ;
  assign n55733 = \pi1153  & ~n53866 ;
  assign n55734 = n51100 & n55608 ;
  assign n55735 = ~\pi1091  & ~\pi1153  ;
  assign n55736 = n50689 & ~n55735 ;
  assign n55737 = ~n55734 & n55736 ;
  assign n55738 = ~n55733 & n55737 ;
  assign n55739 = n55732 & ~n55738 ;
  assign n55740 = ~\pi0057  & n6848 ;
  assign n55741 = \pi1091  & ~\pi1153  ;
  assign n55742 = \pi0219  & n55741 ;
  assign n55743 = ~\pi0253  & ~\pi1091  ;
  assign n55744 = \pi0211  & \pi1091  ;
  assign n55745 = ~n55743 & ~n55744 ;
  assign n55746 = ~n55742 & n55745 ;
  assign n55747 = ~n55740 & n55746 ;
  assign n55748 = \pi0253  & \pi1151  ;
  assign n55749 = ~n55747 & n55748 ;
  assign n55750 = ~n55739 & n55749 ;
  assign n55751 = ~\pi0253  & ~\pi0299  ;
  assign n55752 = ~n12691 & n55751 ;
  assign n55753 = ~\pi0253  & \pi0299  ;
  assign n55754 = ~n12577 & n55753 ;
  assign n55755 = ~n55752 & ~n55754 ;
  assign n55756 = ~n55712 & ~n55755 ;
  assign n55757 = ~\pi0057  & ~n55743 ;
  assign n55758 = n6848 & n55757 ;
  assign n55759 = ~n55756 & n55758 ;
  assign n55760 = \pi1151  & ~n55747 ;
  assign n55761 = ~n55759 & n55760 ;
  assign n55762 = \pi0219  & \pi1091  ;
  assign n55763 = ~n50625 & n55762 ;
  assign n55764 = \pi0219  & ~n55743 ;
  assign n55765 = ~n55763 & n55764 ;
  assign n55766 = ~n9948 & n55765 ;
  assign n55767 = \pi1091  & \pi1153  ;
  assign n55768 = ~\pi0057  & n55767 ;
  assign n55769 = n6848 & n55768 ;
  assign n55770 = n55690 & n55769 ;
  assign n55771 = \pi0253  & ~\pi1091  ;
  assign n55772 = ~\pi1151  & ~n55771 ;
  assign n55773 = ~n55770 & n55772 ;
  assign n55774 = ~n55766 & n55773 ;
  assign n55775 = ~n55761 & ~n55774 ;
  assign n55776 = ~n55750 & n55775 ;
  assign n55777 = n55728 & ~n55776 ;
  assign n55778 = ~n50432 & n55767 ;
  assign n55779 = n51001 & n53866 ;
  assign n55780 = n50689 & ~n55779 ;
  assign n55781 = ~n55778 & n55780 ;
  assign n55782 = ~n50363 & n53829 ;
  assign n55783 = n50371 & n55782 ;
  assign n55784 = \pi0211  & ~n53896 ;
  assign n55785 = ~n55783 & n55784 ;
  assign n55786 = ~\pi0253  & ~n55785 ;
  assign n55787 = ~n55781 & n55786 ;
  assign n55788 = n13645 & n51100 ;
  assign n55789 = ~n55735 & ~n55788 ;
  assign n55790 = n50689 & n53829 ;
  assign n55791 = ~n50371 & n55790 ;
  assign n55792 = ~n52096 & ~n55791 ;
  assign n55793 = n55789 & ~n55792 ;
  assign n55794 = n13647 & n53829 ;
  assign n55795 = ~n50373 & n55794 ;
  assign n55796 = \pi0253  & ~n55795 ;
  assign n55797 = ~n55793 & n55796 ;
  assign n55798 = ~n55787 & ~n55797 ;
  assign n55799 = ~n13647 & ~n50689 ;
  assign n55800 = ~n55771 & n55799 ;
  assign n55801 = ~n55783 & n55800 ;
  assign n55802 = n51966 & ~n53905 ;
  assign n55803 = ~n55801 & n55802 ;
  assign n55804 = ~n55798 & n55803 ;
  assign n55805 = ~n55743 & ~n55763 ;
  assign n55806 = ~n9948 & n55805 ;
  assign n55807 = \pi1091  & ~\pi1151  ;
  assign n55808 = n12577 & n55807 ;
  assign n55809 = n55806 & ~n55808 ;
  assign n55810 = ~n53905 & n55809 ;
  assign n55811 = \pi1152  & n55741 ;
  assign n55812 = \pi1152  & ~n55771 ;
  assign n55813 = n55711 & n55812 ;
  assign n55814 = ~n55811 & ~n55813 ;
  assign n55815 = n55713 & ~n55814 ;
  assign n55816 = n51996 & ~n55743 ;
  assign n55817 = n6848 & n55816 ;
  assign n55818 = \pi1152  & ~n55817 ;
  assign n55819 = ~n53905 & ~n55818 ;
  assign n55820 = ~n55815 & n55819 ;
  assign n55821 = ~n55810 & ~n55820 ;
  assign n55822 = ~\pi0230  & n55821 ;
  assign n55823 = ~n55804 & n55822 ;
  assign n55824 = ~n55777 & ~n55823 ;
  assign n55825 = ~n55727 & n55824 ;
  assign n55826 = \pi1153  & ~n53664 ;
  assign n55827 = ~n53803 & n55826 ;
  assign n55828 = \pi0219  & \pi1153  ;
  assign n55829 = \pi0219  & n53597 ;
  assign n55830 = ~n55828 & ~n55829 ;
  assign n55831 = n53586 & ~n55828 ;
  assign n55832 = ~n53585 & n55831 ;
  assign n55833 = ~n55830 & ~n55832 ;
  assign n55834 = ~n55827 & n55833 ;
  assign n55835 = ~n53575 & n53750 ;
  assign n55836 = \pi0211  & n53561 ;
  assign n55837 = ~n53559 & n55836 ;
  assign n55838 = n53568 & ~n55837 ;
  assign n55839 = ~n53587 & ~n55838 ;
  assign n55840 = n55833 & n55839 ;
  assign n55841 = n55835 & n55840 ;
  assign n55842 = ~n55834 & ~n55841 ;
  assign n55843 = \pi0253  & ~n55842 ;
  assign n55844 = ~\pi0219  & ~n53556 ;
  assign n55845 = ~n55838 & n55844 ;
  assign n55846 = ~n53587 & n55845 ;
  assign n55847 = \pi1153  & n53569 ;
  assign n55848 = n51033 & ~n53585 ;
  assign n55849 = ~n55847 & ~n55848 ;
  assign n55850 = \pi0253  & n55849 ;
  assign n55851 = n55846 & n55850 ;
  assign n55852 = n55740 & ~n55851 ;
  assign n55853 = ~n55843 & n55852 ;
  assign n55854 = \pi0253  & ~n53590 ;
  assign n55855 = \pi0219  & n55854 ;
  assign n55856 = ~\pi1091  & n55854 ;
  assign n55857 = n53555 & n55856 ;
  assign n55858 = ~n55855 & ~n55857 ;
  assign n55859 = ~\pi0211  & n53561 ;
  assign n55860 = ~n53559 & n55859 ;
  assign n55861 = \pi0211  & \pi0273  ;
  assign n55862 = n53934 & n55861 ;
  assign n55863 = \pi0219  & ~n55862 ;
  assign n55864 = ~n55860 & n55863 ;
  assign n55865 = \pi0219  & ~\pi0253  ;
  assign n55866 = ~\pi0253  & n53542 ;
  assign n55867 = n53540 & n55866 ;
  assign n55868 = ~n55865 & ~n55867 ;
  assign n55869 = ~n55864 & ~n55868 ;
  assign n55870 = n55858 & ~n55869 ;
  assign n55871 = ~n9948 & ~n55763 ;
  assign n55872 = ~n55870 & n55871 ;
  assign n55873 = ~\pi0219  & n53542 ;
  assign n55874 = n53540 & n55873 ;
  assign n55875 = ~n53711 & ~n55874 ;
  assign n55876 = ~n53556 & ~n55875 ;
  assign n55877 = ~\pi0219  & n53561 ;
  assign n55878 = ~n9948 & n55877 ;
  assign n55879 = ~n53559 & n55878 ;
  assign n55880 = ~n55876 & n55879 ;
  assign n55881 = ~n55872 & ~n55880 ;
  assign n55882 = \pi1151  & n55881 ;
  assign n55883 = ~n55853 & n55882 ;
  assign n55884 = ~\pi0211  & ~n53564 ;
  assign n55885 = ~\pi0211  & n53538 ;
  assign n55886 = ~n53553 & n55885 ;
  assign n55887 = ~n55884 & ~n55886 ;
  assign n55888 = ~n53776 & ~n55887 ;
  assign n55889 = n53565 & n53677 ;
  assign n55890 = ~n53591 & ~n55889 ;
  assign n55891 = ~n55888 & ~n55890 ;
  assign n55892 = ~\pi1153  & ~n53770 ;
  assign n55893 = \pi0219  & ~n55892 ;
  assign n55894 = ~n55891 & n55893 ;
  assign n55895 = \pi1153  & ~n53569 ;
  assign n55896 = ~n53566 & n55895 ;
  assign n55897 = ~\pi1153  & ~n53569 ;
  assign n55898 = ~n53677 & n55897 ;
  assign n55899 = ~\pi0219  & ~n55898 ;
  assign n55900 = ~n55896 & n55899 ;
  assign n55901 = ~n53616 & ~n55888 ;
  assign n55902 = n55844 & ~n55901 ;
  assign n55903 = ~n55900 & n55902 ;
  assign n55904 = ~n55894 & ~n55903 ;
  assign n55905 = ~n53702 & ~n55904 ;
  assign n55906 = ~\pi0253  & \pi1151  ;
  assign n55907 = ~n55880 & n55906 ;
  assign n55908 = ~n55872 & n55907 ;
  assign n55909 = ~n55905 & n55908 ;
  assign n55910 = ~n55883 & ~n55909 ;
  assign n55911 = ~n53554 & n53586 ;
  assign n55912 = \pi0219  & ~n55911 ;
  assign n55913 = ~n55892 & n55912 ;
  assign n55914 = ~n55891 & n55913 ;
  assign n55915 = ~n52725 & ~n55874 ;
  assign n55916 = ~n53586 & ~n55915 ;
  assign n55917 = n53538 & ~n55915 ;
  assign n55918 = ~n53553 & n55917 ;
  assign n55919 = ~n55916 & ~n55918 ;
  assign n55920 = ~\pi1153  & ~n53577 ;
  assign n55921 = ~n53645 & n55920 ;
  assign n55922 = ~n53702 & ~n55921 ;
  assign n55923 = ~n55919 & n55922 ;
  assign n55924 = ~\pi0253  & ~n55923 ;
  assign n55925 = ~n55914 & n55924 ;
  assign n55926 = n55835 & n55839 ;
  assign n55927 = ~\pi1153  & ~n53591 ;
  assign n55928 = ~n53677 & n55927 ;
  assign n55929 = ~n55741 & ~n55928 ;
  assign n55930 = ~\pi0219  & ~n53569 ;
  assign n55931 = n53591 & ~n55930 ;
  assign n55932 = ~n53611 & ~n55931 ;
  assign n55933 = n55929 & ~n55932 ;
  assign n55934 = ~n55926 & n55933 ;
  assign n55935 = \pi0253  & ~n55934 ;
  assign n55936 = ~n55925 & ~n55935 ;
  assign n55937 = n9948 & n55936 ;
  assign n55938 = ~\pi1151  & ~n55872 ;
  assign n55939 = ~n55937 & n55938 ;
  assign n55940 = n55910 & ~n55939 ;
  assign n55941 = ~\pi1152  & ~n55940 ;
  assign n55942 = \pi1151  & ~n55880 ;
  assign n55943 = ~n55872 & n55942 ;
  assign n55944 = ~n53554 & n55831 ;
  assign n55945 = ~n55830 & ~n55944 ;
  assign n55946 = ~\pi1153  & n55945 ;
  assign n55947 = n55839 & n55945 ;
  assign n55948 = n55835 & n55947 ;
  assign n55949 = ~n55946 & ~n55948 ;
  assign n55950 = ~n53575 & ~n53581 ;
  assign n55951 = \pi1153  & ~n55950 ;
  assign n55952 = ~\pi0219  & \pi1153  ;
  assign n55953 = n55919 & ~n55952 ;
  assign n55954 = ~n55951 & ~n55953 ;
  assign n55955 = \pi0253  & ~n55954 ;
  assign n55956 = n55949 & n55955 ;
  assign n55957 = \pi0219  & n55892 ;
  assign n55958 = \pi0219  & ~n55888 ;
  assign n55959 = ~n55890 & n55958 ;
  assign n55960 = ~n55957 & ~n55959 ;
  assign n55961 = ~\pi0253  & ~n55900 ;
  assign n55962 = n55960 & n55961 ;
  assign n55963 = ~n55956 & ~n55962 ;
  assign n55964 = n9948 & ~n55963 ;
  assign n55965 = n55943 & ~n55964 ;
  assign n55966 = ~n53569 & ~n53611 ;
  assign n55967 = ~\pi1153  & ~n55966 ;
  assign n55968 = ~n53566 & n55839 ;
  assign n55969 = ~n55967 & n55968 ;
  assign n55970 = ~\pi0219  & ~n55969 ;
  assign n55971 = n55960 & ~n55970 ;
  assign n55972 = \pi0219  & n53586 ;
  assign n55973 = ~n53585 & n55972 ;
  assign n55974 = ~\pi0057  & ~\pi0253  ;
  assign n55975 = n6848 & n55974 ;
  assign n55976 = ~n55973 & n55975 ;
  assign n55977 = n55971 & n55976 ;
  assign n55978 = \pi1153  & ~n53814 ;
  assign n55979 = ~n55926 & n55978 ;
  assign n55980 = ~n53575 & n55829 ;
  assign n55981 = ~n55979 & n55980 ;
  assign n55982 = ~n53612 & ~n55967 ;
  assign n55983 = n55902 & ~n55982 ;
  assign n55984 = ~\pi0057  & \pi0253  ;
  assign n55985 = n6848 & n55984 ;
  assign n55986 = ~n55983 & n55985 ;
  assign n55987 = ~n55981 & n55986 ;
  assign n55988 = ~n55977 & ~n55987 ;
  assign n55989 = ~\pi1151  & n55988 ;
  assign n55990 = ~n55965 & ~n55989 ;
  assign n55991 = ~\pi0219  & ~n53543 ;
  assign n55992 = ~n55860 & n55991 ;
  assign n55993 = n55844 & ~n55992 ;
  assign n55994 = n52628 & n53567 ;
  assign n55995 = ~n55993 & n55994 ;
  assign n55996 = ~n55872 & ~n55995 ;
  assign n55997 = \pi1152  & n55996 ;
  assign n55998 = ~n55990 & n55997 ;
  assign n55999 = ~n55941 & ~n55998 ;
  assign n56000 = n53905 & ~n55727 ;
  assign n56001 = n55999 & n56000 ;
  assign n56002 = ~n55825 & ~n56001 ;
  assign n56003 = ~n53618 & ~n53645 ;
  assign n56004 = ~\pi1154  & ~n56003 ;
  assign n56005 = ~\pi1153  & ~n55838 ;
  assign n56006 = ~n53587 & n56005 ;
  assign n56007 = ~n53566 & n56006 ;
  assign n56008 = ~\pi1154  & n55966 ;
  assign n56009 = n56007 & n56008 ;
  assign n56010 = ~n56004 & ~n56009 ;
  assign n56011 = \pi1154  & ~n53578 ;
  assign n56012 = ~n53553 & n56011 ;
  assign n56013 = ~n50416 & ~n56012 ;
  assign n56014 = n55839 & ~n56013 ;
  assign n56015 = ~n55951 & n56014 ;
  assign n56016 = ~\pi0219  & \pi0254  ;
  assign n56017 = ~n56015 & n56016 ;
  assign n56018 = n56010 & n56017 ;
  assign n56019 = ~n53578 & n53597 ;
  assign n56020 = ~n53553 & n56019 ;
  assign n56021 = ~n53775 & ~n56020 ;
  assign n56022 = \pi1154  & ~n56021 ;
  assign n56023 = ~n53566 & n56022 ;
  assign n56024 = ~n53678 & ~n56023 ;
  assign n56025 = n52001 & ~n53543 ;
  assign n56026 = ~n53564 & ~n56025 ;
  assign n56027 = n53538 & ~n56025 ;
  assign n56028 = ~n53553 & n56027 ;
  assign n56029 = ~n56026 & ~n56028 ;
  assign n56030 = ~\pi1153  & n56029 ;
  assign n56031 = ~\pi0254  & ~n56030 ;
  assign n56032 = ~\pi0219  & n56031 ;
  assign n56033 = ~n56024 & n56032 ;
  assign n56034 = \pi0253  & ~n56033 ;
  assign n56035 = ~n56018 & n56034 ;
  assign n56036 = \pi1153  & n43637 ;
  assign n56037 = ~n44032 & n50609 ;
  assign n56038 = ~n56036 & n56037 ;
  assign n56039 = ~\pi1154  & ~n51110 ;
  assign n56040 = ~n51038 & ~n56039 ;
  assign n56041 = ~n56038 & n56040 ;
  assign n56042 = ~\pi0211  & \pi1091  ;
  assign n56043 = \pi1154  & n56042 ;
  assign n56044 = ~n55762 & ~n56043 ;
  assign n56045 = ~n56041 & ~n56044 ;
  assign n56046 = \pi1154  & ~n44032 ;
  assign n56047 = n55744 & n56046 ;
  assign n56048 = ~\pi0219  & ~n51940 ;
  assign n56049 = n56047 & n56048 ;
  assign n56050 = ~n55734 & ~n55735 ;
  assign n56051 = ~\pi1153  & ~\pi1154  ;
  assign n56052 = \pi0199  & ~\pi1154  ;
  assign n56053 = n53829 & n56052 ;
  assign n56054 = ~n56051 & ~n56053 ;
  assign n56055 = n56050 & ~n56054 ;
  assign n56056 = ~\pi0219  & ~n52230 ;
  assign n56057 = ~n12691 & n52725 ;
  assign n56058 = ~n56056 & ~n56057 ;
  assign n56059 = n56055 & ~n56058 ;
  assign n56060 = ~n56049 & ~n56059 ;
  assign n56061 = ~n56045 & n56060 ;
  assign n56062 = ~\pi0253  & \pi0254  ;
  assign n56063 = ~n56061 & n56062 ;
  assign n56064 = ~\pi0254  & ~\pi1091  ;
  assign n56065 = ~\pi0253  & n56064 ;
  assign n56066 = ~\pi0200  & \pi1154  ;
  assign n56067 = ~\pi0219  & ~n56066 ;
  assign n56068 = n13558 & n56067 ;
  assign n56069 = ~\pi0219  & ~n52000 ;
  assign n56070 = n51176 & n56069 ;
  assign n56071 = ~n56068 & ~n56070 ;
  assign n56072 = \pi1154  & ~n55711 ;
  assign n56073 = \pi0219  & ~n51110 ;
  assign n56074 = ~n56072 & n56073 ;
  assign n56075 = n56071 & ~n56074 ;
  assign n56076 = ~\pi0253  & ~\pi0254  ;
  assign n56077 = ~n56075 & n56076 ;
  assign n56078 = ~n56065 & ~n56077 ;
  assign n56079 = n9948 & n56078 ;
  assign n56080 = ~n56063 & n56079 ;
  assign n56081 = ~n56035 & n56080 ;
  assign n56082 = n53804 & ~n55926 ;
  assign n56083 = \pi1154  & n55839 ;
  assign n56084 = n55835 & n56083 ;
  assign n56085 = ~n50510 & ~n56084 ;
  assign n56086 = ~n56082 & ~n56085 ;
  assign n56087 = \pi1153  & n53776 ;
  assign n56088 = ~\pi1154  & n53597 ;
  assign n56089 = ~n50460 & ~n56088 ;
  assign n56090 = ~n50460 & n53586 ;
  assign n56091 = ~n53585 & n56090 ;
  assign n56092 = ~n56089 & ~n56091 ;
  assign n56093 = ~n56087 & n56092 ;
  assign n56094 = \pi0254  & ~n56093 ;
  assign n56095 = ~n56086 & n56094 ;
  assign n56096 = ~\pi0299  & ~n53585 ;
  assign n56097 = ~\pi1153  & ~n53664 ;
  assign n56098 = ~n53662 & n56097 ;
  assign n56099 = ~n56096 & ~n56098 ;
  assign n56100 = n53770 & n56099 ;
  assign n56101 = n53554 & ~n53591 ;
  assign n56102 = n53610 & n53743 ;
  assign n56103 = ~n56101 & ~n56102 ;
  assign n56104 = ~\pi1154  & n56103 ;
  assign n56105 = ~n56100 & n56104 ;
  assign n56106 = ~\pi1153  & n53776 ;
  assign n56107 = ~n53566 & ~n56021 ;
  assign n56108 = ~n56106 & n56107 ;
  assign n56109 = n50627 & ~n53563 ;
  assign n56110 = ~n56108 & n56109 ;
  assign n56111 = \pi1153  & ~n53591 ;
  assign n56112 = ~n53566 & n56111 ;
  assign n56113 = n50609 & n53744 ;
  assign n56114 = ~n56112 & n56113 ;
  assign n56115 = ~\pi0254  & ~n56114 ;
  assign n56116 = ~n56110 & n56115 ;
  assign n56117 = ~n56105 & n56116 ;
  assign n56118 = ~n56095 & ~n56117 ;
  assign n56119 = \pi0219  & n56080 ;
  assign n56120 = ~n56118 & n56119 ;
  assign n56121 = ~n56081 & ~n56120 ;
  assign n56122 = ~\pi0254  & ~n56075 ;
  assign n56123 = n9948 & ~n56064 ;
  assign n56124 = ~n56122 & n56123 ;
  assign n56125 = ~n50627 & n55762 ;
  assign n56126 = ~n50945 & n53909 ;
  assign n56127 = ~n56064 & ~n56126 ;
  assign n56128 = ~n56125 & n56127 ;
  assign n56129 = ~n9948 & n56128 ;
  assign n56130 = ~\pi0211  & n53909 ;
  assign n56131 = ~n9948 & n56130 ;
  assign n56132 = \pi1152  & ~n56131 ;
  assign n56133 = ~n56129 & n56132 ;
  assign n56134 = ~n56124 & n56133 ;
  assign n56135 = \pi0254  & n56133 ;
  assign n56136 = ~n56061 & n56135 ;
  assign n56137 = ~n56134 & ~n56136 ;
  assign n56138 = ~n53905 & n56137 ;
  assign n56139 = ~\pi0230  & ~n56138 ;
  assign n56140 = ~\pi0211  & n51036 ;
  assign n56141 = n53866 & n56140 ;
  assign n56142 = ~n50627 & ~n56141 ;
  assign n56143 = ~n51001 & n53829 ;
  assign n56144 = n50371 & n56143 ;
  assign n56145 = \pi1154  & ~n56144 ;
  assign n56146 = ~\pi0219  & ~n56145 ;
  assign n56147 = ~n56142 & n56146 ;
  assign n56148 = \pi0199  & n55741 ;
  assign n56149 = n44032 & n56148 ;
  assign n56150 = ~n55778 & ~n56149 ;
  assign n56151 = \pi0211  & ~n56051 ;
  assign n56152 = ~n56053 & n56151 ;
  assign n56153 = ~\pi0219  & n56152 ;
  assign n56154 = ~n56150 & n56153 ;
  assign n56155 = ~n50384 & n55741 ;
  assign n56156 = n50627 & ~n56155 ;
  assign n56157 = ~n55778 & n56156 ;
  assign n56158 = \pi0219  & \pi1154  ;
  assign n56159 = \pi0219  & n51036 ;
  assign n56160 = n53866 & n56159 ;
  assign n56161 = ~n56158 & ~n56160 ;
  assign n56162 = n50609 & ~n56144 ;
  assign n56163 = ~n56161 & ~n56162 ;
  assign n56164 = ~n56157 & n56163 ;
  assign n56165 = ~n56154 & ~n56164 ;
  assign n56166 = ~n56147 & n56165 ;
  assign n56167 = ~\pi0254  & ~n56166 ;
  assign n56168 = \pi1091  & ~n13647 ;
  assign n56169 = ~n51034 & n56168 ;
  assign n56170 = ~\pi1154  & ~n56169 ;
  assign n56171 = \pi1091  & n55799 ;
  assign n56172 = ~n51585 & n56171 ;
  assign n56173 = ~n50371 & n53829 ;
  assign n56174 = \pi1153  & ~n56173 ;
  assign n56175 = n50383 & n51100 ;
  assign n56176 = ~n55735 & ~n56175 ;
  assign n56177 = n55799 & n56176 ;
  assign n56178 = ~n56174 & n56177 ;
  assign n56179 = ~n56172 & ~n56178 ;
  assign n56180 = n53884 & ~n55792 ;
  assign n56181 = \pi1154  & ~n56180 ;
  assign n56182 = n56179 & n56181 ;
  assign n56183 = ~n56170 & ~n56182 ;
  assign n56184 = n13647 & n56176 ;
  assign n56185 = ~n56174 & n56184 ;
  assign n56186 = \pi1091  & ~\pi1154  ;
  assign n56187 = n13647 & n56186 ;
  assign n56188 = n51178 & n56187 ;
  assign n56189 = \pi0254  & ~n56188 ;
  assign n56190 = ~n56185 & n56189 ;
  assign n56191 = ~n56183 & n56190 ;
  assign n56192 = ~n56167 & ~n56191 ;
  assign n56193 = n9948 & ~n56192 ;
  assign n56194 = ~\pi1152  & ~n56129 ;
  assign n56195 = ~\pi0230  & n56194 ;
  assign n56196 = ~n56193 & n56195 ;
  assign n56197 = ~n56139 & ~n56196 ;
  assign n56198 = ~\pi0253  & ~n56128 ;
  assign n56199 = ~n9948 & ~n56198 ;
  assign n56200 = ~n56131 & ~n56199 ;
  assign n56201 = ~\pi0219  & ~n55767 ;
  assign n56202 = ~n53543 & n56201 ;
  assign n56203 = ~n55860 & n56202 ;
  assign n56204 = ~\pi0254  & ~n56125 ;
  assign n56205 = ~n55864 & n56204 ;
  assign n56206 = ~n56203 & n56205 ;
  assign n56207 = n13647 & n55741 ;
  assign n56208 = \pi0254  & ~n56207 ;
  assign n56209 = ~n56125 & n56208 ;
  assign n56210 = ~n55874 & n56209 ;
  assign n56211 = \pi0253  & ~n56210 ;
  assign n56212 = \pi0219  & n53561 ;
  assign n56213 = ~n53559 & n56212 ;
  assign n56214 = ~\pi0211  & ~n53937 ;
  assign n56215 = \pi0253  & ~n56214 ;
  assign n56216 = n56213 & n56215 ;
  assign n56217 = ~n56211 & ~n56216 ;
  assign n56218 = ~n56206 & ~n56217 ;
  assign n56219 = ~n56200 & ~n56218 ;
  assign n56220 = \pi1152  & ~n56219 ;
  assign n56221 = ~n56197 & n56220 ;
  assign n56222 = n56121 & n56221 ;
  assign n56223 = n13647 & ~n50945 ;
  assign n56224 = ~n51164 & ~n56223 ;
  assign n56225 = ~n55740 & n56224 ;
  assign n56226 = \pi1152  & ~n56225 ;
  assign n56227 = n9948 & n56071 ;
  assign n56228 = \pi0230  & ~n56227 ;
  assign n56229 = \pi0219  & \pi0230  ;
  assign n56230 = ~n56041 & n56229 ;
  assign n56231 = ~n56228 & ~n56230 ;
  assign n56232 = n56226 & ~n56231 ;
  assign n56233 = \pi1154  & ~n51215 ;
  assign n56234 = ~n50432 & n56233 ;
  assign n56235 = ~n51179 & ~n56234 ;
  assign n56236 = n13647 & ~n56235 ;
  assign n56237 = \pi0299  & n50689 ;
  assign n56238 = ~n13647 & n51003 ;
  assign n56239 = ~n56237 & ~n56238 ;
  assign n56240 = ~n51035 & ~n56239 ;
  assign n56241 = ~n56236 & ~n56240 ;
  assign n56242 = n9948 & ~n56241 ;
  assign n56243 = ~\pi0219  & ~n50945 ;
  assign n56244 = ~n51164 & ~n56243 ;
  assign n56245 = ~n9948 & n56244 ;
  assign n56246 = \pi0230  & ~\pi1152  ;
  assign n56247 = ~n56245 & n56246 ;
  assign n56248 = ~n56242 & n56247 ;
  assign n56249 = ~n56232 & ~n56248 ;
  assign n56250 = n53593 & ~n56106 ;
  assign n56251 = n50609 & ~n56250 ;
  assign n56252 = ~\pi1154  & ~n56100 ;
  assign n56253 = \pi0219  & ~n56106 ;
  assign n56254 = n56107 & n56253 ;
  assign n56255 = ~n51164 & ~n56254 ;
  assign n56256 = ~n56252 & ~n56255 ;
  assign n56257 = ~n56251 & n56256 ;
  assign n56258 = n50511 & ~n53573 ;
  assign n56259 = ~n55915 & ~n56258 ;
  assign n56260 = ~n53578 & ~n55915 ;
  assign n56261 = ~n53553 & n56260 ;
  assign n56262 = ~n56259 & ~n56261 ;
  assign n56263 = ~\pi0254  & ~n13647 ;
  assign n56264 = n56262 & n56263 ;
  assign n56265 = ~n55921 & ~n56096 ;
  assign n56266 = n53678 & n56265 ;
  assign n56267 = \pi1154  & ~n53564 ;
  assign n56268 = \pi1154  & n53538 ;
  assign n56269 = ~n53553 & n56268 ;
  assign n56270 = ~n56267 & ~n56269 ;
  assign n56271 = ~n56003 & ~n56270 ;
  assign n56272 = ~\pi0254  & ~n56271 ;
  assign n56273 = ~n56266 & n56272 ;
  assign n56274 = ~n56264 & ~n56273 ;
  assign n56275 = \pi0253  & ~n56274 ;
  assign n56276 = ~n56257 & n56275 ;
  assign n56277 = ~\pi1153  & n53597 ;
  assign n56278 = ~n53611 & n56277 ;
  assign n56279 = n55901 & ~n56278 ;
  assign n56280 = \pi0199  & n50511 ;
  assign n56281 = ~\pi1091  & n50511 ;
  assign n56282 = n53555 & n56281 ;
  assign n56283 = ~n56280 & ~n56282 ;
  assign n56284 = ~n53585 & ~n56283 ;
  assign n56285 = ~\pi0219  & ~n56284 ;
  assign n56286 = ~n56279 & n56285 ;
  assign n56287 = ~\pi1154  & ~n53586 ;
  assign n56288 = ~\pi1154  & n53538 ;
  assign n56289 = ~n53553 & n56288 ;
  assign n56290 = ~n56287 & ~n56289 ;
  assign n56291 = ~n53744 & ~n56290 ;
  assign n56292 = \pi1153  & ~n53573 ;
  assign n56293 = n53564 & n56292 ;
  assign n56294 = ~n53554 & n56293 ;
  assign n56295 = n53750 & ~n56294 ;
  assign n56296 = ~n56291 & ~n56295 ;
  assign n56297 = \pi0219  & ~n53591 ;
  assign n56298 = ~n53611 & n56297 ;
  assign n56299 = ~n51164 & ~n56298 ;
  assign n56300 = ~n56296 & ~n56299 ;
  assign n56301 = ~n56286 & ~n56300 ;
  assign n56302 = n53732 & ~n56301 ;
  assign n56303 = ~\pi0253  & n56192 ;
  assign n56304 = n9948 & n53905 ;
  assign n56305 = ~n56303 & n56304 ;
  assign n56306 = ~n56302 & n56305 ;
  assign n56307 = ~n56276 & n56306 ;
  assign n56308 = \pi1152  & n53905 ;
  assign n56309 = n56213 & ~n56214 ;
  assign n56310 = n56210 & ~n56309 ;
  assign n56311 = \pi0253  & ~n56310 ;
  assign n56312 = \pi0253  & ~n55992 ;
  assign n56313 = n55844 & n56312 ;
  assign n56314 = ~n56311 & ~n56313 ;
  assign n56315 = ~\pi0211  & ~n53543 ;
  assign n56316 = ~\pi0219  & n56315 ;
  assign n56317 = ~\pi0219  & ~\pi1091  ;
  assign n56318 = n53555 & n56317 ;
  assign n56319 = ~n56316 & ~n56318 ;
  assign n56320 = n56206 & n56319 ;
  assign n56321 = ~n56314 & ~n56320 ;
  assign n56322 = n53905 & n56199 ;
  assign n56323 = ~n56321 & n56322 ;
  assign n56324 = ~n56308 & ~n56323 ;
  assign n56325 = ~n56197 & n56324 ;
  assign n56326 = ~n56307 & n56325 ;
  assign n56327 = n56249 & ~n56326 ;
  assign n56328 = ~n56222 & n56327 ;
  assign n56329 = ~\pi0200  & \pi1049  ;
  assign n56330 = \pi0200  & \pi1036  ;
  assign n56331 = ~n56329 & ~n56330 ;
  assign n56332 = ~n55610 & n56331 ;
  assign n56333 = ~\pi0255  & n55610 ;
  assign n56334 = ~n56332 & ~n56333 ;
  assign n56335 = ~\pi0200  & \pi1048  ;
  assign n56336 = \pi0200  & \pi1070  ;
  assign n56337 = ~n56335 & ~n56336 ;
  assign n56338 = ~n55610 & n56337 ;
  assign n56339 = ~\pi0256  & n55610 ;
  assign n56340 = ~n56338 & ~n56339 ;
  assign n56341 = ~\pi0200  & \pi1084  ;
  assign n56342 = \pi0200  & \pi1065  ;
  assign n56343 = ~n56341 & ~n56342 ;
  assign n56344 = ~n55610 & n56343 ;
  assign n56345 = ~\pi0257  & n55610 ;
  assign n56346 = ~n56344 & ~n56345 ;
  assign n56347 = ~\pi0200  & \pi1072  ;
  assign n56348 = \pi0200  & \pi1062  ;
  assign n56349 = ~n56347 & ~n56348 ;
  assign n56350 = ~n55610 & n56349 ;
  assign n56351 = ~\pi0258  & n55610 ;
  assign n56352 = ~n56350 & ~n56351 ;
  assign n56353 = ~\pi0200  & \pi1059  ;
  assign n56354 = \pi0200  & \pi1069  ;
  assign n56355 = ~n56353 & ~n56354 ;
  assign n56356 = ~n55610 & n56355 ;
  assign n56357 = ~\pi0259  & n55610 ;
  assign n56358 = ~n56356 & ~n56357 ;
  assign n56359 = \pi0200  & \pi1067  ;
  assign n56360 = ~\pi0200  & \pi1044  ;
  assign n56361 = ~\pi0199  & ~n56360 ;
  assign n56362 = ~n56359 & n56361 ;
  assign n56363 = ~n55610 & ~n56362 ;
  assign n56364 = \pi0260  & n55610 ;
  assign n56365 = ~n56363 & ~n56364 ;
  assign n56366 = \pi0200  & \pi1040  ;
  assign n56367 = ~\pi0200  & \pi1037  ;
  assign n56368 = ~\pi0199  & ~n56367 ;
  assign n56369 = ~n56366 & n56368 ;
  assign n56370 = ~n55610 & ~n56369 ;
  assign n56371 = \pi0261  & n55610 ;
  assign n56372 = ~n56370 & ~n56371 ;
  assign n56373 = ~\pi0299  & ~n50876 ;
  assign n56374 = ~\pi0228  & ~\pi1093  ;
  assign n56375 = \pi0123  & \pi0228  ;
  assign n56376 = ~n56374 & ~n56375 ;
  assign n56377 = ~\pi0262  & ~n56376 ;
  assign n56378 = ~n56373 & ~n56377 ;
  assign n56379 = ~n53066 & n56378 ;
  assign n56380 = n9948 & ~n56379 ;
  assign n56381 = \pi1093  & \pi1142  ;
  assign n56382 = ~\pi0262  & ~\pi1093  ;
  assign n56383 = ~n56381 & ~n56382 ;
  assign n56384 = ~\pi0228  & ~n56383 ;
  assign n56385 = \pi0123  & \pi0262  ;
  assign n56386 = ~\pi0123  & ~\pi1142  ;
  assign n56387 = \pi0228  & ~n56386 ;
  assign n56388 = ~n56385 & n56387 ;
  assign n56389 = ~n56384 & ~n56388 ;
  assign n56390 = ~n52704 & n56376 ;
  assign n56391 = ~n56389 & ~n56390 ;
  assign n56392 = n13558 & n56376 ;
  assign n56393 = ~n51972 & ~n56392 ;
  assign n56394 = ~n56391 & ~n56393 ;
  assign n56395 = ~n50418 & ~n53066 ;
  assign n56396 = n56389 & ~n56395 ;
  assign n56397 = ~n56394 & ~n56396 ;
  assign n56398 = n56380 & n56397 ;
  assign n56399 = ~n51169 & n56376 ;
  assign n56400 = ~n9948 & ~n56389 ;
  assign n56401 = ~n56399 & n56400 ;
  assign n56402 = ~n56398 & ~n56401 ;
  assign n56403 = ~\pi0211  & ~n50394 ;
  assign n56404 = n51622 & n56403 ;
  assign n56405 = ~n50390 & n50627 ;
  assign n56406 = ~\pi0219  & ~n56405 ;
  assign n56407 = ~n56404 & n56406 ;
  assign n56408 = ~\pi0200  & ~\pi1154  ;
  assign n56409 = ~n50394 & ~n56408 ;
  assign n56410 = n43637 & n56409 ;
  assign n56411 = n50383 & n50475 ;
  assign n56412 = ~n50435 & ~n56411 ;
  assign n56413 = ~n56410 & n56412 ;
  assign n56414 = \pi0211  & ~n56413 ;
  assign n56415 = n56407 & ~n56414 ;
  assign n56416 = ~n56410 & ~n56411 ;
  assign n56417 = \pi1156  & n52000 ;
  assign n56418 = \pi0219  & ~n56417 ;
  assign n56419 = n56416 & n56418 ;
  assign n56420 = n9948 & ~n56419 ;
  assign n56421 = ~n56415 & n56420 ;
  assign n56422 = ~\pi0219  & ~n50613 ;
  assign n56423 = ~n50627 & n56422 ;
  assign n56424 = \pi0219  & ~n50612 ;
  assign n56425 = ~n9948 & ~n56424 ;
  assign n56426 = ~n56423 & n56425 ;
  assign n56427 = \pi0230  & ~n56426 ;
  assign n56428 = ~n56421 & n56427 ;
  assign n56429 = ~n50388 & n56042 ;
  assign n56430 = ~n51019 & n56429 ;
  assign n56431 = ~\pi1156  & ~n56430 ;
  assign n56432 = n50511 & n55608 ;
  assign n56433 = n55744 & ~n56432 ;
  assign n56434 = ~n51307 & n56433 ;
  assign n56435 = ~\pi0219  & ~n56434 ;
  assign n56436 = n56431 & n56435 ;
  assign n56437 = \pi1155  & ~n50840 ;
  assign n56438 = n53866 & ~n56437 ;
  assign n56439 = ~n51585 & n56186 ;
  assign n56440 = ~n56438 & ~n56439 ;
  assign n56441 = ~\pi0211  & ~n56440 ;
  assign n56442 = ~\pi0199  & ~\pi1154  ;
  assign n56443 = n44032 & ~n56442 ;
  assign n56444 = n55744 & ~n56443 ;
  assign n56445 = ~n51307 & n56444 ;
  assign n56446 = ~\pi0219  & \pi1156  ;
  assign n56447 = ~n56445 & n56446 ;
  assign n56448 = ~n56441 & n56447 ;
  assign n56449 = ~n56436 & ~n56448 ;
  assign n56450 = ~n53896 & n56440 ;
  assign n56451 = n50618 & ~n56450 ;
  assign n56452 = ~\pi1154  & ~n50385 ;
  assign n56453 = \pi1091  & n50612 ;
  assign n56454 = n44035 & ~n50387 ;
  assign n56455 = \pi1154  & ~n56454 ;
  assign n56456 = n56453 & ~n56455 ;
  assign n56457 = ~n56452 & n56456 ;
  assign n56458 = \pi1091  & ~n56432 ;
  assign n56459 = ~\pi1156  & ~n50388 ;
  assign n56460 = n56458 & n56459 ;
  assign n56461 = \pi0219  & ~n56460 ;
  assign n56462 = ~n56457 & n56461 ;
  assign n56463 = ~n56451 & n56462 ;
  assign n56464 = n56449 & ~n56463 ;
  assign n56465 = ~\pi0263  & ~n56464 ;
  assign n56466 = \pi0263  & \pi1091  ;
  assign n56467 = ~\pi0299  & ~n50391 ;
  assign n56468 = ~\pi0199  & \pi1154  ;
  assign n56469 = n51621 & ~n56468 ;
  assign n56470 = n56467 & ~n56469 ;
  assign n56471 = n56418 & ~n56470 ;
  assign n56472 = ~n56407 & ~n56471 ;
  assign n56473 = ~\pi1155  & ~n50390 ;
  assign n56474 = n56452 & ~n56473 ;
  assign n56475 = \pi1154  & \pi1155  ;
  assign n56476 = ~n13558 & n56475 ;
  assign n56477 = \pi1154  & n44032 ;
  assign n56478 = \pi1156  & ~n56477 ;
  assign n56479 = ~n56476 & n56478 ;
  assign n56480 = ~n56474 & n56479 ;
  assign n56481 = n53856 & ~n56432 ;
  assign n56482 = ~n51307 & n56481 ;
  assign n56483 = \pi0211  & ~n56482 ;
  assign n56484 = ~n56471 & n56483 ;
  assign n56485 = ~n56480 & n56484 ;
  assign n56486 = ~n56472 & ~n56485 ;
  assign n56487 = n56466 & ~n56486 ;
  assign n56488 = n9948 & ~n56487 ;
  assign n56489 = ~n56465 & n56488 ;
  assign n56490 = n9948 & ~n53905 ;
  assign n56491 = \pi1091  & n56424 ;
  assign n56492 = \pi1091  & ~n50627 ;
  assign n56493 = n56422 & n56492 ;
  assign n56494 = ~n56491 & ~n56493 ;
  assign n56495 = \pi0263  & ~\pi1091  ;
  assign n56496 = ~n53905 & ~n56495 ;
  assign n56497 = n56494 & n56496 ;
  assign n56498 = ~n56490 & ~n56497 ;
  assign n56499 = ~n56489 & ~n56498 ;
  assign n56500 = ~\pi0230  & ~n56499 ;
  assign n56501 = \pi0267  & n53732 ;
  assign n56502 = ~n56495 & ~n56501 ;
  assign n56503 = n53905 & n56502 ;
  assign n56504 = n56494 & n56503 ;
  assign n56505 = ~n56304 & ~n56504 ;
  assign n56506 = \pi0211  & ~n53543 ;
  assign n56507 = ~n53567 & n56506 ;
  assign n56508 = ~\pi0211  & ~n56186 ;
  assign n56509 = ~n50613 & ~n56508 ;
  assign n56510 = ~\pi0219  & n56509 ;
  assign n56511 = ~n55874 & ~n56510 ;
  assign n56512 = ~n56507 & ~n56511 ;
  assign n56513 = ~\pi0263  & ~n56309 ;
  assign n56514 = ~n56512 & n56513 ;
  assign n56515 = \pi0211  & ~n53561 ;
  assign n56516 = \pi0211  & ~\pi1091  ;
  assign n56517 = ~n53558 & n56516 ;
  assign n56518 = ~n56515 & ~n56517 ;
  assign n56519 = ~n50613 & ~n56043 ;
  assign n56520 = n56518 & ~n56519 ;
  assign n56521 = n55991 & ~n56520 ;
  assign n56522 = \pi0263  & ~n55864 ;
  assign n56523 = ~n56521 & n56522 ;
  assign n56524 = ~n56514 & ~n56523 ;
  assign n56525 = ~n50612 & n55762 ;
  assign n56526 = n53905 & ~n56525 ;
  assign n56527 = n56501 & n56526 ;
  assign n56528 = ~n56524 & n56527 ;
  assign n56529 = n56505 & ~n56528 ;
  assign n56530 = n56500 & n56529 ;
  assign n56531 = ~\pi1154  & ~\pi1155  ;
  assign n56532 = ~\pi1154  & ~n53568 ;
  assign n56533 = ~n53575 & n56532 ;
  assign n56534 = ~n56531 & ~n56533 ;
  assign n56535 = ~\pi1156  & n56534 ;
  assign n56536 = ~\pi1091  & ~\pi1155  ;
  assign n56537 = ~n53770 & n56536 ;
  assign n56538 = ~\pi1156  & ~n53678 ;
  assign n56539 = n56537 & n56538 ;
  assign n56540 = ~n56535 & ~n56539 ;
  assign n56541 = \pi1155  & n56003 ;
  assign n56542 = \pi1154  & ~n53619 ;
  assign n56543 = ~n56541 & n56542 ;
  assign n56544 = ~n53575 & n56088 ;
  assign n56545 = ~n56531 & ~n56544 ;
  assign n56546 = ~n56537 & ~n56545 ;
  assign n56547 = ~n56543 & ~n56546 ;
  assign n56548 = ~n56540 & n56547 ;
  assign n56549 = n53750 & ~n56545 ;
  assign n56550 = ~n53619 & n56011 ;
  assign n56551 = ~n56541 & n56550 ;
  assign n56552 = ~n56549 & ~n56551 ;
  assign n56553 = ~\pi1154  & n53640 ;
  assign n56554 = ~n53611 & n56553 ;
  assign n56555 = ~\pi0299  & ~\pi1154  ;
  assign n56556 = ~\pi1154  & n53542 ;
  assign n56557 = n53540 & n56556 ;
  assign n56558 = ~n56555 & ~n56557 ;
  assign n56559 = n53612 & ~n56558 ;
  assign n56560 = ~n56554 & ~n56559 ;
  assign n56561 = \pi1156  & n56560 ;
  assign n56562 = n56552 & n56561 ;
  assign n56563 = ~\pi0211  & ~n56562 ;
  assign n56564 = ~n56548 & n56563 ;
  assign n56565 = \pi1154  & ~n53569 ;
  assign n56566 = ~n53587 & n56565 ;
  assign n56567 = ~n56541 & n56566 ;
  assign n56568 = ~n56540 & ~n56567 ;
  assign n56569 = \pi1156  & ~n56554 ;
  assign n56570 = ~n56559 & n56569 ;
  assign n56571 = ~n56096 & n56565 ;
  assign n56572 = ~n56541 & n56571 ;
  assign n56573 = n56570 & ~n56572 ;
  assign n56574 = \pi0211  & ~n56573 ;
  assign n56575 = ~n56568 & n56574 ;
  assign n56576 = ~\pi0219  & ~n56575 ;
  assign n56577 = ~n56564 & n56576 ;
  assign n56578 = \pi1155  & ~n53573 ;
  assign n56579 = n53564 & n56578 ;
  assign n56580 = ~n53554 & n56579 ;
  assign n56581 = \pi1154  & ~n56580 ;
  assign n56582 = ~n56021 & n56581 ;
  assign n56583 = ~n56546 & ~n56582 ;
  assign n56584 = ~\pi1156  & ~n56583 ;
  assign n56585 = ~n56021 & ~n56096 ;
  assign n56586 = n56581 & n56585 ;
  assign n56587 = n50618 & n56586 ;
  assign n56588 = n50618 & n53750 ;
  assign n56589 = ~n56545 & n56588 ;
  assign n56590 = ~n56587 & ~n56589 ;
  assign n56591 = ~\pi1154  & ~n53591 ;
  assign n56592 = ~n53677 & n56591 ;
  assign n56593 = n53804 & ~n56592 ;
  assign n56594 = n50612 & ~n56580 ;
  assign n56595 = ~n56593 & n56594 ;
  assign n56596 = \pi0219  & ~n56595 ;
  assign n56597 = n56590 & n56596 ;
  assign n56598 = ~n56584 & n56597 ;
  assign n56599 = ~\pi0263  & ~n56598 ;
  assign n56600 = ~n56577 & n56599 ;
  assign n56601 = ~\pi1155  & ~n53660 ;
  assign n56602 = ~n53581 & ~n53677 ;
  assign n56603 = n50608 & n56602 ;
  assign n56604 = ~n56601 & ~n56603 ;
  assign n56605 = n50613 & ~n56096 ;
  assign n56606 = n53678 & n56605 ;
  assign n56607 = \pi1156  & ~n53564 ;
  assign n56608 = \pi1156  & n53538 ;
  assign n56609 = ~n53553 & n56608 ;
  assign n56610 = ~n56607 & ~n56609 ;
  assign n56611 = ~n56003 & ~n56610 ;
  assign n56612 = ~n56606 & ~n56611 ;
  assign n56613 = n56604 & n56612 ;
  assign n56614 = ~\pi1154  & ~n56613 ;
  assign n56615 = ~n53611 & n53713 ;
  assign n56616 = n53570 & ~n53611 ;
  assign n56617 = ~n53566 & n56616 ;
  assign n56618 = ~n56615 & ~n56617 ;
  assign n56619 = ~\pi1156  & n56618 ;
  assign n56620 = \pi0211  & ~\pi1155  ;
  assign n56621 = ~\pi0299  & n56620 ;
  assign n56622 = n53542 & n56620 ;
  assign n56623 = n53540 & n56622 ;
  assign n56624 = ~n56621 & ~n56623 ;
  assign n56625 = ~n53564 & ~n56624 ;
  assign n56626 = n53538 & ~n56624 ;
  assign n56627 = ~n53553 & n56626 ;
  assign n56628 = ~n56625 & ~n56627 ;
  assign n56629 = ~\pi0211  & ~\pi1155  ;
  assign n56630 = ~n53569 & n56629 ;
  assign n56631 = ~n53702 & n56630 ;
  assign n56632 = n56628 & ~n56631 ;
  assign n56633 = ~n53571 & n56632 ;
  assign n56634 = \pi1154  & ~n56633 ;
  assign n56635 = ~n56619 & n56634 ;
  assign n56636 = ~n56614 & ~n56635 ;
  assign n56637 = ~\pi0219  & ~n56636 ;
  assign n56638 = ~n53585 & n56258 ;
  assign n56639 = ~n50612 & ~n53591 ;
  assign n56640 = ~n53587 & n56639 ;
  assign n56641 = ~n53566 & n56640 ;
  assign n56642 = ~n56638 & ~n56641 ;
  assign n56643 = \pi1155  & ~n53591 ;
  assign n56644 = ~n53677 & n56643 ;
  assign n56645 = n53601 & ~n56644 ;
  assign n56646 = ~\pi1156  & n53677 ;
  assign n56647 = \pi0219  & ~n56646 ;
  assign n56648 = ~n56645 & n56647 ;
  assign n56649 = ~n56642 & n56648 ;
  assign n56650 = \pi1154  & ~n56645 ;
  assign n56651 = \pi0219  & n50612 ;
  assign n56652 = n56650 & n56651 ;
  assign n56653 = ~\pi1154  & ~n56021 ;
  assign n56654 = ~n53566 & n56653 ;
  assign n56655 = ~n56531 & ~n56654 ;
  assign n56656 = ~n53702 & ~n53776 ;
  assign n56657 = ~\pi1155  & ~n56656 ;
  assign n56658 = n56651 & ~n56657 ;
  assign n56659 = ~n56655 & n56658 ;
  assign n56660 = ~n56652 & ~n56659 ;
  assign n56661 = ~n56649 & n56660 ;
  assign n56662 = \pi0263  & n56661 ;
  assign n56663 = ~n56637 & n56662 ;
  assign n56664 = n56501 & ~n56663 ;
  assign n56665 = ~n56600 & n56664 ;
  assign n56666 = ~\pi0263  & ~n56501 ;
  assign n56667 = ~n56464 & n56666 ;
  assign n56668 = n56466 & ~n56501 ;
  assign n56669 = ~n56486 & n56668 ;
  assign n56670 = n9948 & ~n56669 ;
  assign n56671 = ~n56667 & n56670 ;
  assign n56672 = n56500 & n56671 ;
  assign n56673 = ~n56665 & n56672 ;
  assign n56674 = ~n56530 & ~n56673 ;
  assign n56675 = ~n56428 & n56674 ;
  assign n56676 = \pi0314  & ~\pi0796  ;
  assign n56677 = ~\pi1091  & ~n56676 ;
  assign n56678 = ~\pi0081  & ~\pi1091  ;
  assign n56679 = n53533 & n56678 ;
  assign n56680 = ~n56677 & ~n56679 ;
  assign n56681 = ~\pi0081  & \pi0264  ;
  assign n56682 = n53533 & n56681 ;
  assign n56683 = \pi0264  & ~\pi0314  ;
  assign n56684 = \pi0200  & ~n56683 ;
  assign n56685 = ~n56682 & n56684 ;
  assign n56686 = ~n56680 & n56685 ;
  assign n56687 = ~\pi0200  & ~n56683 ;
  assign n56688 = ~n56682 & n56687 ;
  assign n56689 = ~n56680 & n56688 ;
  assign n56690 = \pi1091  & \pi1142  ;
  assign n56691 = \pi0200  & n56690 ;
  assign n56692 = \pi1091  & \pi1141  ;
  assign n56693 = ~\pi0200  & n56692 ;
  assign n56694 = ~\pi0199  & ~n56693 ;
  assign n56695 = ~n56691 & n56694 ;
  assign n56696 = ~n56689 & n56695 ;
  assign n56697 = ~n56686 & n56696 ;
  assign n56698 = \pi0314  & ~n53533 ;
  assign n56699 = \pi0264  & ~n56698 ;
  assign n56700 = ~n53533 & n56676 ;
  assign n56701 = ~\pi1091  & ~n56700 ;
  assign n56702 = ~n56699 & n56701 ;
  assign n56703 = \pi1091  & \pi1143  ;
  assign n56704 = ~\pi0200  & n56703 ;
  assign n56705 = \pi0199  & ~n56704 ;
  assign n56706 = ~n56702 & n56705 ;
  assign n56707 = n20516 & ~n56706 ;
  assign n56708 = ~n56697 & n56707 ;
  assign n56709 = \pi0211  & ~n56683 ;
  assign n56710 = ~n56682 & n56709 ;
  assign n56711 = ~n56680 & n56710 ;
  assign n56712 = ~\pi0211  & ~n56683 ;
  assign n56713 = ~n56682 & n56712 ;
  assign n56714 = ~n56680 & n56713 ;
  assign n56715 = \pi0211  & n56690 ;
  assign n56716 = ~\pi0211  & n56692 ;
  assign n56717 = ~\pi0219  & ~n56716 ;
  assign n56718 = ~n56715 & n56717 ;
  assign n56719 = ~n56714 & n56718 ;
  assign n56720 = ~n56711 & n56719 ;
  assign n56721 = \pi0219  & ~n56042 ;
  assign n56722 = ~n51662 & ~n56721 ;
  assign n56723 = ~n56702 & ~n56722 ;
  assign n56724 = ~n20516 & ~n56723 ;
  assign n56725 = ~n56720 & n56724 ;
  assign n56726 = ~n56708 & ~n56725 ;
  assign n56727 = ~\pi0230  & ~n56726 ;
  assign n56728 = ~\pi0211  & \pi1141  ;
  assign n56729 = ~\pi0219  & ~n56728 ;
  assign n56730 = ~n50663 & n56729 ;
  assign n56731 = ~n51662 & ~n56730 ;
  assign n56732 = ~n20516 & ~n56731 ;
  assign n56733 = \pi0230  & ~n20516 ;
  assign n56734 = ~\pi0199  & \pi1141  ;
  assign n56735 = n51717 & ~n56734 ;
  assign n56736 = \pi0230  & ~n50640 ;
  assign n56737 = ~n56735 & n56736 ;
  assign n56738 = ~n56733 & ~n56737 ;
  assign n56739 = ~n56732 & ~n56738 ;
  assign n56740 = ~n56727 & ~n56739 ;
  assign n56741 = \pi0314  & ~\pi0819  ;
  assign n56742 = ~\pi1091  & ~n56741 ;
  assign n56743 = ~n56679 & ~n56742 ;
  assign n56744 = ~\pi0081  & \pi0265  ;
  assign n56745 = n53533 & n56744 ;
  assign n56746 = \pi0265  & ~\pi0314  ;
  assign n56747 = \pi0200  & ~n56746 ;
  assign n56748 = ~n56745 & n56747 ;
  assign n56749 = ~n56743 & n56748 ;
  assign n56750 = ~\pi0200  & ~n56746 ;
  assign n56751 = ~n56745 & n56750 ;
  assign n56752 = ~n56743 & n56751 ;
  assign n56753 = \pi0200  & n56703 ;
  assign n56754 = ~\pi0200  & n56690 ;
  assign n56755 = ~\pi0199  & ~n56754 ;
  assign n56756 = ~n56753 & n56755 ;
  assign n56757 = ~n56752 & n56756 ;
  assign n56758 = ~n56749 & n56757 ;
  assign n56759 = \pi0265  & ~n56698 ;
  assign n56760 = ~n53533 & n56741 ;
  assign n56761 = ~\pi1091  & ~n56760 ;
  assign n56762 = ~n56759 & n56761 ;
  assign n56763 = \pi1091  & \pi1144  ;
  assign n56764 = ~\pi0200  & n56763 ;
  assign n56765 = \pi0199  & ~n56764 ;
  assign n56766 = ~n56762 & n56765 ;
  assign n56767 = n20516 & ~n56766 ;
  assign n56768 = ~n56758 & n56767 ;
  assign n56769 = \pi0211  & ~n56746 ;
  assign n56770 = ~n56745 & n56769 ;
  assign n56771 = ~n56743 & n56770 ;
  assign n56772 = ~\pi0211  & ~n56746 ;
  assign n56773 = ~n56745 & n56772 ;
  assign n56774 = ~n56743 & n56773 ;
  assign n56775 = \pi0211  & n56703 ;
  assign n56776 = ~\pi0211  & n56690 ;
  assign n56777 = ~\pi0219  & ~n56776 ;
  assign n56778 = ~n56775 & n56777 ;
  assign n56779 = ~n56774 & n56778 ;
  assign n56780 = ~n56771 & n56779 ;
  assign n56781 = ~n53464 & ~n56721 ;
  assign n56782 = ~n56762 & ~n56781 ;
  assign n56783 = ~n20516 & ~n56782 ;
  assign n56784 = ~n56780 & n56783 ;
  assign n56785 = ~n56768 & ~n56784 ;
  assign n56786 = ~\pi0230  & ~n56785 ;
  assign n56787 = ~n50639 & n53428 ;
  assign n56788 = ~n50652 & ~n56787 ;
  assign n56789 = n20516 & ~n56788 ;
  assign n56790 = ~\pi0219  & ~n50657 ;
  assign n56791 = ~n50668 & n56790 ;
  assign n56792 = \pi0230  & ~n53464 ;
  assign n56793 = ~n56791 & n56792 ;
  assign n56794 = ~n53960 & ~n56793 ;
  assign n56795 = ~n56789 & ~n56794 ;
  assign n56796 = ~n56786 & ~n56795 ;
  assign n56797 = \pi0314  & ~\pi0948  ;
  assign n56798 = ~n53534 & n56797 ;
  assign n56799 = ~\pi0081  & ~\pi0266  ;
  assign n56800 = n53533 & n56799 ;
  assign n56801 = ~\pi0266  & ~\pi0314  ;
  assign n56802 = ~\pi1091  & ~n56801 ;
  assign n56803 = ~n56800 & n56802 ;
  assign n56804 = ~n56798 & n56803 ;
  assign n56805 = \pi1091  & \pi1135  ;
  assign n56806 = ~\pi0199  & ~n56805 ;
  assign n56807 = ~n56804 & n56806 ;
  assign n56808 = ~\pi0199  & \pi0200  ;
  assign n56809 = \pi0266  & ~\pi1091  ;
  assign n56810 = \pi0314  & ~\pi1091  ;
  assign n56811 = ~n53533 & n56810 ;
  assign n56812 = ~n56809 & ~n56811 ;
  assign n56813 = ~n53533 & n56797 ;
  assign n56814 = \pi0200  & ~n56813 ;
  assign n56815 = ~n56812 & n56814 ;
  assign n56816 = ~n56808 & ~n56815 ;
  assign n56817 = ~n56807 & ~n56816 ;
  assign n56818 = ~\pi0199  & ~n56804 ;
  assign n56819 = \pi1091  & \pi1136  ;
  assign n56820 = \pi0199  & ~n56819 ;
  assign n56821 = ~\pi0200  & ~n56820 ;
  assign n56822 = ~\pi0200  & ~n56813 ;
  assign n56823 = ~n56812 & n56822 ;
  assign n56824 = ~n56821 & ~n56823 ;
  assign n56825 = ~n56818 & ~n56824 ;
  assign n56826 = ~n56817 & ~n56825 ;
  assign n56827 = ~\pi0211  & \pi1136  ;
  assign n56828 = \pi0219  & ~n56827 ;
  assign n56829 = \pi0211  & ~\pi1135  ;
  assign n56830 = ~n12577 & ~n56829 ;
  assign n56831 = ~n56828 & n56830 ;
  assign n56832 = ~n9948 & n56831 ;
  assign n56833 = \pi0230  & ~n56832 ;
  assign n56834 = n20516 & ~n56833 ;
  assign n56835 = \pi0299  & n56831 ;
  assign n56836 = ~\pi0199  & \pi1135  ;
  assign n56837 = n44035 & n56836 ;
  assign n56838 = \pi0199  & \pi1136  ;
  assign n56839 = n44032 & n56838 ;
  assign n56840 = ~n56837 & ~n56839 ;
  assign n56841 = ~n56835 & n56840 ;
  assign n56842 = n9948 & n20516 ;
  assign n56843 = ~n56841 & n56842 ;
  assign n56844 = ~n56834 & ~n56843 ;
  assign n56845 = ~n56826 & ~n56844 ;
  assign n56846 = n9948 & ~n56841 ;
  assign n56847 = n56833 & ~n56846 ;
  assign n56848 = ~\pi1134  & n56847 ;
  assign n56849 = ~n56812 & ~n56813 ;
  assign n56850 = ~n56721 & ~n56828 ;
  assign n56851 = ~n56849 & ~n56850 ;
  assign n56852 = ~n20516 & ~n56851 ;
  assign n56853 = \pi1135  & n55744 ;
  assign n56854 = ~\pi0219  & ~n56853 ;
  assign n56855 = ~n56804 & n56854 ;
  assign n56856 = n56852 & ~n56855 ;
  assign n56857 = ~\pi0230  & ~\pi1134  ;
  assign n56858 = ~n56856 & n56857 ;
  assign n56859 = ~n56848 & ~n56858 ;
  assign n56860 = ~n56845 & ~n56859 ;
  assign n56861 = \pi1091  & ~n56829 ;
  assign n56862 = ~\pi0219  & ~n56861 ;
  assign n56863 = ~n56804 & n56862 ;
  assign n56864 = n56852 & ~n56863 ;
  assign n56865 = ~\pi0230  & \pi1134  ;
  assign n56866 = ~n56864 & n56865 ;
  assign n56867 = ~\pi0199  & \pi1091  ;
  assign n56868 = n56820 & ~n56867 ;
  assign n56869 = ~n56849 & n56868 ;
  assign n56870 = ~\pi0199  & ~n56867 ;
  assign n56871 = ~n56804 & n56870 ;
  assign n56872 = ~n56869 & ~n56871 ;
  assign n56873 = ~\pi0200  & n20515 ;
  assign n56874 = n6848 & n56873 ;
  assign n56875 = n56872 & n56874 ;
  assign n56876 = n20516 & n56817 ;
  assign n56877 = ~n56875 & ~n56876 ;
  assign n56878 = n56866 & n56877 ;
  assign n56879 = n50383 & ~n56838 ;
  assign n56880 = \pi0200  & ~n56836 ;
  assign n56881 = ~n56879 & ~n56880 ;
  assign n56882 = n20516 & n56881 ;
  assign n56883 = \pi0230  & ~n56882 ;
  assign n56884 = ~n56828 & ~n56829 ;
  assign n56885 = ~n20516 & n56884 ;
  assign n56886 = \pi1134  & ~n56885 ;
  assign n56887 = n56883 & n56886 ;
  assign n56888 = ~n56878 & ~n56887 ;
  assign n56889 = ~n56860 & n56888 ;
  assign n56890 = ~\pi0267  & ~n53556 ;
  assign n56891 = ~n55864 & n56890 ;
  assign n56892 = \pi0267  & ~n55874 ;
  assign n56893 = ~n56309 & n56892 ;
  assign n56894 = n53732 & ~n56893 ;
  assign n56895 = ~n56891 & n56894 ;
  assign n56896 = ~n50609 & ~n50625 ;
  assign n56897 = n53909 & n56896 ;
  assign n56898 = ~n50608 & n55762 ;
  assign n56899 = ~n56897 & ~n56898 ;
  assign n56900 = ~\pi0267  & ~\pi1091  ;
  assign n56901 = ~n53732 & n56900 ;
  assign n56902 = n53905 & ~n56901 ;
  assign n56903 = n56899 & n56902 ;
  assign n56904 = ~n56895 & n56903 ;
  assign n56905 = ~n56304 & ~n56904 ;
  assign n56906 = ~n53569 & ~n53587 ;
  assign n56907 = ~n55898 & ~n56906 ;
  assign n56908 = n53756 & ~n56907 ;
  assign n56909 = \pi1154  & ~n56908 ;
  assign n56910 = ~\pi1154  & n56021 ;
  assign n56911 = n55929 & n56910 ;
  assign n56912 = ~\pi1155  & ~n56911 ;
  assign n56913 = ~n56909 & n56912 ;
  assign n56914 = \pi1155  & n55849 ;
  assign n56915 = n53575 & ~n56592 ;
  assign n56916 = n56914 & ~n56915 ;
  assign n56917 = \pi0267  & ~n56916 ;
  assign n56918 = \pi0267  & ~n53814 ;
  assign n56919 = ~n55926 & n56918 ;
  assign n56920 = ~n56917 & ~n56919 ;
  assign n56921 = ~n56913 & ~n56920 ;
  assign n56922 = ~n56098 & ~n56103 ;
  assign n56923 = ~n53744 & ~n55911 ;
  assign n56924 = ~\pi1154  & ~n56923 ;
  assign n56925 = ~n56922 & n56924 ;
  assign n56926 = \pi0211  & n56925 ;
  assign n56927 = ~n53593 & ~n56112 ;
  assign n56928 = \pi0211  & n56475 ;
  assign n56929 = n56927 & n56928 ;
  assign n56930 = ~n56926 & ~n56929 ;
  assign n56931 = \pi1153  & n53597 ;
  assign n56932 = n50608 & ~n56931 ;
  assign n56933 = n53776 & n56932 ;
  assign n56934 = n50608 & n53702 ;
  assign n56935 = ~n56933 & ~n56934 ;
  assign n56936 = ~n56023 & ~n56935 ;
  assign n56937 = ~\pi0267  & ~n56936 ;
  assign n56938 = n53770 & ~n56013 ;
  assign n56939 = ~\pi1155  & ~n56938 ;
  assign n56940 = ~n56922 & n56939 ;
  assign n56941 = n56937 & ~n56940 ;
  assign n56942 = n56930 & n56941 ;
  assign n56943 = ~n56921 & ~n56942 ;
  assign n56944 = \pi0219  & ~n56943 ;
  assign n56945 = ~n56905 & n56944 ;
  assign n56946 = \pi1154  & n53616 ;
  assign n56947 = ~n56908 & n56946 ;
  assign n56948 = \pi1155  & n56021 ;
  assign n56949 = \pi1155  & ~n53554 ;
  assign n56950 = n53565 & n56949 ;
  assign n56951 = ~n56948 & ~n56950 ;
  assign n56952 = \pi1154  & n56951 ;
  assign n56953 = ~n53564 & ~n53568 ;
  assign n56954 = ~n53645 & ~n56953 ;
  assign n56955 = ~n53586 & ~n56558 ;
  assign n56956 = n53538 & ~n56558 ;
  assign n56957 = ~n53553 & n56956 ;
  assign n56958 = ~n56955 & ~n56957 ;
  assign n56959 = \pi1155  & ~n50460 ;
  assign n56960 = n56958 & n56959 ;
  assign n56961 = ~n56954 & ~n56960 ;
  assign n56962 = ~n56952 & ~n56961 ;
  assign n56963 = ~n56947 & n56962 ;
  assign n56964 = n53678 & ~n56096 ;
  assign n56965 = ~\pi1155  & ~n56964 ;
  assign n56966 = ~n56922 & n56965 ;
  assign n56967 = \pi0211  & ~n56966 ;
  assign n56968 = ~n56963 & n56967 ;
  assign n56969 = ~\pi1154  & ~n55922 ;
  assign n56970 = ~n50510 & ~n53569 ;
  assign n56971 = ~n53677 & n56970 ;
  assign n56972 = ~n56051 & ~n56971 ;
  assign n56973 = ~n56969 & ~n56972 ;
  assign n56974 = \pi1153  & ~\pi1155  ;
  assign n56975 = \pi1154  & ~n56974 ;
  assign n56976 = n56602 & n56975 ;
  assign n56977 = ~\pi1155  & ~n56976 ;
  assign n56978 = ~n56973 & n56977 ;
  assign n56979 = ~n53702 & ~n56003 ;
  assign n56980 = \pi1155  & ~n56931 ;
  assign n56981 = \pi1155  & n53564 ;
  assign n56982 = ~n53554 & n56981 ;
  assign n56983 = ~n56980 & ~n56982 ;
  assign n56984 = ~n56979 & ~n56983 ;
  assign n56985 = ~n56976 & n56984 ;
  assign n56986 = ~\pi0211  & ~n56985 ;
  assign n56987 = ~n56978 & n56986 ;
  assign n56988 = ~\pi0267  & ~n56987 ;
  assign n56989 = ~n56968 & n56988 ;
  assign n56990 = ~\pi1154  & ~n55898 ;
  assign n56991 = ~n53569 & ~n56096 ;
  assign n56992 = n53619 & ~n56991 ;
  assign n56993 = n56990 & n56992 ;
  assign n56994 = \pi1155  & n53569 ;
  assign n56995 = n50419 & ~n53585 ;
  assign n56996 = ~n56994 & ~n56995 ;
  assign n56997 = n56990 & ~n56996 ;
  assign n56998 = ~n56993 & ~n56997 ;
  assign n56999 = \pi0211  & ~n56998 ;
  assign n57000 = ~\pi1155  & ~n53568 ;
  assign n57001 = ~n53575 & n57000 ;
  assign n57002 = \pi1154  & ~n57001 ;
  assign n57003 = ~n53702 & n55897 ;
  assign n57004 = \pi1154  & n56003 ;
  assign n57005 = ~n57003 & n57004 ;
  assign n57006 = ~n57002 & ~n57005 ;
  assign n57007 = ~n53568 & n53612 ;
  assign n57008 = n56914 & n57007 ;
  assign n57009 = \pi0211  & ~n57008 ;
  assign n57010 = ~n57006 & n57009 ;
  assign n57011 = ~n56999 & ~n57010 ;
  assign n57012 = \pi1154  & ~n53573 ;
  assign n57013 = n53564 & n57012 ;
  assign n57014 = ~n53554 & n57013 ;
  assign n57015 = \pi1155  & ~n57014 ;
  assign n57016 = ~\pi0211  & ~n57015 ;
  assign n57017 = ~\pi0211  & n53581 ;
  assign n57018 = ~n56278 & n57017 ;
  assign n57019 = ~n57016 & ~n57018 ;
  assign n57020 = \pi0267  & n57019 ;
  assign n57021 = ~\pi1154  & n53619 ;
  assign n57022 = ~n55898 & n57021 ;
  assign n57023 = ~\pi1155  & ~n57022 ;
  assign n57024 = \pi0267  & ~n57005 ;
  assign n57025 = n57023 & n57024 ;
  assign n57026 = ~n57020 & ~n57025 ;
  assign n57027 = n57011 & ~n57026 ;
  assign n57028 = ~n56989 & ~n57027 ;
  assign n57029 = ~\pi0219  & ~n56905 ;
  assign n57030 = n57028 & n57029 ;
  assign n57031 = ~n56945 & ~n57030 ;
  assign n57032 = n53732 & ~n57031 ;
  assign n57033 = ~n51983 & n56186 ;
  assign n57034 = \pi0219  & ~n57033 ;
  assign n57035 = \pi0219  & \pi1155  ;
  assign n57036 = ~n44035 & n57035 ;
  assign n57037 = ~n52037 & n57036 ;
  assign n57038 = ~n57034 & ~n57037 ;
  assign n57039 = \pi1091  & ~n55734 ;
  assign n57040 = n56437 & n57039 ;
  assign n57041 = n43637 & ~n51013 ;
  assign n57042 = \pi1091  & \pi1154  ;
  assign n57043 = ~n57041 & n57042 ;
  assign n57044 = ~n57040 & n57043 ;
  assign n57045 = ~\pi0211  & ~n57044 ;
  assign n57046 = ~n57038 & n57045 ;
  assign n57047 = \pi1091  & ~n51585 ;
  assign n57048 = ~\pi1153  & \pi1155  ;
  assign n57049 = n50419 & n53865 ;
  assign n57050 = ~n57048 & ~n57049 ;
  assign n57051 = \pi1154  & ~n57050 ;
  assign n57052 = n57047 & n57051 ;
  assign n57053 = ~\pi1153  & ~\pi1155  ;
  assign n57054 = n50458 & n53846 ;
  assign n57055 = ~n57053 & ~n57054 ;
  assign n57056 = \pi1154  & ~n55735 ;
  assign n57057 = ~n55788 & n57056 ;
  assign n57058 = ~n57055 & n57057 ;
  assign n57059 = n51215 & n56186 ;
  assign n57060 = ~\pi0299  & n56186 ;
  assign n57061 = ~n50487 & n57060 ;
  assign n57062 = ~n57059 & ~n57061 ;
  assign n57063 = ~n57058 & n57062 ;
  assign n57064 = ~n57052 & n57063 ;
  assign n57065 = n12577 & n57064 ;
  assign n57066 = ~n57046 & ~n57065 ;
  assign n57067 = n50458 & ~n51014 ;
  assign n57068 = ~n50371 & n50419 ;
  assign n57069 = ~n57067 & ~n57068 ;
  assign n57070 = ~n53974 & n57069 ;
  assign n57071 = ~n50370 & n50419 ;
  assign n57072 = ~n51007 & n57071 ;
  assign n57073 = n57042 & ~n57072 ;
  assign n57074 = ~n57070 & n57073 ;
  assign n57075 = ~n50420 & n57033 ;
  assign n57076 = \pi0211  & ~n57075 ;
  assign n57077 = ~n57074 & n57076 ;
  assign n57078 = n57066 & ~n57077 ;
  assign n57079 = \pi0267  & ~n57078 ;
  assign n57080 = ~\pi0299  & n50405 ;
  assign n57081 = n44035 & ~n56468 ;
  assign n57082 = ~n57080 & ~n57081 ;
  assign n57083 = ~n51219 & n57082 ;
  assign n57084 = \pi1091  & n57083 ;
  assign n57085 = ~\pi0211  & ~n57084 ;
  assign n57086 = \pi1091  & ~\pi1155  ;
  assign n57087 = n50609 & ~n57086 ;
  assign n57088 = ~\pi0299  & n50609 ;
  assign n57089 = ~n51014 & n57088 ;
  assign n57090 = ~n57087 & ~n57089 ;
  assign n57091 = ~n57040 & ~n57090 ;
  assign n57092 = ~\pi0219  & ~n57091 ;
  assign n57093 = ~n57085 & n57092 ;
  assign n57094 = n57041 & n57086 ;
  assign n57095 = \pi1154  & ~n57094 ;
  assign n57096 = ~n57040 & n57095 ;
  assign n57097 = \pi1154  & ~n57096 ;
  assign n57098 = ~\pi1155  & ~n50384 ;
  assign n57099 = ~n44035 & n56186 ;
  assign n57100 = ~n52037 & n57099 ;
  assign n57101 = ~n57098 & n57100 ;
  assign n57102 = ~\pi0211  & ~n57101 ;
  assign n57103 = ~n57097 & n57102 ;
  assign n57104 = ~n50840 & n56475 ;
  assign n57105 = ~n51008 & n57104 ;
  assign n57106 = \pi0219  & ~n57105 ;
  assign n57107 = ~n57096 & n57106 ;
  assign n57108 = ~n50689 & ~n57107 ;
  assign n57109 = ~n57103 & ~n57108 ;
  assign n57110 = ~n57093 & ~n57109 ;
  assign n57111 = \pi0211  & ~\pi1154  ;
  assign n57112 = \pi1091  & ~n51001 ;
  assign n57113 = n44032 & n57112 ;
  assign n57114 = n57111 & ~n57113 ;
  assign n57115 = ~\pi0267  & ~n57111 ;
  assign n57116 = n50458 & ~n55608 ;
  assign n57117 = ~\pi0267  & ~n57053 ;
  assign n57118 = ~n57116 & n57117 ;
  assign n57119 = ~n57115 & ~n57118 ;
  assign n57120 = ~n57114 & ~n57119 ;
  assign n57121 = ~n57110 & n57120 ;
  assign n57122 = ~n57079 & ~n57121 ;
  assign n57123 = ~n53732 & ~n57122 ;
  assign n57124 = n9948 & ~n57123 ;
  assign n57125 = ~n56905 & ~n57124 ;
  assign n57126 = ~n53905 & ~n56900 ;
  assign n57127 = n56899 & n57126 ;
  assign n57128 = ~\pi0230  & ~n56490 ;
  assign n57129 = ~n57127 & n57128 ;
  assign n57130 = ~\pi0057  & ~\pi0230  ;
  assign n57131 = n6848 & n57130 ;
  assign n57132 = n57122 & n57131 ;
  assign n57133 = ~n57129 & ~n57132 ;
  assign n57134 = ~n57125 & ~n57133 ;
  assign n57135 = ~n57032 & n57134 ;
  assign n57136 = \pi1155  & n52040 ;
  assign n57137 = ~\pi1154  & ~n51983 ;
  assign n57138 = ~n51924 & ~n57137 ;
  assign n57139 = ~n57136 & ~n57138 ;
  assign n57140 = \pi0219  & ~n51008 ;
  assign n57141 = \pi0211  & ~n57140 ;
  assign n57142 = ~n57139 & n57141 ;
  assign n57143 = ~\pi0219  & ~n57083 ;
  assign n57144 = \pi0219  & ~n50435 ;
  assign n57145 = ~\pi0211  & ~n57144 ;
  assign n57146 = ~n50433 & ~n51007 ;
  assign n57147 = \pi0200  & ~n56468 ;
  assign n57148 = ~\pi0211  & ~n57147 ;
  assign n57149 = n57146 & n57148 ;
  assign n57150 = ~n57145 & ~n57149 ;
  assign n57151 = ~n57143 & ~n57150 ;
  assign n57152 = ~n57142 & ~n57151 ;
  assign n57153 = n9948 & ~n57152 ;
  assign n57154 = \pi0219  & ~n50608 ;
  assign n57155 = ~\pi0219  & ~n50609 ;
  assign n57156 = ~n50625 & n57155 ;
  assign n57157 = ~n57154 & ~n57156 ;
  assign n57158 = ~n9948 & n57157 ;
  assign n57159 = \pi0230  & ~n57158 ;
  assign n57160 = ~n57153 & n57159 ;
  assign n57161 = ~n57135 & ~n57160 ;
  assign n57162 = n43637 & n51996 ;
  assign n57163 = n6848 & n57162 ;
  assign n57164 = ~n20516 & n53137 ;
  assign n57165 = ~n57163 & ~n57164 ;
  assign n57166 = ~\pi0211  & ~n20516 ;
  assign n57167 = ~\pi0057  & n44032 ;
  assign n57168 = n6848 & n57167 ;
  assign n57169 = ~n57166 & ~n57168 ;
  assign n57170 = n57165 & n57169 ;
  assign n57171 = ~\pi0057  & n43637 ;
  assign n57172 = n6848 & n57171 ;
  assign n57173 = ~\pi1152  & ~n57172 ;
  assign n57174 = ~n54850 & n57173 ;
  assign n57175 = \pi0230  & \pi1150  ;
  assign n57176 = ~n57174 & n57175 ;
  assign n57177 = ~n57170 & n57176 ;
  assign n57178 = n9948 & ~n13649 ;
  assign n57179 = n13647 & ~n55740 ;
  assign n57180 = ~n57178 & ~n57179 ;
  assign n57181 = \pi1151  & ~n57180 ;
  assign n57182 = ~\pi1152  & ~n57181 ;
  assign n57183 = ~\pi1151  & n55693 ;
  assign n57184 = ~\pi1150  & ~n57183 ;
  assign n57185 = ~n57182 & n57184 ;
  assign n57186 = ~n20516 & n55799 ;
  assign n57187 = n50432 & n55740 ;
  assign n57188 = ~n57186 & ~n57187 ;
  assign n57189 = n52250 & ~n57188 ;
  assign n57190 = \pi0230  & ~n57189 ;
  assign n57191 = n57185 & n57190 ;
  assign n57192 = ~n57177 & ~n57191 ;
  assign n57193 = \pi0230  & n57192 ;
  assign n57194 = ~n9948 & ~n55864 ;
  assign n57195 = n56319 & n57194 ;
  assign n57196 = ~n9948 & ~n57195 ;
  assign n57197 = \pi0219  & ~n53586 ;
  assign n57198 = \pi0219  & ~n53578 ;
  assign n57199 = ~n53553 & n57198 ;
  assign n57200 = ~n57197 & ~n57199 ;
  assign n57201 = n55888 & ~n57200 ;
  assign n57202 = ~n53591 & ~n57200 ;
  assign n57203 = ~n53566 & n57202 ;
  assign n57204 = ~n57201 & ~n57203 ;
  assign n57205 = ~n53566 & n55846 ;
  assign n57206 = ~n57195 & ~n57205 ;
  assign n57207 = n57204 & n57206 ;
  assign n57208 = ~n57196 & ~n57207 ;
  assign n57209 = \pi1151  & ~n57208 ;
  assign n57210 = ~n53566 & n55930 ;
  assign n57211 = \pi0219  & n55888 ;
  assign n57212 = ~n53566 & n56297 ;
  assign n57213 = ~n57211 & ~n57212 ;
  assign n57214 = ~n57210 & n57213 ;
  assign n57215 = ~\pi0219  & n56954 ;
  assign n57216 = ~n55911 & ~n57215 ;
  assign n57217 = n55740 & n57216 ;
  assign n57218 = ~n57214 & n57217 ;
  assign n57219 = ~n9948 & ~n55991 ;
  assign n57220 = ~n55864 & n57219 ;
  assign n57221 = ~\pi1151  & ~n57220 ;
  assign n57222 = ~n57218 & n57221 ;
  assign n57223 = ~n57209 & ~n57222 ;
  assign n57224 = \pi1152  & n57223 ;
  assign n57225 = n9948 & ~n57205 ;
  assign n57226 = n57204 & n57225 ;
  assign n57227 = ~n53611 & n55930 ;
  assign n57228 = n9948 & n53804 ;
  assign n57229 = ~n57227 & n57228 ;
  assign n57230 = \pi0219  & ~n55740 ;
  assign n57231 = ~n53590 & n57230 ;
  assign n57232 = n52628 & n55875 ;
  assign n57233 = ~\pi1091  & n52628 ;
  assign n57234 = n53555 & n57233 ;
  assign n57235 = ~n57232 & ~n57234 ;
  assign n57236 = ~n57231 & n57235 ;
  assign n57237 = n53117 & n57236 ;
  assign n57238 = ~n53664 & n55740 ;
  assign n57239 = ~n53662 & n57238 ;
  assign n57240 = n55919 & n57239 ;
  assign n57241 = ~n55991 & ~n57231 ;
  assign n57242 = ~\pi1152  & n57241 ;
  assign n57243 = n57236 & n57242 ;
  assign n57244 = ~n57240 & n57243 ;
  assign n57245 = ~n57237 & ~n57244 ;
  assign n57246 = ~n57229 & ~n57245 ;
  assign n57247 = ~n57226 & n57246 ;
  assign n57248 = ~\pi1151  & n57242 ;
  assign n57249 = ~n57240 & n57248 ;
  assign n57250 = ~\pi0268  & ~n57249 ;
  assign n57251 = ~n57247 & n57250 ;
  assign n57252 = ~n57224 & n57251 ;
  assign n57253 = ~n9948 & n56309 ;
  assign n57254 = ~n9948 & ~n55992 ;
  assign n57255 = n55844 & n57254 ;
  assign n57256 = ~n57253 & ~n57255 ;
  assign n57257 = ~n9948 & ~n56309 ;
  assign n57258 = ~n55993 & n57257 ;
  assign n57259 = n53612 & ~n57258 ;
  assign n57260 = n57256 & ~n57259 ;
  assign n57261 = \pi0219  & n53814 ;
  assign n57262 = \pi0219  & n55839 ;
  assign n57263 = n55835 & n57262 ;
  assign n57264 = ~n57261 & ~n57263 ;
  assign n57265 = ~n55902 & n57256 ;
  assign n57266 = n57264 & n57265 ;
  assign n57267 = ~n57260 & ~n57266 ;
  assign n57268 = \pi1151  & n57267 ;
  assign n57269 = n9948 & ~n57227 ;
  assign n57270 = n57264 & n57269 ;
  assign n57271 = ~n55844 & n57257 ;
  assign n57272 = ~\pi1151  & ~n57271 ;
  assign n57273 = ~n57270 & n57272 ;
  assign n57274 = \pi1152  & ~n57273 ;
  assign n57275 = ~n57268 & n57274 ;
  assign n57276 = ~n9948 & ~n56213 ;
  assign n57277 = ~n55993 & n57276 ;
  assign n57278 = n9948 & ~n55980 ;
  assign n57279 = ~n57277 & ~n57278 ;
  assign n57280 = n55844 & ~n57277 ;
  assign n57281 = ~n55901 & n57280 ;
  assign n57282 = ~n57279 & ~n57281 ;
  assign n57283 = \pi1151  & ~n57282 ;
  assign n57284 = n9948 & n55919 ;
  assign n57285 = ~n53567 & ~n55829 ;
  assign n57286 = ~n53567 & n53586 ;
  assign n57287 = ~n53554 & n57286 ;
  assign n57288 = ~n57285 & ~n57287 ;
  assign n57289 = n57284 & ~n57288 ;
  assign n57290 = ~n9948 & ~n55874 ;
  assign n57291 = ~n53567 & n57290 ;
  assign n57292 = ~\pi1151  & ~n57291 ;
  assign n57293 = ~n57289 & n57292 ;
  assign n57294 = ~\pi1152  & ~n57293 ;
  assign n57295 = ~n57283 & n57294 ;
  assign n57296 = \pi0268  & ~n57295 ;
  assign n57297 = ~n57275 & n57296 ;
  assign n57298 = ~n57252 & ~n57297 ;
  assign n57299 = ~\pi1150  & ~n57298 ;
  assign n57300 = \pi0275  & n53903 ;
  assign n57301 = n53120 & ~n56309 ;
  assign n57302 = ~n55876 & n57301 ;
  assign n57303 = ~n53590 & n55839 ;
  assign n57304 = n55835 & n57303 ;
  assign n57305 = ~n53590 & n53803 ;
  assign n57306 = ~\pi1151  & ~n57305 ;
  assign n57307 = ~n57304 & n57306 ;
  assign n57308 = ~n57302 & ~n57307 ;
  assign n57309 = ~n57229 & ~n57302 ;
  assign n57310 = ~n57226 & n57309 ;
  assign n57311 = ~n57308 & ~n57310 ;
  assign n57312 = \pi0268  & ~\pi1151  ;
  assign n57313 = ~n53559 & n55740 ;
  assign n57314 = ~n55926 & n57313 ;
  assign n57315 = n55829 & ~n55911 ;
  assign n57316 = n57284 & ~n57315 ;
  assign n57317 = ~n56309 & n57290 ;
  assign n57318 = ~n57316 & ~n57317 ;
  assign n57319 = \pi0268  & n57318 ;
  assign n57320 = ~n57314 & n57319 ;
  assign n57321 = ~n57312 & ~n57320 ;
  assign n57322 = ~n57311 & ~n57321 ;
  assign n57323 = n51997 & ~n57214 ;
  assign n57324 = ~n55992 & n57194 ;
  assign n57325 = ~n57271 & n57324 ;
  assign n57326 = ~n57195 & ~n57325 ;
  assign n57327 = \pi1151  & ~n57326 ;
  assign n57328 = ~\pi0268  & ~n57327 ;
  assign n57329 = ~n57323 & n57328 ;
  assign n57330 = \pi1152  & ~n57329 ;
  assign n57331 = n9948 & ~n53564 ;
  assign n57332 = n9948 & n53538 ;
  assign n57333 = ~n53553 & n57332 ;
  assign n57334 = ~n57331 & ~n57333 ;
  assign n57335 = n56297 & ~n57334 ;
  assign n57336 = n55844 & ~n57334 ;
  assign n57337 = ~n55901 & n57336 ;
  assign n57338 = ~n57335 & ~n57337 ;
  assign n57339 = n9948 & n55888 ;
  assign n57340 = ~n57324 & ~n57339 ;
  assign n57341 = n57338 & n57340 ;
  assign n57342 = n55194 & ~n57341 ;
  assign n57343 = ~n57330 & ~n57342 ;
  assign n57344 = ~n57322 & ~n57343 ;
  assign n57345 = ~\pi1151  & n57325 ;
  assign n57346 = n9948 & n56297 ;
  assign n57347 = n9948 & n55844 ;
  assign n57348 = ~n55901 & n57347 ;
  assign n57349 = ~n57346 & ~n57348 ;
  assign n57350 = ~n53677 & ~n53702 ;
  assign n57351 = ~\pi1151  & n57350 ;
  assign n57352 = ~n57349 & n57351 ;
  assign n57353 = ~n57345 & ~n57352 ;
  assign n57354 = ~\pi0268  & ~\pi1151  ;
  assign n57355 = n52628 & ~n55874 ;
  assign n57356 = n53567 & n57355 ;
  assign n57357 = n9948 & n53567 ;
  assign n57358 = n55919 & n57357 ;
  assign n57359 = ~n57315 & n57358 ;
  assign n57360 = ~n57356 & ~n57359 ;
  assign n57361 = ~n57240 & n57241 ;
  assign n57362 = ~\pi0268  & ~n57361 ;
  assign n57363 = n57360 & n57362 ;
  assign n57364 = ~n57354 & ~n57363 ;
  assign n57365 = n57353 & ~n57364 ;
  assign n57366 = \pi1151  & n9948 ;
  assign n57367 = n55919 & n57366 ;
  assign n57368 = ~n57315 & n57367 ;
  assign n57369 = \pi1151  & ~n9948 ;
  assign n57370 = ~n55874 & n57369 ;
  assign n57371 = ~n56213 & n57370 ;
  assign n57372 = \pi0268  & ~n57371 ;
  assign n57373 = ~n57368 & n57372 ;
  assign n57374 = ~\pi1152  & ~n57373 ;
  assign n57375 = ~n55876 & n57276 ;
  assign n57376 = n53350 & n57375 ;
  assign n57377 = n53350 & ~n55926 ;
  assign n57378 = n57226 & n57377 ;
  assign n57379 = ~n57376 & ~n57378 ;
  assign n57380 = ~n57374 & n57379 ;
  assign n57381 = ~n57365 & ~n57380 ;
  assign n57382 = \pi1150  & ~n57381 ;
  assign n57383 = ~n57344 & n57382 ;
  assign n57384 = n57300 & ~n57383 ;
  assign n57385 = ~n57299 & n57384 ;
  assign n57386 = \pi1150  & ~n57174 ;
  assign n57387 = ~n57170 & n57386 ;
  assign n57388 = \pi1091  & ~n57387 ;
  assign n57389 = ~\pi0268  & ~\pi1091  ;
  assign n57390 = ~n57300 & ~n57389 ;
  assign n57391 = ~n57388 & n57390 ;
  assign n57392 = ~n57189 & n57390 ;
  assign n57393 = n57185 & n57392 ;
  assign n57394 = ~n57391 & ~n57393 ;
  assign n57395 = n57192 & n57394 ;
  assign n57396 = ~n57385 & n57395 ;
  assign n57397 = ~n57193 & ~n57396 ;
  assign n57398 = \pi1138  & n56042 ;
  assign n57399 = \pi0219  & ~n57398 ;
  assign n57400 = ~n20516 & n57399 ;
  assign n57401 = ~\pi0200  & \pi1091  ;
  assign n57402 = \pi1138  & n57401 ;
  assign n57403 = \pi0199  & ~n57402 ;
  assign n57404 = n20516 & n57403 ;
  assign n57405 = ~n57400 & ~n57404 ;
  assign n57406 = \pi0269  & ~n56698 ;
  assign n57407 = \pi0314  & ~\pi0817  ;
  assign n57408 = ~n53533 & n57407 ;
  assign n57409 = ~\pi1091  & ~n57408 ;
  assign n57410 = ~n57406 & n57409 ;
  assign n57411 = ~n57405 & ~n57410 ;
  assign n57412 = ~\pi0230  & n57411 ;
  assign n57413 = \pi0211  & \pi1137  ;
  assign n57414 = ~n56827 & ~n57413 ;
  assign n57415 = \pi1091  & ~n57414 ;
  assign n57416 = n54850 & ~n57415 ;
  assign n57417 = ~\pi0200  & n56819 ;
  assign n57418 = \pi1137  & n53865 ;
  assign n57419 = ~n57417 & ~n57418 ;
  assign n57420 = n57172 & n57419 ;
  assign n57421 = ~n57416 & ~n57420 ;
  assign n57422 = \pi0269  & ~\pi0314  ;
  assign n57423 = ~\pi0081  & \pi0269  ;
  assign n57424 = n53533 & n57423 ;
  assign n57425 = ~n57422 & ~n57424 ;
  assign n57426 = ~\pi1091  & ~n57407 ;
  assign n57427 = ~n56679 & ~n57426 ;
  assign n57428 = n57425 & ~n57427 ;
  assign n57429 = ~\pi0230  & ~n57428 ;
  assign n57430 = ~n57421 & n57429 ;
  assign n57431 = ~n57412 & ~n57430 ;
  assign n57432 = ~\pi0211  & \pi1138  ;
  assign n57433 = \pi0219  & n57432 ;
  assign n57434 = ~\pi0219  & ~n57414 ;
  assign n57435 = ~n57433 & ~n57434 ;
  assign n57436 = n56733 & n57435 ;
  assign n57437 = ~\pi0199  & \pi1137  ;
  assign n57438 = \pi0200  & ~n57437 ;
  assign n57439 = ~\pi0199  & \pi1136  ;
  assign n57440 = \pi0199  & \pi1138  ;
  assign n57441 = ~\pi0200  & ~n57440 ;
  assign n57442 = ~n57439 & n57441 ;
  assign n57443 = ~n57438 & ~n57442 ;
  assign n57444 = n53960 & ~n57443 ;
  assign n57445 = ~n57436 & ~n57444 ;
  assign n57446 = n57431 & n57445 ;
  assign n57447 = \pi1091  & n56728 ;
  assign n57448 = \pi0219  & ~n57447 ;
  assign n57449 = ~n20516 & n57448 ;
  assign n57450 = \pi0199  & ~n56693 ;
  assign n57451 = n20516 & n57450 ;
  assign n57452 = ~n57449 & ~n57451 ;
  assign n57453 = \pi0270  & ~n56698 ;
  assign n57454 = \pi0314  & ~\pi0805  ;
  assign n57455 = ~n53533 & n57454 ;
  assign n57456 = ~\pi1091  & ~n57455 ;
  assign n57457 = ~n57453 & n57456 ;
  assign n57458 = ~n57452 & ~n57457 ;
  assign n57459 = ~\pi0230  & n57458 ;
  assign n57460 = ~\pi0211  & \pi1139  ;
  assign n57461 = \pi0211  & \pi1140  ;
  assign n57462 = ~n57460 & ~n57461 ;
  assign n57463 = \pi1091  & ~n57462 ;
  assign n57464 = n54850 & ~n57463 ;
  assign n57465 = \pi1140  & n53865 ;
  assign n57466 = \pi1139  & n57401 ;
  assign n57467 = ~n57465 & ~n57466 ;
  assign n57468 = n57172 & n57467 ;
  assign n57469 = ~n57464 & ~n57468 ;
  assign n57470 = \pi0270  & ~\pi0314  ;
  assign n57471 = ~\pi0081  & \pi0270  ;
  assign n57472 = n53533 & n57471 ;
  assign n57473 = ~n57470 & ~n57472 ;
  assign n57474 = ~\pi1091  & ~n57454 ;
  assign n57475 = ~n56679 & ~n57474 ;
  assign n57476 = n57473 & ~n57475 ;
  assign n57477 = ~\pi0230  & ~n57476 ;
  assign n57478 = ~n57469 & n57477 ;
  assign n57479 = ~n57459 & ~n57478 ;
  assign n57480 = \pi0219  & n56728 ;
  assign n57481 = ~\pi0219  & ~n57462 ;
  assign n57482 = ~n57480 & ~n57481 ;
  assign n57483 = n56733 & n57482 ;
  assign n57484 = \pi1140  & n13645 ;
  assign n57485 = \pi0199  & \pi1141  ;
  assign n57486 = ~\pi0199  & \pi1139  ;
  assign n57487 = ~n57485 & ~n57486 ;
  assign n57488 = ~\pi0200  & ~n57487 ;
  assign n57489 = ~n57484 & ~n57488 ;
  assign n57490 = n53960 & n57489 ;
  assign n57491 = ~n57483 & ~n57490 ;
  assign n57492 = n57479 & n57491 ;
  assign n57493 = ~n53540 & n53541 ;
  assign n57494 = n53540 & n53548 ;
  assign n57495 = ~n57493 & ~n57494 ;
  assign n57496 = \pi1091  & n51665 ;
  assign n57497 = \pi1091  & \pi1146  ;
  assign n57498 = ~\pi0219  & ~n57497 ;
  assign n57499 = ~n57496 & n57498 ;
  assign n57500 = n57495 & n57499 ;
  assign n57501 = \pi0271  & \pi1091  ;
  assign n57502 = \pi0271  & \pi0276  ;
  assign n57503 = n53545 & n57502 ;
  assign n57504 = ~n57501 & ~n57503 ;
  assign n57505 = ~\pi0271  & ~n53937 ;
  assign n57506 = n57504 & ~n57505 ;
  assign n57507 = \pi0219  & ~n57506 ;
  assign n57508 = n12577 & n57497 ;
  assign n57509 = ~n57496 & n57508 ;
  assign n57510 = ~n57507 & ~n57509 ;
  assign n57511 = ~n57500 & n57510 ;
  assign n57512 = ~\pi0211  & \pi1147  ;
  assign n57513 = n55762 & n57512 ;
  assign n57514 = ~\pi0230  & ~n57513 ;
  assign n57515 = ~n20516 & n57514 ;
  assign n57516 = ~n57511 & n57515 ;
  assign n57517 = ~\pi0199  & ~n57497 ;
  assign n57518 = ~n53548 & n57517 ;
  assign n57519 = n53540 & n57518 ;
  assign n57520 = ~n53541 & n57517 ;
  assign n57521 = ~n53540 & n57520 ;
  assign n57522 = ~n57519 & ~n57521 ;
  assign n57523 = \pi0200  & ~n57522 ;
  assign n57524 = n50370 & ~n57506 ;
  assign n57525 = ~n57523 & ~n57524 ;
  assign n57526 = ~\pi0230  & n20515 ;
  assign n57527 = n6848 & n57526 ;
  assign n57528 = ~n57525 & n57527 ;
  assign n57529 = \pi0199  & ~n57506 ;
  assign n57530 = \pi1091  & \pi1145  ;
  assign n57531 = ~n53548 & ~n57530 ;
  assign n57532 = n53540 & n57531 ;
  assign n57533 = ~n53541 & ~n57530 ;
  assign n57534 = ~n53540 & n57533 ;
  assign n57535 = ~n57532 & ~n57534 ;
  assign n57536 = n12691 & ~n57535 ;
  assign n57537 = ~n57529 & ~n57536 ;
  assign n57538 = \pi1147  & n53846 ;
  assign n57539 = n57527 & ~n57538 ;
  assign n57540 = ~n57537 & n57539 ;
  assign n57541 = ~n57528 & ~n57540 ;
  assign n57542 = ~n57516 & n57541 ;
  assign n57543 = ~n51665 & n54456 ;
  assign n57544 = \pi0219  & ~n57512 ;
  assign n57545 = ~n9948 & ~n57544 ;
  assign n57546 = ~n57543 & n57545 ;
  assign n57547 = \pi0230  & ~n57546 ;
  assign n57548 = \pi1147  & n55690 ;
  assign n57549 = n13647 & n52535 ;
  assign n57550 = n12577 & n51630 ;
  assign n57551 = ~n57549 & ~n57550 ;
  assign n57552 = n44032 & n51721 ;
  assign n57553 = ~n52554 & ~n57552 ;
  assign n57554 = n57551 & n57553 ;
  assign n57555 = ~n57548 & n57554 ;
  assign n57556 = n55740 & ~n57555 ;
  assign n57557 = n57547 & ~n57556 ;
  assign n57558 = n57542 & ~n57557 ;
  assign n57559 = \pi1150  & ~n57341 ;
  assign n57560 = ~n57349 & n57350 ;
  assign n57561 = ~\pi1149  & ~n57325 ;
  assign n57562 = ~n57560 & n57561 ;
  assign n57563 = ~n54729 & ~n57562 ;
  assign n57564 = ~n57559 & ~n57563 ;
  assign n57565 = \pi1150  & ~n57326 ;
  assign n57566 = ~\pi0057  & \pi1150  ;
  assign n57567 = n6848 & n57566 ;
  assign n57568 = ~n57214 & n57567 ;
  assign n57569 = ~n57565 & ~n57568 ;
  assign n57570 = \pi1149  & ~n57361 ;
  assign n57571 = n57360 & n57570 ;
  assign n57572 = ~n54594 & ~n57571 ;
  assign n57573 = n57569 & ~n57572 ;
  assign n57574 = \pi1148  & ~n57573 ;
  assign n57575 = ~n57564 & n57574 ;
  assign n57576 = ~\pi1150  & n57241 ;
  assign n57577 = ~n57240 & n57576 ;
  assign n57578 = ~\pi1149  & ~\pi1150  ;
  assign n57579 = ~n57577 & n57578 ;
  assign n57580 = ~\pi1148  & ~n57579 ;
  assign n57581 = \pi0283  & ~n57580 ;
  assign n57582 = ~\pi1149  & ~n57220 ;
  assign n57583 = ~n57577 & n57582 ;
  assign n57584 = \pi0283  & n57583 ;
  assign n57585 = ~n57218 & n57584 ;
  assign n57586 = ~n57581 & ~n57585 ;
  assign n57587 = \pi1150  & ~n57196 ;
  assign n57588 = ~n57207 & n57587 ;
  assign n57589 = \pi1149  & ~n57588 ;
  assign n57590 = ~\pi1150  & ~n57231 ;
  assign n57591 = n57235 & n57590 ;
  assign n57592 = ~n57229 & n57591 ;
  assign n57593 = ~n57226 & n57592 ;
  assign n57594 = \pi0283  & ~n57593 ;
  assign n57595 = n57589 & n57594 ;
  assign n57596 = n57586 & ~n57595 ;
  assign n57597 = ~n57575 & ~n57596 ;
  assign n57598 = n54953 & ~n55693 ;
  assign n57599 = ~n52685 & ~n57598 ;
  assign n57600 = n53356 & n57180 ;
  assign n57601 = n54594 & ~n57188 ;
  assign n57602 = \pi1091  & ~n57601 ;
  assign n57603 = ~n57600 & n57602 ;
  assign n57604 = ~n57599 & n57603 ;
  assign n57605 = ~n9948 & n12577 ;
  assign n57606 = ~n15354 & ~n57605 ;
  assign n57607 = ~n57169 & ~n57606 ;
  assign n57608 = ~n20516 & n54680 ;
  assign n57609 = n44032 & n57566 ;
  assign n57610 = n6848 & n57609 ;
  assign n57611 = ~\pi1149  & ~n57610 ;
  assign n57612 = ~n57608 & n57611 ;
  assign n57613 = ~n57607 & n57612 ;
  assign n57614 = n20515 & ~n50370 ;
  assign n57615 = n6848 & n57614 ;
  assign n57616 = \pi1150  & n57615 ;
  assign n57617 = \pi1150  & ~n50713 ;
  assign n57618 = ~n20516 & n57617 ;
  assign n57619 = ~n57616 & ~n57618 ;
  assign n57620 = \pi1149  & ~n57172 ;
  assign n57621 = ~n54850 & n57620 ;
  assign n57622 = n57619 & n57621 ;
  assign n57623 = \pi1091  & \pi1148  ;
  assign n57624 = ~n57622 & n57623 ;
  assign n57625 = ~n57613 & n57624 ;
  assign n57626 = ~\pi0283  & ~n57625 ;
  assign n57627 = ~n57604 & n57626 ;
  assign n57628 = ~\pi0272  & ~n57627 ;
  assign n57629 = ~n57597 & n57628 ;
  assign n57630 = ~n57226 & ~n57229 ;
  assign n57631 = \pi1150  & ~n57305 ;
  assign n57632 = ~n57304 & n57631 ;
  assign n57633 = ~n57630 & n57632 ;
  assign n57634 = ~\pi1150  & n57375 ;
  assign n57635 = ~\pi1150  & ~n55926 ;
  assign n57636 = n57226 & n57635 ;
  assign n57637 = ~n57634 & ~n57636 ;
  assign n57638 = \pi1150  & ~n9948 ;
  assign n57639 = ~n56309 & n57638 ;
  assign n57640 = ~n55876 & n57639 ;
  assign n57641 = ~\pi1149  & ~n57640 ;
  assign n57642 = n57637 & n57641 ;
  assign n57643 = ~n57633 & n57642 ;
  assign n57644 = ~\pi1150  & n9948 ;
  assign n57645 = n55919 & n57644 ;
  assign n57646 = ~n57315 & n57645 ;
  assign n57647 = ~\pi1150  & ~n9948 ;
  assign n57648 = ~n55874 & n57647 ;
  assign n57649 = ~n56213 & n57648 ;
  assign n57650 = \pi1149  & ~n57649 ;
  assign n57651 = ~n57646 & n57650 ;
  assign n57652 = \pi1148  & ~n57651 ;
  assign n57653 = ~n57314 & n57318 ;
  assign n57654 = \pi1148  & \pi1150  ;
  assign n57655 = ~n57653 & n57654 ;
  assign n57656 = ~n57652 & ~n57655 ;
  assign n57657 = ~n57643 & ~n57656 ;
  assign n57658 = \pi0283  & \pi1148  ;
  assign n57659 = \pi1150  & n57271 ;
  assign n57660 = \pi1150  & n57269 ;
  assign n57661 = n57264 & n57660 ;
  assign n57662 = ~n57659 & ~n57661 ;
  assign n57663 = ~\pi1149  & ~n57291 ;
  assign n57664 = ~n57289 & n57663 ;
  assign n57665 = ~n54729 & ~n57664 ;
  assign n57666 = \pi0283  & ~n57665 ;
  assign n57667 = n57662 & n57666 ;
  assign n57668 = ~n57658 & ~n57667 ;
  assign n57669 = \pi1150  & ~n57267 ;
  assign n57670 = ~\pi1150  & n57282 ;
  assign n57671 = \pi0283  & \pi1149  ;
  assign n57672 = ~n57670 & n57671 ;
  assign n57673 = ~n57669 & n57672 ;
  assign n57674 = n57668 & ~n57673 ;
  assign n57675 = ~n57657 & ~n57674 ;
  assign n57676 = ~n20516 & n56168 ;
  assign n57677 = n53851 & n55740 ;
  assign n57678 = ~n57676 & ~n57677 ;
  assign n57679 = ~\pi1150  & ~n57678 ;
  assign n57680 = \pi1091  & \pi1150  ;
  assign n57681 = ~n57188 & n57680 ;
  assign n57682 = ~n57679 & ~n57681 ;
  assign n57683 = n52685 & ~n57682 ;
  assign n57684 = \pi0272  & ~n57683 ;
  assign n57685 = ~n54850 & ~n57172 ;
  assign n57686 = ~n53356 & n57168 ;
  assign n57687 = ~\pi0211  & ~n53356 ;
  assign n57688 = ~n20516 & n57687 ;
  assign n57689 = ~n57686 & ~n57688 ;
  assign n57690 = n57685 & n57689 ;
  assign n57691 = \pi1148  & ~n57690 ;
  assign n57692 = ~n57613 & n57691 ;
  assign n57693 = \pi1091  & ~n52685 ;
  assign n57694 = ~n57598 & n57693 ;
  assign n57695 = ~n57692 & n57694 ;
  assign n57696 = n57684 & ~n57695 ;
  assign n57697 = ~n53903 & ~n57696 ;
  assign n57698 = ~n57675 & ~n57697 ;
  assign n57699 = ~n57629 & ~n57698 ;
  assign n57700 = ~\pi0230  & n57699 ;
  assign n57701 = ~\pi1150  & ~n57180 ;
  assign n57702 = \pi1149  & n57619 ;
  assign n57703 = \pi1149  & ~n57188 ;
  assign n57704 = ~n57702 & ~n57703 ;
  assign n57705 = ~n57701 & ~n57704 ;
  assign n57706 = ~n57599 & ~n57705 ;
  assign n57707 = \pi1148  & ~n57622 ;
  assign n57708 = ~n57613 & n57707 ;
  assign n57709 = \pi0230  & ~n57708 ;
  assign n57710 = ~n57706 & n57709 ;
  assign n57711 = ~n57700 & ~n57710 ;
  assign n57712 = n53540 & n53541 ;
  assign n57713 = ~\pi0211  & n57497 ;
  assign n57714 = ~\pi0219  & \pi0273  ;
  assign n57715 = ~n57713 & n57714 ;
  assign n57716 = n57712 & n57715 ;
  assign n57717 = ~\pi0219  & ~n57713 ;
  assign n57718 = n53551 & n57717 ;
  assign n57719 = ~\pi0219  & ~\pi0273  ;
  assign n57720 = ~n57713 & n57719 ;
  assign n57721 = ~n57712 & n57720 ;
  assign n57722 = ~n57718 & ~n57721 ;
  assign n57723 = ~n57716 & n57722 ;
  assign n57724 = ~\pi0273  & ~n53934 ;
  assign n57725 = ~n53551 & ~n57724 ;
  assign n57726 = \pi0219  & ~n57725 ;
  assign n57727 = ~n9948 & ~n57726 ;
  assign n57728 = n57723 & n57727 ;
  assign n57729 = \pi0299  & ~n57726 ;
  assign n57730 = n57723 & n57729 ;
  assign n57731 = ~\pi0200  & n57497 ;
  assign n57732 = ~\pi0199  & ~n57731 ;
  assign n57733 = ~\pi0273  & n57732 ;
  assign n57734 = ~n57712 & n57733 ;
  assign n57735 = ~\pi0199  & \pi0273  ;
  assign n57736 = ~n57731 & n57735 ;
  assign n57737 = n57712 & n57736 ;
  assign n57738 = ~n57734 & ~n57737 ;
  assign n57739 = n53551 & n57732 ;
  assign n57740 = \pi0199  & \pi0273  ;
  assign n57741 = n53549 & n57740 ;
  assign n57742 = ~n53546 & n57741 ;
  assign n57743 = \pi0199  & ~\pi0273  ;
  assign n57744 = ~n53934 & n57743 ;
  assign n57745 = ~\pi0299  & ~n57744 ;
  assign n57746 = ~n57742 & n57745 ;
  assign n57747 = ~n57739 & n57746 ;
  assign n57748 = n57738 & n57747 ;
  assign n57749 = ~n57730 & ~n57748 ;
  assign n57750 = n52558 & ~n57749 ;
  assign n57751 = ~\pi1148  & ~n57750 ;
  assign n57752 = n53847 & n57525 ;
  assign n57753 = ~n57748 & ~n57752 ;
  assign n57754 = ~\pi0211  & n55762 ;
  assign n57755 = ~n55740 & n57754 ;
  assign n57756 = \pi1148  & ~n57755 ;
  assign n57757 = n53974 & n56042 ;
  assign n57758 = n57756 & ~n57757 ;
  assign n57759 = ~n57730 & n57758 ;
  assign n57760 = n57753 & n57759 ;
  assign n57761 = \pi1148  & ~n55740 ;
  assign n57762 = ~n57755 & n57761 ;
  assign n57763 = ~n57760 & ~n57762 ;
  assign n57764 = ~n57751 & n57763 ;
  assign n57765 = ~n57728 & ~n57764 ;
  assign n57766 = ~\pi0230  & ~n57765 ;
  assign n57767 = \pi1091  & n13648 ;
  assign n57768 = \pi1091  & ~n56096 ;
  assign n57769 = n53770 & n57768 ;
  assign n57770 = ~n57767 & ~n57769 ;
  assign n57771 = \pi1091  & n57276 ;
  assign n57772 = ~n55993 & n57771 ;
  assign n57773 = n57749 & ~n57772 ;
  assign n57774 = n57770 & n57773 ;
  assign n57775 = ~n9948 & ~n57772 ;
  assign n57776 = ~\pi0230  & \pi1147  ;
  assign n57777 = ~n57775 & n57776 ;
  assign n57778 = ~n57774 & n57777 ;
  assign n57779 = ~\pi0219  & ~n53444 ;
  assign n57780 = ~n20516 & n57779 ;
  assign n57781 = ~\pi1146  & n12691 ;
  assign n57782 = n57172 & ~n57781 ;
  assign n57783 = ~n57780 & ~n57782 ;
  assign n57784 = \pi1147  & ~n57783 ;
  assign n57785 = \pi1146  & ~n54322 ;
  assign n57786 = ~n57606 & n57785 ;
  assign n57787 = ~\pi1148  & ~n57786 ;
  assign n57788 = ~n57784 & n57787 ;
  assign n57789 = ~\pi1146  & n12577 ;
  assign n57790 = \pi0211  & ~\pi1147  ;
  assign n57791 = ~n50713 & ~n57790 ;
  assign n57792 = ~n57789 & n57791 ;
  assign n57793 = ~n20516 & n57792 ;
  assign n57794 = ~\pi0199  & \pi1147  ;
  assign n57795 = \pi0200  & ~n57794 ;
  assign n57796 = ~n57781 & ~n57795 ;
  assign n57797 = n20516 & n57796 ;
  assign n57798 = ~n57793 & ~n57797 ;
  assign n57799 = \pi1148  & n57798 ;
  assign n57800 = \pi0230  & ~n57799 ;
  assign n57801 = ~n57788 & n57800 ;
  assign n57802 = ~n57778 & ~n57801 ;
  assign n57803 = ~n57766 & n57802 ;
  assign n57804 = \pi0314  & ~\pi0659  ;
  assign n57805 = ~\pi1091  & ~n57804 ;
  assign n57806 = ~n56679 & ~n57805 ;
  assign n57807 = ~\pi0081  & \pi0274  ;
  assign n57808 = n53533 & n57807 ;
  assign n57809 = \pi0274  & ~\pi0314  ;
  assign n57810 = ~\pi0211  & ~n57809 ;
  assign n57811 = ~n57808 & n57810 ;
  assign n57812 = ~n57806 & n57811 ;
  assign n57813 = \pi0211  & ~n57809 ;
  assign n57814 = ~n57808 & n57813 ;
  assign n57815 = ~n57806 & n57814 ;
  assign n57816 = ~\pi0211  & n56703 ;
  assign n57817 = \pi0211  & n56763 ;
  assign n57818 = ~\pi0219  & ~n57817 ;
  assign n57819 = ~n57816 & n57818 ;
  assign n57820 = ~n57815 & n57819 ;
  assign n57821 = ~n57812 & n57820 ;
  assign n57822 = \pi0274  & ~n56698 ;
  assign n57823 = ~n53533 & n57804 ;
  assign n57824 = ~\pi1091  & ~n57823 ;
  assign n57825 = ~n57822 & n57824 ;
  assign n57826 = \pi0219  & ~n57496 ;
  assign n57827 = ~n57825 & n57826 ;
  assign n57828 = ~n20516 & ~n57827 ;
  assign n57829 = ~n57821 & n57828 ;
  assign n57830 = ~\pi0230  & ~n20516 ;
  assign n57831 = ~\pi0200  & n57530 ;
  assign n57832 = \pi0199  & ~n57831 ;
  assign n57833 = ~\pi0230  & n57832 ;
  assign n57834 = ~n57825 & n57833 ;
  assign n57835 = ~n57830 & ~n57834 ;
  assign n57836 = ~\pi0230  & ~n56704 ;
  assign n57837 = \pi0200  & n56763 ;
  assign n57838 = ~\pi0199  & ~n57837 ;
  assign n57839 = n57806 & n57838 ;
  assign n57840 = ~n57808 & ~n57809 ;
  assign n57841 = n57838 & ~n57840 ;
  assign n57842 = ~n57839 & ~n57841 ;
  assign n57843 = n57836 & ~n57842 ;
  assign n57844 = n57835 & ~n57843 ;
  assign n57845 = ~n57829 & ~n57844 ;
  assign n57846 = ~n50701 & ~n52920 ;
  assign n57847 = ~\pi0219  & ~n50661 ;
  assign n57848 = ~n51666 & n57847 ;
  assign n57849 = ~n57846 & ~n57848 ;
  assign n57850 = ~\pi0299  & ~n51723 ;
  assign n57851 = ~n50637 & n52517 ;
  assign n57852 = n57850 & ~n57851 ;
  assign n57853 = ~n57849 & ~n57852 ;
  assign n57854 = n9948 & ~n57853 ;
  assign n57855 = ~n9948 & ~n52824 ;
  assign n57856 = ~n57848 & n57855 ;
  assign n57857 = \pi0230  & ~n57856 ;
  assign n57858 = ~n57854 & n57857 ;
  assign n57859 = ~n57845 & ~n57858 ;
  assign n57860 = n53189 & n57188 ;
  assign n57861 = \pi1150  & ~\pi1151  ;
  assign n57862 = ~n57180 & n57861 ;
  assign n57863 = ~n57860 & ~n57862 ;
  assign n57864 = n53397 & ~n55693 ;
  assign n57865 = ~\pi1149  & ~n57864 ;
  assign n57866 = n57863 & n57865 ;
  assign n57867 = \pi1151  & n57168 ;
  assign n57868 = ~\pi0211  & \pi1151  ;
  assign n57869 = ~n20516 & n57868 ;
  assign n57870 = ~n57867 & ~n57869 ;
  assign n57871 = n57621 & n57870 ;
  assign n57872 = n53356 & ~n57168 ;
  assign n57873 = ~n57166 & n57872 ;
  assign n57874 = ~n57871 & ~n57873 ;
  assign n57875 = \pi0230  & n57874 ;
  assign n57876 = ~n57866 & n57875 ;
  assign n57877 = ~n57323 & ~n57327 ;
  assign n57878 = ~\pi0275  & \pi1151  ;
  assign n57879 = ~\pi0275  & ~n57361 ;
  assign n57880 = n57360 & n57879 ;
  assign n57881 = ~n57878 & ~n57880 ;
  assign n57882 = n57877 & ~n57881 ;
  assign n57883 = n55568 & n55919 ;
  assign n57884 = ~n57315 & n57883 ;
  assign n57885 = n53120 & ~n55874 ;
  assign n57886 = ~n56213 & n57885 ;
  assign n57887 = \pi0275  & ~n57886 ;
  assign n57888 = ~n57884 & n57887 ;
  assign n57889 = ~\pi1151  & n57888 ;
  assign n57890 = n57318 & n57888 ;
  assign n57891 = ~n57314 & n57890 ;
  assign n57892 = ~n57889 & ~n57891 ;
  assign n57893 = \pi1150  & n57892 ;
  assign n57894 = ~n57882 & n57893 ;
  assign n57895 = \pi1151  & ~n57305 ;
  assign n57896 = ~n57304 & n57895 ;
  assign n57897 = ~n57630 & n57896 ;
  assign n57898 = ~\pi1151  & n57375 ;
  assign n57899 = ~\pi1151  & ~n55926 ;
  assign n57900 = n57226 & n57899 ;
  assign n57901 = ~n57898 & ~n57900 ;
  assign n57902 = ~n56309 & n57369 ;
  assign n57903 = ~n55876 & n57902 ;
  assign n57904 = \pi0275  & ~n57903 ;
  assign n57905 = n57901 & n57904 ;
  assign n57906 = ~n57897 & n57905 ;
  assign n57907 = ~\pi0275  & ~n57325 ;
  assign n57908 = ~n57560 & n57907 ;
  assign n57909 = ~\pi1150  & ~n57878 ;
  assign n57910 = ~n57908 & n57909 ;
  assign n57911 = n53397 & ~n57341 ;
  assign n57912 = ~n57910 & ~n57911 ;
  assign n57913 = ~n57906 & ~n57912 ;
  assign n57914 = ~n57894 & ~n57913 ;
  assign n57915 = \pi1149  & ~n57914 ;
  assign n57916 = ~n57229 & n57236 ;
  assign n57917 = ~n57226 & n57916 ;
  assign n57918 = ~\pi1151  & ~n57917 ;
  assign n57919 = ~n57588 & ~n57861 ;
  assign n57920 = ~n57918 & ~n57919 ;
  assign n57921 = \pi1151  & ~n57220 ;
  assign n57922 = ~n57218 & n57921 ;
  assign n57923 = ~n53397 & ~n57577 ;
  assign n57924 = ~n57922 & ~n57923 ;
  assign n57925 = ~n57920 & ~n57924 ;
  assign n57926 = ~\pi0275  & n57925 ;
  assign n57927 = ~\pi0275  & ~\pi1149  ;
  assign n57928 = \pi1151  & ~n57271 ;
  assign n57929 = ~n57270 & n57928 ;
  assign n57930 = ~\pi1150  & ~n57293 ;
  assign n57931 = ~\pi1149  & n57930 ;
  assign n57932 = ~n57929 & n57931 ;
  assign n57933 = ~n57927 & ~n57932 ;
  assign n57934 = ~\pi1151  & ~n57282 ;
  assign n57935 = n54729 & ~n57934 ;
  assign n57936 = ~n57268 & n57935 ;
  assign n57937 = n57933 & ~n57936 ;
  assign n57938 = ~n57926 & ~n57937 ;
  assign n57939 = n53903 & ~n57938 ;
  assign n57940 = ~n57915 & n57939 ;
  assign n57941 = ~n57866 & n57874 ;
  assign n57942 = \pi0230  & ~n57941 ;
  assign n57943 = \pi1149  & n57870 ;
  assign n57944 = ~n57607 & n57943 ;
  assign n57945 = ~n53356 & ~n57864 ;
  assign n57946 = ~n57944 & ~n57945 ;
  assign n57947 = ~\pi1149  & \pi1151  ;
  assign n57948 = ~n57188 & n57947 ;
  assign n57949 = ~n57871 & ~n57948 ;
  assign n57950 = \pi1150  & n57949 ;
  assign n57951 = \pi1091  & ~n57950 ;
  assign n57952 = ~n57946 & n57951 ;
  assign n57953 = ~\pi1151  & n54729 ;
  assign n57954 = ~n57678 & n57953 ;
  assign n57955 = \pi0275  & ~n57954 ;
  assign n57956 = ~n57952 & n57955 ;
  assign n57957 = ~\pi0275  & \pi1091  ;
  assign n57958 = n57874 & n57957 ;
  assign n57959 = ~n57866 & n57958 ;
  assign n57960 = ~n53903 & ~n57959 ;
  assign n57961 = ~n57956 & n57960 ;
  assign n57962 = ~n57942 & ~n57961 ;
  assign n57963 = ~n57940 & n57962 ;
  assign n57964 = ~n57876 & ~n57963 ;
  assign n57965 = \pi0219  & ~n57713 ;
  assign n57966 = ~n20516 & n57965 ;
  assign n57967 = \pi0199  & ~n57731 ;
  assign n57968 = n20516 & n57967 ;
  assign n57969 = ~n57966 & ~n57968 ;
  assign n57970 = n53545 & n53547 ;
  assign n57971 = n53536 & ~n53545 ;
  assign n57972 = ~n57970 & ~n57971 ;
  assign n57973 = ~n57969 & n57972 ;
  assign n57974 = ~\pi1091  & ~n53540 ;
  assign n57975 = ~\pi0276  & ~n53535 ;
  assign n57976 = ~\pi0081  & ~\pi0276  ;
  assign n57977 = n53533 & n57976 ;
  assign n57978 = ~n57975 & ~n57977 ;
  assign n57979 = ~\pi0230  & n57978 ;
  assign n57980 = n57974 & n57979 ;
  assign n57981 = ~n50658 & ~n52817 ;
  assign n57982 = \pi1091  & ~n57981 ;
  assign n57983 = n54850 & ~n57982 ;
  assign n57984 = \pi1145  & n53865 ;
  assign n57985 = ~n56764 & ~n57984 ;
  assign n57986 = n57172 & n57985 ;
  assign n57987 = ~\pi0230  & ~n57986 ;
  assign n57988 = ~n57983 & n57987 ;
  assign n57989 = ~n57980 & ~n57988 ;
  assign n57990 = ~n57973 & ~n57989 ;
  assign n57991 = ~\pi0219  & ~n57981 ;
  assign n57992 = \pi0219  & n52816 ;
  assign n57993 = ~n20516 & ~n57992 ;
  assign n57994 = ~n57991 & n57993 ;
  assign n57995 = ~n50644 & n54137 ;
  assign n57996 = \pi0230  & ~n52519 ;
  assign n57997 = ~n57995 & n57996 ;
  assign n57998 = ~n56733 & ~n57997 ;
  assign n57999 = ~n57994 & ~n57998 ;
  assign n58000 = ~n57990 & ~n57999 ;
  assign n58001 = \pi0314  & ~\pi0820  ;
  assign n58002 = ~\pi1091  & ~n58001 ;
  assign n58003 = ~n56679 & ~n58002 ;
  assign n58004 = ~\pi0081  & \pi0277  ;
  assign n58005 = n53533 & n58004 ;
  assign n58006 = \pi0277  & ~\pi0314  ;
  assign n58007 = \pi0211  & ~n58006 ;
  assign n58008 = ~n58005 & n58007 ;
  assign n58009 = ~n58003 & n58008 ;
  assign n58010 = ~\pi0211  & ~n58006 ;
  assign n58011 = ~n58005 & n58010 ;
  assign n58012 = ~n58003 & n58011 ;
  assign n58013 = \pi0211  & n56692 ;
  assign n58014 = \pi1091  & \pi1140  ;
  assign n58015 = ~\pi0211  & n58014 ;
  assign n58016 = ~\pi0219  & ~n58015 ;
  assign n58017 = ~n58013 & n58016 ;
  assign n58018 = ~n58012 & n58017 ;
  assign n58019 = ~n58009 & n58018 ;
  assign n58020 = \pi0277  & ~n56698 ;
  assign n58021 = ~n53533 & n58001 ;
  assign n58022 = ~\pi1091  & ~n58021 ;
  assign n58023 = ~n58020 & n58022 ;
  assign n58024 = ~n50669 & ~n56721 ;
  assign n58025 = ~n58023 & ~n58024 ;
  assign n58026 = ~n20516 & ~n58025 ;
  assign n58027 = ~n58019 & n58026 ;
  assign n58028 = \pi0200  & ~n58006 ;
  assign n58029 = ~n58005 & n58028 ;
  assign n58030 = ~n58003 & n58029 ;
  assign n58031 = ~\pi0200  & ~n58006 ;
  assign n58032 = ~n58005 & n58031 ;
  assign n58033 = ~n58003 & n58032 ;
  assign n58034 = \pi0200  & n56692 ;
  assign n58035 = ~\pi0200  & n58014 ;
  assign n58036 = ~\pi0199  & ~n58035 ;
  assign n58037 = ~n58034 & n58036 ;
  assign n58038 = ~n58033 & n58037 ;
  assign n58039 = ~n58030 & n58038 ;
  assign n58040 = \pi0199  & ~n56754 ;
  assign n58041 = ~n58023 & n58040 ;
  assign n58042 = n20516 & ~n58041 ;
  assign n58043 = ~n58039 & n58042 ;
  assign n58044 = ~n58027 & ~n58043 ;
  assign n58045 = ~\pi0230  & ~n58044 ;
  assign n58046 = ~\pi0199  & \pi1140  ;
  assign n58047 = n50636 & ~n58046 ;
  assign n58048 = \pi0200  & ~n56734 ;
  assign n58049 = ~n58047 & ~n58048 ;
  assign n58050 = n20516 & ~n58049 ;
  assign n58051 = ~\pi0211  & \pi1140  ;
  assign n58052 = \pi0211  & \pi1141  ;
  assign n58053 = ~\pi0219  & ~n58052 ;
  assign n58054 = ~n58051 & n58053 ;
  assign n58055 = \pi0230  & ~n50669 ;
  assign n58056 = ~n58054 & n58055 ;
  assign n58057 = ~n53960 & ~n58056 ;
  assign n58058 = ~n58050 & ~n58057 ;
  assign n58059 = ~n58045 & ~n58058 ;
  assign n58060 = \pi0314  & \pi0976  ;
  assign n58061 = ~\pi1091  & ~n58060 ;
  assign n58062 = ~n56679 & ~n58061 ;
  assign n58063 = ~\pi0081  & \pi0278  ;
  assign n58064 = n53533 & n58063 ;
  assign n58065 = \pi0278  & ~\pi0314  ;
  assign n58066 = ~\pi0199  & ~n58065 ;
  assign n58067 = ~n58064 & n58066 ;
  assign n58068 = ~n58062 & n58067 ;
  assign n58069 = \pi1091  & ~\pi1133  ;
  assign n58070 = ~\pi0199  & n58069 ;
  assign n58071 = ~n58068 & ~n58070 ;
  assign n58072 = \pi0278  & ~\pi1091  ;
  assign n58073 = ~n56811 & ~n58072 ;
  assign n58074 = \pi0314  & ~\pi0976  ;
  assign n58075 = ~n53533 & n58074 ;
  assign n58076 = ~\pi0299  & ~n58075 ;
  assign n58077 = ~n58073 & n58076 ;
  assign n58078 = ~n43637 & ~n58077 ;
  assign n58079 = n58071 & ~n58078 ;
  assign n58080 = ~n44032 & ~n58079 ;
  assign n58081 = \pi1091  & ~\pi1132  ;
  assign n58082 = ~\pi0199  & n58081 ;
  assign n58083 = ~\pi0199  & ~n58082 ;
  assign n58084 = ~n58075 & ~n58082 ;
  assign n58085 = ~n58073 & n58084 ;
  assign n58086 = ~n58083 & ~n58085 ;
  assign n58087 = ~n58068 & ~n58086 ;
  assign n58088 = ~\pi0200  & ~n53846 ;
  assign n58089 = ~n58087 & n58088 ;
  assign n58090 = ~n58080 & ~n58089 ;
  assign n58091 = ~n58073 & ~n58075 ;
  assign n58092 = \pi0219  & ~n58091 ;
  assign n58093 = ~\pi0219  & ~n58065 ;
  assign n58094 = ~n58064 & n58093 ;
  assign n58095 = ~n58062 & n58094 ;
  assign n58096 = \pi0211  & ~\pi1133  ;
  assign n58097 = ~\pi0211  & ~\pi1132  ;
  assign n58098 = ~n58096 & ~n58097 ;
  assign n58099 = n53909 & ~n58098 ;
  assign n58100 = \pi0299  & ~n58099 ;
  assign n58101 = ~n58095 & n58100 ;
  assign n58102 = ~n58092 & n58101 ;
  assign n58103 = ~n9948 & ~n58099 ;
  assign n58104 = ~n58095 & n58103 ;
  assign n58105 = ~n58092 & n58104 ;
  assign n58106 = ~\pi0230  & ~n57757 ;
  assign n58107 = ~n57755 & n58106 ;
  assign n58108 = ~n58105 & n58107 ;
  assign n58109 = ~n58102 & n58108 ;
  assign n58110 = ~n58090 & n58109 ;
  assign n58111 = ~\pi0199  & \pi1133  ;
  assign n58112 = \pi0200  & ~n58111 ;
  assign n58113 = ~\pi0299  & ~n58112 ;
  assign n58114 = ~\pi1132  & n55608 ;
  assign n58115 = n58113 & ~n58114 ;
  assign n58116 = n50701 & n58098 ;
  assign n58117 = ~n56237 & ~n58116 ;
  assign n58118 = ~n58115 & n58117 ;
  assign n58119 = n9948 & ~n58118 ;
  assign n58120 = ~n9948 & ~n50713 ;
  assign n58121 = ~\pi0219  & ~n58098 ;
  assign n58122 = n58120 & ~n58121 ;
  assign n58123 = \pi0230  & ~n58122 ;
  assign n58124 = ~n58119 & n58123 ;
  assign n58125 = ~\pi0230  & ~n9948 ;
  assign n58126 = ~n57755 & n58125 ;
  assign n58127 = ~n58105 & n58126 ;
  assign n58128 = ~n58124 & ~n58127 ;
  assign n58129 = ~n58110 & n58128 ;
  assign n58130 = \pi1134  & n58129 ;
  assign n58131 = ~\pi0230  & ~n58105 ;
  assign n58132 = ~n9948 & n58131 ;
  assign n58133 = ~\pi0200  & ~n58087 ;
  assign n58134 = ~n58080 & ~n58133 ;
  assign n58135 = ~n58102 & n58131 ;
  assign n58136 = ~n58134 & n58135 ;
  assign n58137 = ~n58132 & ~n58136 ;
  assign n58138 = n44035 & n58111 ;
  assign n58139 = ~\pi0199  & \pi1132  ;
  assign n58140 = n44032 & n58139 ;
  assign n58141 = ~n58138 & ~n58140 ;
  assign n58142 = ~n58116 & n58141 ;
  assign n58143 = n9948 & ~n58142 ;
  assign n58144 = ~\pi0219  & n58098 ;
  assign n58145 = ~n9948 & n58144 ;
  assign n58146 = \pi0230  & ~n58145 ;
  assign n58147 = ~n58143 & n58146 ;
  assign n58148 = ~\pi1134  & ~n58147 ;
  assign n58149 = n58137 & n58148 ;
  assign n58150 = ~n58130 & ~n58149 ;
  assign n58151 = \pi1135  & n50689 ;
  assign n58152 = \pi1133  & n12577 ;
  assign n58153 = ~n58151 & ~n58152 ;
  assign n58154 = ~n55740 & ~n58153 ;
  assign n58155 = \pi0230  & ~n58154 ;
  assign n58156 = \pi0199  & \pi1135  ;
  assign n58157 = ~n58111 & ~n58156 ;
  assign n58158 = n44032 & ~n58157 ;
  assign n58159 = \pi0299  & ~n58153 ;
  assign n58160 = ~n58158 & ~n58159 ;
  assign n58161 = n55740 & ~n58160 ;
  assign n58162 = n58155 & ~n58161 ;
  assign n58163 = ~\pi1134  & n58162 ;
  assign n58164 = \pi0279  & ~\pi0314  ;
  assign n58165 = ~\pi0081  & \pi0279  ;
  assign n58166 = n53533 & n58165 ;
  assign n58167 = ~n58164 & ~n58166 ;
  assign n58168 = \pi0314  & \pi0958  ;
  assign n58169 = ~\pi1091  & ~n58168 ;
  assign n58170 = ~n56679 & ~n58169 ;
  assign n58171 = n58167 & ~n58170 ;
  assign n58172 = ~n55744 & ~n58069 ;
  assign n58173 = ~n58171 & n58172 ;
  assign n58174 = ~\pi0219  & ~n58173 ;
  assign n58175 = \pi0279  & ~\pi1091  ;
  assign n58176 = ~n56811 & ~n58175 ;
  assign n58177 = \pi0314  & ~\pi0958  ;
  assign n58178 = ~n53533 & n58177 ;
  assign n58179 = ~n58176 & ~n58178 ;
  assign n58180 = \pi1135  & n56042 ;
  assign n58181 = \pi0219  & ~n58180 ;
  assign n58182 = ~n58179 & n58181 ;
  assign n58183 = ~n20516 & ~n58182 ;
  assign n58184 = ~n58174 & n58183 ;
  assign n58185 = ~\pi0230  & ~n58184 ;
  assign n58186 = ~\pi1133  & n57401 ;
  assign n58187 = ~\pi0199  & ~n58186 ;
  assign n58188 = n20516 & n58187 ;
  assign n58189 = ~n58171 & n58188 ;
  assign n58190 = ~n53865 & n58189 ;
  assign n58191 = n50383 & n56805 ;
  assign n58192 = \pi0199  & ~n58178 ;
  assign n58193 = ~n58176 & n58192 ;
  assign n58194 = ~n58191 & ~n58193 ;
  assign n58195 = n20516 & ~n53865 ;
  assign n58196 = ~n58194 & n58195 ;
  assign n58197 = ~n58190 & ~n58196 ;
  assign n58198 = ~\pi1134  & n58197 ;
  assign n58199 = n58185 & n58198 ;
  assign n58200 = ~n58163 & ~n58199 ;
  assign n58201 = ~\pi1133  & n12691 ;
  assign n58202 = ~\pi0200  & \pi1135  ;
  assign n58203 = \pi0199  & ~n58202 ;
  assign n58204 = ~n58201 & ~n58203 ;
  assign n58205 = n20516 & ~n58204 ;
  assign n58206 = ~\pi0211  & ~\pi1133  ;
  assign n58207 = ~\pi0219  & ~n58206 ;
  assign n58208 = ~n58151 & ~n58207 ;
  assign n58209 = ~n20516 & n58208 ;
  assign n58210 = ~n58205 & ~n58209 ;
  assign n58211 = \pi0230  & ~n58210 ;
  assign n58212 = \pi1134  & n58211 ;
  assign n58213 = n53909 & ~n58206 ;
  assign n58214 = ~n20516 & n58213 ;
  assign n58215 = ~\pi0230  & ~n58214 ;
  assign n58216 = ~n58184 & n58215 ;
  assign n58217 = n20516 & ~n58194 ;
  assign n58218 = ~n58189 & ~n58217 ;
  assign n58219 = \pi1134  & n58218 ;
  assign n58220 = n58216 & n58219 ;
  assign n58221 = ~n58212 & ~n58220 ;
  assign n58222 = n58200 & n58221 ;
  assign n58223 = \pi0280  & ~n56698 ;
  assign n58224 = \pi0314  & ~\pi0914  ;
  assign n58225 = ~n53533 & n58224 ;
  assign n58226 = ~\pi1091  & ~n58225 ;
  assign n58227 = ~n58223 & n58226 ;
  assign n58228 = ~\pi0211  & \pi1137  ;
  assign n58229 = \pi0219  & ~n58228 ;
  assign n58230 = ~n56721 & ~n58229 ;
  assign n58231 = ~n58227 & ~n58230 ;
  assign n58232 = ~\pi0211  & \pi1135  ;
  assign n58233 = \pi0211  & \pi1136  ;
  assign n58234 = ~n58232 & ~n58233 ;
  assign n58235 = n53909 & n58234 ;
  assign n58236 = \pi0314  & \pi0914  ;
  assign n58237 = ~n53534 & n58236 ;
  assign n58238 = ~\pi0081  & ~\pi0280  ;
  assign n58239 = n53533 & n58238 ;
  assign n58240 = ~\pi0280  & ~\pi0314  ;
  assign n58241 = ~\pi1091  & ~n58240 ;
  assign n58242 = ~n58239 & n58241 ;
  assign n58243 = ~n58237 & n58242 ;
  assign n58244 = ~\pi0219  & n58243 ;
  assign n58245 = ~n58235 & ~n58244 ;
  assign n58246 = ~n58231 & n58245 ;
  assign n58247 = n57830 & ~n58246 ;
  assign n58248 = ~\pi0199  & n20515 ;
  assign n58249 = n6848 & n58248 ;
  assign n58250 = \pi1137  & n57401 ;
  assign n58251 = n20516 & ~n58250 ;
  assign n58252 = ~n58227 & n58251 ;
  assign n58253 = ~n58249 & ~n58252 ;
  assign n58254 = \pi0200  & \pi1136  ;
  assign n58255 = \pi1091  & ~n58202 ;
  assign n58256 = ~n58254 & n58255 ;
  assign n58257 = ~\pi0199  & ~n58256 ;
  assign n58258 = ~n58243 & n58257 ;
  assign n58259 = ~\pi0230  & ~n58258 ;
  assign n58260 = ~n58253 & n58259 ;
  assign n58261 = \pi0200  & ~n57439 ;
  assign n58262 = \pi0199  & \pi1137  ;
  assign n58263 = ~\pi0200  & ~n56836 ;
  assign n58264 = ~n58262 & n58263 ;
  assign n58265 = ~n58261 & ~n58264 ;
  assign n58266 = n53960 & ~n58265 ;
  assign n58267 = ~\pi0219  & n58234 ;
  assign n58268 = ~n58229 & ~n58267 ;
  assign n58269 = n56733 & ~n58268 ;
  assign n58270 = ~n58266 & ~n58269 ;
  assign n58271 = ~n58260 & n58270 ;
  assign n58272 = ~n58247 & n58271 ;
  assign n58273 = \pi0211  & \pi1138  ;
  assign n58274 = ~n58228 & ~n58273 ;
  assign n58275 = \pi1091  & ~n58274 ;
  assign n58276 = n54850 & ~n58275 ;
  assign n58277 = \pi1138  & n53865 ;
  assign n58278 = ~n58250 & ~n58277 ;
  assign n58279 = n57172 & n58278 ;
  assign n58280 = ~n58276 & ~n58279 ;
  assign n58281 = \pi0281  & ~\pi0314  ;
  assign n58282 = ~\pi0081  & \pi0281  ;
  assign n58283 = n53533 & n58282 ;
  assign n58284 = ~n58281 & ~n58283 ;
  assign n58285 = \pi0314  & ~\pi0830  ;
  assign n58286 = ~\pi1091  & ~n58285 ;
  assign n58287 = ~n56679 & ~n58286 ;
  assign n58288 = n58284 & ~n58287 ;
  assign n58289 = ~\pi0230  & ~n58288 ;
  assign n58290 = ~n58280 & n58289 ;
  assign n58291 = \pi1139  & n56042 ;
  assign n58292 = \pi0219  & ~n58291 ;
  assign n58293 = ~n20516 & n58292 ;
  assign n58294 = \pi0199  & ~n57466 ;
  assign n58295 = n20516 & n58294 ;
  assign n58296 = ~n58293 & ~n58295 ;
  assign n58297 = \pi0281  & ~n56698 ;
  assign n58298 = ~n53533 & n58285 ;
  assign n58299 = ~\pi1091  & ~n58298 ;
  assign n58300 = ~n58297 & n58299 ;
  assign n58301 = ~\pi0230  & ~n58300 ;
  assign n58302 = ~n58296 & n58301 ;
  assign n58303 = \pi0219  & n57460 ;
  assign n58304 = ~\pi0219  & ~n58274 ;
  assign n58305 = ~n58303 & ~n58304 ;
  assign n58306 = n56733 & n58305 ;
  assign n58307 = ~\pi0199  & \pi1138  ;
  assign n58308 = \pi0200  & ~n58307 ;
  assign n58309 = \pi0199  & \pi1139  ;
  assign n58310 = ~\pi0200  & ~n57437 ;
  assign n58311 = ~n58309 & n58310 ;
  assign n58312 = ~n58308 & ~n58311 ;
  assign n58313 = n53960 & ~n58312 ;
  assign n58314 = ~n58306 & ~n58313 ;
  assign n58315 = ~n58302 & n58314 ;
  assign n58316 = ~n58290 & n58315 ;
  assign n58317 = \pi1140  & n56042 ;
  assign n58318 = \pi0219  & ~n58317 ;
  assign n58319 = ~n20516 & n58318 ;
  assign n58320 = \pi0199  & ~n58035 ;
  assign n58321 = n20516 & n58320 ;
  assign n58322 = ~n58319 & ~n58321 ;
  assign n58323 = \pi0282  & ~n56698 ;
  assign n58324 = \pi0314  & ~\pi0836  ;
  assign n58325 = ~n53533 & n58324 ;
  assign n58326 = ~\pi1091  & ~n58325 ;
  assign n58327 = ~n58323 & n58326 ;
  assign n58328 = ~n58322 & ~n58327 ;
  assign n58329 = ~\pi0230  & n58328 ;
  assign n58330 = \pi0211  & \pi1139  ;
  assign n58331 = ~n57432 & ~n58330 ;
  assign n58332 = \pi1091  & ~n58331 ;
  assign n58333 = n54850 & ~n58332 ;
  assign n58334 = \pi1139  & n53865 ;
  assign n58335 = ~n57402 & ~n58334 ;
  assign n58336 = n57172 & n58335 ;
  assign n58337 = ~n58333 & ~n58336 ;
  assign n58338 = \pi0282  & ~\pi0314  ;
  assign n58339 = ~\pi0081  & \pi0282  ;
  assign n58340 = n53533 & n58339 ;
  assign n58341 = ~n58338 & ~n58340 ;
  assign n58342 = ~\pi1091  & ~n58324 ;
  assign n58343 = ~n56679 & ~n58342 ;
  assign n58344 = n58341 & ~n58343 ;
  assign n58345 = ~\pi0230  & ~n58344 ;
  assign n58346 = ~n58337 & n58345 ;
  assign n58347 = ~n58329 & ~n58346 ;
  assign n58348 = \pi0219  & n58051 ;
  assign n58349 = ~\pi0219  & ~n58331 ;
  assign n58350 = ~n58348 & ~n58349 ;
  assign n58351 = n56733 & n58350 ;
  assign n58352 = \pi0200  & ~n57486 ;
  assign n58353 = \pi0199  & \pi1140  ;
  assign n58354 = ~\pi0200  & ~n58307 ;
  assign n58355 = ~n58353 & n58354 ;
  assign n58356 = ~n58352 & ~n58355 ;
  assign n58357 = n53960 & ~n58356 ;
  assign n58358 = ~n58351 & ~n58357 ;
  assign n58359 = n58347 & n58358 ;
  assign n58360 = \pi1147  & ~n57606 ;
  assign n58361 = \pi1149  & ~n55693 ;
  assign n58362 = ~n58360 & ~n58361 ;
  assign n58363 = ~\pi1148  & ~n58362 ;
  assign n58364 = \pi0230  & n58363 ;
  assign n58365 = \pi1147  & n57172 ;
  assign n58366 = ~n20516 & n54642 ;
  assign n58367 = ~n58365 & ~n58366 ;
  assign n58368 = n57180 & n58367 ;
  assign n58369 = ~\pi1149  & n58368 ;
  assign n58370 = \pi1148  & ~n58369 ;
  assign n58371 = n57703 & ~n58360 ;
  assign n58372 = \pi0230  & ~n58371 ;
  assign n58373 = n58370 & n58372 ;
  assign n58374 = ~n58364 & ~n58373 ;
  assign n58375 = n58370 & ~n58371 ;
  assign n58376 = \pi0230  & ~n58363 ;
  assign n58377 = ~n58375 & n58376 ;
  assign n58378 = \pi1147  & ~\pi1148  ;
  assign n58379 = ~\pi1148  & n57241 ;
  assign n58380 = ~n57240 & n58379 ;
  assign n58381 = ~n58378 & ~n58380 ;
  assign n58382 = \pi1147  & ~n57325 ;
  assign n58383 = ~\pi0283  & ~n58382 ;
  assign n58384 = ~\pi0283  & n57350 ;
  assign n58385 = ~n57349 & n58384 ;
  assign n58386 = ~n58383 & ~n58385 ;
  assign n58387 = ~n58381 & ~n58386 ;
  assign n58388 = ~\pi1147  & ~n57917 ;
  assign n58389 = \pi1147  & ~n57361 ;
  assign n58390 = n57360 & n58389 ;
  assign n58391 = ~\pi0283  & \pi1148  ;
  assign n58392 = ~n58390 & n58391 ;
  assign n58393 = ~n58388 & n58392 ;
  assign n58394 = ~n58387 & ~n58393 ;
  assign n58395 = \pi0283  & ~\pi1147  ;
  assign n58396 = n57282 & n58395 ;
  assign n58397 = ~\pi0283  & ~\pi1149  ;
  assign n58398 = n54899 & n55919 ;
  assign n58399 = ~n57315 & n58398 ;
  assign n58400 = \pi1147  & ~n9948 ;
  assign n58401 = ~n55874 & n58400 ;
  assign n58402 = ~n56213 & n58401 ;
  assign n58403 = \pi1148  & ~n58402 ;
  assign n58404 = ~\pi1149  & n58403 ;
  assign n58405 = ~n58399 & n58404 ;
  assign n58406 = ~n58397 & ~n58405 ;
  assign n58407 = ~n58396 & ~n58406 ;
  assign n58408 = \pi1147  & n57375 ;
  assign n58409 = \pi1147  & ~n55926 ;
  assign n58410 = n57226 & n58409 ;
  assign n58411 = ~n58408 & ~n58410 ;
  assign n58412 = ~n52688 & ~n57664 ;
  assign n58413 = ~\pi1148  & ~n58412 ;
  assign n58414 = n58411 & n58413 ;
  assign n58415 = ~n58407 & ~n58414 ;
  assign n58416 = n58394 & ~n58415 ;
  assign n58417 = ~n58377 & ~n58416 ;
  assign n58418 = n58374 & ~n58417 ;
  assign n58419 = ~n57304 & ~n57305 ;
  assign n58420 = ~n55876 & n57257 ;
  assign n58421 = \pi1147  & ~n58420 ;
  assign n58422 = ~n58419 & n58421 ;
  assign n58423 = ~n57229 & n58421 ;
  assign n58424 = ~n57226 & n58423 ;
  assign n58425 = ~n58422 & ~n58424 ;
  assign n58426 = ~\pi1147  & ~n57271 ;
  assign n58427 = ~\pi1148  & ~n58426 ;
  assign n58428 = ~\pi1148  & n57269 ;
  assign n58429 = n57264 & n58428 ;
  assign n58430 = ~n58427 & ~n58429 ;
  assign n58431 = n58425 & ~n58430 ;
  assign n58432 = \pi0283  & n58431 ;
  assign n58433 = ~\pi1147  & n57267 ;
  assign n58434 = \pi1147  & ~n57317 ;
  assign n58435 = ~n57316 & n58434 ;
  assign n58436 = \pi1148  & ~n58435 ;
  assign n58437 = n9948 & ~n53559 ;
  assign n58438 = \pi1148  & n58437 ;
  assign n58439 = ~n55926 & n58438 ;
  assign n58440 = ~n58436 & ~n58439 ;
  assign n58441 = \pi0283  & ~n58440 ;
  assign n58442 = ~n58433 & n58441 ;
  assign n58443 = ~n58432 & ~n58442 ;
  assign n58444 = ~\pi1147  & ~n57208 ;
  assign n58445 = \pi1147  & ~n57195 ;
  assign n58446 = ~n57325 & n58445 ;
  assign n58447 = ~n9948 & n58446 ;
  assign n58448 = ~n57210 & n58446 ;
  assign n58449 = n57213 & n58448 ;
  assign n58450 = ~n58447 & ~n58449 ;
  assign n58451 = \pi1148  & n58450 ;
  assign n58452 = ~n58444 & n58451 ;
  assign n58453 = ~\pi1147  & ~n57220 ;
  assign n58454 = ~n57218 & n58453 ;
  assign n58455 = \pi1147  & ~n57324 ;
  assign n58456 = ~n57339 & n58455 ;
  assign n58457 = n57338 & n58456 ;
  assign n58458 = ~\pi1148  & ~n58457 ;
  assign n58459 = ~n58454 & n58458 ;
  assign n58460 = ~n58452 & ~n58459 ;
  assign n58461 = ~\pi0283  & ~n58460 ;
  assign n58462 = n58443 & ~n58461 ;
  assign n58463 = \pi1149  & n58374 ;
  assign n58464 = n58462 & n58463 ;
  assign n58465 = ~n58418 & ~n58464 ;
  assign n58466 = ~\pi0284  & ~n56376 ;
  assign n58467 = \pi1143  & n56376 ;
  assign n58468 = ~n52683 & n58467 ;
  assign n58469 = ~n58466 & ~n58468 ;
  assign n58470 = \pi0286  & ~n8696 ;
  assign n58471 = n1291 & n58470 ;
  assign n58472 = \pi0288  & \pi0289  ;
  assign n58473 = n58471 & n58472 ;
  assign n58474 = ~n12313 & n58473 ;
  assign n58475 = \pi0285  & n1291 ;
  assign n58476 = ~n12313 & n58475 ;
  assign n58477 = ~n58474 & ~n58476 ;
  assign n58478 = \pi0285  & n58472 ;
  assign n58479 = n58471 & n58478 ;
  assign n58480 = ~n12313 & n58479 ;
  assign n58481 = n9948 & ~n58480 ;
  assign n58482 = ~n58477 & n58481 ;
  assign n58483 = n55740 & n58472 ;
  assign n58484 = n58471 & n58483 ;
  assign n58485 = ~n12313 & n58484 ;
  assign n58486 = ~\pi0286  & \pi1093  ;
  assign n58487 = ~\pi1091  & n58486 ;
  assign n58488 = n8695 & n58487 ;
  assign n58489 = ~\pi0288  & ~\pi0289  ;
  assign n58490 = n58488 & n58489 ;
  assign n58491 = \pi0285  & ~n58490 ;
  assign n58492 = ~n58485 & n58491 ;
  assign n58493 = ~n58482 & ~n58492 ;
  assign n58494 = ~\pi0793  & ~n58493 ;
  assign n58495 = ~\pi0289  & n9248 ;
  assign n58496 = ~\pi0288  & ~n58495 ;
  assign n58497 = ~n1291 & n58488 ;
  assign n58498 = ~n12143 & n58488 ;
  assign n58499 = n12136 & n58498 ;
  assign n58500 = ~n58497 & ~n58499 ;
  assign n58501 = n58496 & ~n58500 ;
  assign n58502 = n9948 & ~n58501 ;
  assign n58503 = n1291 & ~n8696 ;
  assign n58504 = ~\pi0286  & ~n58503 ;
  assign n58505 = ~\pi0286  & ~n12143 ;
  assign n58506 = n12136 & n58505 ;
  assign n58507 = ~n58504 & ~n58506 ;
  assign n58508 = \pi0288  & ~n58471 ;
  assign n58509 = \pi0288  & ~n12143 ;
  assign n58510 = n12136 & n58509 ;
  assign n58511 = ~n58508 & ~n58510 ;
  assign n58512 = n58507 & ~n58511 ;
  assign n58513 = ~n1291 & n8696 ;
  assign n58514 = n8696 & ~n12143 ;
  assign n58515 = n12136 & n58514 ;
  assign n58516 = ~n58513 & ~n58515 ;
  assign n58517 = \pi0286  & n58496 ;
  assign n58518 = n58516 & n58517 ;
  assign n58519 = ~n58512 & ~n58518 ;
  assign n58520 = n58502 & n58519 ;
  assign n58521 = n8696 & n58496 ;
  assign n58522 = \pi0286  & ~n58521 ;
  assign n58523 = ~\pi0286  & ~\pi0288  ;
  assign n58524 = ~n58495 & n58523 ;
  assign n58525 = n8696 & n58524 ;
  assign n58526 = ~n9948 & ~n58525 ;
  assign n58527 = ~n58522 & n58526 ;
  assign n58528 = ~\pi0793  & ~n58527 ;
  assign n58529 = ~n58520 & n58528 ;
  assign n58530 = ~\pi0287  & \pi0457  ;
  assign n58531 = ~\pi0332  & ~n58530 ;
  assign n58532 = \pi0288  & ~n8696 ;
  assign n58533 = ~n58521 & ~n58532 ;
  assign n58534 = ~n11822 & n58533 ;
  assign n58535 = ~n12143 & n58533 ;
  assign n58536 = n12136 & n58535 ;
  assign n58537 = ~n58534 & ~n58536 ;
  assign n58538 = n11822 & ~n58533 ;
  assign n58539 = ~\pi0793  & ~n58538 ;
  assign n58540 = ~\pi0793  & ~n12143 ;
  assign n58541 = n12136 & n58540 ;
  assign n58542 = ~n58539 & ~n58541 ;
  assign n58543 = n58537 & ~n58542 ;
  assign n58544 = n58489 & n58500 ;
  assign n58545 = \pi0285  & ~\pi0289  ;
  assign n58546 = ~\pi0288  & ~n58545 ;
  assign n58547 = ~n58500 & n58546 ;
  assign n58548 = ~n58544 & ~n58547 ;
  assign n58549 = ~\pi0289  & ~n58511 ;
  assign n58550 = ~n58474 & ~n58549 ;
  assign n58551 = n58548 & n58550 ;
  assign n58552 = n9948 & ~n58551 ;
  assign n58553 = ~\pi0288  & n58488 ;
  assign n58554 = \pi0289  & ~n58553 ;
  assign n58555 = ~\pi0288  & n58545 ;
  assign n58556 = n58488 & n58555 ;
  assign n58557 = ~n9948 & ~n58556 ;
  assign n58558 = ~n58554 & n58557 ;
  assign n58559 = ~\pi0793  & ~n58558 ;
  assign n58560 = ~n58552 & n58559 ;
  assign n58561 = ~\pi0290  & \pi0476  ;
  assign n58562 = ~\pi0476  & ~\pi1048  ;
  assign n58563 = ~n58561 & ~n58562 ;
  assign n58564 = ~\pi0291  & \pi0476  ;
  assign n58565 = ~\pi0476  & ~\pi1049  ;
  assign n58566 = ~n58564 & ~n58565 ;
  assign n58567 = ~\pi0292  & \pi0476  ;
  assign n58568 = ~\pi0476  & ~\pi1084  ;
  assign n58569 = ~n58567 & ~n58568 ;
  assign n58570 = ~\pi0293  & \pi0476  ;
  assign n58571 = ~\pi0476  & ~\pi1059  ;
  assign n58572 = ~n58570 & ~n58571 ;
  assign n58573 = ~\pi0294  & \pi0476  ;
  assign n58574 = ~\pi0476  & ~\pi1072  ;
  assign n58575 = ~n58573 & ~n58574 ;
  assign n58576 = ~\pi0295  & \pi0476  ;
  assign n58577 = ~\pi0476  & ~\pi1053  ;
  assign n58578 = ~n58576 & ~n58577 ;
  assign n58579 = ~\pi0296  & \pi0476  ;
  assign n58580 = ~\pi0476  & ~\pi1037  ;
  assign n58581 = ~n58579 & ~n58580 ;
  assign n58582 = ~\pi0297  & \pi0476  ;
  assign n58583 = ~\pi0476  & ~\pi1044  ;
  assign n58584 = ~n58582 & ~n58583 ;
  assign n58585 = ~\pi0478  & \pi1044  ;
  assign n58586 = \pi0298  & \pi0478  ;
  assign n58587 = ~n58585 & ~n58586 ;
  assign n58588 = \pi0039  & ~n13396 ;
  assign n58589 = ~\pi0054  & ~\pi0093  ;
  assign n58590 = n1277 & n58589 ;
  assign n58591 = n1273 & n58590 ;
  assign n58592 = n11858 & n58591 ;
  assign n58593 = n2363 & n2364 ;
  assign n58594 = n1267 & n58593 ;
  assign n58595 = n58592 & n58594 ;
  assign n58596 = ~n15886 & n58595 ;
  assign n58597 = \pi0054  & n11858 ;
  assign n58598 = n1281 & n58597 ;
  assign n58599 = n1259 & n58593 ;
  assign n58600 = n1249 & n58599 ;
  assign n58601 = n58598 & n58600 ;
  assign n58602 = ~\pi0039  & ~n58601 ;
  assign n58603 = ~n58596 & n58602 ;
  assign n58604 = ~n58588 & ~n58603 ;
  assign n58605 = ~\pi0312  & n7672 ;
  assign n58606 = n13455 & n58605 ;
  assign n58607 = n1281 & n58606 ;
  assign n58608 = n1260 & n58607 ;
  assign n58609 = \pi0300  & ~n58608 ;
  assign n58610 = ~\pi0300  & ~\pi0312  ;
  assign n58611 = n13455 & n58610 ;
  assign n58612 = n1281 & n58611 ;
  assign n58613 = n1260 & n58612 ;
  assign n58614 = n7672 & n58613 ;
  assign n58615 = ~\pi0055  & ~n58614 ;
  assign n58616 = ~n58609 & n58615 ;
  assign n58617 = ~\pi0055  & ~\pi0301  ;
  assign n58618 = ~n58614 & n58617 ;
  assign n58619 = ~\pi0300  & \pi0301  ;
  assign n58620 = ~\pi0055  & n58619 ;
  assign n58621 = n58608 & n58620 ;
  assign n58622 = ~n58618 & ~n58621 ;
  assign n58623 = n6456 & n9948 ;
  assign n58624 = n6400 & ~n20516 ;
  assign n58625 = ~n58623 & ~n58624 ;
  assign n58626 = ~\pi1148  & n58625 ;
  assign n58627 = ~\pi0222  & ~\pi0223  ;
  assign n58628 = \pi0937  & ~n58627 ;
  assign n58629 = \pi0273  & n2522 ;
  assign n58630 = ~n58628 & ~n58629 ;
  assign n58631 = ~n2165 & n58630 ;
  assign n58632 = n58623 & n58631 ;
  assign n58633 = ~\pi0215  & ~\pi0273  ;
  assign n58634 = n2291 & n58633 ;
  assign n58635 = ~\pi0216  & \pi0833  ;
  assign n58636 = n6936 & n58635 ;
  assign n58637 = ~\pi0937  & n58636 ;
  assign n58638 = ~n58634 & ~n58637 ;
  assign n58639 = ~n20516 & ~n58638 ;
  assign n58640 = ~n58632 & ~n58639 ;
  assign n58641 = \pi0237  & n58630 ;
  assign n58642 = n58623 & n58641 ;
  assign n58643 = \pi0237  & n2650 ;
  assign n58644 = ~n20516 & n58643 ;
  assign n58645 = ~n58642 & ~n58644 ;
  assign n58646 = n58640 & n58645 ;
  assign n58647 = ~n58626 & n58646 ;
  assign n58648 = ~\pi0478  & \pi1049  ;
  assign n58649 = \pi0303  & \pi0478  ;
  assign n58650 = ~n58648 & ~n58649 ;
  assign n58651 = ~\pi0478  & \pi1048  ;
  assign n58652 = \pi0304  & \pi0478  ;
  assign n58653 = ~n58651 & ~n58652 ;
  assign n58654 = ~\pi0478  & \pi1084  ;
  assign n58655 = \pi0305  & \pi0478  ;
  assign n58656 = ~n58654 & ~n58655 ;
  assign n58657 = ~\pi0478  & \pi1059  ;
  assign n58658 = \pi0306  & \pi0478  ;
  assign n58659 = ~n58657 & ~n58658 ;
  assign n58660 = ~\pi0478  & \pi1053  ;
  assign n58661 = \pi0307  & \pi0478  ;
  assign n58662 = ~n58660 & ~n58661 ;
  assign n58663 = ~\pi0478  & \pi1037  ;
  assign n58664 = \pi0308  & \pi0478  ;
  assign n58665 = ~n58663 & ~n58664 ;
  assign n58666 = ~\pi0478  & \pi1072  ;
  assign n58667 = \pi0309  & \pi0478  ;
  assign n58668 = ~n58666 & ~n58667 ;
  assign n58669 = \pi1147  & n58625 ;
  assign n58670 = ~n6399 & n24388 ;
  assign n58671 = ~n20516 & n58670 ;
  assign n58672 = \pi0934  & ~n1295 ;
  assign n58673 = \pi0271  & n2291 ;
  assign n58674 = ~n58672 & ~n58673 ;
  assign n58675 = n58671 & ~n58674 ;
  assign n58676 = n2650 & ~n20516 ;
  assign n58677 = \pi0222  & ~\pi0934  ;
  assign n58678 = ~\pi0271  & n2522 ;
  assign n58679 = ~n58677 & ~n58678 ;
  assign n58680 = n58623 & n58679 ;
  assign n58681 = ~n58676 & ~n58680 ;
  assign n58682 = ~n58675 & n58681 ;
  assign n58683 = ~n58669 & n58682 ;
  assign n58684 = ~\pi0233  & ~n58683 ;
  assign n58685 = n58623 & ~n58679 ;
  assign n58686 = n2214 & n20516 ;
  assign n58687 = \pi1147  & ~n58686 ;
  assign n58688 = ~n58685 & n58687 ;
  assign n58689 = n58624 & n58674 ;
  assign n58690 = \pi0233  & ~n58689 ;
  assign n58691 = n58688 & n58690 ;
  assign n58692 = ~n2165 & n3058 ;
  assign n58693 = ~n2193 & n58692 ;
  assign n58694 = n9948 & n58693 ;
  assign n58695 = ~n58671 & ~n58694 ;
  assign n58696 = \pi0233  & ~\pi1147  ;
  assign n58697 = ~n58695 & n58696 ;
  assign n58698 = ~n58682 & n58697 ;
  assign n58699 = ~n58691 & ~n58698 ;
  assign n58700 = ~n58684 & n58699 ;
  assign n58701 = ~\pi0055  & ~\pi0311  ;
  assign n58702 = ~n58621 & ~n58701 ;
  assign n58703 = ~\pi0311  & n58620 ;
  assign n58704 = n58608 & n58703 ;
  assign n58705 = ~n58702 & ~n58704 ;
  assign n58706 = n7672 & n13455 ;
  assign n58707 = n1281 & n58706 ;
  assign n58708 = n1260 & n58707 ;
  assign n58709 = ~\pi0055  & \pi0312  ;
  assign n58710 = ~n58708 & n58709 ;
  assign n58711 = ~\pi0055  & ~\pi0312  ;
  assign n58712 = n58708 & n58711 ;
  assign n58713 = ~n58710 & ~n58712 ;
  assign n58714 = ~\pi0313  & \pi0954  ;
  assign n58715 = n1412 & n13153 ;
  assign n58716 = n15949 & n58715 ;
  assign n58717 = ~n15954 & ~n58716 ;
  assign n58718 = ~\pi0314  & n13153 ;
  assign n58719 = n1412 & n58718 ;
  assign n58720 = n15949 & n58719 ;
  assign n58721 = n8604 & ~n58720 ;
  assign n58722 = \pi0313  & \pi0954  ;
  assign n58723 = n11824 & ~n58722 ;
  assign n58724 = ~n58721 & n58723 ;
  assign n58725 = ~n58717 & n58724 ;
  assign n58726 = ~n58714 & ~n58725 ;
  assign n58727 = n17438 & n17439 ;
  assign n58728 = n7265 & n11858 ;
  assign n58729 = n17444 & ~n58728 ;
  assign n58730 = n58727 & n58729 ;
  assign n58731 = ~n2327 & ~n19776 ;
  assign n58732 = \pi0039  & ~n19776 ;
  assign n58733 = n18192 & n58732 ;
  assign n58734 = ~n58731 & ~n58733 ;
  assign n58735 = ~\pi0039  & ~n19776 ;
  assign n58736 = ~n17515 & n58735 ;
  assign n58737 = n17518 & n58735 ;
  assign n58738 = ~n17490 & n58737 ;
  assign n58739 = ~n58736 & ~n58738 ;
  assign n58740 = ~n17444 & ~n58728 ;
  assign n58741 = n58727 & ~n58740 ;
  assign n58742 = ~\pi0087  & n58741 ;
  assign n58743 = n58739 & n58742 ;
  assign n58744 = n58734 & n58743 ;
  assign n58745 = ~n58730 & ~n58744 ;
  assign n58746 = ~\pi0340  & n11822 ;
  assign n58747 = ~n12313 & n58746 ;
  assign n58748 = \pi0315  & ~n58747 ;
  assign n58749 = ~\pi0340  & \pi1080  ;
  assign n58750 = n11822 & n58749 ;
  assign n58751 = ~n12313 & n58750 ;
  assign n58752 = ~n58748 & ~n58751 ;
  assign n58753 = \pi0316  & ~n58747 ;
  assign n58754 = ~\pi0340  & \pi1047  ;
  assign n58755 = n11822 & n58754 ;
  assign n58756 = ~n12313 & n58755 ;
  assign n58757 = ~n58753 & ~n58756 ;
  assign n58758 = ~\pi0330  & n11822 ;
  assign n58759 = ~n12313 & n58758 ;
  assign n58760 = \pi0317  & ~n58759 ;
  assign n58761 = ~\pi0330  & \pi1078  ;
  assign n58762 = n11822 & n58761 ;
  assign n58763 = ~n12313 & n58762 ;
  assign n58764 = ~n58760 & ~n58763 ;
  assign n58765 = ~\pi0341  & n11822 ;
  assign n58766 = ~n12313 & n58765 ;
  assign n58767 = \pi0318  & ~n58766 ;
  assign n58768 = ~\pi0341  & \pi1074  ;
  assign n58769 = n11822 & n58768 ;
  assign n58770 = ~n12313 & n58769 ;
  assign n58771 = ~n58767 & ~n58770 ;
  assign n58772 = \pi0319  & ~n58766 ;
  assign n58773 = ~\pi0341  & \pi1072  ;
  assign n58774 = n11822 & n58773 ;
  assign n58775 = ~n12313 & n58774 ;
  assign n58776 = ~n58772 & ~n58775 ;
  assign n58777 = \pi0320  & ~n58747 ;
  assign n58778 = ~\pi0340  & \pi1048  ;
  assign n58779 = n11822 & n58778 ;
  assign n58780 = ~n12313 & n58779 ;
  assign n58781 = ~n58777 & ~n58780 ;
  assign n58782 = \pi0321  & ~n58747 ;
  assign n58783 = ~\pi0340  & \pi1058  ;
  assign n58784 = n11822 & n58783 ;
  assign n58785 = ~n12313 & n58784 ;
  assign n58786 = ~n58782 & ~n58785 ;
  assign n58787 = \pi0322  & ~n58747 ;
  assign n58788 = ~\pi0340  & \pi1051  ;
  assign n58789 = n11822 & n58788 ;
  assign n58790 = ~n12313 & n58789 ;
  assign n58791 = ~n58787 & ~n58790 ;
  assign n58792 = \pi0323  & ~n58747 ;
  assign n58793 = ~\pi0340  & \pi1065  ;
  assign n58794 = n11822 & n58793 ;
  assign n58795 = ~n12313 & n58794 ;
  assign n58796 = ~n58792 & ~n58795 ;
  assign n58797 = \pi0324  & ~n58766 ;
  assign n58798 = ~\pi0341  & \pi1086  ;
  assign n58799 = n11822 & n58798 ;
  assign n58800 = ~n12313 & n58799 ;
  assign n58801 = ~n58797 & ~n58800 ;
  assign n58802 = \pi0325  & ~n58766 ;
  assign n58803 = ~\pi0341  & \pi1063  ;
  assign n58804 = n11822 & n58803 ;
  assign n58805 = ~n12313 & n58804 ;
  assign n58806 = ~n58802 & ~n58805 ;
  assign n58807 = \pi0326  & ~n58766 ;
  assign n58808 = ~\pi0341  & \pi1057  ;
  assign n58809 = n11822 & n58808 ;
  assign n58810 = ~n12313 & n58809 ;
  assign n58811 = ~n58807 & ~n58810 ;
  assign n58812 = \pi0327  & ~n58747 ;
  assign n58813 = ~\pi0340  & \pi1040  ;
  assign n58814 = n11822 & n58813 ;
  assign n58815 = ~n12313 & n58814 ;
  assign n58816 = ~n58812 & ~n58815 ;
  assign n58817 = \pi0328  & ~n58766 ;
  assign n58818 = ~\pi0341  & \pi1058  ;
  assign n58819 = n11822 & n58818 ;
  assign n58820 = ~n12313 & n58819 ;
  assign n58821 = ~n58817 & ~n58820 ;
  assign n58822 = \pi0329  & ~n58766 ;
  assign n58823 = ~\pi0341  & \pi1043  ;
  assign n58824 = n11822 & n58823 ;
  assign n58825 = ~n12313 & n58824 ;
  assign n58826 = ~n58822 & ~n58825 ;
  assign n58827 = ~\pi0330  & ~n11822 ;
  assign n58828 = ~\pi0330  & ~n12143 ;
  assign n58829 = n12136 & n58828 ;
  assign n58830 = ~n58827 & ~n58829 ;
  assign n58831 = ~n58747 & n58830 ;
  assign n58832 = \pi1092  & ~n6703 ;
  assign n58833 = ~n58831 & n58832 ;
  assign n58834 = ~\pi0331  & ~n11822 ;
  assign n58835 = ~\pi0331  & ~n12143 ;
  assign n58836 = n12136 & n58835 ;
  assign n58837 = ~n58834 & ~n58836 ;
  assign n58838 = ~n58766 & n58837 ;
  assign n58839 = n58832 & ~n58838 ;
  assign n58840 = \pi0039  & \pi0287  ;
  assign n58841 = n1281 & n58840 ;
  assign n58842 = n1260 & n58841 ;
  assign n58843 = ~\pi0038  & ~n58842 ;
  assign n58844 = ~n50141 & ~n58843 ;
  assign n58845 = ~\pi0097  & n13114 ;
  assign n58846 = n1586 & n58845 ;
  assign n58847 = ~n15534 & ~n58846 ;
  assign n58848 = n1718 & ~n58847 ;
  assign n58849 = n1320 & n15535 ;
  assign n58850 = n1266 & n58849 ;
  assign n58851 = n13114 & n58850 ;
  assign n58852 = ~\pi0097  & n58851 ;
  assign n58853 = n1586 & n58852 ;
  assign n58854 = ~\pi0070  & ~n58853 ;
  assign n58855 = ~n58848 & n58854 ;
  assign n58856 = \pi0332  & n10903 ;
  assign n58857 = ~n1864 & n58856 ;
  assign n58858 = ~n58853 & ~n58857 ;
  assign n58859 = n50266 & ~n58858 ;
  assign n58860 = ~n58855 & n58859 ;
  assign n58861 = ~n58844 & ~n58860 ;
  assign n58862 = \pi0333  & ~n58766 ;
  assign n58863 = ~\pi0341  & \pi1040  ;
  assign n58864 = n11822 & n58863 ;
  assign n58865 = ~n12313 & n58864 ;
  assign n58866 = ~n58862 & ~n58865 ;
  assign n58867 = \pi0334  & ~n58766 ;
  assign n58868 = ~\pi0341  & \pi1065  ;
  assign n58869 = n11822 & n58868 ;
  assign n58870 = ~n12313 & n58869 ;
  assign n58871 = ~n58867 & ~n58870 ;
  assign n58872 = \pi0335  & ~n58766 ;
  assign n58873 = ~\pi0341  & \pi1069  ;
  assign n58874 = n11822 & n58873 ;
  assign n58875 = ~n12313 & n58874 ;
  assign n58876 = ~n58872 & ~n58875 ;
  assign n58877 = \pi0336  & ~n58759 ;
  assign n58878 = ~\pi0330  & \pi1070  ;
  assign n58879 = n11822 & n58878 ;
  assign n58880 = ~n12313 & n58879 ;
  assign n58881 = ~n58877 & ~n58880 ;
  assign n58882 = \pi0337  & ~n58759 ;
  assign n58883 = ~\pi0330  & \pi1044  ;
  assign n58884 = n11822 & n58883 ;
  assign n58885 = ~n12313 & n58884 ;
  assign n58886 = ~n58882 & ~n58885 ;
  assign n58887 = \pi0338  & ~n58759 ;
  assign n58888 = ~\pi0330  & \pi1072  ;
  assign n58889 = n11822 & n58888 ;
  assign n58890 = ~n12313 & n58889 ;
  assign n58891 = ~n58887 & ~n58890 ;
  assign n58892 = \pi0339  & ~n58759 ;
  assign n58893 = ~\pi0330  & \pi1086  ;
  assign n58894 = n11822 & n58893 ;
  assign n58895 = ~n12313 & n58894 ;
  assign n58896 = ~n58892 & ~n58895 ;
  assign n58897 = ~\pi0331  & n11822 ;
  assign n58898 = ~n12313 & n58897 ;
  assign n58899 = ~\pi0340  & ~n11822 ;
  assign n58900 = ~\pi0340  & ~n12143 ;
  assign n58901 = n12136 & n58900 ;
  assign n58902 = ~n58899 & ~n58901 ;
  assign n58903 = \pi1091  & \pi1093  ;
  assign n58904 = \pi1092  & ~n58903 ;
  assign n58905 = n58902 & n58904 ;
  assign n58906 = ~n58898 & n58905 ;
  assign n58907 = ~\pi0341  & ~n11822 ;
  assign n58908 = ~\pi0341  & ~n12143 ;
  assign n58909 = n12136 & n58908 ;
  assign n58910 = ~n58907 & ~n58909 ;
  assign n58911 = ~n58759 & n58910 ;
  assign n58912 = n58904 & ~n58911 ;
  assign n58913 = \pi0342  & ~n58747 ;
  assign n58914 = ~\pi0340  & \pi1049  ;
  assign n58915 = n11822 & n58914 ;
  assign n58916 = ~n12313 & n58915 ;
  assign n58917 = ~n58913 & ~n58916 ;
  assign n58918 = \pi0343  & ~n58747 ;
  assign n58919 = ~\pi0340  & \pi1062  ;
  assign n58920 = n11822 & n58919 ;
  assign n58921 = ~n12313 & n58920 ;
  assign n58922 = ~n58918 & ~n58921 ;
  assign n58923 = \pi0344  & ~n58747 ;
  assign n58924 = ~\pi0340  & \pi1069  ;
  assign n58925 = n11822 & n58924 ;
  assign n58926 = ~n12313 & n58925 ;
  assign n58927 = ~n58923 & ~n58926 ;
  assign n58928 = \pi0345  & ~n58747 ;
  assign n58929 = ~\pi0340  & \pi1039  ;
  assign n58930 = n11822 & n58929 ;
  assign n58931 = ~n12313 & n58930 ;
  assign n58932 = ~n58928 & ~n58931 ;
  assign n58933 = \pi0346  & ~n58747 ;
  assign n58934 = ~\pi0340  & \pi1067  ;
  assign n58935 = n11822 & n58934 ;
  assign n58936 = ~n12313 & n58935 ;
  assign n58937 = ~n58933 & ~n58936 ;
  assign n58938 = \pi0347  & ~n58747 ;
  assign n58939 = ~\pi0340  & \pi1055  ;
  assign n58940 = n11822 & n58939 ;
  assign n58941 = ~n12313 & n58940 ;
  assign n58942 = ~n58938 & ~n58941 ;
  assign n58943 = \pi0348  & ~n58747 ;
  assign n58944 = ~\pi0340  & \pi1087  ;
  assign n58945 = n11822 & n58944 ;
  assign n58946 = ~n12313 & n58945 ;
  assign n58947 = ~n58943 & ~n58946 ;
  assign n58948 = \pi0349  & ~n58747 ;
  assign n58949 = ~\pi0340  & \pi1043  ;
  assign n58950 = n11822 & n58949 ;
  assign n58951 = ~n12313 & n58950 ;
  assign n58952 = ~n58948 & ~n58951 ;
  assign n58953 = \pi0350  & ~n58747 ;
  assign n58954 = ~\pi0340  & \pi1035  ;
  assign n58955 = n11822 & n58954 ;
  assign n58956 = ~n12313 & n58955 ;
  assign n58957 = ~n58953 & ~n58956 ;
  assign n58958 = \pi0351  & ~n58747 ;
  assign n58959 = ~\pi0340  & \pi1079  ;
  assign n58960 = n11822 & n58959 ;
  assign n58961 = ~n12313 & n58960 ;
  assign n58962 = ~n58958 & ~n58961 ;
  assign n58963 = \pi0352  & ~n58747 ;
  assign n58964 = ~\pi0340  & \pi1078  ;
  assign n58965 = n11822 & n58964 ;
  assign n58966 = ~n12313 & n58965 ;
  assign n58967 = ~n58963 & ~n58966 ;
  assign n58968 = \pi0353  & ~n58747 ;
  assign n58969 = ~\pi0340  & \pi1063  ;
  assign n58970 = n11822 & n58969 ;
  assign n58971 = ~n12313 & n58970 ;
  assign n58972 = ~n58968 & ~n58971 ;
  assign n58973 = \pi0354  & ~n58747 ;
  assign n58974 = ~\pi0340  & \pi1045  ;
  assign n58975 = n11822 & n58974 ;
  assign n58976 = ~n12313 & n58975 ;
  assign n58977 = ~n58973 & ~n58976 ;
  assign n58978 = \pi0355  & ~n58747 ;
  assign n58979 = ~\pi0340  & \pi1084  ;
  assign n58980 = n11822 & n58979 ;
  assign n58981 = ~n12313 & n58980 ;
  assign n58982 = ~n58978 & ~n58981 ;
  assign n58983 = \pi0356  & ~n58747 ;
  assign n58984 = ~\pi0340  & \pi1081  ;
  assign n58985 = n11822 & n58984 ;
  assign n58986 = ~n12313 & n58985 ;
  assign n58987 = ~n58983 & ~n58986 ;
  assign n58988 = \pi0357  & ~n58747 ;
  assign n58989 = ~\pi0340  & \pi1076  ;
  assign n58990 = n11822 & n58989 ;
  assign n58991 = ~n12313 & n58990 ;
  assign n58992 = ~n58988 & ~n58991 ;
  assign n58993 = \pi0358  & ~n58747 ;
  assign n58994 = ~\pi0340  & \pi1071  ;
  assign n58995 = n11822 & n58994 ;
  assign n58996 = ~n12313 & n58995 ;
  assign n58997 = ~n58993 & ~n58996 ;
  assign n58998 = \pi0359  & ~n58747 ;
  assign n58999 = ~\pi0340  & \pi1068  ;
  assign n59000 = n11822 & n58999 ;
  assign n59001 = ~n12313 & n59000 ;
  assign n59002 = ~n58998 & ~n59001 ;
  assign n59003 = \pi0360  & ~n58747 ;
  assign n59004 = ~\pi0340  & \pi1042  ;
  assign n59005 = n11822 & n59004 ;
  assign n59006 = ~n12313 & n59005 ;
  assign n59007 = ~n59003 & ~n59006 ;
  assign n59008 = \pi0361  & ~n58747 ;
  assign n59009 = ~\pi0340  & \pi1059  ;
  assign n59010 = n11822 & n59009 ;
  assign n59011 = ~n12313 & n59010 ;
  assign n59012 = ~n59008 & ~n59011 ;
  assign n59013 = \pi0362  & ~n58747 ;
  assign n59014 = ~\pi0340  & \pi1070  ;
  assign n59015 = n11822 & n59014 ;
  assign n59016 = ~n12313 & n59015 ;
  assign n59017 = ~n59013 & ~n59016 ;
  assign n59018 = \pi0363  & ~n58759 ;
  assign n59019 = ~\pi0330  & \pi1049  ;
  assign n59020 = n11822 & n59019 ;
  assign n59021 = ~n12313 & n59020 ;
  assign n59022 = ~n59018 & ~n59021 ;
  assign n59023 = \pi0364  & ~n58759 ;
  assign n59024 = ~\pi0330  & \pi1062  ;
  assign n59025 = n11822 & n59024 ;
  assign n59026 = ~n12313 & n59025 ;
  assign n59027 = ~n59023 & ~n59026 ;
  assign n59028 = \pi0365  & ~n58759 ;
  assign n59029 = ~\pi0330  & \pi1065  ;
  assign n59030 = n11822 & n59029 ;
  assign n59031 = ~n12313 & n59030 ;
  assign n59032 = ~n59028 & ~n59031 ;
  assign n59033 = \pi0366  & ~n58759 ;
  assign n59034 = ~\pi0330  & \pi1069  ;
  assign n59035 = n11822 & n59034 ;
  assign n59036 = ~n12313 & n59035 ;
  assign n59037 = ~n59033 & ~n59036 ;
  assign n59038 = \pi0367  & ~n58759 ;
  assign n59039 = ~\pi0330  & \pi1039  ;
  assign n59040 = n11822 & n59039 ;
  assign n59041 = ~n12313 & n59040 ;
  assign n59042 = ~n59038 & ~n59041 ;
  assign n59043 = \pi0368  & ~n58759 ;
  assign n59044 = ~\pi0330  & \pi1067  ;
  assign n59045 = n11822 & n59044 ;
  assign n59046 = ~n12313 & n59045 ;
  assign n59047 = ~n59043 & ~n59046 ;
  assign n59048 = \pi0369  & ~n58759 ;
  assign n59049 = ~\pi0330  & \pi1080  ;
  assign n59050 = n11822 & n59049 ;
  assign n59051 = ~n12313 & n59050 ;
  assign n59052 = ~n59048 & ~n59051 ;
  assign n59053 = \pi0370  & ~n58759 ;
  assign n59054 = ~\pi0330  & \pi1055  ;
  assign n59055 = n11822 & n59054 ;
  assign n59056 = ~n12313 & n59055 ;
  assign n59057 = ~n59053 & ~n59056 ;
  assign n59058 = \pi0371  & ~n58759 ;
  assign n59059 = ~\pi0330  & \pi1051  ;
  assign n59060 = n11822 & n59059 ;
  assign n59061 = ~n12313 & n59060 ;
  assign n59062 = ~n59058 & ~n59061 ;
  assign n59063 = \pi0372  & ~n58759 ;
  assign n59064 = ~\pi0330  & \pi1048  ;
  assign n59065 = n11822 & n59064 ;
  assign n59066 = ~n12313 & n59065 ;
  assign n59067 = ~n59063 & ~n59066 ;
  assign n59068 = \pi0373  & ~n58759 ;
  assign n59069 = ~\pi0330  & \pi1087  ;
  assign n59070 = n11822 & n59069 ;
  assign n59071 = ~n12313 & n59070 ;
  assign n59072 = ~n59068 & ~n59071 ;
  assign n59073 = \pi0374  & ~n58759 ;
  assign n59074 = ~\pi0330  & \pi1035  ;
  assign n59075 = n11822 & n59074 ;
  assign n59076 = ~n12313 & n59075 ;
  assign n59077 = ~n59073 & ~n59076 ;
  assign n59078 = \pi0375  & ~n58759 ;
  assign n59079 = ~\pi0330  & \pi1047  ;
  assign n59080 = n11822 & n59079 ;
  assign n59081 = ~n12313 & n59080 ;
  assign n59082 = ~n59078 & ~n59081 ;
  assign n59083 = \pi0376  & ~n58759 ;
  assign n59084 = ~\pi0330  & \pi1079  ;
  assign n59085 = n11822 & n59084 ;
  assign n59086 = ~n12313 & n59085 ;
  assign n59087 = ~n59083 & ~n59086 ;
  assign n59088 = \pi0377  & ~n58759 ;
  assign n59089 = ~\pi0330  & \pi1074  ;
  assign n59090 = n11822 & n59089 ;
  assign n59091 = ~n12313 & n59090 ;
  assign n59092 = ~n59088 & ~n59091 ;
  assign n59093 = \pi0378  & ~n58759 ;
  assign n59094 = ~\pi0330  & \pi1063  ;
  assign n59095 = n11822 & n59094 ;
  assign n59096 = ~n12313 & n59095 ;
  assign n59097 = ~n59093 & ~n59096 ;
  assign n59098 = \pi0379  & ~n58759 ;
  assign n59099 = ~\pi0330  & \pi1045  ;
  assign n59100 = n11822 & n59099 ;
  assign n59101 = ~n12313 & n59100 ;
  assign n59102 = ~n59098 & ~n59101 ;
  assign n59103 = \pi0380  & ~n58759 ;
  assign n59104 = ~\pi0330  & \pi1084  ;
  assign n59105 = n11822 & n59104 ;
  assign n59106 = ~n12313 & n59105 ;
  assign n59107 = ~n59103 & ~n59106 ;
  assign n59108 = \pi0381  & ~n58759 ;
  assign n59109 = ~\pi0330  & \pi1081  ;
  assign n59110 = n11822 & n59109 ;
  assign n59111 = ~n12313 & n59110 ;
  assign n59112 = ~n59108 & ~n59111 ;
  assign n59113 = \pi0382  & ~n58759 ;
  assign n59114 = ~\pi0330  & \pi1076  ;
  assign n59115 = n11822 & n59114 ;
  assign n59116 = ~n12313 & n59115 ;
  assign n59117 = ~n59113 & ~n59116 ;
  assign n59118 = \pi0383  & ~n58759 ;
  assign n59119 = ~\pi0330  & \pi1071  ;
  assign n59120 = n11822 & n59119 ;
  assign n59121 = ~n12313 & n59120 ;
  assign n59122 = ~n59118 & ~n59121 ;
  assign n59123 = \pi0384  & ~n58759 ;
  assign n59124 = ~\pi0330  & \pi1068  ;
  assign n59125 = n11822 & n59124 ;
  assign n59126 = ~n12313 & n59125 ;
  assign n59127 = ~n59123 & ~n59126 ;
  assign n59128 = \pi0385  & ~n58759 ;
  assign n59129 = ~\pi0330  & \pi1042  ;
  assign n59130 = n11822 & n59129 ;
  assign n59131 = ~n12313 & n59130 ;
  assign n59132 = ~n59128 & ~n59131 ;
  assign n59133 = \pi0386  & ~n58759 ;
  assign n59134 = ~\pi0330  & \pi1059  ;
  assign n59135 = n11822 & n59134 ;
  assign n59136 = ~n12313 & n59135 ;
  assign n59137 = ~n59133 & ~n59136 ;
  assign n59138 = \pi0387  & ~n58759 ;
  assign n59139 = ~\pi0330  & \pi1053  ;
  assign n59140 = n11822 & n59139 ;
  assign n59141 = ~n12313 & n59140 ;
  assign n59142 = ~n59138 & ~n59141 ;
  assign n59143 = \pi0388  & ~n58759 ;
  assign n59144 = ~\pi0330  & \pi1037  ;
  assign n59145 = n11822 & n59144 ;
  assign n59146 = ~n12313 & n59145 ;
  assign n59147 = ~n59143 & ~n59146 ;
  assign n59148 = \pi0389  & ~n58759 ;
  assign n59149 = ~\pi0330  & \pi1036  ;
  assign n59150 = n11822 & n59149 ;
  assign n59151 = ~n12313 & n59150 ;
  assign n59152 = ~n59148 & ~n59151 ;
  assign n59153 = \pi0390  & ~n58766 ;
  assign n59154 = ~\pi0341  & \pi1049  ;
  assign n59155 = n11822 & n59154 ;
  assign n59156 = ~n12313 & n59155 ;
  assign n59157 = ~n59153 & ~n59156 ;
  assign n59158 = \pi0391  & ~n58766 ;
  assign n59159 = ~\pi0341  & \pi1062  ;
  assign n59160 = n11822 & n59159 ;
  assign n59161 = ~n12313 & n59160 ;
  assign n59162 = ~n59158 & ~n59161 ;
  assign n59163 = \pi0392  & ~n58766 ;
  assign n59164 = ~\pi0341  & \pi1039  ;
  assign n59165 = n11822 & n59164 ;
  assign n59166 = ~n12313 & n59165 ;
  assign n59167 = ~n59163 & ~n59166 ;
  assign n59168 = \pi0393  & ~n58766 ;
  assign n59169 = ~\pi0341  & \pi1067  ;
  assign n59170 = n11822 & n59169 ;
  assign n59171 = ~n12313 & n59170 ;
  assign n59172 = ~n59168 & ~n59171 ;
  assign n59173 = \pi0394  & ~n58766 ;
  assign n59174 = ~\pi0341  & \pi1080  ;
  assign n59175 = n11822 & n59174 ;
  assign n59176 = ~n12313 & n59175 ;
  assign n59177 = ~n59173 & ~n59176 ;
  assign n59178 = \pi0395  & ~n58766 ;
  assign n59179 = ~\pi0341  & \pi1055  ;
  assign n59180 = n11822 & n59179 ;
  assign n59181 = ~n12313 & n59180 ;
  assign n59182 = ~n59178 & ~n59181 ;
  assign n59183 = \pi0396  & ~n58766 ;
  assign n59184 = ~\pi0341  & \pi1051  ;
  assign n59185 = n11822 & n59184 ;
  assign n59186 = ~n12313 & n59185 ;
  assign n59187 = ~n59183 & ~n59186 ;
  assign n59188 = \pi0397  & ~n58766 ;
  assign n59189 = ~\pi0341  & \pi1048  ;
  assign n59190 = n11822 & n59189 ;
  assign n59191 = ~n12313 & n59190 ;
  assign n59192 = ~n59188 & ~n59191 ;
  assign n59193 = \pi0398  & ~n58766 ;
  assign n59194 = ~\pi0341  & \pi1087  ;
  assign n59195 = n11822 & n59194 ;
  assign n59196 = ~n12313 & n59195 ;
  assign n59197 = ~n59193 & ~n59196 ;
  assign n59198 = \pi0399  & ~n58766 ;
  assign n59199 = ~\pi0341  & \pi1047  ;
  assign n59200 = n11822 & n59199 ;
  assign n59201 = ~n12313 & n59200 ;
  assign n59202 = ~n59198 & ~n59201 ;
  assign n59203 = \pi0400  & ~n58766 ;
  assign n59204 = ~\pi0341  & \pi1035  ;
  assign n59205 = n11822 & n59204 ;
  assign n59206 = ~n12313 & n59205 ;
  assign n59207 = ~n59203 & ~n59206 ;
  assign n59208 = \pi0401  & ~n58766 ;
  assign n59209 = ~\pi0341  & \pi1079  ;
  assign n59210 = n11822 & n59209 ;
  assign n59211 = ~n12313 & n59210 ;
  assign n59212 = ~n59208 & ~n59211 ;
  assign n59213 = \pi0402  & ~n58766 ;
  assign n59214 = ~\pi0341  & \pi1078  ;
  assign n59215 = n11822 & n59214 ;
  assign n59216 = ~n12313 & n59215 ;
  assign n59217 = ~n59213 & ~n59216 ;
  assign n59218 = \pi0403  & ~n58766 ;
  assign n59219 = ~\pi0341  & \pi1045  ;
  assign n59220 = n11822 & n59219 ;
  assign n59221 = ~n12313 & n59220 ;
  assign n59222 = ~n59218 & ~n59221 ;
  assign n59223 = \pi0404  & ~n58766 ;
  assign n59224 = ~\pi0341  & \pi1084  ;
  assign n59225 = n11822 & n59224 ;
  assign n59226 = ~n12313 & n59225 ;
  assign n59227 = ~n59223 & ~n59226 ;
  assign n59228 = \pi0405  & ~n58766 ;
  assign n59229 = ~\pi0341  & \pi1081  ;
  assign n59230 = n11822 & n59229 ;
  assign n59231 = ~n12313 & n59230 ;
  assign n59232 = ~n59228 & ~n59231 ;
  assign n59233 = \pi0406  & ~n58766 ;
  assign n59234 = ~\pi0341  & \pi1076  ;
  assign n59235 = n11822 & n59234 ;
  assign n59236 = ~n12313 & n59235 ;
  assign n59237 = ~n59233 & ~n59236 ;
  assign n59238 = \pi0407  & ~n58766 ;
  assign n59239 = ~\pi0341  & \pi1071  ;
  assign n59240 = n11822 & n59239 ;
  assign n59241 = ~n12313 & n59240 ;
  assign n59242 = ~n59238 & ~n59241 ;
  assign n59243 = \pi0408  & ~n58766 ;
  assign n59244 = ~\pi0341  & \pi1068  ;
  assign n59245 = n11822 & n59244 ;
  assign n59246 = ~n12313 & n59245 ;
  assign n59247 = ~n59243 & ~n59246 ;
  assign n59248 = \pi0409  & ~n58766 ;
  assign n59249 = ~\pi0341  & \pi1042  ;
  assign n59250 = n11822 & n59249 ;
  assign n59251 = ~n12313 & n59250 ;
  assign n59252 = ~n59248 & ~n59251 ;
  assign n59253 = \pi0410  & ~n58766 ;
  assign n59254 = ~\pi0341  & \pi1059  ;
  assign n59255 = n11822 & n59254 ;
  assign n59256 = ~n12313 & n59255 ;
  assign n59257 = ~n59253 & ~n59256 ;
  assign n59258 = \pi0411  & ~n58766 ;
  assign n59259 = ~\pi0341  & \pi1053  ;
  assign n59260 = n11822 & n59259 ;
  assign n59261 = ~n12313 & n59260 ;
  assign n59262 = ~n59258 & ~n59261 ;
  assign n59263 = \pi0412  & ~n58766 ;
  assign n59264 = ~\pi0341  & \pi1037  ;
  assign n59265 = n11822 & n59264 ;
  assign n59266 = ~n12313 & n59265 ;
  assign n59267 = ~n59263 & ~n59266 ;
  assign n59268 = \pi0413  & ~n58766 ;
  assign n59269 = ~\pi0341  & \pi1036  ;
  assign n59270 = n11822 & n59269 ;
  assign n59271 = ~n12313 & n59270 ;
  assign n59272 = ~n59268 & ~n59271 ;
  assign n59273 = \pi0414  & ~n58898 ;
  assign n59274 = ~\pi0331  & \pi1049  ;
  assign n59275 = n11822 & n59274 ;
  assign n59276 = ~n12313 & n59275 ;
  assign n59277 = ~n59273 & ~n59276 ;
  assign n59278 = \pi0415  & ~n58898 ;
  assign n59279 = ~\pi0331  & \pi1062  ;
  assign n59280 = n11822 & n59279 ;
  assign n59281 = ~n12313 & n59280 ;
  assign n59282 = ~n59278 & ~n59281 ;
  assign n59283 = \pi0416  & ~n58898 ;
  assign n59284 = ~\pi0331  & \pi1069  ;
  assign n59285 = n11822 & n59284 ;
  assign n59286 = ~n12313 & n59285 ;
  assign n59287 = ~n59283 & ~n59286 ;
  assign n59288 = \pi0417  & ~n58898 ;
  assign n59289 = ~\pi0331  & \pi1039  ;
  assign n59290 = n11822 & n59289 ;
  assign n59291 = ~n12313 & n59290 ;
  assign n59292 = ~n59288 & ~n59291 ;
  assign n59293 = \pi0418  & ~n58898 ;
  assign n59294 = ~\pi0331  & \pi1067  ;
  assign n59295 = n11822 & n59294 ;
  assign n59296 = ~n12313 & n59295 ;
  assign n59297 = ~n59293 & ~n59296 ;
  assign n59298 = \pi0419  & ~n58898 ;
  assign n59299 = ~\pi0331  & \pi1080  ;
  assign n59300 = n11822 & n59299 ;
  assign n59301 = ~n12313 & n59300 ;
  assign n59302 = ~n59298 & ~n59301 ;
  assign n59303 = \pi0420  & ~n58898 ;
  assign n59304 = ~\pi0331  & \pi1055  ;
  assign n59305 = n11822 & n59304 ;
  assign n59306 = ~n12313 & n59305 ;
  assign n59307 = ~n59303 & ~n59306 ;
  assign n59308 = \pi0421  & ~n58898 ;
  assign n59309 = ~\pi0331  & \pi1051  ;
  assign n59310 = n11822 & n59309 ;
  assign n59311 = ~n12313 & n59310 ;
  assign n59312 = ~n59308 & ~n59311 ;
  assign n59313 = \pi0422  & ~n58898 ;
  assign n59314 = ~\pi0331  & \pi1048  ;
  assign n59315 = n11822 & n59314 ;
  assign n59316 = ~n12313 & n59315 ;
  assign n59317 = ~n59313 & ~n59316 ;
  assign n59318 = \pi0423  & ~n58898 ;
  assign n59319 = ~\pi0331  & \pi1087  ;
  assign n59320 = n11822 & n59319 ;
  assign n59321 = ~n12313 & n59320 ;
  assign n59322 = ~n59318 & ~n59321 ;
  assign n59323 = \pi0424  & ~n58898 ;
  assign n59324 = ~\pi0331  & \pi1047  ;
  assign n59325 = n11822 & n59324 ;
  assign n59326 = ~n12313 & n59325 ;
  assign n59327 = ~n59323 & ~n59326 ;
  assign n59328 = \pi0425  & ~n58898 ;
  assign n59329 = ~\pi0331  & \pi1035  ;
  assign n59330 = n11822 & n59329 ;
  assign n59331 = ~n12313 & n59330 ;
  assign n59332 = ~n59328 & ~n59331 ;
  assign n59333 = \pi0426  & ~n58898 ;
  assign n59334 = ~\pi0331  & \pi1079  ;
  assign n59335 = n11822 & n59334 ;
  assign n59336 = ~n12313 & n59335 ;
  assign n59337 = ~n59333 & ~n59336 ;
  assign n59338 = \pi0427  & ~n58898 ;
  assign n59339 = ~\pi0331  & \pi1078  ;
  assign n59340 = n11822 & n59339 ;
  assign n59341 = ~n12313 & n59340 ;
  assign n59342 = ~n59338 & ~n59341 ;
  assign n59343 = \pi0428  & ~n58898 ;
  assign n59344 = ~\pi0331  & \pi1045  ;
  assign n59345 = n11822 & n59344 ;
  assign n59346 = ~n12313 & n59345 ;
  assign n59347 = ~n59343 & ~n59346 ;
  assign n59348 = \pi0429  & ~n58898 ;
  assign n59349 = ~\pi0331  & \pi1084  ;
  assign n59350 = n11822 & n59349 ;
  assign n59351 = ~n12313 & n59350 ;
  assign n59352 = ~n59348 & ~n59351 ;
  assign n59353 = \pi0430  & ~n58898 ;
  assign n59354 = ~\pi0331  & \pi1076  ;
  assign n59355 = n11822 & n59354 ;
  assign n59356 = ~n12313 & n59355 ;
  assign n59357 = ~n59353 & ~n59356 ;
  assign n59358 = \pi0431  & ~n58898 ;
  assign n59359 = ~\pi0331  & \pi1071  ;
  assign n59360 = n11822 & n59359 ;
  assign n59361 = ~n12313 & n59360 ;
  assign n59362 = ~n59358 & ~n59361 ;
  assign n59363 = \pi0432  & ~n58898 ;
  assign n59364 = ~\pi0331  & \pi1068  ;
  assign n59365 = n11822 & n59364 ;
  assign n59366 = ~n12313 & n59365 ;
  assign n59367 = ~n59363 & ~n59366 ;
  assign n59368 = \pi0433  & ~n58898 ;
  assign n59369 = ~\pi0331  & \pi1042  ;
  assign n59370 = n11822 & n59369 ;
  assign n59371 = ~n12313 & n59370 ;
  assign n59372 = ~n59368 & ~n59371 ;
  assign n59373 = \pi0434  & ~n58898 ;
  assign n59374 = ~\pi0331  & \pi1059  ;
  assign n59375 = n11822 & n59374 ;
  assign n59376 = ~n12313 & n59375 ;
  assign n59377 = ~n59373 & ~n59376 ;
  assign n59378 = \pi0435  & ~n58898 ;
  assign n59379 = ~\pi0331  & \pi1053  ;
  assign n59380 = n11822 & n59379 ;
  assign n59381 = ~n12313 & n59380 ;
  assign n59382 = ~n59378 & ~n59381 ;
  assign n59383 = \pi0436  & ~n58898 ;
  assign n59384 = ~\pi0331  & \pi1037  ;
  assign n59385 = n11822 & n59384 ;
  assign n59386 = ~n12313 & n59385 ;
  assign n59387 = ~n59383 & ~n59386 ;
  assign n59388 = \pi0437  & ~n58898 ;
  assign n59389 = ~\pi0331  & \pi1070  ;
  assign n59390 = n11822 & n59389 ;
  assign n59391 = ~n12313 & n59390 ;
  assign n59392 = ~n59388 & ~n59391 ;
  assign n59393 = \pi0438  & ~n58898 ;
  assign n59394 = ~\pi0331  & \pi1036  ;
  assign n59395 = n11822 & n59394 ;
  assign n59396 = ~n12313 & n59395 ;
  assign n59397 = ~n59393 & ~n59396 ;
  assign n59398 = \pi0439  & ~n58759 ;
  assign n59399 = ~\pi0330  & \pi1057  ;
  assign n59400 = n11822 & n59399 ;
  assign n59401 = ~n12313 & n59400 ;
  assign n59402 = ~n59398 & ~n59401 ;
  assign n59403 = \pi0440  & ~n58759 ;
  assign n59404 = ~\pi0330  & \pi1043  ;
  assign n59405 = n11822 & n59404 ;
  assign n59406 = ~n12313 & n59405 ;
  assign n59407 = ~n59403 & ~n59406 ;
  assign n59408 = \pi0441  & ~n58747 ;
  assign n59409 = ~\pi0340  & \pi1044  ;
  assign n59410 = n11822 & n59409 ;
  assign n59411 = ~n12313 & n59410 ;
  assign n59412 = ~n59408 & ~n59411 ;
  assign n59413 = \pi0442  & ~n58759 ;
  assign n59414 = ~\pi0330  & \pi1058  ;
  assign n59415 = n11822 & n59414 ;
  assign n59416 = ~n12313 & n59415 ;
  assign n59417 = ~n59413 & ~n59416 ;
  assign n59418 = \pi0443  & ~n58898 ;
  assign n59419 = ~\pi0331  & \pi1044  ;
  assign n59420 = n11822 & n59419 ;
  assign n59421 = ~n12313 & n59420 ;
  assign n59422 = ~n59418 & ~n59421 ;
  assign n59423 = \pi0444  & ~n58898 ;
  assign n59424 = ~\pi0331  & \pi1072  ;
  assign n59425 = n11822 & n59424 ;
  assign n59426 = ~n12313 & n59425 ;
  assign n59427 = ~n59423 & ~n59426 ;
  assign n59428 = \pi0445  & ~n58898 ;
  assign n59429 = ~\pi0331  & \pi1081  ;
  assign n59430 = n11822 & n59429 ;
  assign n59431 = ~n12313 & n59430 ;
  assign n59432 = ~n59428 & ~n59431 ;
  assign n59433 = \pi0446  & ~n58898 ;
  assign n59434 = ~\pi0331  & \pi1086  ;
  assign n59435 = n11822 & n59434 ;
  assign n59436 = ~n12313 & n59435 ;
  assign n59437 = ~n59433 & ~n59436 ;
  assign n59438 = \pi0447  & ~n58759 ;
  assign n59439 = ~\pi0330  & \pi1040  ;
  assign n59440 = n11822 & n59439 ;
  assign n59441 = ~n12313 & n59440 ;
  assign n59442 = ~n59438 & ~n59441 ;
  assign n59443 = \pi0448  & ~n58898 ;
  assign n59444 = ~\pi0331  & \pi1074  ;
  assign n59445 = n11822 & n59444 ;
  assign n59446 = ~n12313 & n59445 ;
  assign n59447 = ~n59443 & ~n59446 ;
  assign n59448 = \pi0449  & ~n58898 ;
  assign n59449 = ~\pi0331  & \pi1057  ;
  assign n59450 = n11822 & n59449 ;
  assign n59451 = ~n12313 & n59450 ;
  assign n59452 = ~n59448 & ~n59451 ;
  assign n59453 = \pi0450  & ~n58747 ;
  assign n59454 = ~\pi0340  & \pi1036  ;
  assign n59455 = n11822 & n59454 ;
  assign n59456 = ~n12313 & n59455 ;
  assign n59457 = ~n59453 & ~n59456 ;
  assign n59458 = \pi0451  & ~n58898 ;
  assign n59459 = ~\pi0331  & \pi1063  ;
  assign n59460 = n11822 & n59459 ;
  assign n59461 = ~n12313 & n59460 ;
  assign n59462 = ~n59458 & ~n59461 ;
  assign n59463 = \pi0452  & ~n58747 ;
  assign n59464 = ~\pi0340  & \pi1053  ;
  assign n59465 = n11822 & n59464 ;
  assign n59466 = ~n12313 & n59465 ;
  assign n59467 = ~n59463 & ~n59466 ;
  assign n59468 = \pi0453  & ~n58898 ;
  assign n59469 = ~\pi0331  & \pi1040  ;
  assign n59470 = n11822 & n59469 ;
  assign n59471 = ~n12313 & n59470 ;
  assign n59472 = ~n59468 & ~n59471 ;
  assign n59473 = \pi0454  & ~n58898 ;
  assign n59474 = ~\pi0331  & \pi1043  ;
  assign n59475 = n11822 & n59474 ;
  assign n59476 = ~n12313 & n59475 ;
  assign n59477 = ~n59473 & ~n59476 ;
  assign n59478 = \pi0455  & ~n58747 ;
  assign n59479 = ~\pi0340  & \pi1037  ;
  assign n59480 = n11822 & n59479 ;
  assign n59481 = ~n12313 & n59480 ;
  assign n59482 = ~n59478 & ~n59481 ;
  assign n59483 = \pi0456  & ~n58766 ;
  assign n59484 = ~\pi0341  & \pi1044  ;
  assign n59485 = n11822 & n59484 ;
  assign n59486 = ~n12313 & n59485 ;
  assign n59487 = ~n59483 & ~n59486 ;
  assign n59488 = ~\pi0599  & \pi0810  ;
  assign n59489 = \pi0596  & \pi0815  ;
  assign n59490 = ~n59488 & n59489 ;
  assign n59491 = ~\pi0804  & \pi0815  ;
  assign n59492 = \pi0595  & ~n59491 ;
  assign n59493 = ~n59490 & n59492 ;
  assign n59494 = \pi0594  & \pi0600  ;
  assign n59495 = \pi0597  & \pi0601  ;
  assign n59496 = n59494 & n59495 ;
  assign n59497 = ~\pi0804  & ~\pi0810  ;
  assign n59498 = ~\pi0595  & ~n59497 ;
  assign n59499 = \pi0605  & ~n59498 ;
  assign n59500 = n59496 & n59499 ;
  assign n59501 = ~n59493 & n59500 ;
  assign n59502 = ~\pi0601  & ~n59497 ;
  assign n59503 = \pi0600  & ~\pi0810  ;
  assign n59504 = \pi0804  & ~n59503 ;
  assign n59505 = ~n59502 & ~n59504 ;
  assign n59506 = \pi0605  & ~\pi0815  ;
  assign n59507 = n59505 & n59506 ;
  assign n59508 = \pi0804  & ~\pi0815  ;
  assign n59509 = ~n59503 & n59508 ;
  assign n59510 = \pi0990  & n59494 ;
  assign n59511 = n59509 & n59510 ;
  assign n59512 = ~n59507 & ~n59511 ;
  assign n59513 = ~n59501 & n59512 ;
  assign n59514 = \pi0821  & ~n59513 ;
  assign n59515 = \pi0458  & ~n58747 ;
  assign n59516 = ~\pi0340  & \pi1072  ;
  assign n59517 = n11822 & n59516 ;
  assign n59518 = ~n12313 & n59517 ;
  assign n59519 = ~n59515 & ~n59518 ;
  assign n59520 = \pi0459  & ~n58898 ;
  assign n59521 = ~\pi0331  & \pi1058  ;
  assign n59522 = n11822 & n59521 ;
  assign n59523 = ~n12313 & n59522 ;
  assign n59524 = ~n59520 & ~n59523 ;
  assign n59525 = \pi0460  & ~n58747 ;
  assign n59526 = ~\pi0340  & \pi1086  ;
  assign n59527 = n11822 & n59526 ;
  assign n59528 = ~n12313 & n59527 ;
  assign n59529 = ~n59525 & ~n59528 ;
  assign n59530 = \pi0461  & ~n58747 ;
  assign n59531 = ~\pi0340  & \pi1057  ;
  assign n59532 = n11822 & n59531 ;
  assign n59533 = ~n12313 & n59532 ;
  assign n59534 = ~n59530 & ~n59533 ;
  assign n59535 = \pi0462  & ~n58747 ;
  assign n59536 = ~\pi0340  & \pi1074  ;
  assign n59537 = n11822 & n59536 ;
  assign n59538 = ~n12313 & n59537 ;
  assign n59539 = ~n59535 & ~n59538 ;
  assign n59540 = \pi0463  & ~n58766 ;
  assign n59541 = ~\pi0341  & \pi1070  ;
  assign n59542 = n11822 & n59541 ;
  assign n59543 = ~n12313 & n59542 ;
  assign n59544 = ~n59540 & ~n59543 ;
  assign n59545 = \pi0464  & ~n58898 ;
  assign n59546 = ~\pi0331  & \pi1065  ;
  assign n59547 = n11822 & n59546 ;
  assign n59548 = ~n12313 & n59547 ;
  assign n59549 = ~n59545 & ~n59548 ;
  assign n59550 = ~\pi0224  & ~\pi0299  ;
  assign n59551 = n58627 & n59550 ;
  assign n59552 = ~n13622 & ~n59551 ;
  assign n59553 = ~\pi0243  & \pi1157  ;
  assign n59554 = \pi0926  & n59553 ;
  assign n59555 = ~n59552 & n59554 ;
  assign n59556 = n9948 & ~n59555 ;
  assign n59557 = ~n13578 & ~n13582 ;
  assign n59558 = ~\pi0243  & ~n59557 ;
  assign n59559 = \pi0299  & n1295 ;
  assign n59560 = ~\pi0299  & n58627 ;
  assign n59561 = ~n59559 & ~n59560 ;
  assign n59562 = ~n59553 & ~n59561 ;
  assign n59563 = ~\pi1157  & ~n2256 ;
  assign n59564 = \pi0221  & ~\pi1157  ;
  assign n59565 = ~n1220 & n59564 ;
  assign n59566 = ~n59563 & ~n59565 ;
  assign n59567 = ~n6456 & ~n59566 ;
  assign n59568 = ~n59562 & ~n59567 ;
  assign n59569 = ~n6452 & ~n6456 ;
  assign n59570 = ~\pi0926  & ~n59569 ;
  assign n59571 = n59568 & ~n59570 ;
  assign n59572 = ~n59558 & ~n59571 ;
  assign n59573 = n59556 & ~n59572 ;
  assign n59574 = \pi0215  & \pi1157  ;
  assign n59575 = \pi0221  & \pi1157  ;
  assign n59576 = ~n1220 & n59575 ;
  assign n59577 = ~n59574 & ~n59576 ;
  assign n59578 = \pi0926  & n58636 ;
  assign n59579 = ~\pi0215  & ~\pi0243  ;
  assign n59580 = n2291 & n59579 ;
  assign n59581 = ~n59578 & ~n59580 ;
  assign n59582 = n59577 & n59581 ;
  assign n59583 = ~n55740 & ~n59582 ;
  assign n59584 = ~n59573 & ~n59583 ;
  assign n59585 = n9948 & ~n59561 ;
  assign n59586 = n1295 & ~n55740 ;
  assign n59587 = ~n59585 & ~n59586 ;
  assign n59588 = ~\pi0275  & ~n59587 ;
  assign n59589 = \pi0943  & \pi1151  ;
  assign n59590 = n2650 & n59589 ;
  assign n59591 = ~n20516 & n59590 ;
  assign n59592 = n2214 & n59589 ;
  assign n59593 = n20516 & n59592 ;
  assign n59594 = ~n59591 & ~n59593 ;
  assign n59595 = ~n59588 & n59594 ;
  assign n59596 = ~\pi0215  & n2291 ;
  assign n59597 = ~n55740 & ~n59596 ;
  assign n59598 = n55740 & n59557 ;
  assign n59599 = ~n59597 & ~n59598 ;
  assign n59600 = ~\pi0943  & ~\pi1151  ;
  assign n59601 = ~n59599 & n59600 ;
  assign n59602 = \pi0943  & ~\pi1151  ;
  assign n59603 = n58695 & n59602 ;
  assign n59604 = ~n59601 & ~n59603 ;
  assign n59605 = ~\pi0943  & ~n59599 ;
  assign n59606 = ~n58625 & n59605 ;
  assign n59607 = n59604 & ~n59606 ;
  assign n59608 = n59595 & n59607 ;
  assign n59609 = ~n6702 & n50325 ;
  assign n59610 = \pi0040  & \pi1001  ;
  assign n59611 = n55622 & n59610 ;
  assign n59612 = ~\pi0287  & n59611 ;
  assign n59613 = ~n59609 & n59612 ;
  assign n59614 = ~n11822 & ~n59613 ;
  assign n59615 = ~\pi0098  & ~n1535 ;
  assign n59616 = ~\pi0102  & ~n15845 ;
  assign n59617 = n13028 & n13426 ;
  assign n59618 = ~n59616 & n59617 ;
  assign n59619 = n59615 & n59618 ;
  assign n59620 = n59612 & ~n59619 ;
  assign n59621 = n13028 & ~n59612 ;
  assign n59622 = n13426 & n59621 ;
  assign n59623 = ~n59616 & n59622 ;
  assign n59624 = n59615 & n59623 ;
  assign n59625 = ~n8628 & ~n59624 ;
  assign n59626 = ~n59620 & n59625 ;
  assign n59627 = n8628 & ~n59619 ;
  assign n59628 = \pi1091  & ~n59627 ;
  assign n59629 = ~n59626 & n59628 ;
  assign n59630 = n2367 & n12970 ;
  assign n59631 = ~n59629 & n59630 ;
  assign n59632 = ~n59614 & ~n59631 ;
  assign n59633 = ~n9012 & ~n59624 ;
  assign n59634 = ~n59620 & n59633 ;
  assign n59635 = n9012 & ~n59619 ;
  assign n59636 = \pi1093  & ~n59635 ;
  assign n59637 = ~n59634 & n59636 ;
  assign n59638 = ~n6811 & ~n59624 ;
  assign n59639 = ~n59620 & n59638 ;
  assign n59640 = n6811 & ~n59619 ;
  assign n59641 = ~\pi1093  & ~n59640 ;
  assign n59642 = ~n59639 & n59641 ;
  assign n59643 = ~n59637 & ~n59642 ;
  assign n59644 = ~\pi1091  & n11822 ;
  assign n59645 = ~\pi1091  & n59612 ;
  assign n59646 = ~n59609 & n59645 ;
  assign n59647 = ~n59644 & ~n59646 ;
  assign n59648 = ~n59643 & ~n59647 ;
  assign n59649 = ~n59632 & ~n59648 ;
  assign n59650 = n13386 & n13493 ;
  assign n59651 = \pi0038  & ~\pi0057  ;
  assign n59652 = ~\pi0039  & n59651 ;
  assign n59653 = n6848 & n59652 ;
  assign n59654 = ~\pi0024  & n1289 ;
  assign n59655 = n1287 & n59654 ;
  assign n59656 = n59653 & n59655 ;
  assign n59657 = n1281 & n59656 ;
  assign n59658 = n1260 & n59657 ;
  assign n59659 = \pi0468  & ~n59658 ;
  assign n59660 = ~n59650 & ~n59659 ;
  assign n59661 = ~\pi0263  & \pi1156  ;
  assign n59662 = \pi0942  & n59661 ;
  assign n59663 = ~n59552 & n59662 ;
  assign n59664 = n9948 & ~n59663 ;
  assign n59665 = ~\pi0263  & ~n59557 ;
  assign n59666 = n59664 & n59665 ;
  assign n59667 = ~n59561 & ~n59661 ;
  assign n59668 = ~\pi1156  & n59569 ;
  assign n59669 = ~n59667 & ~n59668 ;
  assign n59670 = ~\pi0942  & ~n59569 ;
  assign n59671 = n59664 & ~n59670 ;
  assign n59672 = n59669 & n59671 ;
  assign n59673 = ~n59666 & ~n59672 ;
  assign n59674 = \pi0215  & \pi1156  ;
  assign n59675 = \pi0221  & \pi1156  ;
  assign n59676 = ~n1220 & n59675 ;
  assign n59677 = ~n59674 & ~n59676 ;
  assign n59678 = \pi0942  & n58636 ;
  assign n59679 = ~\pi0215  & ~\pi0263  ;
  assign n59680 = n2291 & n59679 ;
  assign n59681 = ~n59678 & ~n59680 ;
  assign n59682 = n59677 & n59681 ;
  assign n59683 = ~n55740 & ~n59682 ;
  assign n59684 = n59673 & ~n59683 ;
  assign n59685 = \pi0267  & \pi1155  ;
  assign n59686 = \pi0925  & n59685 ;
  assign n59687 = ~n59552 & n59686 ;
  assign n59688 = n9948 & ~n59687 ;
  assign n59689 = \pi0267  & ~n59557 ;
  assign n59690 = n59688 & n59689 ;
  assign n59691 = ~n59561 & ~n59685 ;
  assign n59692 = ~\pi1155  & n59569 ;
  assign n59693 = ~n59691 & ~n59692 ;
  assign n59694 = ~\pi0925  & ~n59569 ;
  assign n59695 = n59688 & ~n59694 ;
  assign n59696 = n59693 & n59695 ;
  assign n59697 = ~n59690 & ~n59696 ;
  assign n59698 = \pi0215  & \pi1155  ;
  assign n59699 = \pi0221  & \pi1155  ;
  assign n59700 = ~n1220 & n59699 ;
  assign n59701 = ~n59698 & ~n59700 ;
  assign n59702 = \pi0925  & n58636 ;
  assign n59703 = ~\pi0215  & \pi0267  ;
  assign n59704 = n2291 & n59703 ;
  assign n59705 = ~n59702 & ~n59704 ;
  assign n59706 = n59701 & n59705 ;
  assign n59707 = ~n55740 & ~n59706 ;
  assign n59708 = n59697 & ~n59707 ;
  assign n59709 = \pi0253  & \pi1153  ;
  assign n59710 = \pi0941  & n59709 ;
  assign n59711 = ~n59552 & n59710 ;
  assign n59712 = n9948 & ~n59711 ;
  assign n59713 = \pi0253  & ~n59557 ;
  assign n59714 = n59712 & n59713 ;
  assign n59715 = ~n59561 & ~n59709 ;
  assign n59716 = ~\pi1153  & n59569 ;
  assign n59717 = ~n59715 & ~n59716 ;
  assign n59718 = ~\pi0941  & ~n59569 ;
  assign n59719 = n59712 & ~n59718 ;
  assign n59720 = n59717 & n59719 ;
  assign n59721 = ~n59714 & ~n59720 ;
  assign n59722 = \pi0215  & \pi1153  ;
  assign n59723 = \pi0221  & \pi1153  ;
  assign n59724 = ~n1220 & n59723 ;
  assign n59725 = ~n59722 & ~n59724 ;
  assign n59726 = \pi0941  & n58636 ;
  assign n59727 = ~\pi0215  & \pi0253  ;
  assign n59728 = n2291 & n59727 ;
  assign n59729 = ~n59726 & ~n59728 ;
  assign n59730 = n59725 & n59729 ;
  assign n59731 = ~n55740 & ~n59730 ;
  assign n59732 = n59721 & ~n59731 ;
  assign n59733 = \pi0254  & \pi1154  ;
  assign n59734 = \pi0923  & n59733 ;
  assign n59735 = ~n59552 & n59734 ;
  assign n59736 = n9948 & ~n59735 ;
  assign n59737 = \pi0254  & ~n59557 ;
  assign n59738 = n59736 & n59737 ;
  assign n59739 = ~n59561 & ~n59733 ;
  assign n59740 = ~\pi1154  & n59569 ;
  assign n59741 = ~n59739 & ~n59740 ;
  assign n59742 = ~\pi0923  & ~n59569 ;
  assign n59743 = n59736 & ~n59742 ;
  assign n59744 = n59741 & n59743 ;
  assign n59745 = ~n59738 & ~n59744 ;
  assign n59746 = \pi0215  & \pi1154  ;
  assign n59747 = \pi0221  & \pi1154  ;
  assign n59748 = ~n1220 & n59747 ;
  assign n59749 = ~n59746 & ~n59748 ;
  assign n59750 = \pi0923  & n58636 ;
  assign n59751 = ~\pi0215  & \pi0254  ;
  assign n59752 = n2291 & n59751 ;
  assign n59753 = ~n59750 & ~n59752 ;
  assign n59754 = n59749 & n59753 ;
  assign n59755 = ~n55740 & ~n59754 ;
  assign n59756 = n59745 & ~n59755 ;
  assign n59757 = ~\pi0268  & ~n59587 ;
  assign n59758 = \pi0922  & \pi1152  ;
  assign n59759 = n2650 & n59758 ;
  assign n59760 = ~n20516 & n59759 ;
  assign n59761 = n2214 & n59758 ;
  assign n59762 = n20516 & n59761 ;
  assign n59763 = ~n59760 & ~n59762 ;
  assign n59764 = ~n59757 & n59763 ;
  assign n59765 = ~\pi0922  & ~\pi1152  ;
  assign n59766 = ~n59599 & n59765 ;
  assign n59767 = \pi0922  & ~\pi1152  ;
  assign n59768 = n58695 & n59767 ;
  assign n59769 = ~n59766 & ~n59768 ;
  assign n59770 = ~\pi0922  & ~n59599 ;
  assign n59771 = ~n58625 & n59770 ;
  assign n59772 = n59769 & ~n59771 ;
  assign n59773 = n59764 & n59772 ;
  assign n59774 = ~\pi0272  & ~n59587 ;
  assign n59775 = \pi0931  & \pi1150  ;
  assign n59776 = n2650 & n59775 ;
  assign n59777 = ~n20516 & n59776 ;
  assign n59778 = n2214 & n59775 ;
  assign n59779 = n20516 & n59778 ;
  assign n59780 = ~n59777 & ~n59779 ;
  assign n59781 = ~n59774 & n59780 ;
  assign n59782 = ~\pi0931  & ~\pi1150  ;
  assign n59783 = ~n59599 & n59782 ;
  assign n59784 = \pi0931  & ~\pi1150  ;
  assign n59785 = n58695 & n59784 ;
  assign n59786 = ~n59783 & ~n59785 ;
  assign n59787 = ~\pi0931  & ~n59599 ;
  assign n59788 = ~n58625 & n59787 ;
  assign n59789 = n59786 & ~n59788 ;
  assign n59790 = n59781 & n59789 ;
  assign n59791 = ~\pi0283  & ~n59587 ;
  assign n59792 = \pi0936  & \pi1149  ;
  assign n59793 = n2650 & n59792 ;
  assign n59794 = ~n20516 & n59793 ;
  assign n59795 = n2214 & n59792 ;
  assign n59796 = n20516 & n59795 ;
  assign n59797 = ~n59794 & ~n59796 ;
  assign n59798 = ~n59791 & n59797 ;
  assign n59799 = ~\pi0936  & ~\pi1149  ;
  assign n59800 = ~n59599 & n59799 ;
  assign n59801 = \pi0936  & ~\pi1149  ;
  assign n59802 = n58695 & n59801 ;
  assign n59803 = ~n59800 & ~n59802 ;
  assign n59804 = ~\pi0936  & ~n59599 ;
  assign n59805 = ~n58625 & n59804 ;
  assign n59806 = n59803 & ~n59805 ;
  assign n59807 = n59798 & n59806 ;
  assign n59808 = n13649 & n15334 ;
  assign n59809 = n11805 & ~n13649 ;
  assign n59810 = n13665 & n59809 ;
  assign n59811 = ~n59808 & ~n59810 ;
  assign n59812 = n1291 & n13042 ;
  assign n59813 = n15340 & n59812 ;
  assign n59814 = ~n59811 & n59813 ;
  assign n59815 = \pi0071  & n13647 ;
  assign n59816 = ~n55740 & n59815 ;
  assign n59817 = \pi0071  & ~\pi0299  ;
  assign n59818 = n13645 & n59817 ;
  assign n59819 = \pi0071  & \pi0299  ;
  assign n59820 = n13647 & n59819 ;
  assign n59821 = ~n59818 & ~n59820 ;
  assign n59822 = ~n59816 & n59821 ;
  assign n59823 = ~n59814 & n59822 ;
  assign n59824 = ~n55740 & ~n59816 ;
  assign n59825 = ~n59823 & ~n59824 ;
  assign n59826 = n11824 & ~n58721 ;
  assign n59827 = ~n58717 & n59826 ;
  assign n59828 = \pi0071  & ~n57606 ;
  assign n59829 = n11822 & ~n12313 ;
  assign n59830 = \pi0481  & ~n44552 ;
  assign n59831 = \pi0248  & n44495 ;
  assign n59832 = n44563 & n59831 ;
  assign n59833 = ~n44546 & n59832 ;
  assign n59834 = ~n59830 & ~n59833 ;
  assign n59835 = \pi0482  & ~n44585 ;
  assign n59836 = \pi0249  & n44573 ;
  assign n59837 = n44563 & n59836 ;
  assign n59838 = ~n44546 & n59837 ;
  assign n59839 = ~n59835 & ~n59838 ;
  assign n59840 = \pi0483  & ~n44789 ;
  assign n59841 = \pi0242  & n44782 ;
  assign n59842 = ~n44593 & n59841 ;
  assign n59843 = n44590 & n59842 ;
  assign n59844 = ~n59840 & ~n59843 ;
  assign n59845 = \pi0484  & ~n44789 ;
  assign n59846 = \pi0249  & n44782 ;
  assign n59847 = ~n44593 & n59846 ;
  assign n59848 = n44590 & n59847 ;
  assign n59849 = ~n59845 & ~n59848 ;
  assign n59850 = \pi0485  & ~n46731 ;
  assign n59851 = \pi0234  & n44573 ;
  assign n59852 = ~n44767 & n59851 ;
  assign n59853 = ~n59850 & ~n59852 ;
  assign n59854 = \pi0486  & ~n46731 ;
  assign n59855 = \pi0244  & n44573 ;
  assign n59856 = ~n44767 & n59855 ;
  assign n59857 = ~n59854 & ~n59856 ;
  assign n59858 = \pi0487  & ~n44552 ;
  assign n59859 = \pi0246  & n44495 ;
  assign n59860 = n44563 & n59859 ;
  assign n59861 = ~n44546 & n59860 ;
  assign n59862 = ~n59858 & ~n59861 ;
  assign n59863 = \pi0488  & ~n44552 ;
  assign n59864 = ~\pi0239  & n44495 ;
  assign n59865 = n44563 & n59864 ;
  assign n59866 = ~n44546 & n59865 ;
  assign n59867 = ~n59863 & ~n59866 ;
  assign n59868 = \pi0489  & ~n46731 ;
  assign n59869 = \pi0242  & n44573 ;
  assign n59870 = ~n44767 & n59869 ;
  assign n59871 = ~n59868 & ~n59870 ;
  assign n59872 = \pi0490  & ~n44789 ;
  assign n59873 = \pi0241  & n44782 ;
  assign n59874 = ~n44767 & n59873 ;
  assign n59875 = ~n59872 & ~n59874 ;
  assign n59876 = \pi0491  & ~n44789 ;
  assign n59877 = \pi0238  & n44782 ;
  assign n59878 = ~n44767 & n59877 ;
  assign n59879 = ~n59876 & ~n59878 ;
  assign n59880 = \pi0492  & ~n44789 ;
  assign n59881 = \pi0240  & n44782 ;
  assign n59882 = ~n44767 & n59881 ;
  assign n59883 = ~n59880 & ~n59882 ;
  assign n59884 = \pi0493  & ~n44789 ;
  assign n59885 = \pi0244  & n44782 ;
  assign n59886 = ~n44767 & n59885 ;
  assign n59887 = ~n59884 & ~n59886 ;
  assign n59888 = \pi0494  & ~n44789 ;
  assign n59889 = ~\pi0239  & n44782 ;
  assign n59890 = ~n44767 & n59889 ;
  assign n59891 = ~n59888 & ~n59890 ;
  assign n59892 = \pi0495  & ~n44789 ;
  assign n59893 = \pi0235  & n44782 ;
  assign n59894 = ~n44767 & n59893 ;
  assign n59895 = ~n59892 & ~n59894 ;
  assign n59896 = \pi0496  & ~n44774 ;
  assign n59897 = \pi0249  & n44556 ;
  assign n59898 = ~n44767 & n59897 ;
  assign n59899 = ~n59896 & ~n59898 ;
  assign n59900 = \pi0497  & ~n44774 ;
  assign n59901 = ~\pi0239  & n44556 ;
  assign n59902 = ~n44767 & n59901 ;
  assign n59903 = ~n59900 & ~n59902 ;
  assign n59904 = \pi0498  & ~n44585 ;
  assign n59905 = \pi0238  & n44573 ;
  assign n59906 = n44563 & n59905 ;
  assign n59907 = ~n44546 & n59906 ;
  assign n59908 = ~n59904 & ~n59907 ;
  assign n59909 = \pi0499  & ~n44774 ;
  assign n59910 = \pi0246  & n44556 ;
  assign n59911 = ~n44767 & n59910 ;
  assign n59912 = ~n59909 & ~n59911 ;
  assign n59913 = \pi0500  & ~n44774 ;
  assign n59914 = \pi0241  & n44556 ;
  assign n59915 = ~n44767 & n59914 ;
  assign n59916 = ~n59913 & ~n59915 ;
  assign n59917 = \pi0501  & ~n44774 ;
  assign n59918 = \pi0248  & n44556 ;
  assign n59919 = ~n44767 & n59918 ;
  assign n59920 = ~n59917 & ~n59919 ;
  assign n59921 = \pi0502  & ~n44774 ;
  assign n59922 = \pi0247  & n44556 ;
  assign n59923 = ~n44767 & n59922 ;
  assign n59924 = ~n59921 & ~n59923 ;
  assign n59925 = \pi0503  & ~n44774 ;
  assign n59926 = \pi0245  & n44556 ;
  assign n59927 = ~n44767 & n59926 ;
  assign n59928 = ~n59925 & ~n59927 ;
  assign n59929 = \pi0504  & ~n44714 ;
  assign n59930 = \pi0242  & n44495 ;
  assign n59931 = ~n44767 & n59930 ;
  assign n59932 = ~n59929 & ~n59931 ;
  assign n59933 = ~n7178 & n20516 ;
  assign n59934 = n44556 & ~n59933 ;
  assign n59935 = ~n44767 & n59934 ;
  assign n59936 = \pi0505  & ~n59935 ;
  assign n59937 = \pi0234  & n44556 ;
  assign n59938 = ~n44767 & n59937 ;
  assign n59939 = ~n59936 & ~n59938 ;
  assign n59940 = \pi0506  & ~n44714 ;
  assign n59941 = \pi0241  & n44495 ;
  assign n59942 = ~n44767 & n59941 ;
  assign n59943 = ~n59940 & ~n59942 ;
  assign n59944 = \pi0507  & ~n44714 ;
  assign n59945 = \pi0238  & n44495 ;
  assign n59946 = ~n44767 & n59945 ;
  assign n59947 = ~n59944 & ~n59946 ;
  assign n59948 = \pi0508  & ~n44714 ;
  assign n59949 = \pi0247  & n44495 ;
  assign n59950 = ~n44767 & n59949 ;
  assign n59951 = ~n59948 & ~n59950 ;
  assign n59952 = \pi0509  & ~n44714 ;
  assign n59953 = \pi0245  & n44495 ;
  assign n59954 = ~n44767 & n59953 ;
  assign n59955 = ~n59952 & ~n59954 ;
  assign n59956 = \pi0510  & ~n44552 ;
  assign n59957 = n44563 & n59930 ;
  assign n59958 = ~n44546 & n59957 ;
  assign n59959 = ~n59956 & ~n59958 ;
  assign n59960 = \pi0511  & ~n44552 ;
  assign n59961 = \pi0234  & n44495 ;
  assign n59962 = n44563 & n59961 ;
  assign n59963 = ~n44546 & n59962 ;
  assign n59964 = ~n59960 & ~n59963 ;
  assign n59965 = \pi0512  & ~n44552 ;
  assign n59966 = \pi0235  & n44495 ;
  assign n59967 = n44563 & n59966 ;
  assign n59968 = ~n44546 & n59967 ;
  assign n59969 = ~n59965 & ~n59968 ;
  assign n59970 = \pi0513  & ~n44552 ;
  assign n59971 = \pi0244  & n44495 ;
  assign n59972 = n44563 & n59971 ;
  assign n59973 = ~n44546 & n59972 ;
  assign n59974 = ~n59970 & ~n59973 ;
  assign n59975 = \pi0514  & ~n44552 ;
  assign n59976 = n44563 & n59953 ;
  assign n59977 = ~n44546 & n59976 ;
  assign n59978 = ~n59975 & ~n59977 ;
  assign n59979 = \pi0515  & ~n44552 ;
  assign n59980 = \pi0240  & n44495 ;
  assign n59981 = n44563 & n59980 ;
  assign n59982 = ~n44546 & n59981 ;
  assign n59983 = ~n59979 & ~n59982 ;
  assign n59984 = \pi0516  & ~n44552 ;
  assign n59985 = n44563 & n59949 ;
  assign n59986 = ~n44546 & n59985 ;
  assign n59987 = ~n59984 & ~n59986 ;
  assign n59988 = \pi0517  & ~n44552 ;
  assign n59989 = n44563 & n59945 ;
  assign n59990 = ~n44546 & n59989 ;
  assign n59991 = ~n59988 & ~n59990 ;
  assign n59992 = \pi0518  & ~n44569 ;
  assign n59993 = n44563 & n59937 ;
  assign n59994 = ~n44546 & n59993 ;
  assign n59995 = ~n59992 & ~n59994 ;
  assign n59996 = \pi0519  & ~n44569 ;
  assign n59997 = n44563 & n59901 ;
  assign n59998 = ~n44546 & n59997 ;
  assign n59999 = ~n59996 & ~n59998 ;
  assign n60000 = \pi0520  & ~n44569 ;
  assign n60001 = n44563 & n59910 ;
  assign n60002 = ~n44546 & n60001 ;
  assign n60003 = ~n60000 & ~n60002 ;
  assign n60004 = \pi0521  & ~n44569 ;
  assign n60005 = n44563 & n59918 ;
  assign n60006 = ~n44546 & n60005 ;
  assign n60007 = ~n60004 & ~n60006 ;
  assign n60008 = \pi0522  & ~n44569 ;
  assign n60009 = \pi0238  & n44556 ;
  assign n60010 = n44563 & n60009 ;
  assign n60011 = ~n44546 & n60010 ;
  assign n60012 = ~n60008 & ~n60011 ;
  assign n60013 = \pi0523  & ~n46793 ;
  assign n60014 = \pi0234  & n44782 ;
  assign n60015 = n44563 & n60014 ;
  assign n60016 = ~n44546 & n60015 ;
  assign n60017 = ~n60013 & ~n60016 ;
  assign n60018 = \pi0524  & ~n46793 ;
  assign n60019 = n44563 & n59889 ;
  assign n60020 = ~n44546 & n60019 ;
  assign n60021 = ~n60018 & ~n60020 ;
  assign n60022 = \pi0525  & ~n46793 ;
  assign n60023 = \pi0245  & n44782 ;
  assign n60024 = n44563 & n60023 ;
  assign n60025 = ~n44546 & n60024 ;
  assign n60026 = ~n60022 & ~n60025 ;
  assign n60027 = \pi0526  & ~n46793 ;
  assign n60028 = \pi0246  & n44782 ;
  assign n60029 = n44563 & n60028 ;
  assign n60030 = ~n44546 & n60029 ;
  assign n60031 = ~n60027 & ~n60030 ;
  assign n60032 = \pi0527  & ~n46793 ;
  assign n60033 = \pi0247  & n44782 ;
  assign n60034 = n44563 & n60033 ;
  assign n60035 = ~n44546 & n60034 ;
  assign n60036 = ~n60032 & ~n60035 ;
  assign n60037 = \pi0528  & ~n46793 ;
  assign n60038 = n44563 & n59846 ;
  assign n60039 = ~n44546 & n60038 ;
  assign n60040 = ~n60037 & ~n60039 ;
  assign n60041 = \pi0529  & ~n46793 ;
  assign n60042 = n44563 & n59877 ;
  assign n60043 = ~n44546 & n60042 ;
  assign n60044 = ~n60041 & ~n60043 ;
  assign n60045 = \pi0530  & ~n46793 ;
  assign n60046 = n44563 & n59881 ;
  assign n60047 = ~n44546 & n60046 ;
  assign n60048 = ~n60045 & ~n60047 ;
  assign n60049 = \pi0531  & ~n44585 ;
  assign n60050 = \pi0235  & n44573 ;
  assign n60051 = n44563 & n60050 ;
  assign n60052 = ~n44546 & n60051 ;
  assign n60053 = ~n60049 & ~n60052 ;
  assign n60054 = \pi0532  & ~n44585 ;
  assign n60055 = \pi0247  & n44573 ;
  assign n60056 = n44563 & n60055 ;
  assign n60057 = ~n44546 & n60056 ;
  assign n60058 = ~n60054 & ~n60057 ;
  assign n60059 = \pi0533  & ~n44714 ;
  assign n60060 = ~n44767 & n59966 ;
  assign n60061 = ~n60059 & ~n60060 ;
  assign n60062 = \pi0534  & ~n44714 ;
  assign n60063 = ~n44767 & n59864 ;
  assign n60064 = ~n60062 & ~n60063 ;
  assign n60065 = \pi0535  & ~n44714 ;
  assign n60066 = ~n44767 & n59980 ;
  assign n60067 = ~n60065 & ~n60066 ;
  assign n60068 = \pi0536  & ~n44714 ;
  assign n60069 = ~n44767 & n59859 ;
  assign n60070 = ~n60068 & ~n60069 ;
  assign n60071 = \pi0537  & ~n44714 ;
  assign n60072 = ~n44767 & n59831 ;
  assign n60073 = ~n60071 & ~n60072 ;
  assign n60074 = \pi0538  & ~n44714 ;
  assign n60075 = \pi0249  & n44495 ;
  assign n60076 = ~n44767 & n60075 ;
  assign n60077 = ~n60074 & ~n60076 ;
  assign n60078 = \pi0539  & ~n44774 ;
  assign n60079 = \pi0242  & n44556 ;
  assign n60080 = ~n44767 & n60079 ;
  assign n60081 = ~n60078 & ~n60080 ;
  assign n60082 = \pi0540  & ~n44774 ;
  assign n60083 = \pi0235  & n44556 ;
  assign n60084 = ~n44767 & n60083 ;
  assign n60085 = ~n60082 & ~n60084 ;
  assign n60086 = \pi0541  & ~n44774 ;
  assign n60087 = \pi0244  & n44556 ;
  assign n60088 = ~n44767 & n60087 ;
  assign n60089 = ~n60086 & ~n60088 ;
  assign n60090 = \pi0542  & ~n44774 ;
  assign n60091 = \pi0240  & n44556 ;
  assign n60092 = ~n44767 & n60091 ;
  assign n60093 = ~n60090 & ~n60092 ;
  assign n60094 = \pi0543  & ~n44774 ;
  assign n60095 = ~n44767 & n60009 ;
  assign n60096 = ~n60094 & ~n60095 ;
  assign n60097 = n44782 & ~n59933 ;
  assign n60098 = ~n44767 & n60097 ;
  assign n60099 = \pi0544  & ~n60098 ;
  assign n60100 = ~n44767 & n60014 ;
  assign n60101 = ~n60099 & ~n60100 ;
  assign n60102 = \pi0545  & ~n44789 ;
  assign n60103 = ~n44767 & n60023 ;
  assign n60104 = ~n60102 & ~n60103 ;
  assign n60105 = \pi0546  & ~n44789 ;
  assign n60106 = ~n44767 & n60028 ;
  assign n60107 = ~n60105 & ~n60106 ;
  assign n60108 = \pi0547  & ~n44789 ;
  assign n60109 = ~n44767 & n60033 ;
  assign n60110 = ~n60108 & ~n60109 ;
  assign n60111 = \pi0548  & ~n44789 ;
  assign n60112 = \pi0248  & n44782 ;
  assign n60113 = ~n44767 & n60112 ;
  assign n60114 = ~n60111 & ~n60113 ;
  assign n60115 = \pi0549  & ~n46731 ;
  assign n60116 = ~n44767 & n60050 ;
  assign n60117 = ~n60115 & ~n60116 ;
  assign n60118 = \pi0550  & ~n46731 ;
  assign n60119 = ~\pi0239  & n44573 ;
  assign n60120 = ~n44767 & n60119 ;
  assign n60121 = ~n60118 & ~n60120 ;
  assign n60122 = \pi0551  & ~n46731 ;
  assign n60123 = \pi0240  & n44573 ;
  assign n60124 = ~n44767 & n60123 ;
  assign n60125 = ~n60122 & ~n60124 ;
  assign n60126 = \pi0552  & ~n46731 ;
  assign n60127 = ~n44767 & n60055 ;
  assign n60128 = ~n60126 & ~n60127 ;
  assign n60129 = \pi0553  & ~n46731 ;
  assign n60130 = \pi0241  & n44573 ;
  assign n60131 = ~n44767 & n60130 ;
  assign n60132 = ~n60129 & ~n60131 ;
  assign n60133 = \pi0554  & ~n46731 ;
  assign n60134 = \pi0248  & n44573 ;
  assign n60135 = ~n44767 & n60134 ;
  assign n60136 = ~n60133 & ~n60135 ;
  assign n60137 = \pi0555  & ~n46731 ;
  assign n60138 = ~n44767 & n59836 ;
  assign n60139 = ~n60137 & ~n60138 ;
  assign n60140 = \pi0556  & ~n44585 ;
  assign n60141 = n44563 & n59869 ;
  assign n60142 = ~n44546 & n60141 ;
  assign n60143 = ~n60140 & ~n60142 ;
  assign n60144 = n44714 & ~n59933 ;
  assign n60145 = \pi0557  & ~n60144 ;
  assign n60146 = ~n44767 & n59961 ;
  assign n60147 = ~n60145 & ~n60146 ;
  assign n60148 = \pi0558  & ~n44714 ;
  assign n60149 = ~n44767 & n59971 ;
  assign n60150 = ~n60148 & ~n60149 ;
  assign n60151 = \pi0559  & ~n44552 ;
  assign n60152 = n44563 & n59941 ;
  assign n60153 = ~n44546 & n60152 ;
  assign n60154 = ~n60151 & ~n60153 ;
  assign n60155 = \pi0560  & ~n44585 ;
  assign n60156 = n44563 & n60123 ;
  assign n60157 = ~n44546 & n60156 ;
  assign n60158 = ~n60155 & ~n60157 ;
  assign n60159 = \pi0561  & ~n44569 ;
  assign n60160 = n44563 & n59922 ;
  assign n60161 = ~n44546 & n60160 ;
  assign n60162 = ~n60159 & ~n60161 ;
  assign n60163 = \pi0562  & ~n44585 ;
  assign n60164 = n44563 & n60130 ;
  assign n60165 = ~n44546 & n60164 ;
  assign n60166 = ~n60163 & ~n60165 ;
  assign n60167 = \pi0563  & ~n46731 ;
  assign n60168 = \pi0246  & n44573 ;
  assign n60169 = ~n44767 & n60168 ;
  assign n60170 = ~n60167 & ~n60169 ;
  assign n60171 = \pi0564  & ~n44585 ;
  assign n60172 = n44563 & n60168 ;
  assign n60173 = ~n44546 & n60172 ;
  assign n60174 = ~n60171 & ~n60173 ;
  assign n60175 = \pi0565  & ~n44585 ;
  assign n60176 = n44563 & n60134 ;
  assign n60177 = ~n44546 & n60176 ;
  assign n60178 = ~n60175 & ~n60177 ;
  assign n60179 = \pi0566  & ~n44585 ;
  assign n60180 = n44563 & n59855 ;
  assign n60181 = ~n44546 & n60180 ;
  assign n60182 = ~n60179 & ~n60181 ;
  assign n60183 = ~\pi0567  & \pi1092  ;
  assign n60184 = ~\pi0230  & ~n60183 ;
  assign n60185 = \pi0603  & n1689 ;
  assign n60186 = n20783 & n60185 ;
  assign n60187 = ~n23880 & n60186 ;
  assign n60188 = ~n20846 & n60187 ;
  assign n60189 = n23832 & n60188 ;
  assign n60190 = ~\pi1093  & n60183 ;
  assign n60191 = \pi1157  & ~n60190 ;
  assign n60192 = ~n60189 & n60191 ;
  assign n60193 = ~n20925 & ~n60192 ;
  assign n60194 = ~\pi1157  & ~n60190 ;
  assign n60195 = \pi0630  & ~n60194 ;
  assign n60196 = \pi0680  & n1689 ;
  assign n60197 = n20854 & n60196 ;
  assign n60198 = ~n20861 & n60197 ;
  assign n60199 = ~n60190 & ~n60198 ;
  assign n60200 = n23885 & ~n60199 ;
  assign n60201 = n23921 & n60200 ;
  assign n60202 = ~n60195 & ~n60201 ;
  assign n60203 = n60193 & ~n60202 ;
  assign n60204 = ~n60189 & n60194 ;
  assign n60205 = ~n22945 & ~n60204 ;
  assign n60206 = ~\pi0630  & ~n60191 ;
  assign n60207 = ~\pi0630  & n23908 ;
  assign n60208 = n60200 & n60207 ;
  assign n60209 = ~n60206 & ~n60208 ;
  assign n60210 = n60205 & ~n60209 ;
  assign n60211 = ~n60203 & ~n60210 ;
  assign n60212 = n32298 & ~n60211 ;
  assign n60213 = n42957 & n60200 ;
  assign n60214 = \pi0629  & n20783 ;
  assign n60215 = n60185 & n60214 ;
  assign n60216 = ~n23880 & n60215 ;
  assign n60217 = \pi1156  & n60216 ;
  assign n60218 = n23832 & n60217 ;
  assign n60219 = ~n60213 & ~n60218 ;
  assign n60220 = n23832 & n60187 ;
  assign n60221 = ~n60200 & ~n60220 ;
  assign n60222 = ~\pi0792  & ~n60221 ;
  assign n60223 = n42949 & n60200 ;
  assign n60224 = ~\pi0629  & n20783 ;
  assign n60225 = n60185 & n60224 ;
  assign n60226 = ~n23880 & n60225 ;
  assign n60227 = n23831 & n60226 ;
  assign n60228 = ~\pi1156  & n21777 ;
  assign n60229 = n60227 & n60228 ;
  assign n60230 = ~n60190 & ~n60229 ;
  assign n60231 = ~n60223 & n60230 ;
  assign n60232 = ~n60222 & n60231 ;
  assign n60233 = n60219 & n60232 ;
  assign n60234 = n30712 & ~n60194 ;
  assign n60235 = ~\pi0630  & ~\pi0647  ;
  assign n60236 = \pi0787  & ~n60235 ;
  assign n60237 = n24994 & ~n60190 ;
  assign n60238 = ~n60236 & ~n60237 ;
  assign n60239 = ~n60234 & ~n60238 ;
  assign n60240 = ~n24761 & ~n60239 ;
  assign n60241 = ~n60233 & n60240 ;
  assign n60242 = \pi0230  & ~\pi0790  ;
  assign n60243 = n26069 & n60200 ;
  assign n60244 = n26080 & n60190 ;
  assign n60245 = n23412 & n26080 ;
  assign n60246 = n21092 & n60245 ;
  assign n60247 = n60220 & n60246 ;
  assign n60248 = ~n60244 & ~n60247 ;
  assign n60249 = n47917 & n60220 ;
  assign n60250 = ~\pi0644  & ~n23316 ;
  assign n60251 = n60190 & n60250 ;
  assign n60252 = \pi0230  & ~n60251 ;
  assign n60253 = ~n60249 & n60252 ;
  assign n60254 = n60248 & n60253 ;
  assign n60255 = ~n60243 & n60254 ;
  assign n60256 = ~n60242 & ~n60255 ;
  assign n60257 = ~n60241 & ~n60256 ;
  assign n60258 = ~n60212 & n60257 ;
  assign n60259 = ~n60184 & ~n60258 ;
  assign n60260 = \pi0568  & ~n44585 ;
  assign n60261 = \pi0245  & n44573 ;
  assign n60262 = n44563 & n60261 ;
  assign n60263 = ~n44546 & n60262 ;
  assign n60264 = ~n60260 & ~n60263 ;
  assign n60265 = \pi0569  & ~n44585 ;
  assign n60266 = n44563 & n60119 ;
  assign n60267 = ~n44546 & n60266 ;
  assign n60268 = ~n60265 & ~n60267 ;
  assign n60269 = \pi0570  & ~n44585 ;
  assign n60270 = n44563 & n59851 ;
  assign n60271 = ~n44546 & n60270 ;
  assign n60272 = ~n60269 & ~n60271 ;
  assign n60273 = \pi0571  & ~n46793 ;
  assign n60274 = n44563 & n59873 ;
  assign n60275 = ~n44546 & n60274 ;
  assign n60276 = ~n60273 & ~n60275 ;
  assign n60277 = \pi0572  & ~n46793 ;
  assign n60278 = n44563 & n59885 ;
  assign n60279 = ~n44546 & n60278 ;
  assign n60280 = ~n60277 & ~n60279 ;
  assign n60281 = \pi0573  & ~n46793 ;
  assign n60282 = n44563 & n59841 ;
  assign n60283 = ~n44546 & n60282 ;
  assign n60284 = ~n60281 & ~n60283 ;
  assign n60285 = \pi0574  & ~n44569 ;
  assign n60286 = n44563 & n59914 ;
  assign n60287 = ~n44546 & n60286 ;
  assign n60288 = ~n60285 & ~n60287 ;
  assign n60289 = \pi0575  & ~n46793 ;
  assign n60290 = n44563 & n59893 ;
  assign n60291 = ~n44546 & n60290 ;
  assign n60292 = ~n60289 & ~n60291 ;
  assign n60293 = \pi0576  & ~n46793 ;
  assign n60294 = n44563 & n60112 ;
  assign n60295 = ~n44546 & n60294 ;
  assign n60296 = ~n60293 & ~n60295 ;
  assign n60297 = \pi0577  & ~n46731 ;
  assign n60298 = ~n44767 & n59905 ;
  assign n60299 = ~n60297 & ~n60298 ;
  assign n60300 = \pi0578  & ~n44569 ;
  assign n60301 = n44563 & n59897 ;
  assign n60302 = ~n44546 & n60301 ;
  assign n60303 = ~n60300 & ~n60302 ;
  assign n60304 = \pi0579  & ~n44552 ;
  assign n60305 = n44563 & n60075 ;
  assign n60306 = ~n44546 & n60305 ;
  assign n60307 = ~n60304 & ~n60306 ;
  assign n60308 = \pi0580  & ~n46731 ;
  assign n60309 = ~n44767 & n60261 ;
  assign n60310 = ~n60308 & ~n60309 ;
  assign n60311 = \pi0581  & ~n44569 ;
  assign n60312 = n44563 & n60083 ;
  assign n60313 = ~n44546 & n60312 ;
  assign n60314 = ~n60311 & ~n60313 ;
  assign n60315 = \pi0582  & ~n44569 ;
  assign n60316 = n44563 & n60091 ;
  assign n60317 = ~n44546 & n60316 ;
  assign n60318 = ~n60315 & ~n60317 ;
  assign n60319 = \pi0584  & ~n44569 ;
  assign n60320 = n44563 & n59926 ;
  assign n60321 = ~n44546 & n60320 ;
  assign n60322 = ~n60319 & ~n60321 ;
  assign n60323 = \pi0585  & ~n44569 ;
  assign n60324 = n44563 & n60087 ;
  assign n60325 = ~n44546 & n60324 ;
  assign n60326 = ~n60323 & ~n60325 ;
  assign n60327 = \pi0586  & ~n44569 ;
  assign n60328 = n44563 & n60079 ;
  assign n60329 = ~n44546 & n60328 ;
  assign n60330 = ~n60327 & ~n60329 ;
  assign n60331 = ~\pi0230  & \pi0587  ;
  assign n60332 = \pi0230  & \pi0603  ;
  assign n60333 = ~n20783 & n60332 ;
  assign n60334 = n23832 & n60333 ;
  assign n60335 = n45843 & n60334 ;
  assign n60336 = ~n60331 & ~n60335 ;
  assign n60337 = ~\pi0123  & n14707 ;
  assign n60338 = ~\pi0588  & ~n60337 ;
  assign n60339 = ~\pi0123  & ~\pi0591  ;
  assign n60340 = n14707 & n60339 ;
  assign n60341 = n58904 & ~n60340 ;
  assign n60342 = ~n60338 & n60341 ;
  assign n60343 = ~\pi0205  & n20516 ;
  assign n60344 = ~\pi0205  & ~n6852 ;
  assign n60345 = ~n6851 & n60344 ;
  assign n60346 = ~n60343 & ~n60345 ;
  assign n60347 = ~n59933 & ~n60346 ;
  assign n60348 = ~\pi0202  & ~n20516 ;
  assign n60349 = n7284 & n60348 ;
  assign n60350 = ~\pi0202  & n20515 ;
  assign n60351 = n6848 & n60350 ;
  assign n60352 = n7343 & n60351 ;
  assign n60353 = ~\pi0233  & ~n60352 ;
  assign n60354 = ~n60349 & n60353 ;
  assign n60355 = ~n60347 & n60354 ;
  assign n60356 = ~\pi0204  & n20516 ;
  assign n60357 = ~\pi0204  & ~n6852 ;
  assign n60358 = ~n6851 & n60357 ;
  assign n60359 = ~n60356 & ~n60358 ;
  assign n60360 = ~n59933 & ~n60359 ;
  assign n60361 = ~\pi0201  & ~n20516 ;
  assign n60362 = n7284 & n60361 ;
  assign n60363 = ~\pi0201  & n20515 ;
  assign n60364 = n6848 & n60363 ;
  assign n60365 = n7343 & n60364 ;
  assign n60366 = \pi0233  & ~n60365 ;
  assign n60367 = ~n60362 & n60366 ;
  assign n60368 = ~n60360 & n60367 ;
  assign n60369 = ~n60355 & ~n60368 ;
  assign n60370 = \pi0237  & ~n60369 ;
  assign n60371 = ~\pi0218  & n20516 ;
  assign n60372 = ~\pi0218  & ~n6852 ;
  assign n60373 = ~n6851 & n60372 ;
  assign n60374 = ~n60371 & ~n60373 ;
  assign n60375 = ~n59933 & ~n60374 ;
  assign n60376 = ~\pi0203  & ~n20516 ;
  assign n60377 = n7284 & n60376 ;
  assign n60378 = ~\pi0203  & n20515 ;
  assign n60379 = n6848 & n60378 ;
  assign n60380 = n7343 & n60379 ;
  assign n60381 = ~\pi0233  & ~n60380 ;
  assign n60382 = ~n60377 & n60381 ;
  assign n60383 = ~n60375 & n60382 ;
  assign n60384 = ~\pi0206  & n20516 ;
  assign n60385 = ~\pi0206  & ~n6852 ;
  assign n60386 = ~n6851 & n60385 ;
  assign n60387 = ~n60384 & ~n60386 ;
  assign n60388 = ~n59933 & ~n60387 ;
  assign n60389 = ~\pi0220  & ~n20516 ;
  assign n60390 = n7284 & n60389 ;
  assign n60391 = ~\pi0220  & n20515 ;
  assign n60392 = n6848 & n60391 ;
  assign n60393 = n7343 & n60392 ;
  assign n60394 = \pi0233  & ~n60393 ;
  assign n60395 = ~n60390 & n60394 ;
  assign n60396 = ~n60388 & n60395 ;
  assign n60397 = ~n60383 & ~n60396 ;
  assign n60398 = ~\pi0237  & ~n60397 ;
  assign n60399 = ~n60370 & ~n60398 ;
  assign n60400 = \pi0590  & ~n60337 ;
  assign n60401 = ~\pi0123  & \pi0588  ;
  assign n60402 = n14707 & n60401 ;
  assign n60403 = n58904 & ~n60402 ;
  assign n60404 = ~n60400 & n60403 ;
  assign n60405 = ~\pi0591  & ~n60337 ;
  assign n60406 = ~\pi0123  & ~\pi0592  ;
  assign n60407 = n14707 & n60406 ;
  assign n60408 = n58904 & ~n60407 ;
  assign n60409 = ~n60405 & n60408 ;
  assign n60410 = ~\pi0592  & ~n60337 ;
  assign n60411 = ~\pi0123  & ~\pi0590  ;
  assign n60412 = n14707 & n60411 ;
  assign n60413 = n58904 & ~n60412 ;
  assign n60414 = ~n60410 & n60413 ;
  assign n60415 = ~\pi0234  & n20516 ;
  assign n60416 = ~\pi0234  & ~n6852 ;
  assign n60417 = ~n6851 & n60416 ;
  assign n60418 = ~n60415 & ~n60417 ;
  assign n60419 = ~n59933 & ~n60418 ;
  assign n60420 = ~\pi0249  & \pi0538  ;
  assign n60421 = \pi0248  & ~\pi0537  ;
  assign n60422 = ~\pi0248  & \pi0537  ;
  assign n60423 = ~n60421 & ~n60422 ;
  assign n60424 = ~n60420 & n60423 ;
  assign n60425 = ~\pi0246  & ~\pi0536  ;
  assign n60426 = \pi0246  & \pi0536  ;
  assign n60427 = ~n60425 & ~n60426 ;
  assign n60428 = \pi0249  & ~\pi0538  ;
  assign n60429 = ~\pi0557  & ~n60428 ;
  assign n60430 = ~n60427 & n60429 ;
  assign n60431 = n60424 & n60430 ;
  assign n60432 = n60419 & n60431 ;
  assign n60433 = \pi0234  & n20516 ;
  assign n60434 = \pi0234  & ~n6852 ;
  assign n60435 = ~n6851 & n60434 ;
  assign n60436 = ~n60433 & ~n60435 ;
  assign n60437 = ~n59933 & ~n60436 ;
  assign n60438 = \pi0557  & ~n60428 ;
  assign n60439 = ~n60427 & n60438 ;
  assign n60440 = n60424 & n60439 ;
  assign n60441 = n60437 & n60440 ;
  assign n60442 = ~n60432 & ~n60441 ;
  assign n60443 = ~\pi0241  & ~\pi0506  ;
  assign n60444 = \pi0241  & \pi0506  ;
  assign n60445 = ~n60443 & ~n60444 ;
  assign n60446 = ~\pi0534  & ~n60445 ;
  assign n60447 = ~\pi0240  & ~\pi0535  ;
  assign n60448 = \pi0240  & \pi0535  ;
  assign n60449 = ~n60447 & ~n60448 ;
  assign n60450 = \pi0239  & ~\pi0504  ;
  assign n60451 = ~n60449 & n60450 ;
  assign n60452 = n60446 & n60451 ;
  assign n60453 = ~n60442 & n60452 ;
  assign n60454 = \pi0534  & ~n60445 ;
  assign n60455 = ~\pi0239  & ~\pi0504  ;
  assign n60456 = ~n60449 & n60455 ;
  assign n60457 = n60454 & n60456 ;
  assign n60458 = ~n60442 & n60457 ;
  assign n60459 = ~n60453 & ~n60458 ;
  assign n60460 = ~\pi0242  & ~\pi0533  ;
  assign n60461 = ~n60459 & n60460 ;
  assign n60462 = \pi0239  & \pi0504  ;
  assign n60463 = ~n60449 & n60462 ;
  assign n60464 = n60446 & n60463 ;
  assign n60465 = ~n60442 & n60464 ;
  assign n60466 = ~\pi0239  & \pi0504  ;
  assign n60467 = ~n60449 & n60466 ;
  assign n60468 = n60454 & n60467 ;
  assign n60469 = ~n60442 & n60468 ;
  assign n60470 = ~n60465 & ~n60469 ;
  assign n60471 = \pi0242  & ~\pi0533  ;
  assign n60472 = ~n60470 & n60471 ;
  assign n60473 = ~n60461 & ~n60472 ;
  assign n60474 = ~\pi0235  & ~\pi0558  ;
  assign n60475 = ~n60473 & n60474 ;
  assign n60476 = ~\pi0242  & \pi0533  ;
  assign n60477 = ~n60459 & n60476 ;
  assign n60478 = \pi0242  & \pi0533  ;
  assign n60479 = ~n60470 & n60478 ;
  assign n60480 = ~n60477 & ~n60479 ;
  assign n60481 = \pi0235  & ~\pi0558  ;
  assign n60482 = ~n60480 & n60481 ;
  assign n60483 = ~n60475 & ~n60482 ;
  assign n60484 = ~\pi0244  & \pi0509  ;
  assign n60485 = ~n60483 & n60484 ;
  assign n60486 = ~\pi0235  & \pi0558  ;
  assign n60487 = ~n60473 & n60486 ;
  assign n60488 = \pi0235  & \pi0558  ;
  assign n60489 = ~n60480 & n60488 ;
  assign n60490 = ~n60487 & ~n60489 ;
  assign n60491 = \pi0244  & \pi0509  ;
  assign n60492 = ~n60490 & n60491 ;
  assign n60493 = ~n60485 & ~n60492 ;
  assign n60494 = \pi0245  & \pi0508  ;
  assign n60495 = ~n60493 & n60494 ;
  assign n60496 = ~\pi0244  & ~\pi0509  ;
  assign n60497 = ~n60483 & n60496 ;
  assign n60498 = \pi0244  & ~\pi0509  ;
  assign n60499 = ~n60490 & n60498 ;
  assign n60500 = ~n60497 & ~n60499 ;
  assign n60501 = ~\pi0245  & \pi0508  ;
  assign n60502 = ~n60500 & n60501 ;
  assign n60503 = ~n60495 & ~n60502 ;
  assign n60504 = \pi0247  & n60503 ;
  assign n60505 = ~\pi0234  & ~n20516 ;
  assign n60506 = n7284 & n60505 ;
  assign n60507 = n7343 & n60415 ;
  assign n60508 = ~n60506 & ~n60507 ;
  assign n60509 = ~\pi0249  & \pi0579  ;
  assign n60510 = \pi0246  & ~\pi0487  ;
  assign n60511 = ~\pi0246  & \pi0487  ;
  assign n60512 = ~n60510 & ~n60511 ;
  assign n60513 = ~n60509 & n60512 ;
  assign n60514 = ~\pi0248  & ~\pi0481  ;
  assign n60515 = \pi0248  & \pi0481  ;
  assign n60516 = ~n60514 & ~n60515 ;
  assign n60517 = \pi0249  & ~\pi0579  ;
  assign n60518 = ~\pi0511  & ~n60517 ;
  assign n60519 = ~n60516 & n60518 ;
  assign n60520 = n60513 & n60519 ;
  assign n60521 = ~n60508 & n60520 ;
  assign n60522 = \pi0234  & ~n20516 ;
  assign n60523 = n7284 & n60522 ;
  assign n60524 = n7343 & n60433 ;
  assign n60525 = ~n60523 & ~n60524 ;
  assign n60526 = \pi0511  & ~n60517 ;
  assign n60527 = ~n60516 & n60526 ;
  assign n60528 = n60513 & n60527 ;
  assign n60529 = ~n60525 & n60528 ;
  assign n60530 = ~n60521 & ~n60529 ;
  assign n60531 = ~\pi0241  & ~\pi0559  ;
  assign n60532 = ~\pi0515  & n60531 ;
  assign n60533 = \pi0241  & \pi0559  ;
  assign n60534 = ~\pi0515  & n60533 ;
  assign n60535 = ~n60532 & ~n60534 ;
  assign n60536 = ~n60530 & ~n60535 ;
  assign n60537 = \pi0239  & ~\pi0488  ;
  assign n60538 = ~\pi0239  & \pi0488  ;
  assign n60539 = ~n60537 & ~n60538 ;
  assign n60540 = ~\pi0240  & ~n60539 ;
  assign n60541 = n60536 & n60540 ;
  assign n60542 = \pi0515  & n60531 ;
  assign n60543 = \pi0515  & n60533 ;
  assign n60544 = ~n60542 & ~n60543 ;
  assign n60545 = ~n60530 & ~n60544 ;
  assign n60546 = \pi0240  & ~n60539 ;
  assign n60547 = n60545 & n60546 ;
  assign n60548 = ~n60541 & ~n60547 ;
  assign n60549 = ~\pi0235  & ~\pi0512  ;
  assign n60550 = \pi0235  & \pi0512  ;
  assign n60551 = ~n60549 & ~n60550 ;
  assign n60552 = ~\pi0242  & ~\pi0510  ;
  assign n60553 = \pi0242  & \pi0510  ;
  assign n60554 = ~n60552 & ~n60553 ;
  assign n60555 = ~\pi0244  & ~\pi0513  ;
  assign n60556 = \pi0244  & \pi0513  ;
  assign n60557 = ~n60555 & ~n60556 ;
  assign n60558 = ~n60554 & ~n60557 ;
  assign n60559 = ~n60551 & n60558 ;
  assign n60560 = ~\pi0245  & ~\pi0514  ;
  assign n60561 = \pi0245  & \pi0514  ;
  assign n60562 = ~n60560 & ~n60561 ;
  assign n60563 = \pi0508  & ~n60562 ;
  assign n60564 = n60559 & n60563 ;
  assign n60565 = ~n60548 & n60564 ;
  assign n60566 = ~\pi0247  & ~n60565 ;
  assign n60567 = ~n60504 & ~n60566 ;
  assign n60568 = ~\pi0238  & ~\pi0516  ;
  assign n60569 = n60567 & n60568 ;
  assign n60570 = \pi0245  & n60493 ;
  assign n60571 = ~\pi0514  & n60570 ;
  assign n60572 = ~\pi0244  & n60483 ;
  assign n60573 = ~\pi0558  & ~n60554 ;
  assign n60574 = ~n60551 & n60573 ;
  assign n60575 = ~n60548 & n60574 ;
  assign n60576 = \pi0244  & ~n60575 ;
  assign n60577 = ~n60572 & ~n60576 ;
  assign n60578 = ~\pi0235  & \pi0512  ;
  assign n60579 = n60473 & n60578 ;
  assign n60580 = ~\pi0242  & ~n60459 ;
  assign n60581 = \pi0242  & ~\pi0504  ;
  assign n60582 = ~n60548 & n60581 ;
  assign n60583 = ~n60580 & ~n60582 ;
  assign n60584 = ~\pi0240  & ~n60536 ;
  assign n60585 = ~\pi0515  & ~n60445 ;
  assign n60586 = ~n60442 & n60585 ;
  assign n60587 = \pi0240  & ~n60586 ;
  assign n60588 = ~n60584 & ~n60587 ;
  assign n60589 = ~\pi0534  & \pi0535  ;
  assign n60590 = n60588 & n60589 ;
  assign n60591 = ~\pi0559  & ~n60530 ;
  assign n60592 = ~\pi0241  & ~n60591 ;
  assign n60593 = ~\pi0506  & ~n60442 ;
  assign n60594 = n60592 & ~n60593 ;
  assign n60595 = \pi0559  & ~n60530 ;
  assign n60596 = \pi0241  & ~n60595 ;
  assign n60597 = \pi0506  & ~n60442 ;
  assign n60598 = n60596 & ~n60597 ;
  assign n60599 = ~n60594 & ~n60598 ;
  assign n60600 = \pi0515  & ~n60584 ;
  assign n60601 = n60589 & n60600 ;
  assign n60602 = n60599 & n60601 ;
  assign n60603 = ~n60590 & ~n60602 ;
  assign n60604 = \pi0240  & ~n60545 ;
  assign n60605 = \pi0515  & ~n60445 ;
  assign n60606 = ~n60442 & n60605 ;
  assign n60607 = ~\pi0240  & ~n60606 ;
  assign n60608 = ~n60604 & ~n60607 ;
  assign n60609 = ~\pi0534  & ~\pi0535  ;
  assign n60610 = n60608 & n60609 ;
  assign n60611 = ~\pi0515  & ~n60604 ;
  assign n60612 = n60609 & n60611 ;
  assign n60613 = n60599 & n60612 ;
  assign n60614 = ~n60610 & ~n60613 ;
  assign n60615 = ~\pi0240  & \pi0534  ;
  assign n60616 = n60536 & n60615 ;
  assign n60617 = \pi0240  & \pi0534  ;
  assign n60618 = n60545 & n60617 ;
  assign n60619 = ~n60616 & ~n60618 ;
  assign n60620 = n60537 & n60619 ;
  assign n60621 = n60614 & n60620 ;
  assign n60622 = n60603 & n60621 ;
  assign n60623 = ~n60449 & n60454 ;
  assign n60624 = ~n60442 & n60623 ;
  assign n60625 = ~\pi0239  & ~\pi0488  ;
  assign n60626 = ~n60624 & n60625 ;
  assign n60627 = n60446 & ~n60449 ;
  assign n60628 = ~n60442 & n60627 ;
  assign n60629 = \pi0239  & \pi0488  ;
  assign n60630 = ~n60628 & n60629 ;
  assign n60631 = ~n60626 & ~n60630 ;
  assign n60632 = ~n60622 & n60631 ;
  assign n60633 = \pi0534  & ~\pi0535  ;
  assign n60634 = n60608 & n60633 ;
  assign n60635 = n60611 & n60633 ;
  assign n60636 = n60599 & n60635 ;
  assign n60637 = ~n60634 & ~n60636 ;
  assign n60638 = \pi0534  & \pi0535  ;
  assign n60639 = n60588 & n60638 ;
  assign n60640 = n60600 & n60638 ;
  assign n60641 = n60599 & n60640 ;
  assign n60642 = ~n60639 & ~n60641 ;
  assign n60643 = ~\pi0240  & ~\pi0534  ;
  assign n60644 = n60536 & n60643 ;
  assign n60645 = \pi0240  & ~\pi0534  ;
  assign n60646 = n60545 & n60645 ;
  assign n60647 = ~n60644 & ~n60646 ;
  assign n60648 = n60538 & n60647 ;
  assign n60649 = n60642 & n60648 ;
  assign n60650 = n60637 & n60649 ;
  assign n60651 = ~\pi0242  & n60459 ;
  assign n60652 = \pi0504  & ~n60651 ;
  assign n60653 = ~n60650 & n60652 ;
  assign n60654 = n60632 & n60653 ;
  assign n60655 = n60583 & ~n60654 ;
  assign n60656 = \pi0510  & \pi0533  ;
  assign n60657 = ~n60655 & n60656 ;
  assign n60658 = \pi0242  & ~n60470 ;
  assign n60659 = ~\pi0242  & \pi0504  ;
  assign n60660 = ~n60548 & n60659 ;
  assign n60661 = ~n60658 & ~n60660 ;
  assign n60662 = \pi0242  & n60470 ;
  assign n60663 = ~\pi0504  & ~n60662 ;
  assign n60664 = ~n60650 & n60663 ;
  assign n60665 = n60632 & n60664 ;
  assign n60666 = n60661 & ~n60665 ;
  assign n60667 = ~\pi0510  & \pi0533  ;
  assign n60668 = ~n60666 & n60667 ;
  assign n60669 = ~n60657 & ~n60668 ;
  assign n60670 = ~\pi0533  & ~n60554 ;
  assign n60671 = ~n60548 & n60670 ;
  assign n60672 = n60550 & ~n60671 ;
  assign n60673 = n60669 & n60672 ;
  assign n60674 = ~n60579 & ~n60673 ;
  assign n60675 = \pi0510  & ~\pi0533  ;
  assign n60676 = ~n60655 & n60675 ;
  assign n60677 = ~\pi0510  & ~\pi0533  ;
  assign n60678 = ~n60666 & n60677 ;
  assign n60679 = ~n60676 & ~n60678 ;
  assign n60680 = \pi0533  & ~n60554 ;
  assign n60681 = ~n60548 & n60680 ;
  assign n60682 = n60549 & ~n60681 ;
  assign n60683 = n60679 & n60682 ;
  assign n60684 = \pi0235  & ~\pi0512  ;
  assign n60685 = n60480 & n60684 ;
  assign n60686 = \pi0558  & ~n60572 ;
  assign n60687 = ~n60685 & n60686 ;
  assign n60688 = ~n60683 & n60687 ;
  assign n60689 = n60674 & n60688 ;
  assign n60690 = ~n60577 & ~n60689 ;
  assign n60691 = ~\pi0509  & \pi0513  ;
  assign n60692 = ~n60690 & n60691 ;
  assign n60693 = \pi0244  & n60490 ;
  assign n60694 = \pi0558  & ~n60554 ;
  assign n60695 = ~n60551 & n60694 ;
  assign n60696 = ~n60548 & n60695 ;
  assign n60697 = ~\pi0244  & ~n60696 ;
  assign n60698 = ~n60693 & ~n60697 ;
  assign n60699 = ~\pi0558  & ~n60693 ;
  assign n60700 = ~n60685 & n60699 ;
  assign n60701 = ~n60683 & n60700 ;
  assign n60702 = n60674 & n60701 ;
  assign n60703 = ~n60698 & ~n60702 ;
  assign n60704 = ~\pi0509  & ~\pi0513  ;
  assign n60705 = ~n60703 & n60704 ;
  assign n60706 = ~n60692 & ~n60705 ;
  assign n60707 = \pi0509  & n60559 ;
  assign n60708 = ~n60548 & n60707 ;
  assign n60709 = ~\pi0245  & ~n60708 ;
  assign n60710 = ~\pi0514  & n60709 ;
  assign n60711 = n60706 & n60710 ;
  assign n60712 = ~n60571 & ~n60711 ;
  assign n60713 = \pi0509  & \pi0513  ;
  assign n60714 = ~n60690 & n60713 ;
  assign n60715 = \pi0509  & ~\pi0513  ;
  assign n60716 = ~n60703 & n60715 ;
  assign n60717 = ~n60714 & ~n60716 ;
  assign n60718 = ~\pi0509  & n60559 ;
  assign n60719 = ~n60548 & n60718 ;
  assign n60720 = \pi0245  & ~n60719 ;
  assign n60721 = \pi0514  & n60720 ;
  assign n60722 = n60717 & n60721 ;
  assign n60723 = ~\pi0245  & \pi0514  ;
  assign n60724 = n60500 & n60723 ;
  assign n60725 = ~n60504 & ~n60724 ;
  assign n60726 = ~n60722 & n60725 ;
  assign n60727 = n60712 & n60726 ;
  assign n60728 = ~\pi0508  & n60568 ;
  assign n60729 = n60727 & n60728 ;
  assign n60730 = ~n60569 & ~n60729 ;
  assign n60731 = ~\pi0238  & \pi0516  ;
  assign n60732 = ~\pi0517  & ~n60731 ;
  assign n60733 = ~\pi0245  & ~\pi0508  ;
  assign n60734 = ~n60500 & n60733 ;
  assign n60735 = \pi0245  & ~\pi0508  ;
  assign n60736 = ~n60493 & n60735 ;
  assign n60737 = ~n60734 & ~n60736 ;
  assign n60738 = ~\pi0247  & n60737 ;
  assign n60739 = \pi0508  & ~n60738 ;
  assign n60740 = ~n60724 & n60739 ;
  assign n60741 = ~n60722 & n60740 ;
  assign n60742 = n60712 & n60741 ;
  assign n60743 = ~\pi0508  & ~n60562 ;
  assign n60744 = n60559 & n60743 ;
  assign n60745 = ~n60548 & n60744 ;
  assign n60746 = \pi0247  & ~n60745 ;
  assign n60747 = ~n60738 & ~n60746 ;
  assign n60748 = ~\pi0517  & ~n60747 ;
  assign n60749 = ~n60742 & n60748 ;
  assign n60750 = ~n60732 & ~n60749 ;
  assign n60751 = n60730 & ~n60750 ;
  assign n60752 = ~\pi0238  & ~\pi0247  ;
  assign n60753 = ~n60737 & n60752 ;
  assign n60754 = ~\pi0238  & \pi0247  ;
  assign n60755 = ~n60503 & n60754 ;
  assign n60756 = ~n60753 & ~n60755 ;
  assign n60757 = \pi0238  & ~n60562 ;
  assign n60758 = ~\pi0247  & ~\pi0516  ;
  assign n60759 = \pi0247  & \pi0516  ;
  assign n60760 = ~n60758 & ~n60759 ;
  assign n60761 = n60757 & ~n60760 ;
  assign n60762 = n60559 & n60761 ;
  assign n60763 = ~n60548 & n60762 ;
  assign n60764 = \pi0517  & ~n60763 ;
  assign n60765 = n60756 & n60764 ;
  assign n60766 = ~\pi0507  & ~n60765 ;
  assign n60767 = ~n60751 & n60766 ;
  assign n60768 = \pi0238  & ~\pi0516  ;
  assign n60769 = n60567 & n60768 ;
  assign n60770 = ~\pi0508  & n60768 ;
  assign n60771 = n60727 & n60770 ;
  assign n60772 = ~n60769 & ~n60771 ;
  assign n60773 = \pi0238  & \pi0516  ;
  assign n60774 = \pi0517  & ~n60773 ;
  assign n60775 = \pi0517  & ~n60747 ;
  assign n60776 = ~n60742 & n60775 ;
  assign n60777 = ~n60774 & ~n60776 ;
  assign n60778 = n60772 & ~n60777 ;
  assign n60779 = \pi0238  & ~\pi0247  ;
  assign n60780 = ~n60737 & n60779 ;
  assign n60781 = \pi0238  & \pi0247  ;
  assign n60782 = ~n60503 & n60781 ;
  assign n60783 = ~n60780 & ~n60782 ;
  assign n60784 = ~\pi0238  & ~n60562 ;
  assign n60785 = ~n60760 & n60784 ;
  assign n60786 = n60559 & n60785 ;
  assign n60787 = ~n60548 & n60786 ;
  assign n60788 = ~\pi0517  & ~n60787 ;
  assign n60789 = n60783 & n60788 ;
  assign n60790 = \pi0507  & ~n60789 ;
  assign n60791 = ~n60778 & n60790 ;
  assign n60792 = ~n60767 & ~n60791 ;
  assign n60793 = \pi0233  & ~n60792 ;
  assign n60794 = \pi0249  & ~\pi0578  ;
  assign n60795 = ~\pi0249  & \pi0578  ;
  assign n60796 = ~n60794 & ~n60795 ;
  assign n60797 = \pi0248  & ~\pi0521  ;
  assign n60798 = ~\pi0246  & \pi0520  ;
  assign n60799 = ~n60797 & ~n60798 ;
  assign n60800 = n60796 & n60799 ;
  assign n60801 = ~\pi0248  & \pi0521  ;
  assign n60802 = \pi0246  & ~\pi0520  ;
  assign n60803 = ~n60801 & ~n60802 ;
  assign n60804 = ~\pi0241  & ~\pi0574  ;
  assign n60805 = \pi0241  & \pi0574  ;
  assign n60806 = ~n60804 & ~n60805 ;
  assign n60807 = n60803 & ~n60806 ;
  assign n60808 = n60800 & n60807 ;
  assign n60809 = ~\pi0518  & n60808 ;
  assign n60810 = ~n60508 & n60809 ;
  assign n60811 = \pi0518  & n60808 ;
  assign n60812 = ~n60525 & n60811 ;
  assign n60813 = ~n60810 & ~n60812 ;
  assign n60814 = \pi0239  & ~\pi0519  ;
  assign n60815 = ~\pi0239  & \pi0519  ;
  assign n60816 = ~n60814 & ~n60815 ;
  assign n60817 = \pi0240  & ~\pi0582  ;
  assign n60818 = ~\pi0240  & \pi0582  ;
  assign n60819 = ~n60817 & ~n60818 ;
  assign n60820 = ~n60816 & n60819 ;
  assign n60821 = ~n60813 & n60820 ;
  assign n60822 = ~\pi0242  & ~\pi0586  ;
  assign n60823 = \pi0242  & \pi0586  ;
  assign n60824 = ~n60822 & ~n60823 ;
  assign n60825 = ~\pi0585  & ~n60824 ;
  assign n60826 = ~\pi0235  & ~\pi0581  ;
  assign n60827 = \pi0235  & \pi0581  ;
  assign n60828 = ~n60826 & ~n60827 ;
  assign n60829 = ~\pi0244  & ~\pi0584  ;
  assign n60830 = ~n60828 & n60829 ;
  assign n60831 = n60825 & n60830 ;
  assign n60832 = n60821 & n60831 ;
  assign n60833 = \pi0585  & ~n60824 ;
  assign n60834 = \pi0244  & ~\pi0584  ;
  assign n60835 = ~n60828 & n60834 ;
  assign n60836 = n60833 & n60835 ;
  assign n60837 = n60821 & n60836 ;
  assign n60838 = ~n60832 & ~n60837 ;
  assign n60839 = ~\pi0247  & ~\pi0561  ;
  assign n60840 = \pi0247  & \pi0561  ;
  assign n60841 = ~n60839 & ~n60840 ;
  assign n60842 = ~\pi0245  & ~n60841 ;
  assign n60843 = ~n60838 & n60842 ;
  assign n60844 = ~\pi0244  & \pi0584  ;
  assign n60845 = ~n60828 & n60844 ;
  assign n60846 = n60825 & n60845 ;
  assign n60847 = n60821 & n60846 ;
  assign n60848 = \pi0244  & \pi0584  ;
  assign n60849 = ~n60828 & n60848 ;
  assign n60850 = n60833 & n60849 ;
  assign n60851 = n60821 & n60850 ;
  assign n60852 = ~n60847 & ~n60851 ;
  assign n60853 = \pi0245  & ~n60841 ;
  assign n60854 = ~n60852 & n60853 ;
  assign n60855 = ~n60843 & ~n60854 ;
  assign n60856 = \pi0238  & \pi0522  ;
  assign n60857 = n60855 & n60856 ;
  assign n60858 = \pi0248  & ~\pi0501  ;
  assign n60859 = ~\pi0248  & \pi0501  ;
  assign n60860 = ~n60858 & ~n60859 ;
  assign n60861 = \pi0246  & ~\pi0499  ;
  assign n60862 = ~\pi0249  & \pi0496  ;
  assign n60863 = ~n60861 & ~n60862 ;
  assign n60864 = n60860 & n60863 ;
  assign n60865 = ~\pi0246  & \pi0499  ;
  assign n60866 = \pi0249  & ~\pi0496  ;
  assign n60867 = ~n60865 & ~n60866 ;
  assign n60868 = ~\pi0241  & ~\pi0500  ;
  assign n60869 = \pi0241  & \pi0500  ;
  assign n60870 = ~n60868 & ~n60869 ;
  assign n60871 = n60867 & ~n60870 ;
  assign n60872 = n60864 & n60871 ;
  assign n60873 = ~\pi0505  & n60872 ;
  assign n60874 = n60419 & n60873 ;
  assign n60875 = \pi0505  & n60872 ;
  assign n60876 = n60437 & n60875 ;
  assign n60877 = ~n60874 & ~n60876 ;
  assign n60878 = ~\pi0240  & ~\pi0542  ;
  assign n60879 = \pi0240  & \pi0542  ;
  assign n60880 = ~n60878 & ~n60879 ;
  assign n60881 = \pi0239  & ~\pi0497  ;
  assign n60882 = ~\pi0239  & \pi0497  ;
  assign n60883 = ~n60881 & ~n60882 ;
  assign n60884 = ~n60880 & ~n60883 ;
  assign n60885 = ~n60877 & n60884 ;
  assign n60886 = ~\pi0242  & \pi0539  ;
  assign n60887 = \pi0242  & ~\pi0539  ;
  assign n60888 = ~\pi0540  & ~n60887 ;
  assign n60889 = ~n60886 & n60888 ;
  assign n60890 = n60885 & n60889 ;
  assign n60891 = ~\pi0244  & ~\pi0541  ;
  assign n60892 = \pi0244  & \pi0541  ;
  assign n60893 = ~n60891 & ~n60892 ;
  assign n60894 = ~\pi0235  & ~n60893 ;
  assign n60895 = n60890 & n60894 ;
  assign n60896 = \pi0242  & \pi0540  ;
  assign n60897 = \pi0539  & ~n60896 ;
  assign n60898 = ~\pi0242  & \pi0540  ;
  assign n60899 = ~\pi0539  & ~n60898 ;
  assign n60900 = ~n60897 & ~n60899 ;
  assign n60901 = n60885 & n60900 ;
  assign n60902 = \pi0235  & ~n60893 ;
  assign n60903 = n60901 & n60902 ;
  assign n60904 = ~n60895 & ~n60903 ;
  assign n60905 = ~\pi0245  & ~\pi0503  ;
  assign n60906 = \pi0245  & \pi0503  ;
  assign n60907 = ~n60905 & ~n60906 ;
  assign n60908 = ~\pi0247  & ~\pi0502  ;
  assign n60909 = \pi0247  & \pi0502  ;
  assign n60910 = ~n60908 & ~n60909 ;
  assign n60911 = ~n60907 & ~n60910 ;
  assign n60912 = ~n60904 & n60911 ;
  assign n60913 = ~\pi0238  & \pi0522  ;
  assign n60914 = ~n60912 & n60913 ;
  assign n60915 = ~n60857 & ~n60914 ;
  assign n60916 = \pi0522  & ~\pi0543  ;
  assign n60917 = n60915 & n60916 ;
  assign n60918 = ~\pi0502  & ~n60907 ;
  assign n60919 = \pi0561  & n60918 ;
  assign n60920 = ~n60904 & n60919 ;
  assign n60921 = ~\pi0247  & ~n60920 ;
  assign n60922 = ~\pi0235  & ~n60890 ;
  assign n60923 = ~\pi0540  & ~n60824 ;
  assign n60924 = n60821 & n60923 ;
  assign n60925 = \pi0235  & ~n60924 ;
  assign n60926 = ~n60922 & ~n60925 ;
  assign n60927 = \pi0539  & n60885 ;
  assign n60928 = \pi0242  & ~n60927 ;
  assign n60929 = ~\pi0586  & n60928 ;
  assign n60930 = ~\pi0497  & ~n60880 ;
  assign n60931 = ~n60877 & n60930 ;
  assign n60932 = \pi0239  & ~n60931 ;
  assign n60933 = ~\pi0239  & n60813 ;
  assign n60934 = ~\pi0240  & ~\pi0582  ;
  assign n60935 = ~\pi0497  & n60934 ;
  assign n60936 = \pi0240  & \pi0582  ;
  assign n60937 = ~\pi0497  & n60936 ;
  assign n60938 = ~\pi0239  & ~n60937 ;
  assign n60939 = ~n60935 & n60938 ;
  assign n60940 = ~n60933 & ~n60939 ;
  assign n60941 = ~n60932 & n60940 ;
  assign n60942 = \pi0519  & ~\pi0539  ;
  assign n60943 = n60941 & n60942 ;
  assign n60944 = ~\pi0582  & ~n60813 ;
  assign n60945 = ~\pi0240  & ~n60944 ;
  assign n60946 = ~\pi0542  & ~n60877 ;
  assign n60947 = n60945 & ~n60946 ;
  assign n60948 = \pi0582  & ~n60813 ;
  assign n60949 = \pi0240  & ~n60948 ;
  assign n60950 = \pi0542  & ~n60877 ;
  assign n60951 = n60949 & ~n60950 ;
  assign n60952 = ~n60947 & ~n60951 ;
  assign n60953 = n60882 & n60942 ;
  assign n60954 = n60952 & n60953 ;
  assign n60955 = ~n60943 & ~n60954 ;
  assign n60956 = \pi0497  & ~n60880 ;
  assign n60957 = ~n60877 & n60956 ;
  assign n60958 = ~\pi0239  & ~n60957 ;
  assign n60959 = \pi0497  & n60934 ;
  assign n60960 = \pi0497  & n60936 ;
  assign n60961 = ~n60959 & ~n60960 ;
  assign n60962 = ~n60813 & ~n60961 ;
  assign n60963 = \pi0239  & ~n60962 ;
  assign n60964 = ~n60958 & ~n60963 ;
  assign n60965 = ~\pi0519  & ~\pi0539  ;
  assign n60966 = n60964 & n60965 ;
  assign n60967 = n60881 & n60965 ;
  assign n60968 = n60952 & n60967 ;
  assign n60969 = ~n60966 & ~n60968 ;
  assign n60970 = n60955 & n60969 ;
  assign n60971 = \pi0539  & n60821 ;
  assign n60972 = ~\pi0242  & ~n60971 ;
  assign n60973 = ~\pi0586  & n60972 ;
  assign n60974 = n60970 & n60973 ;
  assign n60975 = ~n60929 & ~n60974 ;
  assign n60976 = \pi0519  & \pi0539  ;
  assign n60977 = n60941 & n60976 ;
  assign n60978 = n60882 & n60976 ;
  assign n60979 = n60952 & n60978 ;
  assign n60980 = ~n60977 & ~n60979 ;
  assign n60981 = ~\pi0519  & \pi0539  ;
  assign n60982 = n60964 & n60981 ;
  assign n60983 = n60881 & n60981 ;
  assign n60984 = n60952 & n60983 ;
  assign n60985 = ~n60982 & ~n60984 ;
  assign n60986 = n60980 & n60985 ;
  assign n60987 = ~\pi0539  & n60821 ;
  assign n60988 = \pi0242  & ~n60987 ;
  assign n60989 = \pi0586  & n60988 ;
  assign n60990 = n60986 & n60989 ;
  assign n60991 = ~\pi0539  & n60885 ;
  assign n60992 = ~\pi0242  & \pi0586  ;
  assign n60993 = ~n60991 & n60992 ;
  assign n60994 = \pi0540  & ~n60922 ;
  assign n60995 = ~n60993 & n60994 ;
  assign n60996 = ~n60990 & n60995 ;
  assign n60997 = n60975 & n60996 ;
  assign n60998 = ~n60926 & ~n60997 ;
  assign n60999 = \pi0581  & ~\pi0585  ;
  assign n61000 = ~n60998 & n60999 ;
  assign n61001 = ~\pi0581  & ~\pi0585  ;
  assign n61002 = ~\pi0235  & \pi0585  ;
  assign n61003 = n60890 & n61002 ;
  assign n61004 = \pi0235  & \pi0585  ;
  assign n61005 = n60901 & n61004 ;
  assign n61006 = ~n61003 & ~n61005 ;
  assign n61007 = n60891 & n61006 ;
  assign n61008 = ~n61001 & n61007 ;
  assign n61009 = \pi0235  & ~n60901 ;
  assign n61010 = ~\pi0540  & ~n61009 ;
  assign n61011 = ~n60993 & n61010 ;
  assign n61012 = ~n60990 & n61011 ;
  assign n61013 = n60975 & n61012 ;
  assign n61014 = \pi0540  & ~n60824 ;
  assign n61015 = n60821 & n61014 ;
  assign n61016 = ~\pi0235  & ~n61015 ;
  assign n61017 = ~n61009 & ~n61016 ;
  assign n61018 = n61007 & ~n61017 ;
  assign n61019 = ~n61013 & n61018 ;
  assign n61020 = ~n61008 & ~n61019 ;
  assign n61021 = ~n61000 & ~n61020 ;
  assign n61022 = ~n60828 & n60833 ;
  assign n61023 = n60821 & n61022 ;
  assign n61024 = \pi0244  & ~\pi0541  ;
  assign n61025 = ~n61023 & n61024 ;
  assign n61026 = n60825 & ~n60828 ;
  assign n61027 = n60821 & n61026 ;
  assign n61028 = ~\pi0244  & \pi0541  ;
  assign n61029 = ~n61027 & n61028 ;
  assign n61030 = ~n61025 & ~n61029 ;
  assign n61031 = ~n61021 & n61030 ;
  assign n61032 = ~n61013 & ~n61017 ;
  assign n61033 = ~\pi0581  & \pi0585  ;
  assign n61034 = ~n61032 & n61033 ;
  assign n61035 = \pi0581  & \pi0585  ;
  assign n61036 = ~\pi0235  & ~\pi0585  ;
  assign n61037 = n60890 & n61036 ;
  assign n61038 = \pi0235  & ~\pi0585  ;
  assign n61039 = n60901 & n61038 ;
  assign n61040 = ~n61037 & ~n61039 ;
  assign n61041 = n60892 & n61040 ;
  assign n61042 = ~n61035 & n61041 ;
  assign n61043 = ~n60926 & n61041 ;
  assign n61044 = ~n60997 & n61043 ;
  assign n61045 = ~n61042 & ~n61044 ;
  assign n61046 = ~n61034 & ~n61045 ;
  assign n61047 = ~\pi0245  & n60838 ;
  assign n61048 = \pi0584  & ~n61047 ;
  assign n61049 = ~n61046 & n61048 ;
  assign n61050 = n61031 & n61049 ;
  assign n61051 = ~\pi0245  & ~n60838 ;
  assign n61052 = \pi0245  & ~\pi0584  ;
  assign n61053 = ~n60904 & n61052 ;
  assign n61054 = ~n61051 & ~n61053 ;
  assign n61055 = ~\pi0502  & \pi0503  ;
  assign n61056 = n61054 & n61055 ;
  assign n61057 = ~n61050 & n61056 ;
  assign n61058 = \pi0245  & n60852 ;
  assign n61059 = ~\pi0584  & ~n61058 ;
  assign n61060 = ~n61046 & n61059 ;
  assign n61061 = n61031 & n61060 ;
  assign n61062 = \pi0245  & ~n60852 ;
  assign n61063 = ~\pi0245  & \pi0584  ;
  assign n61064 = ~n60904 & n61063 ;
  assign n61065 = ~n61062 & ~n61064 ;
  assign n61066 = ~\pi0502  & ~\pi0503  ;
  assign n61067 = n61065 & n61066 ;
  assign n61068 = ~n61061 & n61067 ;
  assign n61069 = ~\pi0245  & \pi0502  ;
  assign n61070 = n60838 & n61069 ;
  assign n61071 = \pi0245  & \pi0502  ;
  assign n61072 = n60852 & n61071 ;
  assign n61073 = ~\pi0561  & ~n61072 ;
  assign n61074 = ~n61070 & n61073 ;
  assign n61075 = ~n61068 & n61074 ;
  assign n61076 = ~n61057 & n61075 ;
  assign n61077 = n60921 & ~n61076 ;
  assign n61078 = \pi0502  & ~n60907 ;
  assign n61079 = ~\pi0561  & n61078 ;
  assign n61080 = ~n60904 & n61079 ;
  assign n61081 = \pi0247  & ~n61080 ;
  assign n61082 = \pi0502  & \pi0503  ;
  assign n61083 = n61054 & n61082 ;
  assign n61084 = ~n61050 & n61083 ;
  assign n61085 = \pi0502  & ~\pi0503  ;
  assign n61086 = n61065 & n61085 ;
  assign n61087 = ~n61061 & n61086 ;
  assign n61088 = ~n61084 & ~n61087 ;
  assign n61089 = ~\pi0245  & ~\pi0502  ;
  assign n61090 = n60838 & n61089 ;
  assign n61091 = \pi0245  & ~\pi0502  ;
  assign n61092 = n60852 & n61091 ;
  assign n61093 = \pi0561  & ~n61092 ;
  assign n61094 = ~n61090 & n61093 ;
  assign n61095 = n61088 & n61094 ;
  assign n61096 = n61081 & ~n61095 ;
  assign n61097 = ~n61077 & ~n61096 ;
  assign n61098 = ~\pi0238  & ~\pi0543  ;
  assign n61099 = n60915 & n61098 ;
  assign n61100 = n61097 & n61099 ;
  assign n61101 = ~n60917 & ~n61100 ;
  assign n61102 = ~\pi0238  & ~\pi0522  ;
  assign n61103 = n60855 & n61102 ;
  assign n61104 = \pi0238  & ~\pi0522  ;
  assign n61105 = ~n60912 & n61104 ;
  assign n61106 = ~n61103 & ~n61105 ;
  assign n61107 = ~\pi0522  & \pi0543  ;
  assign n61108 = n61106 & n61107 ;
  assign n61109 = \pi0238  & \pi0543  ;
  assign n61110 = n61106 & n61109 ;
  assign n61111 = n61097 & n61110 ;
  assign n61112 = ~n61108 & ~n61111 ;
  assign n61113 = n61101 & n61112 ;
  assign n61114 = ~\pi0233  & ~n61113 ;
  assign n61115 = \pi0237  & ~n61114 ;
  assign n61116 = ~n60793 & n61115 ;
  assign n61117 = ~\pi0239  & ~\pi0550  ;
  assign n61118 = \pi0239  & \pi0550  ;
  assign n61119 = ~n61117 & ~n61118 ;
  assign n61120 = ~\pi0249  & \pi0555  ;
  assign n61121 = \pi0242  & ~\pi0489  ;
  assign n61122 = ~n61120 & ~n61121 ;
  assign n61123 = n61119 & n61122 ;
  assign n61124 = ~\pi0248  & \pi0554  ;
  assign n61125 = ~\pi0240  & \pi0551  ;
  assign n61126 = ~n61124 & ~n61125 ;
  assign n61127 = n61123 & n61126 ;
  assign n61128 = ~\pi0246  & \pi0563  ;
  assign n61129 = \pi0241  & ~\pi0553  ;
  assign n61130 = ~n61128 & ~n61129 ;
  assign n61131 = ~\pi0242  & \pi0489  ;
  assign n61132 = \pi0240  & ~\pi0551  ;
  assign n61133 = ~n61131 & ~n61132 ;
  assign n61134 = n61130 & n61133 ;
  assign n61135 = \pi0249  & ~\pi0555  ;
  assign n61136 = \pi0248  & ~\pi0554  ;
  assign n61137 = ~n61135 & ~n61136 ;
  assign n61138 = ~\pi0241  & \pi0553  ;
  assign n61139 = \pi0246  & ~\pi0563  ;
  assign n61140 = ~n61138 & ~n61139 ;
  assign n61141 = n61137 & n61140 ;
  assign n61142 = n61134 & n61141 ;
  assign n61143 = n61127 & n61142 ;
  assign n61144 = ~\pi0485  & n61143 ;
  assign n61145 = n60419 & n61144 ;
  assign n61146 = \pi0485  & n61143 ;
  assign n61147 = n60437 & n61146 ;
  assign n61148 = ~n61145 & ~n61147 ;
  assign n61149 = ~\pi0235  & ~\pi0549  ;
  assign n61150 = ~\pi0486  & n61149 ;
  assign n61151 = \pi0235  & \pi0549  ;
  assign n61152 = ~\pi0486  & n61151 ;
  assign n61153 = ~n61150 & ~n61152 ;
  assign n61154 = ~n61148 & ~n61153 ;
  assign n61155 = ~\pi0245  & ~\pi0580  ;
  assign n61156 = \pi0245  & \pi0580  ;
  assign n61157 = ~n61155 & ~n61156 ;
  assign n61158 = ~\pi0244  & ~n61157 ;
  assign n61159 = n61154 & n61158 ;
  assign n61160 = \pi0486  & n61149 ;
  assign n61161 = \pi0486  & n61151 ;
  assign n61162 = ~n61160 & ~n61161 ;
  assign n61163 = ~n61148 & ~n61162 ;
  assign n61164 = \pi0244  & ~n61157 ;
  assign n61165 = n61163 & n61164 ;
  assign n61166 = ~n61159 & ~n61165 ;
  assign n61167 = \pi0552  & ~n61166 ;
  assign n61168 = \pi0247  & ~n61167 ;
  assign n61169 = \pi0242  & ~\pi0556  ;
  assign n61170 = ~\pi0242  & \pi0556  ;
  assign n61171 = ~n61169 & ~n61170 ;
  assign n61172 = ~\pi0248  & \pi0565  ;
  assign n61173 = ~\pi0239  & ~\pi0569  ;
  assign n61174 = ~n61172 & ~n61173 ;
  assign n61175 = n61171 & n61174 ;
  assign n61176 = ~\pi0246  & \pi0564  ;
  assign n61177 = ~\pi0241  & \pi0562  ;
  assign n61178 = ~n61176 & ~n61177 ;
  assign n61179 = n61175 & n61178 ;
  assign n61180 = ~\pi0240  & \pi0560  ;
  assign n61181 = \pi0249  & ~\pi0482  ;
  assign n61182 = ~n61180 & ~n61181 ;
  assign n61183 = \pi0239  & \pi0569  ;
  assign n61184 = \pi0241  & ~\pi0562  ;
  assign n61185 = ~n61183 & ~n61184 ;
  assign n61186 = n61182 & n61185 ;
  assign n61187 = \pi0248  & ~\pi0565  ;
  assign n61188 = \pi0246  & ~\pi0564  ;
  assign n61189 = ~n61187 & ~n61188 ;
  assign n61190 = ~\pi0249  & \pi0482  ;
  assign n61191 = \pi0240  & ~\pi0560  ;
  assign n61192 = ~n61190 & ~n61191 ;
  assign n61193 = n61189 & n61192 ;
  assign n61194 = n61186 & n61193 ;
  assign n61195 = n61179 & n61194 ;
  assign n61196 = ~\pi0570  & n61195 ;
  assign n61197 = ~n60508 & n61196 ;
  assign n61198 = \pi0570  & n61195 ;
  assign n61199 = ~n60525 & n61198 ;
  assign n61200 = ~n61197 & ~n61199 ;
  assign n61201 = ~\pi0235  & ~\pi0531  ;
  assign n61202 = \pi0235  & \pi0531  ;
  assign n61203 = ~n61201 & ~n61202 ;
  assign n61204 = \pi0568  & ~n61203 ;
  assign n61205 = ~\pi0244  & ~\pi0566  ;
  assign n61206 = \pi0244  & \pi0566  ;
  assign n61207 = ~n61205 & ~n61206 ;
  assign n61208 = \pi0245  & \pi0552  ;
  assign n61209 = ~n61207 & n61208 ;
  assign n61210 = n61204 & n61209 ;
  assign n61211 = ~n61200 & n61210 ;
  assign n61212 = ~\pi0568  & ~n61203 ;
  assign n61213 = ~\pi0245  & \pi0552  ;
  assign n61214 = ~n61207 & n61213 ;
  assign n61215 = n61212 & n61214 ;
  assign n61216 = ~n61200 & n61215 ;
  assign n61217 = ~\pi0247  & ~n61216 ;
  assign n61218 = ~n61211 & n61217 ;
  assign n61219 = ~n61168 & ~n61218 ;
  assign n61220 = ~\pi0244  & ~n61154 ;
  assign n61221 = ~\pi0486  & ~n61203 ;
  assign n61222 = ~n61200 & n61221 ;
  assign n61223 = \pi0244  & ~n61222 ;
  assign n61224 = ~n61220 & ~n61223 ;
  assign n61225 = \pi0566  & ~\pi0568  ;
  assign n61226 = n61224 & n61225 ;
  assign n61227 = ~\pi0549  & ~n61148 ;
  assign n61228 = ~\pi0235  & ~n61227 ;
  assign n61229 = ~\pi0531  & ~n61200 ;
  assign n61230 = n61228 & ~n61229 ;
  assign n61231 = \pi0549  & ~n61148 ;
  assign n61232 = \pi0235  & ~n61231 ;
  assign n61233 = \pi0531  & ~n61200 ;
  assign n61234 = n61232 & ~n61233 ;
  assign n61235 = ~n61230 & ~n61234 ;
  assign n61236 = \pi0486  & ~n61220 ;
  assign n61237 = n61225 & n61236 ;
  assign n61238 = n61235 & n61237 ;
  assign n61239 = ~n61226 & ~n61238 ;
  assign n61240 = \pi0244  & ~n61163 ;
  assign n61241 = \pi0486  & ~n61203 ;
  assign n61242 = ~n61200 & n61241 ;
  assign n61243 = ~\pi0244  & ~n61242 ;
  assign n61244 = ~n61240 & ~n61243 ;
  assign n61245 = ~\pi0566  & ~\pi0568  ;
  assign n61246 = n61244 & n61245 ;
  assign n61247 = ~\pi0486  & ~n61240 ;
  assign n61248 = n61245 & n61247 ;
  assign n61249 = n61235 & n61248 ;
  assign n61250 = ~n61246 & ~n61249 ;
  assign n61251 = ~\pi0244  & \pi0568  ;
  assign n61252 = n61154 & n61251 ;
  assign n61253 = \pi0244  & \pi0568  ;
  assign n61254 = n61163 & n61253 ;
  assign n61255 = ~n61252 & ~n61254 ;
  assign n61256 = n61155 & n61255 ;
  assign n61257 = n61250 & n61256 ;
  assign n61258 = n61239 & n61257 ;
  assign n61259 = n61204 & ~n61207 ;
  assign n61260 = ~n61200 & n61259 ;
  assign n61261 = \pi0245  & ~\pi0580  ;
  assign n61262 = ~n61260 & n61261 ;
  assign n61263 = ~n61207 & n61212 ;
  assign n61264 = ~n61200 & n61263 ;
  assign n61265 = ~\pi0245  & \pi0580  ;
  assign n61266 = ~n61264 & n61265 ;
  assign n61267 = ~n61262 & ~n61266 ;
  assign n61268 = ~n61258 & n61267 ;
  assign n61269 = ~\pi0566  & \pi0568  ;
  assign n61270 = n61244 & n61269 ;
  assign n61271 = n61247 & n61269 ;
  assign n61272 = n61235 & n61271 ;
  assign n61273 = ~n61270 & ~n61272 ;
  assign n61274 = \pi0566  & \pi0568  ;
  assign n61275 = n61224 & n61274 ;
  assign n61276 = n61236 & n61274 ;
  assign n61277 = n61235 & n61276 ;
  assign n61278 = ~n61275 & ~n61277 ;
  assign n61279 = ~\pi0244  & ~\pi0568  ;
  assign n61280 = n61154 & n61279 ;
  assign n61281 = \pi0244  & ~\pi0568  ;
  assign n61282 = n61163 & n61281 ;
  assign n61283 = ~n61280 & ~n61282 ;
  assign n61284 = n61156 & n61283 ;
  assign n61285 = n61278 & n61284 ;
  assign n61286 = n61273 & n61285 ;
  assign n61287 = ~\pi0552  & ~n61168 ;
  assign n61288 = ~n61286 & n61287 ;
  assign n61289 = n61268 & n61288 ;
  assign n61290 = ~n61219 & ~n61289 ;
  assign n61291 = ~\pi0238  & ~\pi0532  ;
  assign n61292 = ~n61290 & n61291 ;
  assign n61293 = ~\pi0238  & \pi0532  ;
  assign n61294 = ~\pi0577  & ~n61293 ;
  assign n61295 = \pi0247  & \pi0552  ;
  assign n61296 = ~n61286 & n61295 ;
  assign n61297 = n61268 & n61296 ;
  assign n61298 = ~\pi0552  & ~n61166 ;
  assign n61299 = ~\pi0247  & ~n61298 ;
  assign n61300 = \pi0245  & ~\pi0552  ;
  assign n61301 = ~n61207 & n61300 ;
  assign n61302 = n61204 & n61301 ;
  assign n61303 = ~n61200 & n61302 ;
  assign n61304 = ~\pi0245  & ~\pi0552  ;
  assign n61305 = ~n61207 & n61304 ;
  assign n61306 = n61212 & n61305 ;
  assign n61307 = ~n61200 & n61306 ;
  assign n61308 = \pi0247  & ~n61307 ;
  assign n61309 = ~n61303 & n61308 ;
  assign n61310 = ~n61299 & ~n61309 ;
  assign n61311 = ~\pi0577  & ~n61310 ;
  assign n61312 = ~n61297 & n61311 ;
  assign n61313 = ~n61294 & ~n61312 ;
  assign n61314 = ~n61292 & ~n61313 ;
  assign n61315 = \pi0238  & \pi0552  ;
  assign n61316 = \pi0247  & n61315 ;
  assign n61317 = ~n60779 & ~n61316 ;
  assign n61318 = \pi0552  & ~n61316 ;
  assign n61319 = ~n61317 & ~n61318 ;
  assign n61320 = ~n61166 & n61319 ;
  assign n61321 = ~\pi0247  & ~\pi0532  ;
  assign n61322 = \pi0247  & \pi0532  ;
  assign n61323 = ~n61321 & ~n61322 ;
  assign n61324 = ~\pi0245  & ~n61323 ;
  assign n61325 = n61264 & n61324 ;
  assign n61326 = \pi0245  & ~n61323 ;
  assign n61327 = n61260 & n61326 ;
  assign n61328 = ~n61325 & ~n61327 ;
  assign n61329 = ~\pi0238  & ~n61328 ;
  assign n61330 = ~n61320 & ~n61329 ;
  assign n61331 = \pi0577  & n61330 ;
  assign n61332 = ~\pi0498  & ~n61331 ;
  assign n61333 = ~n61314 & n61332 ;
  assign n61334 = \pi0238  & ~\pi0532  ;
  assign n61335 = ~n61290 & n61334 ;
  assign n61336 = \pi0238  & \pi0532  ;
  assign n61337 = \pi0577  & ~n61336 ;
  assign n61338 = \pi0577  & ~n61310 ;
  assign n61339 = ~n61297 & n61338 ;
  assign n61340 = ~n61337 & ~n61339 ;
  assign n61341 = ~n61335 & ~n61340 ;
  assign n61342 = \pi0247  & ~\pi0552  ;
  assign n61343 = ~\pi0247  & \pi0552  ;
  assign n61344 = ~\pi0238  & ~n61343 ;
  assign n61345 = ~n61342 & n61344 ;
  assign n61346 = ~n61166 & n61345 ;
  assign n61347 = \pi0238  & ~n61328 ;
  assign n61348 = ~n61346 & ~n61347 ;
  assign n61349 = ~\pi0577  & n61348 ;
  assign n61350 = \pi0498  & ~n61349 ;
  assign n61351 = ~n61341 & n61350 ;
  assign n61352 = ~n61333 & ~n61351 ;
  assign n61353 = ~\pi0233  & ~n61352 ;
  assign n61354 = ~\pi0233  & ~n61353 ;
  assign n61355 = ~\pi0246  & \pi0546  ;
  assign n61356 = \pi0249  & ~\pi0484  ;
  assign n61357 = ~\pi0249  & \pi0484  ;
  assign n61358 = ~n61356 & ~n61357 ;
  assign n61359 = ~n61355 & n61358 ;
  assign n61360 = ~\pi0248  & ~\pi0548  ;
  assign n61361 = \pi0248  & \pi0548  ;
  assign n61362 = ~n61360 & ~n61361 ;
  assign n61363 = \pi0246  & ~\pi0546  ;
  assign n61364 = ~\pi0544  & ~n61363 ;
  assign n61365 = ~n61362 & n61364 ;
  assign n61366 = n61359 & n61365 ;
  assign n61367 = n60419 & n61366 ;
  assign n61368 = \pi0544  & ~n61363 ;
  assign n61369 = ~n61362 & n61368 ;
  assign n61370 = n61359 & n61369 ;
  assign n61371 = n60437 & n61370 ;
  assign n61372 = ~n61367 & ~n61371 ;
  assign n61373 = ~\pi0241  & ~\pi0490  ;
  assign n61374 = \pi0241  & \pi0490  ;
  assign n61375 = ~n61373 & ~n61374 ;
  assign n61376 = ~\pi0494  & ~n61375 ;
  assign n61377 = ~\pi0240  & ~\pi0492  ;
  assign n61378 = \pi0240  & \pi0492  ;
  assign n61379 = ~n61377 & ~n61378 ;
  assign n61380 = \pi0239  & ~\pi0483  ;
  assign n61381 = ~n61379 & n61380 ;
  assign n61382 = n61376 & n61381 ;
  assign n61383 = ~n61372 & n61382 ;
  assign n61384 = \pi0494  & ~n61375 ;
  assign n61385 = ~\pi0239  & ~\pi0483  ;
  assign n61386 = ~n61379 & n61385 ;
  assign n61387 = n61384 & n61386 ;
  assign n61388 = ~n61372 & n61387 ;
  assign n61389 = ~n61383 & ~n61388 ;
  assign n61390 = ~\pi0242  & ~\pi0495  ;
  assign n61391 = ~n61389 & n61390 ;
  assign n61392 = \pi0239  & \pi0483  ;
  assign n61393 = ~n61379 & n61392 ;
  assign n61394 = n61376 & n61393 ;
  assign n61395 = ~n61372 & n61394 ;
  assign n61396 = ~\pi0239  & \pi0483  ;
  assign n61397 = ~n61379 & n61396 ;
  assign n61398 = n61384 & n61397 ;
  assign n61399 = ~n61372 & n61398 ;
  assign n61400 = ~n61395 & ~n61399 ;
  assign n61401 = \pi0242  & ~\pi0495  ;
  assign n61402 = ~n61400 & n61401 ;
  assign n61403 = ~n61391 & ~n61402 ;
  assign n61404 = ~\pi0244  & ~\pi0493  ;
  assign n61405 = \pi0244  & \pi0493  ;
  assign n61406 = ~n61404 & ~n61405 ;
  assign n61407 = ~\pi0235  & ~n61406 ;
  assign n61408 = ~n61403 & n61407 ;
  assign n61409 = ~\pi0242  & \pi0495  ;
  assign n61410 = ~n61389 & n61409 ;
  assign n61411 = \pi0242  & \pi0495  ;
  assign n61412 = ~n61400 & n61411 ;
  assign n61413 = ~n61410 & ~n61412 ;
  assign n61414 = \pi0235  & ~n61406 ;
  assign n61415 = ~n61413 & n61414 ;
  assign n61416 = ~n61408 & ~n61415 ;
  assign n61417 = ~\pi0245  & ~\pi0547  ;
  assign n61418 = ~\pi0545  & n61417 ;
  assign n61419 = \pi0245  & ~\pi0547  ;
  assign n61420 = \pi0545  & n61419 ;
  assign n61421 = ~n61418 & ~n61420 ;
  assign n61422 = ~n61416 & ~n61421 ;
  assign n61423 = ~\pi0247  & \pi0527  ;
  assign n61424 = ~n61422 & n61423 ;
  assign n61425 = ~\pi0545  & ~n61416 ;
  assign n61426 = ~\pi0245  & ~n61425 ;
  assign n61427 = ~\pi0246  & \pi0526  ;
  assign n61428 = \pi0249  & ~\pi0528  ;
  assign n61429 = ~\pi0249  & \pi0528  ;
  assign n61430 = ~n61428 & ~n61429 ;
  assign n61431 = ~n61427 & n61430 ;
  assign n61432 = ~\pi0248  & ~\pi0576  ;
  assign n61433 = \pi0248  & \pi0576  ;
  assign n61434 = ~n61432 & ~n61433 ;
  assign n61435 = \pi0246  & ~\pi0526  ;
  assign n61436 = ~\pi0523  & ~n61435 ;
  assign n61437 = ~n61434 & n61436 ;
  assign n61438 = n61431 & n61437 ;
  assign n61439 = ~n60508 & n61438 ;
  assign n61440 = \pi0523  & ~n61435 ;
  assign n61441 = ~n61434 & n61440 ;
  assign n61442 = n61431 & n61441 ;
  assign n61443 = ~n60525 & n61442 ;
  assign n61444 = ~n61439 & ~n61443 ;
  assign n61445 = ~\pi0241  & ~\pi0571  ;
  assign n61446 = \pi0530  & n61445 ;
  assign n61447 = \pi0241  & \pi0571  ;
  assign n61448 = \pi0530  & n61447 ;
  assign n61449 = ~n61446 & ~n61448 ;
  assign n61450 = ~n61444 & ~n61449 ;
  assign n61451 = \pi0239  & ~\pi0524  ;
  assign n61452 = ~\pi0239  & \pi0524  ;
  assign n61453 = ~n61451 & ~n61452 ;
  assign n61454 = \pi0240  & ~n61453 ;
  assign n61455 = n61450 & n61454 ;
  assign n61456 = ~\pi0530  & n61445 ;
  assign n61457 = ~\pi0530  & n61447 ;
  assign n61458 = ~n61456 & ~n61457 ;
  assign n61459 = ~n61444 & ~n61458 ;
  assign n61460 = ~\pi0240  & ~n61453 ;
  assign n61461 = n61459 & n61460 ;
  assign n61462 = ~n61455 & ~n61461 ;
  assign n61463 = ~\pi0242  & ~\pi0573  ;
  assign n61464 = \pi0242  & \pi0573  ;
  assign n61465 = ~n61463 & ~n61464 ;
  assign n61466 = \pi0572  & ~n61465 ;
  assign n61467 = ~\pi0235  & ~\pi0575  ;
  assign n61468 = \pi0235  & \pi0575  ;
  assign n61469 = ~n61467 & ~n61468 ;
  assign n61470 = \pi0244  & ~\pi0545  ;
  assign n61471 = ~n61469 & n61470 ;
  assign n61472 = n61466 & n61471 ;
  assign n61473 = ~n61462 & n61472 ;
  assign n61474 = ~\pi0572  & ~n61465 ;
  assign n61475 = ~\pi0244  & ~\pi0545  ;
  assign n61476 = ~n61469 & n61475 ;
  assign n61477 = n61474 & n61476 ;
  assign n61478 = ~n61462 & n61477 ;
  assign n61479 = \pi0245  & ~n61478 ;
  assign n61480 = ~n61473 & n61479 ;
  assign n61481 = ~n61426 & ~n61480 ;
  assign n61482 = ~\pi0235  & n61403 ;
  assign n61483 = ~\pi0495  & ~n61465 ;
  assign n61484 = ~n61462 & n61483 ;
  assign n61485 = \pi0235  & ~n61484 ;
  assign n61486 = ~n61482 & ~n61485 ;
  assign n61487 = \pi0242  & n61400 ;
  assign n61488 = ~\pi0573  & n61487 ;
  assign n61489 = n61376 & ~n61379 ;
  assign n61490 = ~n61372 & n61489 ;
  assign n61491 = \pi0239  & ~n61490 ;
  assign n61492 = ~\pi0240  & ~\pi0494  ;
  assign n61493 = n61459 & n61492 ;
  assign n61494 = \pi0240  & ~\pi0494  ;
  assign n61495 = n61450 & n61494 ;
  assign n61496 = ~\pi0239  & ~n61495 ;
  assign n61497 = ~n61493 & n61496 ;
  assign n61498 = ~n61491 & ~n61497 ;
  assign n61499 = ~\pi0483  & \pi0524  ;
  assign n61500 = n61498 & n61499 ;
  assign n61501 = \pi0492  & n61459 ;
  assign n61502 = ~\pi0240  & ~n61501 ;
  assign n61503 = ~\pi0492  & ~\pi0530  ;
  assign n61504 = ~\pi0492  & ~n61375 ;
  assign n61505 = ~n61372 & n61504 ;
  assign n61506 = ~n61503 & ~n61505 ;
  assign n61507 = n61502 & n61506 ;
  assign n61508 = ~\pi0571  & ~n61444 ;
  assign n61509 = ~\pi0241  & ~n61508 ;
  assign n61510 = ~\pi0490  & ~n61372 ;
  assign n61511 = n61509 & ~n61510 ;
  assign n61512 = \pi0571  & ~n61444 ;
  assign n61513 = \pi0241  & ~n61512 ;
  assign n61514 = \pi0490  & ~n61372 ;
  assign n61515 = n61513 & ~n61514 ;
  assign n61516 = ~n61511 & ~n61515 ;
  assign n61517 = ~\pi0530  & n61502 ;
  assign n61518 = ~n61516 & n61517 ;
  assign n61519 = ~n61507 & ~n61518 ;
  assign n61520 = ~\pi0492  & n61450 ;
  assign n61521 = \pi0240  & ~n61520 ;
  assign n61522 = \pi0492  & \pi0530  ;
  assign n61523 = \pi0492  & ~n61375 ;
  assign n61524 = ~n61372 & n61523 ;
  assign n61525 = ~n61522 & ~n61524 ;
  assign n61526 = n61521 & n61525 ;
  assign n61527 = \pi0530  & n61521 ;
  assign n61528 = ~n61516 & n61527 ;
  assign n61529 = ~n61526 & ~n61528 ;
  assign n61530 = n61519 & n61529 ;
  assign n61531 = ~\pi0239  & \pi0494  ;
  assign n61532 = n61499 & n61531 ;
  assign n61533 = n61530 & n61532 ;
  assign n61534 = ~n61500 & ~n61533 ;
  assign n61535 = ~n61379 & n61384 ;
  assign n61536 = ~n61372 & n61535 ;
  assign n61537 = ~\pi0239  & ~n61536 ;
  assign n61538 = ~\pi0240  & \pi0494  ;
  assign n61539 = n61459 & n61538 ;
  assign n61540 = \pi0240  & \pi0494  ;
  assign n61541 = n61450 & n61540 ;
  assign n61542 = \pi0239  & ~n61541 ;
  assign n61543 = ~n61539 & n61542 ;
  assign n61544 = ~n61537 & ~n61543 ;
  assign n61545 = ~\pi0483  & ~\pi0524  ;
  assign n61546 = n61544 & n61545 ;
  assign n61547 = \pi0239  & ~\pi0494  ;
  assign n61548 = n61545 & n61547 ;
  assign n61549 = n61530 & n61548 ;
  assign n61550 = ~n61546 & ~n61549 ;
  assign n61551 = n61534 & n61550 ;
  assign n61552 = \pi0483  & ~n61462 ;
  assign n61553 = ~\pi0242  & ~n61552 ;
  assign n61554 = ~\pi0573  & n61553 ;
  assign n61555 = n61551 & n61554 ;
  assign n61556 = ~n61488 & ~n61555 ;
  assign n61557 = \pi0483  & \pi0524  ;
  assign n61558 = n61498 & n61557 ;
  assign n61559 = n61531 & n61557 ;
  assign n61560 = n61530 & n61559 ;
  assign n61561 = ~n61558 & ~n61560 ;
  assign n61562 = \pi0483  & ~\pi0524  ;
  assign n61563 = n61544 & n61562 ;
  assign n61564 = n61547 & n61562 ;
  assign n61565 = n61530 & n61564 ;
  assign n61566 = ~n61563 & ~n61565 ;
  assign n61567 = n61561 & n61566 ;
  assign n61568 = ~\pi0483  & ~n61462 ;
  assign n61569 = \pi0242  & ~n61568 ;
  assign n61570 = \pi0573  & n61569 ;
  assign n61571 = n61567 & n61570 ;
  assign n61572 = ~\pi0242  & \pi0573  ;
  assign n61573 = n61389 & n61572 ;
  assign n61574 = \pi0495  & ~n61482 ;
  assign n61575 = ~n61573 & n61574 ;
  assign n61576 = ~n61571 & n61575 ;
  assign n61577 = n61556 & n61576 ;
  assign n61578 = ~n61486 & ~n61577 ;
  assign n61579 = ~\pi0572  & \pi0575  ;
  assign n61580 = ~n61578 & n61579 ;
  assign n61581 = ~\pi0572  & ~\pi0575  ;
  assign n61582 = ~\pi0235  & \pi0572  ;
  assign n61583 = ~n61403 & n61582 ;
  assign n61584 = \pi0235  & \pi0572  ;
  assign n61585 = ~n61413 & n61584 ;
  assign n61586 = ~n61583 & ~n61585 ;
  assign n61587 = n61404 & n61586 ;
  assign n61588 = ~n61581 & n61587 ;
  assign n61589 = \pi0235  & n61413 ;
  assign n61590 = ~\pi0495  & ~n61589 ;
  assign n61591 = ~n61573 & n61590 ;
  assign n61592 = ~n61571 & n61591 ;
  assign n61593 = n61556 & n61592 ;
  assign n61594 = \pi0495  & ~n61465 ;
  assign n61595 = ~n61462 & n61594 ;
  assign n61596 = ~\pi0235  & ~n61595 ;
  assign n61597 = ~n61589 & ~n61596 ;
  assign n61598 = n61587 & ~n61597 ;
  assign n61599 = ~n61593 & n61598 ;
  assign n61600 = ~n61588 & ~n61599 ;
  assign n61601 = ~n61580 & ~n61600 ;
  assign n61602 = n61466 & ~n61469 ;
  assign n61603 = ~n61462 & n61602 ;
  assign n61604 = \pi0244  & ~\pi0493  ;
  assign n61605 = ~n61603 & n61604 ;
  assign n61606 = ~n61469 & n61474 ;
  assign n61607 = ~n61462 & n61606 ;
  assign n61608 = ~\pi0244  & \pi0493  ;
  assign n61609 = ~n61607 & n61608 ;
  assign n61610 = ~n61605 & ~n61609 ;
  assign n61611 = ~n61601 & n61610 ;
  assign n61612 = ~n61593 & ~n61597 ;
  assign n61613 = \pi0572  & ~\pi0575  ;
  assign n61614 = ~n61612 & n61613 ;
  assign n61615 = \pi0572  & \pi0575  ;
  assign n61616 = ~\pi0235  & ~\pi0572  ;
  assign n61617 = ~n61403 & n61616 ;
  assign n61618 = \pi0235  & ~\pi0572  ;
  assign n61619 = ~n61413 & n61618 ;
  assign n61620 = ~n61617 & ~n61619 ;
  assign n61621 = n61405 & n61620 ;
  assign n61622 = ~n61615 & n61621 ;
  assign n61623 = ~n61486 & n61621 ;
  assign n61624 = ~n61577 & n61623 ;
  assign n61625 = ~n61622 & ~n61624 ;
  assign n61626 = ~n61614 & ~n61625 ;
  assign n61627 = \pi0245  & \pi0545  ;
  assign n61628 = ~n61626 & n61627 ;
  assign n61629 = n61611 & n61628 ;
  assign n61630 = ~n61481 & ~n61629 ;
  assign n61631 = \pi0525  & \pi0547  ;
  assign n61632 = ~n61630 & n61631 ;
  assign n61633 = \pi0545  & ~n61416 ;
  assign n61634 = \pi0245  & ~n61633 ;
  assign n61635 = \pi0244  & \pi0545  ;
  assign n61636 = ~n61469 & n61635 ;
  assign n61637 = n61466 & n61636 ;
  assign n61638 = ~n61462 & n61637 ;
  assign n61639 = ~\pi0244  & \pi0545  ;
  assign n61640 = ~n61469 & n61639 ;
  assign n61641 = n61474 & n61640 ;
  assign n61642 = ~n61462 & n61641 ;
  assign n61643 = ~\pi0245  & ~n61642 ;
  assign n61644 = ~n61638 & n61643 ;
  assign n61645 = ~n61634 & ~n61644 ;
  assign n61646 = ~\pi0545  & ~n61634 ;
  assign n61647 = ~n61626 & n61646 ;
  assign n61648 = n61611 & n61647 ;
  assign n61649 = ~n61645 & ~n61648 ;
  assign n61650 = ~\pi0525  & \pi0547  ;
  assign n61651 = ~n61649 & n61650 ;
  assign n61652 = ~n61632 & ~n61651 ;
  assign n61653 = ~\pi0245  & ~\pi0525  ;
  assign n61654 = \pi0245  & \pi0525  ;
  assign n61655 = ~n61653 & ~n61654 ;
  assign n61656 = ~\pi0244  & ~n61655 ;
  assign n61657 = n61606 & n61656 ;
  assign n61658 = ~n61462 & n61657 ;
  assign n61659 = \pi0244  & ~n61655 ;
  assign n61660 = n61602 & n61659 ;
  assign n61661 = ~n61462 & n61660 ;
  assign n61662 = ~n61658 & ~n61661 ;
  assign n61663 = ~\pi0547  & ~n61662 ;
  assign n61664 = \pi0247  & \pi0527  ;
  assign n61665 = ~n61663 & n61664 ;
  assign n61666 = n61652 & n61665 ;
  assign n61667 = ~n61424 & ~n61666 ;
  assign n61668 = \pi0525  & ~\pi0547  ;
  assign n61669 = ~n61630 & n61668 ;
  assign n61670 = ~\pi0525  & ~\pi0547  ;
  assign n61671 = ~n61649 & n61670 ;
  assign n61672 = ~n61669 & ~n61671 ;
  assign n61673 = \pi0547  & ~n61662 ;
  assign n61674 = ~\pi0247  & ~\pi0527  ;
  assign n61675 = ~n61673 & n61674 ;
  assign n61676 = n61672 & n61675 ;
  assign n61677 = ~\pi0245  & \pi0547  ;
  assign n61678 = ~\pi0545  & n61677 ;
  assign n61679 = \pi0245  & \pi0547  ;
  assign n61680 = \pi0545  & n61679 ;
  assign n61681 = ~n61678 & ~n61680 ;
  assign n61682 = ~n61416 & ~n61681 ;
  assign n61683 = \pi0247  & ~\pi0527  ;
  assign n61684 = ~n61682 & n61683 ;
  assign n61685 = n60752 & n61422 ;
  assign n61686 = n60754 & n61682 ;
  assign n61687 = ~n61685 & ~n61686 ;
  assign n61688 = ~n61664 & ~n61674 ;
  assign n61689 = \pi0238  & ~n61688 ;
  assign n61690 = ~n61662 & n61689 ;
  assign n61691 = \pi0529  & ~n61690 ;
  assign n61692 = n61687 & n61691 ;
  assign n61693 = ~\pi0238  & ~\pi0491  ;
  assign n61694 = ~n61692 & n61693 ;
  assign n61695 = ~n61684 & n61694 ;
  assign n61696 = ~n61676 & n61695 ;
  assign n61697 = n61667 & n61696 ;
  assign n61698 = n61687 & ~n61690 ;
  assign n61699 = ~\pi0491  & \pi0529  ;
  assign n61700 = ~n61698 & n61699 ;
  assign n61701 = n60779 & n61422 ;
  assign n61702 = n60781 & n61682 ;
  assign n61703 = ~n61701 & ~n61702 ;
  assign n61704 = ~\pi0238  & ~n61688 ;
  assign n61705 = ~n61662 & n61704 ;
  assign n61706 = n61703 & ~n61705 ;
  assign n61707 = \pi0491  & ~\pi0529  ;
  assign n61708 = ~n61706 & n61707 ;
  assign n61709 = ~n61700 & ~n61708 ;
  assign n61710 = ~n61697 & n61709 ;
  assign n61711 = ~\pi0529  & ~n61705 ;
  assign n61712 = n61703 & n61711 ;
  assign n61713 = \pi0238  & \pi0491  ;
  assign n61714 = ~n61712 & n61713 ;
  assign n61715 = ~n61684 & n61714 ;
  assign n61716 = ~n61676 & n61715 ;
  assign n61717 = n61667 & n61716 ;
  assign n61718 = ~n61353 & ~n61717 ;
  assign n61719 = n61710 & n61718 ;
  assign n61720 = ~n61354 & ~n61719 ;
  assign n61721 = ~\pi0237  & ~n61720 ;
  assign n61722 = ~n61116 & ~n61721 ;
  assign n61723 = ~\pi0806  & \pi0990  ;
  assign n61724 = n59494 & n61723 ;
  assign n61725 = ~\pi0332  & \pi0600  ;
  assign n61726 = n61723 & n61725 ;
  assign n61727 = ~\pi0332  & \pi0594  ;
  assign n61728 = ~n61726 & ~n61727 ;
  assign n61729 = ~n61724 & ~n61728 ;
  assign n61730 = \pi0605  & ~\pi0806  ;
  assign n61731 = \pi0595  & n61730 ;
  assign n61732 = n59496 & n61731 ;
  assign n61733 = ~\pi0332  & \pi0595  ;
  assign n61734 = ~\pi0332  & n61730 ;
  assign n61735 = n59496 & n61734 ;
  assign n61736 = ~n61733 & ~n61735 ;
  assign n61737 = ~n61732 & ~n61736 ;
  assign n61738 = ~\pi0332  & \pi0596  ;
  assign n61739 = ~\pi0332  & ~\pi0806  ;
  assign n61740 = \pi0990  & n61739 ;
  assign n61741 = \pi0595  & \pi0597  ;
  assign n61742 = n59494 & n61741 ;
  assign n61743 = n61740 & n61742 ;
  assign n61744 = ~n61738 & ~n61743 ;
  assign n61745 = \pi0596  & \pi0990  ;
  assign n61746 = n61739 & n61745 ;
  assign n61747 = n61742 & n61746 ;
  assign n61748 = ~n61744 & ~n61747 ;
  assign n61749 = ~\pi0332  & \pi0597  ;
  assign n61750 = ~n61724 & n61749 ;
  assign n61751 = ~\pi0332  & ~\pi0597  ;
  assign n61752 = n61724 & n61751 ;
  assign n61753 = ~n61750 & ~n61752 ;
  assign n61754 = ~\pi0057  & \pi0947  ;
  assign n61755 = ~\pi0882  & n61754 ;
  assign n61756 = n6848 & n61755 ;
  assign n61757 = \pi0598  & ~n61756 ;
  assign n61758 = \pi0740  & \pi0780  ;
  assign n61759 = n6712 & n61758 ;
  assign n61760 = ~n61757 & ~n61759 ;
  assign n61761 = ~\pi0332  & \pi0599  ;
  assign n61762 = ~n61747 & ~n61761 ;
  assign n61763 = \pi0599  & n61747 ;
  assign n61764 = ~n61762 & ~n61763 ;
  assign n61765 = ~n61725 & ~n61740 ;
  assign n61766 = ~n61726 & ~n61765 ;
  assign n61767 = ~\pi0601  & \pi0806  ;
  assign n61768 = ~\pi0806  & ~\pi0989  ;
  assign n61769 = ~\pi0332  & ~n61768 ;
  assign n61770 = ~n61767 & n61769 ;
  assign n61771 = ~\pi0230  & \pi0602  ;
  assign n61772 = \pi0230  & ~n23907 ;
  assign n61773 = \pi0790  & n23317 ;
  assign n61774 = ~n23942 & ~n61773 ;
  assign n61775 = n61772 & n61774 ;
  assign n61776 = n23885 & n61775 ;
  assign n61777 = n24915 & n61776 ;
  assign n61778 = ~n61771 & ~n61777 ;
  assign n61779 = ~\pi0980  & \pi1038  ;
  assign n61780 = \pi1060  & n61779 ;
  assign n61781 = \pi0832  & ~\pi1061  ;
  assign n61782 = \pi0952  & n61781 ;
  assign n61783 = n61780 & n61782 ;
  assign n61784 = ~\pi0603  & ~n61783 ;
  assign n61785 = \pi1060  & ~\pi1100  ;
  assign n61786 = n61779 & n61785 ;
  assign n61787 = n61782 & n61786 ;
  assign n61788 = ~\pi0966  & ~n61787 ;
  assign n61789 = ~n61784 & n61788 ;
  assign n61790 = \pi0871  & \pi0966  ;
  assign n61791 = \pi0872  & \pi0966  ;
  assign n61792 = ~n61790 & ~n61791 ;
  assign n61793 = ~n61789 & n61792 ;
  assign n61794 = ~\pi0662  & \pi0823  ;
  assign n61795 = n6708 & n61794 ;
  assign n61796 = ~\pi0779  & n61795 ;
  assign n61797 = ~\pi0299  & \pi0983  ;
  assign n61798 = \pi0907  & n61797 ;
  assign n61799 = \pi0604  & ~n61798 ;
  assign n61800 = ~n61795 & n61799 ;
  assign n61801 = ~n61796 & ~n61800 ;
  assign n61802 = ~\pi0332  & \pi0605  ;
  assign n61803 = ~n61739 & ~n61802 ;
  assign n61804 = ~n61730 & ~n61803 ;
  assign n61805 = \pi1060  & ~\pi1104  ;
  assign n61806 = ~\pi0966  & n61805 ;
  assign n61807 = n61782 & n61806 ;
  assign n61808 = n61779 & n61807 ;
  assign n61809 = ~\pi0606  & ~\pi0966  ;
  assign n61810 = ~n61783 & n61809 ;
  assign n61811 = ~n61808 & ~n61810 ;
  assign n61812 = ~\pi0837  & \pi0966  ;
  assign n61813 = n61811 & ~n61812 ;
  assign n61814 = ~\pi0607  & ~n61783 ;
  assign n61815 = \pi1060  & ~\pi1107  ;
  assign n61816 = n61779 & n61815 ;
  assign n61817 = n61782 & n61816 ;
  assign n61818 = ~\pi0966  & ~n61817 ;
  assign n61819 = ~n61814 & n61818 ;
  assign n61820 = ~\pi0608  & ~n61783 ;
  assign n61821 = \pi1060  & ~\pi1116  ;
  assign n61822 = n61779 & n61821 ;
  assign n61823 = n61782 & n61822 ;
  assign n61824 = ~\pi0966  & ~n61823 ;
  assign n61825 = ~n61820 & n61824 ;
  assign n61826 = ~\pi0609  & ~n61783 ;
  assign n61827 = \pi1060  & ~\pi1118  ;
  assign n61828 = n61779 & n61827 ;
  assign n61829 = n61782 & n61828 ;
  assign n61830 = ~\pi0966  & ~n61829 ;
  assign n61831 = ~n61826 & n61830 ;
  assign n61832 = ~\pi0610  & ~n61783 ;
  assign n61833 = \pi1060  & ~\pi1113  ;
  assign n61834 = n61779 & n61833 ;
  assign n61835 = n61782 & n61834 ;
  assign n61836 = ~\pi0966  & ~n61835 ;
  assign n61837 = ~n61832 & n61836 ;
  assign n61838 = ~\pi0611  & ~n61783 ;
  assign n61839 = \pi1060  & ~\pi1114  ;
  assign n61840 = n61779 & n61839 ;
  assign n61841 = n61782 & n61840 ;
  assign n61842 = ~\pi0966  & ~n61841 ;
  assign n61843 = ~n61838 & n61842 ;
  assign n61844 = ~\pi0612  & ~n61783 ;
  assign n61845 = \pi1060  & ~\pi1111  ;
  assign n61846 = n61779 & n61845 ;
  assign n61847 = n61782 & n61846 ;
  assign n61848 = ~\pi0966  & ~n61847 ;
  assign n61849 = ~n61844 & n61848 ;
  assign n61850 = ~\pi0613  & ~n61783 ;
  assign n61851 = \pi1060  & ~\pi1115  ;
  assign n61852 = n61779 & n61851 ;
  assign n61853 = n61782 & n61852 ;
  assign n61854 = ~\pi0966  & ~n61853 ;
  assign n61855 = ~n61850 & n61854 ;
  assign n61856 = ~\pi0614  & ~n61783 ;
  assign n61857 = \pi1060  & ~\pi1102  ;
  assign n61858 = n61779 & n61857 ;
  assign n61859 = n61782 & n61858 ;
  assign n61860 = ~\pi0966  & ~n61859 ;
  assign n61861 = ~n61856 & n61860 ;
  assign n61862 = ~n61790 & ~n61861 ;
  assign n61863 = ~\pi0057  & \pi0907  ;
  assign n61864 = ~\pi0882  & n61863 ;
  assign n61865 = n6848 & n61864 ;
  assign n61866 = ~\pi0615  & ~n61865 ;
  assign n61867 = \pi0779  & \pi0797  ;
  assign n61868 = n6709 & n61867 ;
  assign n61869 = ~n61866 & ~n61868 ;
  assign n61870 = ~\pi0616  & ~n61783 ;
  assign n61871 = \pi1060  & ~\pi1101  ;
  assign n61872 = n61779 & n61871 ;
  assign n61873 = n61782 & n61872 ;
  assign n61874 = ~\pi0966  & ~n61873 ;
  assign n61875 = ~n61870 & n61874 ;
  assign n61876 = ~n61791 & ~n61875 ;
  assign n61877 = \pi1060  & ~\pi1105  ;
  assign n61878 = ~\pi0966  & n61877 ;
  assign n61879 = n61782 & n61878 ;
  assign n61880 = n61779 & n61879 ;
  assign n61881 = ~\pi0617  & ~\pi0966  ;
  assign n61882 = ~n61783 & n61881 ;
  assign n61883 = ~n61880 & ~n61882 ;
  assign n61884 = ~\pi0850  & \pi0966  ;
  assign n61885 = n61883 & ~n61884 ;
  assign n61886 = ~\pi0618  & ~n61783 ;
  assign n61887 = \pi1060  & ~\pi1117  ;
  assign n61888 = n61779 & n61887 ;
  assign n61889 = n61782 & n61888 ;
  assign n61890 = ~\pi0966  & ~n61889 ;
  assign n61891 = ~n61886 & n61890 ;
  assign n61892 = ~\pi0619  & ~n61783 ;
  assign n61893 = \pi1060  & ~\pi1122  ;
  assign n61894 = n61779 & n61893 ;
  assign n61895 = n61782 & n61894 ;
  assign n61896 = ~\pi0966  & ~n61895 ;
  assign n61897 = ~n61892 & n61896 ;
  assign n61898 = ~\pi0620  & ~n61783 ;
  assign n61899 = \pi1060  & ~\pi1112  ;
  assign n61900 = n61779 & n61899 ;
  assign n61901 = n61782 & n61900 ;
  assign n61902 = ~\pi0966  & ~n61901 ;
  assign n61903 = ~n61898 & n61902 ;
  assign n61904 = ~\pi0621  & ~n61783 ;
  assign n61905 = \pi1060  & ~\pi1108  ;
  assign n61906 = n61779 & n61905 ;
  assign n61907 = n61782 & n61906 ;
  assign n61908 = ~\pi0966  & ~n61907 ;
  assign n61909 = ~n61904 & n61908 ;
  assign n61910 = ~\pi0622  & ~n61783 ;
  assign n61911 = \pi1060  & ~\pi1109  ;
  assign n61912 = n61779 & n61911 ;
  assign n61913 = n61782 & n61912 ;
  assign n61914 = ~\pi0966  & ~n61913 ;
  assign n61915 = ~n61910 & n61914 ;
  assign n61916 = ~\pi0623  & ~n61783 ;
  assign n61917 = \pi1060  & ~\pi1106  ;
  assign n61918 = n61779 & n61917 ;
  assign n61919 = n61782 & n61918 ;
  assign n61920 = ~\pi0966  & ~n61919 ;
  assign n61921 = ~n61916 & n61920 ;
  assign n61922 = ~\pi0616  & \pi0831  ;
  assign n61923 = n21369 & n61922 ;
  assign n61924 = ~\pi0780  & n61923 ;
  assign n61925 = \pi0947  & n61797 ;
  assign n61926 = \pi0624  & ~n61925 ;
  assign n61927 = ~n61923 & n61926 ;
  assign n61928 = ~n61924 & ~n61927 ;
  assign n61929 = ~\pi1054  & \pi1066  ;
  assign n61930 = \pi1088  & n61929 ;
  assign n61931 = \pi0832  & ~\pi0973  ;
  assign n61932 = ~\pi0953  & n61931 ;
  assign n61933 = n61930 & n61932 ;
  assign n61934 = ~\pi0625  & ~n61933 ;
  assign n61935 = ~\pi0953  & ~\pi1116  ;
  assign n61936 = n61931 & n61935 ;
  assign n61937 = n61930 & n61936 ;
  assign n61938 = ~\pi0962  & ~n61937 ;
  assign n61939 = ~n61934 & n61938 ;
  assign n61940 = ~\pi0626  & ~n61783 ;
  assign n61941 = \pi1060  & ~\pi1121  ;
  assign n61942 = n61779 & n61941 ;
  assign n61943 = n61782 & n61942 ;
  assign n61944 = ~\pi0966  & ~n61943 ;
  assign n61945 = ~n61940 & n61944 ;
  assign n61946 = ~\pi0627  & ~n61933 ;
  assign n61947 = ~\pi0953  & ~\pi1117  ;
  assign n61948 = n61931 & n61947 ;
  assign n61949 = n61930 & n61948 ;
  assign n61950 = ~\pi0962  & ~n61949 ;
  assign n61951 = ~n61946 & n61950 ;
  assign n61952 = ~\pi0628  & ~n61933 ;
  assign n61953 = ~\pi0953  & ~\pi1119  ;
  assign n61954 = n61931 & n61953 ;
  assign n61955 = n61930 & n61954 ;
  assign n61956 = ~\pi0962  & ~n61955 ;
  assign n61957 = ~n61952 & n61956 ;
  assign n61958 = ~\pi0629  & ~n61783 ;
  assign n61959 = \pi1060  & ~\pi1119  ;
  assign n61960 = n61779 & n61959 ;
  assign n61961 = n61782 & n61960 ;
  assign n61962 = ~\pi0966  & ~n61961 ;
  assign n61963 = ~n61958 & n61962 ;
  assign n61964 = ~\pi0630  & ~n61783 ;
  assign n61965 = \pi1060  & ~\pi1120  ;
  assign n61966 = n61779 & n61965 ;
  assign n61967 = n61782 & n61966 ;
  assign n61968 = ~\pi0966  & ~n61967 ;
  assign n61969 = ~n61964 & n61968 ;
  assign n61970 = \pi0631  & ~n61933 ;
  assign n61971 = ~\pi0953  & ~\pi1113  ;
  assign n61972 = n61931 & n61971 ;
  assign n61973 = n61930 & n61972 ;
  assign n61974 = ~\pi0962  & ~n61973 ;
  assign n61975 = ~n61970 & n61974 ;
  assign n61976 = \pi0632  & ~n61933 ;
  assign n61977 = ~\pi0953  & ~\pi1115  ;
  assign n61978 = n61931 & n61977 ;
  assign n61979 = n61930 & n61978 ;
  assign n61980 = ~\pi0962  & ~n61979 ;
  assign n61981 = ~n61976 & n61980 ;
  assign n61982 = ~\pi0633  & ~n61783 ;
  assign n61983 = \pi1060  & ~\pi1110  ;
  assign n61984 = n61779 & n61983 ;
  assign n61985 = n61782 & n61984 ;
  assign n61986 = ~\pi0966  & ~n61985 ;
  assign n61987 = ~n61982 & n61986 ;
  assign n61988 = ~\pi0634  & ~n61933 ;
  assign n61989 = ~\pi0953  & ~\pi1110  ;
  assign n61990 = n61931 & n61989 ;
  assign n61991 = n61930 & n61990 ;
  assign n61992 = ~\pi0962  & ~n61991 ;
  assign n61993 = ~n61988 & n61992 ;
  assign n61994 = \pi0635  & ~n61933 ;
  assign n61995 = ~\pi0953  & ~\pi1112  ;
  assign n61996 = n61931 & n61995 ;
  assign n61997 = n61930 & n61996 ;
  assign n61998 = ~\pi0962  & ~n61997 ;
  assign n61999 = ~n61994 & n61998 ;
  assign n62000 = ~\pi0636  & ~n61783 ;
  assign n62001 = \pi1060  & ~\pi1127  ;
  assign n62002 = n61779 & n62001 ;
  assign n62003 = n61782 & n62002 ;
  assign n62004 = ~\pi0966  & ~n62003 ;
  assign n62005 = ~n62000 & n62004 ;
  assign n62006 = ~\pi0637  & ~n61933 ;
  assign n62007 = ~\pi0953  & ~\pi1105  ;
  assign n62008 = n61931 & n62007 ;
  assign n62009 = n61930 & n62008 ;
  assign n62010 = ~\pi0962  & ~n62009 ;
  assign n62011 = ~n62006 & n62010 ;
  assign n62012 = ~\pi0638  & ~n61933 ;
  assign n62013 = ~\pi0953  & ~\pi1107  ;
  assign n62014 = n61931 & n62013 ;
  assign n62015 = n61930 & n62014 ;
  assign n62016 = ~\pi0962  & ~n62015 ;
  assign n62017 = ~n62012 & n62016 ;
  assign n62018 = ~\pi0639  & ~n61933 ;
  assign n62019 = ~\pi0953  & ~\pi1109  ;
  assign n62020 = n61931 & n62019 ;
  assign n62021 = n61930 & n62020 ;
  assign n62022 = ~\pi0962  & ~n62021 ;
  assign n62023 = ~n62018 & n62022 ;
  assign n62024 = ~\pi0640  & ~n61783 ;
  assign n62025 = \pi1060  & ~\pi1128  ;
  assign n62026 = n61779 & n62025 ;
  assign n62027 = n61782 & n62026 ;
  assign n62028 = ~\pi0966  & ~n62027 ;
  assign n62029 = ~n62024 & n62028 ;
  assign n62030 = ~\pi0641  & ~n61933 ;
  assign n62031 = ~\pi0953  & ~\pi1121  ;
  assign n62032 = n61931 & n62031 ;
  assign n62033 = n61930 & n62032 ;
  assign n62034 = ~\pi0962  & ~n62033 ;
  assign n62035 = ~n62030 & n62034 ;
  assign n62036 = ~\pi0642  & ~n61783 ;
  assign n62037 = \pi1060  & ~\pi1103  ;
  assign n62038 = n61779 & n62037 ;
  assign n62039 = n61782 & n62038 ;
  assign n62040 = ~\pi0966  & ~n62039 ;
  assign n62041 = ~n62036 & n62040 ;
  assign n62042 = ~\pi0643  & ~n61933 ;
  assign n62043 = ~\pi0953  & ~\pi1104  ;
  assign n62044 = n61931 & n62043 ;
  assign n62045 = n61930 & n62044 ;
  assign n62046 = ~\pi0962  & ~n62045 ;
  assign n62047 = ~n62042 & n62046 ;
  assign n62048 = ~\pi0644  & ~n61783 ;
  assign n62049 = \pi1060  & ~\pi1123  ;
  assign n62050 = n61779 & n62049 ;
  assign n62051 = n61782 & n62050 ;
  assign n62052 = ~\pi0966  & ~n62051 ;
  assign n62053 = ~n62048 & n62052 ;
  assign n62054 = ~\pi0645  & ~n61783 ;
  assign n62055 = \pi1060  & ~\pi1125  ;
  assign n62056 = n61779 & n62055 ;
  assign n62057 = n61782 & n62056 ;
  assign n62058 = ~\pi0966  & ~n62057 ;
  assign n62059 = ~n62054 & n62058 ;
  assign n62060 = \pi0646  & ~n61933 ;
  assign n62061 = ~\pi0953  & ~\pi1114  ;
  assign n62062 = n61931 & n62061 ;
  assign n62063 = n61930 & n62062 ;
  assign n62064 = ~\pi0962  & ~n62063 ;
  assign n62065 = ~n62060 & n62064 ;
  assign n62066 = ~\pi0647  & ~n61933 ;
  assign n62067 = ~\pi0953  & ~\pi1120  ;
  assign n62068 = n61931 & n62067 ;
  assign n62069 = n61930 & n62068 ;
  assign n62070 = ~\pi0962  & ~n62069 ;
  assign n62071 = ~n62066 & n62070 ;
  assign n62072 = ~\pi0648  & ~n61933 ;
  assign n62073 = ~\pi0953  & ~\pi1122  ;
  assign n62074 = n61931 & n62073 ;
  assign n62075 = n61930 & n62074 ;
  assign n62076 = ~\pi0962  & ~n62075 ;
  assign n62077 = ~n62072 & n62076 ;
  assign n62078 = \pi0649  & ~n61933 ;
  assign n62079 = ~\pi0953  & ~\pi1126  ;
  assign n62080 = n61931 & n62079 ;
  assign n62081 = n61930 & n62080 ;
  assign n62082 = ~\pi0962  & ~n62081 ;
  assign n62083 = ~n62078 & n62082 ;
  assign n62084 = \pi0650  & ~n61933 ;
  assign n62085 = ~\pi0953  & ~\pi1127  ;
  assign n62086 = n61931 & n62085 ;
  assign n62087 = n61930 & n62086 ;
  assign n62088 = ~\pi0962  & ~n62087 ;
  assign n62089 = ~n62084 & n62088 ;
  assign n62090 = ~\pi0651  & ~n61783 ;
  assign n62091 = \pi1060  & ~\pi1130  ;
  assign n62092 = n61779 & n62091 ;
  assign n62093 = n61782 & n62092 ;
  assign n62094 = ~\pi0966  & ~n62093 ;
  assign n62095 = ~n62090 & n62094 ;
  assign n62096 = ~\pi0652  & ~n61783 ;
  assign n62097 = \pi1060  & ~\pi1131  ;
  assign n62098 = n61779 & n62097 ;
  assign n62099 = n61782 & n62098 ;
  assign n62100 = ~\pi0966  & ~n62099 ;
  assign n62101 = ~n62096 & n62100 ;
  assign n62102 = ~\pi0653  & ~n61783 ;
  assign n62103 = \pi1060  & ~\pi1129  ;
  assign n62104 = n61779 & n62103 ;
  assign n62105 = n61782 & n62104 ;
  assign n62106 = ~\pi0966  & ~n62105 ;
  assign n62107 = ~n62102 & n62106 ;
  assign n62108 = \pi0654  & ~n61933 ;
  assign n62109 = ~\pi0953  & ~\pi1130  ;
  assign n62110 = n61931 & n62109 ;
  assign n62111 = n61930 & n62110 ;
  assign n62112 = ~\pi0962  & ~n62111 ;
  assign n62113 = ~n62108 & n62112 ;
  assign n62114 = \pi0655  & ~n61933 ;
  assign n62115 = ~\pi0953  & ~\pi1124  ;
  assign n62116 = n61931 & n62115 ;
  assign n62117 = n61930 & n62116 ;
  assign n62118 = ~\pi0962  & ~n62117 ;
  assign n62119 = ~n62114 & n62118 ;
  assign n62120 = ~\pi0656  & ~n61783 ;
  assign n62121 = \pi1060  & ~\pi1126  ;
  assign n62122 = n61779 & n62121 ;
  assign n62123 = n61782 & n62122 ;
  assign n62124 = ~\pi0966  & ~n62123 ;
  assign n62125 = ~n62120 & n62124 ;
  assign n62126 = \pi0657  & ~n61933 ;
  assign n62127 = ~\pi0953  & ~\pi1131  ;
  assign n62128 = n61931 & n62127 ;
  assign n62129 = n61930 & n62128 ;
  assign n62130 = ~\pi0962  & ~n62129 ;
  assign n62131 = ~n62126 & n62130 ;
  assign n62132 = ~\pi0658  & ~n61783 ;
  assign n62133 = \pi1060  & ~\pi1124  ;
  assign n62134 = n61779 & n62133 ;
  assign n62135 = n61782 & n62134 ;
  assign n62136 = ~\pi0966  & ~n62135 ;
  assign n62137 = ~n62132 & n62136 ;
  assign n62138 = \pi0266  & \pi0992  ;
  assign n62139 = ~\pi0269  & ~\pi0280  ;
  assign n62140 = n62138 & n62139 ;
  assign n62141 = ~\pi0270  & ~\pi0277  ;
  assign n62142 = ~\pi0281  & ~\pi0282  ;
  assign n62143 = n62141 & n62142 ;
  assign n62144 = ~\pi0264  & ~\pi0274  ;
  assign n62145 = ~\pi0265  & n62144 ;
  assign n62146 = n62143 & n62145 ;
  assign n62147 = n62140 & n62146 ;
  assign n62148 = n62140 & n62143 ;
  assign n62149 = ~\pi0264  & ~\pi0265  ;
  assign n62150 = n62148 & n62149 ;
  assign n62151 = \pi0274  & ~n62150 ;
  assign n62152 = ~n62147 & ~n62151 ;
  assign n62153 = ~\pi0660  & ~n61933 ;
  assign n62154 = ~\pi0953  & ~\pi1118  ;
  assign n62155 = n61931 & n62154 ;
  assign n62156 = n61930 & n62155 ;
  assign n62157 = ~\pi0962  & ~n62156 ;
  assign n62158 = ~n62153 & n62157 ;
  assign n62159 = ~\pi0661  & ~n61933 ;
  assign n62160 = ~\pi0953  & ~\pi1101  ;
  assign n62161 = n61931 & n62160 ;
  assign n62162 = n61930 & n62161 ;
  assign n62163 = ~\pi0962  & ~n62162 ;
  assign n62164 = ~n62159 & n62163 ;
  assign n62165 = ~\pi0662  & ~n61933 ;
  assign n62166 = ~\pi0953  & ~\pi1102  ;
  assign n62167 = n61931 & n62166 ;
  assign n62168 = n61930 & n62167 ;
  assign n62169 = ~\pi0962  & ~n62168 ;
  assign n62170 = ~n62165 & n62169 ;
  assign n62171 = ~\pi0591  & \pi0592  ;
  assign n62172 = \pi0365  & n62171 ;
  assign n62173 = \pi0334  & \pi0591  ;
  assign n62174 = ~\pi0592  & n62173 ;
  assign n62175 = ~n62172 & ~n62174 ;
  assign n62176 = ~\pi0590  & ~n62175 ;
  assign n62177 = \pi0199  & ~\pi1065  ;
  assign n62178 = ~\pi0223  & ~\pi0224  ;
  assign n62179 = ~\pi0199  & ~\pi0257  ;
  assign n62180 = ~n62178 & ~n62179 ;
  assign n62181 = ~n62177 & n62180 ;
  assign n62182 = \pi0590  & ~\pi0591  ;
  assign n62183 = \pi0323  & ~\pi0592  ;
  assign n62184 = n62182 & n62183 ;
  assign n62185 = ~\pi0588  & ~n62184 ;
  assign n62186 = ~n62181 & n62185 ;
  assign n62187 = ~n62176 & n62186 ;
  assign n62188 = n10003 & n62181 ;
  assign n62189 = \pi0464  & ~\pi0592  ;
  assign n62190 = n9927 & n62189 ;
  assign n62191 = \pi0588  & ~n62190 ;
  assign n62192 = n10003 & n62178 ;
  assign n62193 = ~n62191 & n62192 ;
  assign n62194 = ~n62188 & ~n62193 ;
  assign n62195 = ~n62187 & ~n62194 ;
  assign n62196 = ~\pi1137  & ~\pi1138  ;
  assign n62197 = ~\pi1134  & n62196 ;
  assign n62198 = ~\pi0634  & \pi1136  ;
  assign n62199 = ~\pi0784  & ~\pi1136  ;
  assign n62200 = \pi1135  & ~n62199 ;
  assign n62201 = ~n62198 & n62200 ;
  assign n62202 = ~\pi0633  & \pi1136  ;
  assign n62203 = ~\pi0815  & ~\pi1136  ;
  assign n62204 = ~\pi1135  & ~n62203 ;
  assign n62205 = ~n62202 & n62204 ;
  assign n62206 = ~n62201 & ~n62205 ;
  assign n62207 = n62197 & ~n62206 ;
  assign n62208 = \pi1135  & ~\pi1136  ;
  assign n62209 = \pi1134  & n62196 ;
  assign n62210 = ~n62208 & n62209 ;
  assign n62211 = \pi1135  & n62196 ;
  assign n62212 = ~\pi0766  & \pi1136  ;
  assign n62213 = ~n62211 & n62212 ;
  assign n62214 = ~\pi0855  & ~\pi1136  ;
  assign n62215 = ~\pi0700  & \pi1135  ;
  assign n62216 = ~n62214 & ~n62215 ;
  assign n62217 = ~n62213 & n62216 ;
  assign n62218 = n62210 & n62217 ;
  assign n62219 = ~n62207 & ~n62218 ;
  assign n62220 = ~n10003 & ~n62219 ;
  assign n62221 = ~n62195 & ~n62220 ;
  assign n62222 = \pi0404  & n15247 ;
  assign n62223 = ~\pi0590  & \pi0592  ;
  assign n62224 = ~\pi0588  & ~n62223 ;
  assign n62225 = ~n62222 & n62224 ;
  assign n62226 = \pi0380  & ~\pi0591  ;
  assign n62227 = \pi0592  & ~n62226 ;
  assign n62228 = ~n62225 & ~n62227 ;
  assign n62229 = \pi0199  & ~\pi1084  ;
  assign n62230 = ~\pi0199  & ~\pi0292  ;
  assign n62231 = ~n62178 & ~n62230 ;
  assign n62232 = ~n62229 & n62231 ;
  assign n62233 = \pi0355  & ~\pi0592  ;
  assign n62234 = n62182 & n62233 ;
  assign n62235 = ~n62232 & ~n62234 ;
  assign n62236 = ~n62228 & n62235 ;
  assign n62237 = n10003 & n62232 ;
  assign n62238 = \pi0429  & ~\pi0592  ;
  assign n62239 = n9927 & n62238 ;
  assign n62240 = \pi0588  & ~n62239 ;
  assign n62241 = n62192 & ~n62240 ;
  assign n62242 = ~n62237 & ~n62241 ;
  assign n62243 = ~n62236 & ~n62242 ;
  assign n62244 = \pi0785  & \pi1135  ;
  assign n62245 = \pi0811  & ~\pi1135  ;
  assign n62246 = ~n62244 & ~n62245 ;
  assign n62247 = ~\pi1136  & n62246 ;
  assign n62248 = \pi0662  & \pi1135  ;
  assign n62249 = \pi0614  & ~\pi1135  ;
  assign n62250 = \pi1136  & ~n62249 ;
  assign n62251 = ~n62248 & n62250 ;
  assign n62252 = ~n62247 & ~n62251 ;
  assign n62253 = ~\pi1134  & ~n62252 ;
  assign n62254 = ~\pi0727  & \pi1135  ;
  assign n62255 = ~\pi0772  & ~\pi1135  ;
  assign n62256 = ~n62254 & ~n62255 ;
  assign n62257 = \pi1136  & n62256 ;
  assign n62258 = ~\pi1135  & ~\pi1136  ;
  assign n62259 = \pi0872  & n62258 ;
  assign n62260 = \pi1134  & ~n62259 ;
  assign n62261 = ~n62257 & n62260 ;
  assign n62262 = ~n10003 & n62196 ;
  assign n62263 = ~n62261 & n62262 ;
  assign n62264 = ~n62253 & n62263 ;
  assign n62265 = ~n62243 & ~n62264 ;
  assign n62266 = ~\pi0665  & ~n61933 ;
  assign n62267 = ~\pi0953  & ~\pi1108  ;
  assign n62268 = n61931 & n62267 ;
  assign n62269 = n61930 & n62268 ;
  assign n62270 = ~\pi0962  & ~n62269 ;
  assign n62271 = ~n62266 & n62270 ;
  assign n62272 = ~\pi0638  & \pi1135  ;
  assign n62273 = ~\pi0607  & ~\pi1135  ;
  assign n62274 = ~n62272 & ~n62273 ;
  assign n62275 = \pi1136  & n62274 ;
  assign n62276 = \pi0799  & ~\pi1135  ;
  assign n62277 = ~\pi0790  & \pi1135  ;
  assign n62278 = ~n62276 & ~n62277 ;
  assign n62279 = ~\pi1136  & n62278 ;
  assign n62280 = ~n62275 & ~n62279 ;
  assign n62281 = n62197 & ~n62280 ;
  assign n62282 = ~\pi0764  & \pi1136  ;
  assign n62283 = ~n62211 & n62282 ;
  assign n62284 = ~\pi0691  & \pi1135  ;
  assign n62285 = ~\pi0873  & ~\pi1136  ;
  assign n62286 = ~n62284 & ~n62285 ;
  assign n62287 = ~n62283 & n62286 ;
  assign n62288 = n62210 & n62287 ;
  assign n62289 = ~n62281 & ~n62288 ;
  assign n62290 = ~n10003 & ~n62289 ;
  assign n62291 = \pi0456  & n15247 ;
  assign n62292 = n62224 & ~n62291 ;
  assign n62293 = \pi0337  & ~\pi0591  ;
  assign n62294 = \pi0592  & ~n62293 ;
  assign n62295 = ~n62292 & ~n62294 ;
  assign n62296 = \pi0199  & ~\pi1044  ;
  assign n62297 = ~\pi0199  & ~\pi0297  ;
  assign n62298 = ~n62178 & ~n62297 ;
  assign n62299 = ~n62296 & n62298 ;
  assign n62300 = \pi0441  & ~\pi0592  ;
  assign n62301 = n62182 & n62300 ;
  assign n62302 = ~n62299 & ~n62301 ;
  assign n62303 = ~n62295 & n62302 ;
  assign n62304 = n10003 & n62299 ;
  assign n62305 = \pi0443  & ~\pi0592  ;
  assign n62306 = n9927 & n62305 ;
  assign n62307 = \pi0588  & ~n62306 ;
  assign n62308 = n62192 & ~n62307 ;
  assign n62309 = ~n62304 & ~n62308 ;
  assign n62310 = ~n62303 & ~n62309 ;
  assign n62311 = ~n62290 & ~n62310 ;
  assign n62312 = \pi0319  & n15247 ;
  assign n62313 = n62224 & ~n62312 ;
  assign n62314 = \pi0338  & ~\pi0591  ;
  assign n62315 = \pi0592  & ~n62314 ;
  assign n62316 = ~n62313 & ~n62315 ;
  assign n62317 = \pi0199  & ~\pi1072  ;
  assign n62318 = ~\pi0199  & ~\pi0294  ;
  assign n62319 = ~n62178 & ~n62318 ;
  assign n62320 = ~n62317 & n62319 ;
  assign n62321 = \pi0458  & ~\pi0592  ;
  assign n62322 = n62182 & n62321 ;
  assign n62323 = ~n62320 & ~n62322 ;
  assign n62324 = ~n62316 & n62323 ;
  assign n62325 = n10003 & n62320 ;
  assign n62326 = \pi0444  & ~\pi0592  ;
  assign n62327 = n9927 & n62326 ;
  assign n62328 = \pi0588  & ~n62327 ;
  assign n62329 = n62192 & ~n62328 ;
  assign n62330 = ~n62325 & ~n62329 ;
  assign n62331 = ~n62324 & ~n62330 ;
  assign n62332 = \pi0681  & \pi1136  ;
  assign n62333 = \pi0792  & ~\pi1136  ;
  assign n62334 = \pi1135  & ~n62333 ;
  assign n62335 = ~n62332 & n62334 ;
  assign n62336 = \pi0642  & \pi1136  ;
  assign n62337 = ~\pi0809  & ~\pi1136  ;
  assign n62338 = ~\pi1135  & ~n62337 ;
  assign n62339 = ~n62336 & n62338 ;
  assign n62340 = ~n62335 & ~n62339 ;
  assign n62341 = ~\pi1134  & ~n62340 ;
  assign n62342 = ~\pi0699  & \pi1135  ;
  assign n62343 = ~\pi0763  & ~\pi1135  ;
  assign n62344 = ~n62342 & ~n62343 ;
  assign n62345 = \pi1136  & n62344 ;
  assign n62346 = \pi0871  & n62258 ;
  assign n62347 = \pi1134  & ~n62346 ;
  assign n62348 = ~n62345 & n62347 ;
  assign n62349 = n62262 & ~n62348 ;
  assign n62350 = ~n62341 & n62349 ;
  assign n62351 = ~n62331 & ~n62350 ;
  assign n62352 = ~\pi0680  & \pi1135  ;
  assign n62353 = ~\pi0603  & ~\pi1135  ;
  assign n62354 = ~n62352 & ~n62353 ;
  assign n62355 = \pi1136  & n62354 ;
  assign n62356 = ~\pi0778  & \pi1135  ;
  assign n62357 = ~\pi0981  & ~\pi1135  ;
  assign n62358 = ~n62356 & ~n62357 ;
  assign n62359 = ~\pi1136  & n62358 ;
  assign n62360 = ~n62355 & ~n62359 ;
  assign n62361 = n62197 & ~n62360 ;
  assign n62362 = ~\pi0759  & \pi1136  ;
  assign n62363 = ~n62211 & n62362 ;
  assign n62364 = ~\pi0696  & \pi1135  ;
  assign n62365 = ~\pi0837  & ~\pi1136  ;
  assign n62366 = ~n62364 & ~n62365 ;
  assign n62367 = ~n62363 & n62366 ;
  assign n62368 = n62210 & n62367 ;
  assign n62369 = ~n62361 & ~n62368 ;
  assign n62370 = ~n10003 & ~n62369 ;
  assign n62371 = \pi0390  & n15247 ;
  assign n62372 = n62224 & ~n62371 ;
  assign n62373 = \pi0363  & ~\pi0591  ;
  assign n62374 = \pi0592  & ~n62373 ;
  assign n62375 = ~n62372 & ~n62374 ;
  assign n62376 = \pi0199  & ~\pi1049  ;
  assign n62377 = ~\pi0199  & ~\pi0291  ;
  assign n62378 = ~n62178 & ~n62377 ;
  assign n62379 = ~n62376 & n62378 ;
  assign n62380 = \pi0342  & ~\pi0592  ;
  assign n62381 = n62182 & n62380 ;
  assign n62382 = ~n62379 & ~n62381 ;
  assign n62383 = ~n62375 & n62382 ;
  assign n62384 = n10003 & n62379 ;
  assign n62385 = \pi0414  & ~\pi0592  ;
  assign n62386 = n9927 & n62385 ;
  assign n62387 = \pi0588  & ~n62386 ;
  assign n62388 = n62192 & ~n62387 ;
  assign n62389 = ~n62384 & ~n62388 ;
  assign n62390 = ~n62383 & ~n62389 ;
  assign n62391 = ~n62370 & ~n62390 ;
  assign n62392 = \pi0669  & ~n61933 ;
  assign n62393 = ~\pi0953  & ~\pi1125  ;
  assign n62394 = n61931 & n62393 ;
  assign n62395 = n61930 & n62394 ;
  assign n62396 = ~\pi0962  & ~n62395 ;
  assign n62397 = ~n62392 & n62396 ;
  assign n62398 = \pi0364  & n62171 ;
  assign n62399 = \pi0391  & \pi0591  ;
  assign n62400 = ~\pi0592  & n62399 ;
  assign n62401 = ~n62398 & ~n62400 ;
  assign n62402 = ~\pi0590  & ~n62401 ;
  assign n62403 = \pi0199  & ~\pi1062  ;
  assign n62404 = ~\pi0199  & ~\pi0258  ;
  assign n62405 = ~n62178 & ~n62404 ;
  assign n62406 = ~n62403 & n62405 ;
  assign n62407 = \pi0343  & ~\pi0592  ;
  assign n62408 = n62182 & n62407 ;
  assign n62409 = ~\pi0588  & ~n62408 ;
  assign n62410 = ~n62406 & n62409 ;
  assign n62411 = ~n62402 & n62410 ;
  assign n62412 = n10003 & n62406 ;
  assign n62413 = \pi0415  & ~\pi0592  ;
  assign n62414 = n9927 & n62413 ;
  assign n62415 = \pi0588  & ~n62414 ;
  assign n62416 = n62192 & ~n62415 ;
  assign n62417 = ~n62412 & ~n62416 ;
  assign n62418 = ~n62411 & ~n62417 ;
  assign n62419 = \pi0695  & \pi1135  ;
  assign n62420 = ~\pi1134  & ~n62419 ;
  assign n62421 = ~\pi0612  & ~\pi1135  ;
  assign n62422 = \pi1136  & ~n62421 ;
  assign n62423 = n62420 & n62422 ;
  assign n62424 = n62262 & n62423 ;
  assign n62425 = \pi0723  & \pi1135  ;
  assign n62426 = ~\pi0852  & ~\pi1136  ;
  assign n62427 = ~n62425 & ~n62426 ;
  assign n62428 = n62210 & n62427 ;
  assign n62429 = \pi0745  & \pi1136  ;
  assign n62430 = ~n62211 & n62429 ;
  assign n62431 = ~n10003 & ~n62430 ;
  assign n62432 = n62428 & n62431 ;
  assign n62433 = ~n62424 & ~n62432 ;
  assign n62434 = ~n62418 & n62433 ;
  assign n62435 = \pi0447  & n62171 ;
  assign n62436 = \pi0333  & \pi0591  ;
  assign n62437 = ~\pi0592  & n62436 ;
  assign n62438 = ~n62435 & ~n62437 ;
  assign n62439 = ~\pi0590  & ~n62438 ;
  assign n62440 = \pi0199  & ~\pi1040  ;
  assign n62441 = ~\pi0199  & ~\pi0261  ;
  assign n62442 = ~n62178 & ~n62441 ;
  assign n62443 = ~n62440 & n62442 ;
  assign n62444 = \pi0327  & ~\pi0592  ;
  assign n62445 = n62182 & n62444 ;
  assign n62446 = ~\pi0588  & ~n62445 ;
  assign n62447 = ~n62443 & n62446 ;
  assign n62448 = ~n62439 & n62447 ;
  assign n62449 = n10003 & n62443 ;
  assign n62450 = \pi0453  & ~\pi0592  ;
  assign n62451 = n9927 & n62450 ;
  assign n62452 = \pi0588  & ~n62451 ;
  assign n62453 = n62192 & ~n62452 ;
  assign n62454 = ~n62449 & ~n62453 ;
  assign n62455 = ~n62448 & ~n62454 ;
  assign n62456 = \pi0646  & \pi1135  ;
  assign n62457 = ~\pi1134  & ~n62456 ;
  assign n62458 = ~\pi0611  & ~\pi1135  ;
  assign n62459 = \pi1136  & ~n62458 ;
  assign n62460 = n62457 & n62459 ;
  assign n62461 = n62262 & n62460 ;
  assign n62462 = \pi0724  & \pi1135  ;
  assign n62463 = ~\pi0865  & ~\pi1136  ;
  assign n62464 = ~n62462 & ~n62463 ;
  assign n62465 = n62210 & n62464 ;
  assign n62466 = \pi0741  & \pi1136  ;
  assign n62467 = ~n62211 & n62466 ;
  assign n62468 = ~n10003 & ~n62467 ;
  assign n62469 = n62465 & n62468 ;
  assign n62470 = ~n62461 & ~n62469 ;
  assign n62471 = ~n62455 & n62470 ;
  assign n62472 = ~\pi0661  & \pi1135  ;
  assign n62473 = ~\pi0616  & ~\pi1135  ;
  assign n62474 = ~n62472 & ~n62473 ;
  assign n62475 = \pi1136  & n62474 ;
  assign n62476 = ~\pi0781  & \pi1135  ;
  assign n62477 = ~\pi0808  & ~\pi1135  ;
  assign n62478 = ~n62476 & ~n62477 ;
  assign n62479 = ~\pi1136  & n62478 ;
  assign n62480 = ~n62475 & ~n62479 ;
  assign n62481 = n62197 & ~n62480 ;
  assign n62482 = ~\pi0758  & \pi1136  ;
  assign n62483 = ~n62211 & n62482 ;
  assign n62484 = ~\pi0736  & \pi1135  ;
  assign n62485 = ~\pi0850  & ~\pi1136  ;
  assign n62486 = ~n62484 & ~n62485 ;
  assign n62487 = ~n62483 & n62486 ;
  assign n62488 = n62210 & n62487 ;
  assign n62489 = ~n62481 & ~n62488 ;
  assign n62490 = ~n10003 & ~n62489 ;
  assign n62491 = \pi0397  & n15247 ;
  assign n62492 = n62224 & ~n62491 ;
  assign n62493 = \pi0372  & ~\pi0591  ;
  assign n62494 = \pi0592  & ~n62493 ;
  assign n62495 = ~n62492 & ~n62494 ;
  assign n62496 = \pi0199  & ~\pi1048  ;
  assign n62497 = ~\pi0199  & ~\pi0290  ;
  assign n62498 = ~n62178 & ~n62497 ;
  assign n62499 = ~n62496 & n62498 ;
  assign n62500 = \pi0320  & ~\pi0592  ;
  assign n62501 = n62182 & n62500 ;
  assign n62502 = ~n62499 & ~n62501 ;
  assign n62503 = ~n62495 & n62502 ;
  assign n62504 = n10003 & n62499 ;
  assign n62505 = \pi0422  & ~\pi0592  ;
  assign n62506 = n9927 & n62505 ;
  assign n62507 = \pi0588  & ~n62506 ;
  assign n62508 = n62192 & ~n62507 ;
  assign n62509 = ~n62504 & ~n62508 ;
  assign n62510 = ~n62503 & ~n62509 ;
  assign n62511 = ~n62490 & ~n62510 ;
  assign n62512 = ~\pi0637  & \pi1135  ;
  assign n62513 = ~\pi0617  & ~\pi1135  ;
  assign n62514 = ~n62512 & ~n62513 ;
  assign n62515 = \pi1136  & n62514 ;
  assign n62516 = \pi0814  & ~\pi1135  ;
  assign n62517 = ~\pi0788  & \pi1135  ;
  assign n62518 = ~n62516 & ~n62517 ;
  assign n62519 = ~\pi1136  & n62518 ;
  assign n62520 = ~n62515 & ~n62519 ;
  assign n62521 = n62197 & ~n62520 ;
  assign n62522 = ~\pi0749  & \pi1136  ;
  assign n62523 = ~n62211 & n62522 ;
  assign n62524 = ~\pi0706  & \pi1135  ;
  assign n62525 = ~\pi0866  & ~\pi1136  ;
  assign n62526 = ~n62524 & ~n62525 ;
  assign n62527 = ~n62523 & n62526 ;
  assign n62528 = n62210 & n62527 ;
  assign n62529 = ~n62521 & ~n62528 ;
  assign n62530 = ~n10003 & ~n62529 ;
  assign n62531 = \pi0411  & n15247 ;
  assign n62532 = n62224 & ~n62531 ;
  assign n62533 = \pi0387  & ~\pi0591  ;
  assign n62534 = \pi0592  & ~n62533 ;
  assign n62535 = ~n62532 & ~n62534 ;
  assign n62536 = \pi0199  & ~\pi1053  ;
  assign n62537 = ~\pi0199  & ~\pi0295  ;
  assign n62538 = ~n62178 & ~n62537 ;
  assign n62539 = ~n62536 & n62538 ;
  assign n62540 = \pi0452  & ~\pi0592  ;
  assign n62541 = n62182 & n62540 ;
  assign n62542 = ~n62539 & ~n62541 ;
  assign n62543 = ~n62535 & n62542 ;
  assign n62544 = n10003 & n62539 ;
  assign n62545 = \pi0435  & ~\pi0592  ;
  assign n62546 = n9927 & n62545 ;
  assign n62547 = \pi0588  & ~n62546 ;
  assign n62548 = n62192 & ~n62547 ;
  assign n62549 = ~n62544 & ~n62548 ;
  assign n62550 = ~n62543 & ~n62549 ;
  assign n62551 = ~n62530 & ~n62550 ;
  assign n62552 = \pi0336  & n62171 ;
  assign n62553 = \pi0463  & \pi0591  ;
  assign n62554 = ~\pi0592  & n62553 ;
  assign n62555 = ~n62552 & ~n62554 ;
  assign n62556 = ~\pi0590  & ~n62555 ;
  assign n62557 = \pi0199  & ~\pi1070  ;
  assign n62558 = ~\pi0199  & ~\pi0256  ;
  assign n62559 = ~n62178 & ~n62558 ;
  assign n62560 = ~n62557 & n62559 ;
  assign n62561 = \pi0362  & ~\pi0592  ;
  assign n62562 = n62182 & n62561 ;
  assign n62563 = ~\pi0588  & ~n62562 ;
  assign n62564 = ~n62560 & n62563 ;
  assign n62565 = ~n62556 & n62564 ;
  assign n62566 = n10003 & n62560 ;
  assign n62567 = \pi0437  & ~\pi0592  ;
  assign n62568 = n9927 & n62567 ;
  assign n62569 = \pi0588  & ~n62568 ;
  assign n62570 = n62192 & ~n62569 ;
  assign n62571 = ~n62566 & ~n62570 ;
  assign n62572 = ~n62565 & ~n62571 ;
  assign n62573 = \pi0783  & \pi1135  ;
  assign n62574 = \pi0804  & ~\pi1135  ;
  assign n62575 = ~n62573 & ~n62574 ;
  assign n62576 = ~\pi1136  & n62575 ;
  assign n62577 = \pi0639  & \pi1135  ;
  assign n62578 = \pi0622  & ~\pi1135  ;
  assign n62579 = \pi1136  & ~n62578 ;
  assign n62580 = ~n62577 & n62579 ;
  assign n62581 = ~n62576 & ~n62580 ;
  assign n62582 = ~\pi1134  & ~n62581 ;
  assign n62583 = ~\pi0735  & \pi1135  ;
  assign n62584 = ~\pi0743  & ~\pi1135  ;
  assign n62585 = ~n62583 & ~n62584 ;
  assign n62586 = \pi1136  & n62585 ;
  assign n62587 = \pi0859  & n62258 ;
  assign n62588 = \pi1134  & ~n62587 ;
  assign n62589 = ~n62586 & n62588 ;
  assign n62590 = n62262 & ~n62589 ;
  assign n62591 = ~n62582 & n62590 ;
  assign n62592 = ~n62572 & ~n62591 ;
  assign n62593 = \pi0876  & n62258 ;
  assign n62594 = ~\pi0730  & \pi1135  ;
  assign n62595 = ~\pi0748  & ~\pi1135  ;
  assign n62596 = ~n62594 & ~n62595 ;
  assign n62597 = \pi1136  & n62596 ;
  assign n62598 = ~n62593 & ~n62597 ;
  assign n62599 = n62209 & ~n62598 ;
  assign n62600 = ~\pi0710  & \pi1135  ;
  assign n62601 = \pi1136  & ~n62600 ;
  assign n62602 = ~\pi0803  & ~\pi1135  ;
  assign n62603 = \pi0789  & n62208 ;
  assign n62604 = ~n62602 & ~n62603 ;
  assign n62605 = ~n62601 & n62604 ;
  assign n62606 = ~\pi0623  & \pi1136  ;
  assign n62607 = ~n62211 & n62606 ;
  assign n62608 = n62197 & ~n62607 ;
  assign n62609 = ~n62605 & n62608 ;
  assign n62610 = ~n62599 & ~n62609 ;
  assign n62611 = ~n10003 & ~n62610 ;
  assign n62612 = \pi0412  & n15247 ;
  assign n62613 = n62224 & ~n62612 ;
  assign n62614 = \pi0388  & ~\pi0591  ;
  assign n62615 = \pi0592  & ~n62614 ;
  assign n62616 = ~n62613 & ~n62615 ;
  assign n62617 = \pi0199  & ~\pi1037  ;
  assign n62618 = ~\pi0199  & ~\pi0296  ;
  assign n62619 = ~n62178 & ~n62618 ;
  assign n62620 = ~n62617 & n62619 ;
  assign n62621 = \pi0455  & ~\pi0592  ;
  assign n62622 = n62182 & n62621 ;
  assign n62623 = ~n62620 & ~n62622 ;
  assign n62624 = ~n62616 & n62623 ;
  assign n62625 = n10003 & n62620 ;
  assign n62626 = \pi0436  & ~\pi0592  ;
  assign n62627 = n9927 & n62626 ;
  assign n62628 = \pi0588  & ~n62627 ;
  assign n62629 = n62192 & ~n62628 ;
  assign n62630 = ~n62625 & ~n62629 ;
  assign n62631 = ~n62624 & ~n62630 ;
  assign n62632 = ~n62611 & ~n62631 ;
  assign n62633 = ~\pi0643  & \pi1135  ;
  assign n62634 = ~\pi0606  & ~\pi1135  ;
  assign n62635 = ~n62633 & ~n62634 ;
  assign n62636 = \pi1136  & n62635 ;
  assign n62637 = \pi0812  & ~\pi1135  ;
  assign n62638 = ~\pi0787  & \pi1135  ;
  assign n62639 = ~n62637 & ~n62638 ;
  assign n62640 = ~\pi1136  & n62639 ;
  assign n62641 = ~n62636 & ~n62640 ;
  assign n62642 = n62197 & ~n62641 ;
  assign n62643 = ~\pi0746  & \pi1136  ;
  assign n62644 = ~n62211 & n62643 ;
  assign n62645 = ~\pi0729  & \pi1135  ;
  assign n62646 = ~\pi0881  & ~\pi1136  ;
  assign n62647 = ~n62645 & ~n62646 ;
  assign n62648 = ~n62644 & n62647 ;
  assign n62649 = n62210 & n62648 ;
  assign n62650 = ~n62642 & ~n62649 ;
  assign n62651 = ~n10003 & ~n62650 ;
  assign n62652 = \pi0410  & n15247 ;
  assign n62653 = n62224 & ~n62652 ;
  assign n62654 = \pi0386  & ~\pi0591  ;
  assign n62655 = \pi0592  & ~n62654 ;
  assign n62656 = ~n62653 & ~n62655 ;
  assign n62657 = \pi0199  & ~\pi1059  ;
  assign n62658 = ~\pi0199  & ~\pi0293  ;
  assign n62659 = ~n62178 & ~n62658 ;
  assign n62660 = ~n62657 & n62659 ;
  assign n62661 = \pi0361  & ~\pi0592  ;
  assign n62662 = n62182 & n62661 ;
  assign n62663 = ~n62660 & ~n62662 ;
  assign n62664 = ~n62656 & n62663 ;
  assign n62665 = n10003 & n62660 ;
  assign n62666 = \pi0434  & ~\pi0592  ;
  assign n62667 = n9927 & n62666 ;
  assign n62668 = \pi0588  & ~n62667 ;
  assign n62669 = n62192 & ~n62668 ;
  assign n62670 = ~n62665 & ~n62669 ;
  assign n62671 = ~n62664 & ~n62670 ;
  assign n62672 = ~n62651 & ~n62671 ;
  assign n62673 = \pi0366  & n62171 ;
  assign n62674 = \pi0335  & \pi0591  ;
  assign n62675 = ~\pi0592  & n62674 ;
  assign n62676 = ~n62673 & ~n62675 ;
  assign n62677 = ~\pi0590  & ~n62676 ;
  assign n62678 = \pi0199  & ~\pi1069  ;
  assign n62679 = ~\pi0199  & ~\pi0259  ;
  assign n62680 = ~n62178 & ~n62679 ;
  assign n62681 = ~n62678 & n62680 ;
  assign n62682 = \pi0344  & ~\pi0592  ;
  assign n62683 = n62182 & n62682 ;
  assign n62684 = ~\pi0588  & ~n62683 ;
  assign n62685 = ~n62681 & n62684 ;
  assign n62686 = ~n62677 & n62685 ;
  assign n62687 = n10003 & n62681 ;
  assign n62688 = \pi0416  & ~\pi0592  ;
  assign n62689 = n9927 & n62688 ;
  assign n62690 = \pi0588  & ~n62689 ;
  assign n62691 = n62192 & ~n62690 ;
  assign n62692 = ~n62687 & ~n62691 ;
  assign n62693 = ~n62686 & ~n62692 ;
  assign n62694 = \pi0635  & \pi1135  ;
  assign n62695 = ~\pi1134  & ~n62694 ;
  assign n62696 = ~\pi0620  & ~\pi1135  ;
  assign n62697 = \pi1136  & ~n62696 ;
  assign n62698 = n62695 & n62697 ;
  assign n62699 = n62262 & n62698 ;
  assign n62700 = \pi0704  & \pi1135  ;
  assign n62701 = ~\pi0870  & ~\pi1136  ;
  assign n62702 = ~n62700 & ~n62701 ;
  assign n62703 = n62210 & n62702 ;
  assign n62704 = \pi0742  & \pi1136  ;
  assign n62705 = ~n62211 & n62704 ;
  assign n62706 = ~n10003 & ~n62705 ;
  assign n62707 = n62703 & n62706 ;
  assign n62708 = ~n62699 & ~n62707 ;
  assign n62709 = ~n62693 & n62708 ;
  assign n62710 = \pi0368  & n62171 ;
  assign n62711 = \pi0393  & \pi0591  ;
  assign n62712 = ~\pi0592  & n62711 ;
  assign n62713 = ~n62710 & ~n62712 ;
  assign n62714 = ~\pi0590  & ~n62713 ;
  assign n62715 = \pi0199  & ~\pi1067  ;
  assign n62716 = ~\pi0199  & ~\pi0260  ;
  assign n62717 = ~n62178 & ~n62716 ;
  assign n62718 = ~n62715 & n62717 ;
  assign n62719 = \pi0346  & ~\pi0592  ;
  assign n62720 = n62182 & n62719 ;
  assign n62721 = ~\pi0588  & ~n62720 ;
  assign n62722 = ~n62718 & n62721 ;
  assign n62723 = ~n62714 & n62722 ;
  assign n62724 = n10003 & n62718 ;
  assign n62725 = \pi0418  & ~\pi0592  ;
  assign n62726 = n9927 & n62725 ;
  assign n62727 = \pi0588  & ~n62726 ;
  assign n62728 = n62192 & ~n62727 ;
  assign n62729 = ~n62724 & ~n62728 ;
  assign n62730 = ~n62723 & ~n62729 ;
  assign n62731 = \pi0632  & \pi1135  ;
  assign n62732 = ~\pi1134  & ~n62731 ;
  assign n62733 = ~\pi0613  & ~\pi1135  ;
  assign n62734 = \pi1136  & ~n62733 ;
  assign n62735 = n62732 & n62734 ;
  assign n62736 = n62262 & n62735 ;
  assign n62737 = \pi0688  & \pi1135  ;
  assign n62738 = ~\pi0856  & ~\pi1136  ;
  assign n62739 = ~n62737 & ~n62738 ;
  assign n62740 = n62210 & n62739 ;
  assign n62741 = \pi0760  & \pi1136  ;
  assign n62742 = ~n62211 & n62741 ;
  assign n62743 = ~n10003 & ~n62742 ;
  assign n62744 = n62740 & n62743 ;
  assign n62745 = ~n62736 & ~n62744 ;
  assign n62746 = ~n62730 & n62745 ;
  assign n62747 = \pi0389  & n62171 ;
  assign n62748 = \pi0413  & \pi0591  ;
  assign n62749 = ~\pi0592  & n62748 ;
  assign n62750 = ~n62747 & ~n62749 ;
  assign n62751 = ~\pi0590  & ~n62750 ;
  assign n62752 = \pi0199  & ~\pi1036  ;
  assign n62753 = ~\pi0199  & ~\pi0255  ;
  assign n62754 = ~n62178 & ~n62753 ;
  assign n62755 = ~n62752 & n62754 ;
  assign n62756 = \pi0450  & ~\pi0592  ;
  assign n62757 = n62182 & n62756 ;
  assign n62758 = ~\pi0588  & ~n62757 ;
  assign n62759 = ~n62755 & n62758 ;
  assign n62760 = ~n62751 & n62759 ;
  assign n62761 = n10003 & n62755 ;
  assign n62762 = \pi0438  & ~\pi0592  ;
  assign n62763 = n9927 & n62762 ;
  assign n62764 = \pi0588  & ~n62763 ;
  assign n62765 = n62192 & ~n62764 ;
  assign n62766 = ~n62761 & ~n62765 ;
  assign n62767 = ~n62760 & ~n62766 ;
  assign n62768 = ~\pi0665  & \pi1136  ;
  assign n62769 = ~\pi0791  & ~\pi1136  ;
  assign n62770 = \pi1135  & ~n62769 ;
  assign n62771 = ~n62768 & n62770 ;
  assign n62772 = ~\pi0621  & \pi1136  ;
  assign n62773 = ~\pi0810  & ~\pi1136  ;
  assign n62774 = ~\pi1135  & ~n62773 ;
  assign n62775 = ~n62772 & n62774 ;
  assign n62776 = ~n62771 & ~n62775 ;
  assign n62777 = n62197 & ~n62776 ;
  assign n62778 = ~\pi0739  & \pi1136  ;
  assign n62779 = ~n62211 & n62778 ;
  assign n62780 = ~\pi0874  & ~\pi1136  ;
  assign n62781 = ~\pi0690  & \pi1135  ;
  assign n62782 = ~n62780 & ~n62781 ;
  assign n62783 = ~n62779 & n62782 ;
  assign n62784 = n62210 & n62783 ;
  assign n62785 = ~n62777 & ~n62784 ;
  assign n62786 = ~n10003 & ~n62785 ;
  assign n62787 = ~n62767 & ~n62786 ;
  assign n62788 = ~\pi0680  & ~n61933 ;
  assign n62789 = ~\pi0953  & ~\pi1100  ;
  assign n62790 = n61931 & n62789 ;
  assign n62791 = n61930 & n62790 ;
  assign n62792 = ~\pi0962  & ~n62791 ;
  assign n62793 = ~n62788 & n62792 ;
  assign n62794 = ~\pi0681  & ~n61933 ;
  assign n62795 = ~\pi0953  & ~\pi1103  ;
  assign n62796 = n61931 & n62795 ;
  assign n62797 = n61930 & n62796 ;
  assign n62798 = ~\pi0962  & ~n62797 ;
  assign n62799 = ~n62794 & n62798 ;
  assign n62800 = \pi0367  & n62171 ;
  assign n62801 = \pi0392  & \pi0591  ;
  assign n62802 = ~\pi0592  & n62801 ;
  assign n62803 = ~n62800 & ~n62802 ;
  assign n62804 = ~\pi0590  & ~n62803 ;
  assign n62805 = \pi0199  & ~\pi1039  ;
  assign n62806 = ~\pi0199  & ~\pi0251  ;
  assign n62807 = ~n62178 & ~n62806 ;
  assign n62808 = ~n62805 & n62807 ;
  assign n62809 = \pi0345  & ~\pi0592  ;
  assign n62810 = n62182 & n62809 ;
  assign n62811 = ~\pi0588  & ~n62810 ;
  assign n62812 = ~n62808 & n62811 ;
  assign n62813 = ~n62804 & n62812 ;
  assign n62814 = n10003 & n62808 ;
  assign n62815 = \pi0417  & ~\pi0592  ;
  assign n62816 = n9927 & n62815 ;
  assign n62817 = \pi0588  & ~n62816 ;
  assign n62818 = n62192 & ~n62817 ;
  assign n62819 = ~n62814 & ~n62818 ;
  assign n62820 = ~n62813 & ~n62819 ;
  assign n62821 = \pi0631  & \pi1135  ;
  assign n62822 = ~\pi1134  & ~n62821 ;
  assign n62823 = ~\pi0610  & ~\pi1135  ;
  assign n62824 = \pi1136  & ~n62823 ;
  assign n62825 = n62822 & n62824 ;
  assign n62826 = n62262 & n62825 ;
  assign n62827 = \pi0686  & \pi1135  ;
  assign n62828 = ~\pi0848  & ~\pi1136  ;
  assign n62829 = ~n62827 & ~n62828 ;
  assign n62830 = n62210 & n62829 ;
  assign n62831 = \pi0757  & \pi1136  ;
  assign n62832 = ~n62211 & n62831 ;
  assign n62833 = ~n10003 & ~n62832 ;
  assign n62834 = n62830 & n62833 ;
  assign n62835 = ~n62826 & ~n62834 ;
  assign n62836 = ~n62820 & n62835 ;
  assign n62837 = \pi0953  & n61931 ;
  assign n62838 = n61930 & n62837 ;
  assign n62839 = \pi0684  & ~n62838 ;
  assign n62840 = \pi0953  & ~\pi1130  ;
  assign n62841 = n61931 & n62840 ;
  assign n62842 = n61930 & n62841 ;
  assign n62843 = ~\pi0962  & ~n62842 ;
  assign n62844 = ~n62839 & n62843 ;
  assign n62845 = \pi0406  & ~\pi0592  ;
  assign n62846 = ~\pi0588  & \pi0591  ;
  assign n62847 = n62845 & n62846 ;
  assign n62848 = ~\pi0590  & n62847 ;
  assign n62849 = \pi0590  & ~\pi0592  ;
  assign n62850 = \pi0357  & n62849 ;
  assign n62851 = \pi0382  & n62223 ;
  assign n62852 = ~n62850 & ~n62851 ;
  assign n62853 = n9763 & ~n62852 ;
  assign n62854 = ~n62848 & ~n62853 ;
  assign n62855 = \pi0199  & ~\pi1076  ;
  assign n62856 = ~n62178 & ~n62855 ;
  assign n62857 = ~n56362 & n62856 ;
  assign n62858 = \pi0588  & ~\pi0590  ;
  assign n62859 = \pi0430  & n15292 ;
  assign n62860 = n62858 & n62859 ;
  assign n62861 = ~n62857 & ~n62860 ;
  assign n62862 = n62854 & n62861 ;
  assign n62863 = ~n62178 & n62855 ;
  assign n62864 = ~n56359 & ~n62178 ;
  assign n62865 = n56361 & n62864 ;
  assign n62866 = ~n62863 & ~n62865 ;
  assign n62867 = n10003 & n62866 ;
  assign n62868 = ~n62862 & n62867 ;
  assign n62869 = \pi0860  & n62258 ;
  assign n62870 = \pi0728  & \pi1135  ;
  assign n62871 = \pi0744  & ~\pi1135  ;
  assign n62872 = ~n62870 & ~n62871 ;
  assign n62873 = \pi1136  & n62872 ;
  assign n62874 = ~n62869 & ~n62873 ;
  assign n62875 = n62209 & ~n62874 ;
  assign n62876 = \pi1136  & ~n62196 ;
  assign n62877 = ~\pi1134  & ~n62876 ;
  assign n62878 = \pi0657  & \pi1135  ;
  assign n62879 = ~\pi0652  & ~\pi1135  ;
  assign n62880 = ~n62878 & ~n62879 ;
  assign n62881 = \pi1136  & n62880 ;
  assign n62882 = \pi0813  & n62258 ;
  assign n62883 = n62196 & n62882 ;
  assign n62884 = ~n62881 & ~n62883 ;
  assign n62885 = n62877 & ~n62884 ;
  assign n62886 = ~n62875 & ~n62885 ;
  assign n62887 = ~n10003 & ~n62886 ;
  assign n62888 = ~n62868 & ~n62887 ;
  assign n62889 = \pi0686  & ~n62838 ;
  assign n62890 = \pi0953  & ~\pi1113  ;
  assign n62891 = n61931 & n62890 ;
  assign n62892 = n61930 & n62891 ;
  assign n62893 = ~\pi0962  & ~n62892 ;
  assign n62894 = ~n62889 & n62893 ;
  assign n62895 = ~\pi0687  & ~n62838 ;
  assign n62896 = \pi0953  & ~\pi1127  ;
  assign n62897 = n61931 & n62896 ;
  assign n62898 = n61930 & n62897 ;
  assign n62899 = ~\pi0962  & ~n62898 ;
  assign n62900 = ~n62895 & n62899 ;
  assign n62901 = \pi0688  & ~n62838 ;
  assign n62902 = \pi0953  & ~\pi1115  ;
  assign n62903 = n61931 & n62902 ;
  assign n62904 = n61930 & n62903 ;
  assign n62905 = ~\pi0962  & ~n62904 ;
  assign n62906 = ~n62901 & n62905 ;
  assign n62907 = \pi0401  & ~\pi0592  ;
  assign n62908 = n62846 & n62907 ;
  assign n62909 = ~\pi0590  & n62908 ;
  assign n62910 = \pi0351  & n62849 ;
  assign n62911 = \pi0376  & n62223 ;
  assign n62912 = ~n62910 & ~n62911 ;
  assign n62913 = n9763 & ~n62912 ;
  assign n62914 = ~n62909 & ~n62913 ;
  assign n62915 = ~\pi0199  & n56331 ;
  assign n62916 = \pi0199  & ~\pi1079  ;
  assign n62917 = ~n62178 & ~n62916 ;
  assign n62918 = ~n62915 & n62917 ;
  assign n62919 = \pi0426  & n62858 ;
  assign n62920 = n15292 & n62919 ;
  assign n62921 = ~n62918 & ~n62920 ;
  assign n62922 = n62914 & n62921 ;
  assign n62923 = ~n62178 & n62916 ;
  assign n62924 = ~\pi0199  & ~n62178 ;
  assign n62925 = n56331 & n62924 ;
  assign n62926 = ~n62923 & ~n62925 ;
  assign n62927 = n10003 & n62926 ;
  assign n62928 = ~n62922 & n62927 ;
  assign n62929 = \pi0798  & n62258 ;
  assign n62930 = \pi0655  & \pi1135  ;
  assign n62931 = ~\pi0658  & ~\pi1135  ;
  assign n62932 = ~n62930 & ~n62931 ;
  assign n62933 = \pi1136  & n62932 ;
  assign n62934 = ~n62929 & ~n62933 ;
  assign n62935 = n62197 & ~n62934 ;
  assign n62936 = \pi0752  & \pi1136  ;
  assign n62937 = ~n62211 & n62936 ;
  assign n62938 = ~\pi0703  & \pi1135  ;
  assign n62939 = ~\pi0843  & ~\pi1136  ;
  assign n62940 = ~n62938 & ~n62939 ;
  assign n62941 = ~n62937 & n62940 ;
  assign n62942 = n62210 & n62941 ;
  assign n62943 = ~n62935 & ~n62942 ;
  assign n62944 = ~n10003 & ~n62943 ;
  assign n62945 = ~n62928 & ~n62944 ;
  assign n62946 = ~\pi0690  & ~n62838 ;
  assign n62947 = \pi0953  & ~\pi1108  ;
  assign n62948 = n61931 & n62947 ;
  assign n62949 = n61930 & n62948 ;
  assign n62950 = ~\pi0962  & ~n62949 ;
  assign n62951 = ~n62946 & n62950 ;
  assign n62952 = ~\pi0691  & ~n62838 ;
  assign n62953 = \pi0953  & ~\pi1107  ;
  assign n62954 = n61931 & n62953 ;
  assign n62955 = n61930 & n62954 ;
  assign n62956 = ~\pi0962  & ~n62955 ;
  assign n62957 = ~n62952 & n62956 ;
  assign n62958 = \pi0402  & ~\pi0592  ;
  assign n62959 = n62846 & n62958 ;
  assign n62960 = ~\pi0590  & n62959 ;
  assign n62961 = \pi0352  & n62849 ;
  assign n62962 = \pi0317  & n62223 ;
  assign n62963 = ~n62961 & ~n62962 ;
  assign n62964 = n9763 & ~n62963 ;
  assign n62965 = ~n62960 & ~n62964 ;
  assign n62966 = ~\pi0199  & n56343 ;
  assign n62967 = \pi0199  & ~\pi1078  ;
  assign n62968 = ~n62178 & ~n62967 ;
  assign n62969 = ~n62966 & n62968 ;
  assign n62970 = \pi0427  & n62858 ;
  assign n62971 = n15292 & n62970 ;
  assign n62972 = ~n62969 & ~n62971 ;
  assign n62973 = n62965 & n62972 ;
  assign n62974 = ~n62178 & n62967 ;
  assign n62975 = n56343 & n62924 ;
  assign n62976 = ~n62974 & ~n62975 ;
  assign n62977 = n10003 & n62976 ;
  assign n62978 = ~n62973 & n62977 ;
  assign n62979 = \pi0649  & \pi1135  ;
  assign n62980 = ~\pi0656  & ~\pi1135  ;
  assign n62981 = ~n62979 & ~n62980 ;
  assign n62982 = \pi1136  & n62981 ;
  assign n62983 = \pi0801  & n62258 ;
  assign n62984 = ~\pi1134  & ~n62983 ;
  assign n62985 = ~n62982 & n62984 ;
  assign n62986 = \pi0770  & ~\pi1135  ;
  assign n62987 = ~\pi0726  & \pi1135  ;
  assign n62988 = ~n62986 & ~n62987 ;
  assign n62989 = \pi1136  & n62988 ;
  assign n62990 = \pi0844  & n62258 ;
  assign n62991 = \pi1134  & ~n62990 ;
  assign n62992 = ~n62989 & n62991 ;
  assign n62993 = ~n62985 & ~n62992 ;
  assign n62994 = n62262 & n62993 ;
  assign n62995 = ~n62978 & ~n62994 ;
  assign n62996 = \pi0693  & ~n61933 ;
  assign n62997 = ~\pi0953  & ~\pi1129  ;
  assign n62998 = n61931 & n62997 ;
  assign n62999 = n61930 & n62998 ;
  assign n63000 = ~\pi0962  & ~n62999 ;
  assign n63001 = ~n62996 & n63000 ;
  assign n63002 = \pi0694  & ~n62838 ;
  assign n63003 = \pi0953  & ~\pi1128  ;
  assign n63004 = n61931 & n63003 ;
  assign n63005 = n61930 & n63004 ;
  assign n63006 = ~\pi0962  & ~n63005 ;
  assign n63007 = ~n63002 & n63006 ;
  assign n63008 = \pi0695  & ~n61933 ;
  assign n63009 = ~\pi0953  & ~\pi1111  ;
  assign n63010 = n61931 & n63009 ;
  assign n63011 = n61930 & n63010 ;
  assign n63012 = ~\pi0962  & ~n63011 ;
  assign n63013 = ~n63008 & n63012 ;
  assign n63014 = ~\pi0696  & ~n62838 ;
  assign n63015 = \pi0953  & ~\pi1100  ;
  assign n63016 = n61931 & n63015 ;
  assign n63017 = n61930 & n63016 ;
  assign n63018 = ~\pi0962  & ~n63017 ;
  assign n63019 = ~n63014 & n63018 ;
  assign n63020 = \pi0697  & ~n62838 ;
  assign n63021 = \pi0953  & ~\pi1129  ;
  assign n63022 = n61931 & n63021 ;
  assign n63023 = n61930 & n63022 ;
  assign n63024 = ~\pi0962  & ~n63023 ;
  assign n63025 = ~n63020 & n63024 ;
  assign n63026 = \pi0698  & ~n62838 ;
  assign n63027 = \pi0953  & ~\pi1116  ;
  assign n63028 = n61931 & n63027 ;
  assign n63029 = n61930 & n63028 ;
  assign n63030 = ~\pi0962  & ~n63029 ;
  assign n63031 = ~n63026 & n63030 ;
  assign n63032 = ~\pi0699  & ~n62838 ;
  assign n63033 = \pi0953  & ~\pi1103  ;
  assign n63034 = n61931 & n63033 ;
  assign n63035 = n61930 & n63034 ;
  assign n63036 = ~\pi0962  & ~n63035 ;
  assign n63037 = ~n63032 & n63036 ;
  assign n63038 = ~\pi0700  & ~n62838 ;
  assign n63039 = \pi0953  & ~\pi1110  ;
  assign n63040 = n61931 & n63039 ;
  assign n63041 = n61930 & n63040 ;
  assign n63042 = ~\pi0962  & ~n63041 ;
  assign n63043 = ~n63038 & n63042 ;
  assign n63044 = \pi0701  & ~n62838 ;
  assign n63045 = \pi0953  & ~\pi1123  ;
  assign n63046 = n61931 & n63045 ;
  assign n63047 = n61930 & n63046 ;
  assign n63048 = ~\pi0962  & ~n63047 ;
  assign n63049 = ~n63044 & n63048 ;
  assign n63050 = \pi0702  & ~n62838 ;
  assign n63051 = \pi0953  & ~\pi1117  ;
  assign n63052 = n61931 & n63051 ;
  assign n63053 = n61930 & n63052 ;
  assign n63054 = ~\pi0962  & ~n63053 ;
  assign n63055 = ~n63050 & n63054 ;
  assign n63056 = ~\pi0703  & ~n62838 ;
  assign n63057 = \pi0953  & ~\pi1124  ;
  assign n63058 = n61931 & n63057 ;
  assign n63059 = n61930 & n63058 ;
  assign n63060 = ~\pi0962  & ~n63059 ;
  assign n63061 = ~n63056 & n63060 ;
  assign n63062 = \pi0704  & ~n62838 ;
  assign n63063 = \pi0953  & ~\pi1112  ;
  assign n63064 = n61931 & n63063 ;
  assign n63065 = n61930 & n63064 ;
  assign n63066 = ~\pi0962  & ~n63065 ;
  assign n63067 = ~n63062 & n63066 ;
  assign n63068 = ~\pi0705  & ~n62838 ;
  assign n63069 = \pi0953  & ~\pi1125  ;
  assign n63070 = n61931 & n63069 ;
  assign n63071 = n61930 & n63070 ;
  assign n63072 = ~\pi0962  & ~n63071 ;
  assign n63073 = ~n63068 & n63072 ;
  assign n63074 = ~\pi0706  & ~n62838 ;
  assign n63075 = \pi0953  & ~\pi1105  ;
  assign n63076 = n61931 & n63075 ;
  assign n63077 = n61930 & n63076 ;
  assign n63078 = ~\pi0962  & ~n63077 ;
  assign n63079 = ~n63074 & n63078 ;
  assign n63080 = \pi0347  & \pi0590  ;
  assign n63081 = n15292 & n63080 ;
  assign n63082 = ~\pi0588  & n62178 ;
  assign n63083 = n63081 & n63082 ;
  assign n63084 = \pi0370  & n62171 ;
  assign n63085 = \pi0395  & \pi0591  ;
  assign n63086 = ~\pi0592  & n63085 ;
  assign n63087 = ~n63084 & ~n63086 ;
  assign n63088 = ~\pi0588  & ~\pi0590  ;
  assign n63089 = n62178 & n63088 ;
  assign n63090 = ~n63087 & n63089 ;
  assign n63091 = ~n63083 & ~n63090 ;
  assign n63092 = \pi0420  & \pi0588  ;
  assign n63093 = n62178 & n63092 ;
  assign n63094 = n9928 & n63093 ;
  assign n63095 = n10003 & ~n63094 ;
  assign n63096 = ~\pi0200  & ~\pi0304  ;
  assign n63097 = \pi0200  & ~\pi1048  ;
  assign n63098 = ~n63096 & ~n63097 ;
  assign n63099 = ~\pi0199  & ~n63098 ;
  assign n63100 = \pi0199  & ~\pi1055  ;
  assign n63101 = ~n62178 & ~n63100 ;
  assign n63102 = ~n63099 & n63101 ;
  assign n63103 = n63095 & ~n63102 ;
  assign n63104 = n63091 & n63103 ;
  assign n63105 = \pi0753  & \pi1136  ;
  assign n63106 = ~n62211 & n63105 ;
  assign n63107 = \pi0702  & \pi1135  ;
  assign n63108 = ~\pi0847  & ~\pi1136  ;
  assign n63109 = ~n63107 & ~n63108 ;
  assign n63110 = ~n63106 & n63109 ;
  assign n63111 = n62210 & n63110 ;
  assign n63112 = \pi1136  & n62196 ;
  assign n63113 = ~\pi0618  & ~\pi1135  ;
  assign n63114 = ~\pi0627  & \pi1135  ;
  assign n63115 = ~\pi1134  & ~n63114 ;
  assign n63116 = ~n63113 & n63115 ;
  assign n63117 = n63112 & n63116 ;
  assign n63118 = ~n10003 & ~n63117 ;
  assign n63119 = ~n63111 & n63118 ;
  assign n63120 = ~n63104 & ~n63119 ;
  assign n63121 = ~\pi0592  & n62182 ;
  assign n63122 = \pi0321  & ~\pi0588  ;
  assign n63123 = n62178 & n63122 ;
  assign n63124 = n63121 & n63123 ;
  assign n63125 = n62171 & n62178 ;
  assign n63126 = \pi0442  & n63125 ;
  assign n63127 = ~\pi0592  & n62178 ;
  assign n63128 = \pi0328  & \pi0591  ;
  assign n63129 = n63127 & n63128 ;
  assign n63130 = ~n63126 & ~n63129 ;
  assign n63131 = n9782 & ~n63130 ;
  assign n63132 = ~n63124 & ~n63131 ;
  assign n63133 = ~\pi0200  & ~\pi0305  ;
  assign n63134 = \pi0200  & ~\pi1084  ;
  assign n63135 = ~n63133 & ~n63134 ;
  assign n63136 = ~\pi0199  & ~n63135 ;
  assign n63137 = \pi0199  & ~\pi1058  ;
  assign n63138 = ~n62178 & ~n63137 ;
  assign n63139 = ~n63136 & n63138 ;
  assign n63140 = n15292 & n62178 ;
  assign n63141 = \pi0459  & n62858 ;
  assign n63142 = n63140 & n63141 ;
  assign n63143 = n10003 & ~n63142 ;
  assign n63144 = ~n63139 & n63143 ;
  assign n63145 = n63132 & n63144 ;
  assign n63146 = \pi0754  & \pi1136  ;
  assign n63147 = ~n62211 & n63146 ;
  assign n63148 = ~\pi0857  & ~\pi1136  ;
  assign n63149 = \pi0709  & \pi1135  ;
  assign n63150 = ~n63148 & ~n63149 ;
  assign n63151 = ~n63147 & n63150 ;
  assign n63152 = n62210 & n63151 ;
  assign n63153 = ~\pi0609  & ~\pi1135  ;
  assign n63154 = ~\pi0660  & \pi1135  ;
  assign n63155 = ~\pi1134  & ~n63154 ;
  assign n63156 = ~n63153 & n63155 ;
  assign n63157 = n63112 & n63156 ;
  assign n63158 = ~n10003 & ~n63157 ;
  assign n63159 = ~n63152 & n63158 ;
  assign n63160 = ~n63145 & ~n63159 ;
  assign n63161 = \pi0709  & ~n62838 ;
  assign n63162 = \pi0953  & ~\pi1118  ;
  assign n63163 = n61931 & n63162 ;
  assign n63164 = n61930 & n63163 ;
  assign n63165 = ~\pi0962  & ~n63164 ;
  assign n63166 = ~n63161 & n63165 ;
  assign n63167 = ~\pi0710  & ~n61933 ;
  assign n63168 = ~\pi0953  & ~\pi1106  ;
  assign n63169 = n61931 & n63168 ;
  assign n63170 = n61930 & n63169 ;
  assign n63171 = ~\pi0962  & ~n63170 ;
  assign n63172 = ~n63167 & n63171 ;
  assign n63173 = \pi0348  & ~\pi0588  ;
  assign n63174 = n62178 & n63173 ;
  assign n63175 = n63121 & n63174 ;
  assign n63176 = \pi0373  & n62171 ;
  assign n63177 = \pi0398  & \pi0591  ;
  assign n63178 = ~\pi0592  & n63177 ;
  assign n63179 = ~n63176 & ~n63178 ;
  assign n63180 = n63089 & ~n63179 ;
  assign n63181 = ~n63175 & ~n63180 ;
  assign n63182 = \pi0423  & \pi0588  ;
  assign n63183 = n62178 & n63182 ;
  assign n63184 = n9928 & n63183 ;
  assign n63185 = n10003 & ~n63184 ;
  assign n63186 = ~\pi0200  & ~\pi0306  ;
  assign n63187 = \pi0200  & ~\pi1059  ;
  assign n63188 = ~n63186 & ~n63187 ;
  assign n63189 = ~\pi0199  & ~n63188 ;
  assign n63190 = \pi0199  & ~\pi1087  ;
  assign n63191 = ~n62178 & ~n63190 ;
  assign n63192 = ~n63189 & n63191 ;
  assign n63193 = n63185 & ~n63192 ;
  assign n63194 = n63181 & n63193 ;
  assign n63195 = \pi0755  & \pi1136  ;
  assign n63196 = ~n62211 & n63195 ;
  assign n63197 = \pi0725  & \pi1135  ;
  assign n63198 = ~\pi0858  & ~\pi1136  ;
  assign n63199 = ~n63197 & ~n63198 ;
  assign n63200 = ~n63196 & n63199 ;
  assign n63201 = n62210 & n63200 ;
  assign n63202 = ~\pi0630  & ~\pi1135  ;
  assign n63203 = ~\pi0647  & \pi1135  ;
  assign n63204 = ~\pi1134  & ~n63203 ;
  assign n63205 = ~n63202 & n63204 ;
  assign n63206 = n63112 & n63205 ;
  assign n63207 = ~n10003 & ~n63206 ;
  assign n63208 = ~n63201 & n63207 ;
  assign n63209 = ~n63194 & ~n63208 ;
  assign n63210 = ~\pi0715  & \pi1135  ;
  assign n63211 = ~\pi1134  & ~n63210 ;
  assign n63212 = ~\pi0644  & ~\pi1135  ;
  assign n63213 = \pi1136  & ~n63212 ;
  assign n63214 = n63211 & n63213 ;
  assign n63215 = n62262 & n63214 ;
  assign n63216 = ~\pi0842  & ~\pi1136  ;
  assign n63217 = \pi0701  & \pi1135  ;
  assign n63218 = ~n63216 & ~n63217 ;
  assign n63219 = n62210 & n63218 ;
  assign n63220 = \pi0751  & \pi1136  ;
  assign n63221 = ~n62211 & n63220 ;
  assign n63222 = ~n10003 & ~n63221 ;
  assign n63223 = n63219 & n63222 ;
  assign n63224 = ~n63215 & ~n63223 ;
  assign n63225 = \pi0374  & n62171 ;
  assign n63226 = \pi0400  & \pi0591  ;
  assign n63227 = ~\pi0592  & n63226 ;
  assign n63228 = ~n63225 & ~n63227 ;
  assign n63229 = n9782 & ~n63228 ;
  assign n63230 = \pi0350  & ~\pi0592  ;
  assign n63231 = n62182 & n63230 ;
  assign n63232 = ~\pi0588  & n63231 ;
  assign n63233 = \pi0425  & n62858 ;
  assign n63234 = n15292 & n63233 ;
  assign n63235 = ~n63232 & ~n63234 ;
  assign n63236 = ~n63229 & n63235 ;
  assign n63237 = n62178 & n63236 ;
  assign n63238 = \pi1044  & n13645 ;
  assign n63239 = \pi0298  & n12691 ;
  assign n63240 = \pi0199  & \pi1035  ;
  assign n63241 = ~n62178 & ~n63240 ;
  assign n63242 = ~n63239 & n63241 ;
  assign n63243 = ~n63238 & n63242 ;
  assign n63244 = n10003 & ~n63243 ;
  assign n63245 = ~n63237 & n63244 ;
  assign n63246 = n63224 & ~n63245 ;
  assign n63247 = \pi0322  & ~\pi0588  ;
  assign n63248 = n62178 & n63247 ;
  assign n63249 = n63121 & n63248 ;
  assign n63250 = \pi0371  & n62171 ;
  assign n63251 = \pi0396  & \pi0591  ;
  assign n63252 = ~\pi0592  & n63251 ;
  assign n63253 = ~n63250 & ~n63252 ;
  assign n63254 = n63089 & ~n63253 ;
  assign n63255 = ~n63249 & ~n63254 ;
  assign n63256 = \pi0421  & \pi0588  ;
  assign n63257 = n62178 & n63256 ;
  assign n63258 = n9928 & n63257 ;
  assign n63259 = n10003 & ~n63258 ;
  assign n63260 = ~\pi0200  & ~\pi0309  ;
  assign n63261 = \pi0200  & ~\pi1072  ;
  assign n63262 = ~n63260 & ~n63261 ;
  assign n63263 = ~\pi0199  & ~n63262 ;
  assign n63264 = \pi0199  & ~\pi1051  ;
  assign n63265 = ~n62178 & ~n63264 ;
  assign n63266 = ~n63263 & n63265 ;
  assign n63267 = n63259 & ~n63266 ;
  assign n63268 = n63255 & n63267 ;
  assign n63269 = \pi0756  & \pi1136  ;
  assign n63270 = ~n62211 & n63269 ;
  assign n63271 = \pi0734  & \pi1135  ;
  assign n63272 = ~\pi0854  & ~\pi1136  ;
  assign n63273 = ~n63271 & ~n63272 ;
  assign n63274 = ~n63270 & n63273 ;
  assign n63275 = n62210 & n63274 ;
  assign n63276 = ~\pi0629  & ~\pi1135  ;
  assign n63277 = ~\pi0628  & \pi1135  ;
  assign n63278 = ~\pi1134  & ~n63277 ;
  assign n63279 = ~n63276 & n63278 ;
  assign n63280 = n63112 & n63279 ;
  assign n63281 = ~n10003 & ~n63280 ;
  assign n63282 = ~n63275 & n63281 ;
  assign n63283 = ~n63268 & ~n63282 ;
  assign n63284 = \pi0326  & ~\pi0592  ;
  assign n63285 = n62846 & n63284 ;
  assign n63286 = ~\pi0590  & n63285 ;
  assign n63287 = \pi0461  & n62849 ;
  assign n63288 = \pi0439  & n62223 ;
  assign n63289 = ~n63287 & ~n63288 ;
  assign n63290 = n9763 & ~n63289 ;
  assign n63291 = ~n63286 & ~n63290 ;
  assign n63292 = \pi0199  & ~\pi1057  ;
  assign n63293 = ~n62178 & ~n63292 ;
  assign n63294 = ~n55614 & n63293 ;
  assign n63295 = \pi0449  & n62858 ;
  assign n63296 = n15292 & n63295 ;
  assign n63297 = ~n63294 & ~n63296 ;
  assign n63298 = n63291 & n63297 ;
  assign n63299 = ~n62178 & n63292 ;
  assign n63300 = ~n55611 & ~n62178 ;
  assign n63301 = n55613 & n63300 ;
  assign n63302 = ~n63299 & ~n63301 ;
  assign n63303 = n10003 & n63302 ;
  assign n63304 = ~n63298 & n63303 ;
  assign n63305 = \pi0867  & n62258 ;
  assign n63306 = \pi0697  & \pi1135  ;
  assign n63307 = \pi0762  & ~\pi1135  ;
  assign n63308 = ~n63306 & ~n63307 ;
  assign n63309 = \pi1136  & n63308 ;
  assign n63310 = ~n63305 & ~n63309 ;
  assign n63311 = n62209 & ~n63310 ;
  assign n63312 = \pi0693  & \pi1135  ;
  assign n63313 = ~\pi0653  & ~\pi1135  ;
  assign n63314 = ~n63312 & ~n63313 ;
  assign n63315 = \pi1136  & n63314 ;
  assign n63316 = \pi0816  & n62258 ;
  assign n63317 = n62196 & n63316 ;
  assign n63318 = ~n63315 & ~n63317 ;
  assign n63319 = n62877 & ~n63318 ;
  assign n63320 = ~n63311 & ~n63319 ;
  assign n63321 = ~n10003 & ~n63320 ;
  assign n63322 = ~n63304 & ~n63321 ;
  assign n63323 = ~\pi0715  & ~n61933 ;
  assign n63324 = ~\pi0953  & ~\pi1123  ;
  assign n63325 = n61931 & n63324 ;
  assign n63326 = n61930 & n63325 ;
  assign n63327 = ~\pi0962  & ~n63326 ;
  assign n63328 = ~n63323 & n63327 ;
  assign n63329 = \pi0454  & n62858 ;
  assign n63330 = n63140 & n63329 ;
  assign n63331 = n10003 & ~n63330 ;
  assign n63332 = \pi0440  & n63125 ;
  assign n63333 = \pi0329  & ~\pi0592  ;
  assign n63334 = n62178 & n63333 ;
  assign n63335 = \pi0591  & n63334 ;
  assign n63336 = ~n63332 & ~n63335 ;
  assign n63337 = n9782 & ~n63336 ;
  assign n63338 = \pi0349  & ~\pi0592  ;
  assign n63339 = n62182 & n63338 ;
  assign n63340 = n63082 & n63339 ;
  assign n63341 = ~\pi0200  & ~\pi0307  ;
  assign n63342 = \pi0200  & ~\pi1053  ;
  assign n63343 = ~n63341 & ~n63342 ;
  assign n63344 = ~\pi0199  & ~n63343 ;
  assign n63345 = \pi0199  & ~\pi1043  ;
  assign n63346 = ~n62178 & ~n63345 ;
  assign n63347 = ~n63344 & n63346 ;
  assign n63348 = ~n63340 & ~n63347 ;
  assign n63349 = ~n63337 & n63348 ;
  assign n63350 = n63331 & n63349 ;
  assign n63351 = \pi0761  & \pi1136  ;
  assign n63352 = ~n62211 & n63351 ;
  assign n63353 = ~\pi0845  & ~\pi1136  ;
  assign n63354 = \pi0738  & \pi1135  ;
  assign n63355 = ~n63353 & ~n63354 ;
  assign n63356 = ~n63352 & n63355 ;
  assign n63357 = n62210 & n63356 ;
  assign n63358 = ~\pi0626  & ~\pi1135  ;
  assign n63359 = ~\pi0641  & \pi1135  ;
  assign n63360 = ~\pi1134  & ~n63359 ;
  assign n63361 = ~n63358 & n63360 ;
  assign n63362 = n63112 & n63361 ;
  assign n63363 = ~n10003 & ~n63362 ;
  assign n63364 = ~n63357 & n63363 ;
  assign n63365 = ~n63350 & ~n63364 ;
  assign n63366 = \pi0462  & ~\pi0588  ;
  assign n63367 = n62178 & n63366 ;
  assign n63368 = n63121 & n63367 ;
  assign n63369 = \pi0377  & n62171 ;
  assign n63370 = \pi0318  & \pi0591  ;
  assign n63371 = ~\pi0592  & n63370 ;
  assign n63372 = ~n63369 & ~n63371 ;
  assign n63373 = n63089 & ~n63372 ;
  assign n63374 = ~n63368 & ~n63373 ;
  assign n63375 = \pi0448  & \pi0588  ;
  assign n63376 = n62178 & n63375 ;
  assign n63377 = n9928 & n63376 ;
  assign n63378 = ~\pi0199  & n56337 ;
  assign n63379 = \pi0199  & ~\pi1074  ;
  assign n63380 = ~n62178 & ~n63379 ;
  assign n63381 = ~n63378 & n63380 ;
  assign n63382 = ~n63377 & ~n63381 ;
  assign n63383 = n63374 & n63382 ;
  assign n63384 = n10003 & ~n63383 ;
  assign n63385 = \pi0800  & n62258 ;
  assign n63386 = \pi0669  & \pi1135  ;
  assign n63387 = ~\pi0645  & ~\pi1135  ;
  assign n63388 = ~n63386 & ~n63387 ;
  assign n63389 = \pi1136  & n63388 ;
  assign n63390 = ~n63385 & ~n63389 ;
  assign n63391 = n62197 & ~n63390 ;
  assign n63392 = \pi0768  & \pi1136  ;
  assign n63393 = ~n62211 & n63392 ;
  assign n63394 = ~\pi0839  & ~\pi1136  ;
  assign n63395 = ~\pi0705  & \pi1135  ;
  assign n63396 = ~n63394 & ~n63395 ;
  assign n63397 = ~n63393 & n63396 ;
  assign n63398 = n62210 & n63397 ;
  assign n63399 = ~n63391 & ~n63398 ;
  assign n63400 = ~n10003 & ~n63399 ;
  assign n63401 = ~n63384 & ~n63400 ;
  assign n63402 = \pi0419  & n62858 ;
  assign n63403 = n63140 & n63402 ;
  assign n63404 = n10003 & ~n63403 ;
  assign n63405 = \pi0369  & n63125 ;
  assign n63406 = \pi0394  & ~\pi0592  ;
  assign n63407 = n62178 & n63406 ;
  assign n63408 = \pi0591  & n63407 ;
  assign n63409 = ~n63405 & ~n63408 ;
  assign n63410 = n9782 & ~n63409 ;
  assign n63411 = \pi0315  & ~\pi0592  ;
  assign n63412 = n62182 & n63411 ;
  assign n63413 = n63082 & n63412 ;
  assign n63414 = ~\pi0200  & ~\pi0303  ;
  assign n63415 = \pi0200  & ~\pi1049  ;
  assign n63416 = ~n63414 & ~n63415 ;
  assign n63417 = ~\pi0199  & ~n63416 ;
  assign n63418 = \pi0199  & ~\pi1080  ;
  assign n63419 = ~n62178 & ~n63418 ;
  assign n63420 = ~n63417 & n63419 ;
  assign n63421 = ~n63413 & ~n63420 ;
  assign n63422 = ~n63410 & n63421 ;
  assign n63423 = n63404 & n63422 ;
  assign n63424 = \pi0767  & \pi1136  ;
  assign n63425 = ~n62211 & n63424 ;
  assign n63426 = ~\pi0853  & ~\pi1136  ;
  assign n63427 = \pi0698  & \pi1135  ;
  assign n63428 = ~n63426 & ~n63427 ;
  assign n63429 = ~n63425 & n63428 ;
  assign n63430 = n62210 & n63429 ;
  assign n63431 = ~\pi0608  & ~\pi1135  ;
  assign n63432 = ~\pi0625  & \pi1135  ;
  assign n63433 = ~\pi1134  & ~n63432 ;
  assign n63434 = ~n63431 & n63433 ;
  assign n63435 = n63112 & n63434 ;
  assign n63436 = ~n10003 & ~n63435 ;
  assign n63437 = ~n63430 & n63436 ;
  assign n63438 = ~n63423 & ~n63437 ;
  assign n63439 = \pi0353  & ~\pi0588  ;
  assign n63440 = n62178 & n63439 ;
  assign n63441 = n63121 & n63440 ;
  assign n63442 = \pi0378  & n62171 ;
  assign n63443 = \pi0325  & \pi0591  ;
  assign n63444 = ~\pi0592  & n63443 ;
  assign n63445 = ~n63442 & ~n63444 ;
  assign n63446 = n63089 & ~n63445 ;
  assign n63447 = ~n63441 & ~n63446 ;
  assign n63448 = \pi0451  & \pi0588  ;
  assign n63449 = n62178 & n63448 ;
  assign n63450 = n9928 & n63449 ;
  assign n63451 = ~\pi0199  & n56349 ;
  assign n63452 = \pi0199  & ~\pi1063  ;
  assign n63453 = ~n62178 & ~n63452 ;
  assign n63454 = ~n63451 & n63453 ;
  assign n63455 = ~n63450 & ~n63454 ;
  assign n63456 = n63447 & n63455 ;
  assign n63457 = n10003 & ~n63456 ;
  assign n63458 = \pi0807  & n62258 ;
  assign n63459 = \pi0650  & \pi1135  ;
  assign n63460 = ~\pi0636  & ~\pi1135  ;
  assign n63461 = ~n63459 & ~n63460 ;
  assign n63462 = \pi1136  & n63461 ;
  assign n63463 = ~n63458 & ~n63462 ;
  assign n63464 = n62197 & ~n63463 ;
  assign n63465 = \pi0774  & \pi1136  ;
  assign n63466 = ~n62211 & n63465 ;
  assign n63467 = ~\pi0868  & ~\pi1136  ;
  assign n63468 = ~\pi0687  & \pi1135  ;
  assign n63469 = ~n63467 & ~n63468 ;
  assign n63470 = ~n63466 & n63469 ;
  assign n63471 = n62210 & n63470 ;
  assign n63472 = ~n63464 & ~n63471 ;
  assign n63473 = ~n10003 & ~n63472 ;
  assign n63474 = ~n63457 & ~n63473 ;
  assign n63475 = \pi0405  & ~\pi0592  ;
  assign n63476 = n62846 & n63475 ;
  assign n63477 = ~\pi0590  & n63476 ;
  assign n63478 = \pi0356  & n62849 ;
  assign n63479 = \pi0381  & n62223 ;
  assign n63480 = ~n63478 & ~n63479 ;
  assign n63481 = n9763 & ~n63480 ;
  assign n63482 = ~n63477 & ~n63481 ;
  assign n63483 = \pi0199  & ~\pi1081  ;
  assign n63484 = ~n62178 & ~n63483 ;
  assign n63485 = ~n56369 & n63484 ;
  assign n63486 = \pi0445  & n62858 ;
  assign n63487 = n15292 & n63486 ;
  assign n63488 = ~n63485 & ~n63487 ;
  assign n63489 = n63482 & n63488 ;
  assign n63490 = ~n62178 & n63483 ;
  assign n63491 = ~n56366 & ~n62178 ;
  assign n63492 = n56368 & n63491 ;
  assign n63493 = ~n63490 & ~n63492 ;
  assign n63494 = n10003 & n63493 ;
  assign n63495 = ~n63489 & n63494 ;
  assign n63496 = \pi0880  & n62258 ;
  assign n63497 = \pi0684  & \pi1135  ;
  assign n63498 = \pi0750  & ~\pi1135  ;
  assign n63499 = ~n63497 & ~n63498 ;
  assign n63500 = \pi1136  & n63499 ;
  assign n63501 = ~n63496 & ~n63500 ;
  assign n63502 = n62209 & ~n63501 ;
  assign n63503 = \pi0654  & \pi1135  ;
  assign n63504 = ~\pi0651  & ~\pi1135  ;
  assign n63505 = ~n63503 & ~n63504 ;
  assign n63506 = \pi1136  & n63505 ;
  assign n63507 = \pi0794  & n62258 ;
  assign n63508 = n62196 & n63507 ;
  assign n63509 = ~n63506 & ~n63508 ;
  assign n63510 = n62877 & ~n63509 ;
  assign n63511 = ~n63502 & ~n63510 ;
  assign n63512 = ~n10003 & ~n63511 ;
  assign n63513 = ~n63495 & ~n63512 ;
  assign n63514 = ~\pi0731  & ~\pi0795  ;
  assign n63515 = \pi0731  & \pi0795  ;
  assign n63516 = ~n63514 & ~n63515 ;
  assign n63517 = ~\pi0945  & \pi0988  ;
  assign n63518 = \pi0731  & n63517 ;
  assign n63519 = \pi0721  & ~n63518 ;
  assign n63520 = n63516 & n63519 ;
  assign n63521 = ~\pi0765  & ~\pi0798  ;
  assign n63522 = \pi0765  & \pi0798  ;
  assign n63523 = ~n63521 & ~n63522 ;
  assign n63524 = ~\pi0747  & \pi0807  ;
  assign n63525 = \pi0747  & ~\pi0807  ;
  assign n63526 = ~n63524 & ~n63525 ;
  assign n63527 = ~n63523 & n63526 ;
  assign n63528 = ~\pi0771  & ~\pi0800  ;
  assign n63529 = \pi0771  & \pi0800  ;
  assign n63530 = ~n63528 & ~n63529 ;
  assign n63531 = ~\pi0769  & ~\pi0794  ;
  assign n63532 = \pi0769  & \pi0794  ;
  assign n63533 = ~n63531 & ~n63532 ;
  assign n63534 = ~n63530 & ~n63533 ;
  assign n63535 = n63527 & n63534 ;
  assign n63536 = \pi0721  & \pi0813  ;
  assign n63537 = ~\pi0773  & ~\pi0801  ;
  assign n63538 = \pi0773  & \pi0801  ;
  assign n63539 = ~n63537 & ~n63538 ;
  assign n63540 = n63536 & ~n63539 ;
  assign n63541 = ~\pi0775  & ~\pi0816  ;
  assign n63542 = \pi0775  & \pi0816  ;
  assign n63543 = ~n63541 & ~n63542 ;
  assign n63544 = n63540 & ~n63543 ;
  assign n63545 = n63535 & n63544 ;
  assign n63546 = \pi0731  & \pi0775  ;
  assign n63547 = n63517 & n63546 ;
  assign n63548 = \pi0721  & ~n63547 ;
  assign n63549 = ~n63545 & n63548 ;
  assign n63550 = ~n63520 & ~n63549 ;
  assign n63551 = n63535 & n63540 ;
  assign n63552 = \pi0807  & ~n63523 ;
  assign n63553 = ~\pi0721  & ~\pi0813  ;
  assign n63554 = \pi0794  & \pi0801  ;
  assign n63555 = n63553 & n63554 ;
  assign n63556 = ~n63530 & n63555 ;
  assign n63557 = n63552 & n63556 ;
  assign n63558 = \pi0775  & ~n63557 ;
  assign n63559 = ~n63551 & n63558 ;
  assign n63560 = \pi0775  & ~\pi0816  ;
  assign n63561 = \pi0795  & ~n63560 ;
  assign n63562 = ~n63559 & n63561 ;
  assign n63563 = \pi0747  & \pi0773  ;
  assign n63564 = \pi0769  & \pi0775  ;
  assign n63565 = n63563 & n63564 ;
  assign n63566 = \pi0721  & \pi0731  ;
  assign n63567 = n63517 & n63566 ;
  assign n63568 = ~n63565 & n63567 ;
  assign n63569 = ~\pi0721  & \pi0731  ;
  assign n63570 = n63517 & n63569 ;
  assign n63571 = n63565 & n63570 ;
  assign n63572 = ~n63568 & ~n63571 ;
  assign n63573 = ~n63562 & ~n63572 ;
  assign n63574 = n63550 & ~n63573 ;
  assign n63575 = \pi0732  & ~\pi1134  ;
  assign n63576 = \pi0694  & \pi1134  ;
  assign n63577 = \pi1135  & \pi1136  ;
  assign n63578 = ~n63576 & n63577 ;
  assign n63579 = ~n63575 & n63578 ;
  assign n63580 = \pi0776  & \pi1134  ;
  assign n63581 = ~\pi0640  & ~\pi1134  ;
  assign n63582 = ~n63580 & ~n63581 ;
  assign n63583 = ~\pi1135  & \pi1136  ;
  assign n63584 = n63582 & n63583 ;
  assign n63585 = ~\pi0851  & \pi1134  ;
  assign n63586 = ~\pi0795  & ~\pi1134  ;
  assign n63587 = ~n63585 & ~n63586 ;
  assign n63588 = n62258 & n63587 ;
  assign n63589 = ~n63584 & ~n63588 ;
  assign n63590 = ~n63579 & n63589 ;
  assign n63591 = n62262 & ~n63590 ;
  assign n63592 = \pi0354  & ~\pi0588  ;
  assign n63593 = n62178 & n63592 ;
  assign n63594 = n63121 & n63593 ;
  assign n63595 = \pi0379  & n62171 ;
  assign n63596 = \pi0403  & \pi0591  ;
  assign n63597 = ~\pi0592  & n63596 ;
  assign n63598 = ~n63595 & ~n63597 ;
  assign n63599 = n63089 & ~n63598 ;
  assign n63600 = ~n63594 & ~n63599 ;
  assign n63601 = \pi0428  & \pi0588  ;
  assign n63602 = n62178 & n63601 ;
  assign n63603 = n9928 & n63602 ;
  assign n63604 = ~\pi0199  & n56355 ;
  assign n63605 = \pi0199  & ~\pi1045  ;
  assign n63606 = ~n62178 & ~n63605 ;
  assign n63607 = ~n63604 & n63606 ;
  assign n63608 = ~n63603 & ~n63607 ;
  assign n63609 = n63600 & n63608 ;
  assign n63610 = ~\pi1163  & n9996 ;
  assign n63611 = ~n63609 & n63610 ;
  assign n63612 = ~n63591 & ~n63611 ;
  assign n63613 = \pi0723  & ~n62838 ;
  assign n63614 = \pi0953  & ~\pi1111  ;
  assign n63615 = n61931 & n63614 ;
  assign n63616 = n61930 & n63615 ;
  assign n63617 = ~\pi0962  & ~n63616 ;
  assign n63618 = ~n63613 & n63617 ;
  assign n63619 = \pi0724  & ~n62838 ;
  assign n63620 = \pi0953  & ~\pi1114  ;
  assign n63621 = n61931 & n63620 ;
  assign n63622 = n61930 & n63621 ;
  assign n63623 = ~\pi0962  & ~n63622 ;
  assign n63624 = ~n63619 & n63623 ;
  assign n63625 = \pi0725  & ~n62838 ;
  assign n63626 = \pi0953  & ~\pi1120  ;
  assign n63627 = n61931 & n63626 ;
  assign n63628 = n61930 & n63627 ;
  assign n63629 = ~\pi0962  & ~n63628 ;
  assign n63630 = ~n63625 & n63629 ;
  assign n63631 = ~\pi0726  & ~n62838 ;
  assign n63632 = \pi0953  & ~\pi1126  ;
  assign n63633 = n61931 & n63632 ;
  assign n63634 = n61930 & n63633 ;
  assign n63635 = ~\pi0962  & ~n63634 ;
  assign n63636 = ~n63631 & n63635 ;
  assign n63637 = ~\pi0727  & ~n62838 ;
  assign n63638 = \pi0953  & ~\pi1102  ;
  assign n63639 = n61931 & n63638 ;
  assign n63640 = n61930 & n63639 ;
  assign n63641 = ~\pi0962  & ~n63640 ;
  assign n63642 = ~n63637 & n63641 ;
  assign n63643 = \pi0728  & ~n62838 ;
  assign n63644 = \pi0953  & ~\pi1131  ;
  assign n63645 = n61931 & n63644 ;
  assign n63646 = n61930 & n63645 ;
  assign n63647 = ~\pi0962  & ~n63646 ;
  assign n63648 = ~n63643 & n63647 ;
  assign n63649 = ~\pi0729  & ~n62838 ;
  assign n63650 = \pi0953  & ~\pi1104  ;
  assign n63651 = n61931 & n63650 ;
  assign n63652 = n61930 & n63651 ;
  assign n63653 = ~\pi0962  & ~n63652 ;
  assign n63654 = ~n63649 & n63653 ;
  assign n63655 = ~\pi0730  & ~n62838 ;
  assign n63656 = \pi0953  & ~\pi1106  ;
  assign n63657 = n61931 & n63656 ;
  assign n63658 = n61930 & n63657 ;
  assign n63659 = ~\pi0962  & ~n63658 ;
  assign n63660 = ~n63655 & n63659 ;
  assign n63661 = ~n63536 & ~n63553 ;
  assign n63662 = ~n63539 & ~n63661 ;
  assign n63663 = \pi0795  & ~n63543 ;
  assign n63664 = n63662 & n63663 ;
  assign n63665 = n63535 & n63664 ;
  assign n63666 = \pi0731  & n63665 ;
  assign n63667 = \pi0801  & ~n63533 ;
  assign n63668 = ~\pi0795  & \pi0807  ;
  assign n63669 = ~n63523 & n63668 ;
  assign n63670 = n63667 & n63669 ;
  assign n63671 = ~n63543 & ~n63661 ;
  assign n63672 = ~n63530 & n63671 ;
  assign n63673 = n63670 & n63672 ;
  assign n63674 = n63517 & n63563 ;
  assign n63675 = ~\pi0731  & n63674 ;
  assign n63676 = ~n63673 & n63675 ;
  assign n63677 = \pi0731  & ~n63674 ;
  assign n63678 = ~n63676 & ~n63677 ;
  assign n63679 = ~n63666 & ~n63678 ;
  assign n63680 = \pi0732  & ~n61933 ;
  assign n63681 = ~\pi0953  & ~\pi1128  ;
  assign n63682 = n61931 & n63681 ;
  assign n63683 = n61930 & n63682 ;
  assign n63684 = ~\pi0962  & ~n63683 ;
  assign n63685 = ~n63680 & n63684 ;
  assign n63686 = \pi0316  & ~\pi0592  ;
  assign n63687 = n62182 & n63686 ;
  assign n63688 = n63082 & n63687 ;
  assign n63689 = \pi0375  & n63125 ;
  assign n63690 = \pi0399  & ~\pi0592  ;
  assign n63691 = n62178 & n63690 ;
  assign n63692 = \pi0591  & n63691 ;
  assign n63693 = ~n63689 & ~n63692 ;
  assign n63694 = n9782 & ~n63693 ;
  assign n63695 = ~n63688 & ~n63694 ;
  assign n63696 = ~\pi0200  & ~\pi0308  ;
  assign n63697 = \pi0200  & ~\pi1037  ;
  assign n63698 = ~n63696 & ~n63697 ;
  assign n63699 = ~\pi0199  & ~n63698 ;
  assign n63700 = \pi0199  & ~\pi1047  ;
  assign n63701 = ~n62178 & ~n63700 ;
  assign n63702 = ~n63699 & n63701 ;
  assign n63703 = \pi0424  & n62858 ;
  assign n63704 = n63140 & n63703 ;
  assign n63705 = n10003 & ~n63704 ;
  assign n63706 = ~n63702 & n63705 ;
  assign n63707 = n63695 & n63706 ;
  assign n63708 = \pi0777  & \pi1136  ;
  assign n63709 = ~n62211 & n63708 ;
  assign n63710 = ~\pi0838  & ~\pi1136  ;
  assign n63711 = \pi0737  & \pi1135  ;
  assign n63712 = ~n63710 & ~n63711 ;
  assign n63713 = n62210 & n63712 ;
  assign n63714 = ~n63709 & n63713 ;
  assign n63715 = ~\pi0619  & ~\pi1135  ;
  assign n63716 = ~\pi0648  & \pi1135  ;
  assign n63717 = ~\pi1134  & ~n63716 ;
  assign n63718 = ~n63715 & n63717 ;
  assign n63719 = n63112 & n63718 ;
  assign n63720 = ~n10003 & ~n63719 ;
  assign n63721 = ~n63714 & n63720 ;
  assign n63722 = ~n63707 & ~n63721 ;
  assign n63723 = \pi0734  & ~n62838 ;
  assign n63724 = \pi0953  & ~\pi1119  ;
  assign n63725 = n61931 & n63724 ;
  assign n63726 = n61930 & n63725 ;
  assign n63727 = ~\pi0962  & ~n63726 ;
  assign n63728 = ~n63723 & n63727 ;
  assign n63729 = ~\pi0735  & ~n62838 ;
  assign n63730 = \pi0953  & ~\pi1109  ;
  assign n63731 = n61931 & n63730 ;
  assign n63732 = n61930 & n63731 ;
  assign n63733 = ~\pi0962  & ~n63732 ;
  assign n63734 = ~n63729 & n63733 ;
  assign n63735 = ~\pi0736  & ~n62838 ;
  assign n63736 = \pi0953  & ~\pi1101  ;
  assign n63737 = n61931 & n63736 ;
  assign n63738 = n61930 & n63737 ;
  assign n63739 = ~\pi0962  & ~n63738 ;
  assign n63740 = ~n63735 & n63739 ;
  assign n63741 = \pi0737  & ~n62838 ;
  assign n63742 = \pi0953  & ~\pi1122  ;
  assign n63743 = n61931 & n63742 ;
  assign n63744 = n61930 & n63743 ;
  assign n63745 = ~\pi0962  & ~n63744 ;
  assign n63746 = ~n63741 & n63745 ;
  assign n63747 = \pi0738  & ~n62838 ;
  assign n63748 = \pi0953  & ~\pi1121  ;
  assign n63749 = n61931 & n63748 ;
  assign n63750 = n61930 & n63749 ;
  assign n63751 = ~\pi0962  & ~n63750 ;
  assign n63752 = ~n63747 & n63751 ;
  assign n63753 = ~\pi0952  & n61781 ;
  assign n63754 = n61780 & n63753 ;
  assign n63755 = \pi0739  & ~n63754 ;
  assign n63756 = \pi1060  & \pi1108  ;
  assign n63757 = n61779 & n63756 ;
  assign n63758 = n63753 & n63757 ;
  assign n63759 = ~\pi0966  & ~n63758 ;
  assign n63760 = ~n63755 & n63759 ;
  assign n63761 = ~\pi0741  & ~n63754 ;
  assign n63762 = \pi1060  & \pi1114  ;
  assign n63763 = n61779 & n63762 ;
  assign n63764 = n63753 & n63763 ;
  assign n63765 = ~\pi0966  & ~n63764 ;
  assign n63766 = ~n63761 & n63765 ;
  assign n63767 = ~\pi0742  & ~n63754 ;
  assign n63768 = \pi1060  & \pi1112  ;
  assign n63769 = n61779 & n63768 ;
  assign n63770 = n63753 & n63769 ;
  assign n63771 = ~\pi0966  & ~n63770 ;
  assign n63772 = ~n63767 & n63771 ;
  assign n63773 = \pi0743  & ~n63754 ;
  assign n63774 = \pi1060  & \pi1109  ;
  assign n63775 = n61779 & n63774 ;
  assign n63776 = n63753 & n63775 ;
  assign n63777 = ~\pi0966  & ~n63776 ;
  assign n63778 = ~n63773 & n63777 ;
  assign n63779 = ~\pi0744  & ~n63754 ;
  assign n63780 = \pi1060  & \pi1131  ;
  assign n63781 = n61779 & n63780 ;
  assign n63782 = n63753 & n63781 ;
  assign n63783 = ~\pi0966  & ~n63782 ;
  assign n63784 = ~n63779 & n63783 ;
  assign n63785 = ~\pi0745  & ~n63754 ;
  assign n63786 = \pi1060  & \pi1111  ;
  assign n63787 = n61779 & n63786 ;
  assign n63788 = n63753 & n63787 ;
  assign n63789 = ~\pi0966  & ~n63788 ;
  assign n63790 = ~n63785 & n63789 ;
  assign n63791 = \pi0746  & ~n63754 ;
  assign n63792 = \pi1060  & \pi1104  ;
  assign n63793 = n61779 & n63792 ;
  assign n63794 = n63753 & n63793 ;
  assign n63795 = ~\pi0966  & ~n63794 ;
  assign n63796 = ~n63791 & n63795 ;
  assign n63797 = ~\pi0747  & ~\pi0807  ;
  assign n63798 = \pi0801  & n63797 ;
  assign n63799 = ~n63523 & n63798 ;
  assign n63800 = \pi0773  & n63517 ;
  assign n63801 = ~n63539 & ~n63800 ;
  assign n63802 = n63552 & n63801 ;
  assign n63803 = ~n63799 & ~n63802 ;
  assign n63804 = ~n63516 & n63671 ;
  assign n63805 = n63534 & n63804 ;
  assign n63806 = ~n63803 & n63805 ;
  assign n63807 = ~\pi0747  & ~n63800 ;
  assign n63808 = ~n63674 & ~n63807 ;
  assign n63809 = ~n63806 & n63808 ;
  assign n63810 = \pi0748  & ~n63754 ;
  assign n63811 = \pi1060  & \pi1106  ;
  assign n63812 = n61779 & n63811 ;
  assign n63813 = n63753 & n63812 ;
  assign n63814 = ~\pi0966  & ~n63813 ;
  assign n63815 = ~n63810 & n63814 ;
  assign n63816 = \pi0749  & ~n63754 ;
  assign n63817 = \pi1060  & \pi1105  ;
  assign n63818 = n61779 & n63817 ;
  assign n63819 = n63753 & n63818 ;
  assign n63820 = ~\pi0966  & ~n63819 ;
  assign n63821 = ~n63816 & n63820 ;
  assign n63822 = ~\pi0750  & ~n63754 ;
  assign n63823 = \pi1060  & \pi1130  ;
  assign n63824 = n61779 & n63823 ;
  assign n63825 = n63753 & n63824 ;
  assign n63826 = ~\pi0966  & ~n63825 ;
  assign n63827 = ~n63822 & n63826 ;
  assign n63828 = ~\pi0751  & ~n63754 ;
  assign n63829 = \pi1060  & \pi1123  ;
  assign n63830 = n61779 & n63829 ;
  assign n63831 = n63753 & n63830 ;
  assign n63832 = ~\pi0966  & ~n63831 ;
  assign n63833 = ~n63828 & n63832 ;
  assign n63834 = ~\pi0752  & ~n63754 ;
  assign n63835 = \pi1060  & \pi1124  ;
  assign n63836 = n61779 & n63835 ;
  assign n63837 = n63753 & n63836 ;
  assign n63838 = ~\pi0966  & ~n63837 ;
  assign n63839 = ~n63834 & n63838 ;
  assign n63840 = ~\pi0753  & ~n63754 ;
  assign n63841 = \pi1060  & \pi1117  ;
  assign n63842 = n61779 & n63841 ;
  assign n63843 = n63753 & n63842 ;
  assign n63844 = ~\pi0966  & ~n63843 ;
  assign n63845 = ~n63840 & n63844 ;
  assign n63846 = ~\pi0754  & ~n63754 ;
  assign n63847 = \pi1060  & \pi1118  ;
  assign n63848 = n61779 & n63847 ;
  assign n63849 = n63753 & n63848 ;
  assign n63850 = ~\pi0966  & ~n63849 ;
  assign n63851 = ~n63846 & n63850 ;
  assign n63852 = ~\pi0755  & ~n63754 ;
  assign n63853 = \pi1060  & \pi1120  ;
  assign n63854 = n61779 & n63853 ;
  assign n63855 = n63753 & n63854 ;
  assign n63856 = ~\pi0966  & ~n63855 ;
  assign n63857 = ~n63852 & n63856 ;
  assign n63858 = ~\pi0756  & ~n63754 ;
  assign n63859 = \pi1060  & \pi1119  ;
  assign n63860 = n61779 & n63859 ;
  assign n63861 = n63753 & n63860 ;
  assign n63862 = ~\pi0966  & ~n63861 ;
  assign n63863 = ~n63858 & n63862 ;
  assign n63864 = ~\pi0757  & ~n63754 ;
  assign n63865 = \pi1060  & \pi1113  ;
  assign n63866 = n61779 & n63865 ;
  assign n63867 = n63753 & n63866 ;
  assign n63868 = ~\pi0966  & ~n63867 ;
  assign n63869 = ~n63864 & n63868 ;
  assign n63870 = \pi0758  & ~n63754 ;
  assign n63871 = \pi1060  & \pi1101  ;
  assign n63872 = n61779 & n63871 ;
  assign n63873 = n63753 & n63872 ;
  assign n63874 = ~\pi0966  & ~n63873 ;
  assign n63875 = ~n63870 & n63874 ;
  assign n63876 = \pi0759  & ~n63754 ;
  assign n63877 = \pi1060  & \pi1100  ;
  assign n63878 = n61779 & n63877 ;
  assign n63879 = n63753 & n63878 ;
  assign n63880 = ~\pi0966  & ~n63879 ;
  assign n63881 = ~n63876 & n63880 ;
  assign n63882 = ~\pi0760  & ~n63754 ;
  assign n63883 = \pi1060  & \pi1115  ;
  assign n63884 = n61779 & n63883 ;
  assign n63885 = n63753 & n63884 ;
  assign n63886 = ~\pi0966  & ~n63885 ;
  assign n63887 = ~n63882 & n63886 ;
  assign n63888 = ~\pi0761  & ~n63754 ;
  assign n63889 = \pi1060  & \pi1121  ;
  assign n63890 = n61779 & n63889 ;
  assign n63891 = n63753 & n63890 ;
  assign n63892 = ~\pi0966  & ~n63891 ;
  assign n63893 = ~n63888 & n63892 ;
  assign n63894 = ~\pi0762  & ~n63754 ;
  assign n63895 = \pi1060  & \pi1129  ;
  assign n63896 = n61779 & n63895 ;
  assign n63897 = n63753 & n63896 ;
  assign n63898 = ~\pi0966  & ~n63897 ;
  assign n63899 = ~n63894 & n63898 ;
  assign n63900 = \pi0763  & ~n63754 ;
  assign n63901 = \pi1060  & \pi1103  ;
  assign n63902 = n61779 & n63901 ;
  assign n63903 = n63753 & n63902 ;
  assign n63904 = ~\pi0966  & ~n63903 ;
  assign n63905 = ~n63900 & n63904 ;
  assign n63906 = \pi0764  & ~n63754 ;
  assign n63907 = \pi1060  & \pi1107  ;
  assign n63908 = n61779 & n63907 ;
  assign n63909 = n63753 & n63908 ;
  assign n63910 = ~\pi0966  & ~n63909 ;
  assign n63911 = ~n63906 & n63910 ;
  assign n63912 = ~\pi0765  & \pi0945  ;
  assign n63913 = n63535 & ~n63539 ;
  assign n63914 = \pi0945  & ~n63516 ;
  assign n63915 = n63671 & n63914 ;
  assign n63916 = n63913 & n63915 ;
  assign n63917 = ~n63912 & ~n63916 ;
  assign n63918 = ~\pi0765  & ~n63666 ;
  assign n63919 = ~\pi0945  & ~n63918 ;
  assign n63920 = n63542 & ~n63661 ;
  assign n63921 = ~n63539 & n63920 ;
  assign n63922 = n63535 & n63921 ;
  assign n63923 = ~n63551 & ~n63553 ;
  assign n63924 = ~n63922 & n63923 ;
  assign n63925 = \pi0747  & \pi0807  ;
  assign n63926 = ~n63523 & n63925 ;
  assign n63927 = ~\pi0765  & ~\pi0773  ;
  assign n63928 = ~n63529 & n63927 ;
  assign n63929 = ~n63532 & n63928 ;
  assign n63930 = ~n63926 & n63929 ;
  assign n63931 = n63541 & ~n63930 ;
  assign n63932 = n63913 & n63931 ;
  assign n63933 = \pi0721  & n63541 ;
  assign n63934 = ~n63922 & ~n63933 ;
  assign n63935 = ~n63932 & n63934 ;
  assign n63936 = ~n63924 & ~n63935 ;
  assign n63937 = ~\pi0945  & n63514 ;
  assign n63938 = n63936 & n63937 ;
  assign n63939 = ~n63919 & ~n63938 ;
  assign n63940 = n63917 & n63939 ;
  assign n63941 = \pi0766  & ~n63754 ;
  assign n63942 = \pi1060  & \pi1110  ;
  assign n63943 = n61779 & n63942 ;
  assign n63944 = n63753 & n63943 ;
  assign n63945 = ~\pi0966  & ~n63944 ;
  assign n63946 = ~n63941 & n63945 ;
  assign n63947 = ~\pi0767  & ~n63754 ;
  assign n63948 = \pi1060  & \pi1116  ;
  assign n63949 = n61779 & n63948 ;
  assign n63950 = n63753 & n63949 ;
  assign n63951 = ~\pi0966  & ~n63950 ;
  assign n63952 = ~n63947 & n63951 ;
  assign n63953 = ~\pi0768  & ~n63754 ;
  assign n63954 = \pi1060  & \pi1125  ;
  assign n63955 = n61779 & n63954 ;
  assign n63956 = n63753 & n63955 ;
  assign n63957 = ~\pi0966  & ~n63956 ;
  assign n63958 = ~n63953 & n63957 ;
  assign n63959 = \pi0794  & ~n63530 ;
  assign n63960 = n63671 & n63959 ;
  assign n63961 = ~\pi0775  & \pi0795  ;
  assign n63962 = ~n63539 & n63961 ;
  assign n63963 = n63527 & n63962 ;
  assign n63964 = n63960 & n63963 ;
  assign n63965 = \pi0795  & ~n63539 ;
  assign n63966 = n63920 & n63965 ;
  assign n63967 = n63535 & n63966 ;
  assign n63968 = \pi0775  & n63563 ;
  assign n63969 = ~\pi0769  & ~n63968 ;
  assign n63970 = n63518 & ~n63565 ;
  assign n63971 = ~n63969 & n63970 ;
  assign n63972 = ~n63967 & n63971 ;
  assign n63973 = ~n63964 & n63972 ;
  assign n63974 = ~n63516 & ~n63539 ;
  assign n63975 = n63527 & n63974 ;
  assign n63976 = n63960 & n63975 ;
  assign n63977 = \pi0769  & ~n63518 ;
  assign n63978 = ~n63976 & n63977 ;
  assign n63979 = ~n63973 & ~n63978 ;
  assign n63980 = ~\pi0770  & ~n63754 ;
  assign n63981 = \pi1060  & \pi1126  ;
  assign n63982 = n61779 & n63981 ;
  assign n63983 = n63753 & n63982 ;
  assign n63984 = ~\pi0966  & ~n63983 ;
  assign n63985 = ~n63980 & n63984 ;
  assign n63986 = ~n63542 & ~n63933 ;
  assign n63987 = ~n63932 & n63986 ;
  assign n63988 = n63535 & n63662 ;
  assign n63989 = n63514 & n63988 ;
  assign n63990 = ~n63987 & n63989 ;
  assign n63991 = n63515 & ~n63543 ;
  assign n63992 = n63662 & n63991 ;
  assign n63993 = n63535 & n63992 ;
  assign n63994 = ~\pi0945  & \pi0987  ;
  assign n63995 = ~n63993 & n63994 ;
  assign n63996 = ~n63990 & n63995 ;
  assign n63997 = n63804 & n63913 ;
  assign n63998 = \pi0771  & \pi0945  ;
  assign n63999 = ~n63997 & n63998 ;
  assign n64000 = ~n63996 & ~n63999 ;
  assign n64001 = \pi0772  & ~n63754 ;
  assign n64002 = \pi1060  & \pi1102  ;
  assign n64003 = n61779 & n64002 ;
  assign n64004 = n63753 & n64003 ;
  assign n64005 = ~\pi0966  & ~n64004 ;
  assign n64006 = ~n64001 & n64005 ;
  assign n64007 = ~n63990 & ~n63993 ;
  assign n64008 = n63535 & n63537 ;
  assign n64009 = ~n64007 & n64008 ;
  assign n64010 = \pi0801  & ~n63516 ;
  assign n64011 = n63671 & n64010 ;
  assign n64012 = n63535 & n64011 ;
  assign n64013 = \pi0773  & ~n63517 ;
  assign n64014 = ~n64012 & n64013 ;
  assign n64015 = ~\pi0773  & n63517 ;
  assign n64016 = ~n64014 & ~n64015 ;
  assign n64017 = ~n64009 & ~n64016 ;
  assign n64018 = ~\pi0774  & ~n63754 ;
  assign n64019 = \pi1060  & \pi1127  ;
  assign n64020 = n61779 & n64019 ;
  assign n64021 = n63753 & n64020 ;
  assign n64022 = ~\pi0966  & ~n64021 ;
  assign n64023 = ~n64018 & n64022 ;
  assign n64024 = \pi0765  & \pi0771  ;
  assign n64025 = n63563 & n64024 ;
  assign n64026 = ~n63665 & ~n64025 ;
  assign n64027 = \pi0731  & ~\pi0945  ;
  assign n64028 = \pi0775  & n64027 ;
  assign n64029 = ~n64026 & n64028 ;
  assign n64030 = \pi0775  & ~n63997 ;
  assign n64031 = \pi0801  & ~\pi0816  ;
  assign n64032 = \pi0795  & \pi0800  ;
  assign n64033 = n64031 & n64032 ;
  assign n64034 = ~n63533 & n64033 ;
  assign n64035 = ~\pi0775  & ~n63661 ;
  assign n64036 = n63527 & n64035 ;
  assign n64037 = n64034 & n64036 ;
  assign n64038 = ~\pi0775  & ~n64025 ;
  assign n64039 = n64027 & ~n64038 ;
  assign n64040 = ~n64037 & n64039 ;
  assign n64041 = ~n64030 & ~n64040 ;
  assign n64042 = ~n64029 & ~n64041 ;
  assign n64043 = ~\pi0776  & ~n63754 ;
  assign n64044 = \pi1060  & \pi1128  ;
  assign n64045 = n61779 & n64044 ;
  assign n64046 = n63753 & n64045 ;
  assign n64047 = ~\pi0966  & ~n64046 ;
  assign n64048 = ~n64043 & n64047 ;
  assign n64049 = ~\pi0777  & ~n63754 ;
  assign n64050 = \pi1060  & \pi1122  ;
  assign n64051 = n61779 & n64050 ;
  assign n64052 = n63753 & n64051 ;
  assign n64053 = ~\pi0966  & ~n64052 ;
  assign n64054 = ~n64049 & n64053 ;
  assign n64055 = ~\pi1046  & ~\pi1083  ;
  assign n64056 = \pi1085  & n64055 ;
  assign n64057 = \pi0832  & \pi0956  ;
  assign n64058 = ~\pi0968  & n64057 ;
  assign n64059 = n64056 & n64058 ;
  assign n64060 = \pi0778  & ~n64059 ;
  assign n64061 = \pi1085  & \pi1100  ;
  assign n64062 = n64055 & n64061 ;
  assign n64063 = n64058 & n64062 ;
  assign n64064 = ~n64060 & ~n64063 ;
  assign n64065 = \pi0779  & ~n61865 ;
  assign n64066 = \pi0780  & ~n61756 ;
  assign n64067 = \pi0781  & ~n64059 ;
  assign n64068 = \pi1085  & \pi1101  ;
  assign n64069 = n64055 & n64068 ;
  assign n64070 = n64058 & n64069 ;
  assign n64071 = ~n64067 & ~n64070 ;
  assign n64072 = ~\pi0057  & ~\pi0882  ;
  assign n64073 = n6848 & n64072 ;
  assign n64074 = ~n55622 & ~n61797 ;
  assign n64075 = ~n64073 & n64074 ;
  assign n64076 = \pi0783  & ~n64059 ;
  assign n64077 = \pi1085  & \pi1109  ;
  assign n64078 = n64055 & n64077 ;
  assign n64079 = n64058 & n64078 ;
  assign n64080 = ~n64076 & ~n64079 ;
  assign n64081 = \pi0784  & ~n64059 ;
  assign n64082 = \pi1085  & \pi1110  ;
  assign n64083 = n64055 & n64082 ;
  assign n64084 = n64058 & n64083 ;
  assign n64085 = ~n64081 & ~n64084 ;
  assign n64086 = \pi0785  & ~n64059 ;
  assign n64087 = \pi1085  & \pi1102  ;
  assign n64088 = n64055 & n64087 ;
  assign n64089 = n64058 & n64088 ;
  assign n64090 = ~n64086 & ~n64089 ;
  assign n64091 = \pi0024  & ~\pi0954  ;
  assign n64092 = \pi0786  & \pi0954  ;
  assign n64093 = ~n64091 & ~n64092 ;
  assign n64094 = \pi0787  & ~n64059 ;
  assign n64095 = \pi1085  & \pi1104  ;
  assign n64096 = n64055 & n64095 ;
  assign n64097 = n64058 & n64096 ;
  assign n64098 = ~n64094 & ~n64097 ;
  assign n64099 = \pi0788  & ~n64059 ;
  assign n64100 = \pi1085  & \pi1105  ;
  assign n64101 = n64055 & n64100 ;
  assign n64102 = n64058 & n64101 ;
  assign n64103 = ~n64099 & ~n64102 ;
  assign n64104 = \pi0789  & ~n64059 ;
  assign n64105 = \pi1085  & \pi1106  ;
  assign n64106 = n64055 & n64105 ;
  assign n64107 = n64058 & n64106 ;
  assign n64108 = ~n64104 & ~n64107 ;
  assign n64109 = \pi0790  & ~n64059 ;
  assign n64110 = \pi1085  & \pi1107  ;
  assign n64111 = n64055 & n64110 ;
  assign n64112 = n64058 & n64111 ;
  assign n64113 = ~n64109 & ~n64112 ;
  assign n64114 = \pi0791  & ~n64059 ;
  assign n64115 = \pi1085  & \pi1108  ;
  assign n64116 = n64055 & n64115 ;
  assign n64117 = n64058 & n64116 ;
  assign n64118 = ~n64114 & ~n64117 ;
  assign n64119 = \pi0792  & ~n64059 ;
  assign n64120 = \pi1085  & \pi1103  ;
  assign n64121 = n64055 & n64120 ;
  assign n64122 = n64058 & n64121 ;
  assign n64123 = ~n64119 & ~n64122 ;
  assign n64124 = \pi0968  & \pi1085  ;
  assign n64125 = n64055 & n64124 ;
  assign n64126 = n64057 & n64125 ;
  assign n64127 = \pi0794  & ~n64126 ;
  assign n64128 = \pi0968  & \pi1130  ;
  assign n64129 = n64057 & n64128 ;
  assign n64130 = n64056 & n64129 ;
  assign n64131 = ~n64127 & ~n64130 ;
  assign n64132 = \pi0795  & ~n64126 ;
  assign n64133 = \pi0968  & \pi1128  ;
  assign n64134 = n64057 & n64133 ;
  assign n64135 = n64056 & n64134 ;
  assign n64136 = ~n64132 & ~n64135 ;
  assign n64137 = ~\pi0282  & n62141 ;
  assign n64138 = \pi0278  & \pi0279  ;
  assign n64139 = ~\pi0280  & n64138 ;
  assign n64140 = \pi0266  & ~\pi0269  ;
  assign n64141 = ~\pi0281  & n64140 ;
  assign n64142 = n64139 & n64141 ;
  assign n64143 = n64137 & n64142 ;
  assign n64144 = \pi0264  & ~n64143 ;
  assign n64145 = ~\pi0264  & n64137 ;
  assign n64146 = n64142 & n64145 ;
  assign n64147 = ~n64144 & ~n64146 ;
  assign n64148 = \pi0798  & ~n64126 ;
  assign n64149 = \pi0968  & \pi1124  ;
  assign n64150 = n64057 & n64149 ;
  assign n64151 = n64056 & n64150 ;
  assign n64152 = ~n64148 & ~n64151 ;
  assign n64153 = \pi0799  & ~n64126 ;
  assign n64154 = \pi0968  & ~\pi1107  ;
  assign n64155 = n64057 & n64154 ;
  assign n64156 = n64056 & n64155 ;
  assign n64157 = ~n64153 & ~n64156 ;
  assign n64158 = \pi0800  & ~n64126 ;
  assign n64159 = \pi0968  & \pi1125  ;
  assign n64160 = n64057 & n64159 ;
  assign n64161 = n64056 & n64160 ;
  assign n64162 = ~n64158 & ~n64161 ;
  assign n64163 = \pi0801  & ~n64126 ;
  assign n64164 = \pi0968  & \pi1126  ;
  assign n64165 = n64057 & n64164 ;
  assign n64166 = n64056 & n64165 ;
  assign n64167 = ~n64163 & ~n64166 ;
  assign n64168 = \pi0803  & ~n64126 ;
  assign n64169 = \pi0968  & ~\pi1106  ;
  assign n64170 = n64057 & n64169 ;
  assign n64171 = n64056 & n64170 ;
  assign n64172 = ~n64168 & ~n64171 ;
  assign n64173 = \pi0804  & ~n64126 ;
  assign n64174 = \pi0968  & \pi1109  ;
  assign n64175 = n64057 & n64174 ;
  assign n64176 = n64056 & n64175 ;
  assign n64177 = ~n64173 & ~n64176 ;
  assign n64178 = ~\pi0270  & ~\pi0282  ;
  assign n64179 = ~\pi0281  & n64178 ;
  assign n64180 = n62140 & n64179 ;
  assign n64181 = n62140 & n62142 ;
  assign n64182 = \pi0270  & ~n64181 ;
  assign n64183 = ~n64180 & ~n64182 ;
  assign n64184 = \pi0807  & ~n64126 ;
  assign n64185 = \pi0968  & \pi1127  ;
  assign n64186 = n64057 & n64185 ;
  assign n64187 = n64056 & n64186 ;
  assign n64188 = ~n64184 & ~n64187 ;
  assign n64189 = \pi0808  & ~n64126 ;
  assign n64190 = \pi0968  & \pi1101  ;
  assign n64191 = n64057 & n64190 ;
  assign n64192 = n64056 & n64191 ;
  assign n64193 = ~n64189 & ~n64192 ;
  assign n64194 = \pi0809  & ~n64126 ;
  assign n64195 = \pi0968  & ~\pi1103  ;
  assign n64196 = n64057 & n64195 ;
  assign n64197 = n64056 & n64196 ;
  assign n64198 = ~n64194 & ~n64197 ;
  assign n64199 = \pi0810  & ~n64126 ;
  assign n64200 = \pi0968  & \pi1108  ;
  assign n64201 = n64057 & n64200 ;
  assign n64202 = n64056 & n64201 ;
  assign n64203 = ~n64199 & ~n64202 ;
  assign n64204 = \pi0811  & ~n64126 ;
  assign n64205 = \pi0968  & \pi1102  ;
  assign n64206 = n64057 & n64205 ;
  assign n64207 = n64056 & n64206 ;
  assign n64208 = ~n64204 & ~n64207 ;
  assign n64209 = \pi0812  & ~n64126 ;
  assign n64210 = \pi0968  & ~\pi1104  ;
  assign n64211 = n64057 & n64210 ;
  assign n64212 = n64056 & n64211 ;
  assign n64213 = ~n64209 & ~n64212 ;
  assign n64214 = \pi0813  & ~n64126 ;
  assign n64215 = \pi0968  & \pi1131  ;
  assign n64216 = n64057 & n64215 ;
  assign n64217 = n64056 & n64216 ;
  assign n64218 = ~n64214 & ~n64217 ;
  assign n64219 = \pi0814  & ~n64126 ;
  assign n64220 = \pi0968  & ~\pi1105  ;
  assign n64221 = n64057 & n64220 ;
  assign n64222 = n64056 & n64221 ;
  assign n64223 = ~n64219 & ~n64222 ;
  assign n64224 = \pi0815  & ~n64126 ;
  assign n64225 = \pi0968  & \pi1110  ;
  assign n64226 = n64057 & n64225 ;
  assign n64227 = n64056 & n64226 ;
  assign n64228 = ~n64224 & ~n64227 ;
  assign n64229 = \pi0816  & ~n64126 ;
  assign n64230 = \pi0968  & \pi1129  ;
  assign n64231 = n64057 & n64230 ;
  assign n64232 = n64056 & n64231 ;
  assign n64233 = ~n64229 & ~n64232 ;
  assign n64234 = ~\pi0280  & n62138 ;
  assign n64235 = \pi0269  & ~n64234 ;
  assign n64236 = ~n62140 & ~n64235 ;
  assign n64237 = n10003 & n16862 ;
  assign n64238 = ~n17154 & ~n64237 ;
  assign n64239 = ~\pi0264  & n62148 ;
  assign n64240 = \pi0265  & ~n64239 ;
  assign n64241 = ~n62150 & ~n64240 ;
  assign n64242 = \pi0277  & ~n64180 ;
  assign n64243 = ~n62148 & ~n64242 ;
  assign n64244 = ~\pi0811  & ~\pi0893  ;
  assign n64245 = ~\pi0982  & ~n6704 ;
  assign n64246 = n8543 & n10003 ;
  assign n64247 = ~n64245 & ~n64246 ;
  assign n64248 = n6809 & ~n64247 ;
  assign n64249 = \pi0123  & ~\pi0223  ;
  assign n64250 = n2165 & n64249 ;
  assign n64251 = ~\pi1127  & ~\pi1131  ;
  assign n64252 = ~n64250 & ~n64251 ;
  assign n64253 = ~\pi0825  & n64250 ;
  assign n64254 = ~n64252 & ~n64253 ;
  assign n64255 = \pi1127  & \pi1131  ;
  assign n64256 = ~n64250 & n64255 ;
  assign n64257 = ~n64254 & ~n64256 ;
  assign n64258 = \pi1124  & ~\pi1130  ;
  assign n64259 = ~\pi1124  & \pi1130  ;
  assign n64260 = ~n64258 & ~n64259 ;
  assign n64261 = ~\pi1128  & ~\pi1129  ;
  assign n64262 = \pi1128  & \pi1129  ;
  assign n64263 = ~n64261 & ~n64262 ;
  assign n64264 = ~\pi1125  & ~\pi1126  ;
  assign n64265 = \pi1125  & \pi1126  ;
  assign n64266 = ~n64264 & ~n64265 ;
  assign n64267 = ~n64263 & ~n64266 ;
  assign n64268 = n64263 & n64266 ;
  assign n64269 = ~n64267 & ~n64268 ;
  assign n64270 = n64260 & ~n64269 ;
  assign n64271 = ~n64260 & n64269 ;
  assign n64272 = ~n64270 & ~n64271 ;
  assign n64273 = ~n64257 & ~n64272 ;
  assign n64274 = ~n64256 & n64260 ;
  assign n64275 = n64269 & n64274 ;
  assign n64276 = ~n64256 & ~n64260 ;
  assign n64277 = ~n64269 & n64276 ;
  assign n64278 = ~n64275 & ~n64277 ;
  assign n64279 = ~n64250 & n64251 ;
  assign n64280 = ~n64253 & ~n64279 ;
  assign n64281 = ~n64278 & n64280 ;
  assign n64282 = ~n64273 & ~n64281 ;
  assign n64283 = ~\pi1122  & ~\pi1123  ;
  assign n64284 = ~n64250 & ~n64283 ;
  assign n64285 = ~\pi0826  & n64250 ;
  assign n64286 = ~n64284 & ~n64285 ;
  assign n64287 = \pi1122  & \pi1123  ;
  assign n64288 = ~n64250 & n64287 ;
  assign n64289 = ~n64286 & ~n64288 ;
  assign n64290 = \pi1118  & ~\pi1119  ;
  assign n64291 = ~\pi1118  & \pi1119  ;
  assign n64292 = ~n64290 & ~n64291 ;
  assign n64293 = ~\pi1120  & ~\pi1121  ;
  assign n64294 = \pi1120  & \pi1121  ;
  assign n64295 = ~n64293 & ~n64294 ;
  assign n64296 = ~\pi1116  & ~\pi1117  ;
  assign n64297 = \pi1116  & \pi1117  ;
  assign n64298 = ~n64296 & ~n64297 ;
  assign n64299 = ~n64295 & ~n64298 ;
  assign n64300 = n64295 & n64298 ;
  assign n64301 = ~n64299 & ~n64300 ;
  assign n64302 = n64292 & ~n64301 ;
  assign n64303 = ~n64292 & n64301 ;
  assign n64304 = ~n64302 & ~n64303 ;
  assign n64305 = ~n64289 & ~n64304 ;
  assign n64306 = ~n64288 & n64292 ;
  assign n64307 = n64301 & n64306 ;
  assign n64308 = ~n64288 & ~n64292 ;
  assign n64309 = ~n64301 & n64308 ;
  assign n64310 = ~n64307 & ~n64309 ;
  assign n64311 = ~n64250 & n64283 ;
  assign n64312 = ~n64285 & ~n64311 ;
  assign n64313 = ~n64310 & n64312 ;
  assign n64314 = ~n64305 & ~n64313 ;
  assign n64315 = ~\pi1100  & ~\pi1107  ;
  assign n64316 = ~n64250 & ~n64315 ;
  assign n64317 = ~\pi0827  & n64250 ;
  assign n64318 = ~n64316 & ~n64317 ;
  assign n64319 = \pi1100  & \pi1107  ;
  assign n64320 = ~n64250 & n64319 ;
  assign n64321 = ~n64318 & ~n64320 ;
  assign n64322 = \pi1103  & ~\pi1105  ;
  assign n64323 = ~\pi1103  & \pi1105  ;
  assign n64324 = ~n64322 & ~n64323 ;
  assign n64325 = ~\pi1101  & ~\pi1102  ;
  assign n64326 = \pi1101  & \pi1102  ;
  assign n64327 = ~n64325 & ~n64326 ;
  assign n64328 = ~\pi1104  & ~\pi1106  ;
  assign n64329 = \pi1104  & \pi1106  ;
  assign n64330 = ~n64328 & ~n64329 ;
  assign n64331 = ~n64327 & ~n64330 ;
  assign n64332 = n64327 & n64330 ;
  assign n64333 = ~n64331 & ~n64332 ;
  assign n64334 = n64324 & ~n64333 ;
  assign n64335 = ~n64324 & n64333 ;
  assign n64336 = ~n64334 & ~n64335 ;
  assign n64337 = ~n64321 & ~n64336 ;
  assign n64338 = ~n64320 & n64324 ;
  assign n64339 = n64333 & n64338 ;
  assign n64340 = ~n64320 & ~n64324 ;
  assign n64341 = ~n64333 & n64340 ;
  assign n64342 = ~n64339 & ~n64341 ;
  assign n64343 = ~n64250 & n64315 ;
  assign n64344 = ~n64317 & ~n64343 ;
  assign n64345 = ~n64342 & n64344 ;
  assign n64346 = ~n64337 & ~n64345 ;
  assign n64347 = ~\pi1114  & ~\pi1115  ;
  assign n64348 = ~n64250 & ~n64347 ;
  assign n64349 = ~\pi0828  & n64250 ;
  assign n64350 = ~n64348 & ~n64349 ;
  assign n64351 = \pi1114  & \pi1115  ;
  assign n64352 = ~n64250 & n64351 ;
  assign n64353 = ~n64350 & ~n64352 ;
  assign n64354 = \pi1110  & ~\pi1111  ;
  assign n64355 = ~\pi1110  & \pi1111  ;
  assign n64356 = ~n64354 & ~n64355 ;
  assign n64357 = ~\pi1112  & ~\pi1113  ;
  assign n64358 = \pi1112  & \pi1113  ;
  assign n64359 = ~n64357 & ~n64358 ;
  assign n64360 = ~\pi1108  & ~\pi1109  ;
  assign n64361 = \pi1108  & \pi1109  ;
  assign n64362 = ~n64360 & ~n64361 ;
  assign n64363 = ~n64359 & ~n64362 ;
  assign n64364 = n64359 & n64362 ;
  assign n64365 = ~n64363 & ~n64364 ;
  assign n64366 = n64356 & ~n64365 ;
  assign n64367 = ~n64356 & n64365 ;
  assign n64368 = ~n64366 & ~n64367 ;
  assign n64369 = ~n64353 & ~n64368 ;
  assign n64370 = ~n64352 & n64356 ;
  assign n64371 = n64365 & n64370 ;
  assign n64372 = ~n64352 & ~n64356 ;
  assign n64373 = ~n64365 & n64372 ;
  assign n64374 = ~n64371 & ~n64373 ;
  assign n64375 = ~n64250 & n64347 ;
  assign n64376 = ~n64349 & ~n64375 ;
  assign n64377 = ~n64374 & n64376 ;
  assign n64378 = ~n64369 & ~n64377 ;
  assign n64379 = ~\pi0951  & \pi1092  ;
  assign n64380 = \pi1092  & n6703 ;
  assign n64381 = n63610 & n64380 ;
  assign n64382 = ~n64379 & ~n64381 ;
  assign n64383 = n64139 & n64140 ;
  assign n64384 = \pi0281  & ~n64383 ;
  assign n64385 = ~n64142 & ~n64384 ;
  assign n64386 = ~\pi0832  & \pi1091  ;
  assign n64387 = \pi1162  & n64386 ;
  assign n64388 = n10011 & n64387 ;
  assign n64389 = \pi0833  & ~n1689 ;
  assign n64390 = ~n1695 & ~n64389 ;
  assign n64391 = \pi0946  & n1689 ;
  assign n64392 = ~\pi0281  & n62140 ;
  assign n64393 = \pi0282  & ~n64392 ;
  assign n64394 = ~n64181 & ~n64393 ;
  assign n64395 = ~\pi0955  & \pi1049  ;
  assign n64396 = \pi0837  & \pi0955  ;
  assign n64397 = ~n64395 & ~n64396 ;
  assign n64398 = ~\pi0955  & \pi1047  ;
  assign n64399 = \pi0838  & \pi0955  ;
  assign n64400 = ~n64398 & ~n64399 ;
  assign n64401 = ~\pi0955  & \pi1074  ;
  assign n64402 = \pi0839  & \pi0955  ;
  assign n64403 = ~n64401 & ~n64402 ;
  assign n64404 = \pi0840  & ~n1689 ;
  assign n64405 = \pi1196  & n1689 ;
  assign n64406 = ~n64404 & ~n64405 ;
  assign n64407 = ~\pi0033  & n11102 ;
  assign n64408 = ~\pi0955  & \pi1035  ;
  assign n64409 = \pi0842  & \pi0955  ;
  assign n64410 = ~n64408 & ~n64409 ;
  assign n64411 = ~\pi0955  & \pi1079  ;
  assign n64412 = \pi0843  & \pi0955  ;
  assign n64413 = ~n64411 & ~n64412 ;
  assign n64414 = ~\pi0955  & \pi1078  ;
  assign n64415 = \pi0844  & \pi0955  ;
  assign n64416 = ~n64414 & ~n64415 ;
  assign n64417 = ~\pi0955  & \pi1043  ;
  assign n64418 = \pi0845  & \pi0955  ;
  assign n64419 = ~n64417 & ~n64418 ;
  assign n64420 = \pi0846  & ~n56376 ;
  assign n64421 = \pi1134  & n56376 ;
  assign n64422 = ~n64420 & ~n64421 ;
  assign n64423 = ~\pi0955  & \pi1055  ;
  assign n64424 = \pi0847  & \pi0955  ;
  assign n64425 = ~n64423 & ~n64424 ;
  assign n64426 = ~\pi0955  & \pi1039  ;
  assign n64427 = \pi0848  & \pi0955  ;
  assign n64428 = ~n64426 & ~n64427 ;
  assign n64429 = \pi0849  & ~n1689 ;
  assign n64430 = \pi1198  & n1689 ;
  assign n64431 = ~n64429 & ~n64430 ;
  assign n64432 = ~\pi0955  & \pi1048  ;
  assign n64433 = \pi0850  & \pi0955  ;
  assign n64434 = ~n64432 & ~n64433 ;
  assign n64435 = ~\pi0955  & \pi1045  ;
  assign n64436 = \pi0851  & \pi0955  ;
  assign n64437 = ~n64435 & ~n64436 ;
  assign n64438 = ~\pi0955  & \pi1062  ;
  assign n64439 = \pi0852  & \pi0955  ;
  assign n64440 = ~n64438 & ~n64439 ;
  assign n64441 = ~\pi0955  & \pi1080  ;
  assign n64442 = \pi0853  & \pi0955  ;
  assign n64443 = ~n64441 & ~n64442 ;
  assign n64444 = ~\pi0955  & \pi1051  ;
  assign n64445 = \pi0854  & \pi0955  ;
  assign n64446 = ~n64444 & ~n64445 ;
  assign n64447 = ~\pi0955  & \pi1065  ;
  assign n64448 = \pi0855  & \pi0955  ;
  assign n64449 = ~n64447 & ~n64448 ;
  assign n64450 = ~\pi0955  & \pi1067  ;
  assign n64451 = \pi0856  & \pi0955  ;
  assign n64452 = ~n64450 & ~n64451 ;
  assign n64453 = ~\pi0955  & \pi1058  ;
  assign n64454 = \pi0857  & \pi0955  ;
  assign n64455 = ~n64453 & ~n64454 ;
  assign n64456 = ~\pi0955  & \pi1087  ;
  assign n64457 = \pi0858  & \pi0955  ;
  assign n64458 = ~n64456 & ~n64457 ;
  assign n64459 = ~\pi0955  & \pi1070  ;
  assign n64460 = \pi0859  & \pi0955  ;
  assign n64461 = ~n64459 & ~n64460 ;
  assign n64462 = ~\pi0955  & \pi1076  ;
  assign n64463 = \pi0860  & \pi0955  ;
  assign n64464 = ~n64462 & ~n64463 ;
  assign n64465 = \pi1093  & \pi1141  ;
  assign n64466 = \pi0861  & ~\pi1093  ;
  assign n64467 = ~n64465 & ~n64466 ;
  assign n64468 = ~\pi0228  & ~n64467 ;
  assign n64469 = \pi0123  & ~\pi0861  ;
  assign n64470 = ~\pi0123  & ~\pi1141  ;
  assign n64471 = \pi0228  & ~n64470 ;
  assign n64472 = ~n64469 & n64471 ;
  assign n64473 = ~n64468 & ~n64472 ;
  assign n64474 = \pi0862  & ~n56376 ;
  assign n64475 = \pi1139  & n56376 ;
  assign n64476 = ~n64474 & ~n64475 ;
  assign n64477 = \pi0863  & ~n1689 ;
  assign n64478 = \pi1199  & n1689 ;
  assign n64479 = ~n64477 & ~n64478 ;
  assign n64480 = \pi0864  & ~n1689 ;
  assign n64481 = \pi1197  & n1689 ;
  assign n64482 = ~n64480 & ~n64481 ;
  assign n64483 = ~\pi0955  & \pi1040  ;
  assign n64484 = \pi0865  & \pi0955  ;
  assign n64485 = ~n64483 & ~n64484 ;
  assign n64486 = ~\pi0955  & \pi1053  ;
  assign n64487 = \pi0866  & \pi0955  ;
  assign n64488 = ~n64486 & ~n64487 ;
  assign n64489 = ~\pi0955  & \pi1057  ;
  assign n64490 = \pi0867  & \pi0955  ;
  assign n64491 = ~n64489 & ~n64490 ;
  assign n64492 = ~\pi0955  & \pi1063  ;
  assign n64493 = \pi0868  & \pi0955  ;
  assign n64494 = ~n64492 & ~n64493 ;
  assign n64495 = \pi1093  & \pi1140  ;
  assign n64496 = \pi0869  & ~\pi1093  ;
  assign n64497 = ~n64495 & ~n64496 ;
  assign n64498 = ~\pi0228  & ~n64497 ;
  assign n64499 = \pi0123  & ~\pi0869  ;
  assign n64500 = ~\pi0123  & ~\pi1140  ;
  assign n64501 = \pi0228  & ~n64500 ;
  assign n64502 = ~n64499 & n64501 ;
  assign n64503 = ~n64498 & ~n64502 ;
  assign n64504 = ~\pi0955  & \pi1069  ;
  assign n64505 = \pi0870  & \pi0955  ;
  assign n64506 = ~n64504 & ~n64505 ;
  assign n64507 = ~\pi0955  & \pi1072  ;
  assign n64508 = \pi0871  & \pi0955  ;
  assign n64509 = ~n64507 & ~n64508 ;
  assign n64510 = ~\pi0955  & \pi1084  ;
  assign n64511 = \pi0872  & \pi0955  ;
  assign n64512 = ~n64510 & ~n64511 ;
  assign n64513 = ~\pi0955  & \pi1044  ;
  assign n64514 = \pi0873  & \pi0955  ;
  assign n64515 = ~n64513 & ~n64514 ;
  assign n64516 = ~\pi0955  & \pi1036  ;
  assign n64517 = \pi0874  & \pi0955  ;
  assign n64518 = ~n64516 & ~n64517 ;
  assign n64519 = \pi1093  & ~\pi1136  ;
  assign n64520 = ~\pi0875  & ~\pi1093  ;
  assign n64521 = ~n64519 & ~n64520 ;
  assign n64522 = ~\pi0228  & ~n64521 ;
  assign n64523 = \pi0123  & \pi0875  ;
  assign n64524 = ~\pi0123  & \pi1136  ;
  assign n64525 = \pi0228  & ~n64524 ;
  assign n64526 = ~n64523 & n64525 ;
  assign n64527 = ~n64522 & ~n64526 ;
  assign n64528 = ~\pi0955  & \pi1037  ;
  assign n64529 = \pi0876  & \pi0955  ;
  assign n64530 = ~n64528 & ~n64529 ;
  assign n64531 = \pi1093  & \pi1138  ;
  assign n64532 = \pi0877  & ~\pi1093  ;
  assign n64533 = ~n64531 & ~n64532 ;
  assign n64534 = ~\pi0228  & ~n64533 ;
  assign n64535 = \pi0123  & ~\pi0877  ;
  assign n64536 = ~\pi0123  & ~\pi1138  ;
  assign n64537 = \pi0228  & ~n64536 ;
  assign n64538 = ~n64535 & n64537 ;
  assign n64539 = ~n64534 & ~n64538 ;
  assign n64540 = \pi1093  & \pi1137  ;
  assign n64541 = \pi0878  & ~\pi1093  ;
  assign n64542 = ~n64540 & ~n64541 ;
  assign n64543 = ~\pi0228  & ~n64542 ;
  assign n64544 = \pi0123  & ~\pi0878  ;
  assign n64545 = ~\pi0123  & ~\pi1137  ;
  assign n64546 = \pi0228  & ~n64545 ;
  assign n64547 = ~n64544 & n64546 ;
  assign n64548 = ~n64543 & ~n64547 ;
  assign n64549 = \pi1093  & \pi1135  ;
  assign n64550 = \pi0879  & ~\pi1093  ;
  assign n64551 = ~n64549 & ~n64550 ;
  assign n64552 = ~\pi0228  & ~n64551 ;
  assign n64553 = \pi0123  & ~\pi0879  ;
  assign n64554 = ~\pi0123  & ~\pi1135  ;
  assign n64555 = \pi0228  & ~n64554 ;
  assign n64556 = ~n64553 & n64555 ;
  assign n64557 = ~n64552 & ~n64556 ;
  assign n64558 = ~\pi0955  & \pi1081  ;
  assign n64559 = \pi0880  & \pi0955  ;
  assign n64560 = ~n64558 & ~n64559 ;
  assign n64561 = ~\pi0955  & \pi1059  ;
  assign n64562 = \pi0881  & \pi0955  ;
  assign n64563 = ~n64561 & ~n64562 ;
  assign n64564 = \pi1107  & ~n64250 ;
  assign n64565 = ~\pi0883  & n64250 ;
  assign n64566 = ~n64564 & ~n64565 ;
  assign n64567 = \pi1124  & ~n64250 ;
  assign n64568 = ~\pi0884  & n64250 ;
  assign n64569 = ~n64567 & ~n64568 ;
  assign n64570 = \pi1125  & ~n64250 ;
  assign n64571 = ~\pi0885  & n64250 ;
  assign n64572 = ~n64570 & ~n64571 ;
  assign n64573 = \pi1109  & ~n64250 ;
  assign n64574 = ~\pi0886  & n64250 ;
  assign n64575 = ~n64573 & ~n64574 ;
  assign n64576 = \pi1100  & ~n64250 ;
  assign n64577 = ~\pi0887  & n64250 ;
  assign n64578 = ~n64576 & ~n64577 ;
  assign n64579 = \pi1120  & ~n64250 ;
  assign n64580 = ~\pi0888  & n64250 ;
  assign n64581 = ~n64579 & ~n64580 ;
  assign n64582 = \pi1103  & ~n64250 ;
  assign n64583 = ~\pi0889  & n64250 ;
  assign n64584 = ~n64582 & ~n64583 ;
  assign n64585 = \pi1126  & ~n64250 ;
  assign n64586 = ~\pi0890  & n64250 ;
  assign n64587 = ~n64585 & ~n64586 ;
  assign n64588 = \pi1116  & ~n64250 ;
  assign n64589 = ~\pi0891  & n64250 ;
  assign n64590 = ~n64588 & ~n64589 ;
  assign n64591 = \pi1101  & ~n64250 ;
  assign n64592 = ~\pi0892  & n64250 ;
  assign n64593 = ~n64591 & ~n64592 ;
  assign n64594 = \pi1119  & ~n64250 ;
  assign n64595 = ~\pi0894  & n64250 ;
  assign n64596 = ~n64594 & ~n64595 ;
  assign n64597 = \pi1113  & ~n64250 ;
  assign n64598 = ~\pi0895  & n64250 ;
  assign n64599 = ~n64597 & ~n64598 ;
  assign n64600 = \pi1118  & ~n64250 ;
  assign n64601 = ~\pi0896  & n64250 ;
  assign n64602 = ~n64600 & ~n64601 ;
  assign n64603 = \pi1129  & ~n64250 ;
  assign n64604 = ~\pi0898  & n64250 ;
  assign n64605 = ~n64603 & ~n64604 ;
  assign n64606 = \pi1115  & ~n64250 ;
  assign n64607 = ~\pi0899  & n64250 ;
  assign n64608 = ~n64606 & ~n64607 ;
  assign n64609 = \pi1110  & ~n64250 ;
  assign n64610 = ~\pi0900  & n64250 ;
  assign n64611 = ~n64609 & ~n64610 ;
  assign n64612 = \pi1111  & ~n64250 ;
  assign n64613 = ~\pi0902  & n64250 ;
  assign n64614 = ~n64612 & ~n64613 ;
  assign n64615 = \pi1121  & ~n64250 ;
  assign n64616 = ~\pi0903  & n64250 ;
  assign n64617 = ~n64615 & ~n64616 ;
  assign n64618 = \pi1127  & ~n64250 ;
  assign n64619 = ~\pi0904  & n64250 ;
  assign n64620 = ~n64618 & ~n64619 ;
  assign n64621 = \pi1131  & ~n64250 ;
  assign n64622 = ~\pi0905  & n64250 ;
  assign n64623 = ~n64621 & ~n64622 ;
  assign n64624 = \pi1128  & ~n64250 ;
  assign n64625 = ~\pi0906  & n64250 ;
  assign n64626 = ~n64624 & ~n64625 ;
  assign n64627 = ~\pi0604  & ~\pi0979  ;
  assign n64628 = \pi0615  & \pi0979  ;
  assign n64629 = ~n64627 & ~n64628 ;
  assign n64630 = \pi0782  & ~n64629 ;
  assign n64631 = ~\pi0782  & ~\pi0907  ;
  assign n64632 = ~\pi0598  & \pi0979  ;
  assign n64633 = ~\pi0624  & ~\pi0979  ;
  assign n64634 = \pi0782  & ~n64633 ;
  assign n64635 = ~n64632 & n64634 ;
  assign n64636 = ~n64631 & ~n64635 ;
  assign n64637 = ~n64630 & n64636 ;
  assign n64638 = \pi1122  & ~n64250 ;
  assign n64639 = ~\pi0908  & n64250 ;
  assign n64640 = ~n64638 & ~n64639 ;
  assign n64641 = \pi1105  & ~n64250 ;
  assign n64642 = ~\pi0909  & n64250 ;
  assign n64643 = ~n64641 & ~n64642 ;
  assign n64644 = \pi1117  & ~n64250 ;
  assign n64645 = ~\pi0910  & n64250 ;
  assign n64646 = ~n64644 & ~n64645 ;
  assign n64647 = \pi1130  & ~n64250 ;
  assign n64648 = ~\pi0911  & n64250 ;
  assign n64649 = ~n64647 & ~n64648 ;
  assign n64650 = \pi1114  & ~n64250 ;
  assign n64651 = ~\pi0912  & n64250 ;
  assign n64652 = ~n64650 & ~n64651 ;
  assign n64653 = \pi1106  & ~n64250 ;
  assign n64654 = ~\pi0913  & n64250 ;
  assign n64655 = ~n64653 & ~n64654 ;
  assign n64656 = \pi0280  & ~n62138 ;
  assign n64657 = ~n64234 & ~n64656 ;
  assign n64658 = \pi1108  & ~n64250 ;
  assign n64659 = ~\pi0915  & n64250 ;
  assign n64660 = ~n64658 & ~n64659 ;
  assign n64661 = \pi1123  & ~n64250 ;
  assign n64662 = ~\pi0916  & n64250 ;
  assign n64663 = ~n64661 & ~n64662 ;
  assign n64664 = \pi1112  & ~n64250 ;
  assign n64665 = ~\pi0917  & n64250 ;
  assign n64666 = ~n64664 & ~n64665 ;
  assign n64667 = \pi1104  & ~n64250 ;
  assign n64668 = ~\pi0918  & n64250 ;
  assign n64669 = ~n64667 & ~n64668 ;
  assign n64670 = \pi1102  & ~n64250 ;
  assign n64671 = ~\pi0919  & n64250 ;
  assign n64672 = ~n64670 & ~n64671 ;
  assign n64673 = \pi1093  & \pi1139  ;
  assign n64674 = \pi0920  & ~\pi1093  ;
  assign n64675 = ~n64673 & ~n64674 ;
  assign n64676 = \pi0921  & ~\pi1093  ;
  assign n64677 = ~n64495 & ~n64676 ;
  assign n64678 = ~\pi0922  & ~\pi1093  ;
  assign n64679 = \pi1093  & ~\pi1152  ;
  assign n64680 = ~n64678 & ~n64679 ;
  assign n64681 = ~\pi0923  & ~\pi1093  ;
  assign n64682 = \pi1093  & ~\pi1154  ;
  assign n64683 = ~n64681 & ~n64682 ;
  assign n64684 = \pi0301  & \pi0311  ;
  assign n64685 = n58610 & n64684 ;
  assign n64686 = ~\pi0925  & ~\pi1093  ;
  assign n64687 = \pi1093  & ~\pi1155  ;
  assign n64688 = ~n64686 & ~n64687 ;
  assign n64689 = ~\pi0926  & ~\pi1093  ;
  assign n64690 = \pi1093  & ~\pi1157  ;
  assign n64691 = ~n64689 & ~n64690 ;
  assign n64692 = ~\pi0927  & ~\pi1093  ;
  assign n64693 = \pi1093  & ~\pi1145  ;
  assign n64694 = ~n64692 & ~n64693 ;
  assign n64695 = ~\pi0928  & ~\pi1093  ;
  assign n64696 = ~n64519 & ~n64695 ;
  assign n64697 = ~\pi0929  & ~\pi1093  ;
  assign n64698 = \pi1093  & ~\pi1144  ;
  assign n64699 = ~n64697 & ~n64698 ;
  assign n64700 = ~\pi0930  & ~\pi1093  ;
  assign n64701 = \pi1093  & ~\pi1134  ;
  assign n64702 = ~n64700 & ~n64701 ;
  assign n64703 = ~\pi0931  & ~\pi1093  ;
  assign n64704 = \pi1093  & ~\pi1150  ;
  assign n64705 = ~n64703 & ~n64704 ;
  assign n64706 = \pi0932  & ~\pi1093  ;
  assign n64707 = ~n56381 & ~n64706 ;
  assign n64708 = \pi0933  & ~\pi1093  ;
  assign n64709 = ~n64540 & ~n64708 ;
  assign n64710 = ~\pi0934  & ~\pi1093  ;
  assign n64711 = \pi1093  & ~\pi1147  ;
  assign n64712 = ~n64710 & ~n64711 ;
  assign n64713 = \pi0935  & ~\pi1093  ;
  assign n64714 = ~n64465 & ~n64713 ;
  assign n64715 = ~\pi0936  & ~\pi1093  ;
  assign n64716 = \pi1093  & ~\pi1149  ;
  assign n64717 = ~n64715 & ~n64716 ;
  assign n64718 = ~\pi0937  & ~\pi1093  ;
  assign n64719 = \pi1093  & ~\pi1148  ;
  assign n64720 = ~n64718 & ~n64719 ;
  assign n64721 = \pi0938  & ~\pi1093  ;
  assign n64722 = ~n64549 & ~n64721 ;
  assign n64723 = ~\pi0939  & ~\pi1093  ;
  assign n64724 = \pi1093  & ~\pi1146  ;
  assign n64725 = ~n64723 & ~n64724 ;
  assign n64726 = \pi0940  & ~\pi1093  ;
  assign n64727 = ~n64531 & ~n64726 ;
  assign n64728 = ~\pi0941  & ~\pi1093  ;
  assign n64729 = \pi1093  & ~\pi1153  ;
  assign n64730 = ~n64728 & ~n64729 ;
  assign n64731 = ~\pi0942  & ~\pi1093  ;
  assign n64732 = \pi1093  & ~\pi1156  ;
  assign n64733 = ~n64731 & ~n64732 ;
  assign n64734 = ~\pi0943  & ~\pi1093  ;
  assign n64735 = \pi1093  & ~\pi1151  ;
  assign n64736 = ~n64734 & ~n64735 ;
  assign n64737 = \pi1093  & \pi1143  ;
  assign n64738 = \pi0944  & ~\pi1093  ;
  assign n64739 = ~n64737 & ~n64738 ;
  assign n64740 = \pi0230  & n1689 ;
  assign n64741 = ~\pi0782  & \pi0947  ;
  assign n64742 = ~n64635 & ~n64741 ;
  assign n64743 = ~\pi0266  & ~\pi0992  ;
  assign n64744 = ~n62138 & ~n64743 ;
  assign n64745 = ~\pi0313  & ~\pi0954  ;
  assign n64746 = \pi0949  & \pi0954  ;
  assign n64747 = ~n64745 & ~n64746 ;
  assign n64748 = n1686 & n1695 ;
  assign n64749 = ~n8543 & n8739 ;
  assign n64750 = \pi0957  & \pi1092  ;
  assign n64751 = ~\pi0031  & ~n64750 ;
  assign n64752 = ~\pi0782  & \pi0960  ;
  assign n64753 = ~\pi0230  & \pi0961  ;
  assign n64754 = ~\pi0782  & \pi0963  ;
  assign n64755 = ~\pi0230  & \pi0967  ;
  assign n64756 = ~\pi0230  & \pi0969  ;
  assign n64757 = ~\pi0782  & \pi0970  ;
  assign n64758 = ~\pi0230  & \pi0971  ;
  assign n64759 = ~\pi0782  & \pi0972  ;
  assign n64760 = ~\pi0230  & \pi0974  ;
  assign n64761 = ~\pi0782  & \pi0975  ;
  assign n64762 = ~\pi0230  & \pi0977  ;
  assign n64763 = ~\pi0782  & \pi0978  ;
  assign n64764 = ~\pi0598  & \pi0615  ;
  assign n64765 = \pi0824  & \pi1092  ;
  assign n64766 = ~\pi0604  & ~\pi0624  ;
  assign \po0000  = \pi0668  ;
  assign \po0001  = \pi0672  ;
  assign \po0002  = \pi0664  ;
  assign \po0003  = \pi0667  ;
  assign \po0004  = \pi0676  ;
  assign \po0005  = \pi0673  ;
  assign \po0006  = \pi0675  ;
  assign \po0007  = \pi0666  ;
  assign \po0008  = \pi0679  ;
  assign \po0009  = \pi0674  ;
  assign \po0010  = \pi0663  ;
  assign \po0011  = \pi0670  ;
  assign \po0012  = \pi0677  ;
  assign \po0013  = \pi0682  ;
  assign \po0014  = \pi0671  ;
  assign \po0015  = \pi0678  ;
  assign \po0016  = \pi0718  ;
  assign \po0017  = \pi0707  ;
  assign \po0018  = \pi0708  ;
  assign \po0019  = \pi0713  ;
  assign \po0020  = \pi0711  ;
  assign \po0021  = \pi0716  ;
  assign \po0022  = \pi0733  ;
  assign \po0023  = \pi0712  ;
  assign \po0024  = \pi0689  ;
  assign \po0025  = \pi0717  ;
  assign \po0026  = \pi0692  ;
  assign \po0027  = \pi0719  ;
  assign \po0028  = \pi0722  ;
  assign \po0029  = \pi0714  ;
  assign \po0030  = \pi0720  ;
  assign \po0031  = \pi0685  ;
  assign \po0032  = \pi0837  ;
  assign \po0033  = \pi0850  ;
  assign \po0034  = \pi0872  ;
  assign \po0035  = \pi0871  ;
  assign \po0036  = \pi0881  ;
  assign \po0037  = \pi0866  ;
  assign \po0038  = \pi0876  ;
  assign \po0039  = \pi0873  ;
  assign \po0040  = \pi0874  ;
  assign \po0041  = \pi0859  ;
  assign \po0042  = \pi0855  ;
  assign \po0043  = \pi0852  ;
  assign \po0044  = \pi0870  ;
  assign \po0045  = \pi0848  ;
  assign \po0046  = \pi0865  ;
  assign \po0047  = \pi0856  ;
  assign \po0048  = \pi0853  ;
  assign \po0049  = \pi0847  ;
  assign \po0050  = \pi0857  ;
  assign \po0051  = \pi0854  ;
  assign \po0052  = \pi0858  ;
  assign \po0053  = \pi0845  ;
  assign \po0054  = \pi0838  ;
  assign \po0055  = \pi0842  ;
  assign \po0056  = \pi0843  ;
  assign \po0057  = \pi0839  ;
  assign \po0058  = \pi0844  ;
  assign \po0059  = \pi0868  ;
  assign \po0060  = \pi0851  ;
  assign \po0061  = \pi0867  ;
  assign \po0062  = \pi0880  ;
  assign \po0063  = \pi0860  ;
  assign \po0064  = \pi1030  ;
  assign \po0065  = \pi1034  ;
  assign \po0066  = \pi1015  ;
  assign \po0067  = \pi1020  ;
  assign \po0068  = \pi1025  ;
  assign \po0069  = \pi1005  ;
  assign \po0070  = \pi0996  ;
  assign \po0071  = \pi1012  ;
  assign \po0072  = \pi0993  ;
  assign \po0073  = \pi1016  ;
  assign \po0074  = \pi1021  ;
  assign \po0075  = \pi1010  ;
  assign \po0076  = \pi1027  ;
  assign \po0077  = \pi1018  ;
  assign \po0078  = \pi1017  ;
  assign \po0079  = \pi1024  ;
  assign \po0080  = \pi1009  ;
  assign \po0081  = \pi1032  ;
  assign \po0082  = \pi1003  ;
  assign \po0083  = \pi0997  ;
  assign \po0084  = \pi1013  ;
  assign \po0085  = \pi1011  ;
  assign \po0086  = \pi1008  ;
  assign \po0087  = \pi1019  ;
  assign \po0088  = \pi1031  ;
  assign \po0089  = \pi1022  ;
  assign \po0090  = \pi1000  ;
  assign \po0091  = \pi1023  ;
  assign \po0092  = \pi1002  ;
  assign \po0093  = \pi1026  ;
  assign \po0094  = \pi1006  ;
  assign \po0095  = \pi0998  ;
  assign \po0096  = \pi0031  ;
  assign \po0097  = \pi0080  ;
  assign \po0098  = \pi0893  ;
  assign \po0099  = \pi0467  ;
  assign \po0100  = \pi0078  ;
  assign \po0101  = \pi0112  ;
  assign \po0102  = \pi0013  ;
  assign \po0103  = \pi0025  ;
  assign \po0104  = \pi0226  ;
  assign \po0105  = \pi0127  ;
  assign \po0106  = \pi0822  ;
  assign \po0107  = \pi0808  ;
  assign \po0108  = \pi0227  ;
  assign \po0109  = \pi0477  ;
  assign \po0110  = \pi0834  ;
  assign \po0111  = \pi0229  ;
  assign \po0112  = \pi0012  ;
  assign \po0113  = \pi0011  ;
  assign \po0114  = \pi0010  ;
  assign \po0115  = \pi0009  ;
  assign \po0116  = \pi0008  ;
  assign \po0117  = \pi0007  ;
  assign \po0118  = \pi0006  ;
  assign \po0119  = \pi0005  ;
  assign \po0120  = \pi0004  ;
  assign \po0121  = \pi0003  ;
  assign \po0122  = \pi0000  ;
  assign \po0123  = \pi0002  ;
  assign \po0124  = \pi0001  ;
  assign \po0125  = \pi0310  ;
  assign \po0126  = \pi0302  ;
  assign \po0127  = \pi0475  ;
  assign \po0128  = \pi0474  ;
  assign \po0129  = \pi0466  ;
  assign \po0130  = \pi0473  ;
  assign \po0131  = \pi0471  ;
  assign \po0132  = \pi0472  ;
  assign \po0133  = \pi0470  ;
  assign \po0134  = \pi0469  ;
  assign \po0135  = \pi0465  ;
  assign \po0136  = \pi1028  ;
  assign \po0137  = \pi1033  ;
  assign \po0138  = \pi0995  ;
  assign \po0139  = \pi0994  ;
  assign \po0140  = \pi0028  ;
  assign \po0141  = \pi0027  ;
  assign \po0142  = \pi0026  ;
  assign \po0143  = \pi0029  ;
  assign \po0144  = \pi0015  ;
  assign \po0145  = \pi0014  ;
  assign \po0146  = \pi0021  ;
  assign \po0147  = \pi0020  ;
  assign \po0148  = \pi0019  ;
  assign \po0149  = \pi0018  ;
  assign \po0150  = \pi0017  ;
  assign \po0151  = \pi0016  ;
  assign \po0152  = \pi1096  ;
  assign \po0153  = n2466 ;
  assign \po0154  = ~n2784 ;
  assign \po0155  = n3042 ;
  assign \po0156  = n3387 ;
  assign \po0157  = ~n3732 ;
  assign \po0158  = n4067 ;
  assign \po0159  = n4397 ;
  assign \po0160  = ~n4735 ;
  assign \po0161  = n5064 ;
  assign \po0162  = n5398 ;
  assign \po0163  = n5747 ;
  assign \po0164  = n6084 ;
  assign \po0165  = ~n6620 ;
  assign \po0166  = ~1'b0 ;
  assign \po0167  = n6846 ;
  assign \po0168  = \pi0228  ;
  assign \po0169  = \pi0022  ;
  assign \po0170  = ~\pi1090  ;
  assign \po0171  = ~n7279 ;
  assign \po0172  = n7485 ;
  assign \po0173  = n7677 ;
  assign \po0174  = n7812 ;
  assign \po0175  = n7943 ;
  assign \po0176  = n8074 ;
  assign \po0177  = n8205 ;
  assign \po0178  = n8346 ;
  assign \po0179  = \pi1089  ;
  assign \po0180  = \pi0023  ;
  assign \po0181  = n6846 ;
  assign \po0182  = n8452 ;
  assign \po0183  = ~n8528 ;
  assign \po0184  = ~n8533 ;
  assign \po0185  = ~n8536 ;
  assign \po0186  = ~n8539 ;
  assign \po0187  = ~n8542 ;
  assign \po0188  = \pi0037  ;
  assign \po0189  = ~n10014 ;
  assign \po0190  = n10102 ;
  assign \po0191  = n11116 ;
  assign \po0192  = n11686 ;
  assign \po0193  = n11802 ;
  assign \po0194  = n11826 ;
  assign \po0195  = ~n11827 ;
  assign \po0196  = n11857 ;
  assign \po0197  = n11964 ;
  assign \po0198  = n11983 ;
  assign \po0199  = ~n12254 ;
  assign \po0200  = ~n12575 ;
  assign \po0201  = ~n12824 ;
  assign \po0202  = ~n12964 ;
  assign \po0203  = n12973 ;
  assign \po0204  = n12999 ;
  assign \po0205  = n13077 ;
  assign \po0206  = n13081 ;
  assign \po0207  = n13106 ;
  assign \po0208  = n13148 ;
  assign \po0209  = n13156 ;
  assign \po0210  = n13385 ;
  assign \po0211  = n13401 ;
  assign \po0212  = n13425 ;
  assign \po0213  = ~n13446 ;
  assign \po0214  = n13461 ;
  assign \po0215  = ~n13472 ;
  assign \po0216  = n13477 ;
  assign \po0217  = ~n13485 ;
  assign \po0218  = n13495 ;
  assign \po0219  = n13505 ;
  assign \po0220  = ~n13512 ;
  assign \po0221  = n13521 ;
  assign \po0222  = n13533 ;
  assign \po0223  = ~n13542 ;
  assign \po0224  = n13565 ;
  assign \po0225  = n13576 ;
  assign \po0226  = n13586 ;
  assign \po0227  = ~n13610 ;
  assign \po0228  = ~n13641 ;
  assign \po0229  = n13680 ;
  assign \po0230  = n13700 ;
  assign \po0231  = n13715 ;
  assign \po0232  = ~n13734 ;
  assign \po0233  = n13747 ;
  assign \po0234  = n14000 ;
  assign \po0235  = n14016 ;
  assign \po0236  = n14018 ;
  assign \po0237  = ~n14693 ;
  assign \po0238  = n15308 ;
  assign \po0239  = n15317 ;
  assign \po0240  = n15331 ;
  assign \po0241  = n15350 ;
  assign \po0242  = n15357 ;
  assign \po0243  = ~n15373 ;
  assign \po0244  = n15383 ;
  assign \po0245  = n15386 ;
  assign \po0246  = n15421 ;
  assign \po0247  = n15434 ;
  assign \po0248  = n15447 ;
  assign \po0249  = n15465 ;
  assign \po0250  = ~n15479 ;
  assign \po0251  = n15493 ;
  assign \po0252  = n15521 ;
  assign \po0253  = n15542 ;
  assign \po0254  = ~n15561 ;
  assign \po0255  = n15576 ;
  assign \po0256  = n15588 ;
  assign \po0257  = ~n15709 ;
  assign \po0258  = n15727 ;
  assign \po0259  = n15840 ;
  assign \po0260  = n15846 ;
  assign \po0261  = n15857 ;
  assign \po0262  = ~n15881 ;
  assign \po0263  = \pi0117  ;
  assign \po0264  = n15905 ;
  assign \po0265  = n15909 ;
  assign \po0266  = n15938 ;
  assign \po0267  = n15944 ;
  assign \po0268  = ~n15959 ;
  assign \po0269  = n15973 ;
  assign \po0270  = ~n15974 ;
  assign \po0271  = n16050 ;
  assign \po0272  = n16123 ;
  assign \po0273  = n16184 ;
  assign \po0274  = n16283 ;
  assign \po0275  = n16310 ;
  assign \po0276  = ~n16771 ;
  assign \po0277  = ~n16853 ;
  assign \po0278  = ~n17415 ;
  assign \po0279  = ~n18046 ;
  assign \po0280  = n18058 ;
  assign \po0281  = ~n18148 ;
  assign \po0282  = ~n18754 ;
  assign \po0283  = ~n19260 ;
  assign \po0284  = n19378 ;
  assign \po0285  = \pi0131  ;
  assign \po0286  = n19412 ;
  assign \po0287  = n19608 ;
  assign \po0288  = n19618 ;
  assign \po0289  = ~n19975 ;
  assign \po0290  = ~n20043 ;
  assign \po0291  = n20190 ;
  assign \po0292  = n20373 ;
  assign \po0293  = n20505 ;
  assign \po0294  = ~n20527 ;
  assign \po0295  = n20675 ;
  assign \po0296  = n20775 ;
  assign \po0297  = n23081 ;
  assign \po0298  = n23775 ;
  assign \po0299  = ~n24821 ;
  assign \po0300  = n25537 ;
  assign \po0301  = ~n26298 ;
  assign \po0302  = ~n26929 ;
  assign \po0303  = ~n27050 ;
  assign \po0304  = n27318 ;
  assign \po0305  = ~n27419 ;
  assign \po0306  = ~n27506 ;
  assign \po0307  = n27588 ;
  assign \po0308  = n27703 ;
  assign \po0309  = n27861 ;
  assign \po0310  = ~n27968 ;
  assign \po0311  = n28047 ;
  assign \po0312  = ~n28123 ;
  assign \po0313  = n28169 ;
  assign \po0314  = n28254 ;
  assign \po0315  = n28334 ;
  assign \po0316  = n28414 ;
  assign \po0317  = ~n28502 ;
  assign \po0318  = n28640 ;
  assign \po0319  = ~n28726 ;
  assign \po0320  = ~n28813 ;
  assign \po0321  = n28873 ;
  assign \po0322  = n28933 ;
  assign \po0323  = n29083 ;
  assign \po0324  = n29146 ;
  assign \po0325  = ~n29247 ;
  assign \po0326  = ~n29348 ;
  assign \po0327  = n29449 ;
  assign \po0328  = ~n29550 ;
  assign \po0329  = ~n29661 ;
  assign \po0330  = ~n30251 ;
  assign \po0331  = n30829 ;
  assign \po0332  = n31421 ;
  assign \po0333  = ~n31957 ;
  assign \po0334  = n32535 ;
  assign \po0335  = n33107 ;
  assign \po0336  = ~n33715 ;
  assign \po0337  = n34286 ;
  assign \po0338  = ~n34864 ;
  assign \po0339  = ~n35442 ;
  assign \po0340  = ~n36019 ;
  assign \po0341  = ~n36593 ;
  assign \po0342  = n37162 ;
  assign \po0343  = ~n37729 ;
  assign \po0344  = ~n38328 ;
  assign \po0345  = ~n38926 ;
  assign \po0346  = n39524 ;
  assign \po0347  = n40098 ;
  assign \po0348  = n40663 ;
  assign \po0349  = n41228 ;
  assign \po0350  = n41807 ;
  assign \po0351  = ~n42353 ;
  assign \po0352  = ~n42437 ;
  assign \po0353  = ~n42551 ;
  assign \po0354  = n42651 ;
  assign \po0355  = n43627 ;
  assign \po0356  = ~n43962 ;
  assign \po0357  = ~n44301 ;
  assign \po0358  = n44555 ;
  assign \po0359  = n44572 ;
  assign \po0360  = n44588 ;
  assign \po0361  = ~n44763 ;
  assign \po0362  = ~n44781 ;
  assign \po0363  = ~n44796 ;
  assign \po0364  = n45533 ;
  assign \po0365  = n45631 ;
  assign \po0366  = ~n45855 ;
  assign \po0367  = ~n46112 ;
  assign \po0368  = ~n46156 ;
  assign \po0369  = ~n46198 ;
  assign \po0370  = n46239 ;
  assign \po0371  = ~n46281 ;
  assign \po0372  = ~n46484 ;
  assign \po0373  = ~n46681 ;
  assign \po0374  = ~n46722 ;
  assign \po0375  = ~n46738 ;
  assign \po0376  = ~n46784 ;
  assign \po0377  = n46796 ;
  assign \po0378  = n46999 ;
  assign \po0379  = ~n47995 ;
  assign \po0380  = n48878 ;
  assign \po0381  = n49764 ;
  assign \po0382  = ~n49981 ;
  assign \po0383  = n50064 ;
  assign \po0384  = ~n50117 ;
  assign \po0385  = ~n50137 ;
  assign \po0386  = \pi0232  ;
  assign \po0387  = ~n50270 ;
  assign \po0388  = \pi0236  ;
  assign \po0389  = n50361 ;
  assign \po0390  = ~n50821 ;
  assign \po0391  = n51258 ;
  assign \po0392  = n51540 ;
  assign \po0393  = n51563 ;
  assign \po0394  = n51911 ;
  assign \po0395  = ~n52380 ;
  assign \po0396  = n52511 ;
  assign \po0397  = n53032 ;
  assign \po0398  = n53426 ;
  assign \po0399  = ~n53532 ;
  assign \po0400  = n53964 ;
  assign \po0401  = ~n54055 ;
  assign \po0402  = ~n54388 ;
  assign \po0403  = ~n54767 ;
  assign \po0404  = n55093 ;
  assign \po0405  = n55331 ;
  assign \po0406  = n55591 ;
  assign \po0407  = ~n55606 ;
  assign \po0408  = ~n55617 ;
  assign \po0409  = ~n55688 ;
  assign \po0410  = ~n56002 ;
  assign \po0411  = n56328 ;
  assign \po0412  = n56334 ;
  assign \po0413  = n56340 ;
  assign \po0414  = n56346 ;
  assign \po0415  = n56352 ;
  assign \po0416  = n56358 ;
  assign \po0417  = ~n56365 ;
  assign \po0418  = ~n56372 ;
  assign \po0419  = ~n56402 ;
  assign \po0420  = n56675 ;
  assign \po0421  = ~n56740 ;
  assign \po0422  = ~n56796 ;
  assign \po0423  = n56889 ;
  assign \po0424  = n57161 ;
  assign \po0425  = n57397 ;
  assign \po0426  = n57446 ;
  assign \po0427  = n57492 ;
  assign \po0428  = n57558 ;
  assign \po0429  = n57711 ;
  assign \po0430  = ~n57803 ;
  assign \po0431  = n57859 ;
  assign \po0432  = ~n57964 ;
  assign \po0433  = ~n58000 ;
  assign \po0434  = ~n58059 ;
  assign \po0435  = ~n58150 ;
  assign \po0436  = n58222 ;
  assign \po0437  = n58272 ;
  assign \po0438  = n58316 ;
  assign \po0439  = n58359 ;
  assign \po0440  = n58465 ;
  assign \po0441  = ~n58469 ;
  assign \po0442  = n58494 ;
  assign \po0443  = n58529 ;
  assign \po0444  = n58531 ;
  assign \po0445  = n58543 ;
  assign \po0446  = n58560 ;
  assign \po0447  = n58563 ;
  assign \po0448  = n58566 ;
  assign \po0449  = n58569 ;
  assign \po0450  = n58572 ;
  assign \po0451  = n58575 ;
  assign \po0452  = n58578 ;
  assign \po0453  = n58581 ;
  assign \po0454  = n58584 ;
  assign \po0455  = ~n58587 ;
  assign \po0456  = n58604 ;
  assign \po0457  = ~n58616 ;
  assign \po0458  = ~n58622 ;
  assign \po0459  = n58647 ;
  assign \po0460  = ~n58650 ;
  assign \po0461  = ~n58653 ;
  assign \po0462  = ~n58656 ;
  assign \po0463  = ~n58659 ;
  assign \po0464  = ~n58662 ;
  assign \po0465  = ~n58665 ;
  assign \po0466  = ~n58668 ;
  assign \po0467  = ~n58700 ;
  assign \po0468  = n58705 ;
  assign \po0469  = ~n58713 ;
  assign \po0470  = ~n58726 ;
  assign \po0471  = ~n58745 ;
  assign \po0472  = ~n58752 ;
  assign \po0473  = ~n58757 ;
  assign \po0474  = ~n58764 ;
  assign \po0475  = ~n58771 ;
  assign \po0476  = ~n58776 ;
  assign \po0477  = ~n58781 ;
  assign \po0478  = ~n58786 ;
  assign \po0479  = ~n58791 ;
  assign \po0480  = ~n58796 ;
  assign \po0481  = ~n58801 ;
  assign \po0482  = ~n58806 ;
  assign \po0483  = ~n58811 ;
  assign \po0484  = ~n58816 ;
  assign \po0485  = ~n58821 ;
  assign \po0486  = ~n58826 ;
  assign \po0487  = n58833 ;
  assign \po0488  = n58839 ;
  assign \po0489  = ~n58861 ;
  assign \po0490  = ~n58866 ;
  assign \po0491  = ~n58871 ;
  assign \po0492  = ~n58876 ;
  assign \po0493  = ~n58881 ;
  assign \po0494  = ~n58886 ;
  assign \po0495  = ~n58891 ;
  assign \po0496  = ~n58896 ;
  assign \po0497  = ~n58906 ;
  assign \po0498  = n58912 ;
  assign \po0499  = ~n58917 ;
  assign \po0500  = ~n58922 ;
  assign \po0501  = ~n58927 ;
  assign \po0502  = ~n58932 ;
  assign \po0503  = ~n58937 ;
  assign \po0504  = ~n58942 ;
  assign \po0505  = ~n58947 ;
  assign \po0506  = ~n58952 ;
  assign \po0507  = ~n58957 ;
  assign \po0508  = ~n58962 ;
  assign \po0509  = ~n58967 ;
  assign \po0510  = ~n58972 ;
  assign \po0511  = ~n58977 ;
  assign \po0512  = ~n58982 ;
  assign \po0513  = ~n58987 ;
  assign \po0514  = ~n58992 ;
  assign \po0515  = ~n58997 ;
  assign \po0516  = ~n59002 ;
  assign \po0517  = ~n59007 ;
  assign \po0518  = ~n59012 ;
  assign \po0519  = ~n59017 ;
  assign \po0520  = ~n59022 ;
  assign \po0521  = ~n59027 ;
  assign \po0522  = ~n59032 ;
  assign \po0523  = ~n59037 ;
  assign \po0524  = ~n59042 ;
  assign \po0525  = ~n59047 ;
  assign \po0526  = ~n59052 ;
  assign \po0527  = ~n59057 ;
  assign \po0528  = ~n59062 ;
  assign \po0529  = ~n59067 ;
  assign \po0530  = ~n59072 ;
  assign \po0531  = ~n59077 ;
  assign \po0532  = ~n59082 ;
  assign \po0533  = ~n59087 ;
  assign \po0534  = ~n59092 ;
  assign \po0535  = ~n59097 ;
  assign \po0536  = ~n59102 ;
  assign \po0537  = ~n59107 ;
  assign \po0538  = ~n59112 ;
  assign \po0539  = ~n59117 ;
  assign \po0540  = ~n59122 ;
  assign \po0541  = ~n59127 ;
  assign \po0542  = ~n59132 ;
  assign \po0543  = ~n59137 ;
  assign \po0544  = ~n59142 ;
  assign \po0545  = ~n59147 ;
  assign \po0546  = ~n59152 ;
  assign \po0547  = ~n59157 ;
  assign \po0548  = ~n59162 ;
  assign \po0549  = ~n59167 ;
  assign \po0550  = ~n59172 ;
  assign \po0551  = ~n59177 ;
  assign \po0552  = ~n59182 ;
  assign \po0553  = ~n59187 ;
  assign \po0554  = ~n59192 ;
  assign \po0555  = ~n59197 ;
  assign \po0556  = ~n59202 ;
  assign \po0557  = ~n59207 ;
  assign \po0558  = ~n59212 ;
  assign \po0559  = ~n59217 ;
  assign \po0560  = ~n59222 ;
  assign \po0561  = ~n59227 ;
  assign \po0562  = ~n59232 ;
  assign \po0563  = ~n59237 ;
  assign \po0564  = ~n59242 ;
  assign \po0565  = ~n59247 ;
  assign \po0566  = ~n59252 ;
  assign \po0567  = ~n59257 ;
  assign \po0568  = ~n59262 ;
  assign \po0569  = ~n59267 ;
  assign \po0570  = ~n59272 ;
  assign \po0571  = ~n59277 ;
  assign \po0572  = ~n59282 ;
  assign \po0573  = ~n59287 ;
  assign \po0574  = ~n59292 ;
  assign \po0575  = ~n59297 ;
  assign \po0576  = ~n59302 ;
  assign \po0577  = ~n59307 ;
  assign \po0578  = ~n59312 ;
  assign \po0579  = ~n59317 ;
  assign \po0580  = ~n59322 ;
  assign \po0581  = ~n59327 ;
  assign \po0582  = ~n59332 ;
  assign \po0583  = ~n59337 ;
  assign \po0584  = ~n59342 ;
  assign \po0585  = ~n59347 ;
  assign \po0586  = ~n59352 ;
  assign \po0587  = ~n59357 ;
  assign \po0588  = ~n59362 ;
  assign \po0589  = ~n59367 ;
  assign \po0590  = ~n59372 ;
  assign \po0591  = ~n59377 ;
  assign \po0592  = ~n59382 ;
  assign \po0593  = ~n59387 ;
  assign \po0594  = ~n59392 ;
  assign \po0595  = ~n59397 ;
  assign \po0596  = ~n59402 ;
  assign \po0597  = ~n59407 ;
  assign \po0598  = ~n59412 ;
  assign \po0599  = ~n59417 ;
  assign \po0600  = ~n59422 ;
  assign \po0601  = ~n59427 ;
  assign \po0602  = ~n59432 ;
  assign \po0603  = ~n59437 ;
  assign \po0604  = ~n59442 ;
  assign \po0605  = ~n59447 ;
  assign \po0606  = ~n59452 ;
  assign \po0607  = ~n59457 ;
  assign \po0608  = ~n59462 ;
  assign \po0609  = ~n59467 ;
  assign \po0610  = ~n59472 ;
  assign \po0611  = ~n59477 ;
  assign \po0612  = ~n59482 ;
  assign \po0613  = ~n59487 ;
  assign \po0614  = n59514 ;
  assign \po0615  = ~n59519 ;
  assign \po0616  = ~n59524 ;
  assign \po0617  = ~n59529 ;
  assign \po0618  = ~n59534 ;
  assign \po0619  = ~n59539 ;
  assign \po0620  = ~n59544 ;
  assign \po0621  = ~n59549 ;
  assign \po0622  = ~n59584 ;
  assign \po0623  = n59608 ;
  assign \po0624  = ~n59649 ;
  assign \po0625  = ~n59660 ;
  assign \po0626  = ~n59684 ;
  assign \po0627  = ~n59708 ;
  assign \po0628  = ~n59732 ;
  assign \po0629  = ~n59756 ;
  assign \po0630  = n59773 ;
  assign \po0631  = n59790 ;
  assign \po0632  = n59807 ;
  assign \po0633  = n59825 ;
  assign \po0634  = ~n59827 ;
  assign \po0635  = n59828 ;
  assign \po0636  = \pi0583  ;
  assign \po0637  = n59829 ;
  assign \po0638  = ~n59834 ;
  assign \po0639  = ~n59839 ;
  assign \po0640  = ~n59844 ;
  assign \po0641  = ~n59849 ;
  assign \po0642  = ~n59853 ;
  assign \po0643  = ~n59857 ;
  assign \po0644  = ~n59862 ;
  assign \po0645  = n59867 ;
  assign \po0646  = ~n59871 ;
  assign \po0647  = ~n59875 ;
  assign \po0648  = ~n59879 ;
  assign \po0649  = ~n59883 ;
  assign \po0650  = ~n59887 ;
  assign \po0651  = n59891 ;
  assign \po0652  = ~n59895 ;
  assign \po0653  = ~n59899 ;
  assign \po0654  = n59903 ;
  assign \po0655  = ~n59908 ;
  assign \po0656  = ~n59912 ;
  assign \po0657  = ~n59916 ;
  assign \po0658  = ~n59920 ;
  assign \po0659  = ~n59924 ;
  assign \po0660  = ~n59928 ;
  assign \po0661  = ~n59932 ;
  assign \po0662  = ~n59939 ;
  assign \po0663  = ~n59943 ;
  assign \po0664  = ~n59947 ;
  assign \po0665  = ~n59951 ;
  assign \po0666  = ~n59955 ;
  assign \po0667  = ~n59959 ;
  assign \po0668  = ~n59964 ;
  assign \po0669  = ~n59969 ;
  assign \po0670  = ~n59974 ;
  assign \po0671  = ~n59978 ;
  assign \po0672  = ~n59983 ;
  assign \po0673  = ~n59987 ;
  assign \po0674  = ~n59991 ;
  assign \po0675  = ~n59995 ;
  assign \po0676  = n59999 ;
  assign \po0677  = ~n60003 ;
  assign \po0678  = ~n60007 ;
  assign \po0679  = ~n60012 ;
  assign \po0680  = ~n60017 ;
  assign \po0681  = n60021 ;
  assign \po0682  = ~n60026 ;
  assign \po0683  = ~n60031 ;
  assign \po0684  = ~n60036 ;
  assign \po0685  = ~n60040 ;
  assign \po0686  = ~n60044 ;
  assign \po0687  = ~n60048 ;
  assign \po0688  = ~n60053 ;
  assign \po0689  = ~n60058 ;
  assign \po0690  = ~n60061 ;
  assign \po0691  = n60064 ;
  assign \po0692  = ~n60067 ;
  assign \po0693  = ~n60070 ;
  assign \po0694  = ~n60073 ;
  assign \po0695  = ~n60077 ;
  assign \po0696  = ~n60081 ;
  assign \po0697  = ~n60085 ;
  assign \po0698  = ~n60089 ;
  assign \po0699  = ~n60093 ;
  assign \po0700  = ~n60096 ;
  assign \po0701  = ~n60101 ;
  assign \po0702  = ~n60104 ;
  assign \po0703  = ~n60107 ;
  assign \po0704  = ~n60110 ;
  assign \po0705  = ~n60114 ;
  assign \po0706  = ~n60117 ;
  assign \po0707  = n60121 ;
  assign \po0708  = ~n60125 ;
  assign \po0709  = ~n60128 ;
  assign \po0710  = ~n60132 ;
  assign \po0711  = ~n60136 ;
  assign \po0712  = ~n60139 ;
  assign \po0713  = ~n60143 ;
  assign \po0714  = ~n60147 ;
  assign \po0715  = ~n60150 ;
  assign \po0716  = ~n60154 ;
  assign \po0717  = ~n60158 ;
  assign \po0718  = ~n60162 ;
  assign \po0719  = ~n60166 ;
  assign \po0720  = ~n60170 ;
  assign \po0721  = ~n60174 ;
  assign \po0722  = ~n60178 ;
  assign \po0723  = ~n60182 ;
  assign \po0724  = n60259 ;
  assign \po0725  = ~n60264 ;
  assign \po0726  = n60268 ;
  assign \po0727  = ~n60272 ;
  assign \po0728  = ~n60276 ;
  assign \po0729  = ~n60280 ;
  assign \po0730  = ~n60284 ;
  assign \po0731  = ~n60288 ;
  assign \po0732  = ~n60292 ;
  assign \po0733  = ~n60296 ;
  assign \po0734  = ~n60299 ;
  assign \po0735  = ~n60303 ;
  assign \po0736  = ~n60307 ;
  assign \po0737  = ~n60310 ;
  assign \po0738  = ~n60314 ;
  assign \po0739  = ~n60318 ;
  assign \po0740  = n8604 ;
  assign \po0741  = ~n60322 ;
  assign \po0742  = ~n60326 ;
  assign \po0743  = ~n60330 ;
  assign \po0744  = ~n60336 ;
  assign \po0745  = n60342 ;
  assign \po0746  = n60399 ;
  assign \po0747  = ~n60404 ;
  assign \po0748  = n60409 ;
  assign \po0749  = n60414 ;
  assign \po0750  = n61722 ;
  assign \po0751  = n61729 ;
  assign \po0752  = n61737 ;
  assign \po0753  = n61748 ;
  assign \po0754  = ~n61753 ;
  assign \po0755  = ~n61760 ;
  assign \po0756  = n61764 ;
  assign \po0757  = n61766 ;
  assign \po0758  = n61770 ;
  assign \po0759  = ~n61778 ;
  assign \po0760  = ~n61793 ;
  assign \po0761  = ~n61801 ;
  assign \po0762  = n61804 ;
  assign \po0763  = n61813 ;
  assign \po0764  = n61819 ;
  assign \po0765  = n61825 ;
  assign \po0766  = n61831 ;
  assign \po0767  = n61837 ;
  assign \po0768  = n61843 ;
  assign \po0769  = n61849 ;
  assign \po0770  = n61855 ;
  assign \po0771  = ~n61862 ;
  assign \po0772  = ~n61869 ;
  assign \po0773  = ~n61876 ;
  assign \po0774  = n61885 ;
  assign \po0775  = n61891 ;
  assign \po0776  = n61897 ;
  assign \po0777  = n61903 ;
  assign \po0778  = n61909 ;
  assign \po0779  = n61915 ;
  assign \po0780  = n61921 ;
  assign \po0781  = ~n61928 ;
  assign \po0782  = n61939 ;
  assign \po0783  = n61945 ;
  assign \po0784  = n61951 ;
  assign \po0785  = n61957 ;
  assign \po0786  = n61963 ;
  assign \po0787  = n61969 ;
  assign \po0788  = n61975 ;
  assign \po0789  = n61981 ;
  assign \po0790  = n61987 ;
  assign \po0791  = n61993 ;
  assign \po0792  = n61999 ;
  assign \po0793  = n62005 ;
  assign \po0794  = n62011 ;
  assign \po0795  = n62017 ;
  assign \po0796  = n62023 ;
  assign \po0797  = n62029 ;
  assign \po0798  = n62035 ;
  assign \po0799  = n62041 ;
  assign \po0800  = n62047 ;
  assign \po0801  = n62053 ;
  assign \po0802  = n62059 ;
  assign \po0803  = n62065 ;
  assign \po0804  = n62071 ;
  assign \po0805  = n62077 ;
  assign \po0806  = n62083 ;
  assign \po0807  = n62089 ;
  assign \po0808  = n62095 ;
  assign \po0809  = n62101 ;
  assign \po0810  = n62107 ;
  assign \po0811  = n62113 ;
  assign \po0812  = n62119 ;
  assign \po0813  = n62125 ;
  assign \po0814  = n62131 ;
  assign \po0815  = n62137 ;
  assign \po0816  = n62152 ;
  assign \po0817  = n62158 ;
  assign \po0818  = n62164 ;
  assign \po0819  = n62170 ;
  assign \po0820  = ~n62221 ;
  assign \po0821  = ~n62265 ;
  assign \po0822  = n62271 ;
  assign \po0823  = ~n62311 ;
  assign \po0824  = ~n62351 ;
  assign \po0825  = ~n62391 ;
  assign \po0826  = n62397 ;
  assign \po0827  = ~n62434 ;
  assign \po0828  = ~n62471 ;
  assign \po0829  = ~n62511 ;
  assign \po0830  = ~n62551 ;
  assign \po0831  = ~n62592 ;
  assign \po0832  = ~n62632 ;
  assign \po0833  = ~n62672 ;
  assign \po0834  = ~n62709 ;
  assign \po0835  = ~n62746 ;
  assign \po0836  = ~n62787 ;
  assign \po0837  = n62793 ;
  assign \po0838  = n62799 ;
  assign \po0839  = ~n62836 ;
  assign \po0840  = ~n13720 ;
  assign \po0841  = n62844 ;
  assign \po0842  = ~n62888 ;
  assign \po0843  = n62894 ;
  assign \po0844  = n62900 ;
  assign \po0845  = n62906 ;
  assign \po0846  = ~n62945 ;
  assign \po0847  = n62951 ;
  assign \po0848  = n62957 ;
  assign \po0849  = ~n62995 ;
  assign \po0850  = n63001 ;
  assign \po0851  = n63007 ;
  assign \po0852  = n63013 ;
  assign \po0853  = n63019 ;
  assign \po0854  = n63025 ;
  assign \po0855  = n63031 ;
  assign \po0856  = n63037 ;
  assign \po0857  = n63043 ;
  assign \po0858  = n63049 ;
  assign \po0859  = n63055 ;
  assign \po0860  = n63061 ;
  assign \po0861  = n63067 ;
  assign \po0862  = n63073 ;
  assign \po0863  = n63079 ;
  assign \po0864  = n63120 ;
  assign \po0865  = n63160 ;
  assign \po0866  = n63166 ;
  assign \po0867  = n63172 ;
  assign \po0868  = n63209 ;
  assign \po0869  = ~n63246 ;
  assign \po0870  = n63283 ;
  assign \po0871  = ~n63322 ;
  assign \po0872  = n63328 ;
  assign \po0873  = n63365 ;
  assign \po0874  = ~n63401 ;
  assign \po0875  = n63438 ;
  assign \po0876  = ~n63474 ;
  assign \po0877  = ~n63513 ;
  assign \po0878  = ~n63574 ;
  assign \po0879  = ~n63612 ;
  assign \po0880  = n63618 ;
  assign \po0881  = n63624 ;
  assign \po0882  = n63630 ;
  assign \po0883  = n63636 ;
  assign \po0884  = n63642 ;
  assign \po0885  = n63648 ;
  assign \po0886  = n63654 ;
  assign \po0887  = n63660 ;
  assign \po0888  = n63679 ;
  assign \po0889  = n63685 ;
  assign \po0890  = n63722 ;
  assign \po0891  = n63728 ;
  assign \po0892  = n63734 ;
  assign \po0893  = n63740 ;
  assign \po0894  = n63746 ;
  assign \po0895  = n63752 ;
  assign \po0896  = ~n63760 ;
  assign \po0897  = n61783 ;
  assign \po0898  = ~n63766 ;
  assign \po0899  = ~n63772 ;
  assign \po0900  = ~n63778 ;
  assign \po0901  = ~n63784 ;
  assign \po0902  = ~n63790 ;
  assign \po0903  = ~n63796 ;
  assign \po0904  = n63809 ;
  assign \po0905  = ~n63815 ;
  assign \po0906  = ~n63821 ;
  assign \po0907  = ~n63827 ;
  assign \po0908  = ~n63833 ;
  assign \po0909  = ~n63839 ;
  assign \po0910  = ~n63845 ;
  assign \po0911  = ~n63851 ;
  assign \po0912  = ~n63857 ;
  assign \po0913  = ~n63863 ;
  assign \po0914  = ~n63869 ;
  assign \po0915  = ~n63875 ;
  assign \po0916  = ~n63881 ;
  assign \po0917  = ~n63887 ;
  assign \po0918  = ~n63893 ;
  assign \po0919  = ~n63899 ;
  assign \po0920  = ~n63905 ;
  assign \po0921  = ~n63911 ;
  assign \po0922  = n63940 ;
  assign \po0923  = ~n63946 ;
  assign \po0924  = ~n63952 ;
  assign \po0925  = ~n63958 ;
  assign \po0926  = ~n63979 ;
  assign \po0927  = ~n63985 ;
  assign \po0928  = ~n64000 ;
  assign \po0929  = ~n64006 ;
  assign \po0930  = n64017 ;
  assign \po0931  = ~n64023 ;
  assign \po0932  = n64042 ;
  assign \po0933  = ~n64048 ;
  assign \po0934  = ~n64054 ;
  assign \po0935  = ~n64064 ;
  assign \po0936  = ~n64065 ;
  assign \po0937  = ~n64066 ;
  assign \po0938  = ~n64071 ;
  assign \po0939  = ~n64075 ;
  assign \po0940  = ~n64080 ;
  assign \po0941  = ~n64085 ;
  assign \po0942  = ~n64090 ;
  assign \po0943  = n64093 ;
  assign \po0944  = ~n64098 ;
  assign \po0945  = ~n64103 ;
  assign \po0946  = ~n64108 ;
  assign \po0947  = ~n64113 ;
  assign \po0948  = ~n64118 ;
  assign \po0949  = ~n64123 ;
  assign \po0950  = ~n59609 ;
  assign \po0951  = ~n64131 ;
  assign \po0952  = ~n64136 ;
  assign \po0953  = n64147 ;
  assign \po0954  = n61933 ;
  assign \po0955  = ~n64152 ;
  assign \po0956  = n64157 ;
  assign \po0957  = ~n64162 ;
  assign \po0958  = ~n64167 ;
  assign \po0959  = n62147 ;
  assign \po0960  = n64172 ;
  assign \po0961  = ~n64177 ;
  assign \po0962  = n64183 ;
  assign \po0963  = ~n64007 ;
  assign \po0964  = ~n64188 ;
  assign \po0965  = ~n64193 ;
  assign \po0966  = n64198 ;
  assign \po0967  = ~n64203 ;
  assign \po0968  = ~n64208 ;
  assign \po0969  = n64213 ;
  assign \po0970  = ~n64218 ;
  assign \po0971  = n64223 ;
  assign \po0972  = ~n64228 ;
  assign \po0973  = ~n64233 ;
  assign \po0974  = n64236 ;
  assign \po0975  = ~n64238 ;
  assign \po0976  = n64241 ;
  assign \po0977  = n64243 ;
  assign \po0978  = n63997 ;
  assign \po0979  = n64244 ;
  assign \po0980  = n62838 ;
  assign \po0981  = n64248 ;
  assign \po0982  = n64282 ;
  assign \po0983  = n64314 ;
  assign \po0984  = n64346 ;
  assign \po0985  = n64378 ;
  assign \po0986  = ~n64382 ;
  assign \po0987  = n64385 ;
  assign \po0988  = n63754 ;
  assign \po0989  = n64388 ;
  assign \po0990  = ~n64390 ;
  assign \po0991  = n64391 ;
  assign \po0992  = n64394 ;
  assign \po0993  = ~n64397 ;
  assign \po0994  = ~n64400 ;
  assign \po0995  = ~n64403 ;
  assign \po0996  = ~n64406 ;
  assign \po0997  = n64407 ;
  assign \po0998  = ~n64410 ;
  assign \po0999  = ~n64413 ;
  assign \po1000  = ~n64416 ;
  assign \po1001  = ~n64419 ;
  assign \po1002  = ~n64422 ;
  assign \po1003  = ~n64425 ;
  assign \po1004  = ~n64428 ;
  assign \po1005  = ~n64431 ;
  assign \po1006  = ~n64434 ;
  assign \po1007  = ~n64437 ;
  assign \po1008  = ~n64440 ;
  assign \po1009  = ~n64443 ;
  assign \po1010  = ~n64446 ;
  assign \po1011  = ~n64449 ;
  assign \po1012  = ~n64452 ;
  assign \po1013  = ~n64455 ;
  assign \po1014  = ~n64458 ;
  assign \po1015  = ~n64461 ;
  assign \po1016  = ~n64464 ;
  assign \po1017  = ~n64473 ;
  assign \po1018  = ~n64476 ;
  assign \po1019  = ~n64479 ;
  assign \po1020  = ~n64482 ;
  assign \po1021  = ~n64485 ;
  assign \po1022  = ~n64488 ;
  assign \po1023  = ~n64491 ;
  assign \po1024  = ~n64494 ;
  assign \po1025  = ~n64503 ;
  assign \po1026  = ~n64506 ;
  assign \po1027  = ~n64509 ;
  assign \po1028  = ~n64512 ;
  assign \po1029  = ~n64515 ;
  assign \po1030  = ~n64518 ;
  assign \po1031  = n64527 ;
  assign \po1032  = ~n64530 ;
  assign \po1033  = ~n64539 ;
  assign \po1034  = ~n64548 ;
  assign \po1035  = ~n64557 ;
  assign \po1036  = ~n64560 ;
  assign \po1037  = ~n64563 ;
  assign \po1038  = ~n9948 ;
  assign \po1039  = ~n64566 ;
  assign \po1040  = ~n64569 ;
  assign \po1041  = ~n64572 ;
  assign \po1042  = ~n64575 ;
  assign \po1043  = ~n64578 ;
  assign \po1044  = ~n64581 ;
  assign \po1045  = ~n64584 ;
  assign \po1046  = ~n64587 ;
  assign \po1047  = ~n64590 ;
  assign \po1048  = ~n64593 ;
  assign \po1049  = ~n1525 ;
  assign \po1050  = ~n64596 ;
  assign \po1051  = ~n64599 ;
  assign \po1052  = ~n64602 ;
  assign \po1053  = \pi0067  ;
  assign \po1054  = ~n64605 ;
  assign \po1055  = ~n64608 ;
  assign \po1056  = ~n64611 ;
  assign \po1057  = ~n6808 ;
  assign \po1058  = ~n64614 ;
  assign \po1059  = ~n64617 ;
  assign \po1060  = ~n64620 ;
  assign \po1061  = ~n64623 ;
  assign \po1062  = ~n64626 ;
  assign \po1063  = n64637 ;
  assign \po1064  = ~n64640 ;
  assign \po1065  = ~n64643 ;
  assign \po1066  = ~n64646 ;
  assign \po1067  = ~n64649 ;
  assign \po1068  = ~n64652 ;
  assign \po1069  = ~n64655 ;
  assign \po1070  = n64657 ;
  assign \po1071  = ~n64660 ;
  assign \po1072  = ~n64663 ;
  assign \po1073  = ~n64666 ;
  assign \po1074  = ~n64669 ;
  assign \po1075  = ~n64672 ;
  assign \po1076  = ~n64675 ;
  assign \po1077  = ~n64677 ;
  assign \po1078  = n64680 ;
  assign \po1079  = n64683 ;
  assign \po1080  = n64685 ;
  assign \po1081  = n64688 ;
  assign \po1082  = n64691 ;
  assign \po1083  = n64694 ;
  assign \po1084  = n64696 ;
  assign \po1085  = n64699 ;
  assign \po1086  = n64702 ;
  assign \po1087  = n64705 ;
  assign \po1088  = ~n64707 ;
  assign \po1089  = ~n64709 ;
  assign \po1090  = n64712 ;
  assign \po1091  = ~n64714 ;
  assign \po1092  = n64717 ;
  assign \po1093  = n64720 ;
  assign \po1094  = ~n64722 ;
  assign \po1095  = n64725 ;
  assign \po1096  = ~n64727 ;
  assign \po1097  = n64730 ;
  assign \po1098  = n64733 ;
  assign \po1099  = n64736 ;
  assign \po1100  = ~n64739 ;
  assign \po1101  = ~n6713 ;
  assign \po1102  = n64740 ;
  assign \po1103  = ~n64742 ;
  assign \po1104  = n64744 ;
  assign \po1105  = ~n64747 ;
  assign \po1106  = n64748 ;
  assign \po1107  = n64749 ;
  assign \po1108  = \pi1134  ;
  assign \po1109  = \pi0964  ;
  assign \po1110  = ~\pi0954  ;
  assign \po1111  = \pi0965  ;
  assign \po1112  = ~n64751 ;
  assign \po1113  = \pi0991  ;
  assign \po1114  = \pi0985  ;
  assign \po1115  = n64752 ;
  assign \po1116  = n64753 ;
  assign \po1117  = \pi1014  ;
  assign \po1118  = n64754 ;
  assign \po1119  = \pi1029  ;
  assign \po1120  = \pi1004  ;
  assign \po1121  = \pi1007  ;
  assign \po1122  = n64755 ;
  assign \po1123  = \pi1135  ;
  assign \po1124  = n64756 ;
  assign \po1125  = n64757 ;
  assign \po1126  = n64758 ;
  assign \po1127  = n64759 ;
  assign \po1128  = n64760 ;
  assign \po1129  = n64761 ;
  assign \po1130  = ~\pi0278  ;
  assign \po1131  = n64762 ;
  assign \po1132  = n64763 ;
  assign \po1133  = ~n64764 ;
  assign \po1134  = \pi1064  ;
  assign \po1135  = n64765 ;
  assign \po1136  = \pi0299  ;
  assign \po1137  = ~n64766 ;
  assign \po1138  = \pi1075  ;
  assign \po1139  = \pi1052  ;
  assign \po1140  = \pi0771  ;
  assign \po1141  = \pi0765  ;
  assign \po1142  = \pi0605  ;
  assign \po1143  = \pi0601  ;
  assign \po1144  = \pi0278  ;
  assign \po1145  = \pi0279  ;
  assign \po1146  = ~\pi0915  ;
  assign \po1147  = ~\pi0825  ;
  assign \po1148  = ~\pi0826  ;
  assign \po1149  = ~\pi0913  ;
  assign \po1150  = ~\pi0894  ;
  assign \po1151  = ~\pi0905  ;
  assign \po1152  = \pi1095  ;
  assign \po1153  = ~\pi0890  ;
  assign \po1154  = \pi1094  ;
  assign \po1155  = ~\pi0906  ;
  assign \po1156  = ~\pi0896  ;
  assign \po1157  = ~\pi0909  ;
  assign \po1158  = ~\pi0911  ;
  assign \po1159  = ~\pi0908  ;
  assign \po1160  = ~\pi0891  ;
  assign \po1161  = ~\pi0902  ;
  assign \po1162  = ~\pi0903  ;
  assign \po1163  = ~\pi0883  ;
  assign \po1164  = ~\pi0888  ;
  assign \po1165  = ~\pi0919  ;
  assign \po1166  = ~\pi0886  ;
  assign \po1167  = ~\pi0912  ;
  assign \po1168  = ~\pi0895  ;
  assign \po1169  = ~\pi0916  ;
  assign \po1170  = ~\pi0889  ;
  assign \po1171  = ~\pi0900  ;
  assign \po1172  = ~\pi0885  ;
  assign \po1173  = ~\pi0904  ;
  assign \po1174  = ~\pi0899  ;
  assign \po1175  = ~\pi0918  ;
  assign \po1176  = ~\pi0898  ;
  assign \po1177  = ~\pi0917  ;
  assign \po1178  = ~\pi0827  ;
  assign \po1179  = ~\pi0887  ;
  assign \po1180  = ~\pi0884  ;
  assign \po1181  = ~\pi0910  ;
  assign \po1182  = ~\pi0828  ;
  assign \po1183  = ~\pi0892  ;
  assign \po1184  = \pi1187  ;
  assign \po1185  = \pi1172  ;
  assign \po1186  = \pi1170  ;
  assign \po1187  = \pi1138  ;
  assign \po1188  = \pi1177  ;
  assign \po1189  = \pi1178  ;
  assign \po1190  = \pi0863  ;
  assign \po1191  = \pi1203  ;
  assign \po1192  = \pi1185  ;
  assign \po1193  = \pi1171  ;
  assign \po1194  = \pi1192  ;
  assign \po1195  = \pi1137  ;
  assign \po1196  = \pi1186  ;
  assign \po1197  = \pi1165  ;
  assign \po1198  = \pi1164  ;
  assign \po1199  = \pi1098  ;
  assign \po1200  = \pi1183  ;
  assign \po1201  = \pi0230  ;
  assign \po1202  = \pi1169  ;
  assign \po1203  = \pi1136  ;
  assign \po1204  = \pi1181  ;
  assign \po1205  = \pi0849  ;
  assign \po1206  = \pi1193  ;
  assign \po1207  = \pi1182  ;
  assign \po1208  = \pi1168  ;
  assign \po1209  = \pi1175  ;
  assign \po1210  = \pi1191  ;
  assign \po1211  = \pi1099  ;
  assign \po1212  = \pi1174  ;
  assign \po1213  = \pi1179  ;
  assign \po1214  = \pi1202  ;
  assign \po1215  = \pi1176  ;
  assign \po1216  = \pi1173  ;
  assign \po1217  = \pi1201  ;
  assign \po1218  = \pi1167  ;
  assign \po1219  = \pi0840  ;
  assign \po1220  = \pi1189  ;
  assign \po1221  = \pi1195  ;
  assign \po1222  = \pi0864  ;
  assign \po1223  = \pi1190  ;
  assign \po1224  = \pi1188  ;
  assign \po1225  = \pi1180  ;
  assign \po1226  = \pi1194  ;
  assign \po1227  = \pi1097  ;
  assign \po1228  = \pi1166  ;
  assign \po1229  = \pi1200  ;
  assign \po1230  = \pi1184  ;
endmodule
