module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, \j0_pad , j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u0_pad , \v0_pad , \w0_pad , \x0_pad , \y0_pad , \z0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u0_pad  ;
	output \v0_pad  ;
	output \w0_pad  ;
	output \x0_pad  ;
	output \y0_pad  ;
	output \z0_pad  ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		p_pad,
		q_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		r_pad,
		u_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		r_pad,
		u_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w37_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		q_pad,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		s_pad,
		_w36_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		o_pad,
		q_pad,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		v_pad,
		_w37_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		v_pad,
		_w37_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		q_pad,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		s_pad,
		_w43_,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		n_pad,
		q_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		w_pad,
		_w45_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		w_pad,
		_w45_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		q_pad,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		s_pad,
		_w50_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		m_pad,
		q_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		x_pad,
		_w51_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		x_pad,
		_w51_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		q_pad,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		s_pad,
		_w57_,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		l_pad,
		q_pad,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		y_pad,
		_w58_,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		y_pad,
		_w58_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w65_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		q_pad,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		s_pad,
		_w64_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w68_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		k_pad,
		q_pad,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		z_pad,
		_w65_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		z_pad,
		_w65_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w72_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		q_pad,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		s_pad,
		_w71_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		j_pad,
		q_pad,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\a0_pad ,
		_w72_,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\a0_pad ,
		_w72_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		q_pad,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		s_pad,
		_w78_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		i_pad,
		q_pad,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\b0_pad ,
		_w79_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\b0_pad ,
		_w79_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		q_pad,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		s_pad,
		_w85_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		h_pad,
		q_pad,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\c0_pad ,
		_w86_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\c0_pad ,
		_w86_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		q_pad,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		s_pad,
		_w92_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		g_pad,
		q_pad,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		\d0_pad ,
		_w93_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\d0_pad ,
		_w93_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		q_pad,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		s_pad,
		_w99_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		f_pad,
		q_pad,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		\e0_pad ,
		_w100_,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\e0_pad ,
		_w100_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w107_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		q_pad,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		s_pad,
		_w106_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		e_pad,
		q_pad,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\f0_pad ,
		_w107_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\f0_pad ,
		_w107_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		q_pad,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		s_pad,
		_w113_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		d_pad,
		q_pad,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\g0_pad ,
		_w114_,
		_w121_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\g0_pad ,
		_w114_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		q_pad,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		s_pad,
		_w120_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w124_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		c_pad,
		q_pad,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\h0_pad ,
		_w121_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\h0_pad ,
		_w121_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		q_pad,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		s_pad,
		_w127_,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w131_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		b_pad,
		q_pad,
		_w134_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		\i0_pad ,
		_w128_,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\i0_pad ,
		_w128_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w135_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		q_pad,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		s_pad,
		_w134_,
		_w139_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		a_pad,
		q_pad,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\j0_pad ,
		_w135_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\j0_pad ,
		_w135_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		q_pad,
		_w142_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		s_pad,
		_w141_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w145_,
		_w146_,
		_w147_
	);
	assign \k0_pad  = _w42_ ;
	assign \l0_pad  = _w49_ ;
	assign \m0_pad  = _w56_ ;
	assign \n0_pad  = _w63_ ;
	assign \o0_pad  = _w70_ ;
	assign \p0_pad  = _w77_ ;
	assign \q0_pad  = _w84_ ;
	assign \r0_pad  = _w91_ ;
	assign \s0_pad  = _w98_ ;
	assign \t0_pad  = _w105_ ;
	assign \u0_pad  = _w112_ ;
	assign \v0_pad  = _w119_ ;
	assign \w0_pad  = _w126_ ;
	assign \x0_pad  = _w133_ ;
	assign \y0_pad  = _w140_ ;
	assign \z0_pad  = _w147_ ;
endmodule;