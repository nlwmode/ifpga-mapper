module top (\g1000_reg/NET0131 , \g1001_reg/NET0131 , \g1002_reg/NET0131 , \g1003_reg/NET0131 , \g1004_reg/NET0131 , \g1005_reg/NET0131 , \g1006_reg/NET0131 , \g1007_reg/NET0131 , \g1008_reg/NET0131 , \g1009_reg/NET0131 , \g1010_reg/NET0131 , \g1011_reg/NET0131 , \g1018_reg/NET0131 , \g101_reg/NET0131 , \g1024_reg/NET0131 , \g1030_reg/NET0131 , \g1033_reg/NET0131 , \g1036_reg/NET0131 , \g1038_reg/NET0131 , \g1040_reg/NET0131 , \g1041_reg/NET0131 , \g1045_reg/NET0131 , \g1048_reg/NET0131 , \g1051_reg/NET0131 , \g1053_reg/NET0131 , \g1055_reg/NET0131 , \g1056_reg/NET0131 , \g105_reg/NET0131 , \g1060_reg/NET0131 , \g1063_reg/NET0131 , \g1066_reg/NET0131 , \g1068_reg/NET0131 , \g1070_reg/NET0131 , \g1071_reg/NET0131 , \g1075_reg/NET0131 , \g1078_reg/NET0131 , \g1081_reg/NET0131 , \g1083_reg/NET0131 , \g1085_reg/NET0131 , \g1088_reg/NET0131 , \g1089_reg/NET0131 , \g1090_reg/NET0131 , \g1091_reg/NET0131 , \g1092_reg/NET0131 , \g1095_reg/NET0131 , \g1098_reg/NET0131 , \g109_reg/NET0131 , \g1101_reg/NET0131 , \g1104_reg/NET0131 , \g1107_reg/NET0131 , \g1110_reg/NET0131 , \g1113_reg/NET0131 , \g1114_reg/NET0131 , \g1115_reg/NET0131 , \g1116_reg/NET0131 , \g1119_reg/NET0131 , \g1122_reg/NET0131 , \g1125_reg/NET0131 , \g1128_reg/NET0131 , \g1131_reg/NET0131 , \g1134_reg/NET0131 , \g1135_reg/NET0131 , \g1136_reg/NET0131 , \g1138_reg/NET0131 , \g113_reg/NET0131 , \g1140_reg/NET0131 , \g1151_reg/NET0131 , \g1164_reg/NET0131 , \g1165_reg/NET0131 , \g1166_reg/NET0131 , \g1167_reg/NET0131 , \g1171_reg/NET0131 , \g1173_reg/NET0131 , \g1174_reg/NET0131 , \g1175_reg/NET0131 , \g1176_reg/NET0131 , \g1177_reg/NET0131 , \g117_reg/NET0131 , \g1180_reg/NET0131 , \g1183_reg/NET0131 , \g1186_reg/NET0131 , \g1192_reg/NET0131 , \g1193_reg/NET0131 , \g1196_reg/NET0131 , \g1210_reg/NET0131 , \g1211_reg/NET0131 , \g1215_reg/NET0131 , \g1216_reg/NET0131 , \g1217_reg/NET0131 , \g1218_reg/NET0131 , \g1219_reg/NET0131 , \g121_reg/NET0131 , \g1220_reg/NET0131 , \g1222_reg/NET0131 , \g1223_reg/NET0131 , \g1224_reg/NET0131 , \g1227_reg/NET0131 , \g1228_reg/NET0131 , \g1230_reg/NET0131 , \g1234_reg/NET0131 , \g1240_reg/NET0131 , \g1243_reg/NET0131 , \g1245_reg/NET0131 , \g1249_pad , \g1251_reg/NET0131 , \g1253_reg/NET0131 , \g1255_reg/NET0131 , \g1257_reg/NET0131 , \g1259_reg/NET0131 , \g125_reg/NET0131 , \g1261_reg/NET0131 , \g1262_reg/NET0131 , \g1263_reg/NET0131 , \g1264_reg/NET0131 , \g1265_reg/NET0131 , \g1266_reg/NET0131 , \g1267_reg/NET0131 , \g1268_reg/NET0131 , \g1269_reg/NET0131 , \g1270_reg/NET0131 , \g1271_reg/NET0131 , \g1272_reg/NET0131 , \g1273_reg/NET0131 , \g1276_reg/NET0131 , \g1279_reg/NET0131 , \g1282_reg/NET0131 , \g1285_reg/NET0131 , \g1288_reg/NET0131 , \g1291_reg/NET0131 , \g1294_reg/NET0131 , \g1297_reg/NET0131 , \g129_reg/NET0131 , \g1300_reg/NET0131 , \g1303_reg/NET0131 , \g1306_reg/NET0131 , \g130_reg/NET0131 , \g1316_reg/NET0131 , \g1319_reg/NET0131 , \g131_reg/NET0131 , \g1326_reg/NET0131 , \g132_reg/NET0131 , \g1332_reg/NET0131 , \g1339_reg/NET0131 , \g133_reg/NET0131 , \g1345_reg/NET0131 , \g1346_reg/NET0131 , \g134_reg/NET0131 , \g1352_reg/NET0131 , \g1358_reg/NET0131 , \g1365_reg/NET0131 , \g1372_reg/NET0131 , \g1378_reg/NET0131 , \g1384_reg/NET0131 , \g1385_reg/NET0131 , \g1386_reg/NET0131 , \g1387_reg/NET0131 , \g1388_reg/NET0131 , \g1389_reg/NET0131 , \g1390_reg/NET0131 , \g1391_reg/NET0131 , \g1392_reg/NET0131 , \g1393_reg/NET0131 , \g1394_reg/NET0131 , \g1395_reg/NET0131 , \g1396_reg/NET0131 , \g1397_reg/NET0131 , \g1398_reg/NET0131 , \g1399_reg/NET0131 , \g1400_reg/NET0131 , \g1401_reg/NET0131 , \g1402_reg/NET0131 , \g1403_reg/NET0131 , \g1404_reg/NET0131 , \g1405_reg/NET0131 , \g1406_reg/NET0131 , \g1407_reg/NET0131 , \g1408_reg/NET0131 , \g1409_reg/NET0131 , \g1410_reg/NET0131 , \g1411_reg/NET0131 , \g1412_reg/NET0131 , \g1413_reg/NET0131 , \g1414_reg/NET0131 , \g1415_reg/NET0131 , \g1416_reg/NET0131 , \g1417_reg/NET0131 , \g1418_reg/NET0131 , \g1419_reg/NET0131 , \g141_reg/NET0131 , \g1420_reg/NET0131 , \g1421_reg/NET0131 , \g1422_reg/NET0131 , \g1423_reg/NET0131 , \g1424_reg/NET0131 , \g1425_reg/NET0131 , \g1426_reg/NET0131 , \g142_reg/NET0131 , \g1430_reg/NET0131 , \g1435_reg/NET0131 , \g1439_reg/NET0131 , \g143_reg/NET0131 , \g1444_reg/NET0131 , \g1448_reg/NET0131 , \g144_reg/NET0131 , \g1453_reg/NET0131 , \g1457_reg/NET0131 , \g145_reg/NET0131 , \g1462_reg/NET0131 , \g1466_reg/NET0131 , \g146_reg/NET0131 , \g1471_reg/NET0131 , \g1476_reg/NET0131 , \g147_reg/NET0131 , \g1481_reg/NET0131 , \g1486_reg/NET0131 , \g148_reg/NET0131 , \g1491_reg/NET0131 , \g1496_reg/NET0131 , \g149_reg/NET0131 , \g1501_reg/NET0131 , \g1506_reg/NET0131 , \g150_reg/NET0131 , \g1511_reg/NET0131 , \g1512_reg/NET0131 , \g1513_reg/NET0131 , \g1514_reg/NET0131 , \g1515_reg/NET0131 , \g1516_reg/NET0131 , \g151_reg/NET0131 , \g1523_reg/NET0131 , \g1524_reg/NET0131 , \g1525_reg/NET0131 , \g1526_reg/NET0131 , \g1527_reg/NET0131 , \g1528_reg/NET0131 , \g1529_reg/NET0131 , \g152_reg/NET0131 , \g1530_reg/NET0131 , \g1531_reg/NET0131 , \g1532_reg/NET0131 , \g1533_reg/NET0131 , \g1534_reg/NET0131 , \g1535_reg/NET0131 , \g1536_reg/NET0131 , \g1537_reg/NET0131 , \g1538_reg/NET0131 , \g1539_reg/NET0131 , \g153_reg/NET0131 , \g1540_reg/NET0131 , \g1541_reg/NET0131 , \g1542_reg/NET0131 , \g1543_reg/NET0131 , \g1544_reg/NET0131 , \g1545_reg/NET0131 , \g1546_reg/NET0131 , \g154_reg/NET0131 , \g1550_reg/NET0131 , \g1551_reg/NET0131 , \g1552_reg/NET0131 , \g1553_reg/NET0131 , \g1554_reg/NET0131 , \g1555_reg/NET0131 , \g1556_reg/NET0131 , \g1557_reg/NET0131 , \g1558_reg/NET0131 , \g1559_reg/NET0131 , \g155_reg/NET0131 , \g1560_reg/NET0131 , \g1561_reg/NET0131 , \g1563_reg/NET0131 , \g1567_reg/NET0131 , \g156_reg/NET0131 , \g1570_reg/NET0131 , \g1573_reg/NET0131 , \g1576_reg/NET0131 , \g1579_reg/NET0131 , \g157_reg/NET0131 , \g1582_reg/NET0131 , \g1585_reg/NET0131 , \g1588_reg/NET0131 , \g158_reg/NET0131 , \g1591_reg/NET0131 , \g1594_reg/NET0131 , \g1597_reg/NET0131 , \g159_reg/NET0131 , \g1600_reg/NET0131 , \g1603_reg/NET0131 , \g1606_reg/NET0131 , \g1609_reg/NET0131 , \g160_reg/NET0131 , \g1612_reg/NET0131 , \g1615_reg/NET0131 , \g1618_reg/NET0131 , \g161_reg/NET0131 , \g1621_reg/NET0131 , \g1624_reg/NET0131 , \g1627_reg/NET0131 , \g16297_pad , \g162_reg/NET0131 , \g1630_reg/NET0131 , \g1633_reg/NET0131 , \g16355_pad , \g1636_reg/NET0131 , \g16399_pad , \g1639_reg/NET0131 , \g163_reg/NET0131 , \g1642_reg/NET0131 , \g16437_pad , \g1645_reg/NET0131 , \g1648_reg/NET0131 , \g164_reg/NET0131 , \g1651_reg/NET0131 , \g1654_reg/NET0131 , \g1660_reg/NET0131 , \g1662_reg/NET0131 , \g1664_reg/NET0131 , \g1666_reg/NET0131 , \g1668_reg/NET0131 , \g1670_reg/NET0131 , \g1672_reg/NET0131 , \g1679_reg/NET0131 , \g1680_reg/NET0131 , \g1686_reg/NET0131 , \g168_reg/NET0131 , \g1693_reg/NET0131 , \g1694_reg/NET0131 , \g1695_reg/NET0131 , \g1696_reg/NET0131 , \g1697_reg/NET0131 , \g1698_reg/NET0131 , \g1699_reg/NET0131 , \g169_reg/NET0131 , \g1700_reg/NET0131 , \g1701_reg/NET0131 , \g1702_reg/NET0131 , \g1703_reg/NET0131 , \g1704_reg/NET0131 , \g1705_reg/NET0131 , \g170_reg/NET0131 , \g171_reg/NET0131 , \g1724_reg/NET0131 , \g1727_reg/NET0131 , \g172_reg/NET0131 , \g1730_reg/NET0131 , \g1732_reg/NET0131 , \g1734_reg/NET0131 , \g1735_reg/NET0131 , \g1739_reg/NET0131 , \g173_reg/NET0131 , \g1742_reg/NET0131 , \g1745_reg/NET0131 , \g1747_reg/NET0131 , \g1749_reg/NET0131 , \g174_reg/NET0131 , \g1750_reg/NET0131 , \g1754_reg/NET0131 , \g1757_reg/NET0131 , \g175_reg/NET0131 , \g1760_reg/NET0131 , \g1762_reg/NET0131 , \g1764_reg/NET0131 , \g1765_reg/NET0131 , \g1769_reg/NET0131 , \g176_reg/NET0131 , \g1772_reg/NET0131 , \g1775_reg/NET0131 , \g1777_reg/NET0131 , \g1779_reg/NET0131 , \g177_reg/NET0131 , \g1783_reg/NET0131 , \g1784_reg/NET0131 , \g1785_reg/NET0131 , \g1789_reg/NET0131 , \g178_reg/NET0131 , \g1792_reg/NET0131 , \g1795_reg/NET0131 , \g1798_reg/NET0131 , \g179_reg/NET0131 , \g1801_reg/NET0131 , \g1804_reg/NET0131 , \g1807_reg/NET0131 , \g1808_reg/NET0131 , \g1809_reg/NET0131 , \g1810_reg/NET0131 , \g1813_reg/NET0131 , \g1816_reg/NET0131 , \g1819_reg/NET0131 , \g1822_reg/NET0131 , \g1825_reg/NET0131 , \g1828_reg/NET0131 , \g1829_reg/NET0131 , \g1830_reg/NET0131 , \g1832_reg/NET0131 , \g1834_reg/NET0131 , \g1845_reg/NET0131 , \g1846_reg/NET0131 , \g1849_reg/NET0131 , \g1852_reg/NET0131 , \g1858_reg/NET0131 , \g1859_reg/NET0131 , \g185_reg/NET0131 , \g1860_reg/NET0131 , \g1861_reg/NET0131 , \g1865_reg/NET0131 , \g1867_reg/NET0131 , \g1868_reg/NET0131 , \g1869_reg/NET0131 , \g186_reg/NET0131 , \g1870_reg/NET0131 , \g1871_reg/NET0131 , \g1874_reg/NET0131 , \g1877_reg/NET0131 , \g1880_reg/NET0131 , \g1886_reg/NET0131 , \g1887_reg/NET0131 , \g189_reg/NET0131 , \g1904_reg/NET0131 , \g1905_reg/NET0131 , \g1909_reg/NET0131 , \g1910_reg/NET0131 , \g1911_reg/NET0131 , \g1912_reg/NET0131 , \g1913_reg/NET0131 , \g1914_reg/NET0131 , \g1916_reg/NET0131 , \g1917_reg/NET0131 , \g1918_reg/NET0131 , \g1921_reg/NET0131 , \g1922_reg/NET0131 , \g1924_reg/NET0131 , \g1928_reg/NET0131 , \g192_reg/NET0131 , \g1939_reg/NET0131 , \g1943_pad , \g1945_reg/NET0131 , \g1947_reg/NET0131 , \g1949_reg/NET0131 , \g1951_reg/NET0131 , \g1953_reg/NET0131 , \g1955_reg/NET0131 , \g1956_reg/NET0131 , \g1957_reg/NET0131 , \g1958_reg/NET0131 , \g1959_reg/NET0131 , \g195_reg/NET0131 , \g1960_reg/NET0131 , \g1961_reg/NET0131 , \g1962_reg/NET0131 , \g1963_reg/NET0131 , \g1964_reg/NET0131 , \g1965_reg/NET0131 , \g1966_reg/NET0131 , \g1967_reg/NET0131 , \g1970_reg/NET0131 , \g1973_reg/NET0131 , \g1976_reg/NET0131 , \g1979_reg/NET0131 , \g1982_reg/NET0131 , \g1985_reg/NET0131 , \g1988_reg/NET0131 , \g198_reg/NET0131 , \g1991_reg/NET0131 , \g1994_reg/NET0131 , \g1997_reg/NET0131 , \g2000_reg/NET0131 , \g201_reg/NET0131 , \g204_reg/NET0131 , \g2078_reg/NET0131 , \g2079_reg/NET0131 , \g207_reg/NET0131 , \g2080_reg/NET0131 , \g2081_reg/NET0131 , \g2082_reg/NET0131 , \g2083_reg/NET0131 , \g2084_reg/NET0131 , \g2085_reg/NET0131 , \g2086_reg/NET0131 , \g2087_reg/NET0131 , \g2088_reg/NET0131 , \g2089_reg/NET0131 , \g2090_reg/NET0131 , \g2091_reg/NET0131 , \g2092_reg/NET0131 , \g2093_reg/NET0131 , \g2094_reg/NET0131 , \g2095_reg/NET0131 , \g2096_reg/NET0131 , \g2097_reg/NET0131 , \g2098_reg/NET0131 , \g2099_reg/NET0131 , \g2100_reg/NET0131 , \g2101_reg/NET0131 , \g2102_reg/NET0131 , \g2103_reg/NET0131 , \g2104_reg/NET0131 , \g2105_reg/NET0131 , \g2106_reg/NET0131 , \g2107_reg/NET0131 , \g2108_reg/NET0131 , \g2109_reg/NET0131 , \g210_reg/NET0131 , \g2110_reg/NET0131 , \g2111_reg/NET0131 , \g2112_reg/NET0131 , \g2113_reg/NET0131 , \g2114_reg/NET0131 , \g2115_reg/NET0131 , \g2116_reg/NET0131 , \g2117_reg/NET0131 , \g2118_reg/NET0131 , \g2119_reg/NET0131 , \g213_reg/NET0131 , \g2165_reg/NET0131 , \g216_reg/NET0131 , \g2170_reg/NET0131 , \g2175_reg/NET0131 , \g2180_reg/NET0131 , \g2185_reg/NET0131 , \g2190_reg/NET0131 , \g2195_reg/NET0131 , \g219_reg/NET0131 , \g2200_reg/NET0131 , \g2205_reg/NET0131 , \g2206_reg/NET0131 , \g2207_reg/NET0131 , \g2208_reg/NET0131 , \g2209_reg/NET0131 , \g2210_reg/NET0131 , \g2217_reg/NET0131 , \g2218_reg/NET0131 , \g2219_reg/NET0131 , \g2220_reg/NET0131 , \g2221_reg/NET0131 , \g2222_reg/NET0131 , \g2223_reg/NET0131 , \g2224_reg/NET0131 , \g2225_reg/NET0131 , \g2226_reg/NET0131 , \g2227_reg/NET0131 , \g2228_reg/NET0131 , \g2229_reg/NET0131 , \g222_reg/NET0131 , \g2230_reg/NET0131 , \g2231_reg/NET0131 , \g2232_reg/NET0131 , \g2233_reg/NET0131 , \g2234_reg/NET0131 , \g2235_reg/NET0131 , \g2236_reg/NET0131 , \g2237_reg/NET0131 , \g2238_reg/NET0131 , \g2239_reg/NET0131 , \g2240_reg/NET0131 , \g2244_reg/NET0131 , \g2245_reg/NET0131 , \g2246_reg/NET0131 , \g2247_reg/NET0131 , \g2248_reg/NET0131 , \g2249_reg/NET0131 , \g2250_reg/NET0131 , \g2251_reg/NET0131 , \g2252_reg/NET0131 , \g2253_reg/NET0131 , \g2254_reg/NET0131 , \g2255_reg/NET0131 , \g225_reg/NET0131 , \g2261_reg/NET0131 , \g2264_reg/NET0131 , \g2267_reg/NET0131 , \g2270_reg/NET0131 , \g2273_reg/NET0131 , \g2276_reg/NET0131 , \g2279_reg/NET0131 , \g2282_reg/NET0131 , \g2285_reg/NET0131 , \g2288_reg/NET0131 , \g228_reg/NET0131 , \g2291_reg/NET0131 , \g2294_reg/NET0131 , \g2297_reg/NET0131 , \g2300_reg/NET0131 , \g2303_reg/NET0131 , \g2306_reg/NET0131 , \g2309_reg/NET0131 , \g2312_reg/NET0131 , \g2315_reg/NET0131 , \g2318_reg/NET0131 , \g231_reg/NET0131 , \g2321_reg/NET0131 , \g2324_reg/NET0131 , \g2327_reg/NET0131 , \g2330_reg/NET0131 , \g2333_reg/NET0131 , \g2336_reg/NET0131 , \g2339_reg/NET0131 , \g2342_reg/NET0131 , \g2345_reg/NET0131 , \g2348_reg/NET0131 , \g234_reg/NET0131 , \g2354_reg/NET0131 , \g2356_reg/NET0131 , \g2358_reg/NET0131 , \g2360_reg/NET0131 , \g2362_reg/NET0131 , \g2364_reg/NET0131 , \g2366_reg/NET0131 , \g2373_reg/NET0131 , \g2374_reg/NET0131 , \g237_reg/NET0131 , \g2380_reg/NET0131 , \g2387_reg/NET0131 , \g2388_reg/NET0131 , \g2389_reg/NET0131 , \g2390_reg/NET0131 , \g2391_reg/NET0131 , \g2392_reg/NET0131 , \g2393_reg/NET0131 , \g2394_reg/NET0131 , \g2395_reg/NET0131 , \g2396_reg/NET0131 , \g2397_reg/NET0131 , \g2398_reg/NET0131 , \g2399_reg/NET0131 , \g240_reg/NET0131 , \g2418_reg/NET0131 , \g2421_reg/NET0131 , \g2424_reg/NET0131 , \g2426_reg/NET0131 , \g2428_reg/NET0131 , \g2429_reg/NET0131 , \g2433_reg/NET0131 , \g2436_reg/NET0131 , \g2439_reg/NET0131 , \g243_reg/NET0131 , \g2441_reg/NET0131 , \g2443_reg/NET0131 , \g2444_reg/NET0131 , \g2448_reg/NET0131 , \g2451_reg/NET0131 , \g2454_reg/NET0131 , \g2456_reg/NET0131 , \g2458_reg/NET0131 , \g2459_reg/NET0131 , \g2463_reg/NET0131 , \g2466_reg/NET0131 , \g2469_reg/NET0131 , \g246_reg/NET0131 , \g2471_reg/NET0131 , \g2473_reg/NET0131 , \g2477_reg/NET0131 , \g2478_reg/NET0131 , \g2479_reg/NET0131 , \g2483_reg/NET0131 , \g2486_reg/NET0131 , \g2489_reg/NET0131 , \g2492_reg/NET0131 , \g2495_reg/NET0131 , \g2498_reg/NET0131 , \g249_reg/NET0131 , \g2501_reg/NET0131 , \g2502_reg/NET0131 , \g2503_reg/NET0131 , \g2504_reg/NET0131 , \g2507_reg/NET0131 , \g2510_reg/NET0131 , \g2513_reg/NET0131 , \g2516_reg/NET0131 , \g2519_reg/NET0131 , \g2522_reg/NET0131 , \g2523_reg/NET0131 , \g2524_reg/NET0131 , \g2526_reg/NET0131 , \g2528_reg/NET0131 , \g252_reg/NET0131 , \g2539_reg/NET0131 , \g2540_reg/NET0131 , \g2543_reg/NET0131 , \g2546_reg/NET0131 , \g2552_reg/NET0131 , \g2553_reg/NET0131 , \g2554_reg/NET0131 , \g2555_reg/NET0131 , \g2559_reg/NET0131 , \g255_reg/NET0131 , \g2561_reg/NET0131 , \g2562_reg/NET0131 , \g2563_reg/NET0131 , \g2564_reg/NET0131 , \g2565_reg/NET0131 , \g2568_reg/NET0131 , \g2571_reg/NET0131 , \g2574_reg/NET0131 , \g2580_reg/NET0131 , \g2581_reg/NET0131 , \g258_reg/NET0131 , \g2598_reg/NET0131 , \g2599_reg/NET0131 , \g2603_reg/NET0131 , \g2604_reg/NET0131 , \g2605_reg/NET0131 , \g2606_reg/NET0131 , \g2607_reg/NET0131 , \g2608_reg/NET0131 , \g2610_reg/NET0131 , \g2611_reg/NET0131 , \g2612_reg/NET0131 , \g2615_reg/NET0131 , \g2616_reg/NET0131 , \g2618_reg/NET0131 , \g261_reg/NET0131 , \g2622_reg/NET0131 , \g2633_reg/NET0131 , \g2637_pad , \g2639_reg/NET0131 , \g2641_reg/NET0131 , \g2643_reg/NET0131 , \g2645_reg/NET0131 , \g2647_reg/NET0131 , \g2649_reg/NET0131 , \g264_reg/NET0131 , \g2650_reg/NET0131 , \g2651_reg/NET0131 , \g2652_reg/NET0131 , \g2653_reg/NET0131 , \g2654_reg/NET0131 , \g2655_reg/NET0131 , \g2656_reg/NET0131 , \g2657_reg/NET0131 , \g2658_reg/NET0131 , \g2659_reg/NET0131 , \g2660_reg/NET0131 , \g2661_reg/NET0131 , \g2664_reg/NET0131 , \g2667_reg/NET0131 , \g2670_reg/NET0131 , \g2673_reg/NET0131 , \g2676_reg/NET0131 , \g2679_reg/NET0131 , \g267_reg/NET0131 , \g2682_reg/NET0131 , \g2685_reg/NET0131 , \g2688_reg/NET0131 , \g2691_reg/NET0131 , \g2694_reg/NET0131 , \g270_reg/NET0131 , \g273_reg/NET0131 , \g2772_reg/NET0131 , \g2773_reg/NET0131 , \g2774_reg/NET0131 , \g2775_reg/NET0131 , \g2776_reg/NET0131 , \g2777_reg/NET0131 , \g2778_reg/NET0131 , \g2779_reg/NET0131 , \g2780_reg/NET0131 , \g2781_reg/NET0131 , \g2782_reg/NET0131 , \g2783_reg/NET0131 , \g2784_reg/NET0131 , \g2785_reg/NET0131 , \g2786_reg/NET0131 , \g2787_reg/NET0131 , \g2788_reg/NET0131 , \g2789_reg/NET0131 , \g2790_reg/NET0131 , \g2791_reg/NET0131 , \g2792_reg/NET0131 , \g2793_reg/NET0131 , \g2794_reg/NET0131 , \g2795_reg/NET0131 , \g2796_reg/NET0131 , \g2797_reg/NET0131 , \g2798_reg/NET0131 , \g2799_reg/NET0131 , \g279_reg/NET0131 , \g2800_reg/NET0131 , \g2801_reg/NET0131 , \g2802_reg/NET0131 , \g2803_reg/NET0131 , \g2804_reg/NET0131 , \g2805_reg/NET0131 , \g2806_reg/NET0131 , \g2807_reg/NET0131 , \g2808_reg/NET0131 , \g2809_reg/NET0131 , \g2810_reg/NET0131 , \g2811_reg/NET0131 , \g2812_reg/NET0131 , \g2813_reg/NET0131 , \g2814_reg/NET0131 , \g2817_reg/NET0131 , \g281_reg/NET0131 , \g283_reg/NET0131 , \g285_reg/NET0131 , \g2874_reg/NET0131 , \g2879_reg/NET0131 , \g287_reg/NET0131 , \g2883_reg/NET0131 , \g2888_reg/NET0131 , \g2892_reg/NET0131 , \g2896_reg/NET0131 , \g289_reg/NET0131 , \g2900_reg/NET0131 , \g2903_reg/NET0131 , \g2908_reg/NET0131 , \g2912_reg/NET0131 , \g2917_reg/NET0131 , \g291_reg/NET0131 , \g2920_reg/NET0131 , \g2924_reg/NET0131 , \g2929_reg/NET0131 , \g2933_reg/NET0131 , \g2934_reg/NET0131 , \g2935_reg/NET0131 , \g2938_reg/NET0131 , \g2941_reg/NET0131 , \g2944_reg/NET0131 , \g2947_reg/NET0131 , \g2950_reg/NET0131 , \g2953_reg/NET0131 , \g2956_reg/NET0131 , \g2959_reg/NET0131 , \g2962_reg/NET0131 , \g2963_reg/NET0131 , \g2966_reg/NET0131 , \g2969_reg/NET0131 , \g2972_reg/NET0131 , \g2975_reg/NET0131 , \g2978_reg/NET0131 , \g2981_reg/NET0131 , \g2984_reg/NET0131 , \g2985_reg/NET0131 , \g2986_reg/NET0131 , \g2987_reg/NET0131 , \g298_reg/NET0131 , \g2990_reg/NET0131 , \g2991_reg/NET0131 , \g2992_reg/NET0131 , \g2993_reg/NET0131 , \g2997_reg/NET0131 , \g2998_reg/NET0131 , \g299_reg/NET0131 , \g3002_reg/NET0131 , \g3006_reg/NET0131 , \g3010_reg/NET0131 , \g3013_reg/NET0131 , \g3018_reg/NET0131 , \g3024_reg/NET0131 , \g3028_reg/NET0131 , \g3032_reg/NET0131 , \g3036_reg/NET0131 , \g3043_reg/NET0131 , \g3044_reg/NET0131 , \g3045_reg/NET0131 , \g3046_reg/NET0131 , \g3047_reg/NET0131 , \g3048_reg/NET0131 , \g3049_reg/NET0131 , \g3050_reg/NET0131 , \g3051_reg/NET0131 , \g3052_reg/NET0131 , \g3053_reg/NET0131 , \g3054_reg/NET0131 , \g3055_reg/NET0131 , \g3056_reg/NET0131 , \g3057_reg/NET0131 , \g3058_reg/NET0131 , \g3059_reg/NET0131 , \g305_reg/NET0131 , \g3060_reg/NET0131 , \g3061_reg/NET0131 , \g3062_reg/NET0131 , \g3063_reg/NET0131 , \g3064_reg/NET0131 , \g3065_reg/NET0131 , \g3066_reg/NET0131 , \g3067_reg/NET0131 , \g3068_reg/NET0131 , \g3069_reg/NET0131 , \g3070_reg/NET0131 , \g3071_reg/NET0131 , \g3072_reg/NET0131 , \g3073_reg/NET0131 , \g3074_reg/NET0131 , \g3075_reg/NET0131 , \g3076_reg/NET0131 , \g3077_reg/NET0131 , \g3078_reg/NET0131 , \g3079_reg/NET0131 , \g3080_reg/NET0131 , \g3083_reg/NET0131 , \g3097_reg/NET0131 , \g3110_reg/NET0131 , \g3114_reg/NET0131 , \g3120_reg/NET0131 , \g312_reg/NET0131 , \g3139_reg/NET0131 , \g313_reg/NET0131 , \g314_reg/NET0131 , \g315_reg/NET0131 , \g316_reg/NET0131 , \g317_reg/NET0131 , \g318_reg/NET0131 , \g319_reg/NET0131 , \g320_reg/NET0131 , \g321_reg/NET0131 , \g3229_pad , \g322_reg/NET0131 , \g3230_pad , \g3231_pad , \g3233_pad , \g3234_pad , \g323_reg/NET0131 , \g324_reg/NET0131 , \g343_reg/NET0131 , \g346_reg/NET0131 , \g349_reg/NET0131 , \g351_reg/NET0131 , \g353_reg/NET0131 , \g354_reg/NET0131 , \g358_reg/NET0131 , \g361_reg/NET0131 , \g364_reg/NET0131 , \g366_reg/NET0131 , \g368_reg/NET0131 , \g369_reg/NET0131 , \g373_reg/NET0131 , \g376_reg/NET0131 , \g379_reg/NET0131 , \g381_reg/NET0131 , \g383_reg/NET0131 , \g384_reg/NET0131 , \g388_reg/NET0131 , \g391_reg/NET0131 , \g394_reg/NET0131 , \g396_reg/NET0131 , \g398_reg/NET0131 , \g402_reg/NET0131 , \g403_reg/NET0131 , \g404_reg/NET0131 , \g408_reg/NET0131 , \g411_reg/NET0131 , \g414_reg/NET0131 , \g417_reg/NET0131 , \g420_reg/NET0131 , \g423_reg/NET0131 , \g426_reg/NET0131 , \g427_reg/NET0131 , \g428_reg/NET0131 , \g429_reg/NET0131 , \g432_reg/NET0131 , \g435_reg/NET0131 , \g438_reg/NET0131 , \g441_reg/NET0131 , \g444_reg/NET0131 , \g447_reg/NET0131 , \g448_reg/NET0131 , \g449_reg/NET0131 , \g451_reg/NET0131 , \g453_reg/NET0131 , \g464_reg/NET0131 , \g465_reg/NET0131 , \g468_reg/NET0131 , \g471_reg/NET0131 , \g477_reg/NET0131 , \g478_reg/NET0131 , \g479_reg/NET0131 , \g480_reg/NET0131 , \g484_reg/NET0131 , \g486_reg/NET0131 , \g487_reg/NET0131 , \g488_reg/NET0131 , \g489_reg/NET0131 , \g490_reg/NET0131 , \g493_reg/NET0131 , \g496_reg/NET0131 , \g499_reg/NET0131 , \g506_reg/NET0131 , \g507_reg/NET0131 , \g51_pad , \g524_reg/NET0131 , \g525_reg/NET0131 , \g529_reg/NET0131 , \g530_reg/NET0131 , \g531_reg/NET0131 , \g532_reg/NET0131 , \g533_reg/NET0131 , \g534_reg/NET0131 , \g536_reg/NET0131 , \g537_reg/NET0131 , \g5388_pad , \g538_reg/NET0131 , \g541_reg/NET0131 , \g542_reg/NET0131 , \g544_reg/NET0131 , \g548_reg/NET0131 , \g559_reg/NET0131 , \g563_pad , \g5657_pad , \g565_reg/NET0131 , \g567_reg/NET0131 , \g569_reg/NET0131 , \g571_reg/NET0131 , \g573_reg/NET0131 , \g575_reg/NET0131 , \g576_reg/NET0131 , \g577_reg/NET0131 , \g578_reg/NET0131 , \g579_reg/NET0131 , \g580_reg/NET0131 , \g581_reg/NET0131 , \g582_reg/NET0131 , \g583_reg/NET0131 , \g584_reg/NET0131 , \g585_reg/NET0131 , \g586_reg/NET0131 , \g587_reg/NET0131 , \g590_reg/NET0131 , \g593_reg/NET0131 , \g596_reg/NET0131 , \g599_reg/NET0131 , \g602_reg/NET0131 , \g605_reg/NET0131 , \g608_reg/NET0131 , \g611_reg/NET0131 , \g614_reg/NET0131 , \g617_reg/NET0131 , \g620_reg/NET0131 , \g698_reg/NET0131 , \g699_reg/NET0131 , \g700_reg/NET0131 , \g701_reg/NET0131 , \g702_reg/NET0131 , \g703_reg/NET0131 , \g704_reg/NET0131 , \g705_reg/NET0131 , \g706_reg/NET0131 , \g707_reg/NET0131 , \g708_reg/NET0131 , \g709_reg/NET0131 , \g710_reg/NET0131 , \g711_reg/NET0131 , \g712_reg/NET0131 , \g713_reg/NET0131 , \g714_reg/NET0131 , \g715_reg/NET0131 , \g716_reg/NET0131 , \g717_reg/NET0131 , \g718_reg/NET0131 , \g719_reg/NET0131 , \g720_reg/NET0131 , \g721_reg/NET0131 , \g722_reg/NET0131 , \g723_reg/NET0131 , \g724_reg/NET0131 , \g725_reg/NET0131 , \g726_reg/NET0131 , \g727_reg/NET0131 , \g728_reg/NET0131 , \g729_reg/NET0131 , \g730_reg/NET0131 , \g731_reg/NET0131 , \g732_reg/NET0131 , \g733_reg/NET0131 , \g734_reg/NET0131 , \g735_reg/NET0131 , \g736_reg/NET0131 , \g737_reg/NET0131 , \g738_reg/NET0131 , \g739_reg/NET0131 , \g785_reg/NET0131 , \g789_reg/NET0131 , \g793_reg/NET0131 , \g7961_pad , \g797_reg/NET0131 , \g801_reg/NET0131 , \g805_reg/NET0131 , \g809_reg/NET0131 , \g813_reg/NET0131 , \g817_reg/NET0131 , \g818_reg/NET0131 , \g819_reg/NET0131 , \g820_reg/NET0131 , \g821_reg/NET0131 , \g822_reg/NET0131 , \g8259_pad , \g8260_pad , \g8261_pad , \g8262_pad , \g8263_pad , \g8264_pad , \g8265_pad , \g8266_pad , \g8268_pad , \g8269_pad , \g8270_pad , \g8271_pad , \g8272_pad , \g8273_pad , \g8274_pad , \g8275_pad , \g829_reg/NET0131 , \g830_reg/NET0131 , \g831_reg/NET0131 , \g832_reg/NET0131 , \g833_reg/NET0131 , \g834_reg/NET0131 , \g835_reg/NET0131 , \g836_reg/NET0131 , \g837_reg/NET0131 , \g838_reg/NET0131 , \g839_reg/NET0131 , \g840_reg/NET0131 , \g841_reg/NET0131 , \g842_reg/NET0131 , \g843_reg/NET0131 , \g844_reg/NET0131 , \g845_reg/NET0131 , \g846_reg/NET0131 , \g847_reg/NET0131 , \g848_reg/NET0131 , \g849_reg/NET0131 , \g850_reg/NET0131 , \g851_reg/NET0131 , \g852_reg/NET0131 , \g856_reg/NET0131 , \g857_reg/NET0131 , \g858_reg/NET0131 , \g859_reg/NET0131 , \g860_reg/NET0131 , \g861_reg/NET0131 , \g862_reg/NET0131 , \g863_reg/NET0131 , \g864_reg/NET0131 , \g865_reg/NET0131 , \g866_reg/NET0131 , \g867_reg/NET0131 , \g873_reg/NET0131 , \g876_reg/NET0131 , \g879_reg/NET0131 , \g882_reg/NET0131 , \g885_reg/NET0131 , \g888_reg/NET0131 , \g891_reg/NET0131 , \g894_reg/NET0131 , \g897_reg/NET0131 , \g900_reg/NET0131 , \g903_reg/NET0131 , \g906_reg/NET0131 , \g909_reg/NET0131 , \g912_reg/NET0131 , \g915_reg/NET0131 , \g918_reg/NET0131 , \g921_reg/NET0131 , \g924_reg/NET0131 , \g927_reg/NET0131 , \g930_reg/NET0131 , \g933_reg/NET0131 , \g936_reg/NET0131 , \g939_reg/NET0131 , \g942_reg/NET0131 , \g945_reg/NET0131 , \g948_reg/NET0131 , \g951_reg/NET0131 , \g954_reg/NET0131 , \g957_reg/NET0131 , \g960_reg/NET0131 , \g966_reg/NET0131 , \g968_reg/NET0131 , \g970_reg/NET0131 , \g972_reg/NET0131 , \g974_reg/NET0131 , \g976_reg/NET0131 , \g978_reg/NET0131 , \g97_reg/NET0131 , \g985_reg/NET0131 , \g986_reg/NET0131 , \g992_reg/NET0131 , \g999_reg/NET0131 , \_al_n0 , \_al_n1 , \g101_reg/P0001 , \g105_reg/P0001 , \g109_reg/P0001 , \g1138_reg/P0001 , \g113_reg/P0001 , \g1140_reg/P0001 , \g117_reg/P0001 , \g121_reg/P0001 , \g125_reg/P0001 , \g1471_reg/P0001 , \g1476_reg/P0001 , \g1481_reg/P0001 , \g1486_reg/P0001 , \g1491_reg/P0001 , \g1496_reg/P0001 , \g1501_reg/P0001 , \g1506_reg/P0001 , \g16496_pad , \g1660_reg/P0001 , \g1662_reg/P0001 , \g1664_reg/P0001 , \g1666_reg/P0001 , \g1668_reg/P0001 , \g1670_reg/P0001 , \g1672_reg/P0001 , \g18/_0_ , \g1832_reg/P0001 , \g1834_reg/P0001 , \g2165_reg/P0001 , \g2170_reg/P0001 , \g2175_reg/P0001 , \g2180_reg/P0001 , \g2185_reg/P0001 , \g2190_reg/P0001 , \g2195_reg/P0001 , \g2200_reg/P0001 , \g2354_reg/P0001 , \g2356_reg/P0001 , \g2358_reg/P0001 , \g2360_reg/P0001 , \g2362_reg/P0001 , \g2364_reg/P0001 , \g2366_reg/P0001 , \g2526_reg/P0001 , \g2528_reg/P0001 , \g25489_pad , \g279_reg/P0001 , \g281_reg/P0001 , \g283_reg/P0001 , \g285_reg/P0001 , \g2879_reg/NET0131_syn_2 , \g287_reg/P0001 , \g289_reg/P0001 , \g291_reg/P0001 , \g451_reg/P0001 , \g453_reg/P0001 , \g59421/_3_ , \g59425/_1_ , \g59435/_0_ , \g59436/_0_ , \g59441/_3_ , \g59442/_0_ , \g59445/_0_ , \g59453/_0_ , \g59462/_3_ , \g59466/_3_ , \g59467/_3_ , \g59468/_3_ , \g59469/_3_ , \g59470/_3_ , \g59471/_3_ , \g59472/_3_ , \g59473/_3_ , \g59489/_0_ , \g59498/_0_ , \g59499/_0_ , \g59500/_0_ , \g59502/_2_ , \g59503/_0_ , \g59505/_2_ , \g59507/_0_ , \g59508/_0_ , \g59533/_3_ , \g59534/_3_ , \g59535/_3_ , \g59536/_3_ , \g59537/_3_ , \g59538/_3_ , \g59539/_3_ , \g59540/_3_ , \g59548/_0_ , \g59550/_0_ , \g59551/_0_ , \g59552/_0_ , \g59554/_0_ , \g59555/_0_ , \g59556/_0_ , \g59557/_0_ , \g59558/_0_ , \g59559/_0_ , \g59560/_0_ , \g59561/_0_ , \g59639/_0_ , \g59694/_2_ , \g59695/_0_ , \g59697/_2_ , \g59698/_0_ , \g59699/_0_ , \g59700/_0_ , \g59705/_0_ , \g59706/_0_ , \g59707/_0_ , \g59708/_0_ , \g59709/_0_ , \g59710/_0_ , \g59711/_0_ , \g59712/_0_ , \g59713/_0_ , \g59714/_0_ , \g59715/_0_ , \g59716/_0_ , \g59717/_0_ , \g59718/_0_ , \g59719/_0_ , \g59720/_0_ , \g59721/_0_ , \g59722/_0_ , \g59723/_0_ , \g59724/_0_ , \g59725/_0_ , \g59726/_0_ , \g59727/_0_ , \g59728/_0_ , \g59729/_0_ , \g59730/_0_ , \g59731/_0_ , \g59732/_0_ , \g59733/_0_ , \g59734/_0_ , \g59735/_0_ , \g59736/_0_ , \g59737/_0_ , \g59738/_0_ , \g59739/_0_ , \g59740/_0_ , \g59741/_0_ , \g59742/_0_ , \g59743/_0_ , \g59744/_0_ , \g59745/_0_ , \g59747/_0_ , \g59748/_0_ , \g59749/_0_ , \g59750/_0_ , \g59751/_0_ , \g59752/_0_ , \g59753/_0_ , \g59754/_0_ , \g59755/_0_ , \g59756/_0_ , \g59757/_0_ , \g59758/_0_ , \g59759/_0_ , \g59760/_0_ , \g59761/_0_ , \g59762/_0_ , \g59763/_0_ , \g59764/_0_ , \g59765/_0_ , \g59766/_0_ , \g59915/_0_ , \g59952/_2_ , \g60046/_0_ , \g60048/_0_ , \g60049/_0_ , \g60051/_0_ , \g60063/_0_ , \g60103/_0_ , \g60104/_0_ , \g60105/_0_ , \g60107/_2_ , \g60108/_0_ , \g60109/_0_ , \g60110/_0_ , \g60112/_2_ , \g60119/_0_ , \g60120/_0_ , \g60121/_0_ , \g60122/_0_ , \g60123/_0_ , \g60124/_0_ , \g60126/_0_ , \g60127/_0_ , \g60128/_0_ , \g60129/_0_ , \g60130/_0_ , \g60135/_0_ , \g60136/_0_ , \g60137/_0_ , \g60138/_0_ , \g60139/_0_ , \g60143/_3_ , \g60144/_0_ , \g60145/_0_ , \g60339/_0_ , \g60404/_0_ , \g60427/_0_ , \g60428/_0_ , \g60429/_0_ , \g60434/_0_ , \g60435/_0_ , \g60437/_0_ , \g60438/_0_ , \g60439/_0_ , \g60440/_0_ , \g60441/_0_ , \g60448/_0_ , \g60451/_0_ , \g60452/_0_ , \g60453/_0_ , \g60459/_0_ , \g60460/_0_ , \g60523/_0_ , \g60534/_0_ , \g60535/_0_ , \g60536/_0_ , \g60585/_0_ , \g60586/_0_ , \g60587/_0_ , \g60588/_0_ , \g60591/_0_ , \g60592/_0_ , \g60599/_0_ , \g60601/_0_ , \g60602/_0_ , \g60603/_0_ , \g60604/_0_ , \g60605/_0_ , \g60606/_0_ , \g60607/_0_ , \g60608/_0_ , \g60609/_0_ , \g60613/_0_ , \g60614/_0_ , \g60615/_0_ , \g60694/_0_ , \g60708/_0_ , \g60709/_0_ , \g60710/_0_ , \g60785/_0_ , \g60787/_0_ , \g60788/_0_ , \g60799/_0_ , \g60801/_0_ , \g60802/_0_ , \g60803/_1__syn_2 , \g60805/_1__syn_2 , \g60806/_1__syn_2 , \g60808/_0_ , \g60810/_0_ , \g60811/_0_ , \g60825/_3_ , \g60896/_0_ , \g60980/_0_ , \g60981/_0_ , \g60985/_0_ , \g60986/_0_ , \g61012/_0_ , \g61013/_0_ , \g61015/_0_ , \g61017/_0_ , \g61122/_0_ , \g61123/_0_ , \g61124/_0_ , \g61125/_0_ , \g61222/_0_ , \g61223/_0_ , \g61224/_0_ , \g61225/_0_ , \g61228/_0_ , \g61229/_0_ , \g61230/_0_ , \g61231/_0_ , \g61281/_0_ , \g61293/_1_ , \g61307/_0__syn_2 , \g61309/_0__syn_2 , \g61310/_0__syn_2 , \g61311/_1_ , \g61312/_1_ , \g61313/_1_ , \g61324/_1_ , \g61325/_1_ , \g61326/_1_ , \g61328/_1_ , \g61329/_1_ , \g61330/_1_ , \g61332/_1_ , \g61333/_1_ , \g61334/_1_ , \g61335/_1_ , \g61336/_0_ , \g61338/_0_ , \g61339/_0_ , \g61340/_0_ , \g61377/_1_ , \g61378/_1_ , \g61379/_1_ , \g61388/_1_ , \g61391/_0_ , \g61394/_1_ , \g61395/_1_ , \g61396/_1_ , \g61398/_1_ , \g61399/_1_ , \g61421/_1_ , \g61422/_1_ , \g61423/_1_ , \g61524/_0_ , \g61525/_0_ , \g61526/_0_ , \g61527/_0_ , \g61528/_0_ , \g61529/_0_ , \g61530/_0_ , \g61531/_0_ , \g61532/_0_ , \g61533/_0_ , \g61534/_0_ , \g61535/_0_ , \g61536/_0_ , \g61537/_0_ , \g61538/_0_ , \g61539/_0_ , \g61540/_0_ , \g61541/_0_ , \g61542/_0_ , \g61543/_0_ , \g61544/_0_ , \g61545/_0_ , \g61546/_0_ , \g61547/_0_ , \g61548/_0_ , \g61549/_0_ , \g61550/_0_ , \g61551/_0_ , \g61552/_0_ , \g61553/_0_ , \g61554/_0_ , \g61555/_0_ , \g61556/_0_ , \g61557/_0_ , \g61558/_0_ , \g61559/_0_ , \g61560/_0_ , \g61561/_0_ , \g61562/_0_ , \g61563/_0_ , \g61564/_0_ , \g61565/_0_ , \g61566/_0_ , \g61620/_0_ , \g61621/_0_ , \g61622/_0_ , \g61623/_0_ , \g61753/_0_ , \g61764/_0_ , \g61786/_0_ , \g61795/_0_ , \g61801/_0_ , \g61803/_0_ , \g61808/_0_ , \g61848/_0_ , \g61850/_0_ , \g61851/_0_ , \g62097/_0_ , \g62102/_0_ , \g62115/_0_ , \g62119/_0_ , \g62130/_1_ , \g62131/_0_ , \g62132/_0_ , \g62139/_1_ , \g62140/_1_ , \g62141/_1_ , \g62144/_0_ , \g62145/_0_ , \g62146/_0_ , \g62147/_0_ , \g62150/_0_ , \g62151/_1_ , \g62152/_0_ , \g62153/_1_ , \g62156/_1_ , \g62157/_0_ , \g62159/_0_ , \g62161/_0_ , \g62187/_1_ , \g62190/_1_ , \g62191/_1_ , \g62192/_1_ , \g62194/_1_ , \g62195/_1_ , \g62196/_1_ , \g62203/_0_ , \g62204/_1_ , \g62207/_0__syn_2 , \g62208/_1_ , \g62209/_1_ , \g62210/_1_ , \g62211/_1_ , \g62212/_1_ , \g62217/_0_ , \g62286/_0_ , \g62287/_0_ , \g62288/_0_ , \g62289/_0_ , \g62290/_0_ , \g62291/_0_ , \g62292/_0_ , \g62435/_0_ , \g62436/_0_ , \g62439/_0_ , \g62456/_0_ , \g62486/_1_ , \g62492/_1_ , \g62494/_0_ , \g62495/_1_ , \g62497/_0_ , \g62537/_0_ , \g62544/_0_ , \g62546/_0_ , \g62547/_0_ , \g62549/_3_ , \g62552/_0_ , \g62554/_0_ , \g62555/_0_ , \g62556/_0_ , \g62558/_0_ , \g62559/_0_ , \g62561/_0_ , \g62562/_0_ , \g62566/_0_ , \g62567/_0_ , \g62568/_0_ , \g62569/_0_ , \g62570/_0_ , \g62571/_0_ , \g62572/_0_ , \g62573/_0_ , \g62574/_0_ , \g62575/_0_ , \g62576/_0_ , \g62577/_0_ , \g62578/_0_ , \g62579/_0_ , \g62580/_0_ , \g62581/_0_ , \g62582/_0_ , \g62583/_0_ , \g62584/_0_ , \g62585/_0_ , \g62586/_0_ , \g62587/_0_ , \g62588/_0_ , \g62589/_0_ , \g62590/_0_ , \g62591/_0_ , \g62592/_0_ , \g62593/_0_ , \g62594/_0_ , \g62595/_0_ , \g62596/_0_ , \g62597/_0_ , \g62602/_0_ , \g62607/_0_ , \g62608/_0_ , \g62609/_0_ , \g62619/_0_ , \g62620/_0_ , \g62621/_0_ , \g62622/_0_ , \g62623/_0_ , \g62624/_0_ , \g62626/_0_ , \g62627/_0_ , \g62628/_0_ , \g62629/_0_ , \g62630/_0_ , \g62631/_0_ , \g62632/_0_ , \g62633/_0_ , \g62634/_0_ , \g62635/_0_ , \g62636/_0_ , \g62637/_0_ , \g62638/_0_ , \g62639/_0_ , \g62640/_0_ , \g62641/_0_ , \g62642/_0_ , \g62643/_0_ , \g62644/_0_ , \g62645/_0_ , \g62646/_0_ , \g62647/_0_ , \g62648/_0_ , \g62649/_0_ , \g62650/_0_ , \g62651/_0_ , \g62652/_0_ , \g62653/_0_ , \g62654/_0_ , \g62655/_0_ , \g62656/_0_ , \g62657/_0_ , \g62658/_0_ , \g62659/_0_ , \g62660/_0_ , \g62661/_0_ , \g62674/_0_ , \g62682/_0_ , \g62683/_0_ , \g62689/_0_ , \g62690/_0_ , \g62691/_0_ , \g62694/_0_ , \g62695/_0_ , \g62696/_0_ , \g62698/_0_ , \g62699/_0_ , \g62700/_0_ , \g62723/_0_ , \g62724/_0_ , \g62725/_0_ , \g62726/_0_ , \g62727/_0_ , \g62728/_0_ , \g62735/_0_ , \g62736/_0_ , \g62737/_0_ , \g62738/_0_ , \g62739/_0_ , \g62740/_0_ , \g62754/_0_ , \g62762/_0_ , \g62763/_0_ , \g62764/_0_ , \g62780/_0_ , \g62781/_0_ , \g62785/_0_ , \g62786/_0_ , \g62787/_0_ , \g62791/_0_ , \g62792/_0_ , \g62794/_0_ , \g62804/_0_ , \g62806/_0_ , \g62807/_0_ , \g62811/_0_ , \g62968/_0_ , \g63005/_0_ , \g63041/_0_ , \g63116/_0_ , \g63157/_0_ , \g63164/_0_ , \g63170/_0_ , \g63189/_0_ , \g63202/_0_ , \g63206/_0_ , \g63207/_0_ , \g63265/_0_ , \g63266/_0_ , \g63269/_0_ , \g63271/_0_ , \g63272/_0_ , \g63273/_0_ , \g63274/_0_ , \g63275/_0_ , \g63276/_0_ , \g63277/_0_ , \g63278/_0_ , \g63280/_0_ , \g63281/_0_ , \g63282/_0_ , \g63283/_0_ , \g63284/_0_ , \g63285/_0_ , \g63286/_0_ , \g63287/_0_ , \g63288/_0_ , \g63289/_0_ , \g63290/_0_ , \g63292/_0_ , \g63293/_0_ , \g63294/_0_ , \g63295/_0_ , \g63296/_0_ , \g63297/_0_ , \g63298/_0_ , \g63299/_0_ , \g63302/_0_ , \g63303/_0_ , \g63304/_0_ , \g63305/_0_ , \g63306/_0_ , \g63307/_0_ , \g63308/_0_ , \g63309/_0_ , \g63310/_0_ , \g63311/_0_ , \g63312/_0_ , \g63313/_0_ , \g63314/_0_ , \g63315/_0_ , \g63316/_0_ , \g63317/_0_ , \g63318/_0_ , \g63319/_0_ , \g63320/_0_ , \g63321/_0_ , \g63322/_0_ , \g63323/_0_ , \g63324/_0_ , \g63325/_0_ , \g63326/_0_ , \g63327/_0_ , \g63328/_0_ , \g63329/_0_ , \g63330/_0_ , \g63331/_0_ , \g63339/_0_ , \g63505/_0_ , \g63525/_0_ , \g63543/_1_ , \g63602/_0_ , \g63653/_0_ , \g63663/_1_ , \g63677/_0_ , \g63694/_0_ , \g63729/_0_ , \g63766/_0_ , \g63771/_1_ , \g63773/_1_ , \g63784/_1_ , \g63964/_0_ , \g63965/_0_ , \g63966/_0_ , \g63967/_0_ , \g64257/_1_ , \g64266/_0_ , \g64275/_0_ , \g64400/_0_ , \g64416/_0_ , \g64470/_3_ , \g64473/_0_ , \g64474/_0_ , \g64475/_0_ , \g64479/_0_ , \g64480/_0_ , \g64481/_0_ , \g64483/_0_ , \g64484/_0_ , \g64485/_0_ , \g64486/_0_ , \g64493/_0_ , \g64494/_0_ , \g64495/_0_ , \g64496/_0_ , \g64505/_3_ , \g64507/_0_ , \g64508/_0_ , \g64510/_0_ , \g64511/_0_ , \g64544/_0_ , \g64545/_0_ , \g64546/_0_ , \g64639/_0_ , \g64641/_0_ , \g64642/_0_ , \g64645/_0_ , \g64650/_0_ , \g64737/_0_ , \g64738/_0_ , \g65066/_0_ , \g65070/_0_ , \g65090/_0_ , \g65102/_0_ , \g65102/_3_ , \g65126/_3_ , \g65147/_3_ , \g65163/_0_ , \g65176/_3_ , \g65178/_0_ , \g65182/_0_ , \g65190/_1_ , \g65191/_0_ , \g65196/_0_ , \g65268/_0_ , \g65275/_0_ , \g65290/_0_ , \g65290/_3_ , \g65291/_0_ , \g65292/_0_ , \g65298/_0_ , \g65298/_3_ , \g65314/_0_ , \g65314/_3_ , \g65319/_3_ , \g65335/_0_ , \g65342/_0_ , \g65348/_0_ , \g65422/_0_ , \g65465/_1_ , \g65469/_1_ , \g65478/_1_ , \g65507/_0_ , \g65548/_0_ , \g65699/_1_ , \g65713/_1_ , \g65835/_0_ , \g65860/_0_ , \g65863/_0_ , \g66094/_1_ , \g66102/_0_ , \g66107/_0_ , \g66130/_3_ , \g66131/_3_ , \g66228/_1_ , \g66348/_1_ , \g66543/_0_ , \g66549/_1_ , \g66640/_3_ , \g66641/_3_ , \g66950/_1_ , \g67111/_0_ , \g67219/_0_ , \g67263/_0_ , \g67909/_1_ , \g68049/_0_ , \g68220/_0_ , \g68413/_0_ , \g68511/_0_ , \g68536/_0_ , \g68543/_1_ , \g68554/_0_ , \g68559/_0_ , \g70915/_0_ , \g71108/_1_ , \g71115/_2_ , \g71244_dup/_0_ , \g71368/_0_ , \g71581/_0_ , \g71720/_0_ , \g785_reg/P0001 , \g789_reg/P0001 , \g797_reg/P0001 , \g809_reg/P0001 , \g813_reg/P0001 , \g966_reg/P0001 , \g968_reg/P0001 , \g970_reg/P0001 , \g972_reg/P0001 , \g974_reg/P0001 , \g976_reg/P0001 , \g978_reg/P0001 );
	input \g1000_reg/NET0131  ;
	input \g1001_reg/NET0131  ;
	input \g1002_reg/NET0131  ;
	input \g1003_reg/NET0131  ;
	input \g1004_reg/NET0131  ;
	input \g1005_reg/NET0131  ;
	input \g1006_reg/NET0131  ;
	input \g1007_reg/NET0131  ;
	input \g1008_reg/NET0131  ;
	input \g1009_reg/NET0131  ;
	input \g1010_reg/NET0131  ;
	input \g1011_reg/NET0131  ;
	input \g1018_reg/NET0131  ;
	input \g101_reg/NET0131  ;
	input \g1024_reg/NET0131  ;
	input \g1030_reg/NET0131  ;
	input \g1033_reg/NET0131  ;
	input \g1036_reg/NET0131  ;
	input \g1038_reg/NET0131  ;
	input \g1040_reg/NET0131  ;
	input \g1041_reg/NET0131  ;
	input \g1045_reg/NET0131  ;
	input \g1048_reg/NET0131  ;
	input \g1051_reg/NET0131  ;
	input \g1053_reg/NET0131  ;
	input \g1055_reg/NET0131  ;
	input \g1056_reg/NET0131  ;
	input \g105_reg/NET0131  ;
	input \g1060_reg/NET0131  ;
	input \g1063_reg/NET0131  ;
	input \g1066_reg/NET0131  ;
	input \g1068_reg/NET0131  ;
	input \g1070_reg/NET0131  ;
	input \g1071_reg/NET0131  ;
	input \g1075_reg/NET0131  ;
	input \g1078_reg/NET0131  ;
	input \g1081_reg/NET0131  ;
	input \g1083_reg/NET0131  ;
	input \g1085_reg/NET0131  ;
	input \g1088_reg/NET0131  ;
	input \g1089_reg/NET0131  ;
	input \g1090_reg/NET0131  ;
	input \g1091_reg/NET0131  ;
	input \g1092_reg/NET0131  ;
	input \g1095_reg/NET0131  ;
	input \g1098_reg/NET0131  ;
	input \g109_reg/NET0131  ;
	input \g1101_reg/NET0131  ;
	input \g1104_reg/NET0131  ;
	input \g1107_reg/NET0131  ;
	input \g1110_reg/NET0131  ;
	input \g1113_reg/NET0131  ;
	input \g1114_reg/NET0131  ;
	input \g1115_reg/NET0131  ;
	input \g1116_reg/NET0131  ;
	input \g1119_reg/NET0131  ;
	input \g1122_reg/NET0131  ;
	input \g1125_reg/NET0131  ;
	input \g1128_reg/NET0131  ;
	input \g1131_reg/NET0131  ;
	input \g1134_reg/NET0131  ;
	input \g1135_reg/NET0131  ;
	input \g1136_reg/NET0131  ;
	input \g1138_reg/NET0131  ;
	input \g113_reg/NET0131  ;
	input \g1140_reg/NET0131  ;
	input \g1151_reg/NET0131  ;
	input \g1164_reg/NET0131  ;
	input \g1165_reg/NET0131  ;
	input \g1166_reg/NET0131  ;
	input \g1167_reg/NET0131  ;
	input \g1171_reg/NET0131  ;
	input \g1173_reg/NET0131  ;
	input \g1174_reg/NET0131  ;
	input \g1175_reg/NET0131  ;
	input \g1176_reg/NET0131  ;
	input \g1177_reg/NET0131  ;
	input \g117_reg/NET0131  ;
	input \g1180_reg/NET0131  ;
	input \g1183_reg/NET0131  ;
	input \g1186_reg/NET0131  ;
	input \g1192_reg/NET0131  ;
	input \g1193_reg/NET0131  ;
	input \g1196_reg/NET0131  ;
	input \g1210_reg/NET0131  ;
	input \g1211_reg/NET0131  ;
	input \g1215_reg/NET0131  ;
	input \g1216_reg/NET0131  ;
	input \g1217_reg/NET0131  ;
	input \g1218_reg/NET0131  ;
	input \g1219_reg/NET0131  ;
	input \g121_reg/NET0131  ;
	input \g1220_reg/NET0131  ;
	input \g1222_reg/NET0131  ;
	input \g1223_reg/NET0131  ;
	input \g1224_reg/NET0131  ;
	input \g1227_reg/NET0131  ;
	input \g1228_reg/NET0131  ;
	input \g1230_reg/NET0131  ;
	input \g1234_reg/NET0131  ;
	input \g1240_reg/NET0131  ;
	input \g1243_reg/NET0131  ;
	input \g1245_reg/NET0131  ;
	input \g1249_pad  ;
	input \g1251_reg/NET0131  ;
	input \g1253_reg/NET0131  ;
	input \g1255_reg/NET0131  ;
	input \g1257_reg/NET0131  ;
	input \g1259_reg/NET0131  ;
	input \g125_reg/NET0131  ;
	input \g1261_reg/NET0131  ;
	input \g1262_reg/NET0131  ;
	input \g1263_reg/NET0131  ;
	input \g1264_reg/NET0131  ;
	input \g1265_reg/NET0131  ;
	input \g1266_reg/NET0131  ;
	input \g1267_reg/NET0131  ;
	input \g1268_reg/NET0131  ;
	input \g1269_reg/NET0131  ;
	input \g1270_reg/NET0131  ;
	input \g1271_reg/NET0131  ;
	input \g1272_reg/NET0131  ;
	input \g1273_reg/NET0131  ;
	input \g1276_reg/NET0131  ;
	input \g1279_reg/NET0131  ;
	input \g1282_reg/NET0131  ;
	input \g1285_reg/NET0131  ;
	input \g1288_reg/NET0131  ;
	input \g1291_reg/NET0131  ;
	input \g1294_reg/NET0131  ;
	input \g1297_reg/NET0131  ;
	input \g129_reg/NET0131  ;
	input \g1300_reg/NET0131  ;
	input \g1303_reg/NET0131  ;
	input \g1306_reg/NET0131  ;
	input \g130_reg/NET0131  ;
	input \g1316_reg/NET0131  ;
	input \g1319_reg/NET0131  ;
	input \g131_reg/NET0131  ;
	input \g1326_reg/NET0131  ;
	input \g132_reg/NET0131  ;
	input \g1332_reg/NET0131  ;
	input \g1339_reg/NET0131  ;
	input \g133_reg/NET0131  ;
	input \g1345_reg/NET0131  ;
	input \g1346_reg/NET0131  ;
	input \g134_reg/NET0131  ;
	input \g1352_reg/NET0131  ;
	input \g1358_reg/NET0131  ;
	input \g1365_reg/NET0131  ;
	input \g1372_reg/NET0131  ;
	input \g1378_reg/NET0131  ;
	input \g1384_reg/NET0131  ;
	input \g1385_reg/NET0131  ;
	input \g1386_reg/NET0131  ;
	input \g1387_reg/NET0131  ;
	input \g1388_reg/NET0131  ;
	input \g1389_reg/NET0131  ;
	input \g1390_reg/NET0131  ;
	input \g1391_reg/NET0131  ;
	input \g1392_reg/NET0131  ;
	input \g1393_reg/NET0131  ;
	input \g1394_reg/NET0131  ;
	input \g1395_reg/NET0131  ;
	input \g1396_reg/NET0131  ;
	input \g1397_reg/NET0131  ;
	input \g1398_reg/NET0131  ;
	input \g1399_reg/NET0131  ;
	input \g1400_reg/NET0131  ;
	input \g1401_reg/NET0131  ;
	input \g1402_reg/NET0131  ;
	input \g1403_reg/NET0131  ;
	input \g1404_reg/NET0131  ;
	input \g1405_reg/NET0131  ;
	input \g1406_reg/NET0131  ;
	input \g1407_reg/NET0131  ;
	input \g1408_reg/NET0131  ;
	input \g1409_reg/NET0131  ;
	input \g1410_reg/NET0131  ;
	input \g1411_reg/NET0131  ;
	input \g1412_reg/NET0131  ;
	input \g1413_reg/NET0131  ;
	input \g1414_reg/NET0131  ;
	input \g1415_reg/NET0131  ;
	input \g1416_reg/NET0131  ;
	input \g1417_reg/NET0131  ;
	input \g1418_reg/NET0131  ;
	input \g1419_reg/NET0131  ;
	input \g141_reg/NET0131  ;
	input \g1420_reg/NET0131  ;
	input \g1421_reg/NET0131  ;
	input \g1422_reg/NET0131  ;
	input \g1423_reg/NET0131  ;
	input \g1424_reg/NET0131  ;
	input \g1425_reg/NET0131  ;
	input \g1426_reg/NET0131  ;
	input \g142_reg/NET0131  ;
	input \g1430_reg/NET0131  ;
	input \g1435_reg/NET0131  ;
	input \g1439_reg/NET0131  ;
	input \g143_reg/NET0131  ;
	input \g1444_reg/NET0131  ;
	input \g1448_reg/NET0131  ;
	input \g144_reg/NET0131  ;
	input \g1453_reg/NET0131  ;
	input \g1457_reg/NET0131  ;
	input \g145_reg/NET0131  ;
	input \g1462_reg/NET0131  ;
	input \g1466_reg/NET0131  ;
	input \g146_reg/NET0131  ;
	input \g1471_reg/NET0131  ;
	input \g1476_reg/NET0131  ;
	input \g147_reg/NET0131  ;
	input \g1481_reg/NET0131  ;
	input \g1486_reg/NET0131  ;
	input \g148_reg/NET0131  ;
	input \g1491_reg/NET0131  ;
	input \g1496_reg/NET0131  ;
	input \g149_reg/NET0131  ;
	input \g1501_reg/NET0131  ;
	input \g1506_reg/NET0131  ;
	input \g150_reg/NET0131  ;
	input \g1511_reg/NET0131  ;
	input \g1512_reg/NET0131  ;
	input \g1513_reg/NET0131  ;
	input \g1514_reg/NET0131  ;
	input \g1515_reg/NET0131  ;
	input \g1516_reg/NET0131  ;
	input \g151_reg/NET0131  ;
	input \g1523_reg/NET0131  ;
	input \g1524_reg/NET0131  ;
	input \g1525_reg/NET0131  ;
	input \g1526_reg/NET0131  ;
	input \g1527_reg/NET0131  ;
	input \g1528_reg/NET0131  ;
	input \g1529_reg/NET0131  ;
	input \g152_reg/NET0131  ;
	input \g1530_reg/NET0131  ;
	input \g1531_reg/NET0131  ;
	input \g1532_reg/NET0131  ;
	input \g1533_reg/NET0131  ;
	input \g1534_reg/NET0131  ;
	input \g1535_reg/NET0131  ;
	input \g1536_reg/NET0131  ;
	input \g1537_reg/NET0131  ;
	input \g1538_reg/NET0131  ;
	input \g1539_reg/NET0131  ;
	input \g153_reg/NET0131  ;
	input \g1540_reg/NET0131  ;
	input \g1541_reg/NET0131  ;
	input \g1542_reg/NET0131  ;
	input \g1543_reg/NET0131  ;
	input \g1544_reg/NET0131  ;
	input \g1545_reg/NET0131  ;
	input \g1546_reg/NET0131  ;
	input \g154_reg/NET0131  ;
	input \g1550_reg/NET0131  ;
	input \g1551_reg/NET0131  ;
	input \g1552_reg/NET0131  ;
	input \g1553_reg/NET0131  ;
	input \g1554_reg/NET0131  ;
	input \g1555_reg/NET0131  ;
	input \g1556_reg/NET0131  ;
	input \g1557_reg/NET0131  ;
	input \g1558_reg/NET0131  ;
	input \g1559_reg/NET0131  ;
	input \g155_reg/NET0131  ;
	input \g1560_reg/NET0131  ;
	input \g1561_reg/NET0131  ;
	input \g1563_reg/NET0131  ;
	input \g1567_reg/NET0131  ;
	input \g156_reg/NET0131  ;
	input \g1570_reg/NET0131  ;
	input \g1573_reg/NET0131  ;
	input \g1576_reg/NET0131  ;
	input \g1579_reg/NET0131  ;
	input \g157_reg/NET0131  ;
	input \g1582_reg/NET0131  ;
	input \g1585_reg/NET0131  ;
	input \g1588_reg/NET0131  ;
	input \g158_reg/NET0131  ;
	input \g1591_reg/NET0131  ;
	input \g1594_reg/NET0131  ;
	input \g1597_reg/NET0131  ;
	input \g159_reg/NET0131  ;
	input \g1600_reg/NET0131  ;
	input \g1603_reg/NET0131  ;
	input \g1606_reg/NET0131  ;
	input \g1609_reg/NET0131  ;
	input \g160_reg/NET0131  ;
	input \g1612_reg/NET0131  ;
	input \g1615_reg/NET0131  ;
	input \g1618_reg/NET0131  ;
	input \g161_reg/NET0131  ;
	input \g1621_reg/NET0131  ;
	input \g1624_reg/NET0131  ;
	input \g1627_reg/NET0131  ;
	input \g16297_pad  ;
	input \g162_reg/NET0131  ;
	input \g1630_reg/NET0131  ;
	input \g1633_reg/NET0131  ;
	input \g16355_pad  ;
	input \g1636_reg/NET0131  ;
	input \g16399_pad  ;
	input \g1639_reg/NET0131  ;
	input \g163_reg/NET0131  ;
	input \g1642_reg/NET0131  ;
	input \g16437_pad  ;
	input \g1645_reg/NET0131  ;
	input \g1648_reg/NET0131  ;
	input \g164_reg/NET0131  ;
	input \g1651_reg/NET0131  ;
	input \g1654_reg/NET0131  ;
	input \g1660_reg/NET0131  ;
	input \g1662_reg/NET0131  ;
	input \g1664_reg/NET0131  ;
	input \g1666_reg/NET0131  ;
	input \g1668_reg/NET0131  ;
	input \g1670_reg/NET0131  ;
	input \g1672_reg/NET0131  ;
	input \g1679_reg/NET0131  ;
	input \g1680_reg/NET0131  ;
	input \g1686_reg/NET0131  ;
	input \g168_reg/NET0131  ;
	input \g1693_reg/NET0131  ;
	input \g1694_reg/NET0131  ;
	input \g1695_reg/NET0131  ;
	input \g1696_reg/NET0131  ;
	input \g1697_reg/NET0131  ;
	input \g1698_reg/NET0131  ;
	input \g1699_reg/NET0131  ;
	input \g169_reg/NET0131  ;
	input \g1700_reg/NET0131  ;
	input \g1701_reg/NET0131  ;
	input \g1702_reg/NET0131  ;
	input \g1703_reg/NET0131  ;
	input \g1704_reg/NET0131  ;
	input \g1705_reg/NET0131  ;
	input \g170_reg/NET0131  ;
	input \g171_reg/NET0131  ;
	input \g1724_reg/NET0131  ;
	input \g1727_reg/NET0131  ;
	input \g172_reg/NET0131  ;
	input \g1730_reg/NET0131  ;
	input \g1732_reg/NET0131  ;
	input \g1734_reg/NET0131  ;
	input \g1735_reg/NET0131  ;
	input \g1739_reg/NET0131  ;
	input \g173_reg/NET0131  ;
	input \g1742_reg/NET0131  ;
	input \g1745_reg/NET0131  ;
	input \g1747_reg/NET0131  ;
	input \g1749_reg/NET0131  ;
	input \g174_reg/NET0131  ;
	input \g1750_reg/NET0131  ;
	input \g1754_reg/NET0131  ;
	input \g1757_reg/NET0131  ;
	input \g175_reg/NET0131  ;
	input \g1760_reg/NET0131  ;
	input \g1762_reg/NET0131  ;
	input \g1764_reg/NET0131  ;
	input \g1765_reg/NET0131  ;
	input \g1769_reg/NET0131  ;
	input \g176_reg/NET0131  ;
	input \g1772_reg/NET0131  ;
	input \g1775_reg/NET0131  ;
	input \g1777_reg/NET0131  ;
	input \g1779_reg/NET0131  ;
	input \g177_reg/NET0131  ;
	input \g1783_reg/NET0131  ;
	input \g1784_reg/NET0131  ;
	input \g1785_reg/NET0131  ;
	input \g1789_reg/NET0131  ;
	input \g178_reg/NET0131  ;
	input \g1792_reg/NET0131  ;
	input \g1795_reg/NET0131  ;
	input \g1798_reg/NET0131  ;
	input \g179_reg/NET0131  ;
	input \g1801_reg/NET0131  ;
	input \g1804_reg/NET0131  ;
	input \g1807_reg/NET0131  ;
	input \g1808_reg/NET0131  ;
	input \g1809_reg/NET0131  ;
	input \g1810_reg/NET0131  ;
	input \g1813_reg/NET0131  ;
	input \g1816_reg/NET0131  ;
	input \g1819_reg/NET0131  ;
	input \g1822_reg/NET0131  ;
	input \g1825_reg/NET0131  ;
	input \g1828_reg/NET0131  ;
	input \g1829_reg/NET0131  ;
	input \g1830_reg/NET0131  ;
	input \g1832_reg/NET0131  ;
	input \g1834_reg/NET0131  ;
	input \g1845_reg/NET0131  ;
	input \g1846_reg/NET0131  ;
	input \g1849_reg/NET0131  ;
	input \g1852_reg/NET0131  ;
	input \g1858_reg/NET0131  ;
	input \g1859_reg/NET0131  ;
	input \g185_reg/NET0131  ;
	input \g1860_reg/NET0131  ;
	input \g1861_reg/NET0131  ;
	input \g1865_reg/NET0131  ;
	input \g1867_reg/NET0131  ;
	input \g1868_reg/NET0131  ;
	input \g1869_reg/NET0131  ;
	input \g186_reg/NET0131  ;
	input \g1870_reg/NET0131  ;
	input \g1871_reg/NET0131  ;
	input \g1874_reg/NET0131  ;
	input \g1877_reg/NET0131  ;
	input \g1880_reg/NET0131  ;
	input \g1886_reg/NET0131  ;
	input \g1887_reg/NET0131  ;
	input \g189_reg/NET0131  ;
	input \g1904_reg/NET0131  ;
	input \g1905_reg/NET0131  ;
	input \g1909_reg/NET0131  ;
	input \g1910_reg/NET0131  ;
	input \g1911_reg/NET0131  ;
	input \g1912_reg/NET0131  ;
	input \g1913_reg/NET0131  ;
	input \g1914_reg/NET0131  ;
	input \g1916_reg/NET0131  ;
	input \g1917_reg/NET0131  ;
	input \g1918_reg/NET0131  ;
	input \g1921_reg/NET0131  ;
	input \g1922_reg/NET0131  ;
	input \g1924_reg/NET0131  ;
	input \g1928_reg/NET0131  ;
	input \g192_reg/NET0131  ;
	input \g1939_reg/NET0131  ;
	input \g1943_pad  ;
	input \g1945_reg/NET0131  ;
	input \g1947_reg/NET0131  ;
	input \g1949_reg/NET0131  ;
	input \g1951_reg/NET0131  ;
	input \g1953_reg/NET0131  ;
	input \g1955_reg/NET0131  ;
	input \g1956_reg/NET0131  ;
	input \g1957_reg/NET0131  ;
	input \g1958_reg/NET0131  ;
	input \g1959_reg/NET0131  ;
	input \g195_reg/NET0131  ;
	input \g1960_reg/NET0131  ;
	input \g1961_reg/NET0131  ;
	input \g1962_reg/NET0131  ;
	input \g1963_reg/NET0131  ;
	input \g1964_reg/NET0131  ;
	input \g1965_reg/NET0131  ;
	input \g1966_reg/NET0131  ;
	input \g1967_reg/NET0131  ;
	input \g1970_reg/NET0131  ;
	input \g1973_reg/NET0131  ;
	input \g1976_reg/NET0131  ;
	input \g1979_reg/NET0131  ;
	input \g1982_reg/NET0131  ;
	input \g1985_reg/NET0131  ;
	input \g1988_reg/NET0131  ;
	input \g198_reg/NET0131  ;
	input \g1991_reg/NET0131  ;
	input \g1994_reg/NET0131  ;
	input \g1997_reg/NET0131  ;
	input \g2000_reg/NET0131  ;
	input \g201_reg/NET0131  ;
	input \g204_reg/NET0131  ;
	input \g2078_reg/NET0131  ;
	input \g2079_reg/NET0131  ;
	input \g207_reg/NET0131  ;
	input \g2080_reg/NET0131  ;
	input \g2081_reg/NET0131  ;
	input \g2082_reg/NET0131  ;
	input \g2083_reg/NET0131  ;
	input \g2084_reg/NET0131  ;
	input \g2085_reg/NET0131  ;
	input \g2086_reg/NET0131  ;
	input \g2087_reg/NET0131  ;
	input \g2088_reg/NET0131  ;
	input \g2089_reg/NET0131  ;
	input \g2090_reg/NET0131  ;
	input \g2091_reg/NET0131  ;
	input \g2092_reg/NET0131  ;
	input \g2093_reg/NET0131  ;
	input \g2094_reg/NET0131  ;
	input \g2095_reg/NET0131  ;
	input \g2096_reg/NET0131  ;
	input \g2097_reg/NET0131  ;
	input \g2098_reg/NET0131  ;
	input \g2099_reg/NET0131  ;
	input \g2100_reg/NET0131  ;
	input \g2101_reg/NET0131  ;
	input \g2102_reg/NET0131  ;
	input \g2103_reg/NET0131  ;
	input \g2104_reg/NET0131  ;
	input \g2105_reg/NET0131  ;
	input \g2106_reg/NET0131  ;
	input \g2107_reg/NET0131  ;
	input \g2108_reg/NET0131  ;
	input \g2109_reg/NET0131  ;
	input \g210_reg/NET0131  ;
	input \g2110_reg/NET0131  ;
	input \g2111_reg/NET0131  ;
	input \g2112_reg/NET0131  ;
	input \g2113_reg/NET0131  ;
	input \g2114_reg/NET0131  ;
	input \g2115_reg/NET0131  ;
	input \g2116_reg/NET0131  ;
	input \g2117_reg/NET0131  ;
	input \g2118_reg/NET0131  ;
	input \g2119_reg/NET0131  ;
	input \g213_reg/NET0131  ;
	input \g2165_reg/NET0131  ;
	input \g216_reg/NET0131  ;
	input \g2170_reg/NET0131  ;
	input \g2175_reg/NET0131  ;
	input \g2180_reg/NET0131  ;
	input \g2185_reg/NET0131  ;
	input \g2190_reg/NET0131  ;
	input \g2195_reg/NET0131  ;
	input \g219_reg/NET0131  ;
	input \g2200_reg/NET0131  ;
	input \g2205_reg/NET0131  ;
	input \g2206_reg/NET0131  ;
	input \g2207_reg/NET0131  ;
	input \g2208_reg/NET0131  ;
	input \g2209_reg/NET0131  ;
	input \g2210_reg/NET0131  ;
	input \g2217_reg/NET0131  ;
	input \g2218_reg/NET0131  ;
	input \g2219_reg/NET0131  ;
	input \g2220_reg/NET0131  ;
	input \g2221_reg/NET0131  ;
	input \g2222_reg/NET0131  ;
	input \g2223_reg/NET0131  ;
	input \g2224_reg/NET0131  ;
	input \g2225_reg/NET0131  ;
	input \g2226_reg/NET0131  ;
	input \g2227_reg/NET0131  ;
	input \g2228_reg/NET0131  ;
	input \g2229_reg/NET0131  ;
	input \g222_reg/NET0131  ;
	input \g2230_reg/NET0131  ;
	input \g2231_reg/NET0131  ;
	input \g2232_reg/NET0131  ;
	input \g2233_reg/NET0131  ;
	input \g2234_reg/NET0131  ;
	input \g2235_reg/NET0131  ;
	input \g2236_reg/NET0131  ;
	input \g2237_reg/NET0131  ;
	input \g2238_reg/NET0131  ;
	input \g2239_reg/NET0131  ;
	input \g2240_reg/NET0131  ;
	input \g2244_reg/NET0131  ;
	input \g2245_reg/NET0131  ;
	input \g2246_reg/NET0131  ;
	input \g2247_reg/NET0131  ;
	input \g2248_reg/NET0131  ;
	input \g2249_reg/NET0131  ;
	input \g2250_reg/NET0131  ;
	input \g2251_reg/NET0131  ;
	input \g2252_reg/NET0131  ;
	input \g2253_reg/NET0131  ;
	input \g2254_reg/NET0131  ;
	input \g2255_reg/NET0131  ;
	input \g225_reg/NET0131  ;
	input \g2261_reg/NET0131  ;
	input \g2264_reg/NET0131  ;
	input \g2267_reg/NET0131  ;
	input \g2270_reg/NET0131  ;
	input \g2273_reg/NET0131  ;
	input \g2276_reg/NET0131  ;
	input \g2279_reg/NET0131  ;
	input \g2282_reg/NET0131  ;
	input \g2285_reg/NET0131  ;
	input \g2288_reg/NET0131  ;
	input \g228_reg/NET0131  ;
	input \g2291_reg/NET0131  ;
	input \g2294_reg/NET0131  ;
	input \g2297_reg/NET0131  ;
	input \g2300_reg/NET0131  ;
	input \g2303_reg/NET0131  ;
	input \g2306_reg/NET0131  ;
	input \g2309_reg/NET0131  ;
	input \g2312_reg/NET0131  ;
	input \g2315_reg/NET0131  ;
	input \g2318_reg/NET0131  ;
	input \g231_reg/NET0131  ;
	input \g2321_reg/NET0131  ;
	input \g2324_reg/NET0131  ;
	input \g2327_reg/NET0131  ;
	input \g2330_reg/NET0131  ;
	input \g2333_reg/NET0131  ;
	input \g2336_reg/NET0131  ;
	input \g2339_reg/NET0131  ;
	input \g2342_reg/NET0131  ;
	input \g2345_reg/NET0131  ;
	input \g2348_reg/NET0131  ;
	input \g234_reg/NET0131  ;
	input \g2354_reg/NET0131  ;
	input \g2356_reg/NET0131  ;
	input \g2358_reg/NET0131  ;
	input \g2360_reg/NET0131  ;
	input \g2362_reg/NET0131  ;
	input \g2364_reg/NET0131  ;
	input \g2366_reg/NET0131  ;
	input \g2373_reg/NET0131  ;
	input \g2374_reg/NET0131  ;
	input \g237_reg/NET0131  ;
	input \g2380_reg/NET0131  ;
	input \g2387_reg/NET0131  ;
	input \g2388_reg/NET0131  ;
	input \g2389_reg/NET0131  ;
	input \g2390_reg/NET0131  ;
	input \g2391_reg/NET0131  ;
	input \g2392_reg/NET0131  ;
	input \g2393_reg/NET0131  ;
	input \g2394_reg/NET0131  ;
	input \g2395_reg/NET0131  ;
	input \g2396_reg/NET0131  ;
	input \g2397_reg/NET0131  ;
	input \g2398_reg/NET0131  ;
	input \g2399_reg/NET0131  ;
	input \g240_reg/NET0131  ;
	input \g2418_reg/NET0131  ;
	input \g2421_reg/NET0131  ;
	input \g2424_reg/NET0131  ;
	input \g2426_reg/NET0131  ;
	input \g2428_reg/NET0131  ;
	input \g2429_reg/NET0131  ;
	input \g2433_reg/NET0131  ;
	input \g2436_reg/NET0131  ;
	input \g2439_reg/NET0131  ;
	input \g243_reg/NET0131  ;
	input \g2441_reg/NET0131  ;
	input \g2443_reg/NET0131  ;
	input \g2444_reg/NET0131  ;
	input \g2448_reg/NET0131  ;
	input \g2451_reg/NET0131  ;
	input \g2454_reg/NET0131  ;
	input \g2456_reg/NET0131  ;
	input \g2458_reg/NET0131  ;
	input \g2459_reg/NET0131  ;
	input \g2463_reg/NET0131  ;
	input \g2466_reg/NET0131  ;
	input \g2469_reg/NET0131  ;
	input \g246_reg/NET0131  ;
	input \g2471_reg/NET0131  ;
	input \g2473_reg/NET0131  ;
	input \g2477_reg/NET0131  ;
	input \g2478_reg/NET0131  ;
	input \g2479_reg/NET0131  ;
	input \g2483_reg/NET0131  ;
	input \g2486_reg/NET0131  ;
	input \g2489_reg/NET0131  ;
	input \g2492_reg/NET0131  ;
	input \g2495_reg/NET0131  ;
	input \g2498_reg/NET0131  ;
	input \g249_reg/NET0131  ;
	input \g2501_reg/NET0131  ;
	input \g2502_reg/NET0131  ;
	input \g2503_reg/NET0131  ;
	input \g2504_reg/NET0131  ;
	input \g2507_reg/NET0131  ;
	input \g2510_reg/NET0131  ;
	input \g2513_reg/NET0131  ;
	input \g2516_reg/NET0131  ;
	input \g2519_reg/NET0131  ;
	input \g2522_reg/NET0131  ;
	input \g2523_reg/NET0131  ;
	input \g2524_reg/NET0131  ;
	input \g2526_reg/NET0131  ;
	input \g2528_reg/NET0131  ;
	input \g252_reg/NET0131  ;
	input \g2539_reg/NET0131  ;
	input \g2540_reg/NET0131  ;
	input \g2543_reg/NET0131  ;
	input \g2546_reg/NET0131  ;
	input \g2552_reg/NET0131  ;
	input \g2553_reg/NET0131  ;
	input \g2554_reg/NET0131  ;
	input \g2555_reg/NET0131  ;
	input \g2559_reg/NET0131  ;
	input \g255_reg/NET0131  ;
	input \g2561_reg/NET0131  ;
	input \g2562_reg/NET0131  ;
	input \g2563_reg/NET0131  ;
	input \g2564_reg/NET0131  ;
	input \g2565_reg/NET0131  ;
	input \g2568_reg/NET0131  ;
	input \g2571_reg/NET0131  ;
	input \g2574_reg/NET0131  ;
	input \g2580_reg/NET0131  ;
	input \g2581_reg/NET0131  ;
	input \g258_reg/NET0131  ;
	input \g2598_reg/NET0131  ;
	input \g2599_reg/NET0131  ;
	input \g2603_reg/NET0131  ;
	input \g2604_reg/NET0131  ;
	input \g2605_reg/NET0131  ;
	input \g2606_reg/NET0131  ;
	input \g2607_reg/NET0131  ;
	input \g2608_reg/NET0131  ;
	input \g2610_reg/NET0131  ;
	input \g2611_reg/NET0131  ;
	input \g2612_reg/NET0131  ;
	input \g2615_reg/NET0131  ;
	input \g2616_reg/NET0131  ;
	input \g2618_reg/NET0131  ;
	input \g261_reg/NET0131  ;
	input \g2622_reg/NET0131  ;
	input \g2633_reg/NET0131  ;
	input \g2637_pad  ;
	input \g2639_reg/NET0131  ;
	input \g2641_reg/NET0131  ;
	input \g2643_reg/NET0131  ;
	input \g2645_reg/NET0131  ;
	input \g2647_reg/NET0131  ;
	input \g2649_reg/NET0131  ;
	input \g264_reg/NET0131  ;
	input \g2650_reg/NET0131  ;
	input \g2651_reg/NET0131  ;
	input \g2652_reg/NET0131  ;
	input \g2653_reg/NET0131  ;
	input \g2654_reg/NET0131  ;
	input \g2655_reg/NET0131  ;
	input \g2656_reg/NET0131  ;
	input \g2657_reg/NET0131  ;
	input \g2658_reg/NET0131  ;
	input \g2659_reg/NET0131  ;
	input \g2660_reg/NET0131  ;
	input \g2661_reg/NET0131  ;
	input \g2664_reg/NET0131  ;
	input \g2667_reg/NET0131  ;
	input \g2670_reg/NET0131  ;
	input \g2673_reg/NET0131  ;
	input \g2676_reg/NET0131  ;
	input \g2679_reg/NET0131  ;
	input \g267_reg/NET0131  ;
	input \g2682_reg/NET0131  ;
	input \g2685_reg/NET0131  ;
	input \g2688_reg/NET0131  ;
	input \g2691_reg/NET0131  ;
	input \g2694_reg/NET0131  ;
	input \g270_reg/NET0131  ;
	input \g273_reg/NET0131  ;
	input \g2772_reg/NET0131  ;
	input \g2773_reg/NET0131  ;
	input \g2774_reg/NET0131  ;
	input \g2775_reg/NET0131  ;
	input \g2776_reg/NET0131  ;
	input \g2777_reg/NET0131  ;
	input \g2778_reg/NET0131  ;
	input \g2779_reg/NET0131  ;
	input \g2780_reg/NET0131  ;
	input \g2781_reg/NET0131  ;
	input \g2782_reg/NET0131  ;
	input \g2783_reg/NET0131  ;
	input \g2784_reg/NET0131  ;
	input \g2785_reg/NET0131  ;
	input \g2786_reg/NET0131  ;
	input \g2787_reg/NET0131  ;
	input \g2788_reg/NET0131  ;
	input \g2789_reg/NET0131  ;
	input \g2790_reg/NET0131  ;
	input \g2791_reg/NET0131  ;
	input \g2792_reg/NET0131  ;
	input \g2793_reg/NET0131  ;
	input \g2794_reg/NET0131  ;
	input \g2795_reg/NET0131  ;
	input \g2796_reg/NET0131  ;
	input \g2797_reg/NET0131  ;
	input \g2798_reg/NET0131  ;
	input \g2799_reg/NET0131  ;
	input \g279_reg/NET0131  ;
	input \g2800_reg/NET0131  ;
	input \g2801_reg/NET0131  ;
	input \g2802_reg/NET0131  ;
	input \g2803_reg/NET0131  ;
	input \g2804_reg/NET0131  ;
	input \g2805_reg/NET0131  ;
	input \g2806_reg/NET0131  ;
	input \g2807_reg/NET0131  ;
	input \g2808_reg/NET0131  ;
	input \g2809_reg/NET0131  ;
	input \g2810_reg/NET0131  ;
	input \g2811_reg/NET0131  ;
	input \g2812_reg/NET0131  ;
	input \g2813_reg/NET0131  ;
	input \g2814_reg/NET0131  ;
	input \g2817_reg/NET0131  ;
	input \g281_reg/NET0131  ;
	input \g283_reg/NET0131  ;
	input \g285_reg/NET0131  ;
	input \g2874_reg/NET0131  ;
	input \g2879_reg/NET0131  ;
	input \g287_reg/NET0131  ;
	input \g2883_reg/NET0131  ;
	input \g2888_reg/NET0131  ;
	input \g2892_reg/NET0131  ;
	input \g2896_reg/NET0131  ;
	input \g289_reg/NET0131  ;
	input \g2900_reg/NET0131  ;
	input \g2903_reg/NET0131  ;
	input \g2908_reg/NET0131  ;
	input \g2912_reg/NET0131  ;
	input \g2917_reg/NET0131  ;
	input \g291_reg/NET0131  ;
	input \g2920_reg/NET0131  ;
	input \g2924_reg/NET0131  ;
	input \g2929_reg/NET0131  ;
	input \g2933_reg/NET0131  ;
	input \g2934_reg/NET0131  ;
	input \g2935_reg/NET0131  ;
	input \g2938_reg/NET0131  ;
	input \g2941_reg/NET0131  ;
	input \g2944_reg/NET0131  ;
	input \g2947_reg/NET0131  ;
	input \g2950_reg/NET0131  ;
	input \g2953_reg/NET0131  ;
	input \g2956_reg/NET0131  ;
	input \g2959_reg/NET0131  ;
	input \g2962_reg/NET0131  ;
	input \g2963_reg/NET0131  ;
	input \g2966_reg/NET0131  ;
	input \g2969_reg/NET0131  ;
	input \g2972_reg/NET0131  ;
	input \g2975_reg/NET0131  ;
	input \g2978_reg/NET0131  ;
	input \g2981_reg/NET0131  ;
	input \g2984_reg/NET0131  ;
	input \g2985_reg/NET0131  ;
	input \g2986_reg/NET0131  ;
	input \g2987_reg/NET0131  ;
	input \g298_reg/NET0131  ;
	input \g2990_reg/NET0131  ;
	input \g2991_reg/NET0131  ;
	input \g2992_reg/NET0131  ;
	input \g2993_reg/NET0131  ;
	input \g2997_reg/NET0131  ;
	input \g2998_reg/NET0131  ;
	input \g299_reg/NET0131  ;
	input \g3002_reg/NET0131  ;
	input \g3006_reg/NET0131  ;
	input \g3010_reg/NET0131  ;
	input \g3013_reg/NET0131  ;
	input \g3018_reg/NET0131  ;
	input \g3024_reg/NET0131  ;
	input \g3028_reg/NET0131  ;
	input \g3032_reg/NET0131  ;
	input \g3036_reg/NET0131  ;
	input \g3043_reg/NET0131  ;
	input \g3044_reg/NET0131  ;
	input \g3045_reg/NET0131  ;
	input \g3046_reg/NET0131  ;
	input \g3047_reg/NET0131  ;
	input \g3048_reg/NET0131  ;
	input \g3049_reg/NET0131  ;
	input \g3050_reg/NET0131  ;
	input \g3051_reg/NET0131  ;
	input \g3052_reg/NET0131  ;
	input \g3053_reg/NET0131  ;
	input \g3054_reg/NET0131  ;
	input \g3055_reg/NET0131  ;
	input \g3056_reg/NET0131  ;
	input \g3057_reg/NET0131  ;
	input \g3058_reg/NET0131  ;
	input \g3059_reg/NET0131  ;
	input \g305_reg/NET0131  ;
	input \g3060_reg/NET0131  ;
	input \g3061_reg/NET0131  ;
	input \g3062_reg/NET0131  ;
	input \g3063_reg/NET0131  ;
	input \g3064_reg/NET0131  ;
	input \g3065_reg/NET0131  ;
	input \g3066_reg/NET0131  ;
	input \g3067_reg/NET0131  ;
	input \g3068_reg/NET0131  ;
	input \g3069_reg/NET0131  ;
	input \g3070_reg/NET0131  ;
	input \g3071_reg/NET0131  ;
	input \g3072_reg/NET0131  ;
	input \g3073_reg/NET0131  ;
	input \g3074_reg/NET0131  ;
	input \g3075_reg/NET0131  ;
	input \g3076_reg/NET0131  ;
	input \g3077_reg/NET0131  ;
	input \g3078_reg/NET0131  ;
	input \g3079_reg/NET0131  ;
	input \g3080_reg/NET0131  ;
	input \g3083_reg/NET0131  ;
	input \g3097_reg/NET0131  ;
	input \g3110_reg/NET0131  ;
	input \g3114_reg/NET0131  ;
	input \g3120_reg/NET0131  ;
	input \g312_reg/NET0131  ;
	input \g3139_reg/NET0131  ;
	input \g313_reg/NET0131  ;
	input \g314_reg/NET0131  ;
	input \g315_reg/NET0131  ;
	input \g316_reg/NET0131  ;
	input \g317_reg/NET0131  ;
	input \g318_reg/NET0131  ;
	input \g319_reg/NET0131  ;
	input \g320_reg/NET0131  ;
	input \g321_reg/NET0131  ;
	input \g3229_pad  ;
	input \g322_reg/NET0131  ;
	input \g3230_pad  ;
	input \g3231_pad  ;
	input \g3233_pad  ;
	input \g3234_pad  ;
	input \g323_reg/NET0131  ;
	input \g324_reg/NET0131  ;
	input \g343_reg/NET0131  ;
	input \g346_reg/NET0131  ;
	input \g349_reg/NET0131  ;
	input \g351_reg/NET0131  ;
	input \g353_reg/NET0131  ;
	input \g354_reg/NET0131  ;
	input \g358_reg/NET0131  ;
	input \g361_reg/NET0131  ;
	input \g364_reg/NET0131  ;
	input \g366_reg/NET0131  ;
	input \g368_reg/NET0131  ;
	input \g369_reg/NET0131  ;
	input \g373_reg/NET0131  ;
	input \g376_reg/NET0131  ;
	input \g379_reg/NET0131  ;
	input \g381_reg/NET0131  ;
	input \g383_reg/NET0131  ;
	input \g384_reg/NET0131  ;
	input \g388_reg/NET0131  ;
	input \g391_reg/NET0131  ;
	input \g394_reg/NET0131  ;
	input \g396_reg/NET0131  ;
	input \g398_reg/NET0131  ;
	input \g402_reg/NET0131  ;
	input \g403_reg/NET0131  ;
	input \g404_reg/NET0131  ;
	input \g408_reg/NET0131  ;
	input \g411_reg/NET0131  ;
	input \g414_reg/NET0131  ;
	input \g417_reg/NET0131  ;
	input \g420_reg/NET0131  ;
	input \g423_reg/NET0131  ;
	input \g426_reg/NET0131  ;
	input \g427_reg/NET0131  ;
	input \g428_reg/NET0131  ;
	input \g429_reg/NET0131  ;
	input \g432_reg/NET0131  ;
	input \g435_reg/NET0131  ;
	input \g438_reg/NET0131  ;
	input \g441_reg/NET0131  ;
	input \g444_reg/NET0131  ;
	input \g447_reg/NET0131  ;
	input \g448_reg/NET0131  ;
	input \g449_reg/NET0131  ;
	input \g451_reg/NET0131  ;
	input \g453_reg/NET0131  ;
	input \g464_reg/NET0131  ;
	input \g465_reg/NET0131  ;
	input \g468_reg/NET0131  ;
	input \g471_reg/NET0131  ;
	input \g477_reg/NET0131  ;
	input \g478_reg/NET0131  ;
	input \g479_reg/NET0131  ;
	input \g480_reg/NET0131  ;
	input \g484_reg/NET0131  ;
	input \g486_reg/NET0131  ;
	input \g487_reg/NET0131  ;
	input \g488_reg/NET0131  ;
	input \g489_reg/NET0131  ;
	input \g490_reg/NET0131  ;
	input \g493_reg/NET0131  ;
	input \g496_reg/NET0131  ;
	input \g499_reg/NET0131  ;
	input \g506_reg/NET0131  ;
	input \g507_reg/NET0131  ;
	input \g51_pad  ;
	input \g524_reg/NET0131  ;
	input \g525_reg/NET0131  ;
	input \g529_reg/NET0131  ;
	input \g530_reg/NET0131  ;
	input \g531_reg/NET0131  ;
	input \g532_reg/NET0131  ;
	input \g533_reg/NET0131  ;
	input \g534_reg/NET0131  ;
	input \g536_reg/NET0131  ;
	input \g537_reg/NET0131  ;
	input \g5388_pad  ;
	input \g538_reg/NET0131  ;
	input \g541_reg/NET0131  ;
	input \g542_reg/NET0131  ;
	input \g544_reg/NET0131  ;
	input \g548_reg/NET0131  ;
	input \g559_reg/NET0131  ;
	input \g563_pad  ;
	input \g5657_pad  ;
	input \g565_reg/NET0131  ;
	input \g567_reg/NET0131  ;
	input \g569_reg/NET0131  ;
	input \g571_reg/NET0131  ;
	input \g573_reg/NET0131  ;
	input \g575_reg/NET0131  ;
	input \g576_reg/NET0131  ;
	input \g577_reg/NET0131  ;
	input \g578_reg/NET0131  ;
	input \g579_reg/NET0131  ;
	input \g580_reg/NET0131  ;
	input \g581_reg/NET0131  ;
	input \g582_reg/NET0131  ;
	input \g583_reg/NET0131  ;
	input \g584_reg/NET0131  ;
	input \g585_reg/NET0131  ;
	input \g586_reg/NET0131  ;
	input \g587_reg/NET0131  ;
	input \g590_reg/NET0131  ;
	input \g593_reg/NET0131  ;
	input \g596_reg/NET0131  ;
	input \g599_reg/NET0131  ;
	input \g602_reg/NET0131  ;
	input \g605_reg/NET0131  ;
	input \g608_reg/NET0131  ;
	input \g611_reg/NET0131  ;
	input \g614_reg/NET0131  ;
	input \g617_reg/NET0131  ;
	input \g620_reg/NET0131  ;
	input \g698_reg/NET0131  ;
	input \g699_reg/NET0131  ;
	input \g700_reg/NET0131  ;
	input \g701_reg/NET0131  ;
	input \g702_reg/NET0131  ;
	input \g703_reg/NET0131  ;
	input \g704_reg/NET0131  ;
	input \g705_reg/NET0131  ;
	input \g706_reg/NET0131  ;
	input \g707_reg/NET0131  ;
	input \g708_reg/NET0131  ;
	input \g709_reg/NET0131  ;
	input \g710_reg/NET0131  ;
	input \g711_reg/NET0131  ;
	input \g712_reg/NET0131  ;
	input \g713_reg/NET0131  ;
	input \g714_reg/NET0131  ;
	input \g715_reg/NET0131  ;
	input \g716_reg/NET0131  ;
	input \g717_reg/NET0131  ;
	input \g718_reg/NET0131  ;
	input \g719_reg/NET0131  ;
	input \g720_reg/NET0131  ;
	input \g721_reg/NET0131  ;
	input \g722_reg/NET0131  ;
	input \g723_reg/NET0131  ;
	input \g724_reg/NET0131  ;
	input \g725_reg/NET0131  ;
	input \g726_reg/NET0131  ;
	input \g727_reg/NET0131  ;
	input \g728_reg/NET0131  ;
	input \g729_reg/NET0131  ;
	input \g730_reg/NET0131  ;
	input \g731_reg/NET0131  ;
	input \g732_reg/NET0131  ;
	input \g733_reg/NET0131  ;
	input \g734_reg/NET0131  ;
	input \g735_reg/NET0131  ;
	input \g736_reg/NET0131  ;
	input \g737_reg/NET0131  ;
	input \g738_reg/NET0131  ;
	input \g739_reg/NET0131  ;
	input \g785_reg/NET0131  ;
	input \g789_reg/NET0131  ;
	input \g793_reg/NET0131  ;
	input \g7961_pad  ;
	input \g797_reg/NET0131  ;
	input \g801_reg/NET0131  ;
	input \g805_reg/NET0131  ;
	input \g809_reg/NET0131  ;
	input \g813_reg/NET0131  ;
	input \g817_reg/NET0131  ;
	input \g818_reg/NET0131  ;
	input \g819_reg/NET0131  ;
	input \g820_reg/NET0131  ;
	input \g821_reg/NET0131  ;
	input \g822_reg/NET0131  ;
	input \g8259_pad  ;
	input \g8260_pad  ;
	input \g8261_pad  ;
	input \g8262_pad  ;
	input \g8263_pad  ;
	input \g8264_pad  ;
	input \g8265_pad  ;
	input \g8266_pad  ;
	input \g8268_pad  ;
	input \g8269_pad  ;
	input \g8270_pad  ;
	input \g8271_pad  ;
	input \g8272_pad  ;
	input \g8273_pad  ;
	input \g8274_pad  ;
	input \g8275_pad  ;
	input \g829_reg/NET0131  ;
	input \g830_reg/NET0131  ;
	input \g831_reg/NET0131  ;
	input \g832_reg/NET0131  ;
	input \g833_reg/NET0131  ;
	input \g834_reg/NET0131  ;
	input \g835_reg/NET0131  ;
	input \g836_reg/NET0131  ;
	input \g837_reg/NET0131  ;
	input \g838_reg/NET0131  ;
	input \g839_reg/NET0131  ;
	input \g840_reg/NET0131  ;
	input \g841_reg/NET0131  ;
	input \g842_reg/NET0131  ;
	input \g843_reg/NET0131  ;
	input \g844_reg/NET0131  ;
	input \g845_reg/NET0131  ;
	input \g846_reg/NET0131  ;
	input \g847_reg/NET0131  ;
	input \g848_reg/NET0131  ;
	input \g849_reg/NET0131  ;
	input \g850_reg/NET0131  ;
	input \g851_reg/NET0131  ;
	input \g852_reg/NET0131  ;
	input \g856_reg/NET0131  ;
	input \g857_reg/NET0131  ;
	input \g858_reg/NET0131  ;
	input \g859_reg/NET0131  ;
	input \g860_reg/NET0131  ;
	input \g861_reg/NET0131  ;
	input \g862_reg/NET0131  ;
	input \g863_reg/NET0131  ;
	input \g864_reg/NET0131  ;
	input \g865_reg/NET0131  ;
	input \g866_reg/NET0131  ;
	input \g867_reg/NET0131  ;
	input \g873_reg/NET0131  ;
	input \g876_reg/NET0131  ;
	input \g879_reg/NET0131  ;
	input \g882_reg/NET0131  ;
	input \g885_reg/NET0131  ;
	input \g888_reg/NET0131  ;
	input \g891_reg/NET0131  ;
	input \g894_reg/NET0131  ;
	input \g897_reg/NET0131  ;
	input \g900_reg/NET0131  ;
	input \g903_reg/NET0131  ;
	input \g906_reg/NET0131  ;
	input \g909_reg/NET0131  ;
	input \g912_reg/NET0131  ;
	input \g915_reg/NET0131  ;
	input \g918_reg/NET0131  ;
	input \g921_reg/NET0131  ;
	input \g924_reg/NET0131  ;
	input \g927_reg/NET0131  ;
	input \g930_reg/NET0131  ;
	input \g933_reg/NET0131  ;
	input \g936_reg/NET0131  ;
	input \g939_reg/NET0131  ;
	input \g942_reg/NET0131  ;
	input \g945_reg/NET0131  ;
	input \g948_reg/NET0131  ;
	input \g951_reg/NET0131  ;
	input \g954_reg/NET0131  ;
	input \g957_reg/NET0131  ;
	input \g960_reg/NET0131  ;
	input \g966_reg/NET0131  ;
	input \g968_reg/NET0131  ;
	input \g970_reg/NET0131  ;
	input \g972_reg/NET0131  ;
	input \g974_reg/NET0131  ;
	input \g976_reg/NET0131  ;
	input \g978_reg/NET0131  ;
	input \g97_reg/NET0131  ;
	input \g985_reg/NET0131  ;
	input \g986_reg/NET0131  ;
	input \g992_reg/NET0131  ;
	input \g999_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g101_reg/P0001  ;
	output \g105_reg/P0001  ;
	output \g109_reg/P0001  ;
	output \g1138_reg/P0001  ;
	output \g113_reg/P0001  ;
	output \g1140_reg/P0001  ;
	output \g117_reg/P0001  ;
	output \g121_reg/P0001  ;
	output \g125_reg/P0001  ;
	output \g1471_reg/P0001  ;
	output \g1476_reg/P0001  ;
	output \g1481_reg/P0001  ;
	output \g1486_reg/P0001  ;
	output \g1491_reg/P0001  ;
	output \g1496_reg/P0001  ;
	output \g1501_reg/P0001  ;
	output \g1506_reg/P0001  ;
	output \g16496_pad  ;
	output \g1660_reg/P0001  ;
	output \g1662_reg/P0001  ;
	output \g1664_reg/P0001  ;
	output \g1666_reg/P0001  ;
	output \g1668_reg/P0001  ;
	output \g1670_reg/P0001  ;
	output \g1672_reg/P0001  ;
	output \g18/_0_  ;
	output \g1832_reg/P0001  ;
	output \g1834_reg/P0001  ;
	output \g2165_reg/P0001  ;
	output \g2170_reg/P0001  ;
	output \g2175_reg/P0001  ;
	output \g2180_reg/P0001  ;
	output \g2185_reg/P0001  ;
	output \g2190_reg/P0001  ;
	output \g2195_reg/P0001  ;
	output \g2200_reg/P0001  ;
	output \g2354_reg/P0001  ;
	output \g2356_reg/P0001  ;
	output \g2358_reg/P0001  ;
	output \g2360_reg/P0001  ;
	output \g2362_reg/P0001  ;
	output \g2364_reg/P0001  ;
	output \g2366_reg/P0001  ;
	output \g2526_reg/P0001  ;
	output \g2528_reg/P0001  ;
	output \g25489_pad  ;
	output \g279_reg/P0001  ;
	output \g281_reg/P0001  ;
	output \g283_reg/P0001  ;
	output \g285_reg/P0001  ;
	output \g2879_reg/NET0131_syn_2  ;
	output \g287_reg/P0001  ;
	output \g289_reg/P0001  ;
	output \g291_reg/P0001  ;
	output \g451_reg/P0001  ;
	output \g453_reg/P0001  ;
	output \g59421/_3_  ;
	output \g59425/_1_  ;
	output \g59435/_0_  ;
	output \g59436/_0_  ;
	output \g59441/_3_  ;
	output \g59442/_0_  ;
	output \g59445/_0_  ;
	output \g59453/_0_  ;
	output \g59462/_3_  ;
	output \g59466/_3_  ;
	output \g59467/_3_  ;
	output \g59468/_3_  ;
	output \g59469/_3_  ;
	output \g59470/_3_  ;
	output \g59471/_3_  ;
	output \g59472/_3_  ;
	output \g59473/_3_  ;
	output \g59489/_0_  ;
	output \g59498/_0_  ;
	output \g59499/_0_  ;
	output \g59500/_0_  ;
	output \g59502/_2_  ;
	output \g59503/_0_  ;
	output \g59505/_2_  ;
	output \g59507/_0_  ;
	output \g59508/_0_  ;
	output \g59533/_3_  ;
	output \g59534/_3_  ;
	output \g59535/_3_  ;
	output \g59536/_3_  ;
	output \g59537/_3_  ;
	output \g59538/_3_  ;
	output \g59539/_3_  ;
	output \g59540/_3_  ;
	output \g59548/_0_  ;
	output \g59550/_0_  ;
	output \g59551/_0_  ;
	output \g59552/_0_  ;
	output \g59554/_0_  ;
	output \g59555/_0_  ;
	output \g59556/_0_  ;
	output \g59557/_0_  ;
	output \g59558/_0_  ;
	output \g59559/_0_  ;
	output \g59560/_0_  ;
	output \g59561/_0_  ;
	output \g59639/_0_  ;
	output \g59694/_2_  ;
	output \g59695/_0_  ;
	output \g59697/_2_  ;
	output \g59698/_0_  ;
	output \g59699/_0_  ;
	output \g59700/_0_  ;
	output \g59705/_0_  ;
	output \g59706/_0_  ;
	output \g59707/_0_  ;
	output \g59708/_0_  ;
	output \g59709/_0_  ;
	output \g59710/_0_  ;
	output \g59711/_0_  ;
	output \g59712/_0_  ;
	output \g59713/_0_  ;
	output \g59714/_0_  ;
	output \g59715/_0_  ;
	output \g59716/_0_  ;
	output \g59717/_0_  ;
	output \g59718/_0_  ;
	output \g59719/_0_  ;
	output \g59720/_0_  ;
	output \g59721/_0_  ;
	output \g59722/_0_  ;
	output \g59723/_0_  ;
	output \g59724/_0_  ;
	output \g59725/_0_  ;
	output \g59726/_0_  ;
	output \g59727/_0_  ;
	output \g59728/_0_  ;
	output \g59729/_0_  ;
	output \g59730/_0_  ;
	output \g59731/_0_  ;
	output \g59732/_0_  ;
	output \g59733/_0_  ;
	output \g59734/_0_  ;
	output \g59735/_0_  ;
	output \g59736/_0_  ;
	output \g59737/_0_  ;
	output \g59738/_0_  ;
	output \g59739/_0_  ;
	output \g59740/_0_  ;
	output \g59741/_0_  ;
	output \g59742/_0_  ;
	output \g59743/_0_  ;
	output \g59744/_0_  ;
	output \g59745/_0_  ;
	output \g59747/_0_  ;
	output \g59748/_0_  ;
	output \g59749/_0_  ;
	output \g59750/_0_  ;
	output \g59751/_0_  ;
	output \g59752/_0_  ;
	output \g59753/_0_  ;
	output \g59754/_0_  ;
	output \g59755/_0_  ;
	output \g59756/_0_  ;
	output \g59757/_0_  ;
	output \g59758/_0_  ;
	output \g59759/_0_  ;
	output \g59760/_0_  ;
	output \g59761/_0_  ;
	output \g59762/_0_  ;
	output \g59763/_0_  ;
	output \g59764/_0_  ;
	output \g59765/_0_  ;
	output \g59766/_0_  ;
	output \g59915/_0_  ;
	output \g59952/_2_  ;
	output \g60046/_0_  ;
	output \g60048/_0_  ;
	output \g60049/_0_  ;
	output \g60051/_0_  ;
	output \g60063/_0_  ;
	output \g60103/_0_  ;
	output \g60104/_0_  ;
	output \g60105/_0_  ;
	output \g60107/_2_  ;
	output \g60108/_0_  ;
	output \g60109/_0_  ;
	output \g60110/_0_  ;
	output \g60112/_2_  ;
	output \g60119/_0_  ;
	output \g60120/_0_  ;
	output \g60121/_0_  ;
	output \g60122/_0_  ;
	output \g60123/_0_  ;
	output \g60124/_0_  ;
	output \g60126/_0_  ;
	output \g60127/_0_  ;
	output \g60128/_0_  ;
	output \g60129/_0_  ;
	output \g60130/_0_  ;
	output \g60135/_0_  ;
	output \g60136/_0_  ;
	output \g60137/_0_  ;
	output \g60138/_0_  ;
	output \g60139/_0_  ;
	output \g60143/_3_  ;
	output \g60144/_0_  ;
	output \g60145/_0_  ;
	output \g60339/_0_  ;
	output \g60404/_0_  ;
	output \g60427/_0_  ;
	output \g60428/_0_  ;
	output \g60429/_0_  ;
	output \g60434/_0_  ;
	output \g60435/_0_  ;
	output \g60437/_0_  ;
	output \g60438/_0_  ;
	output \g60439/_0_  ;
	output \g60440/_0_  ;
	output \g60441/_0_  ;
	output \g60448/_0_  ;
	output \g60451/_0_  ;
	output \g60452/_0_  ;
	output \g60453/_0_  ;
	output \g60459/_0_  ;
	output \g60460/_0_  ;
	output \g60523/_0_  ;
	output \g60534/_0_  ;
	output \g60535/_0_  ;
	output \g60536/_0_  ;
	output \g60585/_0_  ;
	output \g60586/_0_  ;
	output \g60587/_0_  ;
	output \g60588/_0_  ;
	output \g60591/_0_  ;
	output \g60592/_0_  ;
	output \g60599/_0_  ;
	output \g60601/_0_  ;
	output \g60602/_0_  ;
	output \g60603/_0_  ;
	output \g60604/_0_  ;
	output \g60605/_0_  ;
	output \g60606/_0_  ;
	output \g60607/_0_  ;
	output \g60608/_0_  ;
	output \g60609/_0_  ;
	output \g60613/_0_  ;
	output \g60614/_0_  ;
	output \g60615/_0_  ;
	output \g60694/_0_  ;
	output \g60708/_0_  ;
	output \g60709/_0_  ;
	output \g60710/_0_  ;
	output \g60785/_0_  ;
	output \g60787/_0_  ;
	output \g60788/_0_  ;
	output \g60799/_0_  ;
	output \g60801/_0_  ;
	output \g60802/_0_  ;
	output \g60803/_1__syn_2  ;
	output \g60805/_1__syn_2  ;
	output \g60806/_1__syn_2  ;
	output \g60808/_0_  ;
	output \g60810/_0_  ;
	output \g60811/_0_  ;
	output \g60825/_3_  ;
	output \g60896/_0_  ;
	output \g60980/_0_  ;
	output \g60981/_0_  ;
	output \g60985/_0_  ;
	output \g60986/_0_  ;
	output \g61012/_0_  ;
	output \g61013/_0_  ;
	output \g61015/_0_  ;
	output \g61017/_0_  ;
	output \g61122/_0_  ;
	output \g61123/_0_  ;
	output \g61124/_0_  ;
	output \g61125/_0_  ;
	output \g61222/_0_  ;
	output \g61223/_0_  ;
	output \g61224/_0_  ;
	output \g61225/_0_  ;
	output \g61228/_0_  ;
	output \g61229/_0_  ;
	output \g61230/_0_  ;
	output \g61231/_0_  ;
	output \g61281/_0_  ;
	output \g61293/_1_  ;
	output \g61307/_0__syn_2  ;
	output \g61309/_0__syn_2  ;
	output \g61310/_0__syn_2  ;
	output \g61311/_1_  ;
	output \g61312/_1_  ;
	output \g61313/_1_  ;
	output \g61324/_1_  ;
	output \g61325/_1_  ;
	output \g61326/_1_  ;
	output \g61328/_1_  ;
	output \g61329/_1_  ;
	output \g61330/_1_  ;
	output \g61332/_1_  ;
	output \g61333/_1_  ;
	output \g61334/_1_  ;
	output \g61335/_1_  ;
	output \g61336/_0_  ;
	output \g61338/_0_  ;
	output \g61339/_0_  ;
	output \g61340/_0_  ;
	output \g61377/_1_  ;
	output \g61378/_1_  ;
	output \g61379/_1_  ;
	output \g61388/_1_  ;
	output \g61391/_0_  ;
	output \g61394/_1_  ;
	output \g61395/_1_  ;
	output \g61396/_1_  ;
	output \g61398/_1_  ;
	output \g61399/_1_  ;
	output \g61421/_1_  ;
	output \g61422/_1_  ;
	output \g61423/_1_  ;
	output \g61524/_0_  ;
	output \g61525/_0_  ;
	output \g61526/_0_  ;
	output \g61527/_0_  ;
	output \g61528/_0_  ;
	output \g61529/_0_  ;
	output \g61530/_0_  ;
	output \g61531/_0_  ;
	output \g61532/_0_  ;
	output \g61533/_0_  ;
	output \g61534/_0_  ;
	output \g61535/_0_  ;
	output \g61536/_0_  ;
	output \g61537/_0_  ;
	output \g61538/_0_  ;
	output \g61539/_0_  ;
	output \g61540/_0_  ;
	output \g61541/_0_  ;
	output \g61542/_0_  ;
	output \g61543/_0_  ;
	output \g61544/_0_  ;
	output \g61545/_0_  ;
	output \g61546/_0_  ;
	output \g61547/_0_  ;
	output \g61548/_0_  ;
	output \g61549/_0_  ;
	output \g61550/_0_  ;
	output \g61551/_0_  ;
	output \g61552/_0_  ;
	output \g61553/_0_  ;
	output \g61554/_0_  ;
	output \g61555/_0_  ;
	output \g61556/_0_  ;
	output \g61557/_0_  ;
	output \g61558/_0_  ;
	output \g61559/_0_  ;
	output \g61560/_0_  ;
	output \g61561/_0_  ;
	output \g61562/_0_  ;
	output \g61563/_0_  ;
	output \g61564/_0_  ;
	output \g61565/_0_  ;
	output \g61566/_0_  ;
	output \g61620/_0_  ;
	output \g61621/_0_  ;
	output \g61622/_0_  ;
	output \g61623/_0_  ;
	output \g61753/_0_  ;
	output \g61764/_0_  ;
	output \g61786/_0_  ;
	output \g61795/_0_  ;
	output \g61801/_0_  ;
	output \g61803/_0_  ;
	output \g61808/_0_  ;
	output \g61848/_0_  ;
	output \g61850/_0_  ;
	output \g61851/_0_  ;
	output \g62097/_0_  ;
	output \g62102/_0_  ;
	output \g62115/_0_  ;
	output \g62119/_0_  ;
	output \g62130/_1_  ;
	output \g62131/_0_  ;
	output \g62132/_0_  ;
	output \g62139/_1_  ;
	output \g62140/_1_  ;
	output \g62141/_1_  ;
	output \g62144/_0_  ;
	output \g62145/_0_  ;
	output \g62146/_0_  ;
	output \g62147/_0_  ;
	output \g62150/_0_  ;
	output \g62151/_1_  ;
	output \g62152/_0_  ;
	output \g62153/_1_  ;
	output \g62156/_1_  ;
	output \g62157/_0_  ;
	output \g62159/_0_  ;
	output \g62161/_0_  ;
	output \g62187/_1_  ;
	output \g62190/_1_  ;
	output \g62191/_1_  ;
	output \g62192/_1_  ;
	output \g62194/_1_  ;
	output \g62195/_1_  ;
	output \g62196/_1_  ;
	output \g62203/_0_  ;
	output \g62204/_1_  ;
	output \g62207/_0__syn_2  ;
	output \g62208/_1_  ;
	output \g62209/_1_  ;
	output \g62210/_1_  ;
	output \g62211/_1_  ;
	output \g62212/_1_  ;
	output \g62217/_0_  ;
	output \g62286/_0_  ;
	output \g62287/_0_  ;
	output \g62288/_0_  ;
	output \g62289/_0_  ;
	output \g62290/_0_  ;
	output \g62291/_0_  ;
	output \g62292/_0_  ;
	output \g62435/_0_  ;
	output \g62436/_0_  ;
	output \g62439/_0_  ;
	output \g62456/_0_  ;
	output \g62486/_1_  ;
	output \g62492/_1_  ;
	output \g62494/_0_  ;
	output \g62495/_1_  ;
	output \g62497/_0_  ;
	output \g62537/_0_  ;
	output \g62544/_0_  ;
	output \g62546/_0_  ;
	output \g62547/_0_  ;
	output \g62549/_3_  ;
	output \g62552/_0_  ;
	output \g62554/_0_  ;
	output \g62555/_0_  ;
	output \g62556/_0_  ;
	output \g62558/_0_  ;
	output \g62559/_0_  ;
	output \g62561/_0_  ;
	output \g62562/_0_  ;
	output \g62566/_0_  ;
	output \g62567/_0_  ;
	output \g62568/_0_  ;
	output \g62569/_0_  ;
	output \g62570/_0_  ;
	output \g62571/_0_  ;
	output \g62572/_0_  ;
	output \g62573/_0_  ;
	output \g62574/_0_  ;
	output \g62575/_0_  ;
	output \g62576/_0_  ;
	output \g62577/_0_  ;
	output \g62578/_0_  ;
	output \g62579/_0_  ;
	output \g62580/_0_  ;
	output \g62581/_0_  ;
	output \g62582/_0_  ;
	output \g62583/_0_  ;
	output \g62584/_0_  ;
	output \g62585/_0_  ;
	output \g62586/_0_  ;
	output \g62587/_0_  ;
	output \g62588/_0_  ;
	output \g62589/_0_  ;
	output \g62590/_0_  ;
	output \g62591/_0_  ;
	output \g62592/_0_  ;
	output \g62593/_0_  ;
	output \g62594/_0_  ;
	output \g62595/_0_  ;
	output \g62596/_0_  ;
	output \g62597/_0_  ;
	output \g62602/_0_  ;
	output \g62607/_0_  ;
	output \g62608/_0_  ;
	output \g62609/_0_  ;
	output \g62619/_0_  ;
	output \g62620/_0_  ;
	output \g62621/_0_  ;
	output \g62622/_0_  ;
	output \g62623/_0_  ;
	output \g62624/_0_  ;
	output \g62626/_0_  ;
	output \g62627/_0_  ;
	output \g62628/_0_  ;
	output \g62629/_0_  ;
	output \g62630/_0_  ;
	output \g62631/_0_  ;
	output \g62632/_0_  ;
	output \g62633/_0_  ;
	output \g62634/_0_  ;
	output \g62635/_0_  ;
	output \g62636/_0_  ;
	output \g62637/_0_  ;
	output \g62638/_0_  ;
	output \g62639/_0_  ;
	output \g62640/_0_  ;
	output \g62641/_0_  ;
	output \g62642/_0_  ;
	output \g62643/_0_  ;
	output \g62644/_0_  ;
	output \g62645/_0_  ;
	output \g62646/_0_  ;
	output \g62647/_0_  ;
	output \g62648/_0_  ;
	output \g62649/_0_  ;
	output \g62650/_0_  ;
	output \g62651/_0_  ;
	output \g62652/_0_  ;
	output \g62653/_0_  ;
	output \g62654/_0_  ;
	output \g62655/_0_  ;
	output \g62656/_0_  ;
	output \g62657/_0_  ;
	output \g62658/_0_  ;
	output \g62659/_0_  ;
	output \g62660/_0_  ;
	output \g62661/_0_  ;
	output \g62674/_0_  ;
	output \g62682/_0_  ;
	output \g62683/_0_  ;
	output \g62689/_0_  ;
	output \g62690/_0_  ;
	output \g62691/_0_  ;
	output \g62694/_0_  ;
	output \g62695/_0_  ;
	output \g62696/_0_  ;
	output \g62698/_0_  ;
	output \g62699/_0_  ;
	output \g62700/_0_  ;
	output \g62723/_0_  ;
	output \g62724/_0_  ;
	output \g62725/_0_  ;
	output \g62726/_0_  ;
	output \g62727/_0_  ;
	output \g62728/_0_  ;
	output \g62735/_0_  ;
	output \g62736/_0_  ;
	output \g62737/_0_  ;
	output \g62738/_0_  ;
	output \g62739/_0_  ;
	output \g62740/_0_  ;
	output \g62754/_0_  ;
	output \g62762/_0_  ;
	output \g62763/_0_  ;
	output \g62764/_0_  ;
	output \g62780/_0_  ;
	output \g62781/_0_  ;
	output \g62785/_0_  ;
	output \g62786/_0_  ;
	output \g62787/_0_  ;
	output \g62791/_0_  ;
	output \g62792/_0_  ;
	output \g62794/_0_  ;
	output \g62804/_0_  ;
	output \g62806/_0_  ;
	output \g62807/_0_  ;
	output \g62811/_0_  ;
	output \g62968/_0_  ;
	output \g63005/_0_  ;
	output \g63041/_0_  ;
	output \g63116/_0_  ;
	output \g63157/_0_  ;
	output \g63164/_0_  ;
	output \g63170/_0_  ;
	output \g63189/_0_  ;
	output \g63202/_0_  ;
	output \g63206/_0_  ;
	output \g63207/_0_  ;
	output \g63265/_0_  ;
	output \g63266/_0_  ;
	output \g63269/_0_  ;
	output \g63271/_0_  ;
	output \g63272/_0_  ;
	output \g63273/_0_  ;
	output \g63274/_0_  ;
	output \g63275/_0_  ;
	output \g63276/_0_  ;
	output \g63277/_0_  ;
	output \g63278/_0_  ;
	output \g63280/_0_  ;
	output \g63281/_0_  ;
	output \g63282/_0_  ;
	output \g63283/_0_  ;
	output \g63284/_0_  ;
	output \g63285/_0_  ;
	output \g63286/_0_  ;
	output \g63287/_0_  ;
	output \g63288/_0_  ;
	output \g63289/_0_  ;
	output \g63290/_0_  ;
	output \g63292/_0_  ;
	output \g63293/_0_  ;
	output \g63294/_0_  ;
	output \g63295/_0_  ;
	output \g63296/_0_  ;
	output \g63297/_0_  ;
	output \g63298/_0_  ;
	output \g63299/_0_  ;
	output \g63302/_0_  ;
	output \g63303/_0_  ;
	output \g63304/_0_  ;
	output \g63305/_0_  ;
	output \g63306/_0_  ;
	output \g63307/_0_  ;
	output \g63308/_0_  ;
	output \g63309/_0_  ;
	output \g63310/_0_  ;
	output \g63311/_0_  ;
	output \g63312/_0_  ;
	output \g63313/_0_  ;
	output \g63314/_0_  ;
	output \g63315/_0_  ;
	output \g63316/_0_  ;
	output \g63317/_0_  ;
	output \g63318/_0_  ;
	output \g63319/_0_  ;
	output \g63320/_0_  ;
	output \g63321/_0_  ;
	output \g63322/_0_  ;
	output \g63323/_0_  ;
	output \g63324/_0_  ;
	output \g63325/_0_  ;
	output \g63326/_0_  ;
	output \g63327/_0_  ;
	output \g63328/_0_  ;
	output \g63329/_0_  ;
	output \g63330/_0_  ;
	output \g63331/_0_  ;
	output \g63339/_0_  ;
	output \g63505/_0_  ;
	output \g63525/_0_  ;
	output \g63543/_1_  ;
	output \g63602/_0_  ;
	output \g63653/_0_  ;
	output \g63663/_1_  ;
	output \g63677/_0_  ;
	output \g63694/_0_  ;
	output \g63729/_0_  ;
	output \g63766/_0_  ;
	output \g63771/_1_  ;
	output \g63773/_1_  ;
	output \g63784/_1_  ;
	output \g63964/_0_  ;
	output \g63965/_0_  ;
	output \g63966/_0_  ;
	output \g63967/_0_  ;
	output \g64257/_1_  ;
	output \g64266/_0_  ;
	output \g64275/_0_  ;
	output \g64400/_0_  ;
	output \g64416/_0_  ;
	output \g64470/_3_  ;
	output \g64473/_0_  ;
	output \g64474/_0_  ;
	output \g64475/_0_  ;
	output \g64479/_0_  ;
	output \g64480/_0_  ;
	output \g64481/_0_  ;
	output \g64483/_0_  ;
	output \g64484/_0_  ;
	output \g64485/_0_  ;
	output \g64486/_0_  ;
	output \g64493/_0_  ;
	output \g64494/_0_  ;
	output \g64495/_0_  ;
	output \g64496/_0_  ;
	output \g64505/_3_  ;
	output \g64507/_0_  ;
	output \g64508/_0_  ;
	output \g64510/_0_  ;
	output \g64511/_0_  ;
	output \g64544/_0_  ;
	output \g64545/_0_  ;
	output \g64546/_0_  ;
	output \g64639/_0_  ;
	output \g64641/_0_  ;
	output \g64642/_0_  ;
	output \g64645/_0_  ;
	output \g64650/_0_  ;
	output \g64737/_0_  ;
	output \g64738/_0_  ;
	output \g65066/_0_  ;
	output \g65070/_0_  ;
	output \g65090/_0_  ;
	output \g65102/_0_  ;
	output \g65102/_3_  ;
	output \g65126/_3_  ;
	output \g65147/_3_  ;
	output \g65163/_0_  ;
	output \g65176/_3_  ;
	output \g65178/_0_  ;
	output \g65182/_0_  ;
	output \g65190/_1_  ;
	output \g65191/_0_  ;
	output \g65196/_0_  ;
	output \g65268/_0_  ;
	output \g65275/_0_  ;
	output \g65290/_0_  ;
	output \g65290/_3_  ;
	output \g65291/_0_  ;
	output \g65292/_0_  ;
	output \g65298/_0_  ;
	output \g65298/_3_  ;
	output \g65314/_0_  ;
	output \g65314/_3_  ;
	output \g65319/_3_  ;
	output \g65335/_0_  ;
	output \g65342/_0_  ;
	output \g65348/_0_  ;
	output \g65422/_0_  ;
	output \g65465/_1_  ;
	output \g65469/_1_  ;
	output \g65478/_1_  ;
	output \g65507/_0_  ;
	output \g65548/_0_  ;
	output \g65699/_1_  ;
	output \g65713/_1_  ;
	output \g65835/_0_  ;
	output \g65860/_0_  ;
	output \g65863/_0_  ;
	output \g66094/_1_  ;
	output \g66102/_0_  ;
	output \g66107/_0_  ;
	output \g66130/_3_  ;
	output \g66131/_3_  ;
	output \g66228/_1_  ;
	output \g66348/_1_  ;
	output \g66543/_0_  ;
	output \g66549/_1_  ;
	output \g66640/_3_  ;
	output \g66641/_3_  ;
	output \g66950/_1_  ;
	output \g67111/_0_  ;
	output \g67219/_0_  ;
	output \g67263/_0_  ;
	output \g67909/_1_  ;
	output \g68049/_0_  ;
	output \g68220/_0_  ;
	output \g68413/_0_  ;
	output \g68511/_0_  ;
	output \g68536/_0_  ;
	output \g68543/_1_  ;
	output \g68554/_0_  ;
	output \g68559/_0_  ;
	output \g70915/_0_  ;
	output \g71108/_1_  ;
	output \g71115/_2_  ;
	output \g71244_dup/_0_  ;
	output \g71368/_0_  ;
	output \g71581/_0_  ;
	output \g71720/_0_  ;
	output \g785_reg/P0001  ;
	output \g789_reg/P0001  ;
	output \g797_reg/P0001  ;
	output \g809_reg/P0001  ;
	output \g813_reg/P0001  ;
	output \g966_reg/P0001  ;
	output \g968_reg/P0001  ;
	output \g970_reg/P0001  ;
	output \g972_reg/P0001  ;
	output \g974_reg/P0001  ;
	output \g976_reg/P0001  ;
	output \g978_reg/P0001  ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\g2986_reg/NET0131 ,
		\g5388_pad ,
		_w1180_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\g2987_reg/NET0131 ,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\g2478_reg/NET0131 ,
		\g7961_pad ,
		_w1182_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\g1092_reg/NET0131 ,
		\g2479_reg/NET0131 ,
		_w1183_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\g1088_reg/NET0131 ,
		\g2477_reg/NET0131 ,
		_w1184_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w1182_,
		_w1183_,
		_w1185_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\g1088_reg/NET0131 ,
		\g2220_reg/NET0131 ,
		_w1187_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\g1092_reg/NET0131 ,
		\g2222_reg/NET0131 ,
		_w1188_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\g2221_reg/NET0131 ,
		\g7961_pad ,
		_w1189_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w1187_,
		_w1188_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w1189_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\g2180_reg/NET0131 ,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\g2180_reg/NET0131 ,
		_w1191_,
		_w1193_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w1192_,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\g2233_reg/NET0131 ,
		\g7961_pad ,
		_w1195_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\g1088_reg/NET0131 ,
		\g2232_reg/NET0131 ,
		_w1196_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\g1092_reg/NET0131 ,
		\g2234_reg/NET0131 ,
		_w1197_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w1195_,
		_w1196_,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\g2200_reg/NET0131 ,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\g2200_reg/NET0131 ,
		_w1199_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w1200_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\g1088_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		_w1203_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\g1092_reg/NET0131 ,
		\g2210_reg/NET0131 ,
		_w1204_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\g2209_reg/NET0131 ,
		\g7961_pad ,
		_w1205_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w1203_,
		_w1204_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\g2170_reg/NET0131 ,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\g2170_reg/NET0131 ,
		_w1207_,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w1208_,
		_w1209_,
		_w1210_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\g2230_reg/NET0131 ,
		\g7961_pad ,
		_w1211_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\g1088_reg/NET0131 ,
		\g2229_reg/NET0131 ,
		_w1212_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\g1092_reg/NET0131 ,
		\g2231_reg/NET0131 ,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w1211_,
		_w1212_,
		_w1214_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w1213_,
		_w1214_,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\g2195_reg/NET0131 ,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\g2195_reg/NET0131 ,
		_w1215_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w1216_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\g1092_reg/NET0131 ,
		\g2252_reg/NET0131 ,
		_w1219_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\g2251_reg/NET0131 ,
		\g7961_pad ,
		_w1220_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\g1088_reg/NET0131 ,
		\g2250_reg/NET0131 ,
		_w1221_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w1219_,
		_w1220_,
		_w1222_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\g2236_reg/NET0131 ,
		\g7961_pad ,
		_w1224_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\g1088_reg/NET0131 ,
		\g2235_reg/NET0131 ,
		_w1225_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\g1092_reg/NET0131 ,
		\g2237_reg/NET0131 ,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w1224_,
		_w1225_,
		_w1227_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w1223_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w1223_,
		_w1228_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\g2224_reg/NET0131 ,
		\g7961_pad ,
		_w1232_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\g1088_reg/NET0131 ,
		\g2223_reg/NET0131 ,
		_w1233_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\g1092_reg/NET0131 ,
		\g2225_reg/NET0131 ,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w1232_,
		_w1233_,
		_w1235_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w1234_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\g2185_reg/NET0131 ,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\g2185_reg/NET0131 ,
		_w1236_,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w1237_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\g1092_reg/NET0131 ,
		\g2207_reg/NET0131 ,
		_w1240_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\g1088_reg/NET0131 ,
		\g2205_reg/NET0131 ,
		_w1241_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\g2206_reg/NET0131 ,
		\g7961_pad ,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w1240_,
		_w1241_,
		_w1243_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w1242_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\g2165_reg/NET0131 ,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\g2165_reg/NET0131 ,
		_w1244_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w1245_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\g1092_reg/NET0131 ,
		\g2219_reg/NET0131 ,
		_w1248_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\g1088_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		_w1249_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\g2218_reg/NET0131 ,
		\g7961_pad ,
		_w1250_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w1248_,
		_w1249_,
		_w1251_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w1250_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\g2175_reg/NET0131 ,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\g2175_reg/NET0131 ,
		_w1252_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w1253_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\g1088_reg/NET0131 ,
		\g2226_reg/NET0131 ,
		_w1256_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		\g2227_reg/NET0131 ,
		\g7961_pad ,
		_w1257_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\g1092_reg/NET0131 ,
		\g2228_reg/NET0131 ,
		_w1258_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w1256_,
		_w1257_,
		_w1259_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		\g2190_reg/NET0131 ,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\g2190_reg/NET0131 ,
		_w1260_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w1261_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\g1092_reg/NET0131 ,
		\g2249_reg/NET0131 ,
		_w1264_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\g2248_reg/NET0131 ,
		\g7961_pad ,
		_w1265_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\g1088_reg/NET0131 ,
		\g2247_reg/NET0131 ,
		_w1266_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w1264_,
		_w1265_,
		_w1267_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\g1088_reg/NET0131 ,
		\g2238_reg/NET0131 ,
		_w1269_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\g2239_reg/NET0131 ,
		\g7961_pad ,
		_w1270_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\g1092_reg/NET0131 ,
		\g2240_reg/NET0131 ,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w1269_,
		_w1270_,
		_w1272_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w1271_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w1268_,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w1268_,
		_w1273_,
		_w1275_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w1274_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\g1088_reg/NET0131 ,
		\g2244_reg/NET0131 ,
		_w1277_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		\g2245_reg/NET0131 ,
		\g7961_pad ,
		_w1278_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\g1092_reg/NET0131 ,
		\g2246_reg/NET0131 ,
		_w1279_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w1277_,
		_w1278_,
		_w1280_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w1279_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\g1563_reg/NET0131 ,
		_w1281_,
		_w1282_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w1194_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w1202_,
		_w1210_,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w1218_,
		_w1231_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w1239_,
		_w1247_,
		_w1286_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w1255_,
		_w1263_,
		_w1287_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w1276_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w1285_,
		_w1286_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w1283_,
		_w1284_,
		_w1290_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w1289_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w1288_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w1186_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		\g2393_reg/NET0131 ,
		\g7961_pad ,
		_w1294_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\g1088_reg/NET0131 ,
		\g2395_reg/NET0131 ,
		_w1295_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\g1092_reg/NET0131 ,
		\g2394_reg/NET0131 ,
		_w1296_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w1294_,
		_w1295_,
		_w1297_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w1296_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\g2387_reg/NET0131 ,
		\g7961_pad ,
		_w1299_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\g1092_reg/NET0131 ,
		\g2388_reg/NET0131 ,
		_w1300_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\g1088_reg/NET0131 ,
		\g2389_reg/NET0131 ,
		_w1301_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w1299_,
		_w1300_,
		_w1302_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		_w1301_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w1298_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		\g2390_reg/NET0131 ,
		\g7961_pad ,
		_w1305_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\g1088_reg/NET0131 ,
		\g2392_reg/NET0131 ,
		_w1306_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\g1092_reg/NET0131 ,
		\g2391_reg/NET0131 ,
		_w1307_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w1305_,
		_w1306_,
		_w1308_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w1307_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w1304_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		\g2397_reg/NET0131 ,
		\g7961_pad ,
		_w1311_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		\g1088_reg/NET0131 ,
		\g2396_reg/NET0131 ,
		_w1312_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\g1092_reg/NET0131 ,
		\g2398_reg/NET0131 ,
		_w1313_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w1311_,
		_w1312_,
		_w1314_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w1313_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		_w1292_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		_w1298_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\g1088_reg/NET0131 ,
		\g2348_reg/NET0131 ,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\g1092_reg/NET0131 ,
		\g2345_reg/NET0131 ,
		_w1319_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\g2342_reg/NET0131 ,
		\g7961_pad ,
		_w1320_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w1318_,
		_w1319_,
		_w1321_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		_w1268_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		_w1268_,
		_w1322_,
		_w1324_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\g2324_reg/NET0131 ,
		\g7961_pad ,
		_w1326_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\g1088_reg/NET0131 ,
		\g2330_reg/NET0131 ,
		_w1327_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\g1092_reg/NET0131 ,
		\g2327_reg/NET0131 ,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w1326_,
		_w1327_,
		_w1329_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w1328_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\g2190_reg/NET0131 ,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		\g2190_reg/NET0131 ,
		_w1330_,
		_w1332_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\g2333_reg/NET0131 ,
		\g7961_pad ,
		_w1334_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\g1088_reg/NET0131 ,
		\g2339_reg/NET0131 ,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\g1092_reg/NET0131 ,
		\g2336_reg/NET0131 ,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w1334_,
		_w1335_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w1336_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\g2200_reg/NET0131 ,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\g2200_reg/NET0131 ,
		_w1338_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w1339_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w1333_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\g1092_reg/NET0131 ,
		\g2318_reg/NET0131 ,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\g1088_reg/NET0131 ,
		\g2321_reg/NET0131 ,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\g2315_reg/NET0131 ,
		\g7961_pad ,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w1343_,
		_w1344_,
		_w1346_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w1345_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\g2180_reg/NET0131 ,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\g2180_reg/NET0131 ,
		_w1347_,
		_w1349_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\g1088_reg/NET0131 ,
		\g2312_reg/NET0131 ,
		_w1351_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\g1092_reg/NET0131 ,
		\g2309_reg/NET0131 ,
		_w1352_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\g2306_reg/NET0131 ,
		\g7961_pad ,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w1351_,
		_w1352_,
		_w1354_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\g2170_reg/NET0131 ,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\g2170_reg/NET0131 ,
		_w1355_,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		_w1350_,
		_w1358_,
		_w1359_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w1325_,
		_w1342_,
		_w1360_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w1333_,
		_w1350_,
		_w1362_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w1325_,
		_w1341_,
		_w1363_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w1358_,
		_w1362_,
		_w1364_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		_w1363_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w1325_,
		_w1350_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w1341_,
		_w1358_,
		_w1367_
	);
	LUT2 #(
		.INIT('h2)
	) name188 (
		_w1333_,
		_w1366_,
		_w1368_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w1367_,
		_w1368_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w1361_,
		_w1365_,
		_w1370_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w1369_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\g2279_reg/NET0131 ,
		\g7961_pad ,
		_w1372_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\g1092_reg/NET0131 ,
		\g2282_reg/NET0131 ,
		_w1373_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\g1088_reg/NET0131 ,
		\g2285_reg/NET0131 ,
		_w1374_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w1372_,
		_w1373_,
		_w1375_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\g2185_reg/NET0131 ,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\g2185_reg/NET0131 ,
		_w1376_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w1377_,
		_w1378_,
		_w1379_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\g1088_reg/NET0131 ,
		\g2303_reg/NET0131 ,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\g1092_reg/NET0131 ,
		\g2300_reg/NET0131 ,
		_w1381_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\g2297_reg/NET0131 ,
		\g7961_pad ,
		_w1382_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w1380_,
		_w1381_,
		_w1383_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w1382_,
		_w1383_,
		_w1384_
	);
	LUT2 #(
		.INIT('h2)
	) name205 (
		_w1223_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		_w1223_,
		_w1384_,
		_w1386_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w1385_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\g2288_reg/NET0131 ,
		\g7961_pad ,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		\g1088_reg/NET0131 ,
		\g2294_reg/NET0131 ,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		\g1092_reg/NET0131 ,
		\g2291_reg/NET0131 ,
		_w1390_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w1388_,
		_w1389_,
		_w1391_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w1390_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		\g2195_reg/NET0131 ,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\g2195_reg/NET0131 ,
		_w1392_,
		_w1394_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w1387_,
		_w1395_,
		_w1396_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\g1088_reg/NET0131 ,
		\g2276_reg/NET0131 ,
		_w1397_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\g1092_reg/NET0131 ,
		\g2273_reg/NET0131 ,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\g2270_reg/NET0131 ,
		\g7961_pad ,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w1397_,
		_w1398_,
		_w1400_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		_w1399_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		\g2175_reg/NET0131 ,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\g2175_reg/NET0131 ,
		_w1401_,
		_w1403_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\g2261_reg/NET0131 ,
		\g7961_pad ,
		_w1405_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\g1088_reg/NET0131 ,
		\g2267_reg/NET0131 ,
		_w1406_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		\g1092_reg/NET0131 ,
		\g2264_reg/NET0131 ,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w1405_,
		_w1406_,
		_w1408_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		\g2165_reg/NET0131 ,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		\g2165_reg/NET0131 ,
		_w1409_,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		_w1404_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w1325_,
		_w1379_,
		_w1414_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w1362_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w1367_,
		_w1396_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w1413_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		_w1415_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		_w1371_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		_w1298_,
		_w1419_,
		_w1420_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		_w1395_,
		_w1412_,
		_w1421_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w1387_,
		_w1404_,
		_w1422_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w1379_,
		_w1421_,
		_w1423_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w1379_,
		_w1404_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w1396_,
		_w1412_,
		_w1426_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w1379_,
		_w1395_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w1387_,
		_w1413_,
		_w1429_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w1424_,
		_w1427_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w1430_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w1316_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		_w1281_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h4)
	) name255 (
		_w1420_,
		_w1434_,
		_w1435_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		\g1563_reg/NET0131 ,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w1317_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w1303_,
		_w1437_,
		_w1438_
	);
	LUT2 #(
		.INIT('h2)
	) name259 (
		_w1309_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w1298_,
		_w1419_,
		_w1440_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		_w1432_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		_w1282_,
		_w1309_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w1303_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w1441_,
		_w1443_,
		_w1444_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w1439_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w1293_,
		_w1310_,
		_w1446_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w1445_,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		\g7961_pad ,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		\g2390_reg/NET0131 ,
		\g7961_pad ,
		_w1449_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w1448_,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		\g2984_reg/NET0131 ,
		\g2985_reg/NET0131 ,
		_w1451_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		\g3120_reg/NET0131 ,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\g3139_reg/NET0131 ,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\g2991_reg/NET0131 ,
		\g2992_reg/NET0131 ,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\g3120_reg/NET0131 ,
		_w1454_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w1453_,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		\g3114_reg/NET0131 ,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\g3097_reg/NET0131 ,
		\g3120_reg/NET0131 ,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		\g3139_reg/NET0131 ,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\g3114_reg/NET0131 ,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w1457_,
		_w1460_,
		_w1461_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		\g3230_pad ,
		\g3233_pad ,
		_w1462_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		\g3110_reg/NET0131 ,
		\g3120_reg/NET0131 ,
		_w1463_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		\g3139_reg/NET0131 ,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h4)
	) name285 (
		\g3114_reg/NET0131 ,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		_w1462_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		\g3114_reg/NET0131 ,
		_w1454_,
		_w1467_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		_w1464_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		_w1462_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\g8262_pad ,
		\g8264_pad ,
		_w1470_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		\g8262_pad ,
		\g8264_pad ,
		_w1471_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\g8260_pad ,
		\g8263_pad ,
		_w1473_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\g8260_pad ,
		\g8263_pad ,
		_w1474_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w1473_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\g8266_pad ,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		\g8266_pad ,
		_w1475_,
		_w1477_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w1476_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\g8259_pad ,
		\g8261_pad ,
		_w1479_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		\g8259_pad ,
		\g8261_pad ,
		_w1480_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		\g8265_pad ,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		\g8265_pad ,
		_w1481_,
		_w1483_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w1482_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h2)
	) name305 (
		_w1478_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		_w1478_,
		_w1484_,
		_w1486_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w1485_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		_w1472_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w1472_,
		_w1487_,
		_w1489_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w1488_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		\g2990_reg/NET0131 ,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		\g2990_reg/NET0131 ,
		_w1490_,
		_w1492_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w1491_,
		_w1492_,
		_w1493_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		\g3120_reg/NET0131 ,
		\g3231_pad ,
		_w1494_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		_w1490_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w1490_,
		_w1494_,
		_w1496_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w1495_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\g2987_reg/NET0131 ,
		\g2997_reg/NET0131 ,
		_w1498_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		\g2987_reg/NET0131 ,
		\g3061_reg/NET0131 ,
		_w1499_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w1498_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		\g8274_pad ,
		\g8275_pad ,
		_w1501_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		\g8274_pad ,
		\g8275_pad ,
		_w1502_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w1501_,
		_w1502_,
		_w1503_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		\g8270_pad ,
		\g8271_pad ,
		_w1504_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\g8270_pad ,
		\g8271_pad ,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		\g8273_pad ,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		\g8273_pad ,
		_w1506_,
		_w1508_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		\g8268_pad ,
		\g8269_pad ,
		_w1510_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		\g8268_pad ,
		\g8269_pad ,
		_w1511_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		\g8272_pad ,
		_w1512_,
		_w1513_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		\g8272_pad ,
		_w1512_,
		_w1514_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w1513_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		_w1509_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w1509_,
		_w1515_,
		_w1517_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w1516_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w1503_,
		_w1518_,
		_w1519_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w1503_,
		_w1518_,
		_w1520_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w1519_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		\g3083_reg/NET0131 ,
		_w1521_,
		_w1522_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		\g3083_reg/NET0131 ,
		_w1521_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w1522_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w1494_,
		_w1521_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w1494_,
		_w1521_,
		_w1526_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w1525_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		\g2612_reg/NET0131 ,
		\g3229_pad ,
		_w1528_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\g2574_reg/NET0131 ,
		\g2618_reg/NET0131 ,
		_w1529_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		\g1880_reg/NET0131 ,
		\g1924_reg/NET0131 ,
		_w1530_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\g1186_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w1531_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		\g499_reg/NET0131 ,
		\g544_reg/NET0131 ,
		_w1532_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		\g5657_pad ,
		_w1532_,
		_w1533_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\g1234_reg/NET0131 ,
		\g5657_pad ,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		\g1186_reg/NET0131 ,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w1533_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w1531_,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\g5657_pad ,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		\g1928_reg/NET0131 ,
		\g5657_pad ,
		_w1539_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		\g1880_reg/NET0131 ,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w1538_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w1530_,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\g5657_pad ,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		\g2622_reg/NET0131 ,
		\g5657_pad ,
		_w1544_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		\g2574_reg/NET0131 ,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w1543_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w1529_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\g2633_reg/NET0131 ,
		\g2637_pad ,
		_w1548_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		_w1547_,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w1550_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		\g2599_reg/NET0131 ,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		\g2615_reg/NET0131 ,
		\g3229_pad ,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w1528_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		_w1551_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w1549_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		\g2574_reg/NET0131 ,
		_w1549_,
		_w1556_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		\g1018_reg/NET0131 ,
		\g2798_reg/NET0131 ,
		_w1557_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		\g1024_reg/NET0131 ,
		\g2796_reg/NET0131 ,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		\g2797_reg/NET0131 ,
		\g5657_pad ,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w1557_,
		_w1558_,
		_w1560_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w1559_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\g1024_reg/NET0131 ,
		\g2793_reg/NET0131 ,
		_w1562_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\g1018_reg/NET0131 ,
		\g2795_reg/NET0131 ,
		_w1563_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		\g2794_reg/NET0131 ,
		\g5657_pad ,
		_w1564_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w1562_,
		_w1563_,
		_w1565_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w1564_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		\g1018_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		_w1567_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\g1024_reg/NET0131 ,
		\g2781_reg/NET0131 ,
		_w1568_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		\g2782_reg/NET0131 ,
		\g5657_pad ,
		_w1569_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w1567_,
		_w1568_,
		_w1570_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		\g1024_reg/NET0131 ,
		\g2772_reg/NET0131 ,
		_w1572_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		\g1018_reg/NET0131 ,
		\g2774_reg/NET0131 ,
		_w1573_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		\g2773_reg/NET0131 ,
		\g5657_pad ,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w1572_,
		_w1573_,
		_w1575_
	);
	LUT2 #(
		.INIT('h4)
	) name396 (
		_w1574_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		\g1018_reg/NET0131 ,
		\g2780_reg/NET0131 ,
		_w1577_
	);
	LUT2 #(
		.INIT('h2)
	) name398 (
		\g1024_reg/NET0131 ,
		\g2778_reg/NET0131 ,
		_w1578_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		\g2779_reg/NET0131 ,
		\g5657_pad ,
		_w1579_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w1577_,
		_w1578_,
		_w1580_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		\g1024_reg/NET0131 ,
		\g2790_reg/NET0131 ,
		_w1582_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		\g1018_reg/NET0131 ,
		\g2792_reg/NET0131 ,
		_w1583_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		\g2791_reg/NET0131 ,
		\g5657_pad ,
		_w1584_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w1582_,
		_w1583_,
		_w1585_
	);
	LUT2 #(
		.INIT('h4)
	) name406 (
		_w1584_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		\g1024_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		_w1587_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		\g1018_reg/NET0131 ,
		\g2789_reg/NET0131 ,
		_w1588_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		\g2788_reg/NET0131 ,
		\g5657_pad ,
		_w1589_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w1587_,
		_w1588_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name411 (
		_w1589_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		\g1024_reg/NET0131 ,
		\g2784_reg/NET0131 ,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\g1018_reg/NET0131 ,
		\g2786_reg/NET0131 ,
		_w1593_
	);
	LUT2 #(
		.INIT('h4)
	) name414 (
		\g2785_reg/NET0131 ,
		\g5657_pad ,
		_w1594_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w1592_,
		_w1593_,
		_w1595_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w1594_,
		_w1595_,
		_w1596_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		\g2812_reg/NET0131 ,
		\g5657_pad ,
		_w1597_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\g1024_reg/NET0131 ,
		\g2811_reg/NET0131 ,
		_w1598_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		\g1018_reg/NET0131 ,
		\g2813_reg/NET0131 ,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w1597_,
		_w1598_,
		_w1600_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		\g2806_reg/NET0131 ,
		\g5657_pad ,
		_w1602_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		\g1018_reg/NET0131 ,
		\g2807_reg/NET0131 ,
		_w1603_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		\g1024_reg/NET0131 ,
		\g2805_reg/NET0131 ,
		_w1604_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w1602_,
		_w1603_,
		_w1605_
	);
	LUT2 #(
		.INIT('h4)
	) name426 (
		_w1604_,
		_w1605_,
		_w1606_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		\g1018_reg/NET0131 ,
		\g2801_reg/NET0131 ,
		_w1607_
	);
	LUT2 #(
		.INIT('h2)
	) name428 (
		\g1024_reg/NET0131 ,
		\g2799_reg/NET0131 ,
		_w1608_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		\g2800_reg/NET0131 ,
		\g5657_pad ,
		_w1609_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w1607_,
		_w1608_,
		_w1610_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		\g1024_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		_w1612_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		\g1018_reg/NET0131 ,
		\g2777_reg/NET0131 ,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name434 (
		\g2776_reg/NET0131 ,
		\g5657_pad ,
		_w1614_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w1612_,
		_w1613_,
		_w1615_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		_w1614_,
		_w1615_,
		_w1616_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w1561_,
		_w1566_,
		_w1617_
	);
	LUT2 #(
		.INIT('h4)
	) name438 (
		_w1571_,
		_w1576_,
		_w1618_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w1581_,
		_w1586_,
		_w1619_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w1591_,
		_w1596_,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w1601_,
		_w1606_,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w1611_,
		_w1616_,
		_w1622_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w1621_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w1619_,
		_w1620_,
		_w1624_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		_w1617_,
		_w1618_,
		_w1625_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		_w1624_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w1623_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w1561_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		\g1024_reg/NET0131 ,
		\g2694_reg/NET0131 ,
		_w1629_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\g1018_reg/NET0131 ,
		\g2691_reg/NET0131 ,
		_w1630_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		\g2688_reg/NET0131 ,
		\g5657_pad ,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w1629_,
		_w1630_,
		_w1632_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w1628_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w1628_,
		_w1633_,
		_w1635_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w1634_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w1556_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w1611_,
		_w1627_,
		_w1638_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		\g1024_reg/NET0131 ,
		\g2685_reg/NET0131 ,
		_w1639_
	);
	LUT2 #(
		.INIT('h8)
	) name460 (
		\g1018_reg/NET0131 ,
		\g2682_reg/NET0131 ,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		\g2679_reg/NET0131 ,
		\g5657_pad ,
		_w1641_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w1639_,
		_w1640_,
		_w1642_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		_w1641_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w1638_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		_w1638_,
		_w1643_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w1556_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w1637_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		_w1637_,
		_w1646_,
		_w1649_
	);
	LUT2 #(
		.INIT('h2)
	) name470 (
		\g1243_reg/NET0131 ,
		_w1648_,
		_w1650_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		_w1649_,
		_w1650_,
		_w1651_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		_w1586_,
		_w1633_,
		_w1652_
	);
	LUT2 #(
		.INIT('h2)
	) name473 (
		_w1586_,
		_w1633_,
		_w1653_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w1652_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w1556_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h2)
	) name476 (
		_w1566_,
		_w1643_,
		_w1656_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		_w1566_,
		_w1643_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w1556_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		_w1596_,
		_w1633_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		_w1596_,
		_w1633_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		_w1659_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		_w1556_,
		_w1662_,
		_w1664_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w1658_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w1663_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		_w1591_,
		_w1643_,
		_w1667_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		_w1591_,
		_w1643_,
		_w1668_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w1667_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		_w1556_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		_w1666_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('h4)
	) name492 (
		_w1666_,
		_w1670_,
		_w1672_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w1671_,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w1655_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		_w1655_,
		_w1673_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w1674_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w1616_,
		_w1627_,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w1643_,
		_w1677_,
		_w1678_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		_w1643_,
		_w1677_,
		_w1679_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w1678_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w1556_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w1581_,
		_w1627_,
		_w1682_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w1633_,
		_w1682_,
		_w1683_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		_w1633_,
		_w1682_,
		_w1684_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w1683_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h2)
	) name506 (
		_w1556_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w1571_,
		_w1627_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name508 (
		_w1643_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h2)
	) name509 (
		_w1643_,
		_w1687_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		_w1688_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		_w1686_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		_w1556_,
		_w1690_,
		_w1692_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		_w1685_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w1691_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		_w1576_,
		_w1633_,
		_w1695_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		_w1576_,
		_w1633_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		_w1556_,
		_w1697_,
		_w1698_
	);
	LUT2 #(
		.INIT('h2)
	) name519 (
		_w1694_,
		_w1698_,
		_w1699_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		_w1694_,
		_w1698_,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w1699_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w1681_,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w1681_,
		_w1701_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w1676_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		_w1676_,
		_w1704_,
		_w1706_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		\g1196_reg/NET0131 ,
		_w1705_,
		_w1707_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		_w1706_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w1555_,
		_w1651_,
		_w1709_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		\g2987_reg/NET0131 ,
		\g3070_reg/NET0131 ,
		_w1711_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		\g2987_reg/NET0131 ,
		\g3051_reg/NET0131 ,
		_w1712_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		\g2987_reg/NET0131 ,
		\g3078_reg/NET0131 ,
		_w1714_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		\g2987_reg/NET0131 ,
		\g3060_reg/NET0131 ,
		_w1715_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w1714_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		\g2987_reg/NET0131 ,
		\g3075_reg/NET0131 ,
		_w1717_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		\g2987_reg/NET0131 ,
		\g3057_reg/NET0131 ,
		_w1718_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		_w1717_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		\g2987_reg/NET0131 ,
		\g3076_reg/NET0131 ,
		_w1720_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		\g2987_reg/NET0131 ,
		\g3058_reg/NET0131 ,
		_w1721_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w1720_,
		_w1721_,
		_w1722_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		\g2987_reg/NET0131 ,
		\g3072_reg/NET0131 ,
		_w1723_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		\g2987_reg/NET0131 ,
		\g3053_reg/NET0131 ,
		_w1724_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		_w1723_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\g2987_reg/NET0131 ,
		\g3077_reg/NET0131 ,
		_w1726_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		\g2987_reg/NET0131 ,
		\g3059_reg/NET0131 ,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w1726_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\g2987_reg/NET0131 ,
		\g3074_reg/NET0131 ,
		_w1729_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		\g2987_reg/NET0131 ,
		\g3056_reg/NET0131 ,
		_w1730_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w1729_,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		\g2987_reg/NET0131 ,
		\g3071_reg/NET0131 ,
		_w1732_
	);
	LUT2 #(
		.INIT('h4)
	) name553 (
		\g2987_reg/NET0131 ,
		\g3052_reg/NET0131 ,
		_w1733_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w1732_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name555 (
		\g2987_reg/NET0131 ,
		\g3073_reg/NET0131 ,
		_w1735_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		\g2987_reg/NET0131 ,
		\g3055_reg/NET0131 ,
		_w1736_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w1735_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		\g1939_reg/NET0131 ,
		\g1943_pad ,
		_w1738_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w1542_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		\g1880_reg/NET0131 ,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		\g1994_reg/NET0131 ,
		\g5657_pad ,
		_w1741_
	);
	LUT2 #(
		.INIT('h8)
	) name562 (
		\g1018_reg/NET0131 ,
		\g1997_reg/NET0131 ,
		_w1742_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		\g1024_reg/NET0131 ,
		\g2000_reg/NET0131 ,
		_w1743_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w1741_,
		_w1742_,
		_w1744_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w1743_,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		\g1024_reg/NET0131 ,
		\g2102_reg/NET0131 ,
		_w1746_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		\g1018_reg/NET0131 ,
		\g2104_reg/NET0131 ,
		_w1747_
	);
	LUT2 #(
		.INIT('h4)
	) name568 (
		\g2103_reg/NET0131 ,
		\g5657_pad ,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w1746_,
		_w1747_,
		_w1749_
	);
	LUT2 #(
		.INIT('h4)
	) name570 (
		_w1748_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		\g1018_reg/NET0131 ,
		\g2095_reg/NET0131 ,
		_w1751_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		\g1024_reg/NET0131 ,
		\g2093_reg/NET0131 ,
		_w1752_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		\g2094_reg/NET0131 ,
		\g5657_pad ,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w1751_,
		_w1752_,
		_w1754_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w1753_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		\g1024_reg/NET0131 ,
		\g2078_reg/NET0131 ,
		_w1756_
	);
	LUT2 #(
		.INIT('h2)
	) name577 (
		\g1018_reg/NET0131 ,
		\g2080_reg/NET0131 ,
		_w1757_
	);
	LUT2 #(
		.INIT('h4)
	) name578 (
		\g2079_reg/NET0131 ,
		\g5657_pad ,
		_w1758_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w1756_,
		_w1757_,
		_w1759_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name581 (
		\g1018_reg/NET0131 ,
		\g2092_reg/NET0131 ,
		_w1761_
	);
	LUT2 #(
		.INIT('h2)
	) name582 (
		\g1024_reg/NET0131 ,
		\g2090_reg/NET0131 ,
		_w1762_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		\g2091_reg/NET0131 ,
		\g5657_pad ,
		_w1763_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w1761_,
		_w1762_,
		_w1764_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\g1018_reg/NET0131 ,
		\g2083_reg/NET0131 ,
		_w1766_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		\g1024_reg/NET0131 ,
		\g2081_reg/NET0131 ,
		_w1767_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		\g2082_reg/NET0131 ,
		\g5657_pad ,
		_w1768_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w1766_,
		_w1767_,
		_w1769_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		_w1768_,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		\g1024_reg/NET0131 ,
		\g2087_reg/NET0131 ,
		_w1771_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		\g1018_reg/NET0131 ,
		\g2089_reg/NET0131 ,
		_w1772_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		\g2088_reg/NET0131 ,
		\g5657_pad ,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		_w1771_,
		_w1772_,
		_w1774_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w1773_,
		_w1774_,
		_w1775_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		\g1018_reg/NET0131 ,
		\g2086_reg/NET0131 ,
		_w1776_
	);
	LUT2 #(
		.INIT('h2)
	) name597 (
		\g1024_reg/NET0131 ,
		\g2084_reg/NET0131 ,
		_w1777_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		\g2085_reg/NET0131 ,
		\g5657_pad ,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		_w1776_,
		_w1777_,
		_w1779_
	);
	LUT2 #(
		.INIT('h4)
	) name600 (
		_w1778_,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		\g1018_reg/NET0131 ,
		\g2107_reg/NET0131 ,
		_w1781_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		\g1024_reg/NET0131 ,
		\g2105_reg/NET0131 ,
		_w1782_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		\g2106_reg/NET0131 ,
		\g5657_pad ,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w1781_,
		_w1782_,
		_w1784_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w1783_,
		_w1784_,
		_w1785_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		\g1024_reg/NET0131 ,
		\g2099_reg/NET0131 ,
		_w1786_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		\g1018_reg/NET0131 ,
		\g2101_reg/NET0131 ,
		_w1787_
	);
	LUT2 #(
		.INIT('h4)
	) name608 (
		\g2100_reg/NET0131 ,
		\g5657_pad ,
		_w1788_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w1786_,
		_w1787_,
		_w1789_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w1788_,
		_w1789_,
		_w1790_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		\g2112_reg/NET0131 ,
		\g5657_pad ,
		_w1791_
	);
	LUT2 #(
		.INIT('h2)
	) name612 (
		\g1018_reg/NET0131 ,
		\g2113_reg/NET0131 ,
		_w1792_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		\g1024_reg/NET0131 ,
		\g2111_reg/NET0131 ,
		_w1793_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w1791_,
		_w1792_,
		_w1794_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w1793_,
		_w1794_,
		_w1795_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		\g1018_reg/NET0131 ,
		\g2098_reg/NET0131 ,
		_w1796_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		\g1024_reg/NET0131 ,
		\g2096_reg/NET0131 ,
		_w1797_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		\g2097_reg/NET0131 ,
		\g5657_pad ,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w1796_,
		_w1797_,
		_w1799_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w1798_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h2)
	) name621 (
		\g1024_reg/NET0131 ,
		\g2117_reg/NET0131 ,
		_w1801_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		\g2118_reg/NET0131 ,
		\g5657_pad ,
		_w1802_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		\g1018_reg/NET0131 ,
		\g2119_reg/NET0131 ,
		_w1803_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w1801_,
		_w1802_,
		_w1804_
	);
	LUT2 #(
		.INIT('h4)
	) name625 (
		_w1803_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		_w1750_,
		_w1755_,
		_w1806_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		_w1760_,
		_w1765_,
		_w1807_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w1770_,
		_w1775_,
		_w1808_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w1780_,
		_w1785_,
		_w1809_
	);
	LUT2 #(
		.INIT('h2)
	) name630 (
		_w1790_,
		_w1795_,
		_w1810_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		_w1800_,
		_w1805_,
		_w1811_
	);
	LUT2 #(
		.INIT('h8)
	) name632 (
		_w1810_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		_w1808_,
		_w1809_,
		_w1813_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		_w1806_,
		_w1807_,
		_w1814_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		_w1813_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		_w1812_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		_w1750_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w1745_,
		_w1817_,
		_w1818_
	);
	LUT2 #(
		.INIT('h2)
	) name639 (
		_w1745_,
		_w1817_,
		_w1819_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		_w1818_,
		_w1819_,
		_w1820_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w1740_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		\g1985_reg/NET0131 ,
		\g5657_pad ,
		_w1822_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\g1024_reg/NET0131 ,
		\g1991_reg/NET0131 ,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		\g1018_reg/NET0131 ,
		\g1988_reg/NET0131 ,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w1822_,
		_w1823_,
		_w1825_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w1824_,
		_w1825_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w1785_,
		_w1816_,
		_w1827_
	);
	LUT2 #(
		.INIT('h4)
	) name648 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		_w1826_,
		_w1827_,
		_w1829_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w1828_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		_w1821_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		_w1740_,
		_w1830_,
		_w1832_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		_w1820_,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w1831_,
		_w1833_,
		_w1834_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		\g1243_reg/NET0131 ,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h4)
	) name656 (
		\g1918_reg/NET0131 ,
		\g3229_pad ,
		_w1836_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		\g1905_reg/NET0131 ,
		_w1550_,
		_w1837_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		\g1921_reg/NET0131 ,
		\g3229_pad ,
		_w1838_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w1836_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		_w1837_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w1739_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w1775_,
		_w1816_,
		_w1842_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		_w1826_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w1826_,
		_w1842_,
		_w1844_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		_w1843_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h2)
	) name666 (
		_w1740_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w1780_,
		_w1816_,
		_w1847_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		_w1745_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name669 (
		_w1745_,
		_w1847_,
		_w1849_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w1848_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w1846_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		_w1740_,
		_w1850_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		_w1845_,
		_w1852_,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w1851_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h2)
	) name675 (
		_w1745_,
		_w1760_,
		_w1855_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		_w1745_,
		_w1760_,
		_w1856_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w1855_,
		_w1856_,
		_w1857_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		_w1740_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		_w1854_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w1854_,
		_w1858_,
		_w1860_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w1859_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w1770_,
		_w1816_,
		_w1862_
	);
	LUT2 #(
		.INIT('h4)
	) name683 (
		_w1826_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		_w1826_,
		_w1862_,
		_w1864_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		_w1740_,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w1745_,
		_w1800_,
		_w1867_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		_w1745_,
		_w1800_,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w1867_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w1866_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		_w1740_,
		_w1869_,
		_w1871_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		_w1865_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w1870_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h2)
	) name694 (
		_w1745_,
		_w1765_,
		_w1874_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		_w1745_,
		_w1765_,
		_w1875_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w1874_,
		_w1875_,
		_w1876_
	);
	LUT2 #(
		.INIT('h8)
	) name697 (
		_w1740_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w1755_,
		_w1826_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		_w1755_,
		_w1826_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name700 (
		_w1878_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		_w1877_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		_w1740_,
		_w1880_,
		_w1882_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		_w1876_,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w1881_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		_w1790_,
		_w1826_,
		_w1885_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		_w1790_,
		_w1826_,
		_w1886_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w1885_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w1740_,
		_w1887_,
		_w1888_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		_w1884_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w1884_,
		_w1888_,
		_w1890_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w1889_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w1873_,
		_w1891_,
		_w1892_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w1873_,
		_w1891_,
		_w1893_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w1892_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h2)
	) name715 (
		_w1861_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h4)
	) name716 (
		_w1861_,
		_w1894_,
		_w1896_
	);
	LUT2 #(
		.INIT('h2)
	) name717 (
		\g1196_reg/NET0131 ,
		_w1895_,
		_w1897_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		_w1896_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w1835_,
		_w1841_,
		_w1899_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h4)
	) name721 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w1901_
	);
	LUT2 #(
		.INIT('h2)
	) name722 (
		\g1018_reg/NET0131 ,
		\g2810_reg/NET0131 ,
		_w1902_
	);
	LUT2 #(
		.INIT('h2)
	) name723 (
		\g1024_reg/NET0131 ,
		\g2808_reg/NET0131 ,
		_w1903_
	);
	LUT2 #(
		.INIT('h4)
	) name724 (
		\g2809_reg/NET0131 ,
		\g5657_pad ,
		_w1904_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w1902_,
		_w1903_,
		_w1905_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		_w1904_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h4)
	) name727 (
		_w1627_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		\g2574_reg/NET0131 ,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		_w1549_,
		_w1908_,
		_w1909_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		_w1901_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w1911_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w1551_,
		_w1911_,
		_w1912_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		_w1551_,
		_w1659_,
		_w1913_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w1551_,
		_w1901_,
		_w1914_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		\g2603_reg/NET0131 ,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		_w1549_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w1912_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w1913_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w1910_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h4)
	) name740 (
		_w1551_,
		_w1664_,
		_w1920_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		\g2606_reg/NET0131 ,
		_w1914_,
		_w1921_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		_w1549_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w1912_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h4)
	) name744 (
		_w1920_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		_w1910_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w1549_,
		_w1901_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name747 (
		_w1692_,
		_w1914_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		\g2607_reg/NET0131 ,
		_w1914_,
		_w1928_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		_w1549_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w1912_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		_w1927_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w1926_,
		_w1931_,
		_w1932_
	);
	LUT2 #(
		.INIT('h2)
	) name753 (
		_w1549_,
		_w1908_,
		_w1933_
	);
	LUT2 #(
		.INIT('h2)
	) name754 (
		_w1901_,
		_w1933_,
		_w1934_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		\g2605_reg/NET0131 ,
		_w1914_,
		_w1935_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		_w1549_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w1551_,
		_w1670_,
		_w1937_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w1912_,
		_w1936_,
		_w1938_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		_w1937_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w1934_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h8)
	) name761 (
		_w1686_,
		_w1914_,
		_w1941_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		\g2608_reg/NET0131 ,
		_w1914_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		_w1549_,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w1912_,
		_w1943_,
		_w1944_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		_w1941_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		_w1926_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		\g2604_reg/NET0131 ,
		_w1914_,
		_w1947_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		_w1549_,
		_w1947_,
		_w1948_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		_w1551_,
		_w1655_,
		_w1949_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w1912_,
		_w1948_,
		_w1950_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w1934_,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w1647_,
		_w1901_,
		_w1953_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w1551_,
		_w1681_,
		_w1954_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		\g2610_reg/NET0131 ,
		_w1914_,
		_w1955_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		_w1549_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w1912_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		_w1954_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		_w1953_,
		_w1958_,
		_w1959_
	);
	LUT2 #(
		.INIT('h4)
	) name780 (
		_w1637_,
		_w1901_,
		_w1960_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w1551_,
		_w1698_,
		_w1961_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		\g2611_reg/NET0131 ,
		_w1914_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		_w1549_,
		_w1962_,
		_w1963_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w1912_,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h4)
	) name785 (
		_w1961_,
		_w1964_,
		_w1965_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		_w1960_,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		\g2987_reg/NET0131 ,
		\g3067_reg/NET0131 ,
		_w1967_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		\g2987_reg/NET0131 ,
		\g3048_reg/NET0131 ,
		_w1968_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w1967_,
		_w1968_,
		_w1969_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		\g2987_reg/NET0131 ,
		\g3068_reg/NET0131 ,
		_w1970_
	);
	LUT2 #(
		.INIT('h4)
	) name791 (
		\g2987_reg/NET0131 ,
		\g3049_reg/NET0131 ,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w1970_,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		\g2987_reg/NET0131 ,
		\g3069_reg/NET0131 ,
		_w1973_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		\g2987_reg/NET0131 ,
		\g3050_reg/NET0131 ,
		_w1974_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		\g2987_reg/NET0131 ,
		\g3065_reg/NET0131 ,
		_w1976_
	);
	LUT2 #(
		.INIT('h4)
	) name797 (
		\g2987_reg/NET0131 ,
		\g3046_reg/NET0131 ,
		_w1977_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		_w1976_,
		_w1977_,
		_w1978_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		\g2987_reg/NET0131 ,
		\g3064_reg/NET0131 ,
		_w1979_
	);
	LUT2 #(
		.INIT('h4)
	) name800 (
		\g2987_reg/NET0131 ,
		\g3045_reg/NET0131 ,
		_w1980_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w1979_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\g2987_reg/NET0131 ,
		\g3063_reg/NET0131 ,
		_w1982_
	);
	LUT2 #(
		.INIT('h4)
	) name803 (
		\g2987_reg/NET0131 ,
		\g3044_reg/NET0131 ,
		_w1983_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w1982_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		\g2987_reg/NET0131 ,
		\g3062_reg/NET0131 ,
		_w1985_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		\g2987_reg/NET0131 ,
		\g3043_reg/NET0131 ,
		_w1986_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w1985_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\g2987_reg/NET0131 ,
		\g3066_reg/NET0131 ,
		_w1988_
	);
	LUT2 #(
		.INIT('h4)
	) name809 (
		\g2987_reg/NET0131 ,
		\g3047_reg/NET0131 ,
		_w1989_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w1988_,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		\g2373_reg/NET0131 ,
		\g2374_reg/NET0131 ,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		\g1092_reg/NET0131 ,
		\g2380_reg/NET0131 ,
		_w1992_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		\g1679_reg/NET0131 ,
		\g1680_reg/NET0131 ,
		_w1993_
	);
	LUT2 #(
		.INIT('h1)
	) name814 (
		\g1092_reg/NET0131 ,
		\g1686_reg/NET0131 ,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		\g985_reg/NET0131 ,
		\g986_reg/NET0131 ,
		_w1995_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		\g1092_reg/NET0131 ,
		\g992_reg/NET0131 ,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		\g298_reg/NET0131 ,
		\g299_reg/NET0131 ,
		_w1997_
	);
	LUT2 #(
		.INIT('h2)
	) name818 (
		\g1092_reg/NET0131 ,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		\g986_reg/NET0131 ,
		_w1996_,
		_w1999_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		_w1998_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w1995_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		\g1092_reg/NET0131 ,
		_w2001_,
		_w2002_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		\g1680_reg/NET0131 ,
		_w1994_,
		_w2003_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		_w2002_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		_w1993_,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h8)
	) name826 (
		\g1092_reg/NET0131 ,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		\g2374_reg/NET0131 ,
		_w1992_,
		_w2007_
	);
	LUT2 #(
		.INIT('h4)
	) name828 (
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1991_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h2)
	) name830 (
		\g1088_reg/NET0131 ,
		\g317_reg/NET0131 ,
		_w2010_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		\g1092_reg/NET0131 ,
		\g316_reg/NET0131 ,
		_w2011_
	);
	LUT2 #(
		.INIT('h4)
	) name832 (
		\g315_reg/NET0131 ,
		\g7961_pad ,
		_w2012_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w2010_,
		_w2011_,
		_w2013_
	);
	LUT2 #(
		.INIT('h4)
	) name834 (
		_w2012_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		\g312_reg/NET0131 ,
		\g7961_pad ,
		_w2015_
	);
	LUT2 #(
		.INIT('h2)
	) name836 (
		\g1092_reg/NET0131 ,
		\g313_reg/NET0131 ,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		\g1088_reg/NET0131 ,
		\g314_reg/NET0131 ,
		_w2017_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w2015_,
		_w2016_,
		_w2018_
	);
	LUT2 #(
		.INIT('h4)
	) name839 (
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		\g318_reg/NET0131 ,
		\g7961_pad ,
		_w2020_
	);
	LUT2 #(
		.INIT('h2)
	) name841 (
		\g1092_reg/NET0131 ,
		\g319_reg/NET0131 ,
		_w2021_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		\g1088_reg/NET0131 ,
		\g320_reg/NET0131 ,
		_w2022_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w2020_,
		_w2021_,
		_w2023_
	);
	LUT2 #(
		.INIT('h4)
	) name844 (
		_w2022_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		\g1092_reg/NET0131 ,
		\g323_reg/NET0131 ,
		_w2025_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		\g322_reg/NET0131 ,
		\g7961_pad ,
		_w2026_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		\g1088_reg/NET0131 ,
		\g321_reg/NET0131 ,
		_w2027_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w2025_,
		_w2026_,
		_w2028_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w2027_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		\g1092_reg/NET0131 ,
		\g173_reg/NET0131 ,
		_w2030_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		\g172_reg/NET0131 ,
		\g7961_pad ,
		_w2031_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		\g1088_reg/NET0131 ,
		\g171_reg/NET0131 ,
		_w2032_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w2030_,
		_w2031_,
		_w2033_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		_w2032_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h2)
	) name855 (
		\g1092_reg/NET0131 ,
		\g164_reg/NET0131 ,
		_w2035_
	);
	LUT2 #(
		.INIT('h2)
	) name856 (
		\g1088_reg/NET0131 ,
		\g162_reg/NET0131 ,
		_w2036_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		\g163_reg/NET0131 ,
		\g7961_pad ,
		_w2037_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		_w2035_,
		_w2036_,
		_w2038_
	);
	LUT2 #(
		.INIT('h4)
	) name859 (
		_w2037_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w2034_,
		_w2039_,
		_w2040_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		_w2034_,
		_w2039_,
		_w2041_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w2040_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h2)
	) name863 (
		\g1092_reg/NET0131 ,
		\g176_reg/NET0131 ,
		_w2043_
	);
	LUT2 #(
		.INIT('h4)
	) name864 (
		\g175_reg/NET0131 ,
		\g7961_pad ,
		_w2044_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		\g1088_reg/NET0131 ,
		\g174_reg/NET0131 ,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		_w2043_,
		_w2044_,
		_w2046_
	);
	LUT2 #(
		.INIT('h4)
	) name867 (
		_w2045_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h2)
	) name868 (
		\g1088_reg/NET0131 ,
		\g159_reg/NET0131 ,
		_w2048_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		\g160_reg/NET0131 ,
		\g7961_pad ,
		_w2049_
	);
	LUT2 #(
		.INIT('h2)
	) name870 (
		\g1092_reg/NET0131 ,
		\g161_reg/NET0131 ,
		_w2050_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w2048_,
		_w2049_,
		_w2051_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w2050_,
		_w2051_,
		_w2052_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		_w2047_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		_w2047_,
		_w2052_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		_w2053_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		\g1092_reg/NET0131 ,
		\g131_reg/NET0131 ,
		_w2056_
	);
	LUT2 #(
		.INIT('h2)
	) name877 (
		\g1088_reg/NET0131 ,
		\g129_reg/NET0131 ,
		_w2057_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		\g130_reg/NET0131 ,
		\g7961_pad ,
		_w2058_
	);
	LUT2 #(
		.INIT('h1)
	) name879 (
		_w2056_,
		_w2057_,
		_w2059_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		_w2058_,
		_w2059_,
		_w2060_
	);
	LUT2 #(
		.INIT('h2)
	) name881 (
		\g97_reg/NET0131 ,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		\g97_reg/NET0131 ,
		_w2060_,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w2061_,
		_w2062_,
		_w2063_
	);
	LUT2 #(
		.INIT('h2)
	) name884 (
		\g1088_reg/NET0131 ,
		\g153_reg/NET0131 ,
		_w2064_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		\g154_reg/NET0131 ,
		\g7961_pad ,
		_w2065_
	);
	LUT2 #(
		.INIT('h2)
	) name886 (
		\g1092_reg/NET0131 ,
		\g155_reg/NET0131 ,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w2064_,
		_w2065_,
		_w2067_
	);
	LUT2 #(
		.INIT('h4)
	) name888 (
		_w2066_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		\g121_reg/NET0131 ,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		\g121_reg/NET0131 ,
		_w2068_,
		_w2070_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w2069_,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('h2)
	) name892 (
		\g1088_reg/NET0131 ,
		\g147_reg/NET0131 ,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		\g1092_reg/NET0131 ,
		\g149_reg/NET0131 ,
		_w2073_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		\g148_reg/NET0131 ,
		\g7961_pad ,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w2072_,
		_w2073_,
		_w2075_
	);
	LUT2 #(
		.INIT('h4)
	) name896 (
		_w2074_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h2)
	) name897 (
		\g113_reg/NET0131 ,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h4)
	) name898 (
		\g113_reg/NET0131 ,
		_w2076_,
		_w2078_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w2077_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		\g1088_reg/NET0131 ,
		\g150_reg/NET0131 ,
		_w2080_
	);
	LUT2 #(
		.INIT('h4)
	) name901 (
		\g151_reg/NET0131 ,
		\g7961_pad ,
		_w2081_
	);
	LUT2 #(
		.INIT('h2)
	) name902 (
		\g1092_reg/NET0131 ,
		\g152_reg/NET0131 ,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w2080_,
		_w2081_,
		_w2083_
	);
	LUT2 #(
		.INIT('h4)
	) name904 (
		_w2082_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\g117_reg/NET0131 ,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h4)
	) name906 (
		\g117_reg/NET0131 ,
		_w2084_,
		_w2086_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w2085_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h2)
	) name908 (
		\g1092_reg/NET0131 ,
		\g143_reg/NET0131 ,
		_w2088_
	);
	LUT2 #(
		.INIT('h2)
	) name909 (
		\g1088_reg/NET0131 ,
		\g141_reg/NET0131 ,
		_w2089_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		\g142_reg/NET0131 ,
		\g7961_pad ,
		_w2090_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w2088_,
		_w2089_,
		_w2091_
	);
	LUT2 #(
		.INIT('h4)
	) name912 (
		_w2090_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h2)
	) name913 (
		\g105_reg/NET0131 ,
		_w2092_,
		_w2093_
	);
	LUT2 #(
		.INIT('h4)
	) name914 (
		\g105_reg/NET0131 ,
		_w2092_,
		_w2094_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w2093_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		\g1092_reg/NET0131 ,
		\g158_reg/NET0131 ,
		_w2096_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		\g157_reg/NET0131 ,
		\g7961_pad ,
		_w2097_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		\g1088_reg/NET0131 ,
		\g156_reg/NET0131 ,
		_w2098_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w2096_,
		_w2097_,
		_w2099_
	);
	LUT2 #(
		.INIT('h4)
	) name920 (
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h2)
	) name921 (
		\g125_reg/NET0131 ,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h4)
	) name922 (
		\g125_reg/NET0131 ,
		_w2100_,
		_w2102_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w2101_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h2)
	) name924 (
		\g1092_reg/NET0131 ,
		\g134_reg/NET0131 ,
		_w2104_
	);
	LUT2 #(
		.INIT('h2)
	) name925 (
		\g1088_reg/NET0131 ,
		\g132_reg/NET0131 ,
		_w2105_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		\g133_reg/NET0131 ,
		\g7961_pad ,
		_w2106_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w2104_,
		_w2105_,
		_w2107_
	);
	LUT2 #(
		.INIT('h4)
	) name928 (
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		\g101_reg/NET0131 ,
		_w2108_,
		_w2109_
	);
	LUT2 #(
		.INIT('h2)
	) name930 (
		\g101_reg/NET0131 ,
		_w2108_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name931 (
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h2)
	) name932 (
		\g1092_reg/NET0131 ,
		\g170_reg/NET0131 ,
		_w2112_
	);
	LUT2 #(
		.INIT('h4)
	) name933 (
		\g169_reg/NET0131 ,
		\g7961_pad ,
		_w2113_
	);
	LUT2 #(
		.INIT('h2)
	) name934 (
		\g1088_reg/NET0131 ,
		\g168_reg/NET0131 ,
		_w2114_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		_w2112_,
		_w2113_,
		_w2115_
	);
	LUT2 #(
		.INIT('h4)
	) name936 (
		_w2114_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h2)
	) name937 (
		\g1563_reg/NET0131 ,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		\g1092_reg/NET0131 ,
		\g146_reg/NET0131 ,
		_w2118_
	);
	LUT2 #(
		.INIT('h4)
	) name939 (
		\g145_reg/NET0131 ,
		\g7961_pad ,
		_w2119_
	);
	LUT2 #(
		.INIT('h2)
	) name940 (
		\g1088_reg/NET0131 ,
		\g144_reg/NET0131 ,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name941 (
		_w2118_,
		_w2119_,
		_w2121_
	);
	LUT2 #(
		.INIT('h4)
	) name942 (
		_w2120_,
		_w2121_,
		_w2122_
	);
	LUT2 #(
		.INIT('h2)
	) name943 (
		\g109_reg/NET0131 ,
		_w2122_,
		_w2123_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		\g109_reg/NET0131 ,
		_w2122_,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w2123_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		_w2042_,
		_w2117_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w2055_,
		_w2063_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w2071_,
		_w2079_,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w2087_,
		_w2095_,
		_w2129_
	);
	LUT2 #(
		.INIT('h1)
	) name950 (
		_w2103_,
		_w2111_,
		_w2130_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w2125_,
		_w2130_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		_w2128_,
		_w2129_,
		_w2132_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		_w2126_,
		_w2127_,
		_w2133_
	);
	LUT2 #(
		.INIT('h8)
	) name954 (
		_w2132_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h8)
	) name955 (
		_w2131_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		_w2029_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h4)
	) name957 (
		_w2024_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		\g1088_reg/NET0131 ,
		\g273_reg/NET0131 ,
		_w2138_
	);
	LUT2 #(
		.INIT('h8)
	) name959 (
		\g1092_reg/NET0131 ,
		\g270_reg/NET0131 ,
		_w2139_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		\g267_reg/NET0131 ,
		\g7961_pad ,
		_w2140_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		_w2138_,
		_w2139_,
		_w2141_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT2 #(
		.INIT('h2)
	) name963 (
		_w2034_,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h4)
	) name964 (
		_w2034_,
		_w2142_,
		_w2144_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w2143_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		\g1092_reg/NET0131 ,
		\g261_reg/NET0131 ,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		\g1088_reg/NET0131 ,
		\g264_reg/NET0131 ,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		\g258_reg/NET0131 ,
		\g7961_pad ,
		_w2148_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		_w2146_,
		_w2147_,
		_w2149_
	);
	LUT2 #(
		.INIT('h4)
	) name970 (
		_w2148_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h2)
	) name971 (
		\g125_reg/NET0131 ,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h4)
	) name972 (
		\g125_reg/NET0131 ,
		_w2150_,
		_w2152_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h2)
	) name974 (
		_w2145_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h8)
	) name975 (
		\g1088_reg/NET0131 ,
		\g228_reg/NET0131 ,
		_w2155_
	);
	LUT2 #(
		.INIT('h8)
	) name976 (
		\g1092_reg/NET0131 ,
		\g225_reg/NET0131 ,
		_w2156_
	);
	LUT2 #(
		.INIT('h8)
	) name977 (
		\g222_reg/NET0131 ,
		\g7961_pad ,
		_w2157_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		_w2155_,
		_w2156_,
		_w2158_
	);
	LUT2 #(
		.INIT('h4)
	) name979 (
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h2)
	) name980 (
		_w2047_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		_w2047_,
		_w2159_,
		_w2161_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		_w2160_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		\g186_reg/NET0131 ,
		\g7961_pad ,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name984 (
		\g1092_reg/NET0131 ,
		\g189_reg/NET0131 ,
		_w2164_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		\g1088_reg/NET0131 ,
		\g192_reg/NET0131 ,
		_w2165_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w2163_,
		_w2164_,
		_w2166_
	);
	LUT2 #(
		.INIT('h4)
	) name987 (
		_w2165_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		\g97_reg/NET0131 ,
		_w2167_,
		_w2168_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		\g97_reg/NET0131 ,
		_w2167_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		_w2168_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		\g1092_reg/NET0131 ,
		\g216_reg/NET0131 ,
		_w2171_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		\g1088_reg/NET0131 ,
		\g219_reg/NET0131 ,
		_w2172_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		\g213_reg/NET0131 ,
		\g7961_pad ,
		_w2173_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w2171_,
		_w2172_,
		_w2174_
	);
	LUT2 #(
		.INIT('h4)
	) name995 (
		_w2173_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		\g121_reg/NET0131 ,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		\g121_reg/NET0131 ,
		_w2175_,
		_w2177_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		_w2176_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h4)
	) name999 (
		_w2170_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		\g231_reg/NET0131 ,
		\g7961_pad ,
		_w2180_
	);
	LUT2 #(
		.INIT('h8)
	) name1001 (
		\g1088_reg/NET0131 ,
		\g237_reg/NET0131 ,
		_w2181_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		\g1092_reg/NET0131 ,
		\g234_reg/NET0131 ,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w2180_,
		_w2181_,
		_w2183_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h2)
	) name1005 (
		\g101_reg/NET0131 ,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h4)
	) name1006 (
		\g101_reg/NET0131 ,
		_w2184_,
		_w2186_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		_w2185_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		\g1088_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w2188_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		\g1092_reg/NET0131 ,
		\g198_reg/NET0131 ,
		_w2189_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		\g195_reg/NET0131 ,
		\g7961_pad ,
		_w2190_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w2188_,
		_w2189_,
		_w2191_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		_w2190_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h2)
	) name1013 (
		\g105_reg/NET0131 ,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h4)
	) name1014 (
		\g105_reg/NET0131 ,
		_w2192_,
		_w2194_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w2193_,
		_w2194_,
		_w2195_
	);
	LUT2 #(
		.INIT('h8)
	) name1016 (
		\g204_reg/NET0131 ,
		\g7961_pad ,
		_w2196_
	);
	LUT2 #(
		.INIT('h8)
	) name1017 (
		\g1092_reg/NET0131 ,
		\g207_reg/NET0131 ,
		_w2197_
	);
	LUT2 #(
		.INIT('h8)
	) name1018 (
		\g1088_reg/NET0131 ,
		\g210_reg/NET0131 ,
		_w2198_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		_w2196_,
		_w2197_,
		_w2199_
	);
	LUT2 #(
		.INIT('h4)
	) name1020 (
		_w2198_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		\g113_reg/NET0131 ,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		\g113_reg/NET0131 ,
		_w2200_,
		_w2202_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w2201_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h4)
	) name1024 (
		_w2195_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		\g249_reg/NET0131 ,
		\g7961_pad ,
		_w2205_
	);
	LUT2 #(
		.INIT('h8)
	) name1026 (
		\g1088_reg/NET0131 ,
		\g255_reg/NET0131 ,
		_w2206_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		\g1092_reg/NET0131 ,
		\g252_reg/NET0131 ,
		_w2207_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		_w2205_,
		_w2206_,
		_w2208_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		_w2207_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h2)
	) name1030 (
		\g117_reg/NET0131 ,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		\g117_reg/NET0131 ,
		_w2209_,
		_w2211_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w2210_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		\g1088_reg/NET0131 ,
		\g246_reg/NET0131 ,
		_w2213_
	);
	LUT2 #(
		.INIT('h8)
	) name1034 (
		\g1092_reg/NET0131 ,
		\g243_reg/NET0131 ,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		\g240_reg/NET0131 ,
		\g7961_pad ,
		_w2215_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w2213_,
		_w2214_,
		_w2216_
	);
	LUT2 #(
		.INIT('h4)
	) name1037 (
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h2)
	) name1038 (
		\g109_reg/NET0131 ,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h4)
	) name1039 (
		\g109_reg/NET0131 ,
		_w2217_,
		_w2219_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w2218_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w2212_,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h2)
	) name1042 (
		_w2162_,
		_w2187_,
		_w2222_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		_w2154_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name1044 (
		_w2179_,
		_w2204_,
		_w2224_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		_w2221_,
		_w2224_,
		_w2225_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		_w2223_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h1)
	) name1047 (
		_w2153_,
		_w2187_,
		_w2227_
	);
	LUT2 #(
		.INIT('h2)
	) name1048 (
		_w2212_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		_w2220_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		_w2153_,
		_w2212_,
		_w2230_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		_w2187_,
		_w2220_,
		_w2231_
	);
	LUT2 #(
		.INIT('h4)
	) name1052 (
		_w2228_,
		_w2231_,
		_w2232_
	);
	LUT2 #(
		.INIT('h1)
	) name1053 (
		_w2145_,
		_w2230_,
		_w2233_
	);
	LUT2 #(
		.INIT('h4)
	) name1054 (
		_w2232_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h4)
	) name1055 (
		_w2154_,
		_w2187_,
		_w2235_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		_w2221_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w2229_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		_w2234_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		_w2226_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name1060 (
		_w2024_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		_w2162_,
		_w2178_,
		_w2241_
	);
	LUT2 #(
		.INIT('h2)
	) name1062 (
		_w2170_,
		_w2204_,
		_w2242_
	);
	LUT2 #(
		.INIT('h4)
	) name1063 (
		_w2241_,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w2178_,
		_w2203_,
		_w2244_
	);
	LUT2 #(
		.INIT('h1)
	) name1065 (
		_w2170_,
		_w2195_,
		_w2245_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		_w2162_,
		_w2244_,
		_w2246_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h2)
	) name1068 (
		_w2162_,
		_w2195_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name1069 (
		_w2179_,
		_w2203_,
		_w2249_
	);
	LUT2 #(
		.INIT('h4)
	) name1070 (
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT2 #(
		.INIT('h1)
	) name1071 (
		_w2243_,
		_w2247_,
		_w2251_
	);
	LUT2 #(
		.INIT('h4)
	) name1072 (
		_w2250_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		_w2136_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h1)
	) name1074 (
		_w2116_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h4)
	) name1075 (
		_w2240_,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h2)
	) name1076 (
		\g1563_reg/NET0131 ,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		_w2137_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h2)
	) name1078 (
		_w2014_,
		_w2019_,
		_w2258_
	);
	LUT2 #(
		.INIT('h4)
	) name1079 (
		_w2257_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		\g403_reg/NET0131 ,
		\g7961_pad ,
		_w2260_
	);
	LUT2 #(
		.INIT('h2)
	) name1081 (
		\g1088_reg/NET0131 ,
		\g402_reg/NET0131 ,
		_w2261_
	);
	LUT2 #(
		.INIT('h2)
	) name1082 (
		\g1092_reg/NET0131 ,
		\g404_reg/NET0131 ,
		_w2262_
	);
	LUT2 #(
		.INIT('h1)
	) name1083 (
		_w2260_,
		_w2261_,
		_w2263_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		_w2262_,
		_w2263_,
		_w2264_
	);
	LUT2 #(
		.INIT('h2)
	) name1085 (
		_w2135_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h8)
	) name1086 (
		_w2019_,
		_w2024_,
		_w2266_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		_w2014_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		_w2024_,
		_w2239_,
		_w2268_
	);
	LUT2 #(
		.INIT('h2)
	) name1089 (
		_w2252_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h4)
	) name1090 (
		_w2019_,
		_w2117_,
		_w2270_
	);
	LUT2 #(
		.INIT('h4)
	) name1091 (
		_w2269_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w2267_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		_w2265_,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w2259_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		\g7961_pad ,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h1)
	) name1096 (
		\g315_reg/NET0131 ,
		\g7961_pad ,
		_w2276_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('h2)
	) name1098 (
		\g1092_reg/NET0131 ,
		_w2274_,
		_w2278_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		\g1092_reg/NET0131 ,
		\g316_reg/NET0131 ,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT2 #(
		.INIT('h2)
	) name1101 (
		\g1088_reg/NET0131 ,
		_w2274_,
		_w2281_
	);
	LUT2 #(
		.INIT('h1)
	) name1102 (
		\g1088_reg/NET0131 ,
		\g317_reg/NET0131 ,
		_w2282_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w2281_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h4)
	) name1104 (
		\g1006_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w2284_
	);
	LUT2 #(
		.INIT('h4)
	) name1105 (
		\g1005_reg/NET0131 ,
		\g7961_pad ,
		_w2285_
	);
	LUT2 #(
		.INIT('h4)
	) name1106 (
		\g1007_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name1107 (
		_w2284_,
		_w2285_,
		_w2287_
	);
	LUT2 #(
		.INIT('h4)
	) name1108 (
		_w2286_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h4)
	) name1109 (
		\g1010_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w2289_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		\g1008_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w2290_
	);
	LUT2 #(
		.INIT('h4)
	) name1111 (
		\g1009_reg/NET0131 ,
		\g7961_pad ,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w2289_,
		_w2290_,
		_w2292_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w2291_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h2)
	) name1114 (
		\g7961_pad ,
		\g860_reg/NET0131 ,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name1115 (
		\g1092_reg/NET0131 ,
		\g861_reg/NET0131 ,
		_w2295_
	);
	LUT2 #(
		.INIT('h2)
	) name1116 (
		\g1088_reg/NET0131 ,
		\g859_reg/NET0131 ,
		_w2296_
	);
	LUT2 #(
		.INIT('h1)
	) name1117 (
		_w2294_,
		_w2295_,
		_w2297_
	);
	LUT2 #(
		.INIT('h4)
	) name1118 (
		_w2296_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h2)
	) name1119 (
		\g1088_reg/NET0131 ,
		\g850_reg/NET0131 ,
		_w2299_
	);
	LUT2 #(
		.INIT('h2)
	) name1120 (
		\g1092_reg/NET0131 ,
		\g852_reg/NET0131 ,
		_w2300_
	);
	LUT2 #(
		.INIT('h2)
	) name1121 (
		\g7961_pad ,
		\g851_reg/NET0131 ,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1122 (
		_w2299_,
		_w2300_,
		_w2302_
	);
	LUT2 #(
		.INIT('h4)
	) name1123 (
		_w2301_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		_w2298_,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('h2)
	) name1125 (
		\g7961_pad ,
		\g842_reg/NET0131 ,
		_w2305_
	);
	LUT2 #(
		.INIT('h2)
	) name1126 (
		\g1092_reg/NET0131 ,
		\g843_reg/NET0131 ,
		_w2306_
	);
	LUT2 #(
		.INIT('h2)
	) name1127 (
		\g1088_reg/NET0131 ,
		\g841_reg/NET0131 ,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w2305_,
		_w2306_,
		_w2308_
	);
	LUT2 #(
		.INIT('h4)
	) name1129 (
		_w2307_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h2)
	) name1130 (
		\g809_reg/NET0131 ,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h4)
	) name1131 (
		\g809_reg/NET0131 ,
		_w2309_,
		_w2311_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w2310_,
		_w2311_,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name1133 (
		_w2298_,
		_w2303_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name1134 (
		\g7961_pad ,
		\g818_reg/NET0131 ,
		_w2314_
	);
	LUT2 #(
		.INIT('h2)
	) name1135 (
		\g1088_reg/NET0131 ,
		\g817_reg/NET0131 ,
		_w2315_
	);
	LUT2 #(
		.INIT('h2)
	) name1136 (
		\g1092_reg/NET0131 ,
		\g819_reg/NET0131 ,
		_w2316_
	);
	LUT2 #(
		.INIT('h1)
	) name1137 (
		_w2314_,
		_w2315_,
		_w2317_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		_w2316_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name1139 (
		\g785_reg/NET0131 ,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h4)
	) name1140 (
		\g785_reg/NET0131 ,
		_w2318_,
		_w2320_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w2319_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('h2)
	) name1142 (
		\g7961_pad ,
		\g821_reg/NET0131 ,
		_w2322_
	);
	LUT2 #(
		.INIT('h2)
	) name1143 (
		\g1092_reg/NET0131 ,
		\g822_reg/NET0131 ,
		_w2323_
	);
	LUT2 #(
		.INIT('h2)
	) name1144 (
		\g1088_reg/NET0131 ,
		\g820_reg/NET0131 ,
		_w2324_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w2322_,
		_w2323_,
		_w2325_
	);
	LUT2 #(
		.INIT('h4)
	) name1146 (
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		\g789_reg/NET0131 ,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		\g7961_pad ,
		\g830_reg/NET0131 ,
		_w2328_
	);
	LUT2 #(
		.INIT('h2)
	) name1149 (
		\g1092_reg/NET0131 ,
		\g831_reg/NET0131 ,
		_w2329_
	);
	LUT2 #(
		.INIT('h2)
	) name1150 (
		\g1088_reg/NET0131 ,
		\g829_reg/NET0131 ,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w2328_,
		_w2329_,
		_w2331_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		_w2330_,
		_w2331_,
		_w2332_
	);
	LUT2 #(
		.INIT('h2)
	) name1153 (
		\g793_reg/NET0131 ,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h4)
	) name1154 (
		\g793_reg/NET0131 ,
		_w2332_,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name1155 (
		_w2333_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		\g7961_pad ,
		\g833_reg/NET0131 ,
		_w2336_
	);
	LUT2 #(
		.INIT('h2)
	) name1157 (
		\g1088_reg/NET0131 ,
		\g832_reg/NET0131 ,
		_w2337_
	);
	LUT2 #(
		.INIT('h2)
	) name1158 (
		\g1092_reg/NET0131 ,
		\g834_reg/NET0131 ,
		_w2338_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		_w2336_,
		_w2337_,
		_w2339_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w2338_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\g797_reg/NET0131 ,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h4)
	) name1162 (
		\g797_reg/NET0131 ,
		_w2340_,
		_w2342_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		\g7961_pad ,
		\g836_reg/NET0131 ,
		_w2344_
	);
	LUT2 #(
		.INIT('h2)
	) name1165 (
		\g1092_reg/NET0131 ,
		\g837_reg/NET0131 ,
		_w2345_
	);
	LUT2 #(
		.INIT('h2)
	) name1166 (
		\g1088_reg/NET0131 ,
		\g835_reg/NET0131 ,
		_w2346_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w2344_,
		_w2345_,
		_w2347_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w2346_,
		_w2347_,
		_w2348_
	);
	LUT2 #(
		.INIT('h2)
	) name1169 (
		\g801_reg/NET0131 ,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h4)
	) name1170 (
		\g801_reg/NET0131 ,
		_w2348_,
		_w2350_
	);
	LUT2 #(
		.INIT('h1)
	) name1171 (
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h2)
	) name1172 (
		\g7961_pad ,
		\g863_reg/NET0131 ,
		_w2352_
	);
	LUT2 #(
		.INIT('h2)
	) name1173 (
		\g1092_reg/NET0131 ,
		\g864_reg/NET0131 ,
		_w2353_
	);
	LUT2 #(
		.INIT('h2)
	) name1174 (
		\g1088_reg/NET0131 ,
		\g862_reg/NET0131 ,
		_w2354_
	);
	LUT2 #(
		.INIT('h1)
	) name1175 (
		_w2352_,
		_w2353_,
		_w2355_
	);
	LUT2 #(
		.INIT('h4)
	) name1176 (
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h2)
	) name1177 (
		\g1092_reg/NET0131 ,
		\g849_reg/NET0131 ,
		_w2357_
	);
	LUT2 #(
		.INIT('h2)
	) name1178 (
		\g1088_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w2358_
	);
	LUT2 #(
		.INIT('h2)
	) name1179 (
		\g7961_pad ,
		\g848_reg/NET0131 ,
		_w2359_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w2357_,
		_w2358_,
		_w2360_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		_w2359_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w2356_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h8)
	) name1183 (
		_w2356_,
		_w2361_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w2362_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h2)
	) name1185 (
		\g1088_reg/NET0131 ,
		\g844_reg/NET0131 ,
		_w2365_
	);
	LUT2 #(
		.INIT('h2)
	) name1186 (
		\g1092_reg/NET0131 ,
		\g846_reg/NET0131 ,
		_w2366_
	);
	LUT2 #(
		.INIT('h2)
	) name1187 (
		\g7961_pad ,
		\g845_reg/NET0131 ,
		_w2367_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		_w2365_,
		_w2366_,
		_w2368_
	);
	LUT2 #(
		.INIT('h4)
	) name1189 (
		_w2367_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h2)
	) name1190 (
		\g813_reg/NET0131 ,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h4)
	) name1191 (
		\g813_reg/NET0131 ,
		_w2369_,
		_w2371_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		_w2370_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h2)
	) name1193 (
		\g1088_reg/NET0131 ,
		\g838_reg/NET0131 ,
		_w2373_
	);
	LUT2 #(
		.INIT('h2)
	) name1194 (
		\g1092_reg/NET0131 ,
		\g840_reg/NET0131 ,
		_w2374_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		\g7961_pad ,
		\g839_reg/NET0131 ,
		_w2375_
	);
	LUT2 #(
		.INIT('h1)
	) name1196 (
		_w2373_,
		_w2374_,
		_w2376_
	);
	LUT2 #(
		.INIT('h4)
	) name1197 (
		_w2375_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		\g805_reg/NET0131 ,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		\g1088_reg/NET0131 ,
		\g856_reg/NET0131 ,
		_w2379_
	);
	LUT2 #(
		.INIT('h2)
	) name1200 (
		\g1092_reg/NET0131 ,
		\g858_reg/NET0131 ,
		_w2380_
	);
	LUT2 #(
		.INIT('h2)
	) name1201 (
		\g7961_pad ,
		\g857_reg/NET0131 ,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w2379_,
		_w2380_,
		_w2382_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w2381_,
		_w2382_,
		_w2383_
	);
	LUT2 #(
		.INIT('h2)
	) name1204 (
		\g1563_reg/NET0131 ,
		_w2383_,
		_w2384_
	);
	LUT2 #(
		.INIT('h1)
	) name1205 (
		\g805_reg/NET0131 ,
		_w2377_,
		_w2385_
	);
	LUT2 #(
		.INIT('h8)
	) name1206 (
		\g789_reg/NET0131 ,
		_w2326_,
		_w2386_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w2304_,
		_w2313_,
		_w2387_
	);
	LUT2 #(
		.INIT('h1)
	) name1208 (
		_w2327_,
		_w2378_,
		_w2388_
	);
	LUT2 #(
		.INIT('h2)
	) name1209 (
		_w2384_,
		_w2385_,
		_w2389_
	);
	LUT2 #(
		.INIT('h4)
	) name1210 (
		_w2386_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h8)
	) name1211 (
		_w2387_,
		_w2388_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w2312_,
		_w2321_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name1213 (
		_w2335_,
		_w2343_,
		_w2393_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w2351_,
		_w2364_,
		_w2394_
	);
	LUT2 #(
		.INIT('h4)
	) name1215 (
		_w2372_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		_w2392_,
		_w2393_,
		_w2396_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		_w2390_,
		_w2391_,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name1218 (
		_w2396_,
		_w2397_,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		_w2395_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h4)
	) name1220 (
		_w2293_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		\g1563_reg/NET0131 ,
		_w2383_,
		_w2401_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		_w2400_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h4)
	) name1223 (
		_w2288_,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		\g1000_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w2404_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		\g7961_pad ,
		\g999_reg/NET0131 ,
		_w2405_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		\g1001_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name1227 (
		_w2404_,
		_w2405_,
		_w2407_
	);
	LUT2 #(
		.INIT('h4)
	) name1228 (
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h4)
	) name1229 (
		\g1004_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w2409_
	);
	LUT2 #(
		.INIT('h4)
	) name1230 (
		\g1002_reg/NET0131 ,
		\g7961_pad ,
		_w2410_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		\g1003_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w2411_
	);
	LUT2 #(
		.INIT('h1)
	) name1232 (
		_w2409_,
		_w2410_,
		_w2412_
	);
	LUT2 #(
		.INIT('h4)
	) name1233 (
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h4)
	) name1234 (
		_w2408_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		\g1088_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w2415_
	);
	LUT2 #(
		.INIT('h8)
	) name1236 (
		\g1092_reg/NET0131 ,
		\g930_reg/NET0131 ,
		_w2416_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		\g7961_pad ,
		\g927_reg/NET0131 ,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		_w2415_,
		_w2416_,
		_w2418_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		\g797_reg/NET0131 ,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		\g797_reg/NET0131 ,
		_w2419_,
		_w2421_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w2420_,
		_w2421_,
		_w2422_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		\g1088_reg/NET0131 ,
		\g960_reg/NET0131 ,
		_w2423_
	);
	LUT2 #(
		.INIT('h8)
	) name1244 (
		\g1092_reg/NET0131 ,
		\g957_reg/NET0131 ,
		_w2424_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		\g7961_pad ,
		\g954_reg/NET0131 ,
		_w2425_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w2423_,
		_w2424_,
		_w2426_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		_w2425_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name1248 (
		_w2298_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h4)
	) name1249 (
		_w2298_,
		_w2427_,
		_w2429_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		_w2422_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h8)
	) name1252 (
		\g7961_pad ,
		\g936_reg/NET0131 ,
		_w2432_
	);
	LUT2 #(
		.INIT('h8)
	) name1253 (
		\g1092_reg/NET0131 ,
		\g939_reg/NET0131 ,
		_w2433_
	);
	LUT2 #(
		.INIT('h8)
	) name1254 (
		\g1088_reg/NET0131 ,
		\g942_reg/NET0131 ,
		_w2434_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w2432_,
		_w2433_,
		_w2435_
	);
	LUT2 #(
		.INIT('h4)
	) name1256 (
		_w2434_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		\g805_reg/NET0131 ,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		\g805_reg/NET0131 ,
		_w2436_,
		_w2438_
	);
	LUT2 #(
		.INIT('h1)
	) name1259 (
		_w2437_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('h8)
	) name1260 (
		\g7961_pad ,
		\g945_reg/NET0131 ,
		_w2440_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		\g1088_reg/NET0131 ,
		\g951_reg/NET0131 ,
		_w2441_
	);
	LUT2 #(
		.INIT('h8)
	) name1262 (
		\g1092_reg/NET0131 ,
		\g948_reg/NET0131 ,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w2440_,
		_w2441_,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		_w2442_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name1265 (
		\g813_reg/NET0131 ,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h8)
	) name1266 (
		\g813_reg/NET0131 ,
		_w2444_,
		_w2446_
	);
	LUT2 #(
		.INIT('h1)
	) name1267 (
		_w2445_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h8)
	) name1268 (
		\g1088_reg/NET0131 ,
		\g924_reg/NET0131 ,
		_w2448_
	);
	LUT2 #(
		.INIT('h8)
	) name1269 (
		\g1092_reg/NET0131 ,
		\g921_reg/NET0131 ,
		_w2449_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		\g7961_pad ,
		\g918_reg/NET0131 ,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w2448_,
		_w2449_,
		_w2451_
	);
	LUT2 #(
		.INIT('h4)
	) name1272 (
		_w2450_,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h1)
	) name1273 (
		\g789_reg/NET0131 ,
		_w2452_,
		_w2453_
	);
	LUT2 #(
		.INIT('h8)
	) name1274 (
		\g789_reg/NET0131 ,
		_w2452_,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		_w2453_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h8)
	) name1276 (
		_w2422_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name1277 (
		_w2430_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h4)
	) name1278 (
		_w2447_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h2)
	) name1279 (
		_w2439_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h8)
	) name1280 (
		_w2447_,
		_w2455_,
		_w2460_
	);
	LUT2 #(
		.INIT('h4)
	) name1281 (
		_w2457_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h1)
	) name1282 (
		_w2431_,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w2459_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name1284 (
		_w2422_,
		_w2439_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name1285 (
		_w2430_,
		_w2447_,
		_w2465_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w2455_,
		_w2464_,
		_w2466_
	);
	LUT2 #(
		.INIT('h4)
	) name1287 (
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		_w2463_,
		_w2467_,
		_w2468_
	);
	LUT2 #(
		.INIT('h2)
	) name1289 (
		_w2384_,
		_w2468_,
		_w2469_
	);
	LUT2 #(
		.INIT('h8)
	) name1290 (
		\g1088_reg/NET0131 ,
		\g888_reg/NET0131 ,
		_w2470_
	);
	LUT2 #(
		.INIT('h8)
	) name1291 (
		\g1092_reg/NET0131 ,
		\g885_reg/NET0131 ,
		_w2471_
	);
	LUT2 #(
		.INIT('h8)
	) name1292 (
		\g7961_pad ,
		\g882_reg/NET0131 ,
		_w2472_
	);
	LUT2 #(
		.INIT('h1)
	) name1293 (
		_w2470_,
		_w2471_,
		_w2473_
	);
	LUT2 #(
		.INIT('h4)
	) name1294 (
		_w2472_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('h1)
	) name1295 (
		\g793_reg/NET0131 ,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		\g793_reg/NET0131 ,
		_w2474_,
		_w2476_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		_w2475_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h8)
	) name1298 (
		\g1088_reg/NET0131 ,
		\g915_reg/NET0131 ,
		_w2478_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		\g1092_reg/NET0131 ,
		\g912_reg/NET0131 ,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name1300 (
		\g7961_pad ,
		\g909_reg/NET0131 ,
		_w2480_
	);
	LUT2 #(
		.INIT('h1)
	) name1301 (
		_w2478_,
		_w2479_,
		_w2481_
	);
	LUT2 #(
		.INIT('h4)
	) name1302 (
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h2)
	) name1303 (
		_w2356_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h4)
	) name1304 (
		_w2356_,
		_w2482_,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w2483_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name1306 (
		_w2477_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		\g7961_pad ,
		\g891_reg/NET0131 ,
		_w2487_
	);
	LUT2 #(
		.INIT('h8)
	) name1308 (
		\g1092_reg/NET0131 ,
		\g894_reg/NET0131 ,
		_w2488_
	);
	LUT2 #(
		.INIT('h8)
	) name1309 (
		\g1088_reg/NET0131 ,
		\g897_reg/NET0131 ,
		_w2489_
	);
	LUT2 #(
		.INIT('h1)
	) name1310 (
		_w2487_,
		_w2488_,
		_w2490_
	);
	LUT2 #(
		.INIT('h4)
	) name1311 (
		_w2489_,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('h1)
	) name1312 (
		\g801_reg/NET0131 ,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h8)
	) name1313 (
		\g801_reg/NET0131 ,
		_w2491_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w2492_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		_w2486_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		\g1092_reg/NET0131 ,
		\g903_reg/NET0131 ,
		_w2496_
	);
	LUT2 #(
		.INIT('h8)
	) name1317 (
		\g1088_reg/NET0131 ,
		\g906_reg/NET0131 ,
		_w2497_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		\g7961_pad ,
		\g900_reg/NET0131 ,
		_w2498_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w2496_,
		_w2497_,
		_w2499_
	);
	LUT2 #(
		.INIT('h4)
	) name1320 (
		_w2498_,
		_w2499_,
		_w2500_
	);
	LUT2 #(
		.INIT('h1)
	) name1321 (
		\g809_reg/NET0131 ,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name1322 (
		\g809_reg/NET0131 ,
		_w2500_,
		_w2502_
	);
	LUT2 #(
		.INIT('h1)
	) name1323 (
		_w2501_,
		_w2502_,
		_w2503_
	);
	LUT2 #(
		.INIT('h2)
	) name1324 (
		_w2495_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h8)
	) name1325 (
		_w2477_,
		_w2494_,
		_w2505_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		\g7961_pad ,
		\g873_reg/NET0131 ,
		_w2506_
	);
	LUT2 #(
		.INIT('h8)
	) name1327 (
		\g1092_reg/NET0131 ,
		\g876_reg/NET0131 ,
		_w2507_
	);
	LUT2 #(
		.INIT('h8)
	) name1328 (
		\g1088_reg/NET0131 ,
		\g879_reg/NET0131 ,
		_w2508_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w2506_,
		_w2507_,
		_w2509_
	);
	LUT2 #(
		.INIT('h4)
	) name1330 (
		_w2508_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		\g785_reg/NET0131 ,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h4)
	) name1332 (
		\g785_reg/NET0131 ,
		_w2510_,
		_w2512_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		_w2511_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		_w2485_,
		_w2503_,
		_w2514_
	);
	LUT2 #(
		.INIT('h4)
	) name1335 (
		_w2495_,
		_w2514_,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1336 (
		_w2505_,
		_w2513_,
		_w2516_
	);
	LUT2 #(
		.INIT('h4)
	) name1337 (
		_w2515_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h2)
	) name1338 (
		_w2477_,
		_w2513_,
		_w2518_
	);
	LUT2 #(
		.INIT('h8)
	) name1339 (
		_w2494_,
		_w2503_,
		_w2519_
	);
	LUT2 #(
		.INIT('h1)
	) name1340 (
		_w2485_,
		_w2518_,
		_w2520_
	);
	LUT2 #(
		.INIT('h4)
	) name1341 (
		_w2519_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w2504_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('h4)
	) name1343 (
		_w2517_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h2)
	) name1344 (
		_w2384_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name1345 (
		_w2400_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		_w2455_,
		_w2485_,
		_w2526_
	);
	LUT2 #(
		.INIT('h8)
	) name1347 (
		_w2464_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		_w2465_,
		_w2518_,
		_w2528_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w2519_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		_w2527_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		_w2383_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h4)
	) name1352 (
		_w2525_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h2)
	) name1353 (
		\g1563_reg/NET0131 ,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h2)
	) name1354 (
		_w2288_,
		_w2469_,
		_w2534_
	);
	LUT2 #(
		.INIT('h4)
	) name1355 (
		_w2533_,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h4)
	) name1356 (
		_w2403_,
		_w2414_,
		_w2536_
	);
	LUT2 #(
		.INIT('h4)
	) name1357 (
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT2 #(
		.INIT('h4)
	) name1358 (
		\g1091_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w2538_
	);
	LUT2 #(
		.INIT('h2)
	) name1359 (
		\g1088_reg/NET0131 ,
		\g1089_reg/NET0131 ,
		_w2539_
	);
	LUT2 #(
		.INIT('h4)
	) name1360 (
		\g1090_reg/NET0131 ,
		\g7961_pad ,
		_w2540_
	);
	LUT2 #(
		.INIT('h1)
	) name1361 (
		_w2538_,
		_w2539_,
		_w2541_
	);
	LUT2 #(
		.INIT('h4)
	) name1362 (
		_w2540_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name1363 (
		_w2399_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		\g1563_reg/NET0131 ,
		_w2531_,
		_w2544_
	);
	LUT2 #(
		.INIT('h8)
	) name1365 (
		_w2288_,
		_w2468_,
		_w2545_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		_w2544_,
		_w2545_,
		_w2546_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w2524_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h1)
	) name1368 (
		_w2408_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		_w2413_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h8)
	) name1370 (
		_w2288_,
		_w2408_,
		_w2550_
	);
	LUT2 #(
		.INIT('h8)
	) name1371 (
		_w2413_,
		_w2550_,
		_w2551_
	);
	LUT2 #(
		.INIT('h1)
	) name1372 (
		_w2543_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h4)
	) name1373 (
		_w2537_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h4)
	) name1374 (
		_w2549_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h2)
	) name1375 (
		\g1092_reg/NET0131 ,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		\g1003_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name1378 (
		\g1092_reg/NET0131 ,
		_w1447_,
		_w2558_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		\g1092_reg/NET0131 ,
		\g2391_reg/NET0131 ,
		_w2559_
	);
	LUT2 #(
		.INIT('h1)
	) name1380 (
		_w2558_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name1381 (
		\g1088_reg/NET0131 ,
		_w1447_,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		\g1088_reg/NET0131 ,
		\g2392_reg/NET0131 ,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name1383 (
		_w2561_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h2)
	) name1384 (
		\g1088_reg/NET0131 ,
		_w2554_,
		_w2564_
	);
	LUT2 #(
		.INIT('h1)
	) name1385 (
		\g1004_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name1386 (
		_w2564_,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h2)
	) name1387 (
		\g7961_pad ,
		_w2554_,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name1388 (
		\g1002_reg/NET0131 ,
		\g7961_pad ,
		_w2568_
	);
	LUT2 #(
		.INIT('h1)
	) name1389 (
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h4)
	) name1390 (
		\g1693_reg/NET0131 ,
		\g7961_pad ,
		_w2570_
	);
	LUT2 #(
		.INIT('h2)
	) name1391 (
		\g1092_reg/NET0131 ,
		\g1694_reg/NET0131 ,
		_w2571_
	);
	LUT2 #(
		.INIT('h2)
	) name1392 (
		\g1088_reg/NET0131 ,
		\g1695_reg/NET0131 ,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		_w2570_,
		_w2571_,
		_w2573_
	);
	LUT2 #(
		.INIT('h4)
	) name1394 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h2)
	) name1395 (
		\g1092_reg/NET0131 ,
		\g1552_reg/NET0131 ,
		_w2575_
	);
	LUT2 #(
		.INIT('h4)
	) name1396 (
		\g1551_reg/NET0131 ,
		\g7961_pad ,
		_w2576_
	);
	LUT2 #(
		.INIT('h2)
	) name1397 (
		\g1088_reg/NET0131 ,
		\g1550_reg/NET0131 ,
		_w2577_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w2575_,
		_w2576_,
		_w2578_
	);
	LUT2 #(
		.INIT('h4)
	) name1399 (
		_w2577_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name1400 (
		\g1563_reg/NET0131 ,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name1401 (
		\g1585_reg/NET0131 ,
		\g7961_pad ,
		_w2581_
	);
	LUT2 #(
		.INIT('h8)
	) name1402 (
		\g1092_reg/NET0131 ,
		\g1588_reg/NET0131 ,
		_w2582_
	);
	LUT2 #(
		.INIT('h8)
	) name1403 (
		\g1088_reg/NET0131 ,
		\g1591_reg/NET0131 ,
		_w2583_
	);
	LUT2 #(
		.INIT('h1)
	) name1404 (
		_w2581_,
		_w2582_,
		_w2584_
	);
	LUT2 #(
		.INIT('h4)
	) name1405 (
		_w2583_,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		\g1491_reg/NET0131 ,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h8)
	) name1407 (
		\g1491_reg/NET0131 ,
		_w2585_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name1408 (
		_w2586_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h8)
	) name1409 (
		\g1088_reg/NET0131 ,
		\g1582_reg/NET0131 ,
		_w2589_
	);
	LUT2 #(
		.INIT('h8)
	) name1410 (
		\g1092_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		\g1576_reg/NET0131 ,
		\g7961_pad ,
		_w2591_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w2589_,
		_w2590_,
		_w2592_
	);
	LUT2 #(
		.INIT('h4)
	) name1413 (
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		\g1481_reg/NET0131 ,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h8)
	) name1415 (
		\g1481_reg/NET0131 ,
		_w2593_,
		_w2595_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		_w2594_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('h8)
	) name1417 (
		_w2588_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h8)
	) name1418 (
		\g1092_reg/NET0131 ,
		\g1597_reg/NET0131 ,
		_w2598_
	);
	LUT2 #(
		.INIT('h8)
	) name1419 (
		\g1088_reg/NET0131 ,
		\g1600_reg/NET0131 ,
		_w2599_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		\g1594_reg/NET0131 ,
		\g7961_pad ,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		_w2598_,
		_w2599_,
		_w2601_
	);
	LUT2 #(
		.INIT('h4)
	) name1422 (
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		\g1501_reg/NET0131 ,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h8)
	) name1424 (
		\g1501_reg/NET0131 ,
		_w2602_,
		_w2604_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		_w2603_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h2)
	) name1426 (
		\g1092_reg/NET0131 ,
		\g1558_reg/NET0131 ,
		_w2606_
	);
	LUT2 #(
		.INIT('h4)
	) name1427 (
		\g1557_reg/NET0131 ,
		\g7961_pad ,
		_w2607_
	);
	LUT2 #(
		.INIT('h2)
	) name1428 (
		\g1088_reg/NET0131 ,
		\g1556_reg/NET0131 ,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name1429 (
		_w2606_,
		_w2607_,
		_w2609_
	);
	LUT2 #(
		.INIT('h4)
	) name1430 (
		_w2608_,
		_w2609_,
		_w2610_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		\g1088_reg/NET0131 ,
		\g1609_reg/NET0131 ,
		_w2611_
	);
	LUT2 #(
		.INIT('h8)
	) name1432 (
		\g1092_reg/NET0131 ,
		\g1606_reg/NET0131 ,
		_w2612_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		\g1603_reg/NET0131 ,
		\g7961_pad ,
		_w2613_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w2611_,
		_w2612_,
		_w2614_
	);
	LUT2 #(
		.INIT('h4)
	) name1435 (
		_w2613_,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h2)
	) name1436 (
		_w2610_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h4)
	) name1437 (
		_w2610_,
		_w2615_,
		_w2617_
	);
	LUT2 #(
		.INIT('h1)
	) name1438 (
		_w2616_,
		_w2617_,
		_w2618_
	);
	LUT2 #(
		.INIT('h8)
	) name1439 (
		_w2605_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h8)
	) name1440 (
		\g1567_reg/NET0131 ,
		\g7961_pad ,
		_w2620_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		\g1088_reg/NET0131 ,
		\g1573_reg/NET0131 ,
		_w2621_
	);
	LUT2 #(
		.INIT('h8)
	) name1442 (
		\g1092_reg/NET0131 ,
		\g1570_reg/NET0131 ,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name1443 (
		_w2620_,
		_w2621_,
		_w2623_
	);
	LUT2 #(
		.INIT('h4)
	) name1444 (
		_w2622_,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('h2)
	) name1445 (
		\g1471_reg/NET0131 ,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h4)
	) name1446 (
		\g1471_reg/NET0131 ,
		_w2624_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name1447 (
		_w2625_,
		_w2626_,
		_w2627_
	);
	LUT2 #(
		.INIT('h4)
	) name1448 (
		_w2597_,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h4)
	) name1449 (
		_w2619_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h8)
	) name1450 (
		_w2588_,
		_w2605_,
		_w2630_
	);
	LUT2 #(
		.INIT('h2)
	) name1451 (
		_w2596_,
		_w2627_,
		_w2631_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		_w2618_,
		_w2630_,
		_w2632_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		_w2631_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h8)
	) name1454 (
		_w2596_,
		_w2618_,
		_w2634_
	);
	LUT2 #(
		.INIT('h2)
	) name1455 (
		_w2605_,
		_w2627_,
		_w2635_
	);
	LUT2 #(
		.INIT('h1)
	) name1456 (
		_w2588_,
		_w2634_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name1457 (
		_w2635_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		_w2629_,
		_w2633_,
		_w2638_
	);
	LUT2 #(
		.INIT('h4)
	) name1459 (
		_w2637_,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h2)
	) name1460 (
		_w2580_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		\g1092_reg/NET0131 ,
		\g1624_reg/NET0131 ,
		_w2641_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		\g1088_reg/NET0131 ,
		\g1627_reg/NET0131 ,
		_w2642_
	);
	LUT2 #(
		.INIT('h8)
	) name1463 (
		\g1621_reg/NET0131 ,
		\g7961_pad ,
		_w2643_
	);
	LUT2 #(
		.INIT('h1)
	) name1464 (
		_w2641_,
		_w2642_,
		_w2644_
	);
	LUT2 #(
		.INIT('h4)
	) name1465 (
		_w2643_,
		_w2644_,
		_w2645_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		\g1486_reg/NET0131 ,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h4)
	) name1467 (
		\g1486_reg/NET0131 ,
		_w2645_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		_w2646_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h8)
	) name1469 (
		\g1630_reg/NET0131 ,
		\g7961_pad ,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name1470 (
		\g1088_reg/NET0131 ,
		\g1636_reg/NET0131 ,
		_w2650_
	);
	LUT2 #(
		.INIT('h8)
	) name1471 (
		\g1092_reg/NET0131 ,
		\g1633_reg/NET0131 ,
		_w2651_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w2649_,
		_w2650_,
		_w2652_
	);
	LUT2 #(
		.INIT('h4)
	) name1473 (
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h2)
	) name1474 (
		\g1496_reg/NET0131 ,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		\g1496_reg/NET0131 ,
		_w2653_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name1476 (
		_w2654_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		_w2648_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h8)
	) name1478 (
		\g1092_reg/NET0131 ,
		\g1642_reg/NET0131 ,
		_w2658_
	);
	LUT2 #(
		.INIT('h8)
	) name1479 (
		\g1088_reg/NET0131 ,
		\g1645_reg/NET0131 ,
		_w2659_
	);
	LUT2 #(
		.INIT('h8)
	) name1480 (
		\g1639_reg/NET0131 ,
		\g7961_pad ,
		_w2660_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w2658_,
		_w2659_,
		_w2661_
	);
	LUT2 #(
		.INIT('h4)
	) name1482 (
		_w2660_,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h1)
	) name1483 (
		\g1506_reg/NET0131 ,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h8)
	) name1484 (
		\g1506_reg/NET0131 ,
		_w2662_,
		_w2664_
	);
	LUT2 #(
		.INIT('h1)
	) name1485 (
		_w2663_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h2)
	) name1486 (
		\g1092_reg/NET0131 ,
		\g1555_reg/NET0131 ,
		_w2666_
	);
	LUT2 #(
		.INIT('h4)
	) name1487 (
		\g1554_reg/NET0131 ,
		\g7961_pad ,
		_w2667_
	);
	LUT2 #(
		.INIT('h2)
	) name1488 (
		\g1088_reg/NET0131 ,
		\g1553_reg/NET0131 ,
		_w2668_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w2666_,
		_w2667_,
		_w2669_
	);
	LUT2 #(
		.INIT('h4)
	) name1490 (
		_w2668_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h8)
	) name1491 (
		\g1088_reg/NET0131 ,
		\g1654_reg/NET0131 ,
		_w2671_
	);
	LUT2 #(
		.INIT('h8)
	) name1492 (
		\g1092_reg/NET0131 ,
		\g1651_reg/NET0131 ,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name1493 (
		\g1648_reg/NET0131 ,
		\g7961_pad ,
		_w2673_
	);
	LUT2 #(
		.INIT('h1)
	) name1494 (
		_w2671_,
		_w2672_,
		_w2674_
	);
	LUT2 #(
		.INIT('h4)
	) name1495 (
		_w2673_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name1496 (
		_w2670_,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h4)
	) name1497 (
		_w2670_,
		_w2675_,
		_w2677_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		_w2676_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h8)
	) name1499 (
		_w2665_,
		_w2678_,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name1500 (
		\g1088_reg/NET0131 ,
		\g1618_reg/NET0131 ,
		_w2680_
	);
	LUT2 #(
		.INIT('h8)
	) name1501 (
		\g1092_reg/NET0131 ,
		\g1615_reg/NET0131 ,
		_w2681_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		\g1612_reg/NET0131 ,
		\g7961_pad ,
		_w2682_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w2680_,
		_w2681_,
		_w2683_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w2682_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		\g1476_reg/NET0131 ,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		\g1476_reg/NET0131 ,
		_w2684_,
		_w2686_
	);
	LUT2 #(
		.INIT('h1)
	) name1507 (
		_w2685_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h4)
	) name1508 (
		_w2627_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		_w2630_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		_w2634_,
		_w2657_,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name1511 (
		_w2679_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h8)
	) name1512 (
		_w2689_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name1513 (
		_w2579_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		\g1563_reg/NET0131 ,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h4)
	) name1515 (
		\g1699_reg/NET0131 ,
		\g7961_pad ,
		_w2695_
	);
	LUT2 #(
		.INIT('h2)
	) name1516 (
		\g1088_reg/NET0131 ,
		\g1701_reg/NET0131 ,
		_w2696_
	);
	LUT2 #(
		.INIT('h2)
	) name1517 (
		\g1092_reg/NET0131 ,
		\g1700_reg/NET0131 ,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name1518 (
		_w2695_,
		_w2696_,
		_w2698_
	);
	LUT2 #(
		.INIT('h4)
	) name1519 (
		_w2697_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name1520 (
		_w2665_,
		_w2687_,
		_w2700_
	);
	LUT2 #(
		.INIT('h2)
	) name1521 (
		_w2656_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1522 (
		_w2648_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		_w2656_,
		_w2665_,
		_w2703_
	);
	LUT2 #(
		.INIT('h4)
	) name1524 (
		_w2648_,
		_w2687_,
		_w2704_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		_w2701_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name1526 (
		_w2678_,
		_w2703_,
		_w2706_
	);
	LUT2 #(
		.INIT('h4)
	) name1527 (
		_w2705_,
		_w2706_,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name1528 (
		_w2657_,
		_w2687_,
		_w2708_
	);
	LUT2 #(
		.INIT('h4)
	) name1529 (
		_w2679_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w2702_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h4)
	) name1531 (
		_w2707_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name1532 (
		_w2699_,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		_w2694_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h1)
	) name1534 (
		_w2640_,
		_w2713_,
		_w2714_
	);
	LUT2 #(
		.INIT('h1)
	) name1535 (
		_w2574_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h2)
	) name1536 (
		\g1088_reg/NET0131 ,
		\g1698_reg/NET0131 ,
		_w2716_
	);
	LUT2 #(
		.INIT('h2)
	) name1537 (
		\g1092_reg/NET0131 ,
		\g1697_reg/NET0131 ,
		_w2717_
	);
	LUT2 #(
		.INIT('h4)
	) name1538 (
		\g1696_reg/NET0131 ,
		\g7961_pad ,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w2716_,
		_w2717_,
		_w2719_
	);
	LUT2 #(
		.INIT('h4)
	) name1540 (
		_w2718_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name1541 (
		_w2715_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h4)
	) name1542 (
		\g1703_reg/NET0131 ,
		\g7961_pad ,
		_w2722_
	);
	LUT2 #(
		.INIT('h2)
	) name1543 (
		\g1092_reg/NET0131 ,
		\g1704_reg/NET0131 ,
		_w2723_
	);
	LUT2 #(
		.INIT('h2)
	) name1544 (
		\g1088_reg/NET0131 ,
		\g1702_reg/NET0131 ,
		_w2724_
	);
	LUT2 #(
		.INIT('h1)
	) name1545 (
		_w2722_,
		_w2723_,
		_w2725_
	);
	LUT2 #(
		.INIT('h4)
	) name1546 (
		_w2724_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h2)
	) name1547 (
		\g1092_reg/NET0131 ,
		\g1525_reg/NET0131 ,
		_w2727_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		\g1524_reg/NET0131 ,
		\g7961_pad ,
		_w2728_
	);
	LUT2 #(
		.INIT('h2)
	) name1549 (
		\g1088_reg/NET0131 ,
		\g1523_reg/NET0131 ,
		_w2729_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		_w2727_,
		_w2728_,
		_w2730_
	);
	LUT2 #(
		.INIT('h4)
	) name1551 (
		_w2729_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name1552 (
		\g1481_reg/NET0131 ,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h4)
	) name1553 (
		\g1481_reg/NET0131 ,
		_w2731_,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w2732_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h4)
	) name1555 (
		\g1527_reg/NET0131 ,
		\g7961_pad ,
		_w2735_
	);
	LUT2 #(
		.INIT('h2)
	) name1556 (
		\g1088_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w2736_
	);
	LUT2 #(
		.INIT('h2)
	) name1557 (
		\g1092_reg/NET0131 ,
		\g1528_reg/NET0131 ,
		_w2737_
	);
	LUT2 #(
		.INIT('h1)
	) name1558 (
		_w2735_,
		_w2736_,
		_w2738_
	);
	LUT2 #(
		.INIT('h4)
	) name1559 (
		_w2737_,
		_w2738_,
		_w2739_
	);
	LUT2 #(
		.INIT('h2)
	) name1560 (
		\g1486_reg/NET0131 ,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h4)
	) name1561 (
		\g1486_reg/NET0131 ,
		_w2739_,
		_w2741_
	);
	LUT2 #(
		.INIT('h1)
	) name1562 (
		_w2740_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h4)
	) name1563 (
		\g1512_reg/NET0131 ,
		\g7961_pad ,
		_w2743_
	);
	LUT2 #(
		.INIT('h2)
	) name1564 (
		\g1088_reg/NET0131 ,
		\g1511_reg/NET0131 ,
		_w2744_
	);
	LUT2 #(
		.INIT('h2)
	) name1565 (
		\g1092_reg/NET0131 ,
		\g1513_reg/NET0131 ,
		_w2745_
	);
	LUT2 #(
		.INIT('h1)
	) name1566 (
		_w2743_,
		_w2744_,
		_w2746_
	);
	LUT2 #(
		.INIT('h4)
	) name1567 (
		_w2745_,
		_w2746_,
		_w2747_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		\g1471_reg/NET0131 ,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h4)
	) name1569 (
		\g1471_reg/NET0131 ,
		_w2747_,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w2748_,
		_w2749_,
		_w2750_
	);
	LUT2 #(
		.INIT('h4)
	) name1571 (
		\g1539_reg/NET0131 ,
		\g7961_pad ,
		_w2751_
	);
	LUT2 #(
		.INIT('h2)
	) name1572 (
		\g1088_reg/NET0131 ,
		\g1538_reg/NET0131 ,
		_w2752_
	);
	LUT2 #(
		.INIT('h2)
	) name1573 (
		\g1092_reg/NET0131 ,
		\g1540_reg/NET0131 ,
		_w2753_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		_w2751_,
		_w2752_,
		_w2754_
	);
	LUT2 #(
		.INIT('h4)
	) name1575 (
		_w2753_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h2)
	) name1576 (
		\g1506_reg/NET0131 ,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h4)
	) name1577 (
		\g1506_reg/NET0131 ,
		_w2755_,
		_w2757_
	);
	LUT2 #(
		.INIT('h1)
	) name1578 (
		_w2756_,
		_w2757_,
		_w2758_
	);
	LUT2 #(
		.INIT('h2)
	) name1579 (
		\g1092_reg/NET0131 ,
		\g1537_reg/NET0131 ,
		_w2759_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		\g1088_reg/NET0131 ,
		\g1535_reg/NET0131 ,
		_w2760_
	);
	LUT2 #(
		.INIT('h4)
	) name1581 (
		\g1536_reg/NET0131 ,
		\g7961_pad ,
		_w2761_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		_w2759_,
		_w2760_,
		_w2762_
	);
	LUT2 #(
		.INIT('h4)
	) name1583 (
		_w2761_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h2)
	) name1584 (
		\g1501_reg/NET0131 ,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name1585 (
		\g1501_reg/NET0131 ,
		_w2763_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		_w2764_,
		_w2765_,
		_w2766_
	);
	LUT2 #(
		.INIT('h2)
	) name1587 (
		\g1088_reg/NET0131 ,
		\g1529_reg/NET0131 ,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name1588 (
		\g1092_reg/NET0131 ,
		\g1531_reg/NET0131 ,
		_w2768_
	);
	LUT2 #(
		.INIT('h4)
	) name1589 (
		\g1530_reg/NET0131 ,
		\g7961_pad ,
		_w2769_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w2767_,
		_w2768_,
		_w2770_
	);
	LUT2 #(
		.INIT('h4)
	) name1591 (
		_w2769_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name1592 (
		\g1491_reg/NET0131 ,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h4)
	) name1593 (
		\g1491_reg/NET0131 ,
		_w2771_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name1594 (
		_w2772_,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h4)
	) name1595 (
		\g1515_reg/NET0131 ,
		\g7961_pad ,
		_w2775_
	);
	LUT2 #(
		.INIT('h2)
	) name1596 (
		\g1088_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		_w2776_
	);
	LUT2 #(
		.INIT('h2)
	) name1597 (
		\g1092_reg/NET0131 ,
		\g1516_reg/NET0131 ,
		_w2777_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w2775_,
		_w2776_,
		_w2778_
	);
	LUT2 #(
		.INIT('h4)
	) name1599 (
		_w2777_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h4)
	) name1600 (
		\g1476_reg/NET0131 ,
		_w2779_,
		_w2780_
	);
	LUT2 #(
		.INIT('h2)
	) name1601 (
		\g1476_reg/NET0131 ,
		_w2779_,
		_w2781_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w2780_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h2)
	) name1603 (
		\g1092_reg/NET0131 ,
		\g1546_reg/NET0131 ,
		_w2783_
	);
	LUT2 #(
		.INIT('h2)
	) name1604 (
		\g1088_reg/NET0131 ,
		\g1544_reg/NET0131 ,
		_w2784_
	);
	LUT2 #(
		.INIT('h4)
	) name1605 (
		\g1545_reg/NET0131 ,
		\g7961_pad ,
		_w2785_
	);
	LUT2 #(
		.INIT('h1)
	) name1606 (
		_w2783_,
		_w2784_,
		_w2786_
	);
	LUT2 #(
		.INIT('h4)
	) name1607 (
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w2670_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		_w2670_,
		_w2787_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w2788_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h2)
	) name1611 (
		\g1092_reg/NET0131 ,
		\g1543_reg/NET0131 ,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name1612 (
		\g1088_reg/NET0131 ,
		\g1541_reg/NET0131 ,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name1613 (
		\g1542_reg/NET0131 ,
		\g7961_pad ,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name1614 (
		_w2791_,
		_w2792_,
		_w2794_
	);
	LUT2 #(
		.INIT('h4)
	) name1615 (
		_w2793_,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h1)
	) name1616 (
		_w2610_,
		_w2795_,
		_w2796_
	);
	LUT2 #(
		.INIT('h8)
	) name1617 (
		_w2610_,
		_w2795_,
		_w2797_
	);
	LUT2 #(
		.INIT('h1)
	) name1618 (
		_w2796_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name1619 (
		\g1092_reg/NET0131 ,
		\g1534_reg/NET0131 ,
		_w2799_
	);
	LUT2 #(
		.INIT('h2)
	) name1620 (
		\g1088_reg/NET0131 ,
		\g1532_reg/NET0131 ,
		_w2800_
	);
	LUT2 #(
		.INIT('h4)
	) name1621 (
		\g1533_reg/NET0131 ,
		\g7961_pad ,
		_w2801_
	);
	LUT2 #(
		.INIT('h1)
	) name1622 (
		_w2799_,
		_w2800_,
		_w2802_
	);
	LUT2 #(
		.INIT('h4)
	) name1623 (
		_w2801_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h2)
	) name1624 (
		\g1496_reg/NET0131 ,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h4)
	) name1625 (
		\g1496_reg/NET0131 ,
		_w2803_,
		_w2805_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		_w2804_,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		_w2580_,
		_w2734_,
		_w2807_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w2742_,
		_w2750_,
		_w2808_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		_w2758_,
		_w2766_,
		_w2809_
	);
	LUT2 #(
		.INIT('h1)
	) name1630 (
		_w2774_,
		_w2782_,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w2790_,
		_w2798_,
		_w2811_
	);
	LUT2 #(
		.INIT('h4)
	) name1632 (
		_w2806_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h8)
	) name1633 (
		_w2809_,
		_w2810_,
		_w2813_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		_w2807_,
		_w2808_,
		_w2814_
	);
	LUT2 #(
		.INIT('h8)
	) name1635 (
		_w2813_,
		_w2814_,
		_w2815_
	);
	LUT2 #(
		.INIT('h8)
	) name1636 (
		_w2812_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h4)
	) name1637 (
		_w2726_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h8)
	) name1638 (
		\g1563_reg/NET0131 ,
		_w2579_,
		_w2818_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w2817_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h4)
	) name1640 (
		_w2699_,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h4)
	) name1641 (
		_w2640_,
		_w2817_,
		_w2821_
	);
	LUT2 #(
		.INIT('h2)
	) name1642 (
		_w2693_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		\g1563_reg/NET0131 ,
		_w2822_,
		_w2823_
	);
	LUT2 #(
		.INIT('h2)
	) name1644 (
		_w2580_,
		_w2711_,
		_w2824_
	);
	LUT2 #(
		.INIT('h2)
	) name1645 (
		_w2699_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h4)
	) name1646 (
		_w2823_,
		_w2825_,
		_w2826_
	);
	LUT2 #(
		.INIT('h4)
	) name1647 (
		_w2574_,
		_w2720_,
		_w2827_
	);
	LUT2 #(
		.INIT('h4)
	) name1648 (
		_w2820_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h4)
	) name1649 (
		_w2826_,
		_w2828_,
		_w2829_
	);
	LUT2 #(
		.INIT('h4)
	) name1650 (
		\g1784_reg/NET0131 ,
		\g7961_pad ,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name1651 (
		\g1092_reg/NET0131 ,
		\g1785_reg/NET0131 ,
		_w2831_
	);
	LUT2 #(
		.INIT('h2)
	) name1652 (
		\g1088_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w2832_
	);
	LUT2 #(
		.INIT('h1)
	) name1653 (
		_w2830_,
		_w2831_,
		_w2833_
	);
	LUT2 #(
		.INIT('h4)
	) name1654 (
		_w2832_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h2)
	) name1655 (
		_w2816_,
		_w2834_,
		_w2835_
	);
	LUT2 #(
		.INIT('h8)
	) name1656 (
		_w2574_,
		_w2699_,
		_w2836_
	);
	LUT2 #(
		.INIT('h8)
	) name1657 (
		_w2720_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		_w2835_,
		_w2837_,
		_w2838_
	);
	LUT2 #(
		.INIT('h4)
	) name1659 (
		_w2721_,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('h4)
	) name1660 (
		_w2829_,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h2)
	) name1661 (
		\g7961_pad ,
		_w2840_,
		_w2841_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		\g1696_reg/NET0131 ,
		\g7961_pad ,
		_w2842_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h2)
	) name1664 (
		\g1092_reg/NET0131 ,
		_w2840_,
		_w2844_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		\g1092_reg/NET0131 ,
		\g1697_reg/NET0131 ,
		_w2845_
	);
	LUT2 #(
		.INIT('h1)
	) name1666 (
		_w2844_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name1667 (
		\g1088_reg/NET0131 ,
		_w2840_,
		_w2847_
	);
	LUT2 #(
		.INIT('h1)
	) name1668 (
		\g1088_reg/NET0131 ,
		\g1698_reg/NET0131 ,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name1669 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w2850_
	);
	LUT2 #(
		.INIT('h4)
	) name1671 (
		_w1537_,
		_w2850_,
		_w2851_
	);
	LUT2 #(
		.INIT('h8)
	) name1672 (
		\g1186_reg/NET0131 ,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h2)
	) name1673 (
		\g1018_reg/NET0131 ,
		\g1410_reg/NET0131 ,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		\g1024_reg/NET0131 ,
		\g1408_reg/NET0131 ,
		_w2854_
	);
	LUT2 #(
		.INIT('h4)
	) name1675 (
		\g1409_reg/NET0131 ,
		\g5657_pad ,
		_w2855_
	);
	LUT2 #(
		.INIT('h1)
	) name1676 (
		_w2853_,
		_w2854_,
		_w2856_
	);
	LUT2 #(
		.INIT('h4)
	) name1677 (
		_w2855_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h2)
	) name1678 (
		\g1024_reg/NET0131 ,
		\g1396_reg/NET0131 ,
		_w2858_
	);
	LUT2 #(
		.INIT('h2)
	) name1679 (
		\g1018_reg/NET0131 ,
		\g1398_reg/NET0131 ,
		_w2859_
	);
	LUT2 #(
		.INIT('h4)
	) name1680 (
		\g1397_reg/NET0131 ,
		\g5657_pad ,
		_w2860_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w2858_,
		_w2859_,
		_w2861_
	);
	LUT2 #(
		.INIT('h4)
	) name1682 (
		_w2860_,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h2)
	) name1683 (
		\g1024_reg/NET0131 ,
		\g1384_reg/NET0131 ,
		_w2863_
	);
	LUT2 #(
		.INIT('h2)
	) name1684 (
		\g1018_reg/NET0131 ,
		\g1386_reg/NET0131 ,
		_w2864_
	);
	LUT2 #(
		.INIT('h4)
	) name1685 (
		\g1385_reg/NET0131 ,
		\g5657_pad ,
		_w2865_
	);
	LUT2 #(
		.INIT('h1)
	) name1686 (
		_w2863_,
		_w2864_,
		_w2866_
	);
	LUT2 #(
		.INIT('h4)
	) name1687 (
		_w2865_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h2)
	) name1688 (
		\g1018_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w2868_
	);
	LUT2 #(
		.INIT('h2)
	) name1689 (
		\g1024_reg/NET0131 ,
		\g1387_reg/NET0131 ,
		_w2869_
	);
	LUT2 #(
		.INIT('h4)
	) name1690 (
		\g1388_reg/NET0131 ,
		\g5657_pad ,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w2868_,
		_w2869_,
		_w2871_
	);
	LUT2 #(
		.INIT('h4)
	) name1692 (
		_w2870_,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h2)
	) name1693 (
		\g1018_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		_w2873_
	);
	LUT2 #(
		.INIT('h2)
	) name1694 (
		\g1024_reg/NET0131 ,
		\g1402_reg/NET0131 ,
		_w2874_
	);
	LUT2 #(
		.INIT('h4)
	) name1695 (
		\g1403_reg/NET0131 ,
		\g5657_pad ,
		_w2875_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w2873_,
		_w2874_,
		_w2876_
	);
	LUT2 #(
		.INIT('h4)
	) name1697 (
		_w2875_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h2)
	) name1698 (
		\g1018_reg/NET0131 ,
		\g1395_reg/NET0131 ,
		_w2878_
	);
	LUT2 #(
		.INIT('h2)
	) name1699 (
		\g1024_reg/NET0131 ,
		\g1393_reg/NET0131 ,
		_w2879_
	);
	LUT2 #(
		.INIT('h4)
	) name1700 (
		\g1394_reg/NET0131 ,
		\g5657_pad ,
		_w2880_
	);
	LUT2 #(
		.INIT('h1)
	) name1701 (
		_w2878_,
		_w2879_,
		_w2881_
	);
	LUT2 #(
		.INIT('h4)
	) name1702 (
		_w2880_,
		_w2881_,
		_w2882_
	);
	LUT2 #(
		.INIT('h2)
	) name1703 (
		\g1024_reg/NET0131 ,
		\g1411_reg/NET0131 ,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name1704 (
		\g1018_reg/NET0131 ,
		\g1413_reg/NET0131 ,
		_w2884_
	);
	LUT2 #(
		.INIT('h4)
	) name1705 (
		\g1412_reg/NET0131 ,
		\g5657_pad ,
		_w2885_
	);
	LUT2 #(
		.INIT('h1)
	) name1706 (
		_w2883_,
		_w2884_,
		_w2886_
	);
	LUT2 #(
		.INIT('h4)
	) name1707 (
		_w2885_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h2)
	) name1708 (
		\g1018_reg/NET0131 ,
		\g1407_reg/NET0131 ,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name1709 (
		\g1024_reg/NET0131 ,
		\g1405_reg/NET0131 ,
		_w2889_
	);
	LUT2 #(
		.INIT('h4)
	) name1710 (
		\g1406_reg/NET0131 ,
		\g5657_pad ,
		_w2890_
	);
	LUT2 #(
		.INIT('h1)
	) name1711 (
		_w2888_,
		_w2889_,
		_w2891_
	);
	LUT2 #(
		.INIT('h4)
	) name1712 (
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h4)
	) name1713 (
		\g1424_reg/NET0131 ,
		\g5657_pad ,
		_w2893_
	);
	LUT2 #(
		.INIT('h2)
	) name1714 (
		\g1024_reg/NET0131 ,
		\g1423_reg/NET0131 ,
		_w2894_
	);
	LUT2 #(
		.INIT('h2)
	) name1715 (
		\g1018_reg/NET0131 ,
		\g1425_reg/NET0131 ,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w2893_,
		_w2894_,
		_w2896_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w2895_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h4)
	) name1718 (
		\g1418_reg/NET0131 ,
		\g5657_pad ,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		\g1018_reg/NET0131 ,
		\g1419_reg/NET0131 ,
		_w2899_
	);
	LUT2 #(
		.INIT('h2)
	) name1720 (
		\g1024_reg/NET0131 ,
		\g1417_reg/NET0131 ,
		_w2900_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		_w2898_,
		_w2899_,
		_w2901_
	);
	LUT2 #(
		.INIT('h4)
	) name1722 (
		_w2900_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h2)
	) name1723 (
		\g1018_reg/NET0131 ,
		\g1401_reg/NET0131 ,
		_w2903_
	);
	LUT2 #(
		.INIT('h2)
	) name1724 (
		\g1024_reg/NET0131 ,
		\g1399_reg/NET0131 ,
		_w2904_
	);
	LUT2 #(
		.INIT('h4)
	) name1725 (
		\g1400_reg/NET0131 ,
		\g5657_pad ,
		_w2905_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w2903_,
		_w2904_,
		_w2906_
	);
	LUT2 #(
		.INIT('h4)
	) name1727 (
		_w2905_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		\g1018_reg/NET0131 ,
		\g1392_reg/NET0131 ,
		_w2908_
	);
	LUT2 #(
		.INIT('h2)
	) name1729 (
		\g1024_reg/NET0131 ,
		\g1390_reg/NET0131 ,
		_w2909_
	);
	LUT2 #(
		.INIT('h4)
	) name1730 (
		\g1391_reg/NET0131 ,
		\g5657_pad ,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name1731 (
		_w2908_,
		_w2909_,
		_w2911_
	);
	LUT2 #(
		.INIT('h4)
	) name1732 (
		_w2910_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h4)
	) name1733 (
		_w2857_,
		_w2862_,
		_w2913_
	);
	LUT2 #(
		.INIT('h2)
	) name1734 (
		_w2867_,
		_w2872_,
		_w2914_
	);
	LUT2 #(
		.INIT('h2)
	) name1735 (
		_w2877_,
		_w2882_,
		_w2915_
	);
	LUT2 #(
		.INIT('h4)
	) name1736 (
		_w2887_,
		_w2892_,
		_w2916_
	);
	LUT2 #(
		.INIT('h1)
	) name1737 (
		_w2897_,
		_w2902_,
		_w2917_
	);
	LUT2 #(
		.INIT('h2)
	) name1738 (
		_w2907_,
		_w2912_,
		_w2918_
	);
	LUT2 #(
		.INIT('h8)
	) name1739 (
		_w2917_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h8)
	) name1740 (
		_w2915_,
		_w2916_,
		_w2920_
	);
	LUT2 #(
		.INIT('h8)
	) name1741 (
		_w2913_,
		_w2914_,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name1742 (
		_w2920_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h8)
	) name1743 (
		_w2919_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w2857_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h8)
	) name1745 (
		\g1018_reg/NET0131 ,
		\g1303_reg/NET0131 ,
		_w2925_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		\g1024_reg/NET0131 ,
		\g1306_reg/NET0131 ,
		_w2926_
	);
	LUT2 #(
		.INIT('h8)
	) name1747 (
		\g1300_reg/NET0131 ,
		\g5657_pad ,
		_w2927_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		_w2925_,
		_w2926_,
		_w2928_
	);
	LUT2 #(
		.INIT('h4)
	) name1749 (
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h2)
	) name1750 (
		_w2924_,
		_w2929_,
		_w2930_
	);
	LUT2 #(
		.INIT('h4)
	) name1751 (
		_w2924_,
		_w2929_,
		_w2931_
	);
	LUT2 #(
		.INIT('h1)
	) name1752 (
		_w2930_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h2)
	) name1753 (
		_w2852_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		\g1291_reg/NET0131 ,
		\g5657_pad ,
		_w2934_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		\g1024_reg/NET0131 ,
		\g1297_reg/NET0131 ,
		_w2935_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		\g1018_reg/NET0131 ,
		\g1294_reg/NET0131 ,
		_w2936_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w2934_,
		_w2935_,
		_w2937_
	);
	LUT2 #(
		.INIT('h4)
	) name1758 (
		_w2936_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w2887_,
		_w2923_,
		_w2939_
	);
	LUT2 #(
		.INIT('h4)
	) name1760 (
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h2)
	) name1761 (
		_w2938_,
		_w2939_,
		_w2941_
	);
	LUT2 #(
		.INIT('h1)
	) name1762 (
		_w2940_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		_w2933_,
		_w2942_,
		_w2943_
	);
	LUT2 #(
		.INIT('h2)
	) name1764 (
		_w2852_,
		_w2942_,
		_w2944_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w2932_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h1)
	) name1766 (
		_w2943_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h2)
	) name1767 (
		\g1243_reg/NET0131 ,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h4)
	) name1768 (
		\g1224_reg/NET0131 ,
		\g3229_pad ,
		_w2948_
	);
	LUT2 #(
		.INIT('h8)
	) name1769 (
		\g1211_reg/NET0131 ,
		_w1550_,
		_w2949_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		\g1227_reg/NET0131 ,
		\g3229_pad ,
		_w2950_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w2948_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h8)
	) name1772 (
		_w2949_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		_w2851_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h2)
	) name1774 (
		_w2867_,
		_w2929_,
		_w2954_
	);
	LUT2 #(
		.INIT('h4)
	) name1775 (
		_w2867_,
		_w2929_,
		_w2955_
	);
	LUT2 #(
		.INIT('h1)
	) name1776 (
		_w2954_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		_w2852_,
		_w2956_,
		_w2957_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w2912_,
		_w2923_,
		_w2958_
	);
	LUT2 #(
		.INIT('h4)
	) name1779 (
		_w2929_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name1780 (
		_w2929_,
		_w2958_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w2959_,
		_w2960_,
		_w2961_
	);
	LUT2 #(
		.INIT('h2)
	) name1782 (
		_w2852_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w2882_,
		_w2923_,
		_w2963_
	);
	LUT2 #(
		.INIT('h4)
	) name1784 (
		_w2938_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h2)
	) name1785 (
		_w2938_,
		_w2963_,
		_w2965_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		_w2964_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h8)
	) name1787 (
		_w2962_,
		_w2966_,
		_w2967_
	);
	LUT2 #(
		.INIT('h2)
	) name1788 (
		_w2852_,
		_w2966_,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		_w2961_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h1)
	) name1790 (
		_w2967_,
		_w2969_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w2872_,
		_w2923_,
		_w2971_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w2938_,
		_w2971_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name1793 (
		_w2938_,
		_w2971_,
		_w2973_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		_w2852_,
		_w2972_,
		_w2974_
	);
	LUT2 #(
		.INIT('h4)
	) name1795 (
		_w2973_,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h2)
	) name1796 (
		_w2970_,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h4)
	) name1797 (
		_w2970_,
		_w2975_,
		_w2977_
	);
	LUT2 #(
		.INIT('h1)
	) name1798 (
		_w2976_,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h8)
	) name1799 (
		_w2957_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name1800 (
		_w2957_,
		_w2978_,
		_w2980_
	);
	LUT2 #(
		.INIT('h1)
	) name1801 (
		_w2979_,
		_w2980_,
		_w2981_
	);
	LUT2 #(
		.INIT('h4)
	) name1802 (
		_w2907_,
		_w2938_,
		_w2982_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		_w2907_,
		_w2938_,
		_w2983_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h8)
	) name1805 (
		_w2852_,
		_w2984_,
		_w2985_
	);
	LUT2 #(
		.INIT('h2)
	) name1806 (
		_w2877_,
		_w2929_,
		_w2986_
	);
	LUT2 #(
		.INIT('h4)
	) name1807 (
		_w2877_,
		_w2929_,
		_w2987_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		_w2852_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h2)
	) name1810 (
		_w2892_,
		_w2938_,
		_w2990_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w2892_,
		_w2938_,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w2990_,
		_w2991_,
		_w2992_
	);
	LUT2 #(
		.INIT('h2)
	) name1813 (
		_w2989_,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		_w2852_,
		_w2992_,
		_w2994_
	);
	LUT2 #(
		.INIT('h4)
	) name1815 (
		_w2988_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h1)
	) name1816 (
		_w2993_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('h2)
	) name1817 (
		_w2862_,
		_w2929_,
		_w2997_
	);
	LUT2 #(
		.INIT('h4)
	) name1818 (
		_w2862_,
		_w2929_,
		_w2998_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		_w2997_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h8)
	) name1820 (
		_w2852_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h2)
	) name1821 (
		_w2996_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h4)
	) name1822 (
		_w2996_,
		_w3000_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name1823 (
		_w3001_,
		_w3002_,
		_w3003_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		_w2985_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h1)
	) name1825 (
		_w2985_,
		_w3003_,
		_w3005_
	);
	LUT2 #(
		.INIT('h1)
	) name1826 (
		_w3004_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h8)
	) name1827 (
		_w2981_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h1)
	) name1828 (
		_w2981_,
		_w3006_,
		_w3008_
	);
	LUT2 #(
		.INIT('h2)
	) name1829 (
		\g1196_reg/NET0131 ,
		_w3007_,
		_w3009_
	);
	LUT2 #(
		.INIT('h4)
	) name1830 (
		_w3008_,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h1)
	) name1831 (
		_w2947_,
		_w2953_,
		_w3011_
	);
	LUT2 #(
		.INIT('h4)
	) name1832 (
		_w3010_,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('h2)
	) name1833 (
		\g1018_reg/NET0131 ,
		\g2116_reg/NET0131 ,
		_w3013_
	);
	LUT2 #(
		.INIT('h2)
	) name1834 (
		\g1024_reg/NET0131 ,
		\g2114_reg/NET0131 ,
		_w3014_
	);
	LUT2 #(
		.INIT('h4)
	) name1835 (
		\g2115_reg/NET0131 ,
		\g5657_pad ,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name1836 (
		_w3013_,
		_w3014_,
		_w3016_
	);
	LUT2 #(
		.INIT('h4)
	) name1837 (
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h4)
	) name1838 (
		_w1816_,
		_w3017_,
		_w3018_
	);
	LUT2 #(
		.INIT('h2)
	) name1839 (
		\g1880_reg/NET0131 ,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h2)
	) name1840 (
		_w1739_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w1901_,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name1842 (
		_w1837_,
		_w1911_,
		_w3022_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w1837_,
		_w1871_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name1844 (
		_w1837_,
		_w1901_,
		_w3024_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		\g1910_reg/NET0131 ,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		_w1739_,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w3022_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h4)
	) name1848 (
		_w3023_,
		_w3027_,
		_w3028_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		_w3021_,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('h8)
	) name1850 (
		_w1739_,
		_w3019_,
		_w3030_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		_w1901_,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		\g1909_reg/NET0131 ,
		_w3024_,
		_w3032_
	);
	LUT2 #(
		.INIT('h8)
	) name1853 (
		_w1739_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h4)
	) name1854 (
		_w1837_,
		_w1888_,
		_w3034_
	);
	LUT2 #(
		.INIT('h1)
	) name1855 (
		_w3022_,
		_w3033_,
		_w3035_
	);
	LUT2 #(
		.INIT('h4)
	) name1856 (
		_w3034_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h1)
	) name1857 (
		_w3031_,
		_w3036_,
		_w3037_
	);
	LUT2 #(
		.INIT('h4)
	) name1858 (
		_w1837_,
		_w1882_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name1859 (
		\g1911_reg/NET0131 ,
		_w3024_,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name1860 (
		_w1739_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name1861 (
		_w3022_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h4)
	) name1862 (
		_w3038_,
		_w3041_,
		_w3042_
	);
	LUT2 #(
		.INIT('h1)
	) name1863 (
		_w3021_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h4)
	) name1864 (
		_w1837_,
		_w1877_,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		\g1912_reg/NET0131 ,
		_w3024_,
		_w3045_
	);
	LUT2 #(
		.INIT('h8)
	) name1866 (
		_w1739_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w3022_,
		_w3046_,
		_w3047_
	);
	LUT2 #(
		.INIT('h4)
	) name1868 (
		_w3044_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w3031_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h4)
	) name1870 (
		_w1739_,
		_w1901_,
		_w3050_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		_w1846_,
		_w3024_,
		_w3051_
	);
	LUT2 #(
		.INIT('h1)
	) name1872 (
		\g1913_reg/NET0131 ,
		_w3024_,
		_w3052_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		_w1739_,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h1)
	) name1874 (
		_w3022_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h4)
	) name1875 (
		_w3051_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		_w3050_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h8)
	) name1877 (
		_w1852_,
		_w3024_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name1878 (
		\g1914_reg/NET0131 ,
		_w3024_,
		_w3058_
	);
	LUT2 #(
		.INIT('h8)
	) name1879 (
		_w1739_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h1)
	) name1880 (
		_w3022_,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h4)
	) name1881 (
		_w3057_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		_w3050_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h8)
	) name1883 (
		_w2238_,
		_w2252_,
		_w3063_
	);
	LUT2 #(
		.INIT('h2)
	) name1884 (
		_w2117_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h4)
	) name1885 (
		_w2019_,
		_w2024_,
		_w3065_
	);
	LUT2 #(
		.INIT('h4)
	) name1886 (
		_w3064_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name1887 (
		_w2014_,
		_w2136_,
		_w3067_
	);
	LUT2 #(
		.INIT('h8)
	) name1888 (
		_w3066_,
		_w3067_,
		_w3068_
	);
	LUT2 #(
		.INIT('h8)
	) name1889 (
		\g1563_reg/NET0131 ,
		_w2116_,
		_w3069_
	);
	LUT2 #(
		.INIT('h2)
	) name1890 (
		_w2014_,
		_w2024_,
		_w3070_
	);
	LUT2 #(
		.INIT('h8)
	) name1891 (
		_w2136_,
		_w3070_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name1892 (
		_w3069_,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h1)
	) name1893 (
		_w2019_,
		_w3072_,
		_w3073_
	);
	LUT2 #(
		.INIT('h1)
	) name1894 (
		_w2265_,
		_w3073_,
		_w3074_
	);
	LUT2 #(
		.INIT('h4)
	) name1895 (
		_w3068_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h4)
	) name1896 (
		_w2014_,
		_w2266_,
		_w3076_
	);
	LUT2 #(
		.INIT('h4)
	) name1897 (
		_w2192_,
		_w3076_,
		_w3077_
	);
	LUT2 #(
		.INIT('h8)
	) name1898 (
		_w2175_,
		_w2209_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		_w2150_,
		_w2167_,
		_w3079_
	);
	LUT2 #(
		.INIT('h8)
	) name1900 (
		_w2200_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h8)
	) name1901 (
		_w3078_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h1)
	) name1902 (
		_w2142_,
		_w2159_,
		_w3082_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w2184_,
		_w2217_,
		_w3083_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h8)
	) name1905 (
		_w3077_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h8)
	) name1906 (
		_w3081_,
		_w3085_,
		_w3086_
	);
	LUT2 #(
		.INIT('h8)
	) name1907 (
		_w2014_,
		_w2184_,
		_w3087_
	);
	LUT2 #(
		.INIT('h8)
	) name1908 (
		_w2142_,
		_w2159_,
		_w3088_
	);
	LUT2 #(
		.INIT('h8)
	) name1909 (
		_w2192_,
		_w2217_,
		_w3089_
	);
	LUT2 #(
		.INIT('h8)
	) name1910 (
		_w3088_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w3087_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name1912 (
		_w3081_,
		_w3091_,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		_w3086_,
		_w3092_,
		_w3093_
	);
	LUT2 #(
		.INIT('h2)
	) name1914 (
		_w2266_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h8)
	) name1915 (
		_w3075_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h4)
	) name1916 (
		_w2014_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h2)
	) name1917 (
		_w3075_,
		_w3086_,
		_w3097_
	);
	LUT2 #(
		.INIT('h1)
	) name1918 (
		\g105_reg/NET0131 ,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		_w3075_,
		_w3094_,
		_w3099_
	);
	LUT2 #(
		.INIT('h1)
	) name1920 (
		_w2014_,
		_w2184_,
		_w3100_
	);
	LUT2 #(
		.INIT('h1)
	) name1921 (
		_w3087_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h4)
	) name1922 (
		_w2014_,
		_w2167_,
		_w3102_
	);
	LUT2 #(
		.INIT('h2)
	) name1923 (
		_w2014_,
		_w2167_,
		_w3103_
	);
	LUT2 #(
		.INIT('h2)
	) name1924 (
		_w2266_,
		_w3102_,
		_w3104_
	);
	LUT2 #(
		.INIT('h4)
	) name1925 (
		_w3103_,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('h4)
	) name1926 (
		_w3101_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h1)
	) name1927 (
		_w2192_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		_w2192_,
		_w3106_,
		_w3108_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		_w3107_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name1930 (
		_w3099_,
		_w3109_,
		_w3110_
	);
	LUT2 #(
		.INIT('h1)
	) name1931 (
		_w3096_,
		_w3098_,
		_w3111_
	);
	LUT2 #(
		.INIT('h4)
	) name1932 (
		_w3110_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		\g7961_pad ,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name1934 (
		\g195_reg/NET0131 ,
		\g7961_pad ,
		_w3114_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w3113_,
		_w3114_,
		_w3115_
	);
	LUT2 #(
		.INIT('h2)
	) name1936 (
		\g1092_reg/NET0131 ,
		_w3112_,
		_w3116_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		\g1092_reg/NET0131 ,
		\g198_reg/NET0131 ,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name1938 (
		_w3116_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h2)
	) name1939 (
		\g1088_reg/NET0131 ,
		_w3112_,
		_w3119_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		\g1088_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name1941 (
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h8)
	) name1942 (
		_w2413_,
		_w2452_,
		_w3122_
	);
	LUT2 #(
		.INIT('h8)
	) name1943 (
		_w2436_,
		_w2500_,
		_w3123_
	);
	LUT2 #(
		.INIT('h8)
	) name1944 (
		_w2444_,
		_w2491_,
		_w3124_
	);
	LUT2 #(
		.INIT('h8)
	) name1945 (
		_w2510_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h8)
	) name1946 (
		_w3123_,
		_w3125_,
		_w3126_
	);
	LUT2 #(
		.INIT('h8)
	) name1947 (
		_w2419_,
		_w2427_,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name1948 (
		_w2474_,
		_w2482_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name1949 (
		_w3127_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h8)
	) name1950 (
		_w3122_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		_w3126_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h4)
	) name1952 (
		_w2413_,
		_w2550_,
		_w3132_
	);
	LUT2 #(
		.INIT('h4)
	) name1953 (
		_w2474_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h1)
	) name1954 (
		_w2419_,
		_w2427_,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name1955 (
		_w2452_,
		_w2482_,
		_w3135_
	);
	LUT2 #(
		.INIT('h8)
	) name1956 (
		_w3134_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		_w3126_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h8)
	) name1958 (
		_w3133_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name1959 (
		_w3131_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h4)
	) name1960 (
		_w2288_,
		_w2413_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name1961 (
		_w2401_,
		_w3140_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name1962 (
		_w2408_,
		_w3141_,
		_w3142_
	);
	LUT2 #(
		.INIT('h4)
	) name1963 (
		_w2402_,
		_w3142_,
		_w3143_
	);
	LUT2 #(
		.INIT('h1)
	) name1964 (
		_w2469_,
		_w2524_,
		_w3144_
	);
	LUT2 #(
		.INIT('h8)
	) name1965 (
		_w2288_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('h8)
	) name1966 (
		_w2400_,
		_w2414_,
		_w3146_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		_w3145_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name1968 (
		_w2543_,
		_w3143_,
		_w3148_
	);
	LUT2 #(
		.INIT('h4)
	) name1969 (
		_w3147_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h2)
	) name1970 (
		_w3132_,
		_w3139_,
		_w3150_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		_w3149_,
		_w3150_,
		_w3151_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		\g793_reg/NET0131 ,
		_w3149_,
		_w3152_
	);
	LUT2 #(
		.INIT('h2)
	) name1973 (
		_w2550_,
		_w3139_,
		_w3153_
	);
	LUT2 #(
		.INIT('h2)
	) name1974 (
		_w3149_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h2)
	) name1975 (
		_w2413_,
		_w2510_,
		_w3155_
	);
	LUT2 #(
		.INIT('h2)
	) name1976 (
		_w2550_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w2452_,
		_w2510_,
		_w3157_
	);
	LUT2 #(
		.INIT('h1)
	) name1978 (
		_w3122_,
		_w3157_,
		_w3158_
	);
	LUT2 #(
		.INIT('h2)
	) name1979 (
		_w3156_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		_w2474_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		_w2474_,
		_w3159_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w3160_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		_w3154_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h1)
	) name1984 (
		_w3151_,
		_w3152_,
		_w3164_
	);
	LUT2 #(
		.INIT('h4)
	) name1985 (
		_w3163_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h2)
	) name1986 (
		\g7961_pad ,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h1)
	) name1987 (
		\g7961_pad ,
		\g882_reg/NET0131 ,
		_w3167_
	);
	LUT2 #(
		.INIT('h1)
	) name1988 (
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		\g1092_reg/NET0131 ,
		_w3165_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		\g1092_reg/NET0131 ,
		\g885_reg/NET0131 ,
		_w3170_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w3169_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h2)
	) name1992 (
		\g1088_reg/NET0131 ,
		_w3165_,
		_w3172_
	);
	LUT2 #(
		.INIT('h1)
	) name1993 (
		\g1088_reg/NET0131 ,
		\g888_reg/NET0131 ,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name1994 (
		_w3172_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name1995 (
		\g789_reg/NET0131 ,
		_w3149_,
		_w3175_
	);
	LUT2 #(
		.INIT('h8)
	) name1996 (
		_w2510_,
		_w2550_,
		_w3176_
	);
	LUT2 #(
		.INIT('h4)
	) name1997 (
		_w2413_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		_w3156_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		_w2452_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		_w2452_,
		_w3178_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name2001 (
		_w3179_,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h8)
	) name2002 (
		_w3154_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		_w3151_,
		_w3175_,
		_w3183_
	);
	LUT2 #(
		.INIT('h4)
	) name2004 (
		_w3182_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h2)
	) name2005 (
		\g7961_pad ,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h1)
	) name2006 (
		\g7961_pad ,
		\g918_reg/NET0131 ,
		_w3186_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		\g1092_reg/NET0131 ,
		_w3184_,
		_w3188_
	);
	LUT2 #(
		.INIT('h1)
	) name2009 (
		\g1092_reg/NET0131 ,
		\g921_reg/NET0131 ,
		_w3189_
	);
	LUT2 #(
		.INIT('h1)
	) name2010 (
		_w3188_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h2)
	) name2011 (
		\g1088_reg/NET0131 ,
		_w3184_,
		_w3191_
	);
	LUT2 #(
		.INIT('h1)
	) name2012 (
		\g1088_reg/NET0131 ,
		\g924_reg/NET0131 ,
		_w3192_
	);
	LUT2 #(
		.INIT('h1)
	) name2013 (
		_w3191_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h1)
	) name2014 (
		\g797_reg/NET0131 ,
		_w3149_,
		_w3194_
	);
	LUT2 #(
		.INIT('h2)
	) name2015 (
		_w2474_,
		_w3132_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w3133_,
		_w3195_,
		_w3196_
	);
	LUT2 #(
		.INIT('h2)
	) name2017 (
		_w3159_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name2018 (
		_w2419_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h8)
	) name2019 (
		_w2419_,
		_w3197_,
		_w3199_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w3198_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		_w3154_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name2022 (
		_w3151_,
		_w3194_,
		_w3202_
	);
	LUT2 #(
		.INIT('h4)
	) name2023 (
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT2 #(
		.INIT('h2)
	) name2024 (
		\g7961_pad ,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h1)
	) name2025 (
		\g7961_pad ,
		\g927_reg/NET0131 ,
		_w3205_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		_w3204_,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('h2)
	) name2027 (
		\g1088_reg/NET0131 ,
		_w3203_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		\g1088_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w3208_
	);
	LUT2 #(
		.INIT('h1)
	) name2029 (
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h2)
	) name2030 (
		\g1092_reg/NET0131 ,
		_w3203_,
		_w3210_
	);
	LUT2 #(
		.INIT('h1)
	) name2031 (
		\g1092_reg/NET0131 ,
		\g930_reg/NET0131 ,
		_w3211_
	);
	LUT2 #(
		.INIT('h1)
	) name2032 (
		_w3210_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h2)
	) name2033 (
		_w2298_,
		_w3149_,
		_w3213_
	);
	LUT2 #(
		.INIT('h4)
	) name2034 (
		_w2500_,
		_w3132_,
		_w3214_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w3123_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		_w2419_,
		_w3132_,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name2037 (
		_w2419_,
		_w3132_,
		_w3217_
	);
	LUT2 #(
		.INIT('h1)
	) name2038 (
		_w3216_,
		_w3217_,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		_w3197_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name2040 (
		_w2491_,
		_w3132_,
		_w3220_
	);
	LUT2 #(
		.INIT('h8)
	) name2041 (
		_w2491_,
		_w3132_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name2042 (
		_w3220_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h8)
	) name2043 (
		_w3219_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h2)
	) name2044 (
		_w2436_,
		_w2491_,
		_w3224_
	);
	LUT2 #(
		.INIT('h2)
	) name2045 (
		_w3223_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('h4)
	) name2046 (
		_w3215_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h1)
	) name2047 (
		_w2444_,
		_w3132_,
		_w3227_
	);
	LUT2 #(
		.INIT('h8)
	) name2048 (
		_w2444_,
		_w3132_,
		_w3228_
	);
	LUT2 #(
		.INIT('h1)
	) name2049 (
		_w3227_,
		_w3228_,
		_w3229_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		_w3226_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('h1)
	) name2051 (
		_w2482_,
		_w3132_,
		_w3231_
	);
	LUT2 #(
		.INIT('h8)
	) name2052 (
		_w2482_,
		_w3132_,
		_w3232_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w3231_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w3230_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h1)
	) name2055 (
		_w2427_,
		_w3234_,
		_w3235_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		_w2427_,
		_w3234_,
		_w3236_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		_w3235_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h8)
	) name2058 (
		_w3154_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w3151_,
		_w3213_,
		_w3239_
	);
	LUT2 #(
		.INIT('h4)
	) name2060 (
		_w3238_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h2)
	) name2061 (
		\g7961_pad ,
		_w3240_,
		_w3241_
	);
	LUT2 #(
		.INIT('h1)
	) name2062 (
		\g7961_pad ,
		\g954_reg/NET0131 ,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		\g1092_reg/NET0131 ,
		_w3240_,
		_w3244_
	);
	LUT2 #(
		.INIT('h1)
	) name2065 (
		\g1092_reg/NET0131 ,
		\g957_reg/NET0131 ,
		_w3245_
	);
	LUT2 #(
		.INIT('h1)
	) name2066 (
		_w3244_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\g1088_reg/NET0131 ,
		_w3240_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name2068 (
		\g1088_reg/NET0131 ,
		\g960_reg/NET0131 ,
		_w3248_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		_w3247_,
		_w3248_,
		_w3249_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		_w2684_,
		_w2720_,
		_w3250_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		_w2593_,
		_w2645_,
		_w3251_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		_w2602_,
		_w2653_,
		_w3252_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		_w2585_,
		_w2624_,
		_w3253_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		_w2662_,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		_w3252_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('h8)
	) name2076 (
		_w2615_,
		_w2675_,
		_w3256_
	);
	LUT2 #(
		.INIT('h8)
	) name2077 (
		_w3250_,
		_w3256_,
		_w3257_
	);
	LUT2 #(
		.INIT('h8)
	) name2078 (
		_w3251_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h8)
	) name2079 (
		_w3255_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('h4)
	) name2080 (
		_w2720_,
		_w2836_,
		_w3260_
	);
	LUT2 #(
		.INIT('h4)
	) name2081 (
		_w2615_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h1)
	) name2082 (
		_w2593_,
		_w2645_,
		_w3262_
	);
	LUT2 #(
		.INIT('h1)
	) name2083 (
		_w2675_,
		_w2684_,
		_w3263_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		_w3262_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		_w3255_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		_w3261_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h1)
	) name2087 (
		_w3259_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('h4)
	) name2088 (
		_w2699_,
		_w2720_,
		_w3268_
	);
	LUT2 #(
		.INIT('h1)
	) name2089 (
		_w2818_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name2090 (
		_w2574_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h4)
	) name2091 (
		_w2819_,
		_w3270_,
		_w3271_
	);
	LUT2 #(
		.INIT('h1)
	) name2092 (
		_w2640_,
		_w2824_,
		_w3272_
	);
	LUT2 #(
		.INIT('h4)
	) name2093 (
		_w2574_,
		_w2699_,
		_w3273_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		_w2816_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h8)
	) name2095 (
		_w3272_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h2)
	) name2096 (
		_w2720_,
		_w2726_,
		_w3276_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h1)
	) name2098 (
		_w2835_,
		_w3271_,
		_w3278_
	);
	LUT2 #(
		.INIT('h4)
	) name2099 (
		_w3277_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		_w3260_,
		_w3267_,
		_w3280_
	);
	LUT2 #(
		.INIT('h8)
	) name2101 (
		_w3279_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h1)
	) name2102 (
		\g1481_reg/NET0131 ,
		_w3279_,
		_w3282_
	);
	LUT2 #(
		.INIT('h2)
	) name2103 (
		_w2836_,
		_w3267_,
		_w3283_
	);
	LUT2 #(
		.INIT('h2)
	) name2104 (
		_w3279_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('h4)
	) name2105 (
		_w2624_,
		_w2720_,
		_w3285_
	);
	LUT2 #(
		.INIT('h2)
	) name2106 (
		_w2836_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w2624_,
		_w2684_,
		_w3287_
	);
	LUT2 #(
		.INIT('h1)
	) name2108 (
		_w3250_,
		_w3287_,
		_w3288_
	);
	LUT2 #(
		.INIT('h2)
	) name2109 (
		_w3286_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w2593_,
		_w3289_,
		_w3290_
	);
	LUT2 #(
		.INIT('h8)
	) name2111 (
		_w2593_,
		_w3289_,
		_w3291_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w3290_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		_w3284_,
		_w3292_,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w3281_,
		_w3282_,
		_w3294_
	);
	LUT2 #(
		.INIT('h4)
	) name2115 (
		_w3293_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h2)
	) name2116 (
		\g7961_pad ,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h1)
	) name2117 (
		\g1576_reg/NET0131 ,
		\g7961_pad ,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2118 (
		_w3296_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h8)
	) name2119 (
		_w1309_,
		_w1355_,
		_w3299_
	);
	LUT2 #(
		.INIT('h8)
	) name2120 (
		_w1338_,
		_w1392_,
		_w3300_
	);
	LUT2 #(
		.INIT('h8)
	) name2121 (
		_w1330_,
		_w1376_,
		_w3301_
	);
	LUT2 #(
		.INIT('h8)
	) name2122 (
		_w1409_,
		_w3301_,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		_w3300_,
		_w3302_,
		_w3303_
	);
	LUT2 #(
		.INIT('h8)
	) name2124 (
		_w1322_,
		_w1347_,
		_w3304_
	);
	LUT2 #(
		.INIT('h8)
	) name2125 (
		_w1384_,
		_w1401_,
		_w3305_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		_w3304_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		_w3299_,
		_w3306_,
		_w3307_
	);
	LUT2 #(
		.INIT('h8)
	) name2128 (
		_w3303_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		_w1304_,
		_w1309_,
		_w3309_
	);
	LUT2 #(
		.INIT('h4)
	) name2130 (
		_w1384_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		_w1322_,
		_w1347_,
		_w3311_
	);
	LUT2 #(
		.INIT('h1)
	) name2132 (
		_w1355_,
		_w1401_,
		_w3312_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		_w3311_,
		_w3312_,
		_w3313_
	);
	LUT2 #(
		.INIT('h8)
	) name2134 (
		_w3303_,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h8)
	) name2135 (
		_w3310_,
		_w3314_,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		_w3308_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		\g1563_reg/NET0131 ,
		_w1281_,
		_w3317_
	);
	LUT2 #(
		.INIT('h4)
	) name2138 (
		_w1303_,
		_w3317_,
		_w3318_
	);
	LUT2 #(
		.INIT('h4)
	) name2139 (
		_w1298_,
		_w1309_,
		_w3319_
	);
	LUT2 #(
		.INIT('h4)
	) name2140 (
		_w1303_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h8)
	) name2141 (
		_w1316_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		_w1371_,
		_w1432_,
		_w3322_
	);
	LUT2 #(
		.INIT('h2)
	) name2143 (
		_w1282_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h2)
	) name2144 (
		_w1298_,
		_w1303_,
		_w3324_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		_w1292_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h4)
	) name2146 (
		_w3323_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h2)
	) name2147 (
		_w1309_,
		_w1315_,
		_w3327_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		_w3326_,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w1293_,
		_w3318_,
		_w3329_
	);
	LUT2 #(
		.INIT('h4)
	) name2150 (
		_w3321_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h4)
	) name2151 (
		_w3328_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		_w3309_,
		_w3316_,
		_w3332_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		_w3331_,
		_w3332_,
		_w3333_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		\g2175_reg/NET0131 ,
		_w3331_,
		_w3334_
	);
	LUT2 #(
		.INIT('h2)
	) name2155 (
		_w1304_,
		_w3316_,
		_w3335_
	);
	LUT2 #(
		.INIT('h2)
	) name2156 (
		_w3331_,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h2)
	) name2157 (
		_w1309_,
		_w1409_,
		_w3337_
	);
	LUT2 #(
		.INIT('h2)
	) name2158 (
		_w1304_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name2159 (
		_w1355_,
		_w1409_,
		_w3339_
	);
	LUT2 #(
		.INIT('h1)
	) name2160 (
		_w3299_,
		_w3339_,
		_w3340_
	);
	LUT2 #(
		.INIT('h2)
	) name2161 (
		_w3338_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h1)
	) name2162 (
		_w1401_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		_w1401_,
		_w3341_,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name2164 (
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT2 #(
		.INIT('h8)
	) name2165 (
		_w3336_,
		_w3344_,
		_w3345_
	);
	LUT2 #(
		.INIT('h1)
	) name2166 (
		_w3333_,
		_w3334_,
		_w3346_
	);
	LUT2 #(
		.INIT('h4)
	) name2167 (
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h2)
	) name2168 (
		\g7961_pad ,
		_w3347_,
		_w3348_
	);
	LUT2 #(
		.INIT('h1)
	) name2169 (
		\g2270_reg/NET0131 ,
		\g7961_pad ,
		_w3349_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h2)
	) name2171 (
		\g1088_reg/NET0131 ,
		_w3347_,
		_w3351_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		\g1088_reg/NET0131 ,
		\g2276_reg/NET0131 ,
		_w3352_
	);
	LUT2 #(
		.INIT('h1)
	) name2173 (
		_w3351_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h2)
	) name2174 (
		\g1092_reg/NET0131 ,
		_w3347_,
		_w3354_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		\g1092_reg/NET0131 ,
		\g2273_reg/NET0131 ,
		_w3355_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h2)
	) name2177 (
		\g1092_reg/NET0131 ,
		_w3295_,
		_w3357_
	);
	LUT2 #(
		.INIT('h1)
	) name2178 (
		\g1092_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		_w3358_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w3357_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		\g2170_reg/NET0131 ,
		_w3331_,
		_w3360_
	);
	LUT2 #(
		.INIT('h2)
	) name2181 (
		_w1304_,
		_w1409_,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w1309_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h2)
	) name2183 (
		_w3338_,
		_w3362_,
		_w3363_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		_w1355_,
		_w3363_,
		_w3364_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		_w1355_,
		_w3363_,
		_w3365_
	);
	LUT2 #(
		.INIT('h1)
	) name2186 (
		_w3364_,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		_w3336_,
		_w3366_,
		_w3367_
	);
	LUT2 #(
		.INIT('h1)
	) name2188 (
		_w3333_,
		_w3360_,
		_w3368_
	);
	LUT2 #(
		.INIT('h4)
	) name2189 (
		_w3367_,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('h2)
	) name2190 (
		\g7961_pad ,
		_w3369_,
		_w3370_
	);
	LUT2 #(
		.INIT('h1)
	) name2191 (
		\g2306_reg/NET0131 ,
		\g7961_pad ,
		_w3371_
	);
	LUT2 #(
		.INIT('h1)
	) name2192 (
		_w3370_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h2)
	) name2193 (
		\g1088_reg/NET0131 ,
		_w3295_,
		_w3373_
	);
	LUT2 #(
		.INIT('h1)
	) name2194 (
		\g1088_reg/NET0131 ,
		\g1582_reg/NET0131 ,
		_w3374_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w3373_,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h2)
	) name2196 (
		\g1092_reg/NET0131 ,
		_w3369_,
		_w3376_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		\g1092_reg/NET0131 ,
		\g2309_reg/NET0131 ,
		_w3377_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		_w3376_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h2)
	) name2199 (
		\g1088_reg/NET0131 ,
		_w3369_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name2200 (
		\g1088_reg/NET0131 ,
		\g2312_reg/NET0131 ,
		_w3380_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w3379_,
		_w3380_,
		_w3381_
	);
	LUT2 #(
		.INIT('h1)
	) name2202 (
		\g2180_reg/NET0131 ,
		_w3331_,
		_w3382_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w1401_,
		_w3309_,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name2204 (
		_w1401_,
		_w3309_,
		_w3384_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		_w3341_,
		_w3383_,
		_w3385_
	);
	LUT2 #(
		.INIT('h4)
	) name2206 (
		_w3384_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		_w1347_,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h8)
	) name2208 (
		_w1347_,
		_w3386_,
		_w3388_
	);
	LUT2 #(
		.INIT('h1)
	) name2209 (
		_w3387_,
		_w3388_,
		_w3389_
	);
	LUT2 #(
		.INIT('h8)
	) name2210 (
		_w3336_,
		_w3389_,
		_w3390_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w3333_,
		_w3382_,
		_w3391_
	);
	LUT2 #(
		.INIT('h4)
	) name2212 (
		_w3390_,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h2)
	) name2213 (
		\g7961_pad ,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h1)
	) name2214 (
		\g2315_reg/NET0131 ,
		\g7961_pad ,
		_w3394_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		_w3393_,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		\g1092_reg/NET0131 ,
		_w3392_,
		_w3396_
	);
	LUT2 #(
		.INIT('h1)
	) name2217 (
		\g1092_reg/NET0131 ,
		\g2318_reg/NET0131 ,
		_w3397_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name2219 (
		\g101_reg/NET0131 ,
		_w3097_,
		_w3399_
	);
	LUT2 #(
		.INIT('h1)
	) name2220 (
		_w2184_,
		_w3105_,
		_w3400_
	);
	LUT2 #(
		.INIT('h8)
	) name2221 (
		_w2184_,
		_w3105_,
		_w3401_
	);
	LUT2 #(
		.INIT('h1)
	) name2222 (
		_w3400_,
		_w3401_,
		_w3402_
	);
	LUT2 #(
		.INIT('h8)
	) name2223 (
		_w3099_,
		_w3402_,
		_w3403_
	);
	LUT2 #(
		.INIT('h1)
	) name2224 (
		_w3096_,
		_w3399_,
		_w3404_
	);
	LUT2 #(
		.INIT('h4)
	) name2225 (
		_w3403_,
		_w3404_,
		_w3405_
	);
	LUT2 #(
		.INIT('h2)
	) name2226 (
		\g7961_pad ,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		\g231_reg/NET0131 ,
		\g7961_pad ,
		_w3407_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT2 #(
		.INIT('h2)
	) name2229 (
		\g1088_reg/NET0131 ,
		_w3392_,
		_w3409_
	);
	LUT2 #(
		.INIT('h1)
	) name2230 (
		\g1088_reg/NET0131 ,
		\g2321_reg/NET0131 ,
		_w3410_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		_w3409_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h2)
	) name2232 (
		_w1268_,
		_w3331_,
		_w3412_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w1338_,
		_w1392_,
		_w3413_
	);
	LUT2 #(
		.INIT('h1)
	) name2234 (
		_w3300_,
		_w3413_,
		_w3414_
	);
	LUT2 #(
		.INIT('h4)
	) name2235 (
		_w1347_,
		_w3309_,
		_w3415_
	);
	LUT2 #(
		.INIT('h1)
	) name2236 (
		_w1376_,
		_w3415_,
		_w3416_
	);
	LUT2 #(
		.INIT('h2)
	) name2237 (
		_w1347_,
		_w3309_,
		_w3417_
	);
	LUT2 #(
		.INIT('h2)
	) name2238 (
		_w1376_,
		_w3417_,
		_w3418_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w3416_,
		_w3418_,
		_w3419_
	);
	LUT2 #(
		.INIT('h8)
	) name2240 (
		_w3386_,
		_w3419_,
		_w3420_
	);
	LUT2 #(
		.INIT('h1)
	) name2241 (
		_w1330_,
		_w3309_,
		_w3421_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		_w1330_,
		_w3309_,
		_w3422_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		_w3421_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h8)
	) name2244 (
		_w3420_,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('h1)
	) name2245 (
		_w1392_,
		_w3309_,
		_w3425_
	);
	LUT2 #(
		.INIT('h8)
	) name2246 (
		_w1392_,
		_w3309_,
		_w3426_
	);
	LUT2 #(
		.INIT('h1)
	) name2247 (
		_w3425_,
		_w3426_,
		_w3427_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		_w3424_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name2249 (
		_w3414_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h2)
	) name2250 (
		_w1384_,
		_w3309_,
		_w3430_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		_w3310_,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		_w3429_,
		_w3431_,
		_w3432_
	);
	LUT2 #(
		.INIT('h1)
	) name2253 (
		_w1322_,
		_w3432_,
		_w3433_
	);
	LUT2 #(
		.INIT('h8)
	) name2254 (
		_w1322_,
		_w3432_,
		_w3434_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w3433_,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		_w3336_,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h1)
	) name2257 (
		_w3333_,
		_w3412_,
		_w3437_
	);
	LUT2 #(
		.INIT('h4)
	) name2258 (
		_w3436_,
		_w3437_,
		_w3438_
	);
	LUT2 #(
		.INIT('h2)
	) name2259 (
		\g7961_pad ,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h1)
	) name2260 (
		\g2342_reg/NET0131 ,
		\g7961_pad ,
		_w3440_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		_w3439_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h2)
	) name2262 (
		\g1092_reg/NET0131 ,
		_w3438_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name2263 (
		\g1092_reg/NET0131 ,
		\g2345_reg/NET0131 ,
		_w3443_
	);
	LUT2 #(
		.INIT('h1)
	) name2264 (
		_w3442_,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h2)
	) name2265 (
		\g1088_reg/NET0131 ,
		_w3438_,
		_w3445_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		\g1088_reg/NET0131 ,
		\g2348_reg/NET0131 ,
		_w3446_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		_w3445_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('h2)
	) name2268 (
		\g1092_reg/NET0131 ,
		_w3405_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name2269 (
		\g1092_reg/NET0131 ,
		\g234_reg/NET0131 ,
		_w3449_
	);
	LUT2 #(
		.INIT('h1)
	) name2270 (
		_w3448_,
		_w3449_,
		_w3450_
	);
	LUT2 #(
		.INIT('h2)
	) name2271 (
		\g1088_reg/NET0131 ,
		_w3405_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name2272 (
		\g1088_reg/NET0131 ,
		\g237_reg/NET0131 ,
		_w3452_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w3451_,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		\g1476_reg/NET0131 ,
		_w3279_,
		_w3454_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		_w2624_,
		_w2836_,
		_w3455_
	);
	LUT2 #(
		.INIT('h4)
	) name2276 (
		_w2720_,
		_w3455_,
		_w3456_
	);
	LUT2 #(
		.INIT('h2)
	) name2277 (
		_w3286_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w2684_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w2684_,
		_w3457_,
		_w3459_
	);
	LUT2 #(
		.INIT('h1)
	) name2280 (
		_w3458_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		_w3284_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w3281_,
		_w3454_,
		_w3462_
	);
	LUT2 #(
		.INIT('h4)
	) name2283 (
		_w3461_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name2284 (
		\g7961_pad ,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h1)
	) name2285 (
		\g1612_reg/NET0131 ,
		\g7961_pad ,
		_w3465_
	);
	LUT2 #(
		.INIT('h1)
	) name2286 (
		_w3464_,
		_w3465_,
		_w3466_
	);
	LUT2 #(
		.INIT('h2)
	) name2287 (
		\g1092_reg/NET0131 ,
		_w3463_,
		_w3467_
	);
	LUT2 #(
		.INIT('h1)
	) name2288 (
		\g1092_reg/NET0131 ,
		\g1615_reg/NET0131 ,
		_w3468_
	);
	LUT2 #(
		.INIT('h1)
	) name2289 (
		_w3467_,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h2)
	) name2290 (
		\g1088_reg/NET0131 ,
		_w3463_,
		_w3470_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		\g1088_reg/NET0131 ,
		\g1618_reg/NET0131 ,
		_w3471_
	);
	LUT2 #(
		.INIT('h1)
	) name2292 (
		_w3470_,
		_w3471_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		\g1486_reg/NET0131 ,
		_w3279_,
		_w3473_
	);
	LUT2 #(
		.INIT('h1)
	) name2294 (
		_w2593_,
		_w3260_,
		_w3474_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		_w2593_,
		_w3260_,
		_w3475_
	);
	LUT2 #(
		.INIT('h2)
	) name2296 (
		_w3289_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h4)
	) name2297 (
		_w3474_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		_w2645_,
		_w3477_,
		_w3478_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		_w2645_,
		_w3477_,
		_w3479_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w3478_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		_w3284_,
		_w3480_,
		_w3481_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		_w3281_,
		_w3473_,
		_w3482_
	);
	LUT2 #(
		.INIT('h4)
	) name2303 (
		_w3481_,
		_w3482_,
		_w3483_
	);
	LUT2 #(
		.INIT('h2)
	) name2304 (
		\g7961_pad ,
		_w3483_,
		_w3484_
	);
	LUT2 #(
		.INIT('h1)
	) name2305 (
		\g1621_reg/NET0131 ,
		\g7961_pad ,
		_w3485_
	);
	LUT2 #(
		.INIT('h1)
	) name2306 (
		_w3484_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h2)
	) name2307 (
		\g1092_reg/NET0131 ,
		_w3483_,
		_w3487_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		\g1092_reg/NET0131 ,
		\g1624_reg/NET0131 ,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		_w3487_,
		_w3488_,
		_w3489_
	);
	LUT2 #(
		.INIT('h2)
	) name2310 (
		_w2192_,
		_w3076_,
		_w3490_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		_w3077_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h2)
	) name2312 (
		_w3106_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		_w2217_,
		_w3492_,
		_w3493_
	);
	LUT2 #(
		.INIT('h8)
	) name2314 (
		_w2217_,
		_w3492_,
		_w3494_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w3493_,
		_w3494_,
		_w3495_
	);
	LUT2 #(
		.INIT('h8)
	) name2316 (
		_w3099_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h8)
	) name2317 (
		_w2014_,
		_w3075_,
		_w3497_
	);
	LUT2 #(
		.INIT('h1)
	) name2318 (
		\g109_reg/NET0131 ,
		_w3099_,
		_w3498_
	);
	LUT2 #(
		.INIT('h4)
	) name2319 (
		_w3497_,
		_w3498_,
		_w3499_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		_w3096_,
		_w3496_,
		_w3500_
	);
	LUT2 #(
		.INIT('h4)
	) name2321 (
		_w3499_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h2)
	) name2322 (
		\g7961_pad ,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		\g240_reg/NET0131 ,
		\g7961_pad ,
		_w3503_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		_w3502_,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h2)
	) name2325 (
		\g1088_reg/NET0131 ,
		_w3483_,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name2326 (
		\g1088_reg/NET0131 ,
		\g1627_reg/NET0131 ,
		_w3506_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w3505_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		\g1092_reg/NET0131 ,
		_w3501_,
		_w3508_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		\g1092_reg/NET0131 ,
		\g243_reg/NET0131 ,
		_w3509_
	);
	LUT2 #(
		.INIT('h1)
	) name2330 (
		_w3508_,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h2)
	) name2331 (
		_w2670_,
		_w3279_,
		_w3511_
	);
	LUT2 #(
		.INIT('h2)
	) name2332 (
		_w2615_,
		_w3260_,
		_w3512_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w3261_,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h4)
	) name2334 (
		_w2602_,
		_w3260_,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name2335 (
		_w3252_,
		_w3514_,
		_w3515_
	);
	LUT2 #(
		.INIT('h4)
	) name2336 (
		_w2645_,
		_w3260_,
		_w3516_
	);
	LUT2 #(
		.INIT('h1)
	) name2337 (
		_w3251_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		_w3476_,
		_w3517_,
		_w3518_
	);
	LUT2 #(
		.INIT('h1)
	) name2339 (
		_w2585_,
		_w3260_,
		_w3519_
	);
	LUT2 #(
		.INIT('h8)
	) name2340 (
		_w2585_,
		_w3260_,
		_w3520_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w3519_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h8)
	) name2342 (
		_w3518_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h8)
	) name2343 (
		_w2653_,
		_w3260_,
		_w3523_
	);
	LUT2 #(
		.INIT('h2)
	) name2344 (
		_w3522_,
		_w3523_,
		_w3524_
	);
	LUT2 #(
		.INIT('h4)
	) name2345 (
		_w3515_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h1)
	) name2346 (
		_w2662_,
		_w3260_,
		_w3526_
	);
	LUT2 #(
		.INIT('h8)
	) name2347 (
		_w2662_,
		_w3260_,
		_w3527_
	);
	LUT2 #(
		.INIT('h1)
	) name2348 (
		_w3526_,
		_w3527_,
		_w3528_
	);
	LUT2 #(
		.INIT('h8)
	) name2349 (
		_w3525_,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('h4)
	) name2350 (
		_w3513_,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h1)
	) name2351 (
		_w2675_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		_w2675_,
		_w3530_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w3531_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h8)
	) name2354 (
		_w3284_,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h1)
	) name2355 (
		_w3281_,
		_w3511_,
		_w3535_
	);
	LUT2 #(
		.INIT('h4)
	) name2356 (
		_w3534_,
		_w3535_,
		_w3536_
	);
	LUT2 #(
		.INIT('h2)
	) name2357 (
		\g1092_reg/NET0131 ,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h1)
	) name2358 (
		\g1092_reg/NET0131 ,
		\g1651_reg/NET0131 ,
		_w3538_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		_w3537_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h2)
	) name2360 (
		\g7961_pad ,
		_w3536_,
		_w3540_
	);
	LUT2 #(
		.INIT('h1)
	) name2361 (
		\g1648_reg/NET0131 ,
		\g7961_pad ,
		_w3541_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w3540_,
		_w3541_,
		_w3542_
	);
	LUT2 #(
		.INIT('h2)
	) name2363 (
		\g1088_reg/NET0131 ,
		_w3536_,
		_w3543_
	);
	LUT2 #(
		.INIT('h1)
	) name2364 (
		\g1088_reg/NET0131 ,
		\g1654_reg/NET0131 ,
		_w3544_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w3543_,
		_w3544_,
		_w3545_
	);
	LUT2 #(
		.INIT('h2)
	) name2366 (
		_w2034_,
		_w3097_,
		_w3546_
	);
	LUT2 #(
		.INIT('h1)
	) name2367 (
		_w2175_,
		_w2209_,
		_w3547_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		_w3078_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		_w2217_,
		_w3076_,
		_w3549_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		_w2217_,
		_w3076_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w3549_,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		_w3492_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h1)
	) name2373 (
		_w2200_,
		_w3076_,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		_w2200_,
		_w3076_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w3553_,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('h8)
	) name2376 (
		_w3552_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w2209_,
		_w3076_,
		_w3557_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		_w2209_,
		_w3076_,
		_w3558_
	);
	LUT2 #(
		.INIT('h1)
	) name2379 (
		_w3557_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		_w3556_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h4)
	) name2381 (
		_w3548_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h1)
	) name2382 (
		_w2150_,
		_w3076_,
		_w3562_
	);
	LUT2 #(
		.INIT('h8)
	) name2383 (
		_w2150_,
		_w3076_,
		_w3563_
	);
	LUT2 #(
		.INIT('h1)
	) name2384 (
		_w3562_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		_w3561_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		_w2159_,
		_w3076_,
		_w3566_
	);
	LUT2 #(
		.INIT('h8)
	) name2387 (
		_w2159_,
		_w3076_,
		_w3567_
	);
	LUT2 #(
		.INIT('h1)
	) name2388 (
		_w3566_,
		_w3567_,
		_w3568_
	);
	LUT2 #(
		.INIT('h8)
	) name2389 (
		_w3565_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h1)
	) name2390 (
		_w2142_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		_w2142_,
		_w3569_,
		_w3571_
	);
	LUT2 #(
		.INIT('h1)
	) name2392 (
		_w3570_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		_w3099_,
		_w3572_,
		_w3573_
	);
	LUT2 #(
		.INIT('h1)
	) name2394 (
		_w3096_,
		_w3546_,
		_w3574_
	);
	LUT2 #(
		.INIT('h4)
	) name2395 (
		_w3573_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		\g7961_pad ,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h1)
	) name2397 (
		\g267_reg/NET0131 ,
		\g7961_pad ,
		_w3577_
	);
	LUT2 #(
		.INIT('h1)
	) name2398 (
		_w3576_,
		_w3577_,
		_w3578_
	);
	LUT2 #(
		.INIT('h2)
	) name2399 (
		\g1092_reg/NET0131 ,
		_w3575_,
		_w3579_
	);
	LUT2 #(
		.INIT('h1)
	) name2400 (
		\g1092_reg/NET0131 ,
		\g270_reg/NET0131 ,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w3579_,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h2)
	) name2402 (
		\g1088_reg/NET0131 ,
		_w3575_,
		_w3582_
	);
	LUT2 #(
		.INIT('h1)
	) name2403 (
		\g1088_reg/NET0131 ,
		\g273_reg/NET0131 ,
		_w3583_
	);
	LUT2 #(
		.INIT('h1)
	) name2404 (
		_w3582_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h4)
	) name2405 (
		_w1832_,
		_w1901_,
		_w3585_
	);
	LUT2 #(
		.INIT('h1)
	) name2406 (
		\g1916_reg/NET0131 ,
		_w3024_,
		_w3586_
	);
	LUT2 #(
		.INIT('h8)
	) name2407 (
		_w1739_,
		_w3586_,
		_w3587_
	);
	LUT2 #(
		.INIT('h4)
	) name2408 (
		_w1837_,
		_w1866_,
		_w3588_
	);
	LUT2 #(
		.INIT('h1)
	) name2409 (
		_w3022_,
		_w3587_,
		_w3589_
	);
	LUT2 #(
		.INIT('h4)
	) name2410 (
		_w3588_,
		_w3589_,
		_w3590_
	);
	LUT2 #(
		.INIT('h1)
	) name2411 (
		_w3585_,
		_w3590_,
		_w3591_
	);
	LUT2 #(
		.INIT('h4)
	) name2412 (
		_w1821_,
		_w1901_,
		_w3592_
	);
	LUT2 #(
		.INIT('h4)
	) name2413 (
		_w1837_,
		_w1858_,
		_w3593_
	);
	LUT2 #(
		.INIT('h1)
	) name2414 (
		\g1917_reg/NET0131 ,
		_w3024_,
		_w3594_
	);
	LUT2 #(
		.INIT('h8)
	) name2415 (
		_w1739_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h1)
	) name2416 (
		_w3022_,
		_w3595_,
		_w3596_
	);
	LUT2 #(
		.INIT('h4)
	) name2417 (
		_w3593_,
		_w3596_,
		_w3597_
	);
	LUT2 #(
		.INIT('h1)
	) name2418 (
		_w3592_,
		_w3597_,
		_w3598_
	);
	LUT2 #(
		.INIT('h2)
	) name2419 (
		_w2356_,
		_w3149_,
		_w3599_
	);
	LUT2 #(
		.INIT('h1)
	) name2420 (
		_w2482_,
		_w3230_,
		_w3600_
	);
	LUT2 #(
		.INIT('h8)
	) name2421 (
		_w2482_,
		_w3230_,
		_w3601_
	);
	LUT2 #(
		.INIT('h1)
	) name2422 (
		_w3600_,
		_w3601_,
		_w3602_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		_w3154_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h1)
	) name2424 (
		_w3151_,
		_w3599_,
		_w3604_
	);
	LUT2 #(
		.INIT('h4)
	) name2425 (
		_w3603_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		\g1088_reg/NET0131 ,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		\g1088_reg/NET0131 ,
		\g915_reg/NET0131 ,
		_w3607_
	);
	LUT2 #(
		.INIT('h1)
	) name2428 (
		_w3606_,
		_w3607_,
		_w3608_
	);
	LUT2 #(
		.INIT('h2)
	) name2429 (
		\g7961_pad ,
		_w3605_,
		_w3609_
	);
	LUT2 #(
		.INIT('h1)
	) name2430 (
		\g7961_pad ,
		\g909_reg/NET0131 ,
		_w3610_
	);
	LUT2 #(
		.INIT('h1)
	) name2431 (
		_w3609_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h2)
	) name2432 (
		\g1092_reg/NET0131 ,
		_w3605_,
		_w3612_
	);
	LUT2 #(
		.INIT('h1)
	) name2433 (
		\g1092_reg/NET0131 ,
		\g912_reg/NET0131 ,
		_w3613_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w3612_,
		_w3613_,
		_w3614_
	);
	LUT2 #(
		.INIT('h2)
	) name2435 (
		_w2047_,
		_w3097_,
		_w3615_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		_w2159_,
		_w3565_,
		_w3616_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		_w2159_,
		_w3565_,
		_w3617_
	);
	LUT2 #(
		.INIT('h1)
	) name2438 (
		_w3616_,
		_w3617_,
		_w3618_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		_w3099_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		_w3096_,
		_w3615_,
		_w3620_
	);
	LUT2 #(
		.INIT('h4)
	) name2441 (
		_w3619_,
		_w3620_,
		_w3621_
	);
	LUT2 #(
		.INIT('h2)
	) name2442 (
		\g7961_pad ,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h1)
	) name2443 (
		\g222_reg/NET0131 ,
		\g7961_pad ,
		_w3623_
	);
	LUT2 #(
		.INIT('h1)
	) name2444 (
		_w3622_,
		_w3623_,
		_w3624_
	);
	LUT2 #(
		.INIT('h2)
	) name2445 (
		\g1092_reg/NET0131 ,
		_w3621_,
		_w3625_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		\g1092_reg/NET0131 ,
		\g225_reg/NET0131 ,
		_w3626_
	);
	LUT2 #(
		.INIT('h1)
	) name2447 (
		_w3625_,
		_w3626_,
		_w3627_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		\g1088_reg/NET0131 ,
		_w3621_,
		_w3628_
	);
	LUT2 #(
		.INIT('h1)
	) name2449 (
		\g1088_reg/NET0131 ,
		\g228_reg/NET0131 ,
		_w3629_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		_w3628_,
		_w3629_,
		_w3630_
	);
	LUT2 #(
		.INIT('h2)
	) name2451 (
		_w1223_,
		_w3331_,
		_w3631_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		_w1384_,
		_w3429_,
		_w3632_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		_w1384_,
		_w3429_,
		_w3633_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		_w3632_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h8)
	) name2455 (
		_w3336_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name2456 (
		_w3333_,
		_w3631_,
		_w3636_
	);
	LUT2 #(
		.INIT('h4)
	) name2457 (
		_w3635_,
		_w3636_,
		_w3637_
	);
	LUT2 #(
		.INIT('h2)
	) name2458 (
		\g7961_pad ,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h1)
	) name2459 (
		\g2297_reg/NET0131 ,
		\g7961_pad ,
		_w3639_
	);
	LUT2 #(
		.INIT('h1)
	) name2460 (
		_w3638_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h2)
	) name2461 (
		\g1092_reg/NET0131 ,
		_w3637_,
		_w3641_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		\g1092_reg/NET0131 ,
		\g2300_reg/NET0131 ,
		_w3642_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w3641_,
		_w3642_,
		_w3643_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		\g1088_reg/NET0131 ,
		_w3637_,
		_w3644_
	);
	LUT2 #(
		.INIT('h1)
	) name2465 (
		\g1088_reg/NET0131 ,
		\g2303_reg/NET0131 ,
		_w3645_
	);
	LUT2 #(
		.INIT('h1)
	) name2466 (
		_w3644_,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h2)
	) name2467 (
		_w2610_,
		_w3279_,
		_w3647_
	);
	LUT2 #(
		.INIT('h1)
	) name2468 (
		_w2615_,
		_w3529_,
		_w3648_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		_w2615_,
		_w3529_,
		_w3649_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		_w3648_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h8)
	) name2471 (
		_w3284_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h1)
	) name2472 (
		_w3281_,
		_w3647_,
		_w3652_
	);
	LUT2 #(
		.INIT('h4)
	) name2473 (
		_w3651_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h2)
	) name2474 (
		\g7961_pad ,
		_w3653_,
		_w3654_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		\g1603_reg/NET0131 ,
		\g7961_pad ,
		_w3655_
	);
	LUT2 #(
		.INIT('h1)
	) name2476 (
		_w3654_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h2)
	) name2477 (
		\g1092_reg/NET0131 ,
		_w3653_,
		_w3657_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		\g1092_reg/NET0131 ,
		\g1606_reg/NET0131 ,
		_w3658_
	);
	LUT2 #(
		.INIT('h1)
	) name2479 (
		_w3657_,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h2)
	) name2480 (
		\g1088_reg/NET0131 ,
		_w3653_,
		_w3660_
	);
	LUT2 #(
		.INIT('h1)
	) name2481 (
		\g1088_reg/NET0131 ,
		\g1609_reg/NET0131 ,
		_w3661_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		_w3660_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h4)
	) name2483 (
		\g499_reg/NET0131 ,
		\g548_reg/NET0131 ,
		_w3663_
	);
	LUT2 #(
		.INIT('h4)
	) name2484 (
		\g5657_pad ,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w1532_,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('h1)
	) name2486 (
		\g559_reg/NET0131 ,
		\g563_pad ,
		_w3666_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		_w3665_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		\g499_reg/NET0131 ,
		_w3667_,
		_w3668_
	);
	LUT2 #(
		.INIT('h8)
	) name2489 (
		\g5657_pad ,
		\g605_reg/NET0131 ,
		_w3669_
	);
	LUT2 #(
		.INIT('h8)
	) name2490 (
		\g1018_reg/NET0131 ,
		\g608_reg/NET0131 ,
		_w3670_
	);
	LUT2 #(
		.INIT('h8)
	) name2491 (
		\g1024_reg/NET0131 ,
		\g611_reg/NET0131 ,
		_w3671_
	);
	LUT2 #(
		.INIT('h1)
	) name2492 (
		_w3669_,
		_w3670_,
		_w3672_
	);
	LUT2 #(
		.INIT('h4)
	) name2493 (
		_w3671_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h2)
	) name2494 (
		\g1024_reg/NET0131 ,
		\g725_reg/NET0131 ,
		_w3674_
	);
	LUT2 #(
		.INIT('h2)
	) name2495 (
		\g1018_reg/NET0131 ,
		\g727_reg/NET0131 ,
		_w3675_
	);
	LUT2 #(
		.INIT('h2)
	) name2496 (
		\g5657_pad ,
		\g726_reg/NET0131 ,
		_w3676_
	);
	LUT2 #(
		.INIT('h1)
	) name2497 (
		_w3674_,
		_w3675_,
		_w3677_
	);
	LUT2 #(
		.INIT('h4)
	) name2498 (
		_w3676_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h2)
	) name2499 (
		\g5657_pad ,
		\g732_reg/NET0131 ,
		_w3679_
	);
	LUT2 #(
		.INIT('h2)
	) name2500 (
		\g1018_reg/NET0131 ,
		\g733_reg/NET0131 ,
		_w3680_
	);
	LUT2 #(
		.INIT('h2)
	) name2501 (
		\g1024_reg/NET0131 ,
		\g731_reg/NET0131 ,
		_w3681_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w3679_,
		_w3680_,
		_w3682_
	);
	LUT2 #(
		.INIT('h4)
	) name2503 (
		_w3681_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h2)
	) name2504 (
		\g1018_reg/NET0131 ,
		\g712_reg/NET0131 ,
		_w3684_
	);
	LUT2 #(
		.INIT('h2)
	) name2505 (
		\g1024_reg/NET0131 ,
		\g710_reg/NET0131 ,
		_w3685_
	);
	LUT2 #(
		.INIT('h2)
	) name2506 (
		\g5657_pad ,
		\g711_reg/NET0131 ,
		_w3686_
	);
	LUT2 #(
		.INIT('h1)
	) name2507 (
		_w3684_,
		_w3685_,
		_w3687_
	);
	LUT2 #(
		.INIT('h4)
	) name2508 (
		_w3686_,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h2)
	) name2509 (
		\g1024_reg/NET0131 ,
		\g716_reg/NET0131 ,
		_w3689_
	);
	LUT2 #(
		.INIT('h2)
	) name2510 (
		\g1018_reg/NET0131 ,
		\g718_reg/NET0131 ,
		_w3690_
	);
	LUT2 #(
		.INIT('h2)
	) name2511 (
		\g5657_pad ,
		\g717_reg/NET0131 ,
		_w3691_
	);
	LUT2 #(
		.INIT('h1)
	) name2512 (
		_w3689_,
		_w3690_,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name2513 (
		_w3691_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h2)
	) name2514 (
		\g1018_reg/NET0131 ,
		\g724_reg/NET0131 ,
		_w3694_
	);
	LUT2 #(
		.INIT('h2)
	) name2515 (
		\g1024_reg/NET0131 ,
		\g722_reg/NET0131 ,
		_w3695_
	);
	LUT2 #(
		.INIT('h2)
	) name2516 (
		\g5657_pad ,
		\g723_reg/NET0131 ,
		_w3696_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w3694_,
		_w3695_,
		_w3697_
	);
	LUT2 #(
		.INIT('h4)
	) name2518 (
		_w3696_,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h2)
	) name2519 (
		\g1024_reg/NET0131 ,
		\g701_reg/NET0131 ,
		_w3699_
	);
	LUT2 #(
		.INIT('h2)
	) name2520 (
		\g1018_reg/NET0131 ,
		\g703_reg/NET0131 ,
		_w3700_
	);
	LUT2 #(
		.INIT('h2)
	) name2521 (
		\g5657_pad ,
		\g702_reg/NET0131 ,
		_w3701_
	);
	LUT2 #(
		.INIT('h1)
	) name2522 (
		_w3699_,
		_w3700_,
		_w3702_
	);
	LUT2 #(
		.INIT('h4)
	) name2523 (
		_w3701_,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h2)
	) name2524 (
		\g1024_reg/NET0131 ,
		\g698_reg/NET0131 ,
		_w3704_
	);
	LUT2 #(
		.INIT('h2)
	) name2525 (
		\g1018_reg/NET0131 ,
		\g700_reg/NET0131 ,
		_w3705_
	);
	LUT2 #(
		.INIT('h2)
	) name2526 (
		\g5657_pad ,
		\g699_reg/NET0131 ,
		_w3706_
	);
	LUT2 #(
		.INIT('h1)
	) name2527 (
		_w3704_,
		_w3705_,
		_w3707_
	);
	LUT2 #(
		.INIT('h4)
	) name2528 (
		_w3706_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h2)
	) name2529 (
		\g1018_reg/NET0131 ,
		\g709_reg/NET0131 ,
		_w3709_
	);
	LUT2 #(
		.INIT('h2)
	) name2530 (
		\g1024_reg/NET0131 ,
		\g707_reg/NET0131 ,
		_w3710_
	);
	LUT2 #(
		.INIT('h2)
	) name2531 (
		\g5657_pad ,
		\g708_reg/NET0131 ,
		_w3711_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		_w3709_,
		_w3710_,
		_w3712_
	);
	LUT2 #(
		.INIT('h4)
	) name2533 (
		_w3711_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h2)
	) name2534 (
		\g1024_reg/NET0131 ,
		\g704_reg/NET0131 ,
		_w3714_
	);
	LUT2 #(
		.INIT('h2)
	) name2535 (
		\g1018_reg/NET0131 ,
		\g706_reg/NET0131 ,
		_w3715_
	);
	LUT2 #(
		.INIT('h2)
	) name2536 (
		\g5657_pad ,
		\g705_reg/NET0131 ,
		_w3716_
	);
	LUT2 #(
		.INIT('h1)
	) name2537 (
		_w3714_,
		_w3715_,
		_w3717_
	);
	LUT2 #(
		.INIT('h4)
	) name2538 (
		_w3716_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h2)
	) name2539 (
		\g1024_reg/NET0131 ,
		\g713_reg/NET0131 ,
		_w3719_
	);
	LUT2 #(
		.INIT('h2)
	) name2540 (
		\g1018_reg/NET0131 ,
		\g715_reg/NET0131 ,
		_w3720_
	);
	LUT2 #(
		.INIT('h2)
	) name2541 (
		\g5657_pad ,
		\g714_reg/NET0131 ,
		_w3721_
	);
	LUT2 #(
		.INIT('h1)
	) name2542 (
		_w3719_,
		_w3720_,
		_w3722_
	);
	LUT2 #(
		.INIT('h4)
	) name2543 (
		_w3721_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		\g1018_reg/NET0131 ,
		\g739_reg/NET0131 ,
		_w3724_
	);
	LUT2 #(
		.INIT('h2)
	) name2545 (
		\g1024_reg/NET0131 ,
		\g737_reg/NET0131 ,
		_w3725_
	);
	LUT2 #(
		.INIT('h2)
	) name2546 (
		\g5657_pad ,
		\g738_reg/NET0131 ,
		_w3726_
	);
	LUT2 #(
		.INIT('h1)
	) name2547 (
		_w3724_,
		_w3725_,
		_w3727_
	);
	LUT2 #(
		.INIT('h4)
	) name2548 (
		_w3726_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h2)
	) name2549 (
		\g1024_reg/NET0131 ,
		\g719_reg/NET0131 ,
		_w3729_
	);
	LUT2 #(
		.INIT('h2)
	) name2550 (
		\g1018_reg/NET0131 ,
		\g721_reg/NET0131 ,
		_w3730_
	);
	LUT2 #(
		.INIT('h2)
	) name2551 (
		\g5657_pad ,
		\g720_reg/NET0131 ,
		_w3731_
	);
	LUT2 #(
		.INIT('h1)
	) name2552 (
		_w3729_,
		_w3730_,
		_w3732_
	);
	LUT2 #(
		.INIT('h4)
	) name2553 (
		_w3731_,
		_w3732_,
		_w3733_
	);
	LUT2 #(
		.INIT('h1)
	) name2554 (
		_w3678_,
		_w3683_,
		_w3734_
	);
	LUT2 #(
		.INIT('h8)
	) name2555 (
		_w3688_,
		_w3693_,
		_w3735_
	);
	LUT2 #(
		.INIT('h1)
	) name2556 (
		_w3698_,
		_w3703_,
		_w3736_
	);
	LUT2 #(
		.INIT('h2)
	) name2557 (
		_w3708_,
		_w3713_,
		_w3737_
	);
	LUT2 #(
		.INIT('h4)
	) name2558 (
		_w3718_,
		_w3723_,
		_w3738_
	);
	LUT2 #(
		.INIT('h4)
	) name2559 (
		_w3728_,
		_w3733_,
		_w3739_
	);
	LUT2 #(
		.INIT('h8)
	) name2560 (
		_w3738_,
		_w3739_,
		_w3740_
	);
	LUT2 #(
		.INIT('h8)
	) name2561 (
		_w3736_,
		_w3737_,
		_w3741_
	);
	LUT2 #(
		.INIT('h8)
	) name2562 (
		_w3734_,
		_w3735_,
		_w3742_
	);
	LUT2 #(
		.INIT('h8)
	) name2563 (
		_w3741_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h8)
	) name2564 (
		_w3740_,
		_w3743_,
		_w3744_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w3678_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('h4)
	) name2566 (
		_w3673_,
		_w3745_,
		_w3746_
	);
	LUT2 #(
		.INIT('h2)
	) name2567 (
		_w3673_,
		_w3745_,
		_w3747_
	);
	LUT2 #(
		.INIT('h1)
	) name2568 (
		_w3746_,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h2)
	) name2569 (
		_w3668_,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h8)
	) name2570 (
		\g5657_pad ,
		\g614_reg/NET0131 ,
		_w3750_
	);
	LUT2 #(
		.INIT('h8)
	) name2571 (
		\g1024_reg/NET0131 ,
		\g620_reg/NET0131 ,
		_w3751_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		\g1018_reg/NET0131 ,
		\g617_reg/NET0131 ,
		_w3752_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		_w3750_,
		_w3751_,
		_w3753_
	);
	LUT2 #(
		.INIT('h4)
	) name2574 (
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT2 #(
		.INIT('h1)
	) name2575 (
		_w3698_,
		_w3744_,
		_w3755_
	);
	LUT2 #(
		.INIT('h4)
	) name2576 (
		_w3754_,
		_w3755_,
		_w3756_
	);
	LUT2 #(
		.INIT('h2)
	) name2577 (
		_w3754_,
		_w3755_,
		_w3757_
	);
	LUT2 #(
		.INIT('h1)
	) name2578 (
		_w3756_,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h8)
	) name2579 (
		_w3749_,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h2)
	) name2580 (
		_w3668_,
		_w3758_,
		_w3760_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		_w3748_,
		_w3760_,
		_w3761_
	);
	LUT2 #(
		.INIT('h1)
	) name2582 (
		_w3759_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		\g1243_reg/NET0131 ,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h2)
	) name2584 (
		\g3229_pad ,
		\g538_reg/NET0131 ,
		_w3764_
	);
	LUT2 #(
		.INIT('h4)
	) name2585 (
		\g499_reg/NET0131 ,
		\g5657_pad ,
		_w3765_
	);
	LUT2 #(
		.INIT('h2)
	) name2586 (
		_w3667_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h8)
	) name2587 (
		\g525_reg/NET0131 ,
		_w1550_,
		_w3767_
	);
	LUT2 #(
		.INIT('h1)
	) name2588 (
		\g3229_pad ,
		\g541_reg/NET0131 ,
		_w3768_
	);
	LUT2 #(
		.INIT('h1)
	) name2589 (
		_w3764_,
		_w3768_,
		_w3769_
	);
	LUT2 #(
		.INIT('h8)
	) name2590 (
		_w3767_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h8)
	) name2591 (
		_w3766_,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h2)
	) name2592 (
		_w3688_,
		_w3754_,
		_w3772_
	);
	LUT2 #(
		.INIT('h4)
	) name2593 (
		_w3688_,
		_w3754_,
		_w3773_
	);
	LUT2 #(
		.INIT('h1)
	) name2594 (
		_w3772_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h8)
	) name2595 (
		_w3668_,
		_w3774_,
		_w3775_
	);
	LUT2 #(
		.INIT('h2)
	) name2596 (
		_w3673_,
		_w3723_,
		_w3776_
	);
	LUT2 #(
		.INIT('h4)
	) name2597 (
		_w3673_,
		_w3723_,
		_w3777_
	);
	LUT2 #(
		.INIT('h1)
	) name2598 (
		_w3776_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h2)
	) name2599 (
		_w3775_,
		_w3778_,
		_w3779_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		_w3668_,
		_w3778_,
		_w3780_
	);
	LUT2 #(
		.INIT('h4)
	) name2601 (
		_w3774_,
		_w3780_,
		_w3781_
	);
	LUT2 #(
		.INIT('h1)
	) name2602 (
		_w3779_,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h2)
	) name2603 (
		_w3673_,
		_w3733_,
		_w3783_
	);
	LUT2 #(
		.INIT('h4)
	) name2604 (
		_w3673_,
		_w3733_,
		_w3784_
	);
	LUT2 #(
		.INIT('h1)
	) name2605 (
		_w3783_,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('h8)
	) name2606 (
		_w3668_,
		_w3785_,
		_w3786_
	);
	LUT2 #(
		.INIT('h2)
	) name2607 (
		_w3693_,
		_w3754_,
		_w3787_
	);
	LUT2 #(
		.INIT('h4)
	) name2608 (
		_w3693_,
		_w3754_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name2609 (
		_w3787_,
		_w3788_,
		_w3789_
	);
	LUT2 #(
		.INIT('h2)
	) name2610 (
		_w3786_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		_w3668_,
		_w3789_,
		_w3791_
	);
	LUT2 #(
		.INIT('h4)
	) name2612 (
		_w3785_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h1)
	) name2613 (
		_w3790_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h2)
	) name2614 (
		_w3708_,
		_w3754_,
		_w3794_
	);
	LUT2 #(
		.INIT('h4)
	) name2615 (
		_w3708_,
		_w3754_,
		_w3795_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w3794_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h8)
	) name2617 (
		_w3668_,
		_w3796_,
		_w3797_
	);
	LUT2 #(
		.INIT('h1)
	) name2618 (
		_w3703_,
		_w3744_,
		_w3798_
	);
	LUT2 #(
		.INIT('h4)
	) name2619 (
		_w3673_,
		_w3798_,
		_w3799_
	);
	LUT2 #(
		.INIT('h2)
	) name2620 (
		_w3673_,
		_w3798_,
		_w3800_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		_w3799_,
		_w3800_,
		_w3801_
	);
	LUT2 #(
		.INIT('h8)
	) name2622 (
		_w3797_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h2)
	) name2623 (
		_w3668_,
		_w3801_,
		_w3803_
	);
	LUT2 #(
		.INIT('h4)
	) name2624 (
		_w3796_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		_w3802_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w3713_,
		_w3744_,
		_w3806_
	);
	LUT2 #(
		.INIT('h4)
	) name2627 (
		_w3673_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h2)
	) name2628 (
		_w3673_,
		_w3806_,
		_w3808_
	);
	LUT2 #(
		.INIT('h1)
	) name2629 (
		_w3807_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h2)
	) name2630 (
		_w3668_,
		_w3809_,
		_w3810_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w3718_,
		_w3744_,
		_w3811_
	);
	LUT2 #(
		.INIT('h4)
	) name2632 (
		_w3754_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h2)
	) name2633 (
		_w3754_,
		_w3811_,
		_w3813_
	);
	LUT2 #(
		.INIT('h1)
	) name2634 (
		_w3812_,
		_w3813_,
		_w3814_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		_w3810_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('h2)
	) name2636 (
		_w3668_,
		_w3814_,
		_w3816_
	);
	LUT2 #(
		.INIT('h8)
	) name2637 (
		_w3809_,
		_w3816_,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w3815_,
		_w3817_,
		_w3818_
	);
	LUT2 #(
		.INIT('h2)
	) name2639 (
		_w3805_,
		_w3818_,
		_w3819_
	);
	LUT2 #(
		.INIT('h4)
	) name2640 (
		_w3805_,
		_w3818_,
		_w3820_
	);
	LUT2 #(
		.INIT('h1)
	) name2641 (
		_w3819_,
		_w3820_,
		_w3821_
	);
	LUT2 #(
		.INIT('h8)
	) name2642 (
		_w3793_,
		_w3821_,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name2643 (
		_w3793_,
		_w3821_,
		_w3823_
	);
	LUT2 #(
		.INIT('h1)
	) name2644 (
		_w3822_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h2)
	) name2645 (
		_w3782_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h4)
	) name2646 (
		_w3782_,
		_w3824_,
		_w3826_
	);
	LUT2 #(
		.INIT('h2)
	) name2647 (
		\g1196_reg/NET0131 ,
		_w3825_,
		_w3827_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		_w3826_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w3763_,
		_w3771_,
		_w3829_
	);
	LUT2 #(
		.INIT('h4)
	) name2650 (
		_w3828_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		_w2014_,
		_w3064_,
		_w3831_
	);
	LUT2 #(
		.INIT('h2)
	) name2652 (
		\g1563_reg/NET0131 ,
		_w3831_,
		_w3832_
	);
	LUT2 #(
		.INIT('h2)
	) name2653 (
		_w2024_,
		_w3832_,
		_w3833_
	);
	LUT2 #(
		.INIT('h4)
	) name2654 (
		_w2024_,
		_w3064_,
		_w3834_
	);
	LUT2 #(
		.INIT('h2)
	) name2655 (
		_w2117_,
		_w2226_,
		_w3835_
	);
	LUT2 #(
		.INIT('h1)
	) name2656 (
		_w3834_,
		_w3835_,
		_w3836_
	);
	LUT2 #(
		.INIT('h1)
	) name2657 (
		_w2014_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w3833_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w2019_,
		_w2265_,
		_w3839_
	);
	LUT2 #(
		.INIT('h4)
	) name2660 (
		_w3838_,
		_w3839_,
		_w3840_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		_w1309_,
		_w3323_,
		_w3841_
	);
	LUT2 #(
		.INIT('h2)
	) name2662 (
		\g1563_reg/NET0131 ,
		_w3841_,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name2663 (
		_w1298_,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name2664 (
		_w1418_,
		_w1442_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name2665 (
		_w3843_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('h1)
	) name2666 (
		_w1293_,
		_w1303_,
		_w3846_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		_w3845_,
		_w3846_,
		_w3847_
	);
	LUT2 #(
		.INIT('h2)
	) name2668 (
		_w2413_,
		_w3144_,
		_w3848_
	);
	LUT2 #(
		.INIT('h2)
	) name2669 (
		\g1563_reg/NET0131 ,
		_w3848_,
		_w3849_
	);
	LUT2 #(
		.INIT('h2)
	) name2670 (
		_w2288_,
		_w3849_,
		_w3850_
	);
	LUT2 #(
		.INIT('h4)
	) name2671 (
		_w2413_,
		_w2544_,
		_w3851_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		_w3850_,
		_w3851_,
		_w3852_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		_w2408_,
		_w2543_,
		_w3853_
	);
	LUT2 #(
		.INIT('h4)
	) name2674 (
		_w3852_,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h2)
	) name2675 (
		_w2720_,
		_w3272_,
		_w3855_
	);
	LUT2 #(
		.INIT('h2)
	) name2676 (
		\g1563_reg/NET0131 ,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		_w2699_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h2)
	) name2678 (
		_w2694_,
		_w2720_,
		_w3858_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w3857_,
		_w3858_,
		_w3859_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w2574_,
		_w2835_,
		_w3860_
	);
	LUT2 #(
		.INIT('h4)
	) name2681 (
		_w3859_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h8)
	) name2682 (
		\g2580_reg/NET0131 ,
		\g2581_reg/NET0131 ,
		_w3862_
	);
	LUT2 #(
		.INIT('h1)
	) name2683 (
		\g1018_reg/NET0131 ,
		\g16437_pad ,
		_w3863_
	);
	LUT2 #(
		.INIT('h8)
	) name2684 (
		\g1886_reg/NET0131 ,
		\g1887_reg/NET0131 ,
		_w3864_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		\g1018_reg/NET0131 ,
		\g16399_pad ,
		_w3865_
	);
	LUT2 #(
		.INIT('h2)
	) name2686 (
		\g1192_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		_w3866_
	);
	LUT2 #(
		.INIT('h4)
	) name2687 (
		\g1018_reg/NET0131 ,
		\g16355_pad ,
		_w3867_
	);
	LUT2 #(
		.INIT('h2)
	) name2688 (
		\g506_reg/NET0131 ,
		\g507_reg/NET0131 ,
		_w3868_
	);
	LUT2 #(
		.INIT('h2)
	) name2689 (
		\g1018_reg/NET0131 ,
		_w3868_,
		_w3869_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		\g1192_reg/NET0131 ,
		_w3867_,
		_w3870_
	);
	LUT2 #(
		.INIT('h4)
	) name2691 (
		_w3869_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h1)
	) name2692 (
		_w3866_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h2)
	) name2693 (
		\g1018_reg/NET0131 ,
		_w3872_,
		_w3873_
	);
	LUT2 #(
		.INIT('h1)
	) name2694 (
		\g1886_reg/NET0131 ,
		_w3865_,
		_w3874_
	);
	LUT2 #(
		.INIT('h4)
	) name2695 (
		_w3873_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h1)
	) name2696 (
		_w3864_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h8)
	) name2697 (
		\g1018_reg/NET0131 ,
		_w3876_,
		_w3877_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		\g2580_reg/NET0131 ,
		_w3863_,
		_w3878_
	);
	LUT2 #(
		.INIT('h4)
	) name2699 (
		_w3877_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h1)
	) name2700 (
		_w3862_,
		_w3879_,
		_w3880_
	);
	LUT2 #(
		.INIT('h2)
	) name2701 (
		\g805_reg/NET0131 ,
		_w3149_,
		_w3881_
	);
	LUT2 #(
		.INIT('h2)
	) name2702 (
		_w2436_,
		_w3223_,
		_w3882_
	);
	LUT2 #(
		.INIT('h4)
	) name2703 (
		_w2436_,
		_w3223_,
		_w3883_
	);
	LUT2 #(
		.INIT('h1)
	) name2704 (
		_w3882_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h8)
	) name2705 (
		_w3154_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w3881_,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w2209_,
		_w3556_,
		_w3887_
	);
	LUT2 #(
		.INIT('h8)
	) name2708 (
		_w2209_,
		_w3556_,
		_w3888_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w3887_,
		_w3888_,
		_w3889_
	);
	LUT2 #(
		.INIT('h8)
	) name2710 (
		_w3099_,
		_w3889_,
		_w3890_
	);
	LUT2 #(
		.INIT('h1)
	) name2711 (
		\g117_reg/NET0131 ,
		_w3075_,
		_w3891_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		_w3095_,
		_w3891_,
		_w3892_
	);
	LUT2 #(
		.INIT('h4)
	) name2713 (
		_w3890_,
		_w3892_,
		_w3893_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		\g1421_reg/NET0131 ,
		\g5657_pad ,
		_w3894_
	);
	LUT2 #(
		.INIT('h2)
	) name2715 (
		\g1024_reg/NET0131 ,
		\g1420_reg/NET0131 ,
		_w3895_
	);
	LUT2 #(
		.INIT('h2)
	) name2716 (
		\g1018_reg/NET0131 ,
		\g1422_reg/NET0131 ,
		_w3896_
	);
	LUT2 #(
		.INIT('h1)
	) name2717 (
		_w3894_,
		_w3895_,
		_w3897_
	);
	LUT2 #(
		.INIT('h4)
	) name2718 (
		_w3896_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		_w2923_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h2)
	) name2720 (
		_w2852_,
		_w3899_,
		_w3900_
	);
	LUT2 #(
		.INIT('h2)
	) name2721 (
		_w1901_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w1911_,
		_w2949_,
		_w3902_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w1901_,
		_w2949_,
		_w3903_
	);
	LUT2 #(
		.INIT('h8)
	) name2724 (
		_w2994_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		\g1215_reg/NET0131 ,
		_w3903_,
		_w3905_
	);
	LUT2 #(
		.INIT('h8)
	) name2726 (
		_w2851_,
		_w3905_,
		_w3906_
	);
	LUT2 #(
		.INIT('h1)
	) name2727 (
		_w3902_,
		_w3906_,
		_w3907_
	);
	LUT2 #(
		.INIT('h4)
	) name2728 (
		_w3904_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w3901_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('h2)
	) name2730 (
		\g1186_reg/NET0131 ,
		_w3899_,
		_w3910_
	);
	LUT2 #(
		.INIT('h2)
	) name2731 (
		_w2851_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h2)
	) name2732 (
		_w1901_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		\g1217_reg/NET0131 ,
		_w3903_,
		_w3913_
	);
	LUT2 #(
		.INIT('h8)
	) name2734 (
		_w2851_,
		_w3913_,
		_w3914_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		_w2949_,
		_w2985_,
		_w3915_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w3902_,
		_w3914_,
		_w3916_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w3915_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h1)
	) name2738 (
		_w3912_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		\g1218_reg/NET0131 ,
		_w3903_,
		_w3919_
	);
	LUT2 #(
		.INIT('h8)
	) name2740 (
		_w2851_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('h4)
	) name2741 (
		_w2949_,
		_w3000_,
		_w3921_
	);
	LUT2 #(
		.INIT('h1)
	) name2742 (
		_w3902_,
		_w3920_,
		_w3922_
	);
	LUT2 #(
		.INIT('h4)
	) name2743 (
		_w3921_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h1)
	) name2744 (
		_w3901_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h2)
	) name2745 (
		_w1901_,
		_w2851_,
		_w3925_
	);
	LUT2 #(
		.INIT('h8)
	) name2746 (
		_w2968_,
		_w3903_,
		_w3926_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		\g1219_reg/NET0131 ,
		_w3903_,
		_w3927_
	);
	LUT2 #(
		.INIT('h8)
	) name2748 (
		_w2851_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w3902_,
		_w3928_,
		_w3929_
	);
	LUT2 #(
		.INIT('h4)
	) name2750 (
		_w3926_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w3925_,
		_w3930_,
		_w3931_
	);
	LUT2 #(
		.INIT('h8)
	) name2752 (
		_w2962_,
		_w3903_,
		_w3932_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		\g1220_reg/NET0131 ,
		_w3903_,
		_w3933_
	);
	LUT2 #(
		.INIT('h8)
	) name2754 (
		_w2851_,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h1)
	) name2755 (
		_w3902_,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('h4)
	) name2756 (
		_w3932_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w3925_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h8)
	) name2758 (
		_w2989_,
		_w3903_,
		_w3938_
	);
	LUT2 #(
		.INIT('h1)
	) name2759 (
		\g1216_reg/NET0131 ,
		_w3903_,
		_w3939_
	);
	LUT2 #(
		.INIT('h8)
	) name2760 (
		_w2851_,
		_w3939_,
		_w3940_
	);
	LUT2 #(
		.INIT('h1)
	) name2761 (
		_w3902_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h4)
	) name2762 (
		_w3938_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w3912_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h2)
	) name2764 (
		\g1496_reg/NET0131 ,
		_w3279_,
		_w3944_
	);
	LUT2 #(
		.INIT('h2)
	) name2765 (
		_w2653_,
		_w3522_,
		_w3945_
	);
	LUT2 #(
		.INIT('h4)
	) name2766 (
		_w2653_,
		_w3522_,
		_w3946_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		_w3945_,
		_w3946_,
		_w3947_
	);
	LUT2 #(
		.INIT('h8)
	) name2768 (
		_w3284_,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		_w3944_,
		_w3948_,
		_w3949_
	);
	LUT2 #(
		.INIT('h1)
	) name2770 (
		_w2167_,
		_w2266_,
		_w3950_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		_w2167_,
		_w2266_,
		_w3951_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w3950_,
		_w3951_,
		_w3952_
	);
	LUT2 #(
		.INIT('h8)
	) name2773 (
		_w3099_,
		_w3952_,
		_w3953_
	);
	LUT2 #(
		.INIT('h1)
	) name2774 (
		\g97_reg/NET0131 ,
		_w3075_,
		_w3954_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		_w3095_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h4)
	) name2776 (
		_w3953_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name2777 (
		_w2200_,
		_w3552_,
		_w3957_
	);
	LUT2 #(
		.INIT('h8)
	) name2778 (
		_w2200_,
		_w3552_,
		_w3958_
	);
	LUT2 #(
		.INIT('h1)
	) name2779 (
		_w3957_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		_w3099_,
		_w3959_,
		_w3960_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		\g113_reg/NET0131 ,
		_w3075_,
		_w3961_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		_w3095_,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('h4)
	) name2783 (
		_w3960_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h2)
	) name2784 (
		\g785_reg/NET0131 ,
		_w3149_,
		_w3964_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w2510_,
		_w2550_,
		_w3965_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w3176_,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h2)
	) name2787 (
		_w3154_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w3964_,
		_w3967_,
		_w3968_
	);
	LUT2 #(
		.INIT('h2)
	) name2789 (
		\g1471_reg/NET0131 ,
		_w3279_,
		_w3969_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		_w2624_,
		_w2836_,
		_w3970_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w3455_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('h2)
	) name2792 (
		_w3284_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h1)
	) name2793 (
		_w3969_,
		_w3972_,
		_w3973_
	);
	LUT2 #(
		.INIT('h2)
	) name2794 (
		\g801_reg/NET0131 ,
		_w3149_,
		_w3974_
	);
	LUT2 #(
		.INIT('h2)
	) name2795 (
		_w2491_,
		_w3219_,
		_w3975_
	);
	LUT2 #(
		.INIT('h4)
	) name2796 (
		_w2491_,
		_w3219_,
		_w3976_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w3975_,
		_w3976_,
		_w3977_
	);
	LUT2 #(
		.INIT('h8)
	) name2798 (
		_w3154_,
		_w3977_,
		_w3978_
	);
	LUT2 #(
		.INIT('h1)
	) name2799 (
		_w3974_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h2)
	) name2800 (
		\g2165_reg/NET0131 ,
		_w3331_,
		_w3980_
	);
	LUT2 #(
		.INIT('h4)
	) name2801 (
		_w1304_,
		_w1409_,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name2802 (
		_w3361_,
		_w3981_,
		_w3982_
	);
	LUT2 #(
		.INIT('h8)
	) name2803 (
		_w3336_,
		_w3982_,
		_w3983_
	);
	LUT2 #(
		.INIT('h1)
	) name2804 (
		_w3980_,
		_w3983_,
		_w3984_
	);
	LUT2 #(
		.INIT('h2)
	) name2805 (
		\g2185_reg/NET0131 ,
		_w3331_,
		_w3985_
	);
	LUT2 #(
		.INIT('h1)
	) name2806 (
		_w3336_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h1)
	) name2807 (
		_w3415_,
		_w3417_,
		_w3987_
	);
	LUT2 #(
		.INIT('h2)
	) name2808 (
		_w3386_,
		_w3987_,
		_w3988_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w1376_,
		_w3988_,
		_w3989_
	);
	LUT2 #(
		.INIT('h8)
	) name2810 (
		_w1376_,
		_w3988_,
		_w3990_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w3989_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h8)
	) name2812 (
		_w3336_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h1)
	) name2813 (
		_w3986_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h2)
	) name2814 (
		\g2195_reg/NET0131 ,
		_w3331_,
		_w3994_
	);
	LUT2 #(
		.INIT('h2)
	) name2815 (
		_w1392_,
		_w3424_,
		_w3995_
	);
	LUT2 #(
		.INIT('h4)
	) name2816 (
		_w1392_,
		_w3424_,
		_w3996_
	);
	LUT2 #(
		.INIT('h1)
	) name2817 (
		_w3995_,
		_w3996_,
		_w3997_
	);
	LUT2 #(
		.INIT('h8)
	) name2818 (
		_w3336_,
		_w3997_,
		_w3998_
	);
	LUT2 #(
		.INIT('h1)
	) name2819 (
		_w3994_,
		_w3998_,
		_w3999_
	);
	LUT2 #(
		.INIT('h2)
	) name2820 (
		\g1491_reg/NET0131 ,
		_w3279_,
		_w4000_
	);
	LUT2 #(
		.INIT('h2)
	) name2821 (
		_w2585_,
		_w3518_,
		_w4001_
	);
	LUT2 #(
		.INIT('h4)
	) name2822 (
		_w2585_,
		_w3518_,
		_w4002_
	);
	LUT2 #(
		.INIT('h1)
	) name2823 (
		_w4001_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		_w3284_,
		_w4003_,
		_w4004_
	);
	LUT2 #(
		.INIT('h1)
	) name2825 (
		_w4000_,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		\g1501_reg/NET0131 ,
		_w3279_,
		_w4006_
	);
	LUT2 #(
		.INIT('h1)
	) name2827 (
		_w2653_,
		_w3260_,
		_w4007_
	);
	LUT2 #(
		.INIT('h2)
	) name2828 (
		_w3524_,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h2)
	) name2829 (
		_w2602_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h4)
	) name2830 (
		_w2602_,
		_w4008_,
		_w4010_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		_w4009_,
		_w4010_,
		_w4011_
	);
	LUT2 #(
		.INIT('h8)
	) name2832 (
		_w3284_,
		_w4011_,
		_w4012_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w4006_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h2)
	) name2834 (
		\g809_reg/NET0131 ,
		_w3149_,
		_w4014_
	);
	LUT2 #(
		.INIT('h1)
	) name2835 (
		_w3154_,
		_w4014_,
		_w4015_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		_w2436_,
		_w3132_,
		_w4016_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		_w3225_,
		_w4016_,
		_w4017_
	);
	LUT2 #(
		.INIT('h1)
	) name2838 (
		_w2500_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('h8)
	) name2839 (
		_w2500_,
		_w4017_,
		_w4019_
	);
	LUT2 #(
		.INIT('h1)
	) name2840 (
		_w4018_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h8)
	) name2841 (
		_w3154_,
		_w4020_,
		_w4021_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w4015_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h2)
	) name2843 (
		\g2200_reg/NET0131 ,
		_w3331_,
		_w4023_
	);
	LUT2 #(
		.INIT('h2)
	) name2844 (
		_w1338_,
		_w3428_,
		_w4024_
	);
	LUT2 #(
		.INIT('h4)
	) name2845 (
		_w1338_,
		_w3428_,
		_w4025_
	);
	LUT2 #(
		.INIT('h1)
	) name2846 (
		_w4024_,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h8)
	) name2847 (
		_w3336_,
		_w4026_,
		_w4027_
	);
	LUT2 #(
		.INIT('h1)
	) name2848 (
		_w4023_,
		_w4027_,
		_w4028_
	);
	LUT2 #(
		.INIT('h2)
	) name2849 (
		\g1506_reg/NET0131 ,
		_w3279_,
		_w4029_
	);
	LUT2 #(
		.INIT('h2)
	) name2850 (
		_w2662_,
		_w3525_,
		_w4030_
	);
	LUT2 #(
		.INIT('h4)
	) name2851 (
		_w2662_,
		_w3525_,
		_w4031_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w4030_,
		_w4031_,
		_w4032_
	);
	LUT2 #(
		.INIT('h8)
	) name2853 (
		_w3284_,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('h1)
	) name2854 (
		_w4029_,
		_w4033_,
		_w4034_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		\g813_reg/NET0131 ,
		_w3149_,
		_w4035_
	);
	LUT2 #(
		.INIT('h2)
	) name2856 (
		_w2444_,
		_w3226_,
		_w4036_
	);
	LUT2 #(
		.INIT('h4)
	) name2857 (
		_w2444_,
		_w3226_,
		_w4037_
	);
	LUT2 #(
		.INIT('h1)
	) name2858 (
		_w4036_,
		_w4037_,
		_w4038_
	);
	LUT2 #(
		.INIT('h8)
	) name2859 (
		_w3154_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w4035_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h2)
	) name2861 (
		\g125_reg/NET0131 ,
		_w3075_,
		_w4041_
	);
	LUT2 #(
		.INIT('h2)
	) name2862 (
		_w2150_,
		_w3561_,
		_w4042_
	);
	LUT2 #(
		.INIT('h4)
	) name2863 (
		_w2150_,
		_w3561_,
		_w4043_
	);
	LUT2 #(
		.INIT('h1)
	) name2864 (
		_w4042_,
		_w4043_,
		_w4044_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		_w3099_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		_w4041_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h2)
	) name2867 (
		_w1901_,
		_w2944_,
		_w4047_
	);
	LUT2 #(
		.INIT('h4)
	) name2868 (
		_w2949_,
		_w2975_,
		_w4048_
	);
	LUT2 #(
		.INIT('h1)
	) name2869 (
		\g1222_reg/NET0131 ,
		_w3903_,
		_w4049_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		_w2851_,
		_w4049_,
		_w4050_
	);
	LUT2 #(
		.INIT('h1)
	) name2871 (
		_w3902_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h4)
	) name2872 (
		_w4048_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h1)
	) name2873 (
		_w4047_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name2874 (
		_w1901_,
		_w2933_,
		_w4054_
	);
	LUT2 #(
		.INIT('h4)
	) name2875 (
		_w2949_,
		_w2957_,
		_w4055_
	);
	LUT2 #(
		.INIT('h1)
	) name2876 (
		\g1223_reg/NET0131 ,
		_w3903_,
		_w4056_
	);
	LUT2 #(
		.INIT('h8)
	) name2877 (
		_w2851_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h1)
	) name2878 (
		_w3902_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h4)
	) name2879 (
		_w4055_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h1)
	) name2880 (
		_w4054_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h1)
	) name2881 (
		_w2019_,
		_w3070_,
		_w4061_
	);
	LUT2 #(
		.INIT('h8)
	) name2882 (
		_w3064_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h1)
	) name2883 (
		_w3076_,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h1)
	) name2884 (
		_w2265_,
		_w4063_,
		_w4064_
	);
	LUT2 #(
		.INIT('h1)
	) name2885 (
		_w2408_,
		_w3140_,
		_w4065_
	);
	LUT2 #(
		.INIT('h4)
	) name2886 (
		_w3144_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w3132_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h1)
	) name2888 (
		_w2543_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h1)
	) name2889 (
		_w1303_,
		_w3319_,
		_w4069_
	);
	LUT2 #(
		.INIT('h8)
	) name2890 (
		_w3323_,
		_w4069_,
		_w4070_
	);
	LUT2 #(
		.INIT('h1)
	) name2891 (
		_w3309_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h1)
	) name2892 (
		_w1293_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h1)
	) name2893 (
		_w2574_,
		_w3268_,
		_w4073_
	);
	LUT2 #(
		.INIT('h4)
	) name2894 (
		_w3272_,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h1)
	) name2895 (
		_w3260_,
		_w4074_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name2896 (
		_w2835_,
		_w4075_,
		_w4076_
	);
	LUT2 #(
		.INIT('h2)
	) name2897 (
		\g1018_reg/NET0131 ,
		\g736_reg/NET0131 ,
		_w4077_
	);
	LUT2 #(
		.INIT('h2)
	) name2898 (
		\g1024_reg/NET0131 ,
		\g734_reg/NET0131 ,
		_w4078_
	);
	LUT2 #(
		.INIT('h2)
	) name2899 (
		\g5657_pad ,
		\g735_reg/NET0131 ,
		_w4079_
	);
	LUT2 #(
		.INIT('h1)
	) name2900 (
		_w4077_,
		_w4078_,
		_w4080_
	);
	LUT2 #(
		.INIT('h4)
	) name2901 (
		_w4079_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h4)
	) name2902 (
		_w3744_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h2)
	) name2903 (
		\g499_reg/NET0131 ,
		_w4082_,
		_w4083_
	);
	LUT2 #(
		.INIT('h2)
	) name2904 (
		_w3766_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h2)
	) name2905 (
		_w1901_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name2906 (
		_w1911_,
		_w3767_,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name2907 (
		_w1901_,
		_w3767_,
		_w4087_
	);
	LUT2 #(
		.INIT('h8)
	) name2908 (
		_w3791_,
		_w4087_,
		_w4088_
	);
	LUT2 #(
		.INIT('h1)
	) name2909 (
		\g530_reg/NET0131 ,
		_w4087_,
		_w4089_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		_w3766_,
		_w4089_,
		_w4090_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w4086_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h4)
	) name2912 (
		_w4088_,
		_w4091_,
		_w4092_
	);
	LUT2 #(
		.INIT('h1)
	) name2913 (
		_w4085_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h8)
	) name2914 (
		_w3780_,
		_w4087_,
		_w4094_
	);
	LUT2 #(
		.INIT('h1)
	) name2915 (
		\g531_reg/NET0131 ,
		_w4087_,
		_w4095_
	);
	LUT2 #(
		.INIT('h8)
	) name2916 (
		_w3766_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name2917 (
		_w4086_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h4)
	) name2918 (
		_w4094_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w4085_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h8)
	) name2920 (
		_w3667_,
		_w4083_,
		_w4100_
	);
	LUT2 #(
		.INIT('h2)
	) name2921 (
		_w1901_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h8)
	) name2922 (
		_w3786_,
		_w4087_,
		_w4102_
	);
	LUT2 #(
		.INIT('h1)
	) name2923 (
		\g529_reg/NET0131 ,
		_w4087_,
		_w4103_
	);
	LUT2 #(
		.INIT('h8)
	) name2924 (
		_w3766_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h1)
	) name2925 (
		_w4086_,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('h4)
	) name2926 (
		_w4102_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h1)
	) name2927 (
		_w4101_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h8)
	) name2928 (
		_w3775_,
		_w4087_,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name2929 (
		\g532_reg/NET0131 ,
		_w4087_,
		_w4109_
	);
	LUT2 #(
		.INIT('h8)
	) name2930 (
		_w3766_,
		_w4109_,
		_w4110_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		_w4086_,
		_w4110_,
		_w4111_
	);
	LUT2 #(
		.INIT('h4)
	) name2932 (
		_w4108_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h1)
	) name2933 (
		_w4101_,
		_w4112_,
		_w4113_
	);
	LUT2 #(
		.INIT('h2)
	) name2934 (
		_w1901_,
		_w3766_,
		_w4114_
	);
	LUT2 #(
		.INIT('h8)
	) name2935 (
		_w3810_,
		_w4087_,
		_w4115_
	);
	LUT2 #(
		.INIT('h1)
	) name2936 (
		\g533_reg/NET0131 ,
		_w4087_,
		_w4116_
	);
	LUT2 #(
		.INIT('h8)
	) name2937 (
		_w3766_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h1)
	) name2938 (
		_w4086_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('h4)
	) name2939 (
		_w4115_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h1)
	) name2940 (
		_w4114_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		_w3816_,
		_w4087_,
		_w4121_
	);
	LUT2 #(
		.INIT('h1)
	) name2942 (
		\g534_reg/NET0131 ,
		_w4087_,
		_w4122_
	);
	LUT2 #(
		.INIT('h8)
	) name2943 (
		_w3766_,
		_w4122_,
		_w4123_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		_w4086_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h4)
	) name2945 (
		_w4121_,
		_w4124_,
		_w4125_
	);
	LUT2 #(
		.INIT('h1)
	) name2946 (
		_w4114_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h4)
	) name2947 (
		\g2993_reg/NET0131 ,
		\g2998_reg/NET0131 ,
		_w4127_
	);
	LUT2 #(
		.INIT('h2)
	) name2948 (
		\g3002_reg/NET0131 ,
		\g3006_reg/NET0131 ,
		_w4128_
	);
	LUT2 #(
		.INIT('h4)
	) name2949 (
		\g3010_reg/NET0131 ,
		\g3013_reg/NET0131 ,
		_w4129_
	);
	LUT2 #(
		.INIT('h8)
	) name2950 (
		\g3024_reg/NET0131 ,
		_w4129_,
		_w4130_
	);
	LUT2 #(
		.INIT('h8)
	) name2951 (
		_w4127_,
		_w4128_,
		_w4131_
	);
	LUT2 #(
		.INIT('h8)
	) name2952 (
		_w4130_,
		_w4131_,
		_w4132_
	);
	LUT2 #(
		.INIT('h8)
	) name2953 (
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		_w4133_
	);
	LUT2 #(
		.INIT('h1)
	) name2954 (
		\g3032_reg/NET0131 ,
		\g3036_reg/NET0131 ,
		_w4134_
	);
	LUT2 #(
		.INIT('h8)
	) name2955 (
		_w4133_,
		_w4134_,
		_w4135_
	);
	LUT2 #(
		.INIT('h8)
	) name2956 (
		_w4132_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h2)
	) name2957 (
		_w2929_,
		_w4136_,
		_w4137_
	);
	LUT2 #(
		.INIT('h2)
	) name2958 (
		\g1018_reg/NET0131 ,
		\g1272_reg/NET0131 ,
		_w4138_
	);
	LUT2 #(
		.INIT('h4)
	) name2959 (
		\g1271_reg/NET0131 ,
		\g5657_pad ,
		_w4139_
	);
	LUT2 #(
		.INIT('h2)
	) name2960 (
		\g1024_reg/NET0131 ,
		\g1270_reg/NET0131 ,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name2961 (
		_w4138_,
		_w4139_,
		_w4141_
	);
	LUT2 #(
		.INIT('h4)
	) name2962 (
		_w4140_,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name2963 (
		\g1024_reg/NET0131 ,
		\g1261_reg/NET0131 ,
		_w4143_
	);
	LUT2 #(
		.INIT('h2)
	) name2964 (
		\g1018_reg/NET0131 ,
		\g1263_reg/NET0131 ,
		_w4144_
	);
	LUT2 #(
		.INIT('h4)
	) name2965 (
		\g1262_reg/NET0131 ,
		\g5657_pad ,
		_w4145_
	);
	LUT2 #(
		.INIT('h1)
	) name2966 (
		_w4143_,
		_w4144_,
		_w4146_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		_w4145_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h2)
	) name2968 (
		_w4142_,
		_w4147_,
		_w4148_
	);
	LUT2 #(
		.INIT('h2)
	) name2969 (
		\g1018_reg/NET0131 ,
		\g1266_reg/NET0131 ,
		_w4149_
	);
	LUT2 #(
		.INIT('h4)
	) name2970 (
		\g1265_reg/NET0131 ,
		\g5657_pad ,
		_w4150_
	);
	LUT2 #(
		.INIT('h2)
	) name2971 (
		\g1024_reg/NET0131 ,
		\g1264_reg/NET0131 ,
		_w4151_
	);
	LUT2 #(
		.INIT('h1)
	) name2972 (
		_w4149_,
		_w4150_,
		_w4152_
	);
	LUT2 #(
		.INIT('h4)
	) name2973 (
		_w4151_,
		_w4152_,
		_w4153_
	);
	LUT2 #(
		.INIT('h8)
	) name2974 (
		\g1066_reg/NET0131 ,
		\g5657_pad ,
		_w4154_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		\g1018_reg/NET0131 ,
		\g1068_reg/NET0131 ,
		_w4155_
	);
	LUT2 #(
		.INIT('h8)
	) name2976 (
		\g1024_reg/NET0131 ,
		\g1070_reg/NET0131 ,
		_w4156_
	);
	LUT2 #(
		.INIT('h1)
	) name2977 (
		_w4154_,
		_w4155_,
		_w4157_
	);
	LUT2 #(
		.INIT('h4)
	) name2978 (
		_w4156_,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h8)
	) name2979 (
		\g1051_reg/NET0131 ,
		\g5657_pad ,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name2980 (
		\g1018_reg/NET0131 ,
		\g1053_reg/NET0131 ,
		_w4160_
	);
	LUT2 #(
		.INIT('h8)
	) name2981 (
		\g1024_reg/NET0131 ,
		\g1055_reg/NET0131 ,
		_w4161_
	);
	LUT2 #(
		.INIT('h1)
	) name2982 (
		_w4159_,
		_w4160_,
		_w4162_
	);
	LUT2 #(
		.INIT('h4)
	) name2983 (
		_w4161_,
		_w4162_,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name2984 (
		_w4158_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h8)
	) name2985 (
		\g1036_reg/NET0131 ,
		\g5657_pad ,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name2986 (
		\g1024_reg/NET0131 ,
		\g1040_reg/NET0131 ,
		_w4166_
	);
	LUT2 #(
		.INIT('h8)
	) name2987 (
		\g1018_reg/NET0131 ,
		\g1038_reg/NET0131 ,
		_w4167_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w4165_,
		_w4166_,
		_w4168_
	);
	LUT2 #(
		.INIT('h4)
	) name2989 (
		_w4167_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('h8)
	) name2990 (
		_w4153_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h8)
	) name2991 (
		_w4164_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		_w4148_,
		_w4171_,
		_w4172_
	);
	LUT2 #(
		.INIT('h4)
	) name2993 (
		\g1268_reg/NET0131 ,
		\g5657_pad ,
		_w4173_
	);
	LUT2 #(
		.INIT('h2)
	) name2994 (
		\g1024_reg/NET0131 ,
		\g1267_reg/NET0131 ,
		_w4174_
	);
	LUT2 #(
		.INIT('h2)
	) name2995 (
		\g1018_reg/NET0131 ,
		\g1269_reg/NET0131 ,
		_w4175_
	);
	LUT2 #(
		.INIT('h1)
	) name2996 (
		_w4173_,
		_w4174_,
		_w4176_
	);
	LUT2 #(
		.INIT('h4)
	) name2997 (
		_w4175_,
		_w4176_,
		_w4177_
	);
	LUT2 #(
		.INIT('h2)
	) name2998 (
		_w4163_,
		_w4177_,
		_w4178_
	);
	LUT2 #(
		.INIT('h2)
	) name2999 (
		_w4147_,
		_w4169_,
		_w4179_
	);
	LUT2 #(
		.INIT('h8)
	) name3000 (
		_w4178_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h8)
	) name3001 (
		_w4147_,
		_w4153_,
		_w4181_
	);
	LUT2 #(
		.INIT('h2)
	) name3002 (
		_w4158_,
		_w4169_,
		_w4182_
	);
	LUT2 #(
		.INIT('h8)
	) name3003 (
		_w4142_,
		_w4181_,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name3004 (
		_w4182_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h8)
	) name3005 (
		_w4163_,
		_w4169_,
		_w4185_
	);
	LUT2 #(
		.INIT('h4)
	) name3006 (
		_w4153_,
		_w4177_,
		_w4186_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		_w4185_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h4)
	) name3008 (
		_w4158_,
		_w4163_,
		_w4188_
	);
	LUT2 #(
		.INIT('h2)
	) name3009 (
		_w4147_,
		_w4153_,
		_w4189_
	);
	LUT2 #(
		.INIT('h8)
	) name3010 (
		_w4188_,
		_w4189_,
		_w4190_
	);
	LUT2 #(
		.INIT('h2)
	) name3011 (
		_w4164_,
		_w4169_,
		_w4191_
	);
	LUT2 #(
		.INIT('h4)
	) name3012 (
		_w4142_,
		_w4191_,
		_w4192_
	);
	LUT2 #(
		.INIT('h8)
	) name3013 (
		_w4158_,
		_w4169_,
		_w4193_
	);
	LUT2 #(
		.INIT('h4)
	) name3014 (
		_w4153_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h8)
	) name3015 (
		_w4153_,
		_w4177_,
		_w4195_
	);
	LUT2 #(
		.INIT('h8)
	) name3016 (
		\g1081_reg/NET0131 ,
		\g5657_pad ,
		_w4196_
	);
	LUT2 #(
		.INIT('h8)
	) name3017 (
		\g1018_reg/NET0131 ,
		\g1083_reg/NET0131 ,
		_w4197_
	);
	LUT2 #(
		.INIT('h8)
	) name3018 (
		\g1011_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		_w4198_
	);
	LUT2 #(
		.INIT('h1)
	) name3019 (
		_w4196_,
		_w4197_,
		_w4199_
	);
	LUT2 #(
		.INIT('h4)
	) name3020 (
		_w4198_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h8)
	) name3021 (
		_w4195_,
		_w4200_,
		_w4201_
	);
	LUT2 #(
		.INIT('h1)
	) name3022 (
		_w4194_,
		_w4201_,
		_w4202_
	);
	LUT2 #(
		.INIT('h1)
	) name3023 (
		_w4147_,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h1)
	) name3024 (
		_w4147_,
		_w4177_,
		_w4204_
	);
	LUT2 #(
		.INIT('h1)
	) name3025 (
		_w4179_,
		_w4204_,
		_w4205_
	);
	LUT2 #(
		.INIT('h1)
	) name3026 (
		_w4163_,
		_w4200_,
		_w4206_
	);
	LUT2 #(
		.INIT('h1)
	) name3027 (
		_w4169_,
		_w4195_,
		_w4207_
	);
	LUT2 #(
		.INIT('h4)
	) name3028 (
		_w4205_,
		_w4206_,
		_w4208_
	);
	LUT2 #(
		.INIT('h4)
	) name3029 (
		_w4207_,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name3030 (
		_w4180_,
		_w4187_,
		_w4210_
	);
	LUT2 #(
		.INIT('h4)
	) name3031 (
		_w4190_,
		_w4210_,
		_w4211_
	);
	LUT2 #(
		.INIT('h1)
	) name3032 (
		_w4172_,
		_w4184_,
		_w4212_
	);
	LUT2 #(
		.INIT('h4)
	) name3033 (
		_w4192_,
		_w4212_,
		_w4213_
	);
	LUT2 #(
		.INIT('h4)
	) name3034 (
		_w4203_,
		_w4211_,
		_w4214_
	);
	LUT2 #(
		.INIT('h4)
	) name3035 (
		_w4209_,
		_w4214_,
		_w4215_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		_w4213_,
		_w4215_,
		_w4216_
	);
	LUT2 #(
		.INIT('h8)
	) name3037 (
		\g1282_reg/NET0131 ,
		\g5657_pad ,
		_w4217_
	);
	LUT2 #(
		.INIT('h8)
	) name3038 (
		\g1024_reg/NET0131 ,
		\g1288_reg/NET0131 ,
		_w4218_
	);
	LUT2 #(
		.INIT('h8)
	) name3039 (
		\g1018_reg/NET0131 ,
		\g1285_reg/NET0131 ,
		_w4219_
	);
	LUT2 #(
		.INIT('h8)
	) name3040 (
		\g1251_reg/NET0131 ,
		\g5657_pad ,
		_w4220_
	);
	LUT2 #(
		.INIT('h8)
	) name3041 (
		\g1024_reg/NET0131 ,
		\g1176_reg/NET0131 ,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name3042 (
		\g1018_reg/NET0131 ,
		\g1253_reg/NET0131 ,
		_w4222_
	);
	LUT2 #(
		.INIT('h1)
	) name3043 (
		_w4220_,
		_w4221_,
		_w4223_
	);
	LUT2 #(
		.INIT('h4)
	) name3044 (
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name3045 (
		\g1228_reg/NET0131 ,
		\g185_reg/NET0131 ,
		_w4225_
	);
	LUT2 #(
		.INIT('h4)
	) name3046 (
		_w4224_,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h1)
	) name3047 (
		_w4217_,
		_w4218_,
		_w4227_
	);
	LUT2 #(
		.INIT('h4)
	) name3048 (
		_w4219_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h4)
	) name3049 (
		_w4226_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h4)
	) name3050 (
		_w4147_,
		_w4153_,
		_w4230_
	);
	LUT2 #(
		.INIT('h8)
	) name3051 (
		_w4185_,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name3052 (
		_w4147_,
		_w4177_,
		_w4232_
	);
	LUT2 #(
		.INIT('h8)
	) name3053 (
		_w4191_,
		_w4232_,
		_w4233_
	);
	LUT2 #(
		.INIT('h1)
	) name3054 (
		_w4142_,
		_w4147_,
		_w4234_
	);
	LUT2 #(
		.INIT('h4)
	) name3055 (
		_w4200_,
		_w4234_,
		_w4235_
	);
	LUT2 #(
		.INIT('h4)
	) name3056 (
		_w4163_,
		_w4195_,
		_w4236_
	);
	LUT2 #(
		.INIT('h2)
	) name3057 (
		_w4142_,
		_w4236_,
		_w4237_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		_w4158_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h2)
	) name3059 (
		_w4169_,
		_w4235_,
		_w4239_
	);
	LUT2 #(
		.INIT('h4)
	) name3060 (
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT2 #(
		.INIT('h8)
	) name3061 (
		_w4186_,
		_w4206_,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name3062 (
		_w4148_,
		_w4188_,
		_w4242_
	);
	LUT2 #(
		.INIT('h1)
	) name3063 (
		_w4169_,
		_w4241_,
		_w4243_
	);
	LUT2 #(
		.INIT('h4)
	) name3064 (
		_w4242_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		_w4240_,
		_w4244_,
		_w4245_
	);
	LUT2 #(
		.INIT('h2)
	) name3066 (
		_w4142_,
		_w4169_,
		_w4246_
	);
	LUT2 #(
		.INIT('h2)
	) name3067 (
		_w4177_,
		_w4246_,
		_w4247_
	);
	LUT2 #(
		.INIT('h2)
	) name3068 (
		_w4200_,
		_w4247_,
		_w4248_
	);
	LUT2 #(
		.INIT('h1)
	) name3069 (
		_w4171_,
		_w4248_,
		_w4249_
	);
	LUT2 #(
		.INIT('h2)
	) name3070 (
		_w4147_,
		_w4249_,
		_w4250_
	);
	LUT2 #(
		.INIT('h4)
	) name3071 (
		_w4147_,
		_w4178_,
		_w4251_
	);
	LUT2 #(
		.INIT('h4)
	) name3072 (
		_w4193_,
		_w4251_,
		_w4252_
	);
	LUT2 #(
		.INIT('h1)
	) name3073 (
		_w4153_,
		_w4178_,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name3074 (
		_w4182_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h1)
	) name3075 (
		_w4231_,
		_w4233_,
		_w4255_
	);
	LUT2 #(
		.INIT('h1)
	) name3076 (
		_w4252_,
		_w4254_,
		_w4256_
	);
	LUT2 #(
		.INIT('h8)
	) name3077 (
		_w4255_,
		_w4256_,
		_w4257_
	);
	LUT2 #(
		.INIT('h4)
	) name3078 (
		_w4250_,
		_w4257_,
		_w4258_
	);
	LUT2 #(
		.INIT('h4)
	) name3079 (
		_w4245_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name3080 (
		_w4229_,
		_w4259_,
		_w4260_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		\g1273_reg/NET0131 ,
		\g5657_pad ,
		_w4261_
	);
	LUT2 #(
		.INIT('h8)
	) name3082 (
		\g1018_reg/NET0131 ,
		\g1276_reg/NET0131 ,
		_w4262_
	);
	LUT2 #(
		.INIT('h8)
	) name3083 (
		\g1024_reg/NET0131 ,
		\g1279_reg/NET0131 ,
		_w4263_
	);
	LUT2 #(
		.INIT('h8)
	) name3084 (
		\g1018_reg/NET0131 ,
		\g1257_reg/NET0131 ,
		_w4264_
	);
	LUT2 #(
		.INIT('h8)
	) name3085 (
		\g1024_reg/NET0131 ,
		\g1259_reg/NET0131 ,
		_w4265_
	);
	LUT2 #(
		.INIT('h8)
	) name3086 (
		\g1255_reg/NET0131 ,
		\g5657_pad ,
		_w4266_
	);
	LUT2 #(
		.INIT('h1)
	) name3087 (
		_w4264_,
		_w4265_,
		_w4267_
	);
	LUT2 #(
		.INIT('h4)
	) name3088 (
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT2 #(
		.INIT('h8)
	) name3089 (
		\g1210_reg/NET0131 ,
		\g185_reg/NET0131 ,
		_w4269_
	);
	LUT2 #(
		.INIT('h4)
	) name3090 (
		_w4268_,
		_w4269_,
		_w4270_
	);
	LUT2 #(
		.INIT('h1)
	) name3091 (
		_w4261_,
		_w4262_,
		_w4271_
	);
	LUT2 #(
		.INIT('h4)
	) name3092 (
		_w4263_,
		_w4271_,
		_w4272_
	);
	LUT2 #(
		.INIT('h4)
	) name3093 (
		_w4270_,
		_w4272_,
		_w4273_
	);
	LUT2 #(
		.INIT('h1)
	) name3094 (
		_w4229_,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h2)
	) name3095 (
		_w4216_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h4)
	) name3096 (
		_w4260_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h2)
	) name3097 (
		_w4136_,
		_w4276_,
		_w4277_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		_w4137_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h2)
	) name3099 (
		\g1024_reg/NET0131 ,
		_w4278_,
		_w4279_
	);
	LUT2 #(
		.INIT('h1)
	) name3100 (
		\g1024_reg/NET0131 ,
		\g1306_reg/NET0131 ,
		_w4280_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w4279_,
		_w4280_,
		_w4281_
	);
	LUT2 #(
		.INIT('h2)
	) name3102 (
		_w1633_,
		_w4136_,
		_w4282_
	);
	LUT2 #(
		.INIT('h2)
	) name3103 (
		\g1018_reg/NET0131 ,
		\g2660_reg/NET0131 ,
		_w4283_
	);
	LUT2 #(
		.INIT('h2)
	) name3104 (
		\g1024_reg/NET0131 ,
		\g2658_reg/NET0131 ,
		_w4284_
	);
	LUT2 #(
		.INIT('h4)
	) name3105 (
		\g2659_reg/NET0131 ,
		\g5657_pad ,
		_w4285_
	);
	LUT2 #(
		.INIT('h1)
	) name3106 (
		_w4283_,
		_w4284_,
		_w4286_
	);
	LUT2 #(
		.INIT('h4)
	) name3107 (
		_w4285_,
		_w4286_,
		_w4287_
	);
	LUT2 #(
		.INIT('h8)
	) name3108 (
		\g2424_reg/NET0131 ,
		\g5657_pad ,
		_w4288_
	);
	LUT2 #(
		.INIT('h8)
	) name3109 (
		\g1024_reg/NET0131 ,
		\g2428_reg/NET0131 ,
		_w4289_
	);
	LUT2 #(
		.INIT('h8)
	) name3110 (
		\g1018_reg/NET0131 ,
		\g2426_reg/NET0131 ,
		_w4290_
	);
	LUT2 #(
		.INIT('h1)
	) name3111 (
		_w4288_,
		_w4289_,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name3112 (
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name3113 (
		\g2439_reg/NET0131 ,
		\g5657_pad ,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name3114 (
		\g1024_reg/NET0131 ,
		\g2443_reg/NET0131 ,
		_w4294_
	);
	LUT2 #(
		.INIT('h8)
	) name3115 (
		\g1018_reg/NET0131 ,
		\g2441_reg/NET0131 ,
		_w4295_
	);
	LUT2 #(
		.INIT('h1)
	) name3116 (
		_w4293_,
		_w4294_,
		_w4296_
	);
	LUT2 #(
		.INIT('h4)
	) name3117 (
		_w4295_,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h8)
	) name3118 (
		\g2454_reg/NET0131 ,
		\g5657_pad ,
		_w4298_
	);
	LUT2 #(
		.INIT('h8)
	) name3119 (
		\g1024_reg/NET0131 ,
		\g2458_reg/NET0131 ,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name3120 (
		\g1018_reg/NET0131 ,
		\g2456_reg/NET0131 ,
		_w4300_
	);
	LUT2 #(
		.INIT('h1)
	) name3121 (
		_w4298_,
		_w4299_,
		_w4301_
	);
	LUT2 #(
		.INIT('h4)
	) name3122 (
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('h1)
	) name3123 (
		_w4297_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h4)
	) name3124 (
		_w4292_,
		_w4303_,
		_w4304_
	);
	LUT2 #(
		.INIT('h4)
	) name3125 (
		_w4287_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name3126 (
		_w4292_,
		_w4302_,
		_w4306_
	);
	LUT2 #(
		.INIT('h2)
	) name3127 (
		\g1018_reg/NET0131 ,
		\g2654_reg/NET0131 ,
		_w4307_
	);
	LUT2 #(
		.INIT('h2)
	) name3128 (
		\g1024_reg/NET0131 ,
		\g2652_reg/NET0131 ,
		_w4308_
	);
	LUT2 #(
		.INIT('h4)
	) name3129 (
		\g2653_reg/NET0131 ,
		\g5657_pad ,
		_w4309_
	);
	LUT2 #(
		.INIT('h1)
	) name3130 (
		_w4307_,
		_w4308_,
		_w4310_
	);
	LUT2 #(
		.INIT('h4)
	) name3131 (
		_w4309_,
		_w4310_,
		_w4311_
	);
	LUT2 #(
		.INIT('h2)
	) name3132 (
		\g1024_reg/NET0131 ,
		\g2649_reg/NET0131 ,
		_w4312_
	);
	LUT2 #(
		.INIT('h2)
	) name3133 (
		\g1018_reg/NET0131 ,
		\g2651_reg/NET0131 ,
		_w4313_
	);
	LUT2 #(
		.INIT('h4)
	) name3134 (
		\g2650_reg/NET0131 ,
		\g5657_pad ,
		_w4314_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		_w4312_,
		_w4313_,
		_w4315_
	);
	LUT2 #(
		.INIT('h4)
	) name3136 (
		_w4314_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h1)
	) name3137 (
		_w4311_,
		_w4316_,
		_w4317_
	);
	LUT2 #(
		.INIT('h8)
	) name3138 (
		_w4306_,
		_w4317_,
		_w4318_
	);
	LUT2 #(
		.INIT('h8)
	) name3139 (
		_w4292_,
		_w4303_,
		_w4319_
	);
	LUT2 #(
		.INIT('h2)
	) name3140 (
		_w4311_,
		_w4316_,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name3141 (
		_w4287_,
		_w4320_,
		_w4321_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		_w4319_,
		_w4321_,
		_w4322_
	);
	LUT2 #(
		.INIT('h4)
	) name3143 (
		_w4292_,
		_w4297_,
		_w4323_
	);
	LUT2 #(
		.INIT('h2)
	) name3144 (
		\g1024_reg/NET0131 ,
		\g2655_reg/NET0131 ,
		_w4324_
	);
	LUT2 #(
		.INIT('h4)
	) name3145 (
		\g2656_reg/NET0131 ,
		\g5657_pad ,
		_w4325_
	);
	LUT2 #(
		.INIT('h2)
	) name3146 (
		\g1018_reg/NET0131 ,
		\g2657_reg/NET0131 ,
		_w4326_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w4324_,
		_w4325_,
		_w4327_
	);
	LUT2 #(
		.INIT('h4)
	) name3148 (
		_w4326_,
		_w4327_,
		_w4328_
	);
	LUT2 #(
		.INIT('h2)
	) name3149 (
		_w4316_,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h8)
	) name3150 (
		_w4323_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h2)
	) name3151 (
		_w4297_,
		_w4302_,
		_w4331_
	);
	LUT2 #(
		.INIT('h4)
	) name3152 (
		_w4311_,
		_w4316_,
		_w4332_
	);
	LUT2 #(
		.INIT('h8)
	) name3153 (
		_w4331_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h4)
	) name3154 (
		_w4292_,
		_w4302_,
		_w4334_
	);
	LUT2 #(
		.INIT('h8)
	) name3155 (
		_w4311_,
		_w4316_,
		_w4335_
	);
	LUT2 #(
		.INIT('h8)
	) name3156 (
		_w4287_,
		_w4335_,
		_w4336_
	);
	LUT2 #(
		.INIT('h8)
	) name3157 (
		_w4334_,
		_w4336_,
		_w4337_
	);
	LUT2 #(
		.INIT('h8)
	) name3158 (
		\g2469_reg/NET0131 ,
		\g5657_pad ,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name3159 (
		\g1024_reg/NET0131 ,
		\g2399_reg/NET0131 ,
		_w4339_
	);
	LUT2 #(
		.INIT('h8)
	) name3160 (
		\g1018_reg/NET0131 ,
		\g2471_reg/NET0131 ,
		_w4340_
	);
	LUT2 #(
		.INIT('h1)
	) name3161 (
		_w4338_,
		_w4339_,
		_w4341_
	);
	LUT2 #(
		.INIT('h4)
	) name3162 (
		_w4340_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h1)
	) name3163 (
		_w4297_,
		_w4342_,
		_w4343_
	);
	LUT2 #(
		.INIT('h4)
	) name3164 (
		_w4292_,
		_w4316_,
		_w4344_
	);
	LUT2 #(
		.INIT('h8)
	) name3165 (
		_w4311_,
		_w4328_,
		_w4345_
	);
	LUT2 #(
		.INIT('h8)
	) name3166 (
		_w4344_,
		_w4345_,
		_w4346_
	);
	LUT2 #(
		.INIT('h2)
	) name3167 (
		_w4292_,
		_w4316_,
		_w4347_
	);
	LUT2 #(
		.INIT('h4)
	) name3168 (
		_w4328_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h1)
	) name3169 (
		_w4346_,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('h2)
	) name3170 (
		_w4343_,
		_w4349_,
		_w4350_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		_w4292_,
		_w4297_,
		_w4351_
	);
	LUT2 #(
		.INIT('h4)
	) name3172 (
		_w4311_,
		_w4351_,
		_w4352_
	);
	LUT2 #(
		.INIT('h8)
	) name3173 (
		_w4320_,
		_w4342_,
		_w4353_
	);
	LUT2 #(
		.INIT('h1)
	) name3174 (
		_w4352_,
		_w4353_,
		_w4354_
	);
	LUT2 #(
		.INIT('h2)
	) name3175 (
		_w4328_,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('h1)
	) name3176 (
		_w4318_,
		_w4330_,
		_w4356_
	);
	LUT2 #(
		.INIT('h4)
	) name3177 (
		_w4333_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h1)
	) name3178 (
		_w4305_,
		_w4322_,
		_w4358_
	);
	LUT2 #(
		.INIT('h4)
	) name3179 (
		_w4337_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h4)
	) name3180 (
		_w4350_,
		_w4357_,
		_w4360_
	);
	LUT2 #(
		.INIT('h4)
	) name3181 (
		_w4355_,
		_w4360_,
		_w4361_
	);
	LUT2 #(
		.INIT('h8)
	) name3182 (
		_w4359_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h8)
	) name3183 (
		\g2670_reg/NET0131 ,
		\g5657_pad ,
		_w4363_
	);
	LUT2 #(
		.INIT('h8)
	) name3184 (
		\g1018_reg/NET0131 ,
		\g2673_reg/NET0131 ,
		_w4364_
	);
	LUT2 #(
		.INIT('h8)
	) name3185 (
		\g1024_reg/NET0131 ,
		\g2676_reg/NET0131 ,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name3186 (
		\g2639_reg/NET0131 ,
		\g5657_pad ,
		_w4366_
	);
	LUT2 #(
		.INIT('h8)
	) name3187 (
		\g1018_reg/NET0131 ,
		\g2641_reg/NET0131 ,
		_w4367_
	);
	LUT2 #(
		.INIT('h8)
	) name3188 (
		\g1024_reg/NET0131 ,
		\g2564_reg/NET0131 ,
		_w4368_
	);
	LUT2 #(
		.INIT('h1)
	) name3189 (
		_w4366_,
		_w4367_,
		_w4369_
	);
	LUT2 #(
		.INIT('h4)
	) name3190 (
		_w4368_,
		_w4369_,
		_w4370_
	);
	LUT2 #(
		.INIT('h8)
	) name3191 (
		\g185_reg/NET0131 ,
		\g2616_reg/NET0131 ,
		_w4371_
	);
	LUT2 #(
		.INIT('h4)
	) name3192 (
		_w4370_,
		_w4371_,
		_w4372_
	);
	LUT2 #(
		.INIT('h1)
	) name3193 (
		_w4363_,
		_w4364_,
		_w4373_
	);
	LUT2 #(
		.INIT('h4)
	) name3194 (
		_w4365_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h4)
	) name3195 (
		_w4372_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h8)
	) name3196 (
		_w4320_,
		_w4351_,
		_w4376_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		_w4316_,
		_w4328_,
		_w4377_
	);
	LUT2 #(
		.INIT('h8)
	) name3198 (
		_w4323_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h4)
	) name3199 (
		_w4342_,
		_w4347_,
		_w4379_
	);
	LUT2 #(
		.INIT('h1)
	) name3200 (
		_w4306_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name3201 (
		_w4287_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h1)
	) name3202 (
		_w4297_,
		_w4311_,
		_w4382_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		_w4334_,
		_w4382_,
		_w4383_
	);
	LUT2 #(
		.INIT('h8)
	) name3204 (
		_w4287_,
		_w4342_,
		_w4384_
	);
	LUT2 #(
		.INIT('h8)
	) name3205 (
		_w4344_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h4)
	) name3206 (
		_w4297_,
		_w4306_,
		_w4386_
	);
	LUT2 #(
		.INIT('h8)
	) name3207 (
		_w4345_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h8)
	) name3208 (
		_w4319_,
		_w4335_,
		_w4388_
	);
	LUT2 #(
		.INIT('h1)
	) name3209 (
		_w4304_,
		_w4342_,
		_w4389_
	);
	LUT2 #(
		.INIT('h2)
	) name3210 (
		_w4329_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name3211 (
		_w4287_,
		_w4316_,
		_w4391_
	);
	LUT2 #(
		.INIT('h4)
	) name3212 (
		_w4292_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h1)
	) name3213 (
		_w4377_,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		_w4331_,
		_w4393_,
		_w4394_
	);
	LUT2 #(
		.INIT('h4)
	) name3215 (
		_w4311_,
		_w4328_,
		_w4395_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		_w4302_,
		_w4343_,
		_w4396_
	);
	LUT2 #(
		.INIT('h4)
	) name3217 (
		_w4292_,
		_w4395_,
		_w4397_
	);
	LUT2 #(
		.INIT('h4)
	) name3218 (
		_w4396_,
		_w4397_,
		_w4398_
	);
	LUT2 #(
		.INIT('h1)
	) name3219 (
		_w4376_,
		_w4378_,
		_w4399_
	);
	LUT2 #(
		.INIT('h1)
	) name3220 (
		_w4383_,
		_w4385_,
		_w4400_
	);
	LUT2 #(
		.INIT('h8)
	) name3221 (
		_w4399_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h1)
	) name3222 (
		_w4387_,
		_w4388_,
		_w4402_
	);
	LUT2 #(
		.INIT('h4)
	) name3223 (
		_w4398_,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('h4)
	) name3224 (
		_w4381_,
		_w4401_,
		_w4404_
	);
	LUT2 #(
		.INIT('h1)
	) name3225 (
		_w4390_,
		_w4394_,
		_w4405_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		_w4404_,
		_w4405_,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name3227 (
		_w4403_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		_w4375_,
		_w4407_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name3229 (
		\g2661_reg/NET0131 ,
		\g5657_pad ,
		_w4409_
	);
	LUT2 #(
		.INIT('h8)
	) name3230 (
		\g1018_reg/NET0131 ,
		\g2664_reg/NET0131 ,
		_w4410_
	);
	LUT2 #(
		.INIT('h8)
	) name3231 (
		\g1024_reg/NET0131 ,
		\g2667_reg/NET0131 ,
		_w4411_
	);
	LUT2 #(
		.INIT('h8)
	) name3232 (
		\g1018_reg/NET0131 ,
		\g2645_reg/NET0131 ,
		_w4412_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		\g1024_reg/NET0131 ,
		\g2647_reg/NET0131 ,
		_w4413_
	);
	LUT2 #(
		.INIT('h8)
	) name3234 (
		\g2643_reg/NET0131 ,
		\g5657_pad ,
		_w4414_
	);
	LUT2 #(
		.INIT('h1)
	) name3235 (
		_w4412_,
		_w4413_,
		_w4415_
	);
	LUT2 #(
		.INIT('h4)
	) name3236 (
		_w4414_,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h8)
	) name3237 (
		\g185_reg/NET0131 ,
		\g2598_reg/NET0131 ,
		_w4417_
	);
	LUT2 #(
		.INIT('h4)
	) name3238 (
		_w4416_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h1)
	) name3239 (
		_w4409_,
		_w4410_,
		_w4419_
	);
	LUT2 #(
		.INIT('h4)
	) name3240 (
		_w4411_,
		_w4419_,
		_w4420_
	);
	LUT2 #(
		.INIT('h4)
	) name3241 (
		_w4418_,
		_w4420_,
		_w4421_
	);
	LUT2 #(
		.INIT('h1)
	) name3242 (
		_w4375_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h2)
	) name3243 (
		_w4362_,
		_w4422_,
		_w4423_
	);
	LUT2 #(
		.INIT('h4)
	) name3244 (
		_w4408_,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h2)
	) name3245 (
		_w4136_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('h1)
	) name3246 (
		_w4282_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h2)
	) name3247 (
		\g5657_pad ,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h1)
	) name3248 (
		\g2688_reg/NET0131 ,
		\g5657_pad ,
		_w4428_
	);
	LUT2 #(
		.INIT('h1)
	) name3249 (
		_w4427_,
		_w4428_,
		_w4429_
	);
	LUT2 #(
		.INIT('h2)
	) name3250 (
		\g1018_reg/NET0131 ,
		_w4426_,
		_w4430_
	);
	LUT2 #(
		.INIT('h1)
	) name3251 (
		\g1018_reg/NET0131 ,
		\g2691_reg/NET0131 ,
		_w4431_
	);
	LUT2 #(
		.INIT('h1)
	) name3252 (
		_w4430_,
		_w4431_,
		_w4432_
	);
	LUT2 #(
		.INIT('h2)
	) name3253 (
		\g1024_reg/NET0131 ,
		_w4426_,
		_w4433_
	);
	LUT2 #(
		.INIT('h1)
	) name3254 (
		\g1024_reg/NET0131 ,
		\g2694_reg/NET0131 ,
		_w4434_
	);
	LUT2 #(
		.INIT('h1)
	) name3255 (
		_w4433_,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('h2)
	) name3256 (
		_w1901_,
		_w3749_,
		_w4436_
	);
	LUT2 #(
		.INIT('h1)
	) name3257 (
		\g536_reg/NET0131 ,
		_w4087_,
		_w4437_
	);
	LUT2 #(
		.INIT('h8)
	) name3258 (
		_w3766_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h8)
	) name3259 (
		_w3803_,
		_w4087_,
		_w4439_
	);
	LUT2 #(
		.INIT('h1)
	) name3260 (
		_w4086_,
		_w4438_,
		_w4440_
	);
	LUT2 #(
		.INIT('h4)
	) name3261 (
		_w4439_,
		_w4440_,
		_w4441_
	);
	LUT2 #(
		.INIT('h1)
	) name3262 (
		_w4436_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h2)
	) name3263 (
		_w1901_,
		_w3760_,
		_w4443_
	);
	LUT2 #(
		.INIT('h1)
	) name3264 (
		\g537_reg/NET0131 ,
		_w4087_,
		_w4444_
	);
	LUT2 #(
		.INIT('h8)
	) name3265 (
		_w3766_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h8)
	) name3266 (
		_w3797_,
		_w4087_,
		_w4446_
	);
	LUT2 #(
		.INIT('h1)
	) name3267 (
		_w4086_,
		_w4445_,
		_w4447_
	);
	LUT2 #(
		.INIT('h4)
	) name3268 (
		_w4446_,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h1)
	) name3269 (
		_w4443_,
		_w4448_,
		_w4449_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w1643_,
		_w4136_,
		_w4450_
	);
	LUT2 #(
		.INIT('h8)
	) name3271 (
		_w4362_,
		_w4421_,
		_w4451_
	);
	LUT2 #(
		.INIT('h2)
	) name3272 (
		_w4136_,
		_w4422_,
		_w4452_
	);
	LUT2 #(
		.INIT('h8)
	) name3273 (
		_w4407_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h4)
	) name3274 (
		_w4451_,
		_w4453_,
		_w4454_
	);
	LUT2 #(
		.INIT('h1)
	) name3275 (
		_w4450_,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('h2)
	) name3276 (
		\g5657_pad ,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h2)
	) name3277 (
		\g2679_reg/NET0131 ,
		\g5657_pad ,
		_w4457_
	);
	LUT2 #(
		.INIT('h1)
	) name3278 (
		_w4456_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h2)
	) name3279 (
		\g1018_reg/NET0131 ,
		_w4455_,
		_w4459_
	);
	LUT2 #(
		.INIT('h4)
	) name3280 (
		\g1018_reg/NET0131 ,
		\g2682_reg/NET0131 ,
		_w4460_
	);
	LUT2 #(
		.INIT('h1)
	) name3281 (
		_w4459_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h2)
	) name3282 (
		\g1024_reg/NET0131 ,
		_w4455_,
		_w4462_
	);
	LUT2 #(
		.INIT('h4)
	) name3283 (
		\g1024_reg/NET0131 ,
		\g2685_reg/NET0131 ,
		_w4463_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		_w4462_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h4)
	) name3285 (
		_w2019_,
		_w3070_,
		_w4465_
	);
	LUT2 #(
		.INIT('h1)
	) name3286 (
		_w3066_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h2)
	) name3287 (
		_w2135_,
		_w4466_,
		_w4467_
	);
	LUT2 #(
		.INIT('h8)
	) name3288 (
		_w1292_,
		_w3320_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name3289 (
		_w3326_,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h1)
	) name3290 (
		_w3140_,
		_w3145_,
		_w4470_
	);
	LUT2 #(
		.INIT('h2)
	) name3291 (
		_w2399_,
		_w2408_,
		_w4471_
	);
	LUT2 #(
		.INIT('h4)
	) name3292 (
		_w4470_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h4)
	) name3293 (
		_w2574_,
		_w3268_,
		_w4473_
	);
	LUT2 #(
		.INIT('h8)
	) name3294 (
		_w2816_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h1)
	) name3295 (
		_w3275_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h4)
	) name3296 (
		\g1345_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		_w4476_
	);
	LUT2 #(
		.INIT('h8)
	) name3297 (
		\g2612_reg/NET0131 ,
		_w4476_,
		_w4477_
	);
	LUT2 #(
		.INIT('h8)
	) name3298 (
		\g5657_pad ,
		_w4477_,
		_w4478_
	);
	LUT2 #(
		.INIT('h2)
	) name3299 (
		\g2809_reg/NET0131 ,
		_w4478_,
		_w4479_
	);
	LUT2 #(
		.INIT('h2)
	) name3300 (
		\g1018_reg/NET0131 ,
		\g2804_reg/NET0131 ,
		_w4480_
	);
	LUT2 #(
		.INIT('h4)
	) name3301 (
		\g2803_reg/NET0131 ,
		\g5657_pad ,
		_w4481_
	);
	LUT2 #(
		.INIT('h2)
	) name3302 (
		\g1024_reg/NET0131 ,
		\g2802_reg/NET0131 ,
		_w4482_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		\g1346_reg/NET0131 ,
		_w1596_,
		_w4483_
	);
	LUT2 #(
		.INIT('h1)
	) name3304 (
		\g1352_reg/NET0131 ,
		_w1586_,
		_w4484_
	);
	LUT2 #(
		.INIT('h8)
	) name3305 (
		\g1352_reg/NET0131 ,
		_w1586_,
		_w4485_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		\g1372_reg/NET0131 ,
		_w1561_,
		_w4486_
	);
	LUT2 #(
		.INIT('h1)
	) name3307 (
		\g1319_reg/NET0131 ,
		_w1616_,
		_w4487_
	);
	LUT2 #(
		.INIT('h8)
	) name3308 (
		\g1339_reg/NET0131 ,
		_w1581_,
		_w4488_
	);
	LUT2 #(
		.INIT('h1)
	) name3309 (
		\g1378_reg/NET0131 ,
		_w1611_,
		_w4489_
	);
	LUT2 #(
		.INIT('h1)
	) name3310 (
		\g1332_reg/NET0131 ,
		_w1571_,
		_w4490_
	);
	LUT2 #(
		.INIT('h8)
	) name3311 (
		\g1319_reg/NET0131 ,
		_w1616_,
		_w4491_
	);
	LUT2 #(
		.INIT('h8)
	) name3312 (
		\g1332_reg/NET0131 ,
		_w1571_,
		_w4492_
	);
	LUT2 #(
		.INIT('h8)
	) name3313 (
		\g1346_reg/NET0131 ,
		_w1596_,
		_w4493_
	);
	LUT2 #(
		.INIT('h1)
	) name3314 (
		\g1326_reg/NET0131 ,
		_w1576_,
		_w4494_
	);
	LUT2 #(
		.INIT('h8)
	) name3315 (
		\g1372_reg/NET0131 ,
		_w1561_,
		_w4495_
	);
	LUT2 #(
		.INIT('h8)
	) name3316 (
		\g1378_reg/NET0131 ,
		_w1611_,
		_w4496_
	);
	LUT2 #(
		.INIT('h1)
	) name3317 (
		\g1339_reg/NET0131 ,
		_w1581_,
		_w4497_
	);
	LUT2 #(
		.INIT('h8)
	) name3318 (
		\g1365_reg/NET0131 ,
		_w1566_,
		_w4498_
	);
	LUT2 #(
		.INIT('h8)
	) name3319 (
		\g1358_reg/NET0131 ,
		_w1591_,
		_w4499_
	);
	LUT2 #(
		.INIT('h8)
	) name3320 (
		\g1326_reg/NET0131 ,
		_w1576_,
		_w4500_
	);
	LUT2 #(
		.INIT('h1)
	) name3321 (
		\g1365_reg/NET0131 ,
		_w1566_,
		_w4501_
	);
	LUT2 #(
		.INIT('h1)
	) name3322 (
		\g1358_reg/NET0131 ,
		_w1591_,
		_w4502_
	);
	LUT2 #(
		.INIT('h1)
	) name3323 (
		_w4483_,
		_w4484_,
		_w4503_
	);
	LUT2 #(
		.INIT('h1)
	) name3324 (
		_w4485_,
		_w4486_,
		_w4504_
	);
	LUT2 #(
		.INIT('h1)
	) name3325 (
		_w4487_,
		_w4488_,
		_w4505_
	);
	LUT2 #(
		.INIT('h1)
	) name3326 (
		_w4489_,
		_w4490_,
		_w4506_
	);
	LUT2 #(
		.INIT('h1)
	) name3327 (
		_w4491_,
		_w4492_,
		_w4507_
	);
	LUT2 #(
		.INIT('h1)
	) name3328 (
		_w4493_,
		_w4494_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name3329 (
		_w4495_,
		_w4496_,
		_w4509_
	);
	LUT2 #(
		.INIT('h1)
	) name3330 (
		_w4497_,
		_w4498_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name3331 (
		_w4499_,
		_w4500_,
		_w4511_
	);
	LUT2 #(
		.INIT('h1)
	) name3332 (
		_w4501_,
		_w4502_,
		_w4512_
	);
	LUT2 #(
		.INIT('h8)
	) name3333 (
		_w4511_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		_w4509_,
		_w4510_,
		_w4514_
	);
	LUT2 #(
		.INIT('h8)
	) name3335 (
		_w4507_,
		_w4508_,
		_w4515_
	);
	LUT2 #(
		.INIT('h8)
	) name3336 (
		_w4505_,
		_w4506_,
		_w4516_
	);
	LUT2 #(
		.INIT('h8)
	) name3337 (
		_w4503_,
		_w4504_,
		_w4517_
	);
	LUT2 #(
		.INIT('h8)
	) name3338 (
		_w4516_,
		_w4517_,
		_w4518_
	);
	LUT2 #(
		.INIT('h8)
	) name3339 (
		_w4514_,
		_w4515_,
		_w4519_
	);
	LUT2 #(
		.INIT('h8)
	) name3340 (
		_w4513_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h8)
	) name3341 (
		_w4518_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h1)
	) name3342 (
		_w4480_,
		_w4481_,
		_w4522_
	);
	LUT2 #(
		.INIT('h4)
	) name3343 (
		_w4482_,
		_w4522_,
		_w4523_
	);
	LUT2 #(
		.INIT('h8)
	) name3344 (
		_w1606_,
		_w4523_,
		_w4524_
	);
	LUT2 #(
		.INIT('h4)
	) name3345 (
		_w4521_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h8)
	) name3346 (
		_w4478_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w4479_,
		_w4526_,
		_w4527_
	);
	LUT2 #(
		.INIT('h8)
	) name3348 (
		\g1018_reg/NET0131 ,
		_w4477_,
		_w4528_
	);
	LUT2 #(
		.INIT('h2)
	) name3349 (
		\g2810_reg/NET0131 ,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h8)
	) name3350 (
		_w4525_,
		_w4528_,
		_w4530_
	);
	LUT2 #(
		.INIT('h1)
	) name3351 (
		_w4529_,
		_w4530_,
		_w4531_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		\g1211_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w4532_
	);
	LUT2 #(
		.INIT('h4)
	) name3353 (
		\g1345_reg/NET0131 ,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h8)
	) name3354 (
		\g1024_reg/NET0131 ,
		_w4533_,
		_w4534_
	);
	LUT2 #(
		.INIT('h2)
	) name3355 (
		\g1420_reg/NET0131 ,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h2)
	) name3356 (
		\g1018_reg/NET0131 ,
		\g1416_reg/NET0131 ,
		_w4536_
	);
	LUT2 #(
		.INIT('h4)
	) name3357 (
		\g1415_reg/NET0131 ,
		\g5657_pad ,
		_w4537_
	);
	LUT2 #(
		.INIT('h2)
	) name3358 (
		\g1024_reg/NET0131 ,
		\g1414_reg/NET0131 ,
		_w4538_
	);
	LUT2 #(
		.INIT('h1)
	) name3359 (
		\g1339_reg/NET0131 ,
		_w2912_,
		_w4539_
	);
	LUT2 #(
		.INIT('h1)
	) name3360 (
		\g1372_reg/NET0131 ,
		_w2857_,
		_w4540_
	);
	LUT2 #(
		.INIT('h8)
	) name3361 (
		\g1372_reg/NET0131 ,
		_w2857_,
		_w4541_
	);
	LUT2 #(
		.INIT('h1)
	) name3362 (
		\g1365_reg/NET0131 ,
		_w2892_,
		_w4542_
	);
	LUT2 #(
		.INIT('h1)
	) name3363 (
		\g1346_reg/NET0131 ,
		_w2862_,
		_w4543_
	);
	LUT2 #(
		.INIT('h8)
	) name3364 (
		\g1319_reg/NET0131 ,
		_w2872_,
		_w4544_
	);
	LUT2 #(
		.INIT('h1)
	) name3365 (
		\g1332_reg/NET0131 ,
		_w2882_,
		_w4545_
	);
	LUT2 #(
		.INIT('h1)
	) name3366 (
		\g1358_reg/NET0131 ,
		_w2907_,
		_w4546_
	);
	LUT2 #(
		.INIT('h8)
	) name3367 (
		\g1346_reg/NET0131 ,
		_w2862_,
		_w4547_
	);
	LUT2 #(
		.INIT('h8)
	) name3368 (
		\g1358_reg/NET0131 ,
		_w2907_,
		_w4548_
	);
	LUT2 #(
		.INIT('h8)
	) name3369 (
		\g1339_reg/NET0131 ,
		_w2912_,
		_w4549_
	);
	LUT2 #(
		.INIT('h1)
	) name3370 (
		\g1326_reg/NET0131 ,
		_w2867_,
		_w4550_
	);
	LUT2 #(
		.INIT('h8)
	) name3371 (
		\g1365_reg/NET0131 ,
		_w2892_,
		_w4551_
	);
	LUT2 #(
		.INIT('h8)
	) name3372 (
		\g1332_reg/NET0131 ,
		_w2882_,
		_w4552_
	);
	LUT2 #(
		.INIT('h1)
	) name3373 (
		\g1319_reg/NET0131 ,
		_w2872_,
		_w4553_
	);
	LUT2 #(
		.INIT('h8)
	) name3374 (
		\g1378_reg/NET0131 ,
		_w2887_,
		_w4554_
	);
	LUT2 #(
		.INIT('h8)
	) name3375 (
		\g1352_reg/NET0131 ,
		_w2877_,
		_w4555_
	);
	LUT2 #(
		.INIT('h8)
	) name3376 (
		\g1326_reg/NET0131 ,
		_w2867_,
		_w4556_
	);
	LUT2 #(
		.INIT('h1)
	) name3377 (
		\g1378_reg/NET0131 ,
		_w2887_,
		_w4557_
	);
	LUT2 #(
		.INIT('h1)
	) name3378 (
		\g1352_reg/NET0131 ,
		_w2877_,
		_w4558_
	);
	LUT2 #(
		.INIT('h1)
	) name3379 (
		_w4539_,
		_w4540_,
		_w4559_
	);
	LUT2 #(
		.INIT('h1)
	) name3380 (
		_w4541_,
		_w4542_,
		_w4560_
	);
	LUT2 #(
		.INIT('h1)
	) name3381 (
		_w4543_,
		_w4544_,
		_w4561_
	);
	LUT2 #(
		.INIT('h1)
	) name3382 (
		_w4545_,
		_w4546_,
		_w4562_
	);
	LUT2 #(
		.INIT('h1)
	) name3383 (
		_w4547_,
		_w4548_,
		_w4563_
	);
	LUT2 #(
		.INIT('h1)
	) name3384 (
		_w4549_,
		_w4550_,
		_w4564_
	);
	LUT2 #(
		.INIT('h1)
	) name3385 (
		_w4551_,
		_w4552_,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w4553_,
		_w4554_,
		_w4566_
	);
	LUT2 #(
		.INIT('h1)
	) name3387 (
		_w4555_,
		_w4556_,
		_w4567_
	);
	LUT2 #(
		.INIT('h1)
	) name3388 (
		_w4557_,
		_w4558_,
		_w4568_
	);
	LUT2 #(
		.INIT('h8)
	) name3389 (
		_w4567_,
		_w4568_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name3390 (
		_w4565_,
		_w4566_,
		_w4570_
	);
	LUT2 #(
		.INIT('h8)
	) name3391 (
		_w4563_,
		_w4564_,
		_w4571_
	);
	LUT2 #(
		.INIT('h8)
	) name3392 (
		_w4561_,
		_w4562_,
		_w4572_
	);
	LUT2 #(
		.INIT('h8)
	) name3393 (
		_w4559_,
		_w4560_,
		_w4573_
	);
	LUT2 #(
		.INIT('h8)
	) name3394 (
		_w4572_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h8)
	) name3395 (
		_w4570_,
		_w4571_,
		_w4575_
	);
	LUT2 #(
		.INIT('h8)
	) name3396 (
		_w4569_,
		_w4575_,
		_w4576_
	);
	LUT2 #(
		.INIT('h8)
	) name3397 (
		_w4574_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w4536_,
		_w4537_,
		_w4578_
	);
	LUT2 #(
		.INIT('h4)
	) name3399 (
		_w4538_,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h8)
	) name3400 (
		_w2902_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h4)
	) name3401 (
		_w4577_,
		_w4580_,
		_w4581_
	);
	LUT2 #(
		.INIT('h8)
	) name3402 (
		_w4534_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name3403 (
		_w4535_,
		_w4582_,
		_w4583_
	);
	LUT2 #(
		.INIT('h8)
	) name3404 (
		\g1018_reg/NET0131 ,
		_w4533_,
		_w4584_
	);
	LUT2 #(
		.INIT('h2)
	) name3405 (
		\g1422_reg/NET0131 ,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h8)
	) name3406 (
		_w4581_,
		_w4584_,
		_w4586_
	);
	LUT2 #(
		.INIT('h1)
	) name3407 (
		_w4585_,
		_w4586_,
		_w4587_
	);
	LUT2 #(
		.INIT('h8)
	) name3408 (
		\g5657_pad ,
		_w4533_,
		_w4588_
	);
	LUT2 #(
		.INIT('h2)
	) name3409 (
		\g1421_reg/NET0131 ,
		_w4588_,
		_w4589_
	);
	LUT2 #(
		.INIT('h8)
	) name3410 (
		_w4581_,
		_w4588_,
		_w4590_
	);
	LUT2 #(
		.INIT('h1)
	) name3411 (
		_w4589_,
		_w4590_,
		_w4591_
	);
	LUT2 #(
		.INIT('h4)
	) name3412 (
		\g1345_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name3413 (
		\g1918_reg/NET0131 ,
		_w4592_,
		_w4593_
	);
	LUT2 #(
		.INIT('h8)
	) name3414 (
		\g1024_reg/NET0131 ,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		\g2114_reg/NET0131 ,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h2)
	) name3416 (
		\g1018_reg/NET0131 ,
		\g2110_reg/NET0131 ,
		_w4596_
	);
	LUT2 #(
		.INIT('h4)
	) name3417 (
		\g2109_reg/NET0131 ,
		\g5657_pad ,
		_w4597_
	);
	LUT2 #(
		.INIT('h2)
	) name3418 (
		\g1024_reg/NET0131 ,
		\g2108_reg/NET0131 ,
		_w4598_
	);
	LUT2 #(
		.INIT('h1)
	) name3419 (
		\g1339_reg/NET0131 ,
		_w1780_,
		_w4599_
	);
	LUT2 #(
		.INIT('h1)
	) name3420 (
		\g1378_reg/NET0131 ,
		_w1785_,
		_w4600_
	);
	LUT2 #(
		.INIT('h8)
	) name3421 (
		\g1378_reg/NET0131 ,
		_w1785_,
		_w4601_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		\g1372_reg/NET0131 ,
		_w1750_,
		_w4602_
	);
	LUT2 #(
		.INIT('h1)
	) name3423 (
		\g1346_reg/NET0131 ,
		_w1765_,
		_w4603_
	);
	LUT2 #(
		.INIT('h8)
	) name3424 (
		\g1319_reg/NET0131 ,
		_w1770_,
		_w4604_
	);
	LUT2 #(
		.INIT('h1)
	) name3425 (
		\g1358_reg/NET0131 ,
		_w1755_,
		_w4605_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		\g1332_reg/NET0131 ,
		_w1775_,
		_w4606_
	);
	LUT2 #(
		.INIT('h8)
	) name3427 (
		\g1346_reg/NET0131 ,
		_w1765_,
		_w4607_
	);
	LUT2 #(
		.INIT('h8)
	) name3428 (
		\g1332_reg/NET0131 ,
		_w1775_,
		_w4608_
	);
	LUT2 #(
		.INIT('h8)
	) name3429 (
		\g1339_reg/NET0131 ,
		_w1780_,
		_w4609_
	);
	LUT2 #(
		.INIT('h1)
	) name3430 (
		\g1326_reg/NET0131 ,
		_w1760_,
		_w4610_
	);
	LUT2 #(
		.INIT('h8)
	) name3431 (
		\g1372_reg/NET0131 ,
		_w1750_,
		_w4611_
	);
	LUT2 #(
		.INIT('h8)
	) name3432 (
		\g1358_reg/NET0131 ,
		_w1755_,
		_w4612_
	);
	LUT2 #(
		.INIT('h1)
	) name3433 (
		\g1319_reg/NET0131 ,
		_w1770_,
		_w4613_
	);
	LUT2 #(
		.INIT('h8)
	) name3434 (
		\g1352_reg/NET0131 ,
		_w1800_,
		_w4614_
	);
	LUT2 #(
		.INIT('h8)
	) name3435 (
		\g1365_reg/NET0131 ,
		_w1790_,
		_w4615_
	);
	LUT2 #(
		.INIT('h8)
	) name3436 (
		\g1326_reg/NET0131 ,
		_w1760_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name3437 (
		\g1352_reg/NET0131 ,
		_w1800_,
		_w4617_
	);
	LUT2 #(
		.INIT('h1)
	) name3438 (
		\g1365_reg/NET0131 ,
		_w1790_,
		_w4618_
	);
	LUT2 #(
		.INIT('h1)
	) name3439 (
		_w4599_,
		_w4600_,
		_w4619_
	);
	LUT2 #(
		.INIT('h1)
	) name3440 (
		_w4601_,
		_w4602_,
		_w4620_
	);
	LUT2 #(
		.INIT('h1)
	) name3441 (
		_w4603_,
		_w4604_,
		_w4621_
	);
	LUT2 #(
		.INIT('h1)
	) name3442 (
		_w4605_,
		_w4606_,
		_w4622_
	);
	LUT2 #(
		.INIT('h1)
	) name3443 (
		_w4607_,
		_w4608_,
		_w4623_
	);
	LUT2 #(
		.INIT('h1)
	) name3444 (
		_w4609_,
		_w4610_,
		_w4624_
	);
	LUT2 #(
		.INIT('h1)
	) name3445 (
		_w4611_,
		_w4612_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name3446 (
		_w4613_,
		_w4614_,
		_w4626_
	);
	LUT2 #(
		.INIT('h1)
	) name3447 (
		_w4615_,
		_w4616_,
		_w4627_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		_w4617_,
		_w4618_,
		_w4628_
	);
	LUT2 #(
		.INIT('h8)
	) name3449 (
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('h8)
	) name3450 (
		_w4625_,
		_w4626_,
		_w4630_
	);
	LUT2 #(
		.INIT('h8)
	) name3451 (
		_w4623_,
		_w4624_,
		_w4631_
	);
	LUT2 #(
		.INIT('h8)
	) name3452 (
		_w4621_,
		_w4622_,
		_w4632_
	);
	LUT2 #(
		.INIT('h8)
	) name3453 (
		_w4619_,
		_w4620_,
		_w4633_
	);
	LUT2 #(
		.INIT('h8)
	) name3454 (
		_w4632_,
		_w4633_,
		_w4634_
	);
	LUT2 #(
		.INIT('h8)
	) name3455 (
		_w4630_,
		_w4631_,
		_w4635_
	);
	LUT2 #(
		.INIT('h8)
	) name3456 (
		_w4629_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h8)
	) name3457 (
		_w4634_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		_w4596_,
		_w4597_,
		_w4638_
	);
	LUT2 #(
		.INIT('h4)
	) name3459 (
		_w4598_,
		_w4638_,
		_w4639_
	);
	LUT2 #(
		.INIT('h8)
	) name3460 (
		_w1795_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h4)
	) name3461 (
		_w4637_,
		_w4640_,
		_w4641_
	);
	LUT2 #(
		.INIT('h8)
	) name3462 (
		_w4594_,
		_w4641_,
		_w4642_
	);
	LUT2 #(
		.INIT('h1)
	) name3463 (
		_w4595_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h4)
	) name3464 (
		\g1345_reg/NET0131 ,
		\g525_reg/NET0131 ,
		_w4644_
	);
	LUT2 #(
		.INIT('h8)
	) name3465 (
		\g538_reg/NET0131 ,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h8)
	) name3466 (
		\g1024_reg/NET0131 ,
		_w4645_,
		_w4646_
	);
	LUT2 #(
		.INIT('h2)
	) name3467 (
		\g734_reg/NET0131 ,
		_w4646_,
		_w4647_
	);
	LUT2 #(
		.INIT('h2)
	) name3468 (
		\g1018_reg/NET0131 ,
		\g730_reg/NET0131 ,
		_w4648_
	);
	LUT2 #(
		.INIT('h2)
	) name3469 (
		\g5657_pad ,
		\g729_reg/NET0131 ,
		_w4649_
	);
	LUT2 #(
		.INIT('h2)
	) name3470 (
		\g1024_reg/NET0131 ,
		\g728_reg/NET0131 ,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name3471 (
		\g1339_reg/NET0131 ,
		_w3718_,
		_w4651_
	);
	LUT2 #(
		.INIT('h1)
	) name3472 (
		\g1378_reg/NET0131 ,
		_w3678_,
		_w4652_
	);
	LUT2 #(
		.INIT('h8)
	) name3473 (
		\g1378_reg/NET0131 ,
		_w3678_,
		_w4653_
	);
	LUT2 #(
		.INIT('h1)
	) name3474 (
		\g1372_reg/NET0131 ,
		_w3698_,
		_w4654_
	);
	LUT2 #(
		.INIT('h1)
	) name3475 (
		\g1326_reg/NET0131 ,
		_w3708_,
		_w4655_
	);
	LUT2 #(
		.INIT('h8)
	) name3476 (
		\g1319_reg/NET0131 ,
		_w3703_,
		_w4656_
	);
	LUT2 #(
		.INIT('h1)
	) name3477 (
		\g1358_reg/NET0131 ,
		_w3723_,
		_w4657_
	);
	LUT2 #(
		.INIT('h1)
	) name3478 (
		\g1352_reg/NET0131 ,
		_w3693_,
		_w4658_
	);
	LUT2 #(
		.INIT('h8)
	) name3479 (
		\g1326_reg/NET0131 ,
		_w3708_,
		_w4659_
	);
	LUT2 #(
		.INIT('h8)
	) name3480 (
		\g1352_reg/NET0131 ,
		_w3693_,
		_w4660_
	);
	LUT2 #(
		.INIT('h8)
	) name3481 (
		\g1339_reg/NET0131 ,
		_w3718_,
		_w4661_
	);
	LUT2 #(
		.INIT('h1)
	) name3482 (
		\g1346_reg/NET0131 ,
		_w3688_,
		_w4662_
	);
	LUT2 #(
		.INIT('h8)
	) name3483 (
		\g1372_reg/NET0131 ,
		_w3698_,
		_w4663_
	);
	LUT2 #(
		.INIT('h8)
	) name3484 (
		\g1358_reg/NET0131 ,
		_w3723_,
		_w4664_
	);
	LUT2 #(
		.INIT('h1)
	) name3485 (
		\g1319_reg/NET0131 ,
		_w3703_,
		_w4665_
	);
	LUT2 #(
		.INIT('h8)
	) name3486 (
		\g1332_reg/NET0131 ,
		_w3713_,
		_w4666_
	);
	LUT2 #(
		.INIT('h8)
	) name3487 (
		\g1365_reg/NET0131 ,
		_w3733_,
		_w4667_
	);
	LUT2 #(
		.INIT('h8)
	) name3488 (
		\g1346_reg/NET0131 ,
		_w3688_,
		_w4668_
	);
	LUT2 #(
		.INIT('h1)
	) name3489 (
		\g1332_reg/NET0131 ,
		_w3713_,
		_w4669_
	);
	LUT2 #(
		.INIT('h1)
	) name3490 (
		\g1365_reg/NET0131 ,
		_w3733_,
		_w4670_
	);
	LUT2 #(
		.INIT('h1)
	) name3491 (
		_w4651_,
		_w4652_,
		_w4671_
	);
	LUT2 #(
		.INIT('h1)
	) name3492 (
		_w4653_,
		_w4654_,
		_w4672_
	);
	LUT2 #(
		.INIT('h1)
	) name3493 (
		_w4655_,
		_w4656_,
		_w4673_
	);
	LUT2 #(
		.INIT('h1)
	) name3494 (
		_w4657_,
		_w4658_,
		_w4674_
	);
	LUT2 #(
		.INIT('h1)
	) name3495 (
		_w4659_,
		_w4660_,
		_w4675_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		_w4661_,
		_w4662_,
		_w4676_
	);
	LUT2 #(
		.INIT('h1)
	) name3497 (
		_w4663_,
		_w4664_,
		_w4677_
	);
	LUT2 #(
		.INIT('h1)
	) name3498 (
		_w4665_,
		_w4666_,
		_w4678_
	);
	LUT2 #(
		.INIT('h1)
	) name3499 (
		_w4667_,
		_w4668_,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name3500 (
		_w4669_,
		_w4670_,
		_w4680_
	);
	LUT2 #(
		.INIT('h8)
	) name3501 (
		_w4679_,
		_w4680_,
		_w4681_
	);
	LUT2 #(
		.INIT('h8)
	) name3502 (
		_w4677_,
		_w4678_,
		_w4682_
	);
	LUT2 #(
		.INIT('h8)
	) name3503 (
		_w4675_,
		_w4676_,
		_w4683_
	);
	LUT2 #(
		.INIT('h8)
	) name3504 (
		_w4673_,
		_w4674_,
		_w4684_
	);
	LUT2 #(
		.INIT('h8)
	) name3505 (
		_w4671_,
		_w4672_,
		_w4685_
	);
	LUT2 #(
		.INIT('h8)
	) name3506 (
		_w4684_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('h8)
	) name3507 (
		_w4682_,
		_w4683_,
		_w4687_
	);
	LUT2 #(
		.INIT('h8)
	) name3508 (
		_w4681_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h8)
	) name3509 (
		_w4686_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h1)
	) name3510 (
		_w4648_,
		_w4649_,
		_w4690_
	);
	LUT2 #(
		.INIT('h4)
	) name3511 (
		_w4650_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h8)
	) name3512 (
		_w3683_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h4)
	) name3513 (
		_w4689_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h8)
	) name3514 (
		_w4646_,
		_w4693_,
		_w4694_
	);
	LUT2 #(
		.INIT('h1)
	) name3515 (
		_w4647_,
		_w4694_,
		_w4695_
	);
	LUT2 #(
		.INIT('h8)
	) name3516 (
		\g5657_pad ,
		_w4645_,
		_w4696_
	);
	LUT2 #(
		.INIT('h2)
	) name3517 (
		\g735_reg/NET0131 ,
		_w4696_,
		_w4697_
	);
	LUT2 #(
		.INIT('h8)
	) name3518 (
		_w4693_,
		_w4696_,
		_w4698_
	);
	LUT2 #(
		.INIT('h1)
	) name3519 (
		_w4697_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h8)
	) name3520 (
		\g1018_reg/NET0131 ,
		_w4645_,
		_w4700_
	);
	LUT2 #(
		.INIT('h2)
	) name3521 (
		\g736_reg/NET0131 ,
		_w4700_,
		_w4701_
	);
	LUT2 #(
		.INIT('h8)
	) name3522 (
		_w4693_,
		_w4700_,
		_w4702_
	);
	LUT2 #(
		.INIT('h1)
	) name3523 (
		_w4701_,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		\g1018_reg/NET0131 ,
		_w4593_,
		_w4704_
	);
	LUT2 #(
		.INIT('h2)
	) name3525 (
		\g2116_reg/NET0131 ,
		_w4704_,
		_w4705_
	);
	LUT2 #(
		.INIT('h8)
	) name3526 (
		_w4641_,
		_w4704_,
		_w4706_
	);
	LUT2 #(
		.INIT('h1)
	) name3527 (
		_w4705_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h8)
	) name3528 (
		\g5657_pad ,
		_w4593_,
		_w4708_
	);
	LUT2 #(
		.INIT('h2)
	) name3529 (
		\g2115_reg/NET0131 ,
		_w4708_,
		_w4709_
	);
	LUT2 #(
		.INIT('h8)
	) name3530 (
		_w4641_,
		_w4708_,
		_w4710_
	);
	LUT2 #(
		.INIT('h1)
	) name3531 (
		_w4709_,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h8)
	) name3532 (
		\g1024_reg/NET0131 ,
		_w4477_,
		_w4712_
	);
	LUT2 #(
		.INIT('h2)
	) name3533 (
		\g2808_reg/NET0131 ,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h8)
	) name3534 (
		_w4525_,
		_w4712_,
		_w4714_
	);
	LUT2 #(
		.INIT('h1)
	) name3535 (
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT2 #(
		.INIT('h1)
	) name3536 (
		_w1745_,
		_w4136_,
		_w4716_
	);
	LUT2 #(
		.INIT('h8)
	) name3537 (
		\g1760_reg/NET0131 ,
		\g5657_pad ,
		_w4717_
	);
	LUT2 #(
		.INIT('h8)
	) name3538 (
		\g1024_reg/NET0131 ,
		\g1764_reg/NET0131 ,
		_w4718_
	);
	LUT2 #(
		.INIT('h8)
	) name3539 (
		\g1018_reg/NET0131 ,
		\g1762_reg/NET0131 ,
		_w4719_
	);
	LUT2 #(
		.INIT('h1)
	) name3540 (
		_w4717_,
		_w4718_,
		_w4720_
	);
	LUT2 #(
		.INIT('h4)
	) name3541 (
		_w4719_,
		_w4720_,
		_w4721_
	);
	LUT2 #(
		.INIT('h8)
	) name3542 (
		\g1730_reg/NET0131 ,
		\g5657_pad ,
		_w4722_
	);
	LUT2 #(
		.INIT('h8)
	) name3543 (
		\g1024_reg/NET0131 ,
		\g1734_reg/NET0131 ,
		_w4723_
	);
	LUT2 #(
		.INIT('h8)
	) name3544 (
		\g1018_reg/NET0131 ,
		\g1732_reg/NET0131 ,
		_w4724_
	);
	LUT2 #(
		.INIT('h1)
	) name3545 (
		_w4722_,
		_w4723_,
		_w4725_
	);
	LUT2 #(
		.INIT('h4)
	) name3546 (
		_w4724_,
		_w4725_,
		_w4726_
	);
	LUT2 #(
		.INIT('h8)
	) name3547 (
		_w4721_,
		_w4726_,
		_w4727_
	);
	LUT2 #(
		.INIT('h2)
	) name3548 (
		\g1018_reg/NET0131 ,
		\g1960_reg/NET0131 ,
		_w4728_
	);
	LUT2 #(
		.INIT('h2)
	) name3549 (
		\g1024_reg/NET0131 ,
		\g1958_reg/NET0131 ,
		_w4729_
	);
	LUT2 #(
		.INIT('h4)
	) name3550 (
		\g1959_reg/NET0131 ,
		\g5657_pad ,
		_w4730_
	);
	LUT2 #(
		.INIT('h1)
	) name3551 (
		_w4728_,
		_w4729_,
		_w4731_
	);
	LUT2 #(
		.INIT('h4)
	) name3552 (
		_w4730_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h2)
	) name3553 (
		\g1018_reg/NET0131 ,
		\g1957_reg/NET0131 ,
		_w4733_
	);
	LUT2 #(
		.INIT('h2)
	) name3554 (
		\g1024_reg/NET0131 ,
		\g1955_reg/NET0131 ,
		_w4734_
	);
	LUT2 #(
		.INIT('h4)
	) name3555 (
		\g1956_reg/NET0131 ,
		\g5657_pad ,
		_w4735_
	);
	LUT2 #(
		.INIT('h1)
	) name3556 (
		_w4733_,
		_w4734_,
		_w4736_
	);
	LUT2 #(
		.INIT('h4)
	) name3557 (
		_w4735_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h1)
	) name3558 (
		_w4732_,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h8)
	) name3559 (
		_w4727_,
		_w4738_,
		_w4739_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		\g1745_reg/NET0131 ,
		\g5657_pad ,
		_w4740_
	);
	LUT2 #(
		.INIT('h8)
	) name3561 (
		\g1024_reg/NET0131 ,
		\g1749_reg/NET0131 ,
		_w4741_
	);
	LUT2 #(
		.INIT('h8)
	) name3562 (
		\g1018_reg/NET0131 ,
		\g1747_reg/NET0131 ,
		_w4742_
	);
	LUT2 #(
		.INIT('h1)
	) name3563 (
		_w4740_,
		_w4741_,
		_w4743_
	);
	LUT2 #(
		.INIT('h4)
	) name3564 (
		_w4742_,
		_w4743_,
		_w4744_
	);
	LUT2 #(
		.INIT('h2)
	) name3565 (
		\g1018_reg/NET0131 ,
		\g1963_reg/NET0131 ,
		_w4745_
	);
	LUT2 #(
		.INIT('h4)
	) name3566 (
		\g1962_reg/NET0131 ,
		\g5657_pad ,
		_w4746_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		\g1024_reg/NET0131 ,
		\g1961_reg/NET0131 ,
		_w4747_
	);
	LUT2 #(
		.INIT('h1)
	) name3568 (
		_w4745_,
		_w4746_,
		_w4748_
	);
	LUT2 #(
		.INIT('h4)
	) name3569 (
		_w4747_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h2)
	) name3570 (
		_w4737_,
		_w4749_,
		_w4750_
	);
	LUT2 #(
		.INIT('h1)
	) name3571 (
		_w4726_,
		_w4750_,
		_w4751_
	);
	LUT2 #(
		.INIT('h4)
	) name3572 (
		_w4732_,
		_w4749_,
		_w4752_
	);
	LUT2 #(
		.INIT('h2)
	) name3573 (
		_w4726_,
		_w4752_,
		_w4753_
	);
	LUT2 #(
		.INIT('h2)
	) name3574 (
		_w4744_,
		_w4751_,
		_w4754_
	);
	LUT2 #(
		.INIT('h4)
	) name3575 (
		_w4753_,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h2)
	) name3576 (
		\g1018_reg/NET0131 ,
		\g1966_reg/NET0131 ,
		_w4756_
	);
	LUT2 #(
		.INIT('h4)
	) name3577 (
		\g1965_reg/NET0131 ,
		\g5657_pad ,
		_w4757_
	);
	LUT2 #(
		.INIT('h2)
	) name3578 (
		\g1024_reg/NET0131 ,
		\g1964_reg/NET0131 ,
		_w4758_
	);
	LUT2 #(
		.INIT('h1)
	) name3579 (
		_w4756_,
		_w4757_,
		_w4759_
	);
	LUT2 #(
		.INIT('h4)
	) name3580 (
		_w4758_,
		_w4759_,
		_w4760_
	);
	LUT2 #(
		.INIT('h1)
	) name3581 (
		_w4726_,
		_w4760_,
		_w4761_
	);
	LUT2 #(
		.INIT('h1)
	) name3582 (
		_w4744_,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h4)
	) name3583 (
		_w4732_,
		_w4737_,
		_w4763_
	);
	LUT2 #(
		.INIT('h2)
	) name3584 (
		_w4744_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h1)
	) name3585 (
		_w4721_,
		_w4762_,
		_w4765_
	);
	LUT2 #(
		.INIT('h4)
	) name3586 (
		_w4764_,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h8)
	) name3587 (
		_w4732_,
		_w4749_,
		_w4767_
	);
	LUT2 #(
		.INIT('h1)
	) name3588 (
		_w4726_,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('h8)
	) name3589 (
		\g1775_reg/NET0131 ,
		\g5657_pad ,
		_w4769_
	);
	LUT2 #(
		.INIT('h8)
	) name3590 (
		\g1024_reg/NET0131 ,
		\g1705_reg/NET0131 ,
		_w4770_
	);
	LUT2 #(
		.INIT('h8)
	) name3591 (
		\g1018_reg/NET0131 ,
		\g1777_reg/NET0131 ,
		_w4771_
	);
	LUT2 #(
		.INIT('h1)
	) name3592 (
		_w4769_,
		_w4770_,
		_w4772_
	);
	LUT2 #(
		.INIT('h4)
	) name3593 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h1)
	) name3594 (
		_w4744_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h4)
	) name3595 (
		_w4726_,
		_w4737_,
		_w4775_
	);
	LUT2 #(
		.INIT('h1)
	) name3596 (
		_w4737_,
		_w4749_,
		_w4776_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w4775_,
		_w4776_,
		_w4777_
	);
	LUT2 #(
		.INIT('h4)
	) name3598 (
		_w4768_,
		_w4774_,
		_w4778_
	);
	LUT2 #(
		.INIT('h4)
	) name3599 (
		_w4777_,
		_w4778_,
		_w4779_
	);
	LUT2 #(
		.INIT('h2)
	) name3600 (
		_w4721_,
		_w4726_,
		_w4780_
	);
	LUT2 #(
		.INIT('h8)
	) name3601 (
		_w4732_,
		_w4737_,
		_w4781_
	);
	LUT2 #(
		.INIT('h8)
	) name3602 (
		_w4760_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('h8)
	) name3603 (
		_w4780_,
		_w4782_,
		_w4783_
	);
	LUT2 #(
		.INIT('h4)
	) name3604 (
		_w4721_,
		_w4726_,
		_w4784_
	);
	LUT2 #(
		.INIT('h4)
	) name3605 (
		_w4744_,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h2)
	) name3606 (
		_w4732_,
		_w4737_,
		_w4786_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		_w4760_,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('h8)
	) name3608 (
		_w4785_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h8)
	) name3609 (
		_w4749_,
		_w4773_,
		_w4789_
	);
	LUT2 #(
		.INIT('h8)
	) name3610 (
		_w4786_,
		_w4789_,
		_w4790_
	);
	LUT2 #(
		.INIT('h1)
	) name3611 (
		_w4739_,
		_w4790_,
		_w4791_
	);
	LUT2 #(
		.INIT('h4)
	) name3612 (
		_w4783_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h4)
	) name3613 (
		_w4788_,
		_w4792_,
		_w4793_
	);
	LUT2 #(
		.INIT('h1)
	) name3614 (
		_w4755_,
		_w4766_,
		_w4794_
	);
	LUT2 #(
		.INIT('h4)
	) name3615 (
		_w4779_,
		_w4794_,
		_w4795_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		_w4793_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h8)
	) name3617 (
		_w4781_,
		_w4785_,
		_w4797_
	);
	LUT2 #(
		.INIT('h1)
	) name3618 (
		_w4727_,
		_w4749_,
		_w4798_
	);
	LUT2 #(
		.INIT('h1)
	) name3619 (
		_w4721_,
		_w4726_,
		_w4799_
	);
	LUT2 #(
		.INIT('h8)
	) name3620 (
		_w4760_,
		_w4799_,
		_w4800_
	);
	LUT2 #(
		.INIT('h1)
	) name3621 (
		_w4798_,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h2)
	) name3622 (
		_w4744_,
		_w4801_,
		_w4802_
	);
	LUT2 #(
		.INIT('h2)
	) name3623 (
		_w4726_,
		_w4760_,
		_w4803_
	);
	LUT2 #(
		.INIT('h4)
	) name3624 (
		_w4773_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h1)
	) name3625 (
		_w4802_,
		_w4804_,
		_w4805_
	);
	LUT2 #(
		.INIT('h1)
	) name3626 (
		_w4737_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h8)
	) name3627 (
		_w4750_,
		_w4799_,
		_w4807_
	);
	LUT2 #(
		.INIT('h8)
	) name3628 (
		_w4727_,
		_w4767_,
		_w4808_
	);
	LUT2 #(
		.INIT('h4)
	) name3629 (
		_w4732_,
		_w4780_,
		_w4809_
	);
	LUT2 #(
		.INIT('h1)
	) name3630 (
		_w4807_,
		_w4808_,
		_w4810_
	);
	LUT2 #(
		.INIT('h4)
	) name3631 (
		_w4809_,
		_w4810_,
		_w4811_
	);
	LUT2 #(
		.INIT('h1)
	) name3632 (
		_w4744_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h8)
	) name3633 (
		_w4760_,
		_w4775_,
		_w4813_
	);
	LUT2 #(
		.INIT('h1)
	) name3634 (
		_w4750_,
		_w4813_,
		_w4814_
	);
	LUT2 #(
		.INIT('h2)
	) name3635 (
		_w4773_,
		_w4814_,
		_w4815_
	);
	LUT2 #(
		.INIT('h2)
	) name3636 (
		_w4721_,
		_w4760_,
		_w4816_
	);
	LUT2 #(
		.INIT('h8)
	) name3637 (
		_w4744_,
		_w4786_,
		_w4817_
	);
	LUT2 #(
		.INIT('h1)
	) name3638 (
		_w4816_,
		_w4817_,
		_w4818_
	);
	LUT2 #(
		.INIT('h2)
	) name3639 (
		_w4726_,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h1)
	) name3640 (
		_w4721_,
		_w4774_,
		_w4820_
	);
	LUT2 #(
		.INIT('h4)
	) name3641 (
		_w4726_,
		_w4752_,
		_w4821_
	);
	LUT2 #(
		.INIT('h4)
	) name3642 (
		_w4820_,
		_w4821_,
		_w4822_
	);
	LUT2 #(
		.INIT('h1)
	) name3643 (
		_w4797_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h4)
	) name3644 (
		_w4815_,
		_w4823_,
		_w4824_
	);
	LUT2 #(
		.INIT('h4)
	) name3645 (
		_w4819_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h4)
	) name3646 (
		_w4812_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h4)
	) name3647 (
		_w4806_,
		_w4826_,
		_w4827_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		\g1976_reg/NET0131 ,
		\g5657_pad ,
		_w4828_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		\g1024_reg/NET0131 ,
		\g1982_reg/NET0131 ,
		_w4829_
	);
	LUT2 #(
		.INIT('h8)
	) name3650 (
		\g1018_reg/NET0131 ,
		\g1979_reg/NET0131 ,
		_w4830_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		\g1945_reg/NET0131 ,
		\g5657_pad ,
		_w4831_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		\g1024_reg/NET0131 ,
		\g1870_reg/NET0131 ,
		_w4832_
	);
	LUT2 #(
		.INIT('h8)
	) name3653 (
		\g1018_reg/NET0131 ,
		\g1947_reg/NET0131 ,
		_w4833_
	);
	LUT2 #(
		.INIT('h1)
	) name3654 (
		_w4831_,
		_w4832_,
		_w4834_
	);
	LUT2 #(
		.INIT('h4)
	) name3655 (
		_w4833_,
		_w4834_,
		_w4835_
	);
	LUT2 #(
		.INIT('h8)
	) name3656 (
		\g185_reg/NET0131 ,
		\g1922_reg/NET0131 ,
		_w4836_
	);
	LUT2 #(
		.INIT('h4)
	) name3657 (
		_w4835_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h1)
	) name3658 (
		_w4828_,
		_w4829_,
		_w4838_
	);
	LUT2 #(
		.INIT('h4)
	) name3659 (
		_w4830_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h4)
	) name3660 (
		_w4837_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h8)
	) name3661 (
		_w4827_,
		_w4840_,
		_w4841_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		\g1967_reg/NET0131 ,
		\g5657_pad ,
		_w4842_
	);
	LUT2 #(
		.INIT('h8)
	) name3663 (
		\g1018_reg/NET0131 ,
		\g1970_reg/NET0131 ,
		_w4843_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		\g1024_reg/NET0131 ,
		\g1973_reg/NET0131 ,
		_w4844_
	);
	LUT2 #(
		.INIT('h8)
	) name3665 (
		\g1018_reg/NET0131 ,
		\g1951_reg/NET0131 ,
		_w4845_
	);
	LUT2 #(
		.INIT('h8)
	) name3666 (
		\g1024_reg/NET0131 ,
		\g1953_reg/NET0131 ,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name3667 (
		\g1949_reg/NET0131 ,
		\g5657_pad ,
		_w4847_
	);
	LUT2 #(
		.INIT('h1)
	) name3668 (
		_w4845_,
		_w4846_,
		_w4848_
	);
	LUT2 #(
		.INIT('h4)
	) name3669 (
		_w4847_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h8)
	) name3670 (
		\g185_reg/NET0131 ,
		\g1904_reg/NET0131 ,
		_w4850_
	);
	LUT2 #(
		.INIT('h4)
	) name3671 (
		_w4849_,
		_w4850_,
		_w4851_
	);
	LUT2 #(
		.INIT('h1)
	) name3672 (
		_w4842_,
		_w4843_,
		_w4852_
	);
	LUT2 #(
		.INIT('h4)
	) name3673 (
		_w4844_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h4)
	) name3674 (
		_w4851_,
		_w4853_,
		_w4854_
	);
	LUT2 #(
		.INIT('h1)
	) name3675 (
		_w4840_,
		_w4854_,
		_w4855_
	);
	LUT2 #(
		.INIT('h2)
	) name3676 (
		_w4136_,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h8)
	) name3677 (
		_w4796_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('h4)
	) name3678 (
		_w4841_,
		_w4857_,
		_w4858_
	);
	LUT2 #(
		.INIT('h1)
	) name3679 (
		_w4716_,
		_w4858_,
		_w4859_
	);
	LUT2 #(
		.INIT('h1)
	) name3680 (
		_w3754_,
		_w4136_,
		_w4860_
	);
	LUT2 #(
		.INIT('h8)
	) name3681 (
		\g364_reg/NET0131 ,
		\g5657_pad ,
		_w4861_
	);
	LUT2 #(
		.INIT('h8)
	) name3682 (
		\g1024_reg/NET0131 ,
		\g368_reg/NET0131 ,
		_w4862_
	);
	LUT2 #(
		.INIT('h8)
	) name3683 (
		\g1018_reg/NET0131 ,
		\g366_reg/NET0131 ,
		_w4863_
	);
	LUT2 #(
		.INIT('h1)
	) name3684 (
		_w4861_,
		_w4862_,
		_w4864_
	);
	LUT2 #(
		.INIT('h4)
	) name3685 (
		_w4863_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('h8)
	) name3686 (
		\g379_reg/NET0131 ,
		\g5657_pad ,
		_w4866_
	);
	LUT2 #(
		.INIT('h8)
	) name3687 (
		\g1024_reg/NET0131 ,
		\g383_reg/NET0131 ,
		_w4867_
	);
	LUT2 #(
		.INIT('h8)
	) name3688 (
		\g1018_reg/NET0131 ,
		\g381_reg/NET0131 ,
		_w4868_
	);
	LUT2 #(
		.INIT('h1)
	) name3689 (
		_w4866_,
		_w4867_,
		_w4869_
	);
	LUT2 #(
		.INIT('h4)
	) name3690 (
		_w4868_,
		_w4869_,
		_w4870_
	);
	LUT2 #(
		.INIT('h2)
	) name3691 (
		_w4865_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		\g1018_reg/NET0131 ,
		\g580_reg/NET0131 ,
		_w4872_
	);
	LUT2 #(
		.INIT('h2)
	) name3693 (
		\g5657_pad ,
		\g579_reg/NET0131 ,
		_w4873_
	);
	LUT2 #(
		.INIT('h2)
	) name3694 (
		\g1024_reg/NET0131 ,
		\g578_reg/NET0131 ,
		_w4874_
	);
	LUT2 #(
		.INIT('h1)
	) name3695 (
		_w4872_,
		_w4873_,
		_w4875_
	);
	LUT2 #(
		.INIT('h4)
	) name3696 (
		_w4874_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h2)
	) name3697 (
		\g1024_reg/NET0131 ,
		\g575_reg/NET0131 ,
		_w4877_
	);
	LUT2 #(
		.INIT('h2)
	) name3698 (
		\g1018_reg/NET0131 ,
		\g577_reg/NET0131 ,
		_w4878_
	);
	LUT2 #(
		.INIT('h2)
	) name3699 (
		\g5657_pad ,
		\g576_reg/NET0131 ,
		_w4879_
	);
	LUT2 #(
		.INIT('h1)
	) name3700 (
		_w4877_,
		_w4878_,
		_w4880_
	);
	LUT2 #(
		.INIT('h4)
	) name3701 (
		_w4879_,
		_w4880_,
		_w4881_
	);
	LUT2 #(
		.INIT('h4)
	) name3702 (
		_w4876_,
		_w4881_,
		_w4882_
	);
	LUT2 #(
		.INIT('h8)
	) name3703 (
		_w4871_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h8)
	) name3704 (
		\g349_reg/NET0131 ,
		\g5657_pad ,
		_w4884_
	);
	LUT2 #(
		.INIT('h8)
	) name3705 (
		\g1024_reg/NET0131 ,
		\g353_reg/NET0131 ,
		_w4885_
	);
	LUT2 #(
		.INIT('h8)
	) name3706 (
		\g1018_reg/NET0131 ,
		\g351_reg/NET0131 ,
		_w4886_
	);
	LUT2 #(
		.INIT('h1)
	) name3707 (
		_w4884_,
		_w4885_,
		_w4887_
	);
	LUT2 #(
		.INIT('h4)
	) name3708 (
		_w4886_,
		_w4887_,
		_w4888_
	);
	LUT2 #(
		.INIT('h1)
	) name3709 (
		_w4876_,
		_w4881_,
		_w4889_
	);
	LUT2 #(
		.INIT('h8)
	) name3710 (
		_w4870_,
		_w4888_,
		_w4890_
	);
	LUT2 #(
		.INIT('h8)
	) name3711 (
		_w4889_,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h2)
	) name3712 (
		_w4870_,
		_w4888_,
		_w4892_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		_w4876_,
		_w4881_,
		_w4893_
	);
	LUT2 #(
		.INIT('h2)
	) name3714 (
		\g1018_reg/NET0131 ,
		\g586_reg/NET0131 ,
		_w4894_
	);
	LUT2 #(
		.INIT('h2)
	) name3715 (
		\g1024_reg/NET0131 ,
		\g584_reg/NET0131 ,
		_w4895_
	);
	LUT2 #(
		.INIT('h2)
	) name3716 (
		\g5657_pad ,
		\g585_reg/NET0131 ,
		_w4896_
	);
	LUT2 #(
		.INIT('h1)
	) name3717 (
		_w4894_,
		_w4895_,
		_w4897_
	);
	LUT2 #(
		.INIT('h4)
	) name3718 (
		_w4896_,
		_w4897_,
		_w4898_
	);
	LUT2 #(
		.INIT('h8)
	) name3719 (
		_w4893_,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		_w4892_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h1)
	) name3721 (
		_w4865_,
		_w4888_,
		_w4901_
	);
	LUT2 #(
		.INIT('h4)
	) name3722 (
		_w4870_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('h4)
	) name3723 (
		_w4898_,
		_w4902_,
		_w4903_
	);
	LUT2 #(
		.INIT('h4)
	) name3724 (
		_w4865_,
		_w4888_,
		_w4904_
	);
	LUT2 #(
		.INIT('h4)
	) name3725 (
		_w4870_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h2)
	) name3726 (
		_w4876_,
		_w4881_,
		_w4906_
	);
	LUT2 #(
		.INIT('h8)
	) name3727 (
		_w4898_,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		_w4905_,
		_w4907_,
		_w4908_
	);
	LUT2 #(
		.INIT('h8)
	) name3729 (
		\g394_reg/NET0131 ,
		\g5657_pad ,
		_w4909_
	);
	LUT2 #(
		.INIT('h8)
	) name3730 (
		\g1024_reg/NET0131 ,
		\g324_reg/NET0131 ,
		_w4910_
	);
	LUT2 #(
		.INIT('h8)
	) name3731 (
		\g1018_reg/NET0131 ,
		\g396_reg/NET0131 ,
		_w4911_
	);
	LUT2 #(
		.INIT('h1)
	) name3732 (
		_w4909_,
		_w4910_,
		_w4912_
	);
	LUT2 #(
		.INIT('h4)
	) name3733 (
		_w4911_,
		_w4912_,
		_w4913_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\g1018_reg/NET0131 ,
		\g583_reg/NET0131 ,
		_w4914_
	);
	LUT2 #(
		.INIT('h2)
	) name3735 (
		\g5657_pad ,
		\g582_reg/NET0131 ,
		_w4915_
	);
	LUT2 #(
		.INIT('h2)
	) name3736 (
		\g1024_reg/NET0131 ,
		\g581_reg/NET0131 ,
		_w4916_
	);
	LUT2 #(
		.INIT('h1)
	) name3737 (
		_w4914_,
		_w4915_,
		_w4917_
	);
	LUT2 #(
		.INIT('h4)
	) name3738 (
		_w4916_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h1)
	) name3739 (
		_w4881_,
		_w4918_,
		_w4919_
	);
	LUT2 #(
		.INIT('h2)
	) name3740 (
		_w4904_,
		_w4913_,
		_w4920_
	);
	LUT2 #(
		.INIT('h8)
	) name3741 (
		_w4919_,
		_w4920_,
		_w4921_
	);
	LUT2 #(
		.INIT('h2)
	) name3742 (
		_w4881_,
		_w4918_,
		_w4922_
	);
	LUT2 #(
		.INIT('h2)
	) name3743 (
		_w4865_,
		_w4888_,
		_w4923_
	);
	LUT2 #(
		.INIT('h8)
	) name3744 (
		_w4922_,
		_w4923_,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name3745 (
		_w4865_,
		_w4888_,
		_w4925_
	);
	LUT2 #(
		.INIT('h4)
	) name3746 (
		_w4876_,
		_w4925_,
		_w4926_
	);
	LUT2 #(
		.INIT('h2)
	) name3747 (
		_w4901_,
		_w4913_,
		_w4927_
	);
	LUT2 #(
		.INIT('h8)
	) name3748 (
		_w4893_,
		_w4927_,
		_w4928_
	);
	LUT2 #(
		.INIT('h8)
	) name3749 (
		_w4906_,
		_w4913_,
		_w4929_
	);
	LUT2 #(
		.INIT('h1)
	) name3750 (
		_w4926_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h4)
	) name3751 (
		_w4928_,
		_w4930_,
		_w4931_
	);
	LUT2 #(
		.INIT('h2)
	) name3752 (
		_w4918_,
		_w4931_,
		_w4932_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w4883_,
		_w4891_,
		_w4933_
	);
	LUT2 #(
		.INIT('h4)
	) name3754 (
		_w4924_,
		_w4933_,
		_w4934_
	);
	LUT2 #(
		.INIT('h1)
	) name3755 (
		_w4900_,
		_w4903_,
		_w4935_
	);
	LUT2 #(
		.INIT('h1)
	) name3756 (
		_w4908_,
		_w4921_,
		_w4936_
	);
	LUT2 #(
		.INIT('h8)
	) name3757 (
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('h8)
	) name3758 (
		_w4934_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h4)
	) name3759 (
		_w4932_,
		_w4938_,
		_w4939_
	);
	LUT2 #(
		.INIT('h8)
	) name3760 (
		\g5657_pad ,
		\g596_reg/NET0131 ,
		_w4940_
	);
	LUT2 #(
		.INIT('h8)
	) name3761 (
		\g1018_reg/NET0131 ,
		\g599_reg/NET0131 ,
		_w4941_
	);
	LUT2 #(
		.INIT('h8)
	) name3762 (
		\g1024_reg/NET0131 ,
		\g602_reg/NET0131 ,
		_w4942_
	);
	LUT2 #(
		.INIT('h8)
	) name3763 (
		\g5657_pad ,
		\g565_reg/NET0131 ,
		_w4943_
	);
	LUT2 #(
		.INIT('h8)
	) name3764 (
		\g1024_reg/NET0131 ,
		\g489_reg/NET0131 ,
		_w4944_
	);
	LUT2 #(
		.INIT('h8)
	) name3765 (
		\g1018_reg/NET0131 ,
		\g567_reg/NET0131 ,
		_w4945_
	);
	LUT2 #(
		.INIT('h1)
	) name3766 (
		_w4943_,
		_w4944_,
		_w4946_
	);
	LUT2 #(
		.INIT('h4)
	) name3767 (
		_w4945_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h8)
	) name3768 (
		\g185_reg/NET0131 ,
		\g542_reg/NET0131 ,
		_w4948_
	);
	LUT2 #(
		.INIT('h4)
	) name3769 (
		_w4947_,
		_w4948_,
		_w4949_
	);
	LUT2 #(
		.INIT('h1)
	) name3770 (
		_w4940_,
		_w4941_,
		_w4950_
	);
	LUT2 #(
		.INIT('h4)
	) name3771 (
		_w4942_,
		_w4950_,
		_w4951_
	);
	LUT2 #(
		.INIT('h4)
	) name3772 (
		_w4949_,
		_w4951_,
		_w4952_
	);
	LUT2 #(
		.INIT('h4)
	) name3773 (
		_w4876_,
		_w4918_,
		_w4953_
	);
	LUT2 #(
		.INIT('h1)
	) name3774 (
		_w4892_,
		_w4927_,
		_w4954_
	);
	LUT2 #(
		.INIT('h2)
	) name3775 (
		_w4953_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h8)
	) name3776 (
		_w4893_,
		_w4905_,
		_w4956_
	);
	LUT2 #(
		.INIT('h1)
	) name3777 (
		_w4902_,
		_w4913_,
		_w4957_
	);
	LUT2 #(
		.INIT('h2)
	) name3778 (
		_w4922_,
		_w4957_,
		_w4958_
	);
	LUT2 #(
		.INIT('h4)
	) name3779 (
		_w4888_,
		_w4898_,
		_w4959_
	);
	LUT2 #(
		.INIT('h2)
	) name3780 (
		_w4918_,
		_w4959_,
		_w4960_
	);
	LUT2 #(
		.INIT('h2)
	) name3781 (
		_w4871_,
		_w4881_,
		_w4961_
	);
	LUT2 #(
		.INIT('h4)
	) name3782 (
		_w4960_,
		_w4961_,
		_w4962_
	);
	LUT2 #(
		.INIT('h8)
	) name3783 (
		_w4906_,
		_w4925_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name3784 (
		_w4881_,
		_w4913_,
		_w4964_
	);
	LUT2 #(
		.INIT('h1)
	) name3785 (
		_w4870_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h1)
	) name3786 (
		_w4898_,
		_w4965_,
		_w4966_
	);
	LUT2 #(
		.INIT('h4)
	) name3787 (
		_w4865_,
		_w4870_,
		_w4967_
	);
	LUT2 #(
		.INIT('h8)
	) name3788 (
		_w4876_,
		_w4918_,
		_w4968_
	);
	LUT2 #(
		.INIT('h8)
	) name3789 (
		_w4967_,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name3790 (
		_w4966_,
		_w4969_,
		_w4970_
	);
	LUT2 #(
		.INIT('h2)
	) name3791 (
		_w4888_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h8)
	) name3792 (
		_w4919_,
		_w4923_,
		_w4972_
	);
	LUT2 #(
		.INIT('h8)
	) name3793 (
		_w4881_,
		_w4913_,
		_w4973_
	);
	LUT2 #(
		.INIT('h8)
	) name3794 (
		_w4959_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h2)
	) name3795 (
		_w4870_,
		_w4876_,
		_w4975_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		_w4901_,
		_w4975_,
		_w4976_
	);
	LUT2 #(
		.INIT('h1)
	) name3797 (
		_w4963_,
		_w4972_,
		_w4977_
	);
	LUT2 #(
		.INIT('h1)
	) name3798 (
		_w4974_,
		_w4976_,
		_w4978_
	);
	LUT2 #(
		.INIT('h8)
	) name3799 (
		_w4977_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h1)
	) name3800 (
		_w4956_,
		_w4962_,
		_w4980_
	);
	LUT2 #(
		.INIT('h8)
	) name3801 (
		_w4979_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w4955_,
		_w4958_,
		_w4982_
	);
	LUT2 #(
		.INIT('h8)
	) name3803 (
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h4)
	) name3804 (
		_w4971_,
		_w4983_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name3805 (
		_w4952_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('h8)
	) name3806 (
		\g5657_pad ,
		\g587_reg/NET0131 ,
		_w4986_
	);
	LUT2 #(
		.INIT('h8)
	) name3807 (
		\g1024_reg/NET0131 ,
		\g593_reg/NET0131 ,
		_w4987_
	);
	LUT2 #(
		.INIT('h8)
	) name3808 (
		\g1018_reg/NET0131 ,
		\g590_reg/NET0131 ,
		_w4988_
	);
	LUT2 #(
		.INIT('h8)
	) name3809 (
		\g1018_reg/NET0131 ,
		\g571_reg/NET0131 ,
		_w4989_
	);
	LUT2 #(
		.INIT('h8)
	) name3810 (
		\g1024_reg/NET0131 ,
		\g573_reg/NET0131 ,
		_w4990_
	);
	LUT2 #(
		.INIT('h8)
	) name3811 (
		\g5657_pad ,
		\g569_reg/NET0131 ,
		_w4991_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w4989_,
		_w4990_,
		_w4992_
	);
	LUT2 #(
		.INIT('h4)
	) name3813 (
		_w4991_,
		_w4992_,
		_w4993_
	);
	LUT2 #(
		.INIT('h8)
	) name3814 (
		\g185_reg/NET0131 ,
		\g524_reg/NET0131 ,
		_w4994_
	);
	LUT2 #(
		.INIT('h4)
	) name3815 (
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h1)
	) name3816 (
		_w4986_,
		_w4987_,
		_w4996_
	);
	LUT2 #(
		.INIT('h4)
	) name3817 (
		_w4988_,
		_w4996_,
		_w4997_
	);
	LUT2 #(
		.INIT('h4)
	) name3818 (
		_w4995_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w4952_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h2)
	) name3820 (
		_w4136_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h8)
	) name3821 (
		_w4939_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h4)
	) name3822 (
		_w4985_,
		_w5001_,
		_w5002_
	);
	LUT2 #(
		.INIT('h1)
	) name3823 (
		_w4860_,
		_w5002_,
		_w5003_
	);
	LUT2 #(
		.INIT('h4)
	) name3824 (
		\g1092_reg/NET0131 ,
		\g299_reg/NET0131 ,
		_w5004_
	);
	LUT2 #(
		.INIT('h8)
	) name3825 (
		\g305_reg/NET0131 ,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h1)
	) name3826 (
		_w1997_,
		_w5005_,
		_w5006_
	);
	LUT2 #(
		.INIT('h1)
	) name3827 (
		_w1826_,
		_w4136_,
		_w5007_
	);
	LUT2 #(
		.INIT('h8)
	) name3828 (
		_w4796_,
		_w4854_,
		_w5008_
	);
	LUT2 #(
		.INIT('h8)
	) name3829 (
		_w4827_,
		_w4856_,
		_w5009_
	);
	LUT2 #(
		.INIT('h4)
	) name3830 (
		_w5008_,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		_w5007_,
		_w5010_,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name3832 (
		_w2938_,
		_w4136_,
		_w5012_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		_w4216_,
		_w4273_,
		_w5013_
	);
	LUT2 #(
		.INIT('h2)
	) name3834 (
		_w4136_,
		_w4274_,
		_w5014_
	);
	LUT2 #(
		.INIT('h8)
	) name3835 (
		_w4259_,
		_w5014_,
		_w5015_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		_w5013_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h1)
	) name3837 (
		_w5012_,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h1)
	) name3838 (
		_w3673_,
		_w4136_,
		_w5018_
	);
	LUT2 #(
		.INIT('h8)
	) name3839 (
		_w4939_,
		_w4998_,
		_w5019_
	);
	LUT2 #(
		.INIT('h8)
	) name3840 (
		_w4984_,
		_w5000_,
		_w5020_
	);
	LUT2 #(
		.INIT('h4)
	) name3841 (
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		_w5018_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h8)
	) name3843 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w5023_
	);
	LUT2 #(
		.INIT('h1)
	) name3844 (
		_w2116_,
		_w2226_,
		_w5024_
	);
	LUT2 #(
		.INIT('h1)
	) name3845 (
		_w4465_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h2)
	) name3846 (
		_w5023_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h8)
	) name3847 (
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w5027_
	);
	LUT2 #(
		.INIT('h4)
	) name3848 (
		_w5025_,
		_w5027_,
		_w5028_
	);
	LUT2 #(
		.INIT('h8)
	) name3849 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w5029_
	);
	LUT2 #(
		.INIT('h4)
	) name3850 (
		_w5025_,
		_w5029_,
		_w5030_
	);
	LUT2 #(
		.INIT('h1)
	) name3851 (
		_w1281_,
		_w1418_,
		_w5031_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		_w3320_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h2)
	) name3853 (
		_w5023_,
		_w5032_,
		_w5033_
	);
	LUT2 #(
		.INIT('h2)
	) name3854 (
		_w5027_,
		_w5032_,
		_w5034_
	);
	LUT2 #(
		.INIT('h2)
	) name3855 (
		_w5029_,
		_w5032_,
		_w5035_
	);
	LUT2 #(
		.INIT('h4)
	) name3856 (
		_w2408_,
		_w3140_,
		_w5036_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w2531_,
		_w5036_,
		_w5037_
	);
	LUT2 #(
		.INIT('h2)
	) name3858 (
		_w5023_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h2)
	) name3859 (
		_w5027_,
		_w5037_,
		_w5039_
	);
	LUT2 #(
		.INIT('h2)
	) name3860 (
		_w5029_,
		_w5037_,
		_w5040_
	);
	LUT2 #(
		.INIT('h1)
	) name3861 (
		_w2693_,
		_w4473_,
		_w5041_
	);
	LUT2 #(
		.INIT('h2)
	) name3862 (
		_w5023_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h2)
	) name3863 (
		_w5027_,
		_w5041_,
		_w5043_
	);
	LUT2 #(
		.INIT('h2)
	) name3864 (
		_w5029_,
		_w5041_,
		_w5044_
	);
	LUT2 #(
		.INIT('h8)
	) name3865 (
		\g1018_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		_w5045_
	);
	LUT2 #(
		.INIT('h2)
	) name3866 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w5046_
	);
	LUT2 #(
		.INIT('h8)
	) name3867 (
		\g1326_reg/NET0131 ,
		_w5046_,
		_w5047_
	);
	LUT2 #(
		.INIT('h8)
	) name3868 (
		\g1319_reg/NET0131 ,
		_w5047_,
		_w5048_
	);
	LUT2 #(
		.INIT('h8)
	) name3869 (
		\g1339_reg/NET0131 ,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h8)
	) name3870 (
		\g1332_reg/NET0131 ,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h8)
	) name3871 (
		\g1346_reg/NET0131 ,
		_w5050_,
		_w5051_
	);
	LUT2 #(
		.INIT('h8)
	) name3872 (
		\g1358_reg/NET0131 ,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h8)
	) name3873 (
		\g1352_reg/NET0131 ,
		_w5052_,
		_w5053_
	);
	LUT2 #(
		.INIT('h8)
	) name3874 (
		\g1365_reg/NET0131 ,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		\g1372_reg/NET0131 ,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name3876 (
		\g1378_reg/NET0131 ,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h8)
	) name3877 (
		\g1378_reg/NET0131 ,
		_w5055_,
		_w5057_
	);
	LUT2 #(
		.INIT('h1)
	) name3878 (
		_w5045_,
		_w5056_,
		_w5058_
	);
	LUT2 #(
		.INIT('h4)
	) name3879 (
		_w5057_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h8)
	) name3880 (
		\g1095_reg/NET0131 ,
		\g7961_pad ,
		_w5060_
	);
	LUT2 #(
		.INIT('h8)
	) name3881 (
		\g1088_reg/NET0131 ,
		\g1101_reg/NET0131 ,
		_w5061_
	);
	LUT2 #(
		.INIT('h8)
	) name3882 (
		\g1092_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		_w5062_
	);
	LUT2 #(
		.INIT('h1)
	) name3883 (
		_w5060_,
		_w5061_,
		_w5063_
	);
	LUT2 #(
		.INIT('h4)
	) name3884 (
		_w5062_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h4)
	) name3885 (
		\g1114_reg/NET0131 ,
		\g7961_pad ,
		_w5065_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		\g1092_reg/NET0131 ,
		\g1115_reg/NET0131 ,
		_w5066_
	);
	LUT2 #(
		.INIT('h2)
	) name3887 (
		\g1088_reg/NET0131 ,
		\g1113_reg/NET0131 ,
		_w5067_
	);
	LUT2 #(
		.INIT('h1)
	) name3888 (
		_w5065_,
		_w5066_,
		_w5068_
	);
	LUT2 #(
		.INIT('h4)
	) name3889 (
		_w5067_,
		_w5068_,
		_w5069_
	);
	LUT2 #(
		.INIT('h1)
	) name3890 (
		_w5064_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h8)
	) name3891 (
		\g1563_reg/NET0131 ,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h8)
	) name3892 (
		\g1104_reg/NET0131 ,
		\g7961_pad ,
		_w5072_
	);
	LUT2 #(
		.INIT('h8)
	) name3893 (
		\g1088_reg/NET0131 ,
		\g1110_reg/NET0131 ,
		_w5073_
	);
	LUT2 #(
		.INIT('h8)
	) name3894 (
		\g1092_reg/NET0131 ,
		\g1107_reg/NET0131 ,
		_w5074_
	);
	LUT2 #(
		.INIT('h1)
	) name3895 (
		_w5072_,
		_w5073_,
		_w5075_
	);
	LUT2 #(
		.INIT('h4)
	) name3896 (
		_w5074_,
		_w5075_,
		_w5076_
	);
	LUT2 #(
		.INIT('h1)
	) name3897 (
		_w5071_,
		_w5076_,
		_w5077_
	);
	LUT2 #(
		.INIT('h1)
	) name3898 (
		_w2383_,
		_w5070_,
		_w5078_
	);
	LUT2 #(
		.INIT('h8)
	) name3899 (
		\g801_reg/NET0131 ,
		\g813_reg/NET0131 ,
		_w5079_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		\g785_reg/NET0131 ,
		\g789_reg/NET0131 ,
		_w5080_
	);
	LUT2 #(
		.INIT('h8)
	) name3901 (
		\g793_reg/NET0131 ,
		\g797_reg/NET0131 ,
		_w5081_
	);
	LUT2 #(
		.INIT('h8)
	) name3902 (
		\g805_reg/NET0131 ,
		\g809_reg/NET0131 ,
		_w5082_
	);
	LUT2 #(
		.INIT('h8)
	) name3903 (
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h8)
	) name3904 (
		_w5079_,
		_w5080_,
		_w5084_
	);
	LUT2 #(
		.INIT('h8)
	) name3905 (
		_w5083_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h1)
	) name3906 (
		_w2298_,
		_w2356_,
		_w5086_
	);
	LUT2 #(
		.INIT('h8)
	) name3907 (
		_w5085_,
		_w5086_,
		_w5087_
	);
	LUT2 #(
		.INIT('h2)
	) name3908 (
		\g1563_reg/NET0131 ,
		_w5078_,
		_w5088_
	);
	LUT2 #(
		.INIT('h8)
	) name3909 (
		_w5087_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h1)
	) name3910 (
		_w5077_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h8)
	) name3911 (
		\g408_reg/NET0131 ,
		\g7961_pad ,
		_w5091_
	);
	LUT2 #(
		.INIT('h8)
	) name3912 (
		\g1088_reg/NET0131 ,
		\g414_reg/NET0131 ,
		_w5092_
	);
	LUT2 #(
		.INIT('h8)
	) name3913 (
		\g1092_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w5093_
	);
	LUT2 #(
		.INIT('h1)
	) name3914 (
		_w5091_,
		_w5092_,
		_w5094_
	);
	LUT2 #(
		.INIT('h4)
	) name3915 (
		_w5093_,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h4)
	) name3916 (
		\g427_reg/NET0131 ,
		\g7961_pad ,
		_w5096_
	);
	LUT2 #(
		.INIT('h2)
	) name3917 (
		\g1092_reg/NET0131 ,
		\g428_reg/NET0131 ,
		_w5097_
	);
	LUT2 #(
		.INIT('h2)
	) name3918 (
		\g1088_reg/NET0131 ,
		\g426_reg/NET0131 ,
		_w5098_
	);
	LUT2 #(
		.INIT('h1)
	) name3919 (
		_w5096_,
		_w5097_,
		_w5099_
	);
	LUT2 #(
		.INIT('h4)
	) name3920 (
		_w5098_,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('h1)
	) name3921 (
		_w5095_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name3922 (
		\g1563_reg/NET0131 ,
		_w5101_,
		_w5102_
	);
	LUT2 #(
		.INIT('h8)
	) name3923 (
		\g417_reg/NET0131 ,
		\g7961_pad ,
		_w5103_
	);
	LUT2 #(
		.INIT('h8)
	) name3924 (
		\g1088_reg/NET0131 ,
		\g423_reg/NET0131 ,
		_w5104_
	);
	LUT2 #(
		.INIT('h8)
	) name3925 (
		\g1092_reg/NET0131 ,
		\g420_reg/NET0131 ,
		_w5105_
	);
	LUT2 #(
		.INIT('h1)
	) name3926 (
		_w5103_,
		_w5104_,
		_w5106_
	);
	LUT2 #(
		.INIT('h4)
	) name3927 (
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h1)
	) name3928 (
		_w5102_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h1)
	) name3929 (
		_w2116_,
		_w5101_,
		_w5109_
	);
	LUT2 #(
		.INIT('h8)
	) name3930 (
		\g113_reg/NET0131 ,
		\g125_reg/NET0131 ,
		_w5110_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		\g101_reg/NET0131 ,
		\g105_reg/NET0131 ,
		_w5111_
	);
	LUT2 #(
		.INIT('h8)
	) name3932 (
		\g109_reg/NET0131 ,
		\g117_reg/NET0131 ,
		_w5112_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		\g121_reg/NET0131 ,
		\g97_reg/NET0131 ,
		_w5113_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		_w5112_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h8)
	) name3935 (
		_w5110_,
		_w5111_,
		_w5115_
	);
	LUT2 #(
		.INIT('h8)
	) name3936 (
		_w5114_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w2034_,
		_w2047_,
		_w5117_
	);
	LUT2 #(
		.INIT('h8)
	) name3938 (
		_w5116_,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h2)
	) name3939 (
		\g1563_reg/NET0131 ,
		_w5109_,
		_w5119_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		_w5118_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h1)
	) name3941 (
		_w5108_,
		_w5120_,
		_w5121_
	);
	LUT2 #(
		.INIT('h8)
	) name3942 (
		\g2483_reg/NET0131 ,
		\g7961_pad ,
		_w5122_
	);
	LUT2 #(
		.INIT('h8)
	) name3943 (
		\g1088_reg/NET0131 ,
		\g2489_reg/NET0131 ,
		_w5123_
	);
	LUT2 #(
		.INIT('h8)
	) name3944 (
		\g1092_reg/NET0131 ,
		\g2486_reg/NET0131 ,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name3945 (
		_w5122_,
		_w5123_,
		_w5125_
	);
	LUT2 #(
		.INIT('h4)
	) name3946 (
		_w5124_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h4)
	) name3947 (
		\g2502_reg/NET0131 ,
		\g7961_pad ,
		_w5127_
	);
	LUT2 #(
		.INIT('h2)
	) name3948 (
		\g1092_reg/NET0131 ,
		\g2503_reg/NET0131 ,
		_w5128_
	);
	LUT2 #(
		.INIT('h2)
	) name3949 (
		\g1088_reg/NET0131 ,
		\g2501_reg/NET0131 ,
		_w5129_
	);
	LUT2 #(
		.INIT('h1)
	) name3950 (
		_w5127_,
		_w5128_,
		_w5130_
	);
	LUT2 #(
		.INIT('h4)
	) name3951 (
		_w5129_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h1)
	) name3952 (
		_w5126_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('h8)
	) name3953 (
		\g1563_reg/NET0131 ,
		_w5132_,
		_w5133_
	);
	LUT2 #(
		.INIT('h8)
	) name3954 (
		\g2492_reg/NET0131 ,
		\g7961_pad ,
		_w5134_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		\g1088_reg/NET0131 ,
		\g2498_reg/NET0131 ,
		_w5135_
	);
	LUT2 #(
		.INIT('h8)
	) name3956 (
		\g1092_reg/NET0131 ,
		\g2495_reg/NET0131 ,
		_w5136_
	);
	LUT2 #(
		.INIT('h1)
	) name3957 (
		_w5134_,
		_w5135_,
		_w5137_
	);
	LUT2 #(
		.INIT('h4)
	) name3958 (
		_w5136_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name3959 (
		_w5133_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h1)
	) name3960 (
		_w1281_,
		_w5132_,
		_w5140_
	);
	LUT2 #(
		.INIT('h8)
	) name3961 (
		\g2185_reg/NET0131 ,
		\g2200_reg/NET0131 ,
		_w5141_
	);
	LUT2 #(
		.INIT('h8)
	) name3962 (
		\g2165_reg/NET0131 ,
		\g2170_reg/NET0131 ,
		_w5142_
	);
	LUT2 #(
		.INIT('h8)
	) name3963 (
		\g2175_reg/NET0131 ,
		\g2180_reg/NET0131 ,
		_w5143_
	);
	LUT2 #(
		.INIT('h8)
	) name3964 (
		\g2190_reg/NET0131 ,
		\g2195_reg/NET0131 ,
		_w5144_
	);
	LUT2 #(
		.INIT('h8)
	) name3965 (
		_w5143_,
		_w5144_,
		_w5145_
	);
	LUT2 #(
		.INIT('h8)
	) name3966 (
		_w5141_,
		_w5142_,
		_w5146_
	);
	LUT2 #(
		.INIT('h8)
	) name3967 (
		_w5145_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h1)
	) name3968 (
		_w1223_,
		_w1268_,
		_w5148_
	);
	LUT2 #(
		.INIT('h8)
	) name3969 (
		_w5147_,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h2)
	) name3970 (
		\g1563_reg/NET0131 ,
		_w5140_,
		_w5150_
	);
	LUT2 #(
		.INIT('h8)
	) name3971 (
		_w5149_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h1)
	) name3972 (
		_w5139_,
		_w5151_,
		_w5152_
	);
	LUT2 #(
		.INIT('h4)
	) name3973 (
		\g1808_reg/NET0131 ,
		\g7961_pad ,
		_w5153_
	);
	LUT2 #(
		.INIT('h2)
	) name3974 (
		\g1092_reg/NET0131 ,
		\g1809_reg/NET0131 ,
		_w5154_
	);
	LUT2 #(
		.INIT('h2)
	) name3975 (
		\g1088_reg/NET0131 ,
		\g1807_reg/NET0131 ,
		_w5155_
	);
	LUT2 #(
		.INIT('h1)
	) name3976 (
		_w5153_,
		_w5154_,
		_w5156_
	);
	LUT2 #(
		.INIT('h4)
	) name3977 (
		_w5155_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h8)
	) name3978 (
		\g1789_reg/NET0131 ,
		\g7961_pad ,
		_w5158_
	);
	LUT2 #(
		.INIT('h8)
	) name3979 (
		\g1088_reg/NET0131 ,
		\g1795_reg/NET0131 ,
		_w5159_
	);
	LUT2 #(
		.INIT('h8)
	) name3980 (
		\g1092_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		_w5160_
	);
	LUT2 #(
		.INIT('h1)
	) name3981 (
		_w5158_,
		_w5159_,
		_w5161_
	);
	LUT2 #(
		.INIT('h4)
	) name3982 (
		_w5160_,
		_w5161_,
		_w5162_
	);
	LUT2 #(
		.INIT('h1)
	) name3983 (
		_w5157_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h8)
	) name3984 (
		\g1563_reg/NET0131 ,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h8)
	) name3985 (
		\g1798_reg/NET0131 ,
		\g7961_pad ,
		_w5165_
	);
	LUT2 #(
		.INIT('h8)
	) name3986 (
		\g1088_reg/NET0131 ,
		\g1804_reg/NET0131 ,
		_w5166_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		\g1092_reg/NET0131 ,
		\g1801_reg/NET0131 ,
		_w5167_
	);
	LUT2 #(
		.INIT('h1)
	) name3988 (
		_w5165_,
		_w5166_,
		_w5168_
	);
	LUT2 #(
		.INIT('h4)
	) name3989 (
		_w5167_,
		_w5168_,
		_w5169_
	);
	LUT2 #(
		.INIT('h1)
	) name3990 (
		_w5164_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h1)
	) name3991 (
		_w2579_,
		_w5163_,
		_w5171_
	);
	LUT2 #(
		.INIT('h8)
	) name3992 (
		\g1491_reg/NET0131 ,
		\g1506_reg/NET0131 ,
		_w5172_
	);
	LUT2 #(
		.INIT('h8)
	) name3993 (
		\g1471_reg/NET0131 ,
		\g1476_reg/NET0131 ,
		_w5173_
	);
	LUT2 #(
		.INIT('h8)
	) name3994 (
		\g1481_reg/NET0131 ,
		\g1486_reg/NET0131 ,
		_w5174_
	);
	LUT2 #(
		.INIT('h8)
	) name3995 (
		\g1496_reg/NET0131 ,
		\g1501_reg/NET0131 ,
		_w5175_
	);
	LUT2 #(
		.INIT('h8)
	) name3996 (
		_w5174_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('h8)
	) name3997 (
		_w5172_,
		_w5173_,
		_w5177_
	);
	LUT2 #(
		.INIT('h8)
	) name3998 (
		_w5176_,
		_w5177_,
		_w5178_
	);
	LUT2 #(
		.INIT('h1)
	) name3999 (
		_w2610_,
		_w2670_,
		_w5179_
	);
	LUT2 #(
		.INIT('h8)
	) name4000 (
		_w5178_,
		_w5179_,
		_w5180_
	);
	LUT2 #(
		.INIT('h2)
	) name4001 (
		\g1563_reg/NET0131 ,
		_w5171_,
		_w5181_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		_w5180_,
		_w5181_,
		_w5182_
	);
	LUT2 #(
		.INIT('h1)
	) name4003 (
		_w5170_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('h8)
	) name4004 (
		_w2399_,
		_w2542_,
		_w5184_
	);
	LUT2 #(
		.INIT('h8)
	) name4005 (
		_w2135_,
		_w2264_,
		_w5185_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		_w1186_,
		_w1292_,
		_w5186_
	);
	LUT2 #(
		.INIT('h8)
	) name4007 (
		_w2816_,
		_w2834_,
		_w5187_
	);
	LUT2 #(
		.INIT('h1)
	) name4008 (
		\g1563_reg/NET0131 ,
		_w5064_,
		_w5188_
	);
	LUT2 #(
		.INIT('h2)
	) name4009 (
		_w5076_,
		_w5087_,
		_w5189_
	);
	LUT2 #(
		.INIT('h4)
	) name4010 (
		_w2383_,
		_w5076_,
		_w5190_
	);
	LUT2 #(
		.INIT('h2)
	) name4011 (
		_w5087_,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h2)
	) name4012 (
		\g1563_reg/NET0131 ,
		_w5189_,
		_w5192_
	);
	LUT2 #(
		.INIT('h4)
	) name4013 (
		_w5191_,
		_w5192_,
		_w5193_
	);
	LUT2 #(
		.INIT('h4)
	) name4014 (
		_w5070_,
		_w5193_,
		_w5194_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w5188_,
		_w5194_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name4016 (
		\g1563_reg/NET0131 ,
		_w5095_,
		_w5196_
	);
	LUT2 #(
		.INIT('h2)
	) name4017 (
		_w5107_,
		_w5118_,
		_w5197_
	);
	LUT2 #(
		.INIT('h4)
	) name4018 (
		_w2116_,
		_w5107_,
		_w5198_
	);
	LUT2 #(
		.INIT('h2)
	) name4019 (
		_w5118_,
		_w5198_,
		_w5199_
	);
	LUT2 #(
		.INIT('h2)
	) name4020 (
		\g1563_reg/NET0131 ,
		_w5197_,
		_w5200_
	);
	LUT2 #(
		.INIT('h4)
	) name4021 (
		_w5199_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h4)
	) name4022 (
		_w5101_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w5196_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h1)
	) name4024 (
		\g1563_reg/NET0131 ,
		_w5126_,
		_w5204_
	);
	LUT2 #(
		.INIT('h2)
	) name4025 (
		_w5138_,
		_w5149_,
		_w5205_
	);
	LUT2 #(
		.INIT('h4)
	) name4026 (
		_w1281_,
		_w5138_,
		_w5206_
	);
	LUT2 #(
		.INIT('h2)
	) name4027 (
		_w5149_,
		_w5206_,
		_w5207_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		\g1563_reg/NET0131 ,
		_w5205_,
		_w5208_
	);
	LUT2 #(
		.INIT('h4)
	) name4029 (
		_w5207_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h4)
	) name4030 (
		_w5132_,
		_w5209_,
		_w5210_
	);
	LUT2 #(
		.INIT('h1)
	) name4031 (
		_w5204_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name4032 (
		\g1563_reg/NET0131 ,
		_w5162_,
		_w5212_
	);
	LUT2 #(
		.INIT('h2)
	) name4033 (
		_w5169_,
		_w5180_,
		_w5213_
	);
	LUT2 #(
		.INIT('h4)
	) name4034 (
		_w2579_,
		_w5169_,
		_w5214_
	);
	LUT2 #(
		.INIT('h2)
	) name4035 (
		_w5180_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h2)
	) name4036 (
		\g1563_reg/NET0131 ,
		_w5213_,
		_w5216_
	);
	LUT2 #(
		.INIT('h4)
	) name4037 (
		_w5215_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h4)
	) name4038 (
		_w5163_,
		_w5217_,
		_w5218_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		_w5212_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('h1)
	) name4040 (
		_w4136_,
		_w4854_,
		_w5220_
	);
	LUT2 #(
		.INIT('h1)
	) name4041 (
		_w4136_,
		_w4840_,
		_w5221_
	);
	LUT2 #(
		.INIT('h1)
	) name4042 (
		_w4136_,
		_w4998_,
		_w5222_
	);
	LUT2 #(
		.INIT('h1)
	) name4043 (
		_w4136_,
		_w4952_,
		_w5223_
	);
	LUT2 #(
		.INIT('h1)
	) name4044 (
		_w4136_,
		_w4273_,
		_w5224_
	);
	LUT2 #(
		.INIT('h1)
	) name4045 (
		_w4136_,
		_w4229_,
		_w5225_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		_w4136_,
		_w4421_,
		_w5226_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		_w4136_,
		_w4375_,
		_w5227_
	);
	LUT2 #(
		.INIT('h1)
	) name4048 (
		\g1372_reg/NET0131 ,
		_w5054_,
		_w5228_
	);
	LUT2 #(
		.INIT('h1)
	) name4049 (
		_w5045_,
		_w5055_,
		_w5229_
	);
	LUT2 #(
		.INIT('h4)
	) name4050 (
		_w5228_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h4)
	) name4051 (
		_w1451_,
		_w1465_,
		_w5231_
	);
	LUT2 #(
		.INIT('h2)
	) name4052 (
		_w1462_,
		_w5231_,
		_w5232_
	);
	LUT2 #(
		.INIT('h8)
	) name4053 (
		\g1088_reg/NET0131 ,
		_w5194_,
		_w5233_
	);
	LUT2 #(
		.INIT('h8)
	) name4054 (
		\g7961_pad ,
		_w5194_,
		_w5234_
	);
	LUT2 #(
		.INIT('h8)
	) name4055 (
		\g1092_reg/NET0131 ,
		_w5194_,
		_w5235_
	);
	LUT2 #(
		.INIT('h8)
	) name4056 (
		\g1088_reg/NET0131 ,
		_w5202_,
		_w5236_
	);
	LUT2 #(
		.INIT('h8)
	) name4057 (
		\g7961_pad ,
		_w5202_,
		_w5237_
	);
	LUT2 #(
		.INIT('h8)
	) name4058 (
		\g1092_reg/NET0131 ,
		_w5202_,
		_w5238_
	);
	LUT2 #(
		.INIT('h8)
	) name4059 (
		\g1088_reg/NET0131 ,
		_w5210_,
		_w5239_
	);
	LUT2 #(
		.INIT('h8)
	) name4060 (
		\g7961_pad ,
		_w5210_,
		_w5240_
	);
	LUT2 #(
		.INIT('h8)
	) name4061 (
		\g1092_reg/NET0131 ,
		_w5210_,
		_w5241_
	);
	LUT2 #(
		.INIT('h8)
	) name4062 (
		\g1088_reg/NET0131 ,
		_w5218_,
		_w5242_
	);
	LUT2 #(
		.INIT('h8)
	) name4063 (
		\g7961_pad ,
		_w5218_,
		_w5243_
	);
	LUT2 #(
		.INIT('h8)
	) name4064 (
		\g1092_reg/NET0131 ,
		_w5218_,
		_w5244_
	);
	LUT2 #(
		.INIT('h8)
	) name4065 (
		_w2266_,
		_w3092_,
		_w5245_
	);
	LUT2 #(
		.INIT('h1)
	) name4066 (
		\g1448_reg/NET0131 ,
		_w2200_,
		_w5246_
	);
	LUT2 #(
		.INIT('h2)
	) name4067 (
		\g1444_reg/NET0131 ,
		_w2209_,
		_w5247_
	);
	LUT2 #(
		.INIT('h4)
	) name4068 (
		\g1444_reg/NET0131 ,
		_w2209_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name4069 (
		_w5247_,
		_w5248_,
		_w5249_
	);
	LUT2 #(
		.INIT('h1)
	) name4070 (
		\g1466_reg/NET0131 ,
		_w2167_,
		_w5250_
	);
	LUT2 #(
		.INIT('h8)
	) name4071 (
		\g1435_reg/NET0131 ,
		_w2150_,
		_w5251_
	);
	LUT2 #(
		.INIT('h8)
	) name4072 (
		\g1466_reg/NET0131 ,
		_w2167_,
		_w5252_
	);
	LUT2 #(
		.INIT('h1)
	) name4073 (
		\g1435_reg/NET0131 ,
		_w2150_,
		_w5253_
	);
	LUT2 #(
		.INIT('h1)
	) name4074 (
		\g1426_reg/NET0131 ,
		_w2142_,
		_w5254_
	);
	LUT2 #(
		.INIT('h8)
	) name4075 (
		\g1426_reg/NET0131 ,
		_w2142_,
		_w5255_
	);
	LUT2 #(
		.INIT('h2)
	) name4076 (
		\g1462_reg/NET0131 ,
		_w2184_,
		_w5256_
	);
	LUT2 #(
		.INIT('h4)
	) name4077 (
		\g1462_reg/NET0131 ,
		_w2184_,
		_w5257_
	);
	LUT2 #(
		.INIT('h1)
	) name4078 (
		_w5256_,
		_w5257_,
		_w5258_
	);
	LUT2 #(
		.INIT('h1)
	) name4079 (
		\g2896_reg/NET0131 ,
		\g2900_reg/NET0131 ,
		_w5259_
	);
	LUT2 #(
		.INIT('h1)
	) name4080 (
		\g2892_reg/NET0131 ,
		\g2903_reg/NET0131 ,
		_w5260_
	);
	LUT2 #(
		.INIT('h4)
	) name4081 (
		\g2908_reg/NET0131 ,
		_w5260_,
		_w5261_
	);
	LUT2 #(
		.INIT('h8)
	) name4082 (
		_w5259_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h4)
	) name4083 (
		_w2014_,
		_w2019_,
		_w5263_
	);
	LUT2 #(
		.INIT('h4)
	) name4084 (
		_w2024_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h1)
	) name4085 (
		_w5262_,
		_w5264_,
		_w5265_
	);
	LUT2 #(
		.INIT('h1)
	) name4086 (
		\g1457_reg/NET0131 ,
		_w2192_,
		_w5266_
	);
	LUT2 #(
		.INIT('h8)
	) name4087 (
		\g1457_reg/NET0131 ,
		_w2192_,
		_w5267_
	);
	LUT2 #(
		.INIT('h8)
	) name4088 (
		\g1448_reg/NET0131 ,
		_w2200_,
		_w5268_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		\g1453_reg/NET0131 ,
		_w2217_,
		_w5269_
	);
	LUT2 #(
		.INIT('h2)
	) name4090 (
		\g1430_reg/NET0131 ,
		_w2159_,
		_w5270_
	);
	LUT2 #(
		.INIT('h4)
	) name4091 (
		\g1430_reg/NET0131 ,
		_w2159_,
		_w5271_
	);
	LUT2 #(
		.INIT('h1)
	) name4092 (
		_w5270_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h8)
	) name4093 (
		\g1439_reg/NET0131 ,
		_w2175_,
		_w5273_
	);
	LUT2 #(
		.INIT('h1)
	) name4094 (
		\g1439_reg/NET0131 ,
		_w2175_,
		_w5274_
	);
	LUT2 #(
		.INIT('h1)
	) name4095 (
		\g1453_reg/NET0131 ,
		_w2217_,
		_w5275_
	);
	LUT2 #(
		.INIT('h1)
	) name4096 (
		_w5246_,
		_w5250_,
		_w5276_
	);
	LUT2 #(
		.INIT('h1)
	) name4097 (
		_w5251_,
		_w5252_,
		_w5277_
	);
	LUT2 #(
		.INIT('h1)
	) name4098 (
		_w5253_,
		_w5254_,
		_w5278_
	);
	LUT2 #(
		.INIT('h1)
	) name4099 (
		_w5255_,
		_w5266_,
		_w5279_
	);
	LUT2 #(
		.INIT('h1)
	) name4100 (
		_w5267_,
		_w5268_,
		_w5280_
	);
	LUT2 #(
		.INIT('h1)
	) name4101 (
		_w5269_,
		_w5273_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name4102 (
		_w5274_,
		_w5275_,
		_w5282_
	);
	LUT2 #(
		.INIT('h8)
	) name4103 (
		_w5281_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h8)
	) name4104 (
		_w5279_,
		_w5280_,
		_w5284_
	);
	LUT2 #(
		.INIT('h8)
	) name4105 (
		_w5277_,
		_w5278_,
		_w5285_
	);
	LUT2 #(
		.INIT('h4)
	) name4106 (
		_w5249_,
		_w5276_,
		_w5286_
	);
	LUT2 #(
		.INIT('h1)
	) name4107 (
		_w5258_,
		_w5272_,
		_w5287_
	);
	LUT2 #(
		.INIT('h8)
	) name4108 (
		_w5286_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		_w5284_,
		_w5285_,
		_w5289_
	);
	LUT2 #(
		.INIT('h8)
	) name4110 (
		_w5265_,
		_w5283_,
		_w5290_
	);
	LUT2 #(
		.INIT('h8)
	) name4111 (
		_w5289_,
		_w5290_,
		_w5291_
	);
	LUT2 #(
		.INIT('h8)
	) name4112 (
		_w5288_,
		_w5291_,
		_w5292_
	);
	LUT2 #(
		.INIT('h1)
	) name4113 (
		_w5245_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h8)
	) name4114 (
		_w2550_,
		_w3131_,
		_w5294_
	);
	LUT2 #(
		.INIT('h1)
	) name4115 (
		\g1453_reg/NET0131 ,
		_w2419_,
		_w5295_
	);
	LUT2 #(
		.INIT('h1)
	) name4116 (
		\g1444_reg/NET0131 ,
		_w2436_,
		_w5296_
	);
	LUT2 #(
		.INIT('h1)
	) name4117 (
		\g1462_reg/NET0131 ,
		_w2452_,
		_w5297_
	);
	LUT2 #(
		.INIT('h1)
	) name4118 (
		\g1466_reg/NET0131 ,
		_w2510_,
		_w5298_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		\g1435_reg/NET0131 ,
		_w2444_,
		_w5299_
	);
	LUT2 #(
		.INIT('h1)
	) name4120 (
		\g1435_reg/NET0131 ,
		_w2444_,
		_w5300_
	);
	LUT2 #(
		.INIT('h8)
	) name4121 (
		\g1430_reg/NET0131 ,
		_w2482_,
		_w5301_
	);
	LUT2 #(
		.INIT('h8)
	) name4122 (
		\g1448_reg/NET0131 ,
		_w2491_,
		_w5302_
	);
	LUT2 #(
		.INIT('h8)
	) name4123 (
		\g1426_reg/NET0131 ,
		_w2427_,
		_w5303_
	);
	LUT2 #(
		.INIT('h8)
	) name4124 (
		\g1453_reg/NET0131 ,
		_w2419_,
		_w5304_
	);
	LUT2 #(
		.INIT('h1)
	) name4125 (
		\g1439_reg/NET0131 ,
		_w2500_,
		_w5305_
	);
	LUT2 #(
		.INIT('h1)
	) name4126 (
		\g1448_reg/NET0131 ,
		_w2491_,
		_w5306_
	);
	LUT2 #(
		.INIT('h8)
	) name4127 (
		\g1444_reg/NET0131 ,
		_w2436_,
		_w5307_
	);
	LUT2 #(
		.INIT('h4)
	) name4128 (
		_w2288_,
		_w2408_,
		_w5308_
	);
	LUT2 #(
		.INIT('h4)
	) name4129 (
		_w2413_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h1)
	) name4130 (
		_w5262_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h1)
	) name4131 (
		\g1426_reg/NET0131 ,
		_w2427_,
		_w5311_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		\g1430_reg/NET0131 ,
		_w2482_,
		_w5312_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		\g1457_reg/NET0131 ,
		_w2474_,
		_w5313_
	);
	LUT2 #(
		.INIT('h8)
	) name4134 (
		\g1439_reg/NET0131 ,
		_w2500_,
		_w5314_
	);
	LUT2 #(
		.INIT('h8)
	) name4135 (
		\g1457_reg/NET0131 ,
		_w2474_,
		_w5315_
	);
	LUT2 #(
		.INIT('h8)
	) name4136 (
		\g1462_reg/NET0131 ,
		_w2452_,
		_w5316_
	);
	LUT2 #(
		.INIT('h8)
	) name4137 (
		\g1466_reg/NET0131 ,
		_w2510_,
		_w5317_
	);
	LUT2 #(
		.INIT('h1)
	) name4138 (
		_w5295_,
		_w5296_,
		_w5318_
	);
	LUT2 #(
		.INIT('h1)
	) name4139 (
		_w5297_,
		_w5298_,
		_w5319_
	);
	LUT2 #(
		.INIT('h1)
	) name4140 (
		_w5299_,
		_w5300_,
		_w5320_
	);
	LUT2 #(
		.INIT('h1)
	) name4141 (
		_w5301_,
		_w5302_,
		_w5321_
	);
	LUT2 #(
		.INIT('h1)
	) name4142 (
		_w5303_,
		_w5304_,
		_w5322_
	);
	LUT2 #(
		.INIT('h1)
	) name4143 (
		_w5305_,
		_w5306_,
		_w5323_
	);
	LUT2 #(
		.INIT('h1)
	) name4144 (
		_w5307_,
		_w5311_,
		_w5324_
	);
	LUT2 #(
		.INIT('h1)
	) name4145 (
		_w5312_,
		_w5313_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name4146 (
		_w5314_,
		_w5315_,
		_w5326_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w5316_,
		_w5317_,
		_w5327_
	);
	LUT2 #(
		.INIT('h8)
	) name4148 (
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h8)
	) name4149 (
		_w5324_,
		_w5325_,
		_w5329_
	);
	LUT2 #(
		.INIT('h8)
	) name4150 (
		_w5322_,
		_w5323_,
		_w5330_
	);
	LUT2 #(
		.INIT('h8)
	) name4151 (
		_w5320_,
		_w5321_,
		_w5331_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		_w5318_,
		_w5319_,
		_w5332_
	);
	LUT2 #(
		.INIT('h8)
	) name4153 (
		_w5331_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h8)
	) name4154 (
		_w5329_,
		_w5330_,
		_w5334_
	);
	LUT2 #(
		.INIT('h8)
	) name4155 (
		_w5310_,
		_w5328_,
		_w5335_
	);
	LUT2 #(
		.INIT('h8)
	) name4156 (
		_w5334_,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h8)
	) name4157 (
		_w5333_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h1)
	) name4158 (
		_w5294_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h8)
	) name4159 (
		_w1304_,
		_w3308_,
		_w5339_
	);
	LUT2 #(
		.INIT('h1)
	) name4160 (
		\g1462_reg/NET0131 ,
		_w1355_,
		_w5340_
	);
	LUT2 #(
		.INIT('h1)
	) name4161 (
		\g1435_reg/NET0131 ,
		_w1338_,
		_w5341_
	);
	LUT2 #(
		.INIT('h4)
	) name4162 (
		_w1298_,
		_w1303_,
		_w5342_
	);
	LUT2 #(
		.INIT('h4)
	) name4163 (
		_w1309_,
		_w5342_,
		_w5343_
	);
	LUT2 #(
		.INIT('h1)
	) name4164 (
		_w5262_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h8)
	) name4165 (
		\g1444_reg/NET0131 ,
		_w1330_,
		_w5345_
	);
	LUT2 #(
		.INIT('h1)
	) name4166 (
		\g1453_reg/NET0131 ,
		_w1347_,
		_w5346_
	);
	LUT2 #(
		.INIT('h8)
	) name4167 (
		\g1435_reg/NET0131 ,
		_w1338_,
		_w5347_
	);
	LUT2 #(
		.INIT('h8)
	) name4168 (
		\g1453_reg/NET0131 ,
		_w1347_,
		_w5348_
	);
	LUT2 #(
		.INIT('h1)
	) name4169 (
		\g1466_reg/NET0131 ,
		_w1409_,
		_w5349_
	);
	LUT2 #(
		.INIT('h1)
	) name4170 (
		\g1430_reg/NET0131 ,
		_w1384_,
		_w5350_
	);
	LUT2 #(
		.INIT('h8)
	) name4171 (
		\g1457_reg/NET0131 ,
		_w1401_,
		_w5351_
	);
	LUT2 #(
		.INIT('h8)
	) name4172 (
		\g1426_reg/NET0131 ,
		_w1322_,
		_w5352_
	);
	LUT2 #(
		.INIT('h1)
	) name4173 (
		\g1457_reg/NET0131 ,
		_w1401_,
		_w5353_
	);
	LUT2 #(
		.INIT('h1)
	) name4174 (
		\g1444_reg/NET0131 ,
		_w1330_,
		_w5354_
	);
	LUT2 #(
		.INIT('h8)
	) name4175 (
		\g1439_reg/NET0131 ,
		_w1392_,
		_w5355_
	);
	LUT2 #(
		.INIT('h1)
	) name4176 (
		\g1426_reg/NET0131 ,
		_w1322_,
		_w5356_
	);
	LUT2 #(
		.INIT('h1)
	) name4177 (
		\g1439_reg/NET0131 ,
		_w1392_,
		_w5357_
	);
	LUT2 #(
		.INIT('h8)
	) name4178 (
		\g1430_reg/NET0131 ,
		_w1384_,
		_w5358_
	);
	LUT2 #(
		.INIT('h8)
	) name4179 (
		\g1462_reg/NET0131 ,
		_w1355_,
		_w5359_
	);
	LUT2 #(
		.INIT('h8)
	) name4180 (
		\g1466_reg/NET0131 ,
		_w1409_,
		_w5360_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		\g1448_reg/NET0131 ,
		_w1376_,
		_w5361_
	);
	LUT2 #(
		.INIT('h8)
	) name4182 (
		\g1448_reg/NET0131 ,
		_w1376_,
		_w5362_
	);
	LUT2 #(
		.INIT('h1)
	) name4183 (
		_w5340_,
		_w5341_,
		_w5363_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		_w5345_,
		_w5346_,
		_w5364_
	);
	LUT2 #(
		.INIT('h1)
	) name4185 (
		_w5347_,
		_w5348_,
		_w5365_
	);
	LUT2 #(
		.INIT('h1)
	) name4186 (
		_w5349_,
		_w5350_,
		_w5366_
	);
	LUT2 #(
		.INIT('h1)
	) name4187 (
		_w5351_,
		_w5352_,
		_w5367_
	);
	LUT2 #(
		.INIT('h1)
	) name4188 (
		_w5353_,
		_w5354_,
		_w5368_
	);
	LUT2 #(
		.INIT('h1)
	) name4189 (
		_w5355_,
		_w5356_,
		_w5369_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		_w5357_,
		_w5358_,
		_w5370_
	);
	LUT2 #(
		.INIT('h1)
	) name4191 (
		_w5359_,
		_w5360_,
		_w5371_
	);
	LUT2 #(
		.INIT('h1)
	) name4192 (
		_w5361_,
		_w5362_,
		_w5372_
	);
	LUT2 #(
		.INIT('h8)
	) name4193 (
		_w5371_,
		_w5372_,
		_w5373_
	);
	LUT2 #(
		.INIT('h8)
	) name4194 (
		_w5369_,
		_w5370_,
		_w5374_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		_w5367_,
		_w5368_,
		_w5375_
	);
	LUT2 #(
		.INIT('h8)
	) name4196 (
		_w5365_,
		_w5366_,
		_w5376_
	);
	LUT2 #(
		.INIT('h8)
	) name4197 (
		_w5363_,
		_w5364_,
		_w5377_
	);
	LUT2 #(
		.INIT('h8)
	) name4198 (
		_w5376_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h8)
	) name4199 (
		_w5374_,
		_w5375_,
		_w5379_
	);
	LUT2 #(
		.INIT('h8)
	) name4200 (
		_w5344_,
		_w5373_,
		_w5380_
	);
	LUT2 #(
		.INIT('h8)
	) name4201 (
		_w5379_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h8)
	) name4202 (
		_w5378_,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h1)
	) name4203 (
		_w5339_,
		_w5382_,
		_w5383_
	);
	LUT2 #(
		.INIT('h8)
	) name4204 (
		_w2836_,
		_w3259_,
		_w5384_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		\g1430_reg/NET0131 ,
		_w2615_,
		_w5385_
	);
	LUT2 #(
		.INIT('h1)
	) name4206 (
		\g1466_reg/NET0131 ,
		_w2624_,
		_w5386_
	);
	LUT2 #(
		.INIT('h1)
	) name4207 (
		\g1457_reg/NET0131 ,
		_w2593_,
		_w5387_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		\g1444_reg/NET0131 ,
		_w2653_,
		_w5388_
	);
	LUT2 #(
		.INIT('h8)
	) name4209 (
		\g1435_reg/NET0131 ,
		_w2662_,
		_w5389_
	);
	LUT2 #(
		.INIT('h1)
	) name4210 (
		\g1435_reg/NET0131 ,
		_w2662_,
		_w5390_
	);
	LUT2 #(
		.INIT('h8)
	) name4211 (
		\g1453_reg/NET0131 ,
		_w2645_,
		_w5391_
	);
	LUT2 #(
		.INIT('h8)
	) name4212 (
		\g1426_reg/NET0131 ,
		_w2675_,
		_w5392_
	);
	LUT2 #(
		.INIT('h8)
	) name4213 (
		\g1448_reg/NET0131 ,
		_w2585_,
		_w5393_
	);
	LUT2 #(
		.INIT('h8)
	) name4214 (
		\g1430_reg/NET0131 ,
		_w2615_,
		_w5394_
	);
	LUT2 #(
		.INIT('h1)
	) name4215 (
		\g1439_reg/NET0131 ,
		_w2602_,
		_w5395_
	);
	LUT2 #(
		.INIT('h1)
	) name4216 (
		\g1426_reg/NET0131 ,
		_w2675_,
		_w5396_
	);
	LUT2 #(
		.INIT('h8)
	) name4217 (
		\g1466_reg/NET0131 ,
		_w2624_,
		_w5397_
	);
	LUT2 #(
		.INIT('h2)
	) name4218 (
		_w2574_,
		_w2699_,
		_w5398_
	);
	LUT2 #(
		.INIT('h4)
	) name4219 (
		_w2720_,
		_w5398_,
		_w5399_
	);
	LUT2 #(
		.INIT('h1)
	) name4220 (
		_w5262_,
		_w5399_,
		_w5400_
	);
	LUT2 #(
		.INIT('h1)
	) name4221 (
		\g1448_reg/NET0131 ,
		_w2585_,
		_w5401_
	);
	LUT2 #(
		.INIT('h1)
	) name4222 (
		\g1453_reg/NET0131 ,
		_w2645_,
		_w5402_
	);
	LUT2 #(
		.INIT('h1)
	) name4223 (
		\g1462_reg/NET0131 ,
		_w2684_,
		_w5403_
	);
	LUT2 #(
		.INIT('h8)
	) name4224 (
		\g1439_reg/NET0131 ,
		_w2602_,
		_w5404_
	);
	LUT2 #(
		.INIT('h8)
	) name4225 (
		\g1462_reg/NET0131 ,
		_w2684_,
		_w5405_
	);
	LUT2 #(
		.INIT('h8)
	) name4226 (
		\g1457_reg/NET0131 ,
		_w2593_,
		_w5406_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		\g1444_reg/NET0131 ,
		_w2653_,
		_w5407_
	);
	LUT2 #(
		.INIT('h1)
	) name4228 (
		_w5385_,
		_w5386_,
		_w5408_
	);
	LUT2 #(
		.INIT('h1)
	) name4229 (
		_w5387_,
		_w5388_,
		_w5409_
	);
	LUT2 #(
		.INIT('h1)
	) name4230 (
		_w5389_,
		_w5390_,
		_w5410_
	);
	LUT2 #(
		.INIT('h1)
	) name4231 (
		_w5391_,
		_w5392_,
		_w5411_
	);
	LUT2 #(
		.INIT('h1)
	) name4232 (
		_w5393_,
		_w5394_,
		_w5412_
	);
	LUT2 #(
		.INIT('h1)
	) name4233 (
		_w5395_,
		_w5396_,
		_w5413_
	);
	LUT2 #(
		.INIT('h1)
	) name4234 (
		_w5397_,
		_w5401_,
		_w5414_
	);
	LUT2 #(
		.INIT('h1)
	) name4235 (
		_w5402_,
		_w5403_,
		_w5415_
	);
	LUT2 #(
		.INIT('h1)
	) name4236 (
		_w5404_,
		_w5405_,
		_w5416_
	);
	LUT2 #(
		.INIT('h1)
	) name4237 (
		_w5406_,
		_w5407_,
		_w5417_
	);
	LUT2 #(
		.INIT('h8)
	) name4238 (
		_w5416_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('h8)
	) name4239 (
		_w5414_,
		_w5415_,
		_w5419_
	);
	LUT2 #(
		.INIT('h8)
	) name4240 (
		_w5412_,
		_w5413_,
		_w5420_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		_w5410_,
		_w5411_,
		_w5421_
	);
	LUT2 #(
		.INIT('h8)
	) name4242 (
		_w5408_,
		_w5409_,
		_w5422_
	);
	LUT2 #(
		.INIT('h8)
	) name4243 (
		_w5421_,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h8)
	) name4244 (
		_w5419_,
		_w5420_,
		_w5424_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		_w5400_,
		_w5418_,
		_w5425_
	);
	LUT2 #(
		.INIT('h8)
	) name4246 (
		_w5424_,
		_w5425_,
		_w5426_
	);
	LUT2 #(
		.INIT('h8)
	) name4247 (
		_w5423_,
		_w5426_,
		_w5427_
	);
	LUT2 #(
		.INIT('h1)
	) name4248 (
		_w5384_,
		_w5427_,
		_w5428_
	);
	LUT2 #(
		.INIT('h2)
	) name4249 (
		\g1088_reg/NET0131 ,
		\g1559_reg/NET0131 ,
		_w5429_
	);
	LUT2 #(
		.INIT('h4)
	) name4250 (
		\g1560_reg/NET0131 ,
		\g7961_pad ,
		_w5430_
	);
	LUT2 #(
		.INIT('h2)
	) name4251 (
		\g1092_reg/NET0131 ,
		\g1561_reg/NET0131 ,
		_w5431_
	);
	LUT2 #(
		.INIT('h1)
	) name4252 (
		_w5429_,
		_w5430_,
		_w5432_
	);
	LUT2 #(
		.INIT('h4)
	) name4253 (
		_w5431_,
		_w5432_,
		_w5433_
	);
	LUT2 #(
		.INIT('h2)
	) name4254 (
		_w5178_,
		_w5433_,
		_w5434_
	);
	LUT2 #(
		.INIT('h2)
	) name4255 (
		\g1563_reg/NET0131 ,
		_w5434_,
		_w5435_
	);
	LUT2 #(
		.INIT('h8)
	) name4256 (
		\g1088_reg/NET0131 ,
		\g1816_reg/NET0131 ,
		_w5436_
	);
	LUT2 #(
		.INIT('h8)
	) name4257 (
		\g1092_reg/NET0131 ,
		\g1813_reg/NET0131 ,
		_w5437_
	);
	LUT2 #(
		.INIT('h8)
	) name4258 (
		\g1810_reg/NET0131 ,
		\g7961_pad ,
		_w5438_
	);
	LUT2 #(
		.INIT('h1)
	) name4259 (
		_w5436_,
		_w5437_,
		_w5439_
	);
	LUT2 #(
		.INIT('h4)
	) name4260 (
		_w5438_,
		_w5439_,
		_w5440_
	);
	LUT2 #(
		.INIT('h4)
	) name4261 (
		\g1563_reg/NET0131 ,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h1)
	) name4262 (
		_w5435_,
		_w5441_,
		_w5442_
	);
	LUT2 #(
		.INIT('h2)
	) name4263 (
		\g1092_reg/NET0131 ,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h1)
	) name4264 (
		\g1092_reg/NET0131 ,
		\g1813_reg/NET0131 ,
		_w5444_
	);
	LUT2 #(
		.INIT('h1)
	) name4265 (
		_w5443_,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('h2)
	) name4266 (
		\g1088_reg/NET0131 ,
		\g865_reg/NET0131 ,
		_w5446_
	);
	LUT2 #(
		.INIT('h2)
	) name4267 (
		\g7961_pad ,
		\g866_reg/NET0131 ,
		_w5447_
	);
	LUT2 #(
		.INIT('h2)
	) name4268 (
		\g1092_reg/NET0131 ,
		\g867_reg/NET0131 ,
		_w5448_
	);
	LUT2 #(
		.INIT('h1)
	) name4269 (
		_w5446_,
		_w5447_,
		_w5449_
	);
	LUT2 #(
		.INIT('h4)
	) name4270 (
		_w5448_,
		_w5449_,
		_w5450_
	);
	LUT2 #(
		.INIT('h2)
	) name4271 (
		_w5085_,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h2)
	) name4272 (
		\g1563_reg/NET0131 ,
		_w5451_,
		_w5452_
	);
	LUT2 #(
		.INIT('h8)
	) name4273 (
		\g1092_reg/NET0131 ,
		\g1119_reg/NET0131 ,
		_w5453_
	);
	LUT2 #(
		.INIT('h8)
	) name4274 (
		\g1088_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w5454_
	);
	LUT2 #(
		.INIT('h8)
	) name4275 (
		\g1116_reg/NET0131 ,
		\g7961_pad ,
		_w5455_
	);
	LUT2 #(
		.INIT('h1)
	) name4276 (
		_w5453_,
		_w5454_,
		_w5456_
	);
	LUT2 #(
		.INIT('h4)
	) name4277 (
		_w5455_,
		_w5456_,
		_w5457_
	);
	LUT2 #(
		.INIT('h4)
	) name4278 (
		\g1563_reg/NET0131 ,
		_w5457_,
		_w5458_
	);
	LUT2 #(
		.INIT('h1)
	) name4279 (
		_w5452_,
		_w5458_,
		_w5459_
	);
	LUT2 #(
		.INIT('h2)
	) name4280 (
		\g7961_pad ,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h1)
	) name4281 (
		\g1116_reg/NET0131 ,
		\g7961_pad ,
		_w5461_
	);
	LUT2 #(
		.INIT('h1)
	) name4282 (
		_w5460_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('h2)
	) name4283 (
		\g1092_reg/NET0131 ,
		_w5459_,
		_w5463_
	);
	LUT2 #(
		.INIT('h1)
	) name4284 (
		\g1092_reg/NET0131 ,
		\g1119_reg/NET0131 ,
		_w5464_
	);
	LUT2 #(
		.INIT('h1)
	) name4285 (
		_w5463_,
		_w5464_,
		_w5465_
	);
	LUT2 #(
		.INIT('h2)
	) name4286 (
		\g1088_reg/NET0131 ,
		_w5459_,
		_w5466_
	);
	LUT2 #(
		.INIT('h1)
	) name4287 (
		\g1088_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w5467_
	);
	LUT2 #(
		.INIT('h1)
	) name4288 (
		_w5466_,
		_w5467_,
		_w5468_
	);
	LUT2 #(
		.INIT('h4)
	) name4289 (
		\g1829_reg/NET0131 ,
		\g7961_pad ,
		_w5469_
	);
	LUT2 #(
		.INIT('h2)
	) name4290 (
		\g1092_reg/NET0131 ,
		\g1830_reg/NET0131 ,
		_w5470_
	);
	LUT2 #(
		.INIT('h2)
	) name4291 (
		\g1088_reg/NET0131 ,
		\g1828_reg/NET0131 ,
		_w5471_
	);
	LUT2 #(
		.INIT('h1)
	) name4292 (
		_w5469_,
		_w5470_,
		_w5472_
	);
	LUT2 #(
		.INIT('h4)
	) name4293 (
		_w5471_,
		_w5472_,
		_w5473_
	);
	LUT2 #(
		.INIT('h8)
	) name4294 (
		\g1819_reg/NET0131 ,
		\g7961_pad ,
		_w5474_
	);
	LUT2 #(
		.INIT('h8)
	) name4295 (
		\g1088_reg/NET0131 ,
		\g1825_reg/NET0131 ,
		_w5475_
	);
	LUT2 #(
		.INIT('h8)
	) name4296 (
		\g1092_reg/NET0131 ,
		\g1822_reg/NET0131 ,
		_w5476_
	);
	LUT2 #(
		.INIT('h1)
	) name4297 (
		_w5474_,
		_w5475_,
		_w5477_
	);
	LUT2 #(
		.INIT('h4)
	) name4298 (
		_w5476_,
		_w5477_,
		_w5478_
	);
	LUT2 #(
		.INIT('h2)
	) name4299 (
		_w5434_,
		_w5478_,
		_w5479_
	);
	LUT2 #(
		.INIT('h1)
	) name4300 (
		_w5434_,
		_w5440_,
		_w5480_
	);
	LUT2 #(
		.INIT('h8)
	) name4301 (
		_w5440_,
		_w5478_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name4302 (
		_w5480_,
		_w5481_,
		_w5482_
	);
	LUT2 #(
		.INIT('h2)
	) name4303 (
		\g1563_reg/NET0131 ,
		_w5479_,
		_w5483_
	);
	LUT2 #(
		.INIT('h8)
	) name4304 (
		_w5482_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h8)
	) name4305 (
		_w5473_,
		_w5484_,
		_w5485_
	);
	LUT2 #(
		.INIT('h4)
	) name4306 (
		_w5434_,
		_w5478_,
		_w5486_
	);
	LUT2 #(
		.INIT('h2)
	) name4307 (
		\g1563_reg/NET0131 ,
		_w5486_,
		_w5487_
	);
	LUT2 #(
		.INIT('h4)
	) name4308 (
		_w5482_,
		_w5487_,
		_w5488_
	);
	LUT2 #(
		.INIT('h1)
	) name4309 (
		_w5485_,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h2)
	) name4310 (
		\g1088_reg/NET0131 ,
		_w5489_,
		_w5490_
	);
	LUT2 #(
		.INIT('h2)
	) name4311 (
		\g7961_pad ,
		_w5489_,
		_w5491_
	);
	LUT2 #(
		.INIT('h2)
	) name4312 (
		\g1092_reg/NET0131 ,
		_w5489_,
		_w5492_
	);
	LUT2 #(
		.INIT('h4)
	) name4313 (
		\g448_reg/NET0131 ,
		\g7961_pad ,
		_w5493_
	);
	LUT2 #(
		.INIT('h2)
	) name4314 (
		\g1092_reg/NET0131 ,
		\g449_reg/NET0131 ,
		_w5494_
	);
	LUT2 #(
		.INIT('h2)
	) name4315 (
		\g1088_reg/NET0131 ,
		\g447_reg/NET0131 ,
		_w5495_
	);
	LUT2 #(
		.INIT('h1)
	) name4316 (
		_w5493_,
		_w5494_,
		_w5496_
	);
	LUT2 #(
		.INIT('h4)
	) name4317 (
		_w5495_,
		_w5496_,
		_w5497_
	);
	LUT2 #(
		.INIT('h8)
	) name4318 (
		\g429_reg/NET0131 ,
		\g7961_pad ,
		_w5498_
	);
	LUT2 #(
		.INIT('h8)
	) name4319 (
		\g1088_reg/NET0131 ,
		\g435_reg/NET0131 ,
		_w5499_
	);
	LUT2 #(
		.INIT('h8)
	) name4320 (
		\g1092_reg/NET0131 ,
		\g432_reg/NET0131 ,
		_w5500_
	);
	LUT2 #(
		.INIT('h1)
	) name4321 (
		_w5498_,
		_w5499_,
		_w5501_
	);
	LUT2 #(
		.INIT('h4)
	) name4322 (
		_w5500_,
		_w5501_,
		_w5502_
	);
	LUT2 #(
		.INIT('h2)
	) name4323 (
		\g1088_reg/NET0131 ,
		\g177_reg/NET0131 ,
		_w5503_
	);
	LUT2 #(
		.INIT('h4)
	) name4324 (
		\g178_reg/NET0131 ,
		\g7961_pad ,
		_w5504_
	);
	LUT2 #(
		.INIT('h2)
	) name4325 (
		\g1092_reg/NET0131 ,
		\g179_reg/NET0131 ,
		_w5505_
	);
	LUT2 #(
		.INIT('h1)
	) name4326 (
		_w5503_,
		_w5504_,
		_w5506_
	);
	LUT2 #(
		.INIT('h4)
	) name4327 (
		_w5505_,
		_w5506_,
		_w5507_
	);
	LUT2 #(
		.INIT('h2)
	) name4328 (
		_w5116_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h1)
	) name4329 (
		_w5502_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h8)
	) name4330 (
		\g438_reg/NET0131 ,
		\g7961_pad ,
		_w5510_
	);
	LUT2 #(
		.INIT('h8)
	) name4331 (
		\g1088_reg/NET0131 ,
		\g444_reg/NET0131 ,
		_w5511_
	);
	LUT2 #(
		.INIT('h8)
	) name4332 (
		\g1092_reg/NET0131 ,
		\g441_reg/NET0131 ,
		_w5512_
	);
	LUT2 #(
		.INIT('h1)
	) name4333 (
		_w5510_,
		_w5511_,
		_w5513_
	);
	LUT2 #(
		.INIT('h4)
	) name4334 (
		_w5512_,
		_w5513_,
		_w5514_
	);
	LUT2 #(
		.INIT('h4)
	) name4335 (
		_w5502_,
		_w5514_,
		_w5515_
	);
	LUT2 #(
		.INIT('h1)
	) name4336 (
		_w5508_,
		_w5514_,
		_w5516_
	);
	LUT2 #(
		.INIT('h1)
	) name4337 (
		_w5515_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('h2)
	) name4338 (
		\g1563_reg/NET0131 ,
		_w5509_,
		_w5518_
	);
	LUT2 #(
		.INIT('h4)
	) name4339 (
		_w5517_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h8)
	) name4340 (
		_w5497_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h8)
	) name4341 (
		_w5508_,
		_w5514_,
		_w5521_
	);
	LUT2 #(
		.INIT('h1)
	) name4342 (
		_w5509_,
		_w5521_,
		_w5522_
	);
	LUT2 #(
		.INIT('h2)
	) name4343 (
		\g1563_reg/NET0131 ,
		_w5515_,
		_w5523_
	);
	LUT2 #(
		.INIT('h4)
	) name4344 (
		_w5522_,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('h1)
	) name4345 (
		_w5520_,
		_w5524_,
		_w5525_
	);
	LUT2 #(
		.INIT('h2)
	) name4346 (
		\g7961_pad ,
		_w5525_,
		_w5526_
	);
	LUT2 #(
		.INIT('h8)
	) name4347 (
		_w5023_,
		_w5262_,
		_w5527_
	);
	LUT2 #(
		.INIT('h2)
	) name4348 (
		\g1088_reg/NET0131 ,
		_w5262_,
		_w5528_
	);
	LUT2 #(
		.INIT('h8)
	) name4349 (
		\g1466_reg/NET0131 ,
		_w5528_,
		_w5529_
	);
	LUT2 #(
		.INIT('h8)
	) name4350 (
		\g1462_reg/NET0131 ,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h8)
	) name4351 (
		\g1457_reg/NET0131 ,
		_w5530_,
		_w5531_
	);
	LUT2 #(
		.INIT('h8)
	) name4352 (
		\g1453_reg/NET0131 ,
		_w5531_,
		_w5532_
	);
	LUT2 #(
		.INIT('h8)
	) name4353 (
		\g1448_reg/NET0131 ,
		_w5532_,
		_w5533_
	);
	LUT2 #(
		.INIT('h8)
	) name4354 (
		\g1444_reg/NET0131 ,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h8)
	) name4355 (
		\g1439_reg/NET0131 ,
		_w5534_,
		_w5535_
	);
	LUT2 #(
		.INIT('h8)
	) name4356 (
		\g1435_reg/NET0131 ,
		_w5535_,
		_w5536_
	);
	LUT2 #(
		.INIT('h8)
	) name4357 (
		\g1430_reg/NET0131 ,
		_w5536_,
		_w5537_
	);
	LUT2 #(
		.INIT('h1)
	) name4358 (
		\g1426_reg/NET0131 ,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h8)
	) name4359 (
		\g1426_reg/NET0131 ,
		_w5537_,
		_w5539_
	);
	LUT2 #(
		.INIT('h1)
	) name4360 (
		_w5527_,
		_w5538_,
		_w5540_
	);
	LUT2 #(
		.INIT('h4)
	) name4361 (
		_w5539_,
		_w5540_,
		_w5541_
	);
	LUT2 #(
		.INIT('h2)
	) name4362 (
		\g1088_reg/NET0131 ,
		_w5525_,
		_w5542_
	);
	LUT2 #(
		.INIT('h2)
	) name4363 (
		\g1092_reg/NET0131 ,
		_w5525_,
		_w5543_
	);
	LUT2 #(
		.INIT('h4)
	) name4364 (
		\g1135_reg/NET0131 ,
		\g7961_pad ,
		_w5544_
	);
	LUT2 #(
		.INIT('h2)
	) name4365 (
		\g1092_reg/NET0131 ,
		\g1136_reg/NET0131 ,
		_w5545_
	);
	LUT2 #(
		.INIT('h2)
	) name4366 (
		\g1088_reg/NET0131 ,
		\g1134_reg/NET0131 ,
		_w5546_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		_w5544_,
		_w5545_,
		_w5547_
	);
	LUT2 #(
		.INIT('h4)
	) name4368 (
		_w5546_,
		_w5547_,
		_w5548_
	);
	LUT2 #(
		.INIT('h8)
	) name4369 (
		\g1125_reg/NET0131 ,
		\g7961_pad ,
		_w5549_
	);
	LUT2 #(
		.INIT('h8)
	) name4370 (
		\g1088_reg/NET0131 ,
		\g1131_reg/NET0131 ,
		_w5550_
	);
	LUT2 #(
		.INIT('h8)
	) name4371 (
		\g1092_reg/NET0131 ,
		\g1128_reg/NET0131 ,
		_w5551_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w5549_,
		_w5550_,
		_w5552_
	);
	LUT2 #(
		.INIT('h4)
	) name4373 (
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h2)
	) name4374 (
		_w5451_,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h1)
	) name4375 (
		_w5451_,
		_w5457_,
		_w5555_
	);
	LUT2 #(
		.INIT('h8)
	) name4376 (
		_w5457_,
		_w5553_,
		_w5556_
	);
	LUT2 #(
		.INIT('h1)
	) name4377 (
		_w5555_,
		_w5556_,
		_w5557_
	);
	LUT2 #(
		.INIT('h2)
	) name4378 (
		\g1563_reg/NET0131 ,
		_w5554_,
		_w5558_
	);
	LUT2 #(
		.INIT('h8)
	) name4379 (
		_w5557_,
		_w5558_,
		_w5559_
	);
	LUT2 #(
		.INIT('h8)
	) name4380 (
		_w5548_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h4)
	) name4381 (
		_w5451_,
		_w5553_,
		_w5561_
	);
	LUT2 #(
		.INIT('h2)
	) name4382 (
		\g1563_reg/NET0131 ,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h4)
	) name4383 (
		_w5557_,
		_w5562_,
		_w5563_
	);
	LUT2 #(
		.INIT('h1)
	) name4384 (
		_w5560_,
		_w5563_,
		_w5564_
	);
	LUT2 #(
		.INIT('h2)
	) name4385 (
		\g1088_reg/NET0131 ,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h2)
	) name4386 (
		\g7961_pad ,
		_w5564_,
		_w5566_
	);
	LUT2 #(
		.INIT('h2)
	) name4387 (
		\g1092_reg/NET0131 ,
		_w5564_,
		_w5567_
	);
	LUT2 #(
		.INIT('h4)
	) name4388 (
		\g2523_reg/NET0131 ,
		\g7961_pad ,
		_w5568_
	);
	LUT2 #(
		.INIT('h2)
	) name4389 (
		\g1092_reg/NET0131 ,
		\g2524_reg/NET0131 ,
		_w5569_
	);
	LUT2 #(
		.INIT('h2)
	) name4390 (
		\g1088_reg/NET0131 ,
		\g2522_reg/NET0131 ,
		_w5570_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w5568_,
		_w5569_,
		_w5571_
	);
	LUT2 #(
		.INIT('h4)
	) name4392 (
		_w5570_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h8)
	) name4393 (
		\g2504_reg/NET0131 ,
		\g7961_pad ,
		_w5573_
	);
	LUT2 #(
		.INIT('h8)
	) name4394 (
		\g1088_reg/NET0131 ,
		\g2510_reg/NET0131 ,
		_w5574_
	);
	LUT2 #(
		.INIT('h8)
	) name4395 (
		\g1092_reg/NET0131 ,
		\g2507_reg/NET0131 ,
		_w5575_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		_w5573_,
		_w5574_,
		_w5576_
	);
	LUT2 #(
		.INIT('h4)
	) name4397 (
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h2)
	) name4398 (
		\g1092_reg/NET0131 ,
		\g2255_reg/NET0131 ,
		_w5578_
	);
	LUT2 #(
		.INIT('h2)
	) name4399 (
		\g1088_reg/NET0131 ,
		\g2253_reg/NET0131 ,
		_w5579_
	);
	LUT2 #(
		.INIT('h4)
	) name4400 (
		\g2254_reg/NET0131 ,
		\g7961_pad ,
		_w5580_
	);
	LUT2 #(
		.INIT('h1)
	) name4401 (
		_w5578_,
		_w5579_,
		_w5581_
	);
	LUT2 #(
		.INIT('h4)
	) name4402 (
		_w5580_,
		_w5581_,
		_w5582_
	);
	LUT2 #(
		.INIT('h2)
	) name4403 (
		_w5147_,
		_w5582_,
		_w5583_
	);
	LUT2 #(
		.INIT('h1)
	) name4404 (
		_w5577_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h8)
	) name4405 (
		\g2513_reg/NET0131 ,
		\g7961_pad ,
		_w5585_
	);
	LUT2 #(
		.INIT('h8)
	) name4406 (
		\g1088_reg/NET0131 ,
		\g2519_reg/NET0131 ,
		_w5586_
	);
	LUT2 #(
		.INIT('h8)
	) name4407 (
		\g1092_reg/NET0131 ,
		\g2516_reg/NET0131 ,
		_w5587_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		_w5585_,
		_w5586_,
		_w5588_
	);
	LUT2 #(
		.INIT('h4)
	) name4409 (
		_w5587_,
		_w5588_,
		_w5589_
	);
	LUT2 #(
		.INIT('h4)
	) name4410 (
		_w5577_,
		_w5589_,
		_w5590_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w5583_,
		_w5589_,
		_w5591_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w5590_,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('h2)
	) name4413 (
		\g1563_reg/NET0131 ,
		_w5584_,
		_w5593_
	);
	LUT2 #(
		.INIT('h4)
	) name4414 (
		_w5592_,
		_w5593_,
		_w5594_
	);
	LUT2 #(
		.INIT('h8)
	) name4415 (
		_w5572_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('h8)
	) name4416 (
		_w5583_,
		_w5589_,
		_w5596_
	);
	LUT2 #(
		.INIT('h1)
	) name4417 (
		_w5584_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('h2)
	) name4418 (
		\g1563_reg/NET0131 ,
		_w5590_,
		_w5598_
	);
	LUT2 #(
		.INIT('h4)
	) name4419 (
		_w5597_,
		_w5598_,
		_w5599_
	);
	LUT2 #(
		.INIT('h1)
	) name4420 (
		_w5595_,
		_w5599_,
		_w5600_
	);
	LUT2 #(
		.INIT('h2)
	) name4421 (
		\g1088_reg/NET0131 ,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h2)
	) name4422 (
		\g7961_pad ,
		_w5600_,
		_w5602_
	);
	LUT2 #(
		.INIT('h2)
	) name4423 (
		\g1092_reg/NET0131 ,
		_w5600_,
		_w5603_
	);
	LUT2 #(
		.INIT('h1)
	) name4424 (
		_w2551_,
		_w5310_,
		_w5604_
	);
	LUT2 #(
		.INIT('h2)
	) name4425 (
		\g1092_reg/NET0131 ,
		_w5604_,
		_w5605_
	);
	LUT2 #(
		.INIT('h4)
	) name4426 (
		\g1045_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w5606_
	);
	LUT2 #(
		.INIT('h4)
	) name4427 (
		\g1048_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w5607_
	);
	LUT2 #(
		.INIT('h4)
	) name4428 (
		\g1056_reg/NET0131 ,
		\g7961_pad ,
		_w5608_
	);
	LUT2 #(
		.INIT('h1)
	) name4429 (
		_w5606_,
		_w5607_,
		_w5609_
	);
	LUT2 #(
		.INIT('h4)
	) name4430 (
		_w5608_,
		_w5609_,
		_w5610_
	);
	LUT2 #(
		.INIT('h4)
	) name4431 (
		\g1075_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w5611_
	);
	LUT2 #(
		.INIT('h4)
	) name4432 (
		\g1078_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w5612_
	);
	LUT2 #(
		.INIT('h4)
	) name4433 (
		\g1085_reg/NET0131 ,
		\g7961_pad ,
		_w5613_
	);
	LUT2 #(
		.INIT('h1)
	) name4434 (
		_w5611_,
		_w5612_,
		_w5614_
	);
	LUT2 #(
		.INIT('h4)
	) name4435 (
		_w5613_,
		_w5614_,
		_w5615_
	);
	LUT2 #(
		.INIT('h8)
	) name4436 (
		_w5610_,
		_w5615_,
		_w5616_
	);
	LUT2 #(
		.INIT('h4)
	) name4437 (
		\g1030_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w5617_
	);
	LUT2 #(
		.INIT('h4)
	) name4438 (
		\g1033_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w5618_
	);
	LUT2 #(
		.INIT('h4)
	) name4439 (
		\g1041_reg/NET0131 ,
		\g7961_pad ,
		_w5619_
	);
	LUT2 #(
		.INIT('h1)
	) name4440 (
		_w5617_,
		_w5618_,
		_w5620_
	);
	LUT2 #(
		.INIT('h4)
	) name4441 (
		_w5619_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('h2)
	) name4442 (
		\g3229_pad ,
		_w5621_,
		_w5622_
	);
	LUT2 #(
		.INIT('h4)
	) name4443 (
		\g3229_pad ,
		_w5621_,
		_w5623_
	);
	LUT2 #(
		.INIT('h1)
	) name4444 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h1)
	) name4445 (
		_w5616_,
		_w5624_,
		_w5625_
	);
	LUT2 #(
		.INIT('h8)
	) name4446 (
		_w5610_,
		_w5624_,
		_w5626_
	);
	LUT2 #(
		.INIT('h1)
	) name4447 (
		_w5625_,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h2)
	) name4448 (
		_w5605_,
		_w5627_,
		_w5628_
	);
	LUT2 #(
		.INIT('h2)
	) name4449 (
		\g1060_reg/NET0131 ,
		_w5605_,
		_w5629_
	);
	LUT2 #(
		.INIT('h1)
	) name4450 (
		_w5628_,
		_w5629_,
		_w5630_
	);
	LUT2 #(
		.INIT('h2)
	) name4451 (
		\g1088_reg/NET0131 ,
		_w5604_,
		_w5631_
	);
	LUT2 #(
		.INIT('h4)
	) name4452 (
		_w5627_,
		_w5631_,
		_w5632_
	);
	LUT2 #(
		.INIT('h2)
	) name4453 (
		\g1063_reg/NET0131 ,
		_w5631_,
		_w5633_
	);
	LUT2 #(
		.INIT('h1)
	) name4454 (
		_w5632_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h2)
	) name4455 (
		\g7961_pad ,
		_w5604_,
		_w5635_
	);
	LUT2 #(
		.INIT('h4)
	) name4456 (
		_w5627_,
		_w5635_,
		_w5636_
	);
	LUT2 #(
		.INIT('h2)
	) name4457 (
		\g1071_reg/NET0131 ,
		_w5635_,
		_w5637_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w5636_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h8)
	) name4459 (
		\g1871_reg/NET0131 ,
		\g5657_pad ,
		_w5639_
	);
	LUT2 #(
		.INIT('h8)
	) name4460 (
		\g1024_reg/NET0131 ,
		\g1877_reg/NET0131 ,
		_w5640_
	);
	LUT2 #(
		.INIT('h8)
	) name4461 (
		\g1018_reg/NET0131 ,
		\g1874_reg/NET0131 ,
		_w5641_
	);
	LUT2 #(
		.INIT('h1)
	) name4462 (
		_w5639_,
		_w5640_,
		_w5642_
	);
	LUT2 #(
		.INIT('h4)
	) name4463 (
		_w5641_,
		_w5642_,
		_w5643_
	);
	LUT2 #(
		.INIT('h1)
	) name4464 (
		_w1826_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h1)
	) name4465 (
		\g3002_reg/NET0131 ,
		\g3006_reg/NET0131 ,
		_w5645_
	);
	LUT2 #(
		.INIT('h1)
	) name4466 (
		\g3010_reg/NET0131 ,
		\g3013_reg/NET0131 ,
		_w5646_
	);
	LUT2 #(
		.INIT('h4)
	) name4467 (
		\g3024_reg/NET0131 ,
		_w5646_,
		_w5647_
	);
	LUT2 #(
		.INIT('h8)
	) name4468 (
		_w5645_,
		_w5647_,
		_w5648_
	);
	LUT2 #(
		.INIT('h1)
	) name4469 (
		_w5644_,
		_w5648_,
		_w5649_
	);
	LUT2 #(
		.INIT('h2)
	) name4470 (
		\g1196_reg/NET0131 ,
		_w1745_,
		_w5650_
	);
	LUT2 #(
		.INIT('h8)
	) name4471 (
		_w5643_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h1)
	) name4472 (
		_w5649_,
		_w5651_,
		_w5652_
	);
	LUT2 #(
		.INIT('h2)
	) name4473 (
		\g1024_reg/NET0131 ,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('h2)
	) name4474 (
		\g1955_reg/NET0131 ,
		_w5653_,
		_w5654_
	);
	LUT2 #(
		.INIT('h4)
	) name4475 (
		_w4737_,
		_w4760_,
		_w5655_
	);
	LUT2 #(
		.INIT('h1)
	) name4476 (
		_w4752_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h1)
	) name4477 (
		\g3229_pad ,
		_w5656_,
		_w5657_
	);
	LUT2 #(
		.INIT('h2)
	) name4478 (
		_w4760_,
		_w4776_,
		_w5658_
	);
	LUT2 #(
		.INIT('h4)
	) name4479 (
		_w4786_,
		_w5658_,
		_w5659_
	);
	LUT2 #(
		.INIT('h2)
	) name4480 (
		\g3229_pad ,
		_w5659_,
		_w5660_
	);
	LUT2 #(
		.INIT('h1)
	) name4481 (
		_w5657_,
		_w5660_,
		_w5661_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		_w5653_,
		_w5661_,
		_w5662_
	);
	LUT2 #(
		.INIT('h1)
	) name4483 (
		_w5654_,
		_w5662_,
		_w5663_
	);
	LUT2 #(
		.INIT('h2)
	) name4484 (
		\g5657_pad ,
		_w5652_,
		_w5664_
	);
	LUT2 #(
		.INIT('h2)
	) name4485 (
		\g1956_reg/NET0131 ,
		_w5664_,
		_w5665_
	);
	LUT2 #(
		.INIT('h8)
	) name4486 (
		_w5661_,
		_w5664_,
		_w5666_
	);
	LUT2 #(
		.INIT('h1)
	) name4487 (
		_w5665_,
		_w5666_,
		_w5667_
	);
	LUT2 #(
		.INIT('h2)
	) name4488 (
		\g1018_reg/NET0131 ,
		_w5652_,
		_w5668_
	);
	LUT2 #(
		.INIT('h2)
	) name4489 (
		\g1957_reg/NET0131 ,
		_w5668_,
		_w5669_
	);
	LUT2 #(
		.INIT('h8)
	) name4490 (
		_w5661_,
		_w5668_,
		_w5670_
	);
	LUT2 #(
		.INIT('h1)
	) name4491 (
		_w5669_,
		_w5670_,
		_w5671_
	);
	LUT2 #(
		.INIT('h8)
	) name4492 (
		_w2014_,
		_w2266_,
		_w5672_
	);
	LUT2 #(
		.INIT('h1)
	) name4493 (
		_w5265_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h2)
	) name4494 (
		\g1092_reg/NET0131 ,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h2)
	) name4495 (
		\g343_reg/NET0131 ,
		_w5674_,
		_w5675_
	);
	LUT2 #(
		.INIT('h2)
	) name4496 (
		\g1092_reg/NET0131 ,
		\g388_reg/NET0131 ,
		_w5676_
	);
	LUT2 #(
		.INIT('h2)
	) name4497 (
		\g1088_reg/NET0131 ,
		\g391_reg/NET0131 ,
		_w5677_
	);
	LUT2 #(
		.INIT('h4)
	) name4498 (
		\g398_reg/NET0131 ,
		\g7961_pad ,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name4499 (
		_w5676_,
		_w5677_,
		_w5679_
	);
	LUT2 #(
		.INIT('h4)
	) name4500 (
		_w5678_,
		_w5679_,
		_w5680_
	);
	LUT2 #(
		.INIT('h2)
	) name4501 (
		\g1088_reg/NET0131 ,
		\g346_reg/NET0131 ,
		_w5681_
	);
	LUT2 #(
		.INIT('h2)
	) name4502 (
		\g1092_reg/NET0131 ,
		\g343_reg/NET0131 ,
		_w5682_
	);
	LUT2 #(
		.INIT('h4)
	) name4503 (
		\g354_reg/NET0131 ,
		\g7961_pad ,
		_w5683_
	);
	LUT2 #(
		.INIT('h1)
	) name4504 (
		_w5681_,
		_w5682_,
		_w5684_
	);
	LUT2 #(
		.INIT('h4)
	) name4505 (
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT2 #(
		.INIT('h2)
	) name4506 (
		_w5680_,
		_w5685_,
		_w5686_
	);
	LUT2 #(
		.INIT('h2)
	) name4507 (
		\g1092_reg/NET0131 ,
		\g358_reg/NET0131 ,
		_w5687_
	);
	LUT2 #(
		.INIT('h2)
	) name4508 (
		\g1088_reg/NET0131 ,
		\g361_reg/NET0131 ,
		_w5688_
	);
	LUT2 #(
		.INIT('h4)
	) name4509 (
		\g369_reg/NET0131 ,
		\g7961_pad ,
		_w5689_
	);
	LUT2 #(
		.INIT('h1)
	) name4510 (
		_w5687_,
		_w5688_,
		_w5690_
	);
	LUT2 #(
		.INIT('h4)
	) name4511 (
		_w5689_,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('h2)
	) name4512 (
		\g1088_reg/NET0131 ,
		\g376_reg/NET0131 ,
		_w5692_
	);
	LUT2 #(
		.INIT('h4)
	) name4513 (
		\g384_reg/NET0131 ,
		\g7961_pad ,
		_w5693_
	);
	LUT2 #(
		.INIT('h2)
	) name4514 (
		\g1092_reg/NET0131 ,
		\g373_reg/NET0131 ,
		_w5694_
	);
	LUT2 #(
		.INIT('h1)
	) name4515 (
		_w5692_,
		_w5693_,
		_w5695_
	);
	LUT2 #(
		.INIT('h4)
	) name4516 (
		_w5694_,
		_w5695_,
		_w5696_
	);
	LUT2 #(
		.INIT('h4)
	) name4517 (
		_w5691_,
		_w5696_,
		_w5697_
	);
	LUT2 #(
		.INIT('h1)
	) name4518 (
		_w5686_,
		_w5697_,
		_w5698_
	);
	LUT2 #(
		.INIT('h1)
	) name4519 (
		\g3229_pad ,
		_w5698_,
		_w5699_
	);
	LUT2 #(
		.INIT('h1)
	) name4520 (
		_w5685_,
		_w5697_,
		_w5700_
	);
	LUT2 #(
		.INIT('h2)
	) name4521 (
		_w5680_,
		_w5700_,
		_w5701_
	);
	LUT2 #(
		.INIT('h2)
	) name4522 (
		\g3229_pad ,
		_w5701_,
		_w5702_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		_w5699_,
		_w5702_,
		_w5703_
	);
	LUT2 #(
		.INIT('h8)
	) name4524 (
		_w5674_,
		_w5703_,
		_w5704_
	);
	LUT2 #(
		.INIT('h1)
	) name4525 (
		_w5675_,
		_w5704_,
		_w5705_
	);
	LUT2 #(
		.INIT('h2)
	) name4526 (
		\g1088_reg/NET0131 ,
		_w5673_,
		_w5706_
	);
	LUT2 #(
		.INIT('h2)
	) name4527 (
		\g346_reg/NET0131 ,
		_w5706_,
		_w5707_
	);
	LUT2 #(
		.INIT('h8)
	) name4528 (
		_w5703_,
		_w5706_,
		_w5708_
	);
	LUT2 #(
		.INIT('h1)
	) name4529 (
		_w5707_,
		_w5708_,
		_w5709_
	);
	LUT2 #(
		.INIT('h2)
	) name4530 (
		\g7961_pad ,
		_w5673_,
		_w5710_
	);
	LUT2 #(
		.INIT('h2)
	) name4531 (
		\g354_reg/NET0131 ,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h8)
	) name4532 (
		_w5703_,
		_w5710_,
		_w5712_
	);
	LUT2 #(
		.INIT('h1)
	) name4533 (
		_w5711_,
		_w5712_,
		_w5713_
	);
	LUT2 #(
		.INIT('h2)
	) name4534 (
		\g3229_pad ,
		_w5685_,
		_w5714_
	);
	LUT2 #(
		.INIT('h4)
	) name4535 (
		\g3229_pad ,
		_w5685_,
		_w5715_
	);
	LUT2 #(
		.INIT('h1)
	) name4536 (
		_w5714_,
		_w5715_,
		_w5716_
	);
	LUT2 #(
		.INIT('h8)
	) name4537 (
		_w5691_,
		_w5716_,
		_w5717_
	);
	LUT2 #(
		.INIT('h8)
	) name4538 (
		_w5680_,
		_w5691_,
		_w5718_
	);
	LUT2 #(
		.INIT('h1)
	) name4539 (
		_w5716_,
		_w5718_,
		_w5719_
	);
	LUT2 #(
		.INIT('h1)
	) name4540 (
		_w5717_,
		_w5719_,
		_w5720_
	);
	LUT2 #(
		.INIT('h2)
	) name4541 (
		_w5674_,
		_w5720_,
		_w5721_
	);
	LUT2 #(
		.INIT('h2)
	) name4542 (
		\g373_reg/NET0131 ,
		_w5674_,
		_w5722_
	);
	LUT2 #(
		.INIT('h1)
	) name4543 (
		_w5721_,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h2)
	) name4544 (
		_w5706_,
		_w5720_,
		_w5724_
	);
	LUT2 #(
		.INIT('h2)
	) name4545 (
		\g376_reg/NET0131 ,
		_w5706_,
		_w5725_
	);
	LUT2 #(
		.INIT('h1)
	) name4546 (
		_w5724_,
		_w5725_,
		_w5726_
	);
	LUT2 #(
		.INIT('h2)
	) name4547 (
		_w5710_,
		_w5720_,
		_w5727_
	);
	LUT2 #(
		.INIT('h2)
	) name4548 (
		\g384_reg/NET0131 ,
		_w5710_,
		_w5728_
	);
	LUT2 #(
		.INIT('h1)
	) name4549 (
		_w5727_,
		_w5728_,
		_w5729_
	);
	LUT2 #(
		.INIT('h8)
	) name4550 (
		\g490_reg/NET0131 ,
		\g5657_pad ,
		_w5730_
	);
	LUT2 #(
		.INIT('h8)
	) name4551 (
		\g1024_reg/NET0131 ,
		\g496_reg/NET0131 ,
		_w5731_
	);
	LUT2 #(
		.INIT('h8)
	) name4552 (
		\g1018_reg/NET0131 ,
		\g493_reg/NET0131 ,
		_w5732_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w5730_,
		_w5731_,
		_w5733_
	);
	LUT2 #(
		.INIT('h4)
	) name4554 (
		_w5732_,
		_w5733_,
		_w5734_
	);
	LUT2 #(
		.INIT('h1)
	) name4555 (
		_w3673_,
		_w5734_,
		_w5735_
	);
	LUT2 #(
		.INIT('h1)
	) name4556 (
		_w5648_,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h2)
	) name4557 (
		\g1196_reg/NET0131 ,
		_w3754_,
		_w5737_
	);
	LUT2 #(
		.INIT('h8)
	) name4558 (
		_w5734_,
		_w5737_,
		_w5738_
	);
	LUT2 #(
		.INIT('h1)
	) name4559 (
		_w5736_,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h2)
	) name4560 (
		\g1024_reg/NET0131 ,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h2)
	) name4561 (
		\g575_reg/NET0131 ,
		_w5740_,
		_w5741_
	);
	LUT2 #(
		.INIT('h4)
	) name4562 (
		_w4881_,
		_w4898_,
		_w5742_
	);
	LUT2 #(
		.INIT('h1)
	) name4563 (
		_w4953_,
		_w5742_,
		_w5743_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		\g3229_pad ,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h2)
	) name4565 (
		_w4898_,
		_w4906_,
		_w5745_
	);
	LUT2 #(
		.INIT('h4)
	) name4566 (
		_w4919_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h2)
	) name4567 (
		\g3229_pad ,
		_w5746_,
		_w5747_
	);
	LUT2 #(
		.INIT('h1)
	) name4568 (
		_w5744_,
		_w5747_,
		_w5748_
	);
	LUT2 #(
		.INIT('h8)
	) name4569 (
		_w5740_,
		_w5748_,
		_w5749_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		_w5741_,
		_w5749_,
		_w5750_
	);
	LUT2 #(
		.INIT('h2)
	) name4571 (
		\g5657_pad ,
		_w5739_,
		_w5751_
	);
	LUT2 #(
		.INIT('h2)
	) name4572 (
		\g576_reg/NET0131 ,
		_w5751_,
		_w5752_
	);
	LUT2 #(
		.INIT('h8)
	) name4573 (
		_w5748_,
		_w5751_,
		_w5753_
	);
	LUT2 #(
		.INIT('h1)
	) name4574 (
		_w5752_,
		_w5753_,
		_w5754_
	);
	LUT2 #(
		.INIT('h2)
	) name4575 (
		\g1018_reg/NET0131 ,
		_w5739_,
		_w5755_
	);
	LUT2 #(
		.INIT('h2)
	) name4576 (
		\g577_reg/NET0131 ,
		_w5755_,
		_w5756_
	);
	LUT2 #(
		.INIT('h8)
	) name4577 (
		_w5748_,
		_w5755_,
		_w5757_
	);
	LUT2 #(
		.INIT('h1)
	) name4578 (
		_w5756_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h1)
	) name4579 (
		\g1018_reg/NET0131 ,
		\g16297_pad ,
		_w5759_
	);
	LUT2 #(
		.INIT('h4)
	) name4580 (
		\g506_reg/NET0131 ,
		_w5759_,
		_w5760_
	);
	LUT2 #(
		.INIT('h1)
	) name4581 (
		_w3868_,
		_w5760_,
		_w5761_
	);
	LUT2 #(
		.INIT('h8)
	) name4582 (
		\g1177_reg/NET0131 ,
		\g5657_pad ,
		_w5762_
	);
	LUT2 #(
		.INIT('h8)
	) name4583 (
		\g1024_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		_w5763_
	);
	LUT2 #(
		.INIT('h8)
	) name4584 (
		\g1018_reg/NET0131 ,
		\g1180_reg/NET0131 ,
		_w5764_
	);
	LUT2 #(
		.INIT('h1)
	) name4585 (
		_w5762_,
		_w5763_,
		_w5765_
	);
	LUT2 #(
		.INIT('h4)
	) name4586 (
		_w5764_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h1)
	) name4587 (
		_w2938_,
		_w5766_,
		_w5767_
	);
	LUT2 #(
		.INIT('h1)
	) name4588 (
		_w5648_,
		_w5767_,
		_w5768_
	);
	LUT2 #(
		.INIT('h2)
	) name4589 (
		\g1196_reg/NET0131 ,
		_w2929_,
		_w5769_
	);
	LUT2 #(
		.INIT('h8)
	) name4590 (
		_w5766_,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('h1)
	) name4591 (
		_w5768_,
		_w5770_,
		_w5771_
	);
	LUT2 #(
		.INIT('h2)
	) name4592 (
		\g1024_reg/NET0131 ,
		_w5771_,
		_w5772_
	);
	LUT2 #(
		.INIT('h2)
	) name4593 (
		\g1261_reg/NET0131 ,
		_w5772_,
		_w5773_
	);
	LUT2 #(
		.INIT('h1)
	) name4594 (
		_w4148_,
		_w4186_,
		_w5774_
	);
	LUT2 #(
		.INIT('h1)
	) name4595 (
		\g3229_pad ,
		_w5774_,
		_w5775_
	);
	LUT2 #(
		.INIT('h2)
	) name4596 (
		_w4142_,
		_w4204_,
		_w5776_
	);
	LUT2 #(
		.INIT('h4)
	) name4597 (
		_w4230_,
		_w5776_,
		_w5777_
	);
	LUT2 #(
		.INIT('h2)
	) name4598 (
		\g3229_pad ,
		_w5777_,
		_w5778_
	);
	LUT2 #(
		.INIT('h1)
	) name4599 (
		_w5775_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h8)
	) name4600 (
		_w5772_,
		_w5779_,
		_w5780_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		_w5773_,
		_w5780_,
		_w5781_
	);
	LUT2 #(
		.INIT('h2)
	) name4602 (
		\g5657_pad ,
		_w5771_,
		_w5782_
	);
	LUT2 #(
		.INIT('h2)
	) name4603 (
		\g1262_reg/NET0131 ,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h8)
	) name4604 (
		_w5779_,
		_w5782_,
		_w5784_
	);
	LUT2 #(
		.INIT('h1)
	) name4605 (
		_w5783_,
		_w5784_,
		_w5785_
	);
	LUT2 #(
		.INIT('h2)
	) name4606 (
		\g1018_reg/NET0131 ,
		_w5771_,
		_w5786_
	);
	LUT2 #(
		.INIT('h2)
	) name4607 (
		\g1263_reg/NET0131 ,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h8)
	) name4608 (
		_w5779_,
		_w5786_,
		_w5788_
	);
	LUT2 #(
		.INIT('h1)
	) name4609 (
		_w5787_,
		_w5788_,
		_w5789_
	);
	LUT2 #(
		.INIT('h4)
	) name4610 (
		_w4142_,
		_w4153_,
		_w5790_
	);
	LUT2 #(
		.INIT('h1)
	) name4611 (
		_w4189_,
		_w4230_,
		_w5791_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		\g3229_pad ,
		_w5791_,
		_w5792_
	);
	LUT2 #(
		.INIT('h8)
	) name4613 (
		\g3229_pad ,
		_w5791_,
		_w5793_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		_w5790_,
		_w5792_,
		_w5794_
	);
	LUT2 #(
		.INIT('h4)
	) name4615 (
		_w5793_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h2)
	) name4616 (
		_w5772_,
		_w5795_,
		_w5796_
	);
	LUT2 #(
		.INIT('h2)
	) name4617 (
		\g1267_reg/NET0131 ,
		_w5772_,
		_w5797_
	);
	LUT2 #(
		.INIT('h1)
	) name4618 (
		_w5796_,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h1)
	) name4619 (
		_w1310_,
		_w5344_,
		_w5799_
	);
	LUT2 #(
		.INIT('h2)
	) name4620 (
		\g1092_reg/NET0131 ,
		_w5799_,
		_w5800_
	);
	LUT2 #(
		.INIT('h2)
	) name4621 (
		\g2418_reg/NET0131 ,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h2)
	) name4622 (
		\g1092_reg/NET0131 ,
		\g2463_reg/NET0131 ,
		_w5802_
	);
	LUT2 #(
		.INIT('h2)
	) name4623 (
		\g1088_reg/NET0131 ,
		\g2466_reg/NET0131 ,
		_w5803_
	);
	LUT2 #(
		.INIT('h4)
	) name4624 (
		\g2473_reg/NET0131 ,
		\g7961_pad ,
		_w5804_
	);
	LUT2 #(
		.INIT('h1)
	) name4625 (
		_w5802_,
		_w5803_,
		_w5805_
	);
	LUT2 #(
		.INIT('h4)
	) name4626 (
		_w5804_,
		_w5805_,
		_w5806_
	);
	LUT2 #(
		.INIT('h2)
	) name4627 (
		\g1088_reg/NET0131 ,
		\g2421_reg/NET0131 ,
		_w5807_
	);
	LUT2 #(
		.INIT('h2)
	) name4628 (
		\g1092_reg/NET0131 ,
		\g2418_reg/NET0131 ,
		_w5808_
	);
	LUT2 #(
		.INIT('h4)
	) name4629 (
		\g2429_reg/NET0131 ,
		\g7961_pad ,
		_w5809_
	);
	LUT2 #(
		.INIT('h1)
	) name4630 (
		_w5807_,
		_w5808_,
		_w5810_
	);
	LUT2 #(
		.INIT('h4)
	) name4631 (
		_w5809_,
		_w5810_,
		_w5811_
	);
	LUT2 #(
		.INIT('h2)
	) name4632 (
		_w5806_,
		_w5811_,
		_w5812_
	);
	LUT2 #(
		.INIT('h2)
	) name4633 (
		\g1092_reg/NET0131 ,
		\g2433_reg/NET0131 ,
		_w5813_
	);
	LUT2 #(
		.INIT('h2)
	) name4634 (
		\g1088_reg/NET0131 ,
		\g2436_reg/NET0131 ,
		_w5814_
	);
	LUT2 #(
		.INIT('h4)
	) name4635 (
		\g2444_reg/NET0131 ,
		\g7961_pad ,
		_w5815_
	);
	LUT2 #(
		.INIT('h1)
	) name4636 (
		_w5813_,
		_w5814_,
		_w5816_
	);
	LUT2 #(
		.INIT('h4)
	) name4637 (
		_w5815_,
		_w5816_,
		_w5817_
	);
	LUT2 #(
		.INIT('h2)
	) name4638 (
		\g1088_reg/NET0131 ,
		\g2451_reg/NET0131 ,
		_w5818_
	);
	LUT2 #(
		.INIT('h4)
	) name4639 (
		\g2459_reg/NET0131 ,
		\g7961_pad ,
		_w5819_
	);
	LUT2 #(
		.INIT('h2)
	) name4640 (
		\g1092_reg/NET0131 ,
		\g2448_reg/NET0131 ,
		_w5820_
	);
	LUT2 #(
		.INIT('h1)
	) name4641 (
		_w5818_,
		_w5819_,
		_w5821_
	);
	LUT2 #(
		.INIT('h4)
	) name4642 (
		_w5820_,
		_w5821_,
		_w5822_
	);
	LUT2 #(
		.INIT('h4)
	) name4643 (
		_w5817_,
		_w5822_,
		_w5823_
	);
	LUT2 #(
		.INIT('h1)
	) name4644 (
		_w5812_,
		_w5823_,
		_w5824_
	);
	LUT2 #(
		.INIT('h1)
	) name4645 (
		\g3229_pad ,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h1)
	) name4646 (
		_w5811_,
		_w5823_,
		_w5826_
	);
	LUT2 #(
		.INIT('h2)
	) name4647 (
		_w5806_,
		_w5826_,
		_w5827_
	);
	LUT2 #(
		.INIT('h2)
	) name4648 (
		\g3229_pad ,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h1)
	) name4649 (
		_w5825_,
		_w5828_,
		_w5829_
	);
	LUT2 #(
		.INIT('h8)
	) name4650 (
		_w5800_,
		_w5829_,
		_w5830_
	);
	LUT2 #(
		.INIT('h1)
	) name4651 (
		_w5801_,
		_w5830_,
		_w5831_
	);
	LUT2 #(
		.INIT('h2)
	) name4652 (
		_w5782_,
		_w5795_,
		_w5832_
	);
	LUT2 #(
		.INIT('h2)
	) name4653 (
		\g1268_reg/NET0131 ,
		_w5782_,
		_w5833_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w5832_,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		_w5786_,
		_w5795_,
		_w5835_
	);
	LUT2 #(
		.INIT('h2)
	) name4656 (
		\g1269_reg/NET0131 ,
		_w5786_,
		_w5836_
	);
	LUT2 #(
		.INIT('h1)
	) name4657 (
		_w5835_,
		_w5836_,
		_w5837_
	);
	LUT2 #(
		.INIT('h2)
	) name4658 (
		\g1088_reg/NET0131 ,
		_w5799_,
		_w5838_
	);
	LUT2 #(
		.INIT('h2)
	) name4659 (
		\g2421_reg/NET0131 ,
		_w5838_,
		_w5839_
	);
	LUT2 #(
		.INIT('h8)
	) name4660 (
		_w5829_,
		_w5838_,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name4661 (
		_w5839_,
		_w5840_,
		_w5841_
	);
	LUT2 #(
		.INIT('h2)
	) name4662 (
		\g7961_pad ,
		_w5799_,
		_w5842_
	);
	LUT2 #(
		.INIT('h2)
	) name4663 (
		\g2429_reg/NET0131 ,
		_w5842_,
		_w5843_
	);
	LUT2 #(
		.INIT('h8)
	) name4664 (
		_w5829_,
		_w5842_,
		_w5844_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		_w5843_,
		_w5844_,
		_w5845_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		\g3229_pad ,
		_w5811_,
		_w5846_
	);
	LUT2 #(
		.INIT('h4)
	) name4667 (
		\g3229_pad ,
		_w5811_,
		_w5847_
	);
	LUT2 #(
		.INIT('h1)
	) name4668 (
		_w5846_,
		_w5847_,
		_w5848_
	);
	LUT2 #(
		.INIT('h8)
	) name4669 (
		_w5817_,
		_w5848_,
		_w5849_
	);
	LUT2 #(
		.INIT('h8)
	) name4670 (
		_w5806_,
		_w5817_,
		_w5850_
	);
	LUT2 #(
		.INIT('h1)
	) name4671 (
		_w5848_,
		_w5850_,
		_w5851_
	);
	LUT2 #(
		.INIT('h1)
	) name4672 (
		_w5849_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h2)
	) name4673 (
		_w5800_,
		_w5852_,
		_w5853_
	);
	LUT2 #(
		.INIT('h2)
	) name4674 (
		\g2448_reg/NET0131 ,
		_w5800_,
		_w5854_
	);
	LUT2 #(
		.INIT('h1)
	) name4675 (
		_w5853_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h2)
	) name4676 (
		_w5838_,
		_w5852_,
		_w5856_
	);
	LUT2 #(
		.INIT('h2)
	) name4677 (
		\g2451_reg/NET0131 ,
		_w5838_,
		_w5857_
	);
	LUT2 #(
		.INIT('h1)
	) name4678 (
		_w5856_,
		_w5857_,
		_w5858_
	);
	LUT2 #(
		.INIT('h2)
	) name4679 (
		_w5842_,
		_w5852_,
		_w5859_
	);
	LUT2 #(
		.INIT('h2)
	) name4680 (
		\g2459_reg/NET0131 ,
		_w5842_,
		_w5860_
	);
	LUT2 #(
		.INIT('h1)
	) name4681 (
		_w5859_,
		_w5860_,
		_w5861_
	);
	LUT2 #(
		.INIT('h2)
	) name4682 (
		\g1030_reg/NET0131 ,
		_w5605_,
		_w5862_
	);
	LUT2 #(
		.INIT('h4)
	) name4683 (
		\g1063_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w5863_
	);
	LUT2 #(
		.INIT('h4)
	) name4684 (
		\g1071_reg/NET0131 ,
		\g7961_pad ,
		_w5864_
	);
	LUT2 #(
		.INIT('h4)
	) name4685 (
		\g1060_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w5865_
	);
	LUT2 #(
		.INIT('h1)
	) name4686 (
		_w5863_,
		_w5864_,
		_w5866_
	);
	LUT2 #(
		.INIT('h4)
	) name4687 (
		_w5865_,
		_w5866_,
		_w5867_
	);
	LUT2 #(
		.INIT('h4)
	) name4688 (
		_w5610_,
		_w5867_,
		_w5868_
	);
	LUT2 #(
		.INIT('h2)
	) name4689 (
		_w5615_,
		_w5621_,
		_w5869_
	);
	LUT2 #(
		.INIT('h1)
	) name4690 (
		_w5868_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h1)
	) name4691 (
		\g3229_pad ,
		_w5870_,
		_w5871_
	);
	LUT2 #(
		.INIT('h1)
	) name4692 (
		_w5621_,
		_w5868_,
		_w5872_
	);
	LUT2 #(
		.INIT('h2)
	) name4693 (
		_w5615_,
		_w5872_,
		_w5873_
	);
	LUT2 #(
		.INIT('h2)
	) name4694 (
		\g3229_pad ,
		_w5873_,
		_w5874_
	);
	LUT2 #(
		.INIT('h1)
	) name4695 (
		_w5871_,
		_w5874_,
		_w5875_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		_w5605_,
		_w5875_,
		_w5876_
	);
	LUT2 #(
		.INIT('h1)
	) name4697 (
		_w5862_,
		_w5876_,
		_w5877_
	);
	LUT2 #(
		.INIT('h8)
	) name4698 (
		\g2565_reg/NET0131 ,
		\g5657_pad ,
		_w5878_
	);
	LUT2 #(
		.INIT('h8)
	) name4699 (
		\g1024_reg/NET0131 ,
		\g2571_reg/NET0131 ,
		_w5879_
	);
	LUT2 #(
		.INIT('h8)
	) name4700 (
		\g1018_reg/NET0131 ,
		\g2568_reg/NET0131 ,
		_w5880_
	);
	LUT2 #(
		.INIT('h1)
	) name4701 (
		_w5878_,
		_w5879_,
		_w5881_
	);
	LUT2 #(
		.INIT('h4)
	) name4702 (
		_w5880_,
		_w5881_,
		_w5882_
	);
	LUT2 #(
		.INIT('h1)
	) name4703 (
		_w1643_,
		_w5882_,
		_w5883_
	);
	LUT2 #(
		.INIT('h1)
	) name4704 (
		_w5648_,
		_w5883_,
		_w5884_
	);
	LUT2 #(
		.INIT('h2)
	) name4705 (
		\g1196_reg/NET0131 ,
		_w1633_,
		_w5885_
	);
	LUT2 #(
		.INIT('h8)
	) name4706 (
		_w5882_,
		_w5885_,
		_w5886_
	);
	LUT2 #(
		.INIT('h1)
	) name4707 (
		_w5884_,
		_w5886_,
		_w5887_
	);
	LUT2 #(
		.INIT('h2)
	) name4708 (
		\g1024_reg/NET0131 ,
		_w5887_,
		_w5888_
	);
	LUT2 #(
		.INIT('h2)
	) name4709 (
		\g2649_reg/NET0131 ,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h1)
	) name4710 (
		_w4391_,
		_w4395_,
		_w5890_
	);
	LUT2 #(
		.INIT('h1)
	) name4711 (
		\g3229_pad ,
		_w5890_,
		_w5891_
	);
	LUT2 #(
		.INIT('h2)
	) name4712 (
		_w4287_,
		_w4320_,
		_w5892_
	);
	LUT2 #(
		.INIT('h4)
	) name4713 (
		_w4377_,
		_w5892_,
		_w5893_
	);
	LUT2 #(
		.INIT('h2)
	) name4714 (
		\g3229_pad ,
		_w5893_,
		_w5894_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w5891_,
		_w5894_,
		_w5895_
	);
	LUT2 #(
		.INIT('h8)
	) name4716 (
		_w5888_,
		_w5895_,
		_w5896_
	);
	LUT2 #(
		.INIT('h1)
	) name4717 (
		_w5889_,
		_w5896_,
		_w5897_
	);
	LUT2 #(
		.INIT('h1)
	) name4718 (
		_w2837_,
		_w5400_,
		_w5898_
	);
	LUT2 #(
		.INIT('h2)
	) name4719 (
		\g1092_reg/NET0131 ,
		_w5898_,
		_w5899_
	);
	LUT2 #(
		.INIT('h2)
	) name4720 (
		\g1724_reg/NET0131 ,
		_w5899_,
		_w5900_
	);
	LUT2 #(
		.INIT('h2)
	) name4721 (
		\g1092_reg/NET0131 ,
		\g1769_reg/NET0131 ,
		_w5901_
	);
	LUT2 #(
		.INIT('h2)
	) name4722 (
		\g1088_reg/NET0131 ,
		\g1772_reg/NET0131 ,
		_w5902_
	);
	LUT2 #(
		.INIT('h4)
	) name4723 (
		\g1779_reg/NET0131 ,
		\g7961_pad ,
		_w5903_
	);
	LUT2 #(
		.INIT('h1)
	) name4724 (
		_w5901_,
		_w5902_,
		_w5904_
	);
	LUT2 #(
		.INIT('h4)
	) name4725 (
		_w5903_,
		_w5904_,
		_w5905_
	);
	LUT2 #(
		.INIT('h2)
	) name4726 (
		\g1088_reg/NET0131 ,
		\g1727_reg/NET0131 ,
		_w5906_
	);
	LUT2 #(
		.INIT('h2)
	) name4727 (
		\g1092_reg/NET0131 ,
		\g1724_reg/NET0131 ,
		_w5907_
	);
	LUT2 #(
		.INIT('h4)
	) name4728 (
		\g1735_reg/NET0131 ,
		\g7961_pad ,
		_w5908_
	);
	LUT2 #(
		.INIT('h1)
	) name4729 (
		_w5906_,
		_w5907_,
		_w5909_
	);
	LUT2 #(
		.INIT('h4)
	) name4730 (
		_w5908_,
		_w5909_,
		_w5910_
	);
	LUT2 #(
		.INIT('h2)
	) name4731 (
		_w5905_,
		_w5910_,
		_w5911_
	);
	LUT2 #(
		.INIT('h2)
	) name4732 (
		\g1092_reg/NET0131 ,
		\g1739_reg/NET0131 ,
		_w5912_
	);
	LUT2 #(
		.INIT('h2)
	) name4733 (
		\g1088_reg/NET0131 ,
		\g1742_reg/NET0131 ,
		_w5913_
	);
	LUT2 #(
		.INIT('h4)
	) name4734 (
		\g1750_reg/NET0131 ,
		\g7961_pad ,
		_w5914_
	);
	LUT2 #(
		.INIT('h1)
	) name4735 (
		_w5912_,
		_w5913_,
		_w5915_
	);
	LUT2 #(
		.INIT('h4)
	) name4736 (
		_w5914_,
		_w5915_,
		_w5916_
	);
	LUT2 #(
		.INIT('h2)
	) name4737 (
		\g1088_reg/NET0131 ,
		\g1757_reg/NET0131 ,
		_w5917_
	);
	LUT2 #(
		.INIT('h4)
	) name4738 (
		\g1765_reg/NET0131 ,
		\g7961_pad ,
		_w5918_
	);
	LUT2 #(
		.INIT('h2)
	) name4739 (
		\g1092_reg/NET0131 ,
		\g1754_reg/NET0131 ,
		_w5919_
	);
	LUT2 #(
		.INIT('h1)
	) name4740 (
		_w5917_,
		_w5918_,
		_w5920_
	);
	LUT2 #(
		.INIT('h4)
	) name4741 (
		_w5919_,
		_w5920_,
		_w5921_
	);
	LUT2 #(
		.INIT('h4)
	) name4742 (
		_w5916_,
		_w5921_,
		_w5922_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		_w5911_,
		_w5922_,
		_w5923_
	);
	LUT2 #(
		.INIT('h1)
	) name4744 (
		\g3229_pad ,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h1)
	) name4745 (
		_w5910_,
		_w5922_,
		_w5925_
	);
	LUT2 #(
		.INIT('h2)
	) name4746 (
		_w5905_,
		_w5925_,
		_w5926_
	);
	LUT2 #(
		.INIT('h2)
	) name4747 (
		\g3229_pad ,
		_w5926_,
		_w5927_
	);
	LUT2 #(
		.INIT('h1)
	) name4748 (
		_w5924_,
		_w5927_,
		_w5928_
	);
	LUT2 #(
		.INIT('h8)
	) name4749 (
		_w5899_,
		_w5928_,
		_w5929_
	);
	LUT2 #(
		.INIT('h1)
	) name4750 (
		_w5900_,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h2)
	) name4751 (
		\g5657_pad ,
		_w5887_,
		_w5931_
	);
	LUT2 #(
		.INIT('h2)
	) name4752 (
		\g2650_reg/NET0131 ,
		_w5931_,
		_w5932_
	);
	LUT2 #(
		.INIT('h8)
	) name4753 (
		_w5895_,
		_w5931_,
		_w5933_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w5932_,
		_w5933_,
		_w5934_
	);
	LUT2 #(
		.INIT('h2)
	) name4755 (
		\g1018_reg/NET0131 ,
		_w5887_,
		_w5935_
	);
	LUT2 #(
		.INIT('h2)
	) name4756 (
		\g2651_reg/NET0131 ,
		_w5935_,
		_w5936_
	);
	LUT2 #(
		.INIT('h8)
	) name4757 (
		_w5895_,
		_w5935_,
		_w5937_
	);
	LUT2 #(
		.INIT('h1)
	) name4758 (
		_w5936_,
		_w5937_,
		_w5938_
	);
	LUT2 #(
		.INIT('h2)
	) name4759 (
		\g2655_reg/NET0131 ,
		_w5888_,
		_w5939_
	);
	LUT2 #(
		.INIT('h1)
	) name4760 (
		_w4317_,
		_w4336_,
		_w5940_
	);
	LUT2 #(
		.INIT('h1)
	) name4761 (
		\g3229_pad ,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h1)
	) name4762 (
		_w4321_,
		_w4332_,
		_w5942_
	);
	LUT2 #(
		.INIT('h2)
	) name4763 (
		\g3229_pad ,
		_w5942_,
		_w5943_
	);
	LUT2 #(
		.INIT('h1)
	) name4764 (
		_w5941_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h8)
	) name4765 (
		_w5888_,
		_w5944_,
		_w5945_
	);
	LUT2 #(
		.INIT('h1)
	) name4766 (
		_w5939_,
		_w5945_,
		_w5946_
	);
	LUT2 #(
		.INIT('h2)
	) name4767 (
		\g2656_reg/NET0131 ,
		_w5931_,
		_w5947_
	);
	LUT2 #(
		.INIT('h8)
	) name4768 (
		_w5931_,
		_w5944_,
		_w5948_
	);
	LUT2 #(
		.INIT('h1)
	) name4769 (
		_w5947_,
		_w5948_,
		_w5949_
	);
	LUT2 #(
		.INIT('h2)
	) name4770 (
		\g2657_reg/NET0131 ,
		_w5935_,
		_w5950_
	);
	LUT2 #(
		.INIT('h8)
	) name4771 (
		_w5935_,
		_w5944_,
		_w5951_
	);
	LUT2 #(
		.INIT('h1)
	) name4772 (
		_w5950_,
		_w5951_,
		_w5952_
	);
	LUT2 #(
		.INIT('h2)
	) name4773 (
		\g1088_reg/NET0131 ,
		_w5898_,
		_w5953_
	);
	LUT2 #(
		.INIT('h2)
	) name4774 (
		\g1727_reg/NET0131 ,
		_w5953_,
		_w5954_
	);
	LUT2 #(
		.INIT('h8)
	) name4775 (
		_w5928_,
		_w5953_,
		_w5955_
	);
	LUT2 #(
		.INIT('h1)
	) name4776 (
		_w5954_,
		_w5955_,
		_w5956_
	);
	LUT2 #(
		.INIT('h2)
	) name4777 (
		\g7961_pad ,
		_w5898_,
		_w5957_
	);
	LUT2 #(
		.INIT('h2)
	) name4778 (
		\g1735_reg/NET0131 ,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h8)
	) name4779 (
		_w5928_,
		_w5957_,
		_w5959_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		_w5958_,
		_w5959_,
		_w5960_
	);
	LUT2 #(
		.INIT('h2)
	) name4781 (
		\g3229_pad ,
		_w5910_,
		_w5961_
	);
	LUT2 #(
		.INIT('h4)
	) name4782 (
		\g3229_pad ,
		_w5910_,
		_w5962_
	);
	LUT2 #(
		.INIT('h1)
	) name4783 (
		_w5961_,
		_w5962_,
		_w5963_
	);
	LUT2 #(
		.INIT('h8)
	) name4784 (
		_w5916_,
		_w5963_,
		_w5964_
	);
	LUT2 #(
		.INIT('h8)
	) name4785 (
		_w5905_,
		_w5916_,
		_w5965_
	);
	LUT2 #(
		.INIT('h1)
	) name4786 (
		_w5963_,
		_w5965_,
		_w5966_
	);
	LUT2 #(
		.INIT('h1)
	) name4787 (
		_w5964_,
		_w5966_,
		_w5967_
	);
	LUT2 #(
		.INIT('h2)
	) name4788 (
		_w5899_,
		_w5967_,
		_w5968_
	);
	LUT2 #(
		.INIT('h2)
	) name4789 (
		\g1754_reg/NET0131 ,
		_w5899_,
		_w5969_
	);
	LUT2 #(
		.INIT('h1)
	) name4790 (
		_w5968_,
		_w5969_,
		_w5970_
	);
	LUT2 #(
		.INIT('h2)
	) name4791 (
		_w5953_,
		_w5967_,
		_w5971_
	);
	LUT2 #(
		.INIT('h2)
	) name4792 (
		\g1757_reg/NET0131 ,
		_w5953_,
		_w5972_
	);
	LUT2 #(
		.INIT('h1)
	) name4793 (
		_w5971_,
		_w5972_,
		_w5973_
	);
	LUT2 #(
		.INIT('h2)
	) name4794 (
		_w5957_,
		_w5967_,
		_w5974_
	);
	LUT2 #(
		.INIT('h2)
	) name4795 (
		\g1765_reg/NET0131 ,
		_w5957_,
		_w5975_
	);
	LUT2 #(
		.INIT('h1)
	) name4796 (
		_w5974_,
		_w5975_,
		_w5976_
	);
	LUT2 #(
		.INIT('h2)
	) name4797 (
		\g1033_reg/NET0131 ,
		_w5631_,
		_w5977_
	);
	LUT2 #(
		.INIT('h8)
	) name4798 (
		_w5631_,
		_w5875_,
		_w5978_
	);
	LUT2 #(
		.INIT('h1)
	) name4799 (
		_w5977_,
		_w5978_,
		_w5979_
	);
	LUT2 #(
		.INIT('h2)
	) name4800 (
		\g1041_reg/NET0131 ,
		_w5635_,
		_w5980_
	);
	LUT2 #(
		.INIT('h8)
	) name4801 (
		_w5635_,
		_w5875_,
		_w5981_
	);
	LUT2 #(
		.INIT('h1)
	) name4802 (
		_w5980_,
		_w5981_,
		_w5982_
	);
	LUT2 #(
		.INIT('h4)
	) name4803 (
		_w5473_,
		_w5484_,
		_w5983_
	);
	LUT2 #(
		.INIT('h2)
	) name4804 (
		_w5478_,
		_w5983_,
		_w5984_
	);
	LUT2 #(
		.INIT('h4)
	) name4805 (
		_w5478_,
		_w5983_,
		_w5985_
	);
	LUT2 #(
		.INIT('h1)
	) name4806 (
		_w5984_,
		_w5985_,
		_w5986_
	);
	LUT2 #(
		.INIT('h4)
	) name4807 (
		_w5548_,
		_w5559_,
		_w5987_
	);
	LUT2 #(
		.INIT('h2)
	) name4808 (
		_w5553_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h4)
	) name4809 (
		_w5553_,
		_w5987_,
		_w5989_
	);
	LUT2 #(
		.INIT('h1)
	) name4810 (
		_w5988_,
		_w5989_,
		_w5990_
	);
	LUT2 #(
		.INIT('h4)
	) name4811 (
		_w5497_,
		_w5519_,
		_w5991_
	);
	LUT2 #(
		.INIT('h2)
	) name4812 (
		_w5514_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h4)
	) name4813 (
		_w5514_,
		_w5991_,
		_w5993_
	);
	LUT2 #(
		.INIT('h1)
	) name4814 (
		_w5992_,
		_w5993_,
		_w5994_
	);
	LUT2 #(
		.INIT('h4)
	) name4815 (
		_w5572_,
		_w5594_,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name4816 (
		_w5589_,
		_w5995_,
		_w5996_
	);
	LUT2 #(
		.INIT('h4)
	) name4817 (
		_w5589_,
		_w5995_,
		_w5997_
	);
	LUT2 #(
		.INIT('h1)
	) name4818 (
		_w5996_,
		_w5997_,
		_w5998_
	);
	LUT2 #(
		.INIT('h4)
	) name4819 (
		_w5064_,
		_w5069_,
		_w5999_
	);
	LUT2 #(
		.INIT('h8)
	) name4820 (
		_w5193_,
		_w5999_,
		_w6000_
	);
	LUT2 #(
		.INIT('h4)
	) name4821 (
		_w5095_,
		_w5100_,
		_w6001_
	);
	LUT2 #(
		.INIT('h8)
	) name4822 (
		_w5201_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h4)
	) name4823 (
		_w5126_,
		_w5131_,
		_w6003_
	);
	LUT2 #(
		.INIT('h8)
	) name4824 (
		_w5209_,
		_w6003_,
		_w6004_
	);
	LUT2 #(
		.INIT('h2)
	) name4825 (
		_w5157_,
		_w5162_,
		_w6005_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		_w5217_,
		_w6005_,
		_w6006_
	);
	LUT2 #(
		.INIT('h8)
	) name4827 (
		\g3080_reg/NET0131 ,
		_w4132_,
		_w6007_
	);
	LUT2 #(
		.INIT('h8)
	) name4828 (
		\g3018_reg/NET0131 ,
		_w6007_,
		_w6008_
	);
	LUT2 #(
		.INIT('h8)
	) name4829 (
		\g3028_reg/NET0131 ,
		_w6008_,
		_w6009_
	);
	LUT2 #(
		.INIT('h1)
	) name4830 (
		\g3028_reg/NET0131 ,
		_w6008_,
		_w6010_
	);
	LUT2 #(
		.INIT('h4)
	) name4831 (
		\g3028_reg/NET0131 ,
		\g3032_reg/NET0131 ,
		_w6011_
	);
	LUT2 #(
		.INIT('h4)
	) name4832 (
		\g3036_reg/NET0131 ,
		_w6011_,
		_w6012_
	);
	LUT2 #(
		.INIT('h8)
	) name4833 (
		_w6008_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h1)
	) name4834 (
		\g3234_pad ,
		_w6013_,
		_w6014_
	);
	LUT2 #(
		.INIT('h1)
	) name4835 (
		_w6009_,
		_w6010_,
		_w6015_
	);
	LUT2 #(
		.INIT('h8)
	) name4836 (
		_w6014_,
		_w6015_,
		_w6016_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		\g1425_reg/NET0131 ,
		_w4584_,
		_w6017_
	);
	LUT2 #(
		.INIT('h1)
	) name4838 (
		_w5045_,
		_w6017_,
		_w6018_
	);
	LUT2 #(
		.INIT('h1)
	) name4839 (
		\g739_reg/NET0131 ,
		_w4700_,
		_w6019_
	);
	LUT2 #(
		.INIT('h1)
	) name4840 (
		_w5045_,
		_w6019_,
		_w6020_
	);
	LUT2 #(
		.INIT('h2)
	) name4841 (
		\g1563_reg/NET0131 ,
		_w5508_,
		_w6021_
	);
	LUT2 #(
		.INIT('h4)
	) name4842 (
		\g1563_reg/NET0131 ,
		_w5502_,
		_w6022_
	);
	LUT2 #(
		.INIT('h1)
	) name4843 (
		_w6021_,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h2)
	) name4844 (
		\g1563_reg/NET0131 ,
		_w5583_,
		_w6024_
	);
	LUT2 #(
		.INIT('h4)
	) name4845 (
		\g1563_reg/NET0131 ,
		_w5577_,
		_w6025_
	);
	LUT2 #(
		.INIT('h1)
	) name4846 (
		_w6024_,
		_w6025_,
		_w6026_
	);
	LUT2 #(
		.INIT('h1)
	) name4847 (
		\g3036_reg/NET0131 ,
		_w6009_,
		_w6027_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		\g3036_reg/NET0131 ,
		_w6009_,
		_w6028_
	);
	LUT2 #(
		.INIT('h2)
	) name4849 (
		_w6014_,
		_w6027_,
		_w6029_
	);
	LUT2 #(
		.INIT('h4)
	) name4850 (
		_w6028_,
		_w6029_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		\g3032_reg/NET0131 ,
		_w6028_,
		_w6031_
	);
	LUT2 #(
		.INIT('h8)
	) name4852 (
		\g3032_reg/NET0131 ,
		_w6028_,
		_w6032_
	);
	LUT2 #(
		.INIT('h2)
	) name4853 (
		_w6014_,
		_w6031_,
		_w6033_
	);
	LUT2 #(
		.INIT('h4)
	) name4854 (
		_w6032_,
		_w6033_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name4855 (
		\g1365_reg/NET0131 ,
		_w5053_,
		_w6035_
	);
	LUT2 #(
		.INIT('h1)
	) name4856 (
		_w5045_,
		_w5054_,
		_w6036_
	);
	LUT2 #(
		.INIT('h4)
	) name4857 (
		_w6035_,
		_w6036_,
		_w6037_
	);
	LUT2 #(
		.INIT('h1)
	) name4858 (
		\g3018_reg/NET0131 ,
		_w6007_,
		_w6038_
	);
	LUT2 #(
		.INIT('h1)
	) name4859 (
		_w6008_,
		_w6038_,
		_w6039_
	);
	LUT2 #(
		.INIT('h2)
	) name4860 (
		_w6014_,
		_w6039_,
		_w6040_
	);
	LUT2 #(
		.INIT('h1)
	) name4861 (
		\g3234_pad ,
		_w6007_,
		_w6041_
	);
	LUT2 #(
		.INIT('h8)
	) name4862 (
		\g2993_reg/NET0131 ,
		\g2998_reg/NET0131 ,
		_w6042_
	);
	LUT2 #(
		.INIT('h8)
	) name4863 (
		\g3080_reg/NET0131 ,
		_w6042_,
		_w6043_
	);
	LUT2 #(
		.INIT('h8)
	) name4864 (
		\g3006_reg/NET0131 ,
		_w6043_,
		_w6044_
	);
	LUT2 #(
		.INIT('h8)
	) name4865 (
		\g3002_reg/NET0131 ,
		_w6044_,
		_w6045_
	);
	LUT2 #(
		.INIT('h8)
	) name4866 (
		\g3013_reg/NET0131 ,
		_w6045_,
		_w6046_
	);
	LUT2 #(
		.INIT('h8)
	) name4867 (
		\g3010_reg/NET0131 ,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		\g3024_reg/NET0131 ,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h8)
	) name4869 (
		\g3024_reg/NET0131 ,
		_w6047_,
		_w6049_
	);
	LUT2 #(
		.INIT('h2)
	) name4870 (
		_w6041_,
		_w6048_,
		_w6050_
	);
	LUT2 #(
		.INIT('h4)
	) name4871 (
		_w6049_,
		_w6050_,
		_w6051_
	);
	LUT2 #(
		.INIT('h1)
	) name4872 (
		_w4738_,
		_w4782_,
		_w6052_
	);
	LUT2 #(
		.INIT('h1)
	) name4873 (
		\g3229_pad ,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h1)
	) name4874 (
		_w4763_,
		_w4787_,
		_w6054_
	);
	LUT2 #(
		.INIT('h2)
	) name4875 (
		\g3229_pad ,
		_w6054_,
		_w6055_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		_w6053_,
		_w6055_,
		_w6056_
	);
	LUT2 #(
		.INIT('h1)
	) name4877 (
		\g1430_reg/NET0131 ,
		_w5536_,
		_w6057_
	);
	LUT2 #(
		.INIT('h1)
	) name4878 (
		_w5527_,
		_w5537_,
		_w6058_
	);
	LUT2 #(
		.INIT('h4)
	) name4879 (
		_w6057_,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h1)
	) name4880 (
		\g1435_reg/NET0131 ,
		_w5535_,
		_w6060_
	);
	LUT2 #(
		.INIT('h1)
	) name4881 (
		_w5527_,
		_w5536_,
		_w6061_
	);
	LUT2 #(
		.INIT('h4)
	) name4882 (
		_w6060_,
		_w6061_,
		_w6062_
	);
	LUT2 #(
		.INIT('h1)
	) name4883 (
		\g1444_reg/NET0131 ,
		_w5533_,
		_w6063_
	);
	LUT2 #(
		.INIT('h1)
	) name4884 (
		_w5527_,
		_w5534_,
		_w6064_
	);
	LUT2 #(
		.INIT('h4)
	) name4885 (
		_w6063_,
		_w6064_,
		_w6065_
	);
	LUT2 #(
		.INIT('h1)
	) name4886 (
		\g1453_reg/NET0131 ,
		_w5531_,
		_w6066_
	);
	LUT2 #(
		.INIT('h1)
	) name4887 (
		_w5527_,
		_w5532_,
		_w6067_
	);
	LUT2 #(
		.INIT('h4)
	) name4888 (
		_w6066_,
		_w6067_,
		_w6068_
	);
	LUT2 #(
		.INIT('h1)
	) name4889 (
		\g1462_reg/NET0131 ,
		_w5529_,
		_w6069_
	);
	LUT2 #(
		.INIT('h1)
	) name4890 (
		_w5527_,
		_w5530_,
		_w6070_
	);
	LUT2 #(
		.INIT('h4)
	) name4891 (
		_w6069_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('h1)
	) name4892 (
		_w4889_,
		_w4899_,
		_w6072_
	);
	LUT2 #(
		.INIT('h1)
	) name4893 (
		\g3229_pad ,
		_w6072_,
		_w6073_
	);
	LUT2 #(
		.INIT('h1)
	) name4894 (
		_w4882_,
		_w4907_,
		_w6074_
	);
	LUT2 #(
		.INIT('h2)
	) name4895 (
		\g3229_pad ,
		_w6074_,
		_w6075_
	);
	LUT2 #(
		.INIT('h1)
	) name4896 (
		_w6073_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h1)
	) name4897 (
		\g1352_reg/NET0131 ,
		_w5052_,
		_w6077_
	);
	LUT2 #(
		.INIT('h1)
	) name4898 (
		_w5045_,
		_w5053_,
		_w6078_
	);
	LUT2 #(
		.INIT('h4)
	) name4899 (
		_w6077_,
		_w6078_,
		_w6079_
	);
	LUT2 #(
		.INIT('h4)
	) name4900 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		_w6080_
	);
	LUT2 #(
		.INIT('h8)
	) name4901 (
		\g2892_reg/NET0131 ,
		\g2903_reg/NET0131 ,
		_w6081_
	);
	LUT2 #(
		.INIT('h8)
	) name4902 (
		\g2908_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w6082_
	);
	LUT2 #(
		.INIT('h8)
	) name4903 (
		_w6081_,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h8)
	) name4904 (
		_w5259_,
		_w6080_,
		_w6084_
	);
	LUT2 #(
		.INIT('h8)
	) name4905 (
		_w6083_,
		_w6084_,
		_w6085_
	);
	LUT2 #(
		.INIT('h8)
	) name4906 (
		\g2912_reg/NET0131 ,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h4)
	) name4907 (
		\g2917_reg/NET0131 ,
		\g2920_reg/NET0131 ,
		_w6087_
	);
	LUT2 #(
		.INIT('h4)
	) name4908 (
		\g2924_reg/NET0131 ,
		_w6087_,
		_w6088_
	);
	LUT2 #(
		.INIT('h8)
	) name4909 (
		_w6086_,
		_w6088_,
		_w6089_
	);
	LUT2 #(
		.INIT('h1)
	) name4910 (
		\g2814_reg/NET0131 ,
		_w6089_,
		_w6090_
	);
	LUT2 #(
		.INIT('h8)
	) name4911 (
		\g2917_reg/NET0131 ,
		_w6086_,
		_w6091_
	);
	LUT2 #(
		.INIT('h8)
	) name4912 (
		\g2924_reg/NET0131 ,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('h1)
	) name4913 (
		\g2920_reg/NET0131 ,
		_w6092_,
		_w6093_
	);
	LUT2 #(
		.INIT('h8)
	) name4914 (
		\g2920_reg/NET0131 ,
		_w6092_,
		_w6094_
	);
	LUT2 #(
		.INIT('h2)
	) name4915 (
		_w6090_,
		_w6093_,
		_w6095_
	);
	LUT2 #(
		.INIT('h4)
	) name4916 (
		_w6094_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h1)
	) name4917 (
		\g2813_reg/NET0131 ,
		_w4528_,
		_w6097_
	);
	LUT2 #(
		.INIT('h1)
	) name4918 (
		_w5045_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h8)
	) name4919 (
		\g1024_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		_w6099_
	);
	LUT2 #(
		.INIT('h1)
	) name4920 (
		\g1423_reg/NET0131 ,
		_w4534_,
		_w6100_
	);
	LUT2 #(
		.INIT('h1)
	) name4921 (
		_w6099_,
		_w6100_,
		_w6101_
	);
	LUT2 #(
		.INIT('h8)
	) name4922 (
		\g1316_reg/NET0131 ,
		\g5657_pad ,
		_w6102_
	);
	LUT2 #(
		.INIT('h1)
	) name4923 (
		\g1424_reg/NET0131 ,
		_w4588_,
		_w6103_
	);
	LUT2 #(
		.INIT('h1)
	) name4924 (
		_w6102_,
		_w6103_,
		_w6104_
	);
	LUT2 #(
		.INIT('h1)
	) name4925 (
		\g737_reg/NET0131 ,
		_w4646_,
		_w6105_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		_w6099_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name4927 (
		\g2119_reg/NET0131 ,
		_w4704_,
		_w6107_
	);
	LUT2 #(
		.INIT('h1)
	) name4928 (
		_w5045_,
		_w6107_,
		_w6108_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		\g738_reg/NET0131 ,
		_w4696_,
		_w6109_
	);
	LUT2 #(
		.INIT('h1)
	) name4930 (
		_w6102_,
		_w6109_,
		_w6110_
	);
	LUT2 #(
		.INIT('h1)
	) name4931 (
		\g1439_reg/NET0131 ,
		_w5534_,
		_w6111_
	);
	LUT2 #(
		.INIT('h1)
	) name4932 (
		_w5527_,
		_w5535_,
		_w6112_
	);
	LUT2 #(
		.INIT('h4)
	) name4933 (
		_w6111_,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h1)
	) name4934 (
		\g1448_reg/NET0131 ,
		_w5532_,
		_w6114_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w5527_,
		_w5533_,
		_w6115_
	);
	LUT2 #(
		.INIT('h4)
	) name4936 (
		_w6114_,
		_w6115_,
		_w6116_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		\g1466_reg/NET0131 ,
		_w5528_,
		_w6117_
	);
	LUT2 #(
		.INIT('h1)
	) name4938 (
		_w5527_,
		_w5529_,
		_w6118_
	);
	LUT2 #(
		.INIT('h4)
	) name4939 (
		_w6117_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h1)
	) name4940 (
		\g1457_reg/NET0131 ,
		_w5530_,
		_w6120_
	);
	LUT2 #(
		.INIT('h1)
	) name4941 (
		_w5527_,
		_w5531_,
		_w6121_
	);
	LUT2 #(
		.INIT('h4)
	) name4942 (
		_w6120_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h1)
	) name4943 (
		\g1346_reg/NET0131 ,
		_w5050_,
		_w6123_
	);
	LUT2 #(
		.INIT('h1)
	) name4944 (
		_w5045_,
		_w5051_,
		_w6124_
	);
	LUT2 #(
		.INIT('h4)
	) name4945 (
		_w6123_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h1)
	) name4946 (
		\g1358_reg/NET0131 ,
		_w5051_,
		_w6126_
	);
	LUT2 #(
		.INIT('h1)
	) name4947 (
		_w5045_,
		_w5052_,
		_w6127_
	);
	LUT2 #(
		.INIT('h4)
	) name4948 (
		_w6126_,
		_w6127_,
		_w6128_
	);
	LUT2 #(
		.INIT('h4)
	) name4949 (
		\g3229_pad ,
		_w4329_,
		_w6129_
	);
	LUT2 #(
		.INIT('h8)
	) name4950 (
		\g3229_pad ,
		_w4377_,
		_w6130_
	);
	LUT2 #(
		.INIT('h1)
	) name4951 (
		_w4395_,
		_w6129_,
		_w6131_
	);
	LUT2 #(
		.INIT('h4)
	) name4952 (
		_w6130_,
		_w6131_,
		_w6132_
	);
	LUT2 #(
		.INIT('h8)
	) name4953 (
		_w5626_,
		_w5867_,
		_w6133_
	);
	LUT2 #(
		.INIT('h1)
	) name4954 (
		\g3229_pad ,
		_w4786_,
		_w6134_
	);
	LUT2 #(
		.INIT('h2)
	) name4955 (
		\g3229_pad ,
		_w4781_,
		_w6135_
	);
	LUT2 #(
		.INIT('h2)
	) name4956 (
		_w4749_,
		_w6134_,
		_w6136_
	);
	LUT2 #(
		.INIT('h4)
	) name4957 (
		_w6135_,
		_w6136_,
		_w6137_
	);
	LUT2 #(
		.INIT('h8)
	) name4958 (
		_w5696_,
		_w5717_,
		_w6138_
	);
	LUT2 #(
		.INIT('h1)
	) name4959 (
		\g3229_pad ,
		_w4906_,
		_w6139_
	);
	LUT2 #(
		.INIT('h2)
	) name4960 (
		\g3229_pad ,
		_w4893_,
		_w6140_
	);
	LUT2 #(
		.INIT('h2)
	) name4961 (
		_w4918_,
		_w6139_,
		_w6141_
	);
	LUT2 #(
		.INIT('h4)
	) name4962 (
		_w6140_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('h1)
	) name4963 (
		\g3229_pad ,
		_w4230_,
		_w6143_
	);
	LUT2 #(
		.INIT('h2)
	) name4964 (
		\g3229_pad ,
		_w4181_,
		_w6144_
	);
	LUT2 #(
		.INIT('h2)
	) name4965 (
		_w4177_,
		_w6143_,
		_w6145_
	);
	LUT2 #(
		.INIT('h4)
	) name4966 (
		_w6144_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h8)
	) name4967 (
		_w5822_,
		_w5849_,
		_w6147_
	);
	LUT2 #(
		.INIT('h1)
	) name4968 (
		\g3229_pad ,
		_w4320_,
		_w6148_
	);
	LUT2 #(
		.INIT('h2)
	) name4969 (
		\g3229_pad ,
		_w4335_,
		_w6149_
	);
	LUT2 #(
		.INIT('h2)
	) name4970 (
		_w4328_,
		_w6148_,
		_w6150_
	);
	LUT2 #(
		.INIT('h4)
	) name4971 (
		_w6149_,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h8)
	) name4972 (
		_w5921_,
		_w5964_,
		_w6152_
	);
	LUT2 #(
		.INIT('h1)
	) name4973 (
		\g1384_reg/NET0131 ,
		_w4534_,
		_w6153_
	);
	LUT2 #(
		.INIT('h8)
	) name4974 (
		_w4532_,
		_w5047_,
		_w6154_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w6153_,
		_w6154_,
		_w6155_
	);
	LUT2 #(
		.INIT('h2)
	) name4976 (
		\g1385_reg/NET0131 ,
		_w4588_,
		_w6156_
	);
	LUT2 #(
		.INIT('h4)
	) name4977 (
		\g1326_reg/NET0131 ,
		_w4588_,
		_w6157_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w6156_,
		_w6157_,
		_w6158_
	);
	LUT2 #(
		.INIT('h1)
	) name4979 (
		\g2811_reg/NET0131 ,
		_w4712_,
		_w6159_
	);
	LUT2 #(
		.INIT('h1)
	) name4980 (
		_w6099_,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h2)
	) name4981 (
		\g1386_reg/NET0131 ,
		_w4584_,
		_w6161_
	);
	LUT2 #(
		.INIT('h4)
	) name4982 (
		\g1326_reg/NET0131 ,
		_w4584_,
		_w6162_
	);
	LUT2 #(
		.INIT('h1)
	) name4983 (
		_w6161_,
		_w6162_,
		_w6163_
	);
	LUT2 #(
		.INIT('h1)
	) name4984 (
		\g2812_reg/NET0131 ,
		_w4478_,
		_w6164_
	);
	LUT2 #(
		.INIT('h1)
	) name4985 (
		_w6102_,
		_w6164_,
		_w6165_
	);
	LUT2 #(
		.INIT('h2)
	) name4986 (
		\g1387_reg/NET0131 ,
		_w4534_,
		_w6166_
	);
	LUT2 #(
		.INIT('h4)
	) name4987 (
		\g1319_reg/NET0131 ,
		_w4534_,
		_w6167_
	);
	LUT2 #(
		.INIT('h1)
	) name4988 (
		_w6166_,
		_w6167_,
		_w6168_
	);
	LUT2 #(
		.INIT('h2)
	) name4989 (
		\g1388_reg/NET0131 ,
		_w4588_,
		_w6169_
	);
	LUT2 #(
		.INIT('h4)
	) name4990 (
		\g1319_reg/NET0131 ,
		_w4588_,
		_w6170_
	);
	LUT2 #(
		.INIT('h1)
	) name4991 (
		_w6169_,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('h2)
	) name4992 (
		\g1389_reg/NET0131 ,
		_w4584_,
		_w6172_
	);
	LUT2 #(
		.INIT('h4)
	) name4993 (
		\g1319_reg/NET0131 ,
		_w4584_,
		_w6173_
	);
	LUT2 #(
		.INIT('h1)
	) name4994 (
		_w6172_,
		_w6173_,
		_w6174_
	);
	LUT2 #(
		.INIT('h2)
	) name4995 (
		\g1390_reg/NET0131 ,
		_w4534_,
		_w6175_
	);
	LUT2 #(
		.INIT('h4)
	) name4996 (
		\g1339_reg/NET0131 ,
		_w4534_,
		_w6176_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		_w6175_,
		_w6176_,
		_w6177_
	);
	LUT2 #(
		.INIT('h2)
	) name4998 (
		\g1391_reg/NET0131 ,
		_w4588_,
		_w6178_
	);
	LUT2 #(
		.INIT('h4)
	) name4999 (
		\g1339_reg/NET0131 ,
		_w4588_,
		_w6179_
	);
	LUT2 #(
		.INIT('h1)
	) name5000 (
		_w6178_,
		_w6179_,
		_w6180_
	);
	LUT2 #(
		.INIT('h2)
	) name5001 (
		\g1392_reg/NET0131 ,
		_w4584_,
		_w6181_
	);
	LUT2 #(
		.INIT('h4)
	) name5002 (
		\g1339_reg/NET0131 ,
		_w4584_,
		_w6182_
	);
	LUT2 #(
		.INIT('h1)
	) name5003 (
		_w6181_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h2)
	) name5004 (
		\g1393_reg/NET0131 ,
		_w4534_,
		_w6184_
	);
	LUT2 #(
		.INIT('h4)
	) name5005 (
		\g1332_reg/NET0131 ,
		_w4534_,
		_w6185_
	);
	LUT2 #(
		.INIT('h1)
	) name5006 (
		_w6184_,
		_w6185_,
		_w6186_
	);
	LUT2 #(
		.INIT('h2)
	) name5007 (
		\g1394_reg/NET0131 ,
		_w4588_,
		_w6187_
	);
	LUT2 #(
		.INIT('h4)
	) name5008 (
		\g1332_reg/NET0131 ,
		_w4588_,
		_w6188_
	);
	LUT2 #(
		.INIT('h1)
	) name5009 (
		_w6187_,
		_w6188_,
		_w6189_
	);
	LUT2 #(
		.INIT('h2)
	) name5010 (
		\g1395_reg/NET0131 ,
		_w4584_,
		_w6190_
	);
	LUT2 #(
		.INIT('h4)
	) name5011 (
		\g1332_reg/NET0131 ,
		_w4584_,
		_w6191_
	);
	LUT2 #(
		.INIT('h1)
	) name5012 (
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT2 #(
		.INIT('h2)
	) name5013 (
		\g1396_reg/NET0131 ,
		_w4534_,
		_w6193_
	);
	LUT2 #(
		.INIT('h4)
	) name5014 (
		\g1346_reg/NET0131 ,
		_w4534_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name5015 (
		_w6193_,
		_w6194_,
		_w6195_
	);
	LUT2 #(
		.INIT('h2)
	) name5016 (
		\g1397_reg/NET0131 ,
		_w4588_,
		_w6196_
	);
	LUT2 #(
		.INIT('h4)
	) name5017 (
		\g1346_reg/NET0131 ,
		_w4588_,
		_w6197_
	);
	LUT2 #(
		.INIT('h1)
	) name5018 (
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h2)
	) name5019 (
		\g1398_reg/NET0131 ,
		_w4584_,
		_w6199_
	);
	LUT2 #(
		.INIT('h4)
	) name5020 (
		\g1346_reg/NET0131 ,
		_w4584_,
		_w6200_
	);
	LUT2 #(
		.INIT('h1)
	) name5021 (
		_w6199_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h2)
	) name5022 (
		\g1399_reg/NET0131 ,
		_w4534_,
		_w6202_
	);
	LUT2 #(
		.INIT('h4)
	) name5023 (
		\g1358_reg/NET0131 ,
		_w4534_,
		_w6203_
	);
	LUT2 #(
		.INIT('h1)
	) name5024 (
		_w6202_,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h2)
	) name5025 (
		\g1400_reg/NET0131 ,
		_w4588_,
		_w6205_
	);
	LUT2 #(
		.INIT('h4)
	) name5026 (
		\g1358_reg/NET0131 ,
		_w4588_,
		_w6206_
	);
	LUT2 #(
		.INIT('h1)
	) name5027 (
		_w6205_,
		_w6206_,
		_w6207_
	);
	LUT2 #(
		.INIT('h2)
	) name5028 (
		\g1401_reg/NET0131 ,
		_w4584_,
		_w6208_
	);
	LUT2 #(
		.INIT('h4)
	) name5029 (
		\g1358_reg/NET0131 ,
		_w4584_,
		_w6209_
	);
	LUT2 #(
		.INIT('h1)
	) name5030 (
		_w6208_,
		_w6209_,
		_w6210_
	);
	LUT2 #(
		.INIT('h2)
	) name5031 (
		\g1402_reg/NET0131 ,
		_w4534_,
		_w6211_
	);
	LUT2 #(
		.INIT('h4)
	) name5032 (
		\g1352_reg/NET0131 ,
		_w4534_,
		_w6212_
	);
	LUT2 #(
		.INIT('h1)
	) name5033 (
		_w6211_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h2)
	) name5034 (
		\g1403_reg/NET0131 ,
		_w4588_,
		_w6214_
	);
	LUT2 #(
		.INIT('h4)
	) name5035 (
		\g1352_reg/NET0131 ,
		_w4588_,
		_w6215_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		_w6214_,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h2)
	) name5037 (
		\g1404_reg/NET0131 ,
		_w4584_,
		_w6217_
	);
	LUT2 #(
		.INIT('h4)
	) name5038 (
		\g1352_reg/NET0131 ,
		_w4584_,
		_w6218_
	);
	LUT2 #(
		.INIT('h1)
	) name5039 (
		_w6217_,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h2)
	) name5040 (
		\g1405_reg/NET0131 ,
		_w4534_,
		_w6220_
	);
	LUT2 #(
		.INIT('h4)
	) name5041 (
		\g1365_reg/NET0131 ,
		_w4534_,
		_w6221_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		_w6220_,
		_w6221_,
		_w6222_
	);
	LUT2 #(
		.INIT('h2)
	) name5043 (
		\g1406_reg/NET0131 ,
		_w4588_,
		_w6223_
	);
	LUT2 #(
		.INIT('h4)
	) name5044 (
		\g1365_reg/NET0131 ,
		_w4588_,
		_w6224_
	);
	LUT2 #(
		.INIT('h1)
	) name5045 (
		_w6223_,
		_w6224_,
		_w6225_
	);
	LUT2 #(
		.INIT('h2)
	) name5046 (
		\g1407_reg/NET0131 ,
		_w4584_,
		_w6226_
	);
	LUT2 #(
		.INIT('h4)
	) name5047 (
		\g1365_reg/NET0131 ,
		_w4584_,
		_w6227_
	);
	LUT2 #(
		.INIT('h1)
	) name5048 (
		_w6226_,
		_w6227_,
		_w6228_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		\g1408_reg/NET0131 ,
		_w4534_,
		_w6229_
	);
	LUT2 #(
		.INIT('h4)
	) name5050 (
		\g1372_reg/NET0131 ,
		_w4534_,
		_w6230_
	);
	LUT2 #(
		.INIT('h1)
	) name5051 (
		_w6229_,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h2)
	) name5052 (
		\g1409_reg/NET0131 ,
		_w4588_,
		_w6232_
	);
	LUT2 #(
		.INIT('h4)
	) name5053 (
		\g1372_reg/NET0131 ,
		_w4588_,
		_w6233_
	);
	LUT2 #(
		.INIT('h1)
	) name5054 (
		_w6232_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h2)
	) name5055 (
		\g1410_reg/NET0131 ,
		_w4584_,
		_w6235_
	);
	LUT2 #(
		.INIT('h4)
	) name5056 (
		\g1372_reg/NET0131 ,
		_w4584_,
		_w6236_
	);
	LUT2 #(
		.INIT('h1)
	) name5057 (
		_w6235_,
		_w6236_,
		_w6237_
	);
	LUT2 #(
		.INIT('h2)
	) name5058 (
		\g1411_reg/NET0131 ,
		_w4534_,
		_w6238_
	);
	LUT2 #(
		.INIT('h4)
	) name5059 (
		\g1378_reg/NET0131 ,
		_w4534_,
		_w6239_
	);
	LUT2 #(
		.INIT('h1)
	) name5060 (
		_w6238_,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h2)
	) name5061 (
		\g1412_reg/NET0131 ,
		_w4588_,
		_w6241_
	);
	LUT2 #(
		.INIT('h4)
	) name5062 (
		\g1378_reg/NET0131 ,
		_w4588_,
		_w6242_
	);
	LUT2 #(
		.INIT('h1)
	) name5063 (
		_w6241_,
		_w6242_,
		_w6243_
	);
	LUT2 #(
		.INIT('h2)
	) name5064 (
		\g1413_reg/NET0131 ,
		_w4584_,
		_w6244_
	);
	LUT2 #(
		.INIT('h4)
	) name5065 (
		\g1378_reg/NET0131 ,
		_w4584_,
		_w6245_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w6244_,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h2)
	) name5067 (
		\g2232_reg/NET0131 ,
		_w5023_,
		_w6247_
	);
	LUT2 #(
		.INIT('h4)
	) name5068 (
		\g2200_reg/NET0131 ,
		_w5023_,
		_w6248_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w6247_,
		_w6248_,
		_w6249_
	);
	LUT2 #(
		.INIT('h2)
	) name5070 (
		\g1511_reg/NET0131 ,
		_w5023_,
		_w6250_
	);
	LUT2 #(
		.INIT('h4)
	) name5071 (
		\g1471_reg/NET0131 ,
		_w5023_,
		_w6251_
	);
	LUT2 #(
		.INIT('h1)
	) name5072 (
		_w6250_,
		_w6251_,
		_w6252_
	);
	LUT2 #(
		.INIT('h2)
	) name5073 (
		\g1512_reg/NET0131 ,
		_w5027_,
		_w6253_
	);
	LUT2 #(
		.INIT('h4)
	) name5074 (
		\g1471_reg/NET0131 ,
		_w5027_,
		_w6254_
	);
	LUT2 #(
		.INIT('h1)
	) name5075 (
		_w6253_,
		_w6254_,
		_w6255_
	);
	LUT2 #(
		.INIT('h2)
	) name5076 (
		\g1513_reg/NET0131 ,
		_w5029_,
		_w6256_
	);
	LUT2 #(
		.INIT('h4)
	) name5077 (
		\g1471_reg/NET0131 ,
		_w5029_,
		_w6257_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		_w6256_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h2)
	) name5079 (
		\g1529_reg/NET0131 ,
		_w5023_,
		_w6259_
	);
	LUT2 #(
		.INIT('h4)
	) name5080 (
		\g1491_reg/NET0131 ,
		_w5023_,
		_w6260_
	);
	LUT2 #(
		.INIT('h1)
	) name5081 (
		_w6259_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('h2)
	) name5082 (
		\g1531_reg/NET0131 ,
		_w5029_,
		_w6262_
	);
	LUT2 #(
		.INIT('h4)
	) name5083 (
		\g1491_reg/NET0131 ,
		_w5029_,
		_w6263_
	);
	LUT2 #(
		.INIT('h1)
	) name5084 (
		_w6262_,
		_w6263_,
		_w6264_
	);
	LUT2 #(
		.INIT('h2)
	) name5085 (
		\g1530_reg/NET0131 ,
		_w5027_,
		_w6265_
	);
	LUT2 #(
		.INIT('h4)
	) name5086 (
		\g1491_reg/NET0131 ,
		_w5027_,
		_w6266_
	);
	LUT2 #(
		.INIT('h1)
	) name5087 (
		_w6265_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h2)
	) name5088 (
		\g1532_reg/NET0131 ,
		_w5023_,
		_w6268_
	);
	LUT2 #(
		.INIT('h4)
	) name5089 (
		\g1496_reg/NET0131 ,
		_w5023_,
		_w6269_
	);
	LUT2 #(
		.INIT('h1)
	) name5090 (
		_w6268_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h2)
	) name5091 (
		\g1533_reg/NET0131 ,
		_w5027_,
		_w6271_
	);
	LUT2 #(
		.INIT('h4)
	) name5092 (
		\g1496_reg/NET0131 ,
		_w5027_,
		_w6272_
	);
	LUT2 #(
		.INIT('h1)
	) name5093 (
		_w6271_,
		_w6272_,
		_w6273_
	);
	LUT2 #(
		.INIT('h2)
	) name5094 (
		\g1534_reg/NET0131 ,
		_w5029_,
		_w6274_
	);
	LUT2 #(
		.INIT('h4)
	) name5095 (
		\g1496_reg/NET0131 ,
		_w5029_,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		_w6274_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h2)
	) name5097 (
		\g1535_reg/NET0131 ,
		_w5023_,
		_w6277_
	);
	LUT2 #(
		.INIT('h4)
	) name5098 (
		\g1501_reg/NET0131 ,
		_w5023_,
		_w6278_
	);
	LUT2 #(
		.INIT('h1)
	) name5099 (
		_w6277_,
		_w6278_,
		_w6279_
	);
	LUT2 #(
		.INIT('h2)
	) name5100 (
		\g1536_reg/NET0131 ,
		_w5027_,
		_w6280_
	);
	LUT2 #(
		.INIT('h4)
	) name5101 (
		\g1501_reg/NET0131 ,
		_w5027_,
		_w6281_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		_w6280_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h2)
	) name5103 (
		\g1537_reg/NET0131 ,
		_w5029_,
		_w6283_
	);
	LUT2 #(
		.INIT('h4)
	) name5104 (
		\g1501_reg/NET0131 ,
		_w5029_,
		_w6284_
	);
	LUT2 #(
		.INIT('h1)
	) name5105 (
		_w6283_,
		_w6284_,
		_w6285_
	);
	LUT2 #(
		.INIT('h2)
	) name5106 (
		\g1538_reg/NET0131 ,
		_w5023_,
		_w6286_
	);
	LUT2 #(
		.INIT('h4)
	) name5107 (
		\g1506_reg/NET0131 ,
		_w5023_,
		_w6287_
	);
	LUT2 #(
		.INIT('h1)
	) name5108 (
		_w6286_,
		_w6287_,
		_w6288_
	);
	LUT2 #(
		.INIT('h2)
	) name5109 (
		\g1539_reg/NET0131 ,
		_w5027_,
		_w6289_
	);
	LUT2 #(
		.INIT('h4)
	) name5110 (
		\g1506_reg/NET0131 ,
		_w5027_,
		_w6290_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w6289_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h2)
	) name5112 (
		\g698_reg/NET0131 ,
		_w4646_,
		_w6292_
	);
	LUT2 #(
		.INIT('h4)
	) name5113 (
		\g1326_reg/NET0131 ,
		_w4646_,
		_w6293_
	);
	LUT2 #(
		.INIT('h1)
	) name5114 (
		_w6292_,
		_w6293_,
		_w6294_
	);
	LUT2 #(
		.INIT('h2)
	) name5115 (
		\g699_reg/NET0131 ,
		_w4696_,
		_w6295_
	);
	LUT2 #(
		.INIT('h4)
	) name5116 (
		\g1326_reg/NET0131 ,
		_w4696_,
		_w6296_
	);
	LUT2 #(
		.INIT('h1)
	) name5117 (
		_w6295_,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h2)
	) name5118 (
		\g700_reg/NET0131 ,
		_w4700_,
		_w6298_
	);
	LUT2 #(
		.INIT('h4)
	) name5119 (
		\g1326_reg/NET0131 ,
		_w4700_,
		_w6299_
	);
	LUT2 #(
		.INIT('h1)
	) name5120 (
		_w6298_,
		_w6299_,
		_w6300_
	);
	LUT2 #(
		.INIT('h2)
	) name5121 (
		\g701_reg/NET0131 ,
		_w4646_,
		_w6301_
	);
	LUT2 #(
		.INIT('h4)
	) name5122 (
		\g1319_reg/NET0131 ,
		_w4646_,
		_w6302_
	);
	LUT2 #(
		.INIT('h1)
	) name5123 (
		_w6301_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h2)
	) name5124 (
		\g702_reg/NET0131 ,
		_w4696_,
		_w6304_
	);
	LUT2 #(
		.INIT('h4)
	) name5125 (
		\g1319_reg/NET0131 ,
		_w4696_,
		_w6305_
	);
	LUT2 #(
		.INIT('h1)
	) name5126 (
		_w6304_,
		_w6305_,
		_w6306_
	);
	LUT2 #(
		.INIT('h2)
	) name5127 (
		\g703_reg/NET0131 ,
		_w4700_,
		_w6307_
	);
	LUT2 #(
		.INIT('h4)
	) name5128 (
		\g1319_reg/NET0131 ,
		_w4700_,
		_w6308_
	);
	LUT2 #(
		.INIT('h1)
	) name5129 (
		_w6307_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('h2)
	) name5130 (
		\g704_reg/NET0131 ,
		_w4646_,
		_w6310_
	);
	LUT2 #(
		.INIT('h4)
	) name5131 (
		\g1339_reg/NET0131 ,
		_w4646_,
		_w6311_
	);
	LUT2 #(
		.INIT('h1)
	) name5132 (
		_w6310_,
		_w6311_,
		_w6312_
	);
	LUT2 #(
		.INIT('h2)
	) name5133 (
		\g705_reg/NET0131 ,
		_w4696_,
		_w6313_
	);
	LUT2 #(
		.INIT('h4)
	) name5134 (
		\g1339_reg/NET0131 ,
		_w4696_,
		_w6314_
	);
	LUT2 #(
		.INIT('h1)
	) name5135 (
		_w6313_,
		_w6314_,
		_w6315_
	);
	LUT2 #(
		.INIT('h2)
	) name5136 (
		\g706_reg/NET0131 ,
		_w4700_,
		_w6316_
	);
	LUT2 #(
		.INIT('h4)
	) name5137 (
		\g1339_reg/NET0131 ,
		_w4700_,
		_w6317_
	);
	LUT2 #(
		.INIT('h1)
	) name5138 (
		_w6316_,
		_w6317_,
		_w6318_
	);
	LUT2 #(
		.INIT('h2)
	) name5139 (
		\g707_reg/NET0131 ,
		_w4646_,
		_w6319_
	);
	LUT2 #(
		.INIT('h4)
	) name5140 (
		\g1332_reg/NET0131 ,
		_w4646_,
		_w6320_
	);
	LUT2 #(
		.INIT('h1)
	) name5141 (
		_w6319_,
		_w6320_,
		_w6321_
	);
	LUT2 #(
		.INIT('h2)
	) name5142 (
		\g708_reg/NET0131 ,
		_w4696_,
		_w6322_
	);
	LUT2 #(
		.INIT('h4)
	) name5143 (
		\g1332_reg/NET0131 ,
		_w4696_,
		_w6323_
	);
	LUT2 #(
		.INIT('h1)
	) name5144 (
		_w6322_,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h2)
	) name5145 (
		\g709_reg/NET0131 ,
		_w4700_,
		_w6325_
	);
	LUT2 #(
		.INIT('h4)
	) name5146 (
		\g1332_reg/NET0131 ,
		_w4700_,
		_w6326_
	);
	LUT2 #(
		.INIT('h1)
	) name5147 (
		_w6325_,
		_w6326_,
		_w6327_
	);
	LUT2 #(
		.INIT('h2)
	) name5148 (
		\g710_reg/NET0131 ,
		_w4646_,
		_w6328_
	);
	LUT2 #(
		.INIT('h4)
	) name5149 (
		\g1346_reg/NET0131 ,
		_w4646_,
		_w6329_
	);
	LUT2 #(
		.INIT('h1)
	) name5150 (
		_w6328_,
		_w6329_,
		_w6330_
	);
	LUT2 #(
		.INIT('h2)
	) name5151 (
		\g711_reg/NET0131 ,
		_w4696_,
		_w6331_
	);
	LUT2 #(
		.INIT('h4)
	) name5152 (
		\g1346_reg/NET0131 ,
		_w4696_,
		_w6332_
	);
	LUT2 #(
		.INIT('h1)
	) name5153 (
		_w6331_,
		_w6332_,
		_w6333_
	);
	LUT2 #(
		.INIT('h2)
	) name5154 (
		\g712_reg/NET0131 ,
		_w4700_,
		_w6334_
	);
	LUT2 #(
		.INIT('h4)
	) name5155 (
		\g1346_reg/NET0131 ,
		_w4700_,
		_w6335_
	);
	LUT2 #(
		.INIT('h1)
	) name5156 (
		_w6334_,
		_w6335_,
		_w6336_
	);
	LUT2 #(
		.INIT('h2)
	) name5157 (
		\g713_reg/NET0131 ,
		_w4646_,
		_w6337_
	);
	LUT2 #(
		.INIT('h4)
	) name5158 (
		\g1358_reg/NET0131 ,
		_w4646_,
		_w6338_
	);
	LUT2 #(
		.INIT('h1)
	) name5159 (
		_w6337_,
		_w6338_,
		_w6339_
	);
	LUT2 #(
		.INIT('h2)
	) name5160 (
		\g714_reg/NET0131 ,
		_w4696_,
		_w6340_
	);
	LUT2 #(
		.INIT('h4)
	) name5161 (
		\g1358_reg/NET0131 ,
		_w4696_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name5162 (
		_w6340_,
		_w6341_,
		_w6342_
	);
	LUT2 #(
		.INIT('h2)
	) name5163 (
		\g715_reg/NET0131 ,
		_w4700_,
		_w6343_
	);
	LUT2 #(
		.INIT('h4)
	) name5164 (
		\g1358_reg/NET0131 ,
		_w4700_,
		_w6344_
	);
	LUT2 #(
		.INIT('h1)
	) name5165 (
		_w6343_,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h2)
	) name5166 (
		\g716_reg/NET0131 ,
		_w4646_,
		_w6346_
	);
	LUT2 #(
		.INIT('h4)
	) name5167 (
		\g1352_reg/NET0131 ,
		_w4646_,
		_w6347_
	);
	LUT2 #(
		.INIT('h1)
	) name5168 (
		_w6346_,
		_w6347_,
		_w6348_
	);
	LUT2 #(
		.INIT('h2)
	) name5169 (
		\g717_reg/NET0131 ,
		_w4696_,
		_w6349_
	);
	LUT2 #(
		.INIT('h4)
	) name5170 (
		\g1352_reg/NET0131 ,
		_w4696_,
		_w6350_
	);
	LUT2 #(
		.INIT('h1)
	) name5171 (
		_w6349_,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('h2)
	) name5172 (
		\g718_reg/NET0131 ,
		_w4700_,
		_w6352_
	);
	LUT2 #(
		.INIT('h4)
	) name5173 (
		\g1352_reg/NET0131 ,
		_w4700_,
		_w6353_
	);
	LUT2 #(
		.INIT('h1)
	) name5174 (
		_w6352_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h2)
	) name5175 (
		\g719_reg/NET0131 ,
		_w4646_,
		_w6355_
	);
	LUT2 #(
		.INIT('h4)
	) name5176 (
		\g1365_reg/NET0131 ,
		_w4646_,
		_w6356_
	);
	LUT2 #(
		.INIT('h1)
	) name5177 (
		_w6355_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h2)
	) name5178 (
		\g720_reg/NET0131 ,
		_w4696_,
		_w6358_
	);
	LUT2 #(
		.INIT('h4)
	) name5179 (
		\g1365_reg/NET0131 ,
		_w4696_,
		_w6359_
	);
	LUT2 #(
		.INIT('h1)
	) name5180 (
		_w6358_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h2)
	) name5181 (
		\g721_reg/NET0131 ,
		_w4700_,
		_w6361_
	);
	LUT2 #(
		.INIT('h4)
	) name5182 (
		\g1365_reg/NET0131 ,
		_w4700_,
		_w6362_
	);
	LUT2 #(
		.INIT('h1)
	) name5183 (
		_w6361_,
		_w6362_,
		_w6363_
	);
	LUT2 #(
		.INIT('h2)
	) name5184 (
		\g722_reg/NET0131 ,
		_w4646_,
		_w6364_
	);
	LUT2 #(
		.INIT('h4)
	) name5185 (
		\g1372_reg/NET0131 ,
		_w4646_,
		_w6365_
	);
	LUT2 #(
		.INIT('h1)
	) name5186 (
		_w6364_,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h2)
	) name5187 (
		\g723_reg/NET0131 ,
		_w4696_,
		_w6367_
	);
	LUT2 #(
		.INIT('h4)
	) name5188 (
		\g1372_reg/NET0131 ,
		_w4696_,
		_w6368_
	);
	LUT2 #(
		.INIT('h1)
	) name5189 (
		_w6367_,
		_w6368_,
		_w6369_
	);
	LUT2 #(
		.INIT('h2)
	) name5190 (
		\g724_reg/NET0131 ,
		_w4700_,
		_w6370_
	);
	LUT2 #(
		.INIT('h4)
	) name5191 (
		\g1372_reg/NET0131 ,
		_w4700_,
		_w6371_
	);
	LUT2 #(
		.INIT('h1)
	) name5192 (
		_w6370_,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('h2)
	) name5193 (
		\g725_reg/NET0131 ,
		_w4646_,
		_w6373_
	);
	LUT2 #(
		.INIT('h4)
	) name5194 (
		\g1378_reg/NET0131 ,
		_w4646_,
		_w6374_
	);
	LUT2 #(
		.INIT('h1)
	) name5195 (
		_w6373_,
		_w6374_,
		_w6375_
	);
	LUT2 #(
		.INIT('h2)
	) name5196 (
		\g726_reg/NET0131 ,
		_w4696_,
		_w6376_
	);
	LUT2 #(
		.INIT('h4)
	) name5197 (
		\g1378_reg/NET0131 ,
		_w4696_,
		_w6377_
	);
	LUT2 #(
		.INIT('h1)
	) name5198 (
		_w6376_,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h2)
	) name5199 (
		\g727_reg/NET0131 ,
		_w4700_,
		_w6379_
	);
	LUT2 #(
		.INIT('h4)
	) name5200 (
		\g1378_reg/NET0131 ,
		_w4700_,
		_w6380_
	);
	LUT2 #(
		.INIT('h1)
	) name5201 (
		_w6379_,
		_w6380_,
		_w6381_
	);
	LUT2 #(
		.INIT('h1)
	) name5202 (
		\g2118_reg/NET0131 ,
		_w4708_,
		_w6382_
	);
	LUT2 #(
		.INIT('h1)
	) name5203 (
		_w6102_,
		_w6382_,
		_w6383_
	);
	LUT2 #(
		.INIT('h2)
	) name5204 (
		\g2229_reg/NET0131 ,
		_w5023_,
		_w6384_
	);
	LUT2 #(
		.INIT('h4)
	) name5205 (
		\g2195_reg/NET0131 ,
		_w5023_,
		_w6385_
	);
	LUT2 #(
		.INIT('h1)
	) name5206 (
		_w6384_,
		_w6385_,
		_w6386_
	);
	LUT2 #(
		.INIT('h2)
	) name5207 (
		\g1540_reg/NET0131 ,
		_w5029_,
		_w6387_
	);
	LUT2 #(
		.INIT('h4)
	) name5208 (
		\g1506_reg/NET0131 ,
		_w5029_,
		_w6388_
	);
	LUT2 #(
		.INIT('h1)
	) name5209 (
		_w6387_,
		_w6388_,
		_w6389_
	);
	LUT2 #(
		.INIT('h1)
	) name5210 (
		\g2117_reg/NET0131 ,
		_w4594_,
		_w6390_
	);
	LUT2 #(
		.INIT('h1)
	) name5211 (
		_w6099_,
		_w6390_,
		_w6391_
	);
	LUT2 #(
		.INIT('h2)
	) name5212 (
		\g7961_pad ,
		_w2837_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name5213 (
		\g1846_reg/NET0131 ,
		\g7961_pad ,
		_w6393_
	);
	LUT2 #(
		.INIT('h1)
	) name5214 (
		_w6392_,
		_w6393_,
		_w6394_
	);
	LUT2 #(
		.INIT('h2)
	) name5215 (
		\g1092_reg/NET0131 ,
		_w2837_,
		_w6395_
	);
	LUT2 #(
		.INIT('h1)
	) name5216 (
		\g1092_reg/NET0131 ,
		\g1849_reg/NET0131 ,
		_w6396_
	);
	LUT2 #(
		.INIT('h1)
	) name5217 (
		_w6395_,
		_w6396_,
		_w6397_
	);
	LUT2 #(
		.INIT('h2)
	) name5218 (
		\g1088_reg/NET0131 ,
		_w2837_,
		_w6398_
	);
	LUT2 #(
		.INIT('h1)
	) name5219 (
		\g1088_reg/NET0131 ,
		\g1852_reg/NET0131 ,
		_w6399_
	);
	LUT2 #(
		.INIT('h1)
	) name5220 (
		_w6398_,
		_w6399_,
		_w6400_
	);
	LUT2 #(
		.INIT('h2)
	) name5221 (
		\g7961_pad ,
		_w5672_,
		_w6401_
	);
	LUT2 #(
		.INIT('h1)
	) name5222 (
		\g465_reg/NET0131 ,
		\g7961_pad ,
		_w6402_
	);
	LUT2 #(
		.INIT('h1)
	) name5223 (
		_w6401_,
		_w6402_,
		_w6403_
	);
	LUT2 #(
		.INIT('h2)
	) name5224 (
		\g1092_reg/NET0131 ,
		_w5672_,
		_w6404_
	);
	LUT2 #(
		.INIT('h1)
	) name5225 (
		\g1092_reg/NET0131 ,
		\g468_reg/NET0131 ,
		_w6405_
	);
	LUT2 #(
		.INIT('h1)
	) name5226 (
		_w6404_,
		_w6405_,
		_w6406_
	);
	LUT2 #(
		.INIT('h2)
	) name5227 (
		\g1088_reg/NET0131 ,
		_w5672_,
		_w6407_
	);
	LUT2 #(
		.INIT('h1)
	) name5228 (
		\g1088_reg/NET0131 ,
		\g471_reg/NET0131 ,
		_w6408_
	);
	LUT2 #(
		.INIT('h1)
	) name5229 (
		_w6407_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h2)
	) name5230 (
		\g7961_pad ,
		_w1310_,
		_w6410_
	);
	LUT2 #(
		.INIT('h1)
	) name5231 (
		\g2540_reg/NET0131 ,
		\g7961_pad ,
		_w6411_
	);
	LUT2 #(
		.INIT('h1)
	) name5232 (
		_w6410_,
		_w6411_,
		_w6412_
	);
	LUT2 #(
		.INIT('h2)
	) name5233 (
		\g1092_reg/NET0131 ,
		_w1310_,
		_w6413_
	);
	LUT2 #(
		.INIT('h1)
	) name5234 (
		\g1092_reg/NET0131 ,
		\g2543_reg/NET0131 ,
		_w6414_
	);
	LUT2 #(
		.INIT('h1)
	) name5235 (
		_w6413_,
		_w6414_,
		_w6415_
	);
	LUT2 #(
		.INIT('h2)
	) name5236 (
		\g1088_reg/NET0131 ,
		_w1310_,
		_w6416_
	);
	LUT2 #(
		.INIT('h1)
	) name5237 (
		\g1088_reg/NET0131 ,
		\g2546_reg/NET0131 ,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name5238 (
		_w6416_,
		_w6417_,
		_w6418_
	);
	LUT2 #(
		.INIT('h2)
	) name5239 (
		\g847_reg/NET0131 ,
		_w5023_,
		_w6419_
	);
	LUT2 #(
		.INIT('h8)
	) name5240 (
		_w2356_,
		_w5023_,
		_w6420_
	);
	LUT2 #(
		.INIT('h1)
	) name5241 (
		_w6419_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h2)
	) name5242 (
		\g848_reg/NET0131 ,
		_w5027_,
		_w6422_
	);
	LUT2 #(
		.INIT('h8)
	) name5243 (
		_w2356_,
		_w5027_,
		_w6423_
	);
	LUT2 #(
		.INIT('h1)
	) name5244 (
		_w6422_,
		_w6423_,
		_w6424_
	);
	LUT2 #(
		.INIT('h2)
	) name5245 (
		\g849_reg/NET0131 ,
		_w5029_,
		_w6425_
	);
	LUT2 #(
		.INIT('h8)
	) name5246 (
		_w2356_,
		_w5029_,
		_w6426_
	);
	LUT2 #(
		.INIT('h1)
	) name5247 (
		_w6425_,
		_w6426_,
		_w6427_
	);
	LUT2 #(
		.INIT('h2)
	) name5248 (
		\g850_reg/NET0131 ,
		_w5023_,
		_w6428_
	);
	LUT2 #(
		.INIT('h8)
	) name5249 (
		_w2298_,
		_w5023_,
		_w6429_
	);
	LUT2 #(
		.INIT('h1)
	) name5250 (
		_w6428_,
		_w6429_,
		_w6430_
	);
	LUT2 #(
		.INIT('h2)
	) name5251 (
		\g851_reg/NET0131 ,
		_w5027_,
		_w6431_
	);
	LUT2 #(
		.INIT('h8)
	) name5252 (
		_w2298_,
		_w5027_,
		_w6432_
	);
	LUT2 #(
		.INIT('h1)
	) name5253 (
		_w6431_,
		_w6432_,
		_w6433_
	);
	LUT2 #(
		.INIT('h2)
	) name5254 (
		\g852_reg/NET0131 ,
		_w5029_,
		_w6434_
	);
	LUT2 #(
		.INIT('h8)
	) name5255 (
		_w2298_,
		_w5029_,
		_w6435_
	);
	LUT2 #(
		.INIT('h1)
	) name5256 (
		_w6434_,
		_w6435_,
		_w6436_
	);
	LUT2 #(
		.INIT('h2)
	) name5257 (
		\g159_reg/NET0131 ,
		_w5023_,
		_w6437_
	);
	LUT2 #(
		.INIT('h8)
	) name5258 (
		_w2047_,
		_w5023_,
		_w6438_
	);
	LUT2 #(
		.INIT('h1)
	) name5259 (
		_w6437_,
		_w6438_,
		_w6439_
	);
	LUT2 #(
		.INIT('h2)
	) name5260 (
		\g160_reg/NET0131 ,
		_w5027_,
		_w6440_
	);
	LUT2 #(
		.INIT('h8)
	) name5261 (
		_w2047_,
		_w5027_,
		_w6441_
	);
	LUT2 #(
		.INIT('h1)
	) name5262 (
		_w6440_,
		_w6441_,
		_w6442_
	);
	LUT2 #(
		.INIT('h2)
	) name5263 (
		\g161_reg/NET0131 ,
		_w5029_,
		_w6443_
	);
	LUT2 #(
		.INIT('h8)
	) name5264 (
		_w2047_,
		_w5029_,
		_w6444_
	);
	LUT2 #(
		.INIT('h1)
	) name5265 (
		_w6443_,
		_w6444_,
		_w6445_
	);
	LUT2 #(
		.INIT('h2)
	) name5266 (
		\g162_reg/NET0131 ,
		_w5023_,
		_w6446_
	);
	LUT2 #(
		.INIT('h8)
	) name5267 (
		_w2034_,
		_w5023_,
		_w6447_
	);
	LUT2 #(
		.INIT('h1)
	) name5268 (
		_w6446_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h2)
	) name5269 (
		\g163_reg/NET0131 ,
		_w5027_,
		_w6449_
	);
	LUT2 #(
		.INIT('h8)
	) name5270 (
		_w2034_,
		_w5027_,
		_w6450_
	);
	LUT2 #(
		.INIT('h1)
	) name5271 (
		_w6449_,
		_w6450_,
		_w6451_
	);
	LUT2 #(
		.INIT('h2)
	) name5272 (
		\g164_reg/NET0131 ,
		_w5029_,
		_w6452_
	);
	LUT2 #(
		.INIT('h8)
	) name5273 (
		_w2034_,
		_w5029_,
		_w6453_
	);
	LUT2 #(
		.INIT('h1)
	) name5274 (
		_w6452_,
		_w6453_,
		_w6454_
	);
	LUT2 #(
		.INIT('h2)
	) name5275 (
		\g838_reg/NET0131 ,
		_w5023_,
		_w6455_
	);
	LUT2 #(
		.INIT('h4)
	) name5276 (
		\g805_reg/NET0131 ,
		_w5023_,
		_w6456_
	);
	LUT2 #(
		.INIT('h1)
	) name5277 (
		_w6455_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h2)
	) name5278 (
		\g150_reg/NET0131 ,
		_w5023_,
		_w6458_
	);
	LUT2 #(
		.INIT('h4)
	) name5279 (
		\g117_reg/NET0131 ,
		_w5023_,
		_w6459_
	);
	LUT2 #(
		.INIT('h1)
	) name5280 (
		_w6458_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h2)
	) name5281 (
		\g151_reg/NET0131 ,
		_w5027_,
		_w6461_
	);
	LUT2 #(
		.INIT('h4)
	) name5282 (
		\g117_reg/NET0131 ,
		_w5027_,
		_w6462_
	);
	LUT2 #(
		.INIT('h1)
	) name5283 (
		_w6461_,
		_w6462_,
		_w6463_
	);
	LUT2 #(
		.INIT('h2)
	) name5284 (
		\g152_reg/NET0131 ,
		_w5029_,
		_w6464_
	);
	LUT2 #(
		.INIT('h4)
	) name5285 (
		\g117_reg/NET0131 ,
		_w5029_,
		_w6465_
	);
	LUT2 #(
		.INIT('h1)
	) name5286 (
		_w6464_,
		_w6465_,
		_w6466_
	);
	LUT2 #(
		.INIT('h2)
	) name5287 (
		\g839_reg/NET0131 ,
		_w5027_,
		_w6467_
	);
	LUT2 #(
		.INIT('h4)
	) name5288 (
		\g805_reg/NET0131 ,
		_w5027_,
		_w6468_
	);
	LUT2 #(
		.INIT('h1)
	) name5289 (
		_w6467_,
		_w6468_,
		_w6469_
	);
	LUT2 #(
		.INIT('h2)
	) name5290 (
		\g840_reg/NET0131 ,
		_w5029_,
		_w6470_
	);
	LUT2 #(
		.INIT('h4)
	) name5291 (
		\g805_reg/NET0131 ,
		_w5029_,
		_w6471_
	);
	LUT2 #(
		.INIT('h1)
	) name5292 (
		_w6470_,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h2)
	) name5293 (
		\g844_reg/NET0131 ,
		_w5023_,
		_w6473_
	);
	LUT2 #(
		.INIT('h4)
	) name5294 (
		\g813_reg/NET0131 ,
		_w5023_,
		_w6474_
	);
	LUT2 #(
		.INIT('h1)
	) name5295 (
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h2)
	) name5296 (
		\g845_reg/NET0131 ,
		_w5027_,
		_w6476_
	);
	LUT2 #(
		.INIT('h4)
	) name5297 (
		\g813_reg/NET0131 ,
		_w5027_,
		_w6477_
	);
	LUT2 #(
		.INIT('h1)
	) name5298 (
		_w6476_,
		_w6477_,
		_w6478_
	);
	LUT2 #(
		.INIT('h2)
	) name5299 (
		\g846_reg/NET0131 ,
		_w5029_,
		_w6479_
	);
	LUT2 #(
		.INIT('h4)
	) name5300 (
		\g813_reg/NET0131 ,
		_w5029_,
		_w6480_
	);
	LUT2 #(
		.INIT('h1)
	) name5301 (
		_w6479_,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h2)
	) name5302 (
		\g156_reg/NET0131 ,
		_w5023_,
		_w6482_
	);
	LUT2 #(
		.INIT('h4)
	) name5303 (
		\g125_reg/NET0131 ,
		_w5023_,
		_w6483_
	);
	LUT2 #(
		.INIT('h1)
	) name5304 (
		_w6482_,
		_w6483_,
		_w6484_
	);
	LUT2 #(
		.INIT('h2)
	) name5305 (
		\g157_reg/NET0131 ,
		_w5027_,
		_w6485_
	);
	LUT2 #(
		.INIT('h4)
	) name5306 (
		\g125_reg/NET0131 ,
		_w5027_,
		_w6486_
	);
	LUT2 #(
		.INIT('h1)
	) name5307 (
		_w6485_,
		_w6486_,
		_w6487_
	);
	LUT2 #(
		.INIT('h2)
	) name5308 (
		\g158_reg/NET0131 ,
		_w5029_,
		_w6488_
	);
	LUT2 #(
		.INIT('h4)
	) name5309 (
		\g125_reg/NET0131 ,
		_w5029_,
		_w6489_
	);
	LUT2 #(
		.INIT('h1)
	) name5310 (
		_w6488_,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h8)
	) name5311 (
		\g1196_reg/NET0131 ,
		_w1745_,
		_w6491_
	);
	LUT2 #(
		.INIT('h8)
	) name5312 (
		_w5643_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h8)
	) name5313 (
		\g1196_reg/NET0131 ,
		_w3754_,
		_w6493_
	);
	LUT2 #(
		.INIT('h8)
	) name5314 (
		_w5734_,
		_w6493_,
		_w6494_
	);
	LUT2 #(
		.INIT('h8)
	) name5315 (
		\g1196_reg/NET0131 ,
		_w2929_,
		_w6495_
	);
	LUT2 #(
		.INIT('h8)
	) name5316 (
		_w5766_,
		_w6495_,
		_w6496_
	);
	LUT2 #(
		.INIT('h8)
	) name5317 (
		\g1196_reg/NET0131 ,
		_w1633_,
		_w6497_
	);
	LUT2 #(
		.INIT('h8)
	) name5318 (
		_w5882_,
		_w6497_,
		_w6498_
	);
	LUT2 #(
		.INIT('h1)
	) name5319 (
		\g1332_reg/NET0131 ,
		_w5049_,
		_w6499_
	);
	LUT2 #(
		.INIT('h1)
	) name5320 (
		_w5045_,
		_w5050_,
		_w6500_
	);
	LUT2 #(
		.INIT('h4)
	) name5321 (
		_w6499_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h1)
	) name5322 (
		\g3010_reg/NET0131 ,
		_w6046_,
		_w6502_
	);
	LUT2 #(
		.INIT('h2)
	) name5323 (
		_w6041_,
		_w6047_,
		_w6503_
	);
	LUT2 #(
		.INIT('h4)
	) name5324 (
		_w6502_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h1)
	) name5325 (
		_w5696_,
		_w5716_,
		_w6505_
	);
	LUT2 #(
		.INIT('h1)
	) name5326 (
		_w5697_,
		_w6505_,
		_w6506_
	);
	LUT2 #(
		.INIT('h4)
	) name5327 (
		\g3229_pad ,
		_w4750_,
		_w6507_
	);
	LUT2 #(
		.INIT('h8)
	) name5328 (
		\g3229_pad ,
		_w4776_,
		_w6508_
	);
	LUT2 #(
		.INIT('h1)
	) name5329 (
		_w4752_,
		_w6507_,
		_w6509_
	);
	LUT2 #(
		.INIT('h4)
	) name5330 (
		_w6508_,
		_w6509_,
		_w6510_
	);
	LUT2 #(
		.INIT('h4)
	) name5331 (
		\g3229_pad ,
		_w4232_,
		_w6511_
	);
	LUT2 #(
		.INIT('h8)
	) name5332 (
		\g3229_pad ,
		_w4204_,
		_w6512_
	);
	LUT2 #(
		.INIT('h1)
	) name5333 (
		_w4186_,
		_w6511_,
		_w6513_
	);
	LUT2 #(
		.INIT('h4)
	) name5334 (
		_w6512_,
		_w6513_,
		_w6514_
	);
	LUT2 #(
		.INIT('h1)
	) name5335 (
		_w5822_,
		_w5848_,
		_w6515_
	);
	LUT2 #(
		.INIT('h1)
	) name5336 (
		_w5823_,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h4)
	) name5337 (
		\g3229_pad ,
		_w4922_,
		_w6517_
	);
	LUT2 #(
		.INIT('h8)
	) name5338 (
		\g3229_pad ,
		_w4919_,
		_w6518_
	);
	LUT2 #(
		.INIT('h1)
	) name5339 (
		_w4953_,
		_w6517_,
		_w6519_
	);
	LUT2 #(
		.INIT('h4)
	) name5340 (
		_w6518_,
		_w6519_,
		_w6520_
	);
	LUT2 #(
		.INIT('h1)
	) name5341 (
		_w5921_,
		_w5963_,
		_w6521_
	);
	LUT2 #(
		.INIT('h1)
	) name5342 (
		_w5922_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h1)
	) name5343 (
		\g1339_reg/NET0131 ,
		_w5048_,
		_w6523_
	);
	LUT2 #(
		.INIT('h1)
	) name5344 (
		_w5045_,
		_w5049_,
		_w6524_
	);
	LUT2 #(
		.INIT('h4)
	) name5345 (
		_w6523_,
		_w6524_,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name5346 (
		_w5624_,
		_w5867_,
		_w6526_
	);
	LUT2 #(
		.INIT('h1)
	) name5347 (
		_w5868_,
		_w6526_,
		_w6527_
	);
	LUT2 #(
		.INIT('h1)
	) name5348 (
		\g2814_reg/NET0131 ,
		_w6085_,
		_w6528_
	);
	LUT2 #(
		.INIT('h8)
	) name5349 (
		\g2883_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w6529_
	);
	LUT2 #(
		.INIT('h8)
	) name5350 (
		\g2888_reg/NET0131 ,
		_w6529_,
		_w6530_
	);
	LUT2 #(
		.INIT('h8)
	) name5351 (
		\g2896_reg/NET0131 ,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h8)
	) name5352 (
		\g2892_reg/NET0131 ,
		_w6531_,
		_w6532_
	);
	LUT2 #(
		.INIT('h8)
	) name5353 (
		\g2903_reg/NET0131 ,
		_w6532_,
		_w6533_
	);
	LUT2 #(
		.INIT('h8)
	) name5354 (
		\g2900_reg/NET0131 ,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h1)
	) name5355 (
		\g2908_reg/NET0131 ,
		_w6534_,
		_w6535_
	);
	LUT2 #(
		.INIT('h8)
	) name5356 (
		\g2908_reg/NET0131 ,
		_w6534_,
		_w6536_
	);
	LUT2 #(
		.INIT('h2)
	) name5357 (
		_w6528_,
		_w6535_,
		_w6537_
	);
	LUT2 #(
		.INIT('h4)
	) name5358 (
		_w6536_,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h2)
	) name5359 (
		\g2080_reg/NET0131 ,
		_w4704_,
		_w6539_
	);
	LUT2 #(
		.INIT('h4)
	) name5360 (
		\g1326_reg/NET0131 ,
		_w4704_,
		_w6540_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w6539_,
		_w6540_,
		_w6541_
	);
	LUT2 #(
		.INIT('h2)
	) name5362 (
		\g2103_reg/NET0131 ,
		_w4708_,
		_w6542_
	);
	LUT2 #(
		.INIT('h4)
	) name5363 (
		\g1372_reg/NET0131 ,
		_w4708_,
		_w6543_
	);
	LUT2 #(
		.INIT('h1)
	) name5364 (
		_w6542_,
		_w6543_,
		_w6544_
	);
	LUT2 #(
		.INIT('h2)
	) name5365 (
		\g2092_reg/NET0131 ,
		_w4704_,
		_w6545_
	);
	LUT2 #(
		.INIT('h4)
	) name5366 (
		\g1346_reg/NET0131 ,
		_w4704_,
		_w6546_
	);
	LUT2 #(
		.INIT('h1)
	) name5367 (
		_w6545_,
		_w6546_,
		_w6547_
	);
	LUT2 #(
		.INIT('h2)
	) name5368 (
		\g2078_reg/NET0131 ,
		_w4594_,
		_w6548_
	);
	LUT2 #(
		.INIT('h4)
	) name5369 (
		\g1326_reg/NET0131 ,
		_w4594_,
		_w6549_
	);
	LUT2 #(
		.INIT('h1)
	) name5370 (
		_w6548_,
		_w6549_,
		_w6550_
	);
	LUT2 #(
		.INIT('h2)
	) name5371 (
		\g2079_reg/NET0131 ,
		_w4708_,
		_w6551_
	);
	LUT2 #(
		.INIT('h4)
	) name5372 (
		\g1326_reg/NET0131 ,
		_w4708_,
		_w6552_
	);
	LUT2 #(
		.INIT('h1)
	) name5373 (
		_w6551_,
		_w6552_,
		_w6553_
	);
	LUT2 #(
		.INIT('h2)
	) name5374 (
		\g2081_reg/NET0131 ,
		_w4594_,
		_w6554_
	);
	LUT2 #(
		.INIT('h4)
	) name5375 (
		\g1319_reg/NET0131 ,
		_w4594_,
		_w6555_
	);
	LUT2 #(
		.INIT('h1)
	) name5376 (
		_w6554_,
		_w6555_,
		_w6556_
	);
	LUT2 #(
		.INIT('h2)
	) name5377 (
		\g2082_reg/NET0131 ,
		_w4708_,
		_w6557_
	);
	LUT2 #(
		.INIT('h4)
	) name5378 (
		\g1319_reg/NET0131 ,
		_w4708_,
		_w6558_
	);
	LUT2 #(
		.INIT('h1)
	) name5379 (
		_w6557_,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h2)
	) name5380 (
		\g2083_reg/NET0131 ,
		_w4704_,
		_w6560_
	);
	LUT2 #(
		.INIT('h4)
	) name5381 (
		\g1319_reg/NET0131 ,
		_w4704_,
		_w6561_
	);
	LUT2 #(
		.INIT('h1)
	) name5382 (
		_w6560_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h2)
	) name5383 (
		\g2084_reg/NET0131 ,
		_w4594_,
		_w6563_
	);
	LUT2 #(
		.INIT('h4)
	) name5384 (
		\g1339_reg/NET0131 ,
		_w4594_,
		_w6564_
	);
	LUT2 #(
		.INIT('h1)
	) name5385 (
		_w6563_,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h2)
	) name5386 (
		\g2085_reg/NET0131 ,
		_w4708_,
		_w6566_
	);
	LUT2 #(
		.INIT('h4)
	) name5387 (
		\g1339_reg/NET0131 ,
		_w4708_,
		_w6567_
	);
	LUT2 #(
		.INIT('h1)
	) name5388 (
		_w6566_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h2)
	) name5389 (
		\g2087_reg/NET0131 ,
		_w4594_,
		_w6569_
	);
	LUT2 #(
		.INIT('h4)
	) name5390 (
		\g1332_reg/NET0131 ,
		_w4594_,
		_w6570_
	);
	LUT2 #(
		.INIT('h1)
	) name5391 (
		_w6569_,
		_w6570_,
		_w6571_
	);
	LUT2 #(
		.INIT('h2)
	) name5392 (
		\g2089_reg/NET0131 ,
		_w4704_,
		_w6572_
	);
	LUT2 #(
		.INIT('h4)
	) name5393 (
		\g1332_reg/NET0131 ,
		_w4704_,
		_w6573_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		_w6572_,
		_w6573_,
		_w6574_
	);
	LUT2 #(
		.INIT('h2)
	) name5395 (
		\g2093_reg/NET0131 ,
		_w4594_,
		_w6575_
	);
	LUT2 #(
		.INIT('h4)
	) name5396 (
		\g1358_reg/NET0131 ,
		_w4594_,
		_w6576_
	);
	LUT2 #(
		.INIT('h1)
	) name5397 (
		_w6575_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h2)
	) name5398 (
		\g2095_reg/NET0131 ,
		_w4704_,
		_w6578_
	);
	LUT2 #(
		.INIT('h4)
	) name5399 (
		\g1358_reg/NET0131 ,
		_w4704_,
		_w6579_
	);
	LUT2 #(
		.INIT('h1)
	) name5400 (
		_w6578_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h2)
	) name5401 (
		\g2097_reg/NET0131 ,
		_w4708_,
		_w6581_
	);
	LUT2 #(
		.INIT('h4)
	) name5402 (
		\g1352_reg/NET0131 ,
		_w4708_,
		_w6582_
	);
	LUT2 #(
		.INIT('h1)
	) name5403 (
		_w6581_,
		_w6582_,
		_w6583_
	);
	LUT2 #(
		.INIT('h2)
	) name5404 (
		\g2099_reg/NET0131 ,
		_w4594_,
		_w6584_
	);
	LUT2 #(
		.INIT('h4)
	) name5405 (
		\g1365_reg/NET0131 ,
		_w4594_,
		_w6585_
	);
	LUT2 #(
		.INIT('h1)
	) name5406 (
		_w6584_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h2)
	) name5407 (
		\g2100_reg/NET0131 ,
		_w4708_,
		_w6587_
	);
	LUT2 #(
		.INIT('h4)
	) name5408 (
		\g1365_reg/NET0131 ,
		_w4708_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name5409 (
		_w6587_,
		_w6588_,
		_w6589_
	);
	LUT2 #(
		.INIT('h2)
	) name5410 (
		\g2101_reg/NET0131 ,
		_w4704_,
		_w6590_
	);
	LUT2 #(
		.INIT('h4)
	) name5411 (
		\g1365_reg/NET0131 ,
		_w4704_,
		_w6591_
	);
	LUT2 #(
		.INIT('h1)
	) name5412 (
		_w6590_,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h2)
	) name5413 (
		\g2102_reg/NET0131 ,
		_w4594_,
		_w6593_
	);
	LUT2 #(
		.INIT('h4)
	) name5414 (
		\g1372_reg/NET0131 ,
		_w4594_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name5415 (
		_w6593_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h2)
	) name5416 (
		\g2104_reg/NET0131 ,
		_w4704_,
		_w6596_
	);
	LUT2 #(
		.INIT('h4)
	) name5417 (
		\g1372_reg/NET0131 ,
		_w4704_,
		_w6597_
	);
	LUT2 #(
		.INIT('h1)
	) name5418 (
		_w6596_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h2)
	) name5419 (
		\g2106_reg/NET0131 ,
		_w4708_,
		_w6599_
	);
	LUT2 #(
		.INIT('h4)
	) name5420 (
		\g1378_reg/NET0131 ,
		_w4708_,
		_w6600_
	);
	LUT2 #(
		.INIT('h1)
	) name5421 (
		_w6599_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h2)
	) name5422 (
		\g2107_reg/NET0131 ,
		_w4704_,
		_w6602_
	);
	LUT2 #(
		.INIT('h4)
	) name5423 (
		\g1378_reg/NET0131 ,
		_w4704_,
		_w6603_
	);
	LUT2 #(
		.INIT('h1)
	) name5424 (
		_w6602_,
		_w6603_,
		_w6604_
	);
	LUT2 #(
		.INIT('h2)
	) name5425 (
		\g2091_reg/NET0131 ,
		_w4708_,
		_w6605_
	);
	LUT2 #(
		.INIT('h4)
	) name5426 (
		\g1346_reg/NET0131 ,
		_w4708_,
		_w6606_
	);
	LUT2 #(
		.INIT('h1)
	) name5427 (
		_w6605_,
		_w6606_,
		_w6607_
	);
	LUT2 #(
		.INIT('h2)
	) name5428 (
		\g2090_reg/NET0131 ,
		_w4594_,
		_w6608_
	);
	LUT2 #(
		.INIT('h4)
	) name5429 (
		\g1346_reg/NET0131 ,
		_w4594_,
		_w6609_
	);
	LUT2 #(
		.INIT('h1)
	) name5430 (
		_w6608_,
		_w6609_,
		_w6610_
	);
	LUT2 #(
		.INIT('h2)
	) name5431 (
		\g2086_reg/NET0131 ,
		_w4704_,
		_w6611_
	);
	LUT2 #(
		.INIT('h4)
	) name5432 (
		\g1339_reg/NET0131 ,
		_w4704_,
		_w6612_
	);
	LUT2 #(
		.INIT('h1)
	) name5433 (
		_w6611_,
		_w6612_,
		_w6613_
	);
	LUT2 #(
		.INIT('h2)
	) name5434 (
		\g2788_reg/NET0131 ,
		_w4478_,
		_w6614_
	);
	LUT2 #(
		.INIT('h4)
	) name5435 (
		\g1358_reg/NET0131 ,
		_w4478_,
		_w6615_
	);
	LUT2 #(
		.INIT('h1)
	) name5436 (
		_w6614_,
		_w6615_,
		_w6616_
	);
	LUT2 #(
		.INIT('h2)
	) name5437 (
		\g2105_reg/NET0131 ,
		_w4594_,
		_w6617_
	);
	LUT2 #(
		.INIT('h4)
	) name5438 (
		\g1378_reg/NET0131 ,
		_w4594_,
		_w6618_
	);
	LUT2 #(
		.INIT('h1)
	) name5439 (
		_w6617_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('h2)
	) name5440 (
		\g2088_reg/NET0131 ,
		_w4708_,
		_w6620_
	);
	LUT2 #(
		.INIT('h4)
	) name5441 (
		\g1332_reg/NET0131 ,
		_w4708_,
		_w6621_
	);
	LUT2 #(
		.INIT('h1)
	) name5442 (
		_w6620_,
		_w6621_,
		_w6622_
	);
	LUT2 #(
		.INIT('h2)
	) name5443 (
		\g2098_reg/NET0131 ,
		_w4704_,
		_w6623_
	);
	LUT2 #(
		.INIT('h4)
	) name5444 (
		\g1352_reg/NET0131 ,
		_w4704_,
		_w6624_
	);
	LUT2 #(
		.INIT('h1)
	) name5445 (
		_w6623_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h2)
	) name5446 (
		\g2094_reg/NET0131 ,
		_w4708_,
		_w6626_
	);
	LUT2 #(
		.INIT('h4)
	) name5447 (
		\g1358_reg/NET0131 ,
		_w4708_,
		_w6627_
	);
	LUT2 #(
		.INIT('h1)
	) name5448 (
		_w6626_,
		_w6627_,
		_w6628_
	);
	LUT2 #(
		.INIT('h2)
	) name5449 (
		\g2772_reg/NET0131 ,
		_w4712_,
		_w6629_
	);
	LUT2 #(
		.INIT('h4)
	) name5450 (
		\g1326_reg/NET0131 ,
		_w4712_,
		_w6630_
	);
	LUT2 #(
		.INIT('h1)
	) name5451 (
		_w6629_,
		_w6630_,
		_w6631_
	);
	LUT2 #(
		.INIT('h2)
	) name5452 (
		\g2773_reg/NET0131 ,
		_w4478_,
		_w6632_
	);
	LUT2 #(
		.INIT('h4)
	) name5453 (
		\g1326_reg/NET0131 ,
		_w4478_,
		_w6633_
	);
	LUT2 #(
		.INIT('h1)
	) name5454 (
		_w6632_,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h2)
	) name5455 (
		\g2774_reg/NET0131 ,
		_w4528_,
		_w6635_
	);
	LUT2 #(
		.INIT('h4)
	) name5456 (
		\g1326_reg/NET0131 ,
		_w4528_,
		_w6636_
	);
	LUT2 #(
		.INIT('h1)
	) name5457 (
		_w6635_,
		_w6636_,
		_w6637_
	);
	LUT2 #(
		.INIT('h2)
	) name5458 (
		\g2775_reg/NET0131 ,
		_w4712_,
		_w6638_
	);
	LUT2 #(
		.INIT('h4)
	) name5459 (
		\g1319_reg/NET0131 ,
		_w4712_,
		_w6639_
	);
	LUT2 #(
		.INIT('h1)
	) name5460 (
		_w6638_,
		_w6639_,
		_w6640_
	);
	LUT2 #(
		.INIT('h2)
	) name5461 (
		\g2776_reg/NET0131 ,
		_w4478_,
		_w6641_
	);
	LUT2 #(
		.INIT('h4)
	) name5462 (
		\g1319_reg/NET0131 ,
		_w4478_,
		_w6642_
	);
	LUT2 #(
		.INIT('h1)
	) name5463 (
		_w6641_,
		_w6642_,
		_w6643_
	);
	LUT2 #(
		.INIT('h2)
	) name5464 (
		\g2777_reg/NET0131 ,
		_w4528_,
		_w6644_
	);
	LUT2 #(
		.INIT('h4)
	) name5465 (
		\g1319_reg/NET0131 ,
		_w4528_,
		_w6645_
	);
	LUT2 #(
		.INIT('h1)
	) name5466 (
		_w6644_,
		_w6645_,
		_w6646_
	);
	LUT2 #(
		.INIT('h2)
	) name5467 (
		\g2778_reg/NET0131 ,
		_w4712_,
		_w6647_
	);
	LUT2 #(
		.INIT('h4)
	) name5468 (
		\g1339_reg/NET0131 ,
		_w4712_,
		_w6648_
	);
	LUT2 #(
		.INIT('h1)
	) name5469 (
		_w6647_,
		_w6648_,
		_w6649_
	);
	LUT2 #(
		.INIT('h2)
	) name5470 (
		\g2779_reg/NET0131 ,
		_w4478_,
		_w6650_
	);
	LUT2 #(
		.INIT('h4)
	) name5471 (
		\g1339_reg/NET0131 ,
		_w4478_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name5472 (
		_w6650_,
		_w6651_,
		_w6652_
	);
	LUT2 #(
		.INIT('h2)
	) name5473 (
		\g2780_reg/NET0131 ,
		_w4528_,
		_w6653_
	);
	LUT2 #(
		.INIT('h4)
	) name5474 (
		\g1339_reg/NET0131 ,
		_w4528_,
		_w6654_
	);
	LUT2 #(
		.INIT('h1)
	) name5475 (
		_w6653_,
		_w6654_,
		_w6655_
	);
	LUT2 #(
		.INIT('h2)
	) name5476 (
		\g2781_reg/NET0131 ,
		_w4712_,
		_w6656_
	);
	LUT2 #(
		.INIT('h4)
	) name5477 (
		\g1332_reg/NET0131 ,
		_w4712_,
		_w6657_
	);
	LUT2 #(
		.INIT('h1)
	) name5478 (
		_w6656_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h2)
	) name5479 (
		\g2782_reg/NET0131 ,
		_w4478_,
		_w6659_
	);
	LUT2 #(
		.INIT('h4)
	) name5480 (
		\g1332_reg/NET0131 ,
		_w4478_,
		_w6660_
	);
	LUT2 #(
		.INIT('h1)
	) name5481 (
		_w6659_,
		_w6660_,
		_w6661_
	);
	LUT2 #(
		.INIT('h2)
	) name5482 (
		\g2783_reg/NET0131 ,
		_w4528_,
		_w6662_
	);
	LUT2 #(
		.INIT('h4)
	) name5483 (
		\g1332_reg/NET0131 ,
		_w4528_,
		_w6663_
	);
	LUT2 #(
		.INIT('h1)
	) name5484 (
		_w6662_,
		_w6663_,
		_w6664_
	);
	LUT2 #(
		.INIT('h2)
	) name5485 (
		\g2784_reg/NET0131 ,
		_w4712_,
		_w6665_
	);
	LUT2 #(
		.INIT('h4)
	) name5486 (
		\g1346_reg/NET0131 ,
		_w4712_,
		_w6666_
	);
	LUT2 #(
		.INIT('h1)
	) name5487 (
		_w6665_,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h2)
	) name5488 (
		\g2785_reg/NET0131 ,
		_w4478_,
		_w6668_
	);
	LUT2 #(
		.INIT('h4)
	) name5489 (
		\g1346_reg/NET0131 ,
		_w4478_,
		_w6669_
	);
	LUT2 #(
		.INIT('h1)
	) name5490 (
		_w6668_,
		_w6669_,
		_w6670_
	);
	LUT2 #(
		.INIT('h2)
	) name5491 (
		\g2786_reg/NET0131 ,
		_w4528_,
		_w6671_
	);
	LUT2 #(
		.INIT('h4)
	) name5492 (
		\g1346_reg/NET0131 ,
		_w4528_,
		_w6672_
	);
	LUT2 #(
		.INIT('h1)
	) name5493 (
		_w6671_,
		_w6672_,
		_w6673_
	);
	LUT2 #(
		.INIT('h2)
	) name5494 (
		\g2787_reg/NET0131 ,
		_w4712_,
		_w6674_
	);
	LUT2 #(
		.INIT('h4)
	) name5495 (
		\g1358_reg/NET0131 ,
		_w4712_,
		_w6675_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		_w6674_,
		_w6675_,
		_w6676_
	);
	LUT2 #(
		.INIT('h2)
	) name5497 (
		\g2789_reg/NET0131 ,
		_w4528_,
		_w6677_
	);
	LUT2 #(
		.INIT('h4)
	) name5498 (
		\g1358_reg/NET0131 ,
		_w4528_,
		_w6678_
	);
	LUT2 #(
		.INIT('h1)
	) name5499 (
		_w6677_,
		_w6678_,
		_w6679_
	);
	LUT2 #(
		.INIT('h2)
	) name5500 (
		\g2790_reg/NET0131 ,
		_w4712_,
		_w6680_
	);
	LUT2 #(
		.INIT('h4)
	) name5501 (
		\g1352_reg/NET0131 ,
		_w4712_,
		_w6681_
	);
	LUT2 #(
		.INIT('h1)
	) name5502 (
		_w6680_,
		_w6681_,
		_w6682_
	);
	LUT2 #(
		.INIT('h2)
	) name5503 (
		\g2791_reg/NET0131 ,
		_w4478_,
		_w6683_
	);
	LUT2 #(
		.INIT('h4)
	) name5504 (
		\g1352_reg/NET0131 ,
		_w4478_,
		_w6684_
	);
	LUT2 #(
		.INIT('h1)
	) name5505 (
		_w6683_,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('h2)
	) name5506 (
		\g2792_reg/NET0131 ,
		_w4528_,
		_w6686_
	);
	LUT2 #(
		.INIT('h4)
	) name5507 (
		\g1352_reg/NET0131 ,
		_w4528_,
		_w6687_
	);
	LUT2 #(
		.INIT('h1)
	) name5508 (
		_w6686_,
		_w6687_,
		_w6688_
	);
	LUT2 #(
		.INIT('h2)
	) name5509 (
		\g2793_reg/NET0131 ,
		_w4712_,
		_w6689_
	);
	LUT2 #(
		.INIT('h4)
	) name5510 (
		\g1365_reg/NET0131 ,
		_w4712_,
		_w6690_
	);
	LUT2 #(
		.INIT('h1)
	) name5511 (
		_w6689_,
		_w6690_,
		_w6691_
	);
	LUT2 #(
		.INIT('h2)
	) name5512 (
		\g2096_reg/NET0131 ,
		_w4594_,
		_w6692_
	);
	LUT2 #(
		.INIT('h4)
	) name5513 (
		\g1352_reg/NET0131 ,
		_w4594_,
		_w6693_
	);
	LUT2 #(
		.INIT('h1)
	) name5514 (
		_w6692_,
		_w6693_,
		_w6694_
	);
	LUT2 #(
		.INIT('h2)
	) name5515 (
		\g2794_reg/NET0131 ,
		_w4478_,
		_w6695_
	);
	LUT2 #(
		.INIT('h4)
	) name5516 (
		\g1365_reg/NET0131 ,
		_w4478_,
		_w6696_
	);
	LUT2 #(
		.INIT('h1)
	) name5517 (
		_w6695_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h2)
	) name5518 (
		\g2795_reg/NET0131 ,
		_w4528_,
		_w6698_
	);
	LUT2 #(
		.INIT('h4)
	) name5519 (
		\g1365_reg/NET0131 ,
		_w4528_,
		_w6699_
	);
	LUT2 #(
		.INIT('h1)
	) name5520 (
		_w6698_,
		_w6699_,
		_w6700_
	);
	LUT2 #(
		.INIT('h2)
	) name5521 (
		\g2796_reg/NET0131 ,
		_w4712_,
		_w6701_
	);
	LUT2 #(
		.INIT('h4)
	) name5522 (
		\g1372_reg/NET0131 ,
		_w4712_,
		_w6702_
	);
	LUT2 #(
		.INIT('h1)
	) name5523 (
		_w6701_,
		_w6702_,
		_w6703_
	);
	LUT2 #(
		.INIT('h2)
	) name5524 (
		\g2797_reg/NET0131 ,
		_w4478_,
		_w6704_
	);
	LUT2 #(
		.INIT('h4)
	) name5525 (
		\g1372_reg/NET0131 ,
		_w4478_,
		_w6705_
	);
	LUT2 #(
		.INIT('h1)
	) name5526 (
		_w6704_,
		_w6705_,
		_w6706_
	);
	LUT2 #(
		.INIT('h2)
	) name5527 (
		\g2798_reg/NET0131 ,
		_w4528_,
		_w6707_
	);
	LUT2 #(
		.INIT('h4)
	) name5528 (
		\g1372_reg/NET0131 ,
		_w4528_,
		_w6708_
	);
	LUT2 #(
		.INIT('h1)
	) name5529 (
		_w6707_,
		_w6708_,
		_w6709_
	);
	LUT2 #(
		.INIT('h2)
	) name5530 (
		\g2799_reg/NET0131 ,
		_w4712_,
		_w6710_
	);
	LUT2 #(
		.INIT('h4)
	) name5531 (
		\g1378_reg/NET0131 ,
		_w4712_,
		_w6711_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		_w6710_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h2)
	) name5533 (
		\g2800_reg/NET0131 ,
		_w4478_,
		_w6713_
	);
	LUT2 #(
		.INIT('h4)
	) name5534 (
		\g1378_reg/NET0131 ,
		_w4478_,
		_w6714_
	);
	LUT2 #(
		.INIT('h1)
	) name5535 (
		_w6713_,
		_w6714_,
		_w6715_
	);
	LUT2 #(
		.INIT('h2)
	) name5536 (
		\g2801_reg/NET0131 ,
		_w4528_,
		_w6716_
	);
	LUT2 #(
		.INIT('h4)
	) name5537 (
		\g1378_reg/NET0131 ,
		_w4528_,
		_w6717_
	);
	LUT2 #(
		.INIT('h1)
	) name5538 (
		_w6716_,
		_w6717_,
		_w6718_
	);
	LUT2 #(
		.INIT('h2)
	) name5539 (
		\g7961_pad ,
		_w5036_,
		_w6719_
	);
	LUT2 #(
		.INIT('h1)
	) name5540 (
		\g1164_reg/NET0131 ,
		\g7961_pad ,
		_w6720_
	);
	LUT2 #(
		.INIT('h1)
	) name5541 (
		_w6719_,
		_w6720_,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name5542 (
		\g2900_reg/NET0131 ,
		_w6533_,
		_w6722_
	);
	LUT2 #(
		.INIT('h2)
	) name5543 (
		_w6528_,
		_w6534_,
		_w6723_
	);
	LUT2 #(
		.INIT('h4)
	) name5544 (
		_w6722_,
		_w6723_,
		_w6724_
	);
	LUT2 #(
		.INIT('h1)
	) name5545 (
		\g2924_reg/NET0131 ,
		_w6091_,
		_w6725_
	);
	LUT2 #(
		.INIT('h2)
	) name5546 (
		_w6090_,
		_w6092_,
		_w6726_
	);
	LUT2 #(
		.INIT('h4)
	) name5547 (
		_w6725_,
		_w6726_,
		_w6727_
	);
	LUT2 #(
		.INIT('h1)
	) name5548 (
		\g1319_reg/NET0131 ,
		_w5047_,
		_w6728_
	);
	LUT2 #(
		.INIT('h1)
	) name5549 (
		_w5045_,
		_w5048_,
		_w6729_
	);
	LUT2 #(
		.INIT('h4)
	) name5550 (
		_w6728_,
		_w6729_,
		_w6730_
	);
	LUT2 #(
		.INIT('h1)
	) name5551 (
		\g2917_reg/NET0131 ,
		_w6086_,
		_w6731_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		_w6091_,
		_w6731_,
		_w6732_
	);
	LUT2 #(
		.INIT('h8)
	) name5553 (
		_w6090_,
		_w6732_,
		_w6733_
	);
	LUT2 #(
		.INIT('h2)
	) name5554 (
		\g3139_reg/NET0131 ,
		\g3231_pad ,
		_w6734_
	);
	LUT2 #(
		.INIT('h2)
	) name5555 (
		\g2969_reg/NET0131 ,
		\g2972_reg/NET0131 ,
		_w6735_
	);
	LUT2 #(
		.INIT('h4)
	) name5556 (
		\g2969_reg/NET0131 ,
		\g2972_reg/NET0131 ,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name5557 (
		_w6735_,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('h1)
	) name5558 (
		\g2975_reg/NET0131 ,
		\g2978_reg/NET0131 ,
		_w6738_
	);
	LUT2 #(
		.INIT('h8)
	) name5559 (
		\g2975_reg/NET0131 ,
		\g2978_reg/NET0131 ,
		_w6739_
	);
	LUT2 #(
		.INIT('h1)
	) name5560 (
		_w6738_,
		_w6739_,
		_w6740_
	);
	LUT2 #(
		.INIT('h8)
	) name5561 (
		\g2966_reg/NET0131 ,
		_w6740_,
		_w6741_
	);
	LUT2 #(
		.INIT('h1)
	) name5562 (
		\g2966_reg/NET0131 ,
		_w6740_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name5563 (
		_w6741_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h2)
	) name5564 (
		\g2874_reg/NET0131 ,
		\g2981_reg/NET0131 ,
		_w6744_
	);
	LUT2 #(
		.INIT('h4)
	) name5565 (
		\g2874_reg/NET0131 ,
		\g2981_reg/NET0131 ,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name5566 (
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h8)
	) name5567 (
		\g2963_reg/NET0131 ,
		_w6746_,
		_w6747_
	);
	LUT2 #(
		.INIT('h1)
	) name5568 (
		\g2963_reg/NET0131 ,
		_w6746_,
		_w6748_
	);
	LUT2 #(
		.INIT('h1)
	) name5569 (
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h2)
	) name5570 (
		_w6743_,
		_w6749_,
		_w6750_
	);
	LUT2 #(
		.INIT('h4)
	) name5571 (
		_w6743_,
		_w6749_,
		_w6751_
	);
	LUT2 #(
		.INIT('h1)
	) name5572 (
		_w6750_,
		_w6751_,
		_w6752_
	);
	LUT2 #(
		.INIT('h8)
	) name5573 (
		_w6737_,
		_w6752_,
		_w6753_
	);
	LUT2 #(
		.INIT('h1)
	) name5574 (
		_w6737_,
		_w6752_,
		_w6754_
	);
	LUT2 #(
		.INIT('h1)
	) name5575 (
		_w6753_,
		_w6754_,
		_w6755_
	);
	LUT2 #(
		.INIT('h4)
	) name5576 (
		_w6734_,
		_w6755_,
		_w6756_
	);
	LUT2 #(
		.INIT('h2)
	) name5577 (
		_w6734_,
		_w6755_,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name5578 (
		_w6756_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h2)
	) name5579 (
		\g2947_reg/NET0131 ,
		\g2953_reg/NET0131 ,
		_w6759_
	);
	LUT2 #(
		.INIT('h4)
	) name5580 (
		\g2947_reg/NET0131 ,
		\g2953_reg/NET0131 ,
		_w6760_
	);
	LUT2 #(
		.INIT('h1)
	) name5581 (
		_w6759_,
		_w6760_,
		_w6761_
	);
	LUT2 #(
		.INIT('h1)
	) name5582 (
		\g2935_reg/NET0131 ,
		\g2938_reg/NET0131 ,
		_w6762_
	);
	LUT2 #(
		.INIT('h8)
	) name5583 (
		\g2935_reg/NET0131 ,
		\g2938_reg/NET0131 ,
		_w6763_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		_w6762_,
		_w6763_,
		_w6764_
	);
	LUT2 #(
		.INIT('h8)
	) name5585 (
		\g2959_reg/NET0131 ,
		_w6764_,
		_w6765_
	);
	LUT2 #(
		.INIT('h1)
	) name5586 (
		\g2959_reg/NET0131 ,
		_w6764_,
		_w6766_
	);
	LUT2 #(
		.INIT('h1)
	) name5587 (
		_w6765_,
		_w6766_,
		_w6767_
	);
	LUT2 #(
		.INIT('h2)
	) name5588 (
		\g2941_reg/NET0131 ,
		\g2944_reg/NET0131 ,
		_w6768_
	);
	LUT2 #(
		.INIT('h4)
	) name5589 (
		\g2941_reg/NET0131 ,
		\g2944_reg/NET0131 ,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name5590 (
		_w6768_,
		_w6769_,
		_w6770_
	);
	LUT2 #(
		.INIT('h8)
	) name5591 (
		\g2956_reg/NET0131 ,
		_w6770_,
		_w6771_
	);
	LUT2 #(
		.INIT('h1)
	) name5592 (
		\g2956_reg/NET0131 ,
		_w6770_,
		_w6772_
	);
	LUT2 #(
		.INIT('h1)
	) name5593 (
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT2 #(
		.INIT('h2)
	) name5594 (
		_w6767_,
		_w6773_,
		_w6774_
	);
	LUT2 #(
		.INIT('h4)
	) name5595 (
		_w6767_,
		_w6773_,
		_w6775_
	);
	LUT2 #(
		.INIT('h1)
	) name5596 (
		_w6774_,
		_w6775_,
		_w6776_
	);
	LUT2 #(
		.INIT('h8)
	) name5597 (
		_w6761_,
		_w6776_,
		_w6777_
	);
	LUT2 #(
		.INIT('h1)
	) name5598 (
		_w6761_,
		_w6776_,
		_w6778_
	);
	LUT2 #(
		.INIT('h1)
	) name5599 (
		_w6777_,
		_w6778_,
		_w6779_
	);
	LUT2 #(
		.INIT('h4)
	) name5600 (
		_w6734_,
		_w6779_,
		_w6780_
	);
	LUT2 #(
		.INIT('h2)
	) name5601 (
		_w6734_,
		_w6779_,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name5602 (
		_w6780_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h8)
	) name5603 (
		\g2934_reg/NET0131 ,
		_w6779_,
		_w6783_
	);
	LUT2 #(
		.INIT('h1)
	) name5604 (
		\g2934_reg/NET0131 ,
		_w6779_,
		_w6784_
	);
	LUT2 #(
		.INIT('h1)
	) name5605 (
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT2 #(
		.INIT('h8)
	) name5606 (
		\g2962_reg/NET0131 ,
		_w6755_,
		_w6786_
	);
	LUT2 #(
		.INIT('h1)
	) name5607 (
		\g2962_reg/NET0131 ,
		_w6755_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name5608 (
		_w6786_,
		_w6787_,
		_w6788_
	);
	LUT2 #(
		.INIT('h1)
	) name5609 (
		\g2912_reg/NET0131 ,
		_w6085_,
		_w6789_
	);
	LUT2 #(
		.INIT('h1)
	) name5610 (
		_w6086_,
		_w6789_,
		_w6790_
	);
	LUT2 #(
		.INIT('h2)
	) name5611 (
		_w6090_,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h1)
	) name5612 (
		\g3002_reg/NET0131 ,
		_w6044_,
		_w6792_
	);
	LUT2 #(
		.INIT('h1)
	) name5613 (
		_w6045_,
		_w6792_,
		_w6793_
	);
	LUT2 #(
		.INIT('h8)
	) name5614 (
		_w6041_,
		_w6793_,
		_w6794_
	);
	LUT2 #(
		.INIT('h8)
	) name5615 (
		\g2993_reg/NET0131 ,
		\g3080_reg/NET0131 ,
		_w6795_
	);
	LUT2 #(
		.INIT('h1)
	) name5616 (
		\g2998_reg/NET0131 ,
		_w6795_,
		_w6796_
	);
	LUT2 #(
		.INIT('h1)
	) name5617 (
		_w6043_,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h8)
	) name5618 (
		_w6041_,
		_w6797_,
		_w6798_
	);
	LUT2 #(
		.INIT('h1)
	) name5619 (
		\g3234_pad ,
		_w6798_,
		_w6799_
	);
	LUT2 #(
		.INIT('h2)
	) name5620 (
		\g1018_reg/NET0131 ,
		\g1867_reg/NET0131 ,
		_w6800_
	);
	LUT2 #(
		.INIT('h2)
	) name5621 (
		\g1024_reg/NET0131 ,
		\g1868_reg/NET0131 ,
		_w6801_
	);
	LUT2 #(
		.INIT('h4)
	) name5622 (
		\g1869_reg/NET0131 ,
		\g5657_pad ,
		_w6802_
	);
	LUT2 #(
		.INIT('h1)
	) name5623 (
		_w6800_,
		_w6801_,
		_w6803_
	);
	LUT2 #(
		.INIT('h4)
	) name5624 (
		_w6802_,
		_w6803_,
		_w6804_
	);
	LUT2 #(
		.INIT('h2)
	) name5625 (
		\g1018_reg/NET0131 ,
		\g486_reg/NET0131 ,
		_w6805_
	);
	LUT2 #(
		.INIT('h2)
	) name5626 (
		\g1024_reg/NET0131 ,
		\g487_reg/NET0131 ,
		_w6806_
	);
	LUT2 #(
		.INIT('h4)
	) name5627 (
		\g488_reg/NET0131 ,
		\g5657_pad ,
		_w6807_
	);
	LUT2 #(
		.INIT('h1)
	) name5628 (
		_w6805_,
		_w6806_,
		_w6808_
	);
	LUT2 #(
		.INIT('h4)
	) name5629 (
		_w6807_,
		_w6808_,
		_w6809_
	);
	LUT2 #(
		.INIT('h2)
	) name5630 (
		\g1018_reg/NET0131 ,
		\g1858_reg/NET0131 ,
		_w6810_
	);
	LUT2 #(
		.INIT('h2)
	) name5631 (
		\g1024_reg/NET0131 ,
		\g1859_reg/NET0131 ,
		_w6811_
	);
	LUT2 #(
		.INIT('h4)
	) name5632 (
		\g1860_reg/NET0131 ,
		\g5657_pad ,
		_w6812_
	);
	LUT2 #(
		.INIT('h1)
	) name5633 (
		_w6810_,
		_w6811_,
		_w6813_
	);
	LUT2 #(
		.INIT('h4)
	) name5634 (
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h2)
	) name5635 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		_w6815_
	);
	LUT2 #(
		.INIT('h1)
	) name5636 (
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w6816_
	);
	LUT2 #(
		.INIT('h4)
	) name5637 (
		\g2920_reg/NET0131 ,
		\g2924_reg/NET0131 ,
		_w6817_
	);
	LUT2 #(
		.INIT('h8)
	) name5638 (
		_w6816_,
		_w6817_,
		_w6818_
	);
	LUT2 #(
		.INIT('h8)
	) name5639 (
		_w6815_,
		_w6818_,
		_w6819_
	);
	LUT2 #(
		.INIT('h8)
	) name5640 (
		_w5262_,
		_w6819_,
		_w6820_
	);
	LUT2 #(
		.INIT('h8)
	) name5641 (
		\g1088_reg/NET0131 ,
		_w6820_,
		_w6821_
	);
	LUT2 #(
		.INIT('h2)
	) name5642 (
		\g856_reg/NET0131 ,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('h1)
	) name5643 (
		\g805_reg/NET0131 ,
		\g809_reg/NET0131 ,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name5644 (
		_w5079_,
		_w6823_,
		_w6824_
	);
	LUT2 #(
		.INIT('h8)
	) name5645 (
		_w6821_,
		_w6824_,
		_w6825_
	);
	LUT2 #(
		.INIT('h1)
	) name5646 (
		_w6822_,
		_w6825_,
		_w6826_
	);
	LUT2 #(
		.INIT('h8)
	) name5647 (
		\g7961_pad ,
		_w6820_,
		_w6827_
	);
	LUT2 #(
		.INIT('h2)
	) name5648 (
		\g857_reg/NET0131 ,
		_w6827_,
		_w6828_
	);
	LUT2 #(
		.INIT('h8)
	) name5649 (
		_w6824_,
		_w6827_,
		_w6829_
	);
	LUT2 #(
		.INIT('h1)
	) name5650 (
		_w6828_,
		_w6829_,
		_w6830_
	);
	LUT2 #(
		.INIT('h8)
	) name5651 (
		\g1092_reg/NET0131 ,
		_w6820_,
		_w6831_
	);
	LUT2 #(
		.INIT('h2)
	) name5652 (
		\g858_reg/NET0131 ,
		_w6831_,
		_w6832_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		_w6824_,
		_w6831_,
		_w6833_
	);
	LUT2 #(
		.INIT('h1)
	) name5654 (
		_w6832_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h2)
	) name5655 (
		\g1018_reg/NET0131 ,
		\g477_reg/NET0131 ,
		_w6835_
	);
	LUT2 #(
		.INIT('h2)
	) name5656 (
		\g1024_reg/NET0131 ,
		\g478_reg/NET0131 ,
		_w6836_
	);
	LUT2 #(
		.INIT('h4)
	) name5657 (
		\g479_reg/NET0131 ,
		\g5657_pad ,
		_w6837_
	);
	LUT2 #(
		.INIT('h1)
	) name5658 (
		_w6835_,
		_w6836_,
		_w6838_
	);
	LUT2 #(
		.INIT('h4)
	) name5659 (
		_w6837_,
		_w6838_,
		_w6839_
	);
	LUT2 #(
		.INIT('h2)
	) name5660 (
		\g2244_reg/NET0131 ,
		_w6821_,
		_w6840_
	);
	LUT2 #(
		.INIT('h1)
	) name5661 (
		\g2190_reg/NET0131 ,
		\g2195_reg/NET0131 ,
		_w6841_
	);
	LUT2 #(
		.INIT('h8)
	) name5662 (
		_w5141_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h8)
	) name5663 (
		_w6821_,
		_w6842_,
		_w6843_
	);
	LUT2 #(
		.INIT('h1)
	) name5664 (
		_w6840_,
		_w6843_,
		_w6844_
	);
	LUT2 #(
		.INIT('h2)
	) name5665 (
		\g2245_reg/NET0131 ,
		_w6827_,
		_w6845_
	);
	LUT2 #(
		.INIT('h8)
	) name5666 (
		_w6827_,
		_w6842_,
		_w6846_
	);
	LUT2 #(
		.INIT('h1)
	) name5667 (
		_w6845_,
		_w6846_,
		_w6847_
	);
	LUT2 #(
		.INIT('h2)
	) name5668 (
		\g2246_reg/NET0131 ,
		_w6831_,
		_w6848_
	);
	LUT2 #(
		.INIT('h8)
	) name5669 (
		_w6831_,
		_w6842_,
		_w6849_
	);
	LUT2 #(
		.INIT('h1)
	) name5670 (
		_w6848_,
		_w6849_,
		_w6850_
	);
	LUT2 #(
		.INIT('h2)
	) name5671 (
		\g1024_reg/NET0131 ,
		\g1165_reg/NET0131 ,
		_w6851_
	);
	LUT2 #(
		.INIT('h2)
	) name5672 (
		\g1018_reg/NET0131 ,
		\g1164_reg/NET0131 ,
		_w6852_
	);
	LUT2 #(
		.INIT('h4)
	) name5673 (
		\g1166_reg/NET0131 ,
		\g5657_pad ,
		_w6853_
	);
	LUT2 #(
		.INIT('h1)
	) name5674 (
		_w6851_,
		_w6852_,
		_w6854_
	);
	LUT2 #(
		.INIT('h4)
	) name5675 (
		_w6853_,
		_w6854_,
		_w6855_
	);
	LUT2 #(
		.INIT('h2)
	) name5676 (
		\g1018_reg/NET0131 ,
		\g480_reg/NET0131 ,
		_w6856_
	);
	LUT2 #(
		.INIT('h2)
	) name5677 (
		\g1024_reg/NET0131 ,
		\g484_reg/NET0131 ,
		_w6857_
	);
	LUT2 #(
		.INIT('h4)
	) name5678 (
		\g464_reg/NET0131 ,
		\g5657_pad ,
		_w6858_
	);
	LUT2 #(
		.INIT('h1)
	) name5679 (
		_w6856_,
		_w6857_,
		_w6859_
	);
	LUT2 #(
		.INIT('h4)
	) name5680 (
		_w6858_,
		_w6859_,
		_w6860_
	);
	LUT2 #(
		.INIT('h2)
	) name5681 (
		\g1018_reg/NET0131 ,
		\g1167_reg/NET0131 ,
		_w6861_
	);
	LUT2 #(
		.INIT('h2)
	) name5682 (
		\g1024_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		_w6862_
	);
	LUT2 #(
		.INIT('h4)
	) name5683 (
		\g1151_reg/NET0131 ,
		\g5657_pad ,
		_w6863_
	);
	LUT2 #(
		.INIT('h1)
	) name5684 (
		_w6861_,
		_w6862_,
		_w6864_
	);
	LUT2 #(
		.INIT('h4)
	) name5685 (
		_w6863_,
		_w6864_,
		_w6865_
	);
	LUT2 #(
		.INIT('h2)
	) name5686 (
		\g1018_reg/NET0131 ,
		\g1173_reg/NET0131 ,
		_w6866_
	);
	LUT2 #(
		.INIT('h2)
	) name5687 (
		\g1024_reg/NET0131 ,
		\g1174_reg/NET0131 ,
		_w6867_
	);
	LUT2 #(
		.INIT('h4)
	) name5688 (
		\g1175_reg/NET0131 ,
		\g5657_pad ,
		_w6868_
	);
	LUT2 #(
		.INIT('h1)
	) name5689 (
		_w6866_,
		_w6867_,
		_w6869_
	);
	LUT2 #(
		.INIT('h4)
	) name5690 (
		_w6868_,
		_w6869_,
		_w6870_
	);
	LUT2 #(
		.INIT('h1)
	) name5691 (
		\g2993_reg/NET0131 ,
		\g3080_reg/NET0131 ,
		_w6871_
	);
	LUT2 #(
		.INIT('h1)
	) name5692 (
		\g3234_pad ,
		_w6795_,
		_w6872_
	);
	LUT2 #(
		.INIT('h4)
	) name5693 (
		_w6871_,
		_w6872_,
		_w6873_
	);
	LUT2 #(
		.INIT('h2)
	) name5694 (
		\g1018_reg/NET0131 ,
		\g2552_reg/NET0131 ,
		_w6874_
	);
	LUT2 #(
		.INIT('h2)
	) name5695 (
		\g1024_reg/NET0131 ,
		\g2553_reg/NET0131 ,
		_w6875_
	);
	LUT2 #(
		.INIT('h4)
	) name5696 (
		\g2554_reg/NET0131 ,
		\g5657_pad ,
		_w6876_
	);
	LUT2 #(
		.INIT('h1)
	) name5697 (
		_w6874_,
		_w6875_,
		_w6877_
	);
	LUT2 #(
		.INIT('h4)
	) name5698 (
		_w6876_,
		_w6877_,
		_w6878_
	);
	LUT2 #(
		.INIT('h2)
	) name5699 (
		\g1018_reg/NET0131 ,
		\g2555_reg/NET0131 ,
		_w6879_
	);
	LUT2 #(
		.INIT('h2)
	) name5700 (
		\g1024_reg/NET0131 ,
		\g2559_reg/NET0131 ,
		_w6880_
	);
	LUT2 #(
		.INIT('h4)
	) name5701 (
		\g2539_reg/NET0131 ,
		\g5657_pad ,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name5702 (
		_w6879_,
		_w6880_,
		_w6882_
	);
	LUT2 #(
		.INIT('h4)
	) name5703 (
		_w6881_,
		_w6882_,
		_w6883_
	);
	LUT2 #(
		.INIT('h2)
	) name5704 (
		\g1018_reg/NET0131 ,
		\g2561_reg/NET0131 ,
		_w6884_
	);
	LUT2 #(
		.INIT('h2)
	) name5705 (
		\g1024_reg/NET0131 ,
		\g2562_reg/NET0131 ,
		_w6885_
	);
	LUT2 #(
		.INIT('h4)
	) name5706 (
		\g2563_reg/NET0131 ,
		\g5657_pad ,
		_w6886_
	);
	LUT2 #(
		.INIT('h1)
	) name5707 (
		_w6884_,
		_w6885_,
		_w6887_
	);
	LUT2 #(
		.INIT('h4)
	) name5708 (
		_w6886_,
		_w6887_,
		_w6888_
	);
	LUT2 #(
		.INIT('h2)
	) name5709 (
		\g1018_reg/NET0131 ,
		\g1861_reg/NET0131 ,
		_w6889_
	);
	LUT2 #(
		.INIT('h2)
	) name5710 (
		\g1024_reg/NET0131 ,
		\g1865_reg/NET0131 ,
		_w6890_
	);
	LUT2 #(
		.INIT('h4)
	) name5711 (
		\g1845_reg/NET0131 ,
		\g5657_pad ,
		_w6891_
	);
	LUT2 #(
		.INIT('h1)
	) name5712 (
		_w6889_,
		_w6890_,
		_w6892_
	);
	LUT2 #(
		.INIT('h4)
	) name5713 (
		_w6891_,
		_w6892_,
		_w6893_
	);
	LUT2 #(
		.INIT('h4)
	) name5714 (
		_w5147_,
		_w6821_,
		_w6894_
	);
	LUT2 #(
		.INIT('h2)
	) name5715 (
		\g2253_reg/NET0131 ,
		_w6821_,
		_w6895_
	);
	LUT2 #(
		.INIT('h1)
	) name5716 (
		_w6894_,
		_w6895_,
		_w6896_
	);
	LUT2 #(
		.INIT('h4)
	) name5717 (
		_w5147_,
		_w6827_,
		_w6897_
	);
	LUT2 #(
		.INIT('h2)
	) name5718 (
		\g2254_reg/NET0131 ,
		_w6827_,
		_w6898_
	);
	LUT2 #(
		.INIT('h1)
	) name5719 (
		_w6897_,
		_w6898_,
		_w6899_
	);
	LUT2 #(
		.INIT('h4)
	) name5720 (
		_w5147_,
		_w6831_,
		_w6900_
	);
	LUT2 #(
		.INIT('h2)
	) name5721 (
		\g2255_reg/NET0131 ,
		_w6831_,
		_w6901_
	);
	LUT2 #(
		.INIT('h1)
	) name5722 (
		_w6900_,
		_w6901_,
		_w6902_
	);
	LUT2 #(
		.INIT('h1)
	) name5723 (
		\g3006_reg/NET0131 ,
		_w6043_,
		_w6903_
	);
	LUT2 #(
		.INIT('h1)
	) name5724 (
		_w6044_,
		_w6903_,
		_w6904_
	);
	LUT2 #(
		.INIT('h8)
	) name5725 (
		_w6041_,
		_w6904_,
		_w6905_
	);
	LUT2 #(
		.INIT('h1)
	) name5726 (
		\g2883_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w6906_
	);
	LUT2 #(
		.INIT('h1)
	) name5727 (
		_w6529_,
		_w6906_,
		_w6907_
	);
	LUT2 #(
		.INIT('h2)
	) name5728 (
		_w6528_,
		_w6907_,
		_w6908_
	);
	LUT2 #(
		.INIT('h1)
	) name5729 (
		\g2892_reg/NET0131 ,
		_w6531_,
		_w6909_
	);
	LUT2 #(
		.INIT('h2)
	) name5730 (
		_w6528_,
		_w6532_,
		_w6910_
	);
	LUT2 #(
		.INIT('h4)
	) name5731 (
		_w6909_,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('h1)
	) name5732 (
		\g2903_reg/NET0131 ,
		_w6532_,
		_w6912_
	);
	LUT2 #(
		.INIT('h2)
	) name5733 (
		_w6528_,
		_w6533_,
		_w6913_
	);
	LUT2 #(
		.INIT('h4)
	) name5734 (
		_w6912_,
		_w6913_,
		_w6914_
	);
	LUT2 #(
		.INIT('h1)
	) name5735 (
		\g3013_reg/NET0131 ,
		_w6045_,
		_w6915_
	);
	LUT2 #(
		.INIT('h2)
	) name5736 (
		_w6041_,
		_w6046_,
		_w6916_
	);
	LUT2 #(
		.INIT('h4)
	) name5737 (
		_w6915_,
		_w6916_,
		_w6917_
	);
	LUT2 #(
		.INIT('h1)
	) name5738 (
		\g1326_reg/NET0131 ,
		_w5046_,
		_w6918_
	);
	LUT2 #(
		.INIT('h1)
	) name5739 (
		_w5045_,
		_w5047_,
		_w6919_
	);
	LUT2 #(
		.INIT('h4)
	) name5740 (
		_w6918_,
		_w6919_,
		_w6920_
	);
	LUT2 #(
		.INIT('h1)
	) name5741 (
		\g2888_reg/NET0131 ,
		_w6529_,
		_w6921_
	);
	LUT2 #(
		.INIT('h1)
	) name5742 (
		_w6530_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h8)
	) name5743 (
		_w6528_,
		_w6922_,
		_w6923_
	);
	LUT2 #(
		.INIT('h1)
	) name5744 (
		\g2896_reg/NET0131 ,
		_w6530_,
		_w6924_
	);
	LUT2 #(
		.INIT('h1)
	) name5745 (
		_w6531_,
		_w6924_,
		_w6925_
	);
	LUT2 #(
		.INIT('h8)
	) name5746 (
		_w6528_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h1)
	) name5747 (
		\g2933_reg/NET0131 ,
		\g51_pad ,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name5748 (
		\g3079_reg/NET0131 ,
		\g3234_pad ,
		_w6928_
	);
	LUT2 #(
		.INIT('h2)
	) name5749 (
		\g1024_reg/NET0131 ,
		_w5648_,
		_w6929_
	);
	LUT2 #(
		.INIT('h1)
	) name5750 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w6930_
	);
	LUT2 #(
		.INIT('h1)
	) name5751 (
		_w6929_,
		_w6930_,
		_w6931_
	);
	LUT2 #(
		.INIT('h2)
	) name5752 (
		\g1024_reg/NET0131 ,
		\g1240_reg/NET0131 ,
		_w6932_
	);
	LUT2 #(
		.INIT('h4)
	) name5753 (
		\g1024_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w6933_
	);
	LUT2 #(
		.INIT('h1)
	) name5754 (
		_w6932_,
		_w6933_,
		_w6934_
	);
	LUT2 #(
		.INIT('h4)
	) name5755 (
		\g291_reg/NET0131 ,
		\g3229_pad ,
		_w6935_
	);
	LUT2 #(
		.INIT('h2)
	) name5756 (
		\g305_reg/NET0131 ,
		\g3229_pad ,
		_w6936_
	);
	LUT2 #(
		.INIT('h1)
	) name5757 (
		_w6935_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h2)
	) name5758 (
		\g3229_pad ,
		\g978_reg/NET0131 ,
		_w6938_
	);
	LUT2 #(
		.INIT('h4)
	) name5759 (
		\g3229_pad ,
		\g992_reg/NET0131 ,
		_w6939_
	);
	LUT2 #(
		.INIT('h1)
	) name5760 (
		_w6938_,
		_w6939_,
		_w6940_
	);
	LUT2 #(
		.INIT('h2)
	) name5761 (
		\g2814_reg/NET0131 ,
		\g2929_reg/NET0131 ,
		_w6941_
	);
	LUT2 #(
		.INIT('h2)
	) name5762 (
		\g2879_reg/NET0131 ,
		_w6941_,
		_w6942_
	);
	LUT2 #(
		.INIT('h4)
	) name5763 (
		\g1672_reg/NET0131 ,
		\g3229_pad ,
		_w6943_
	);
	LUT2 #(
		.INIT('h2)
	) name5764 (
		\g1686_reg/NET0131 ,
		\g3229_pad ,
		_w6944_
	);
	LUT2 #(
		.INIT('h1)
	) name5765 (
		_w6943_,
		_w6944_,
		_w6945_
	);
	LUT2 #(
		.INIT('h4)
	) name5766 (
		\g2366_reg/NET0131 ,
		\g3229_pad ,
		_w6946_
	);
	LUT2 #(
		.INIT('h2)
	) name5767 (
		\g2380_reg/NET0131 ,
		\g3229_pad ,
		_w6947_
	);
	LUT2 #(
		.INIT('h1)
	) name5768 (
		_w6946_,
		_w6947_,
		_w6948_
	);
	LUT2 #(
		.INIT('h2)
	) name5769 (
		\g2817_reg/NET0131 ,
		\g51_pad ,
		_w6949_
	);
	LUT2 #(
		.INIT('h2)
	) name5770 (
		\g3054_reg/NET0131 ,
		\g3234_pad ,
		_w6950_
	);
	LUT2 #(
		.INIT('h1)
	) name5771 (
		\g117_reg/NET0131 ,
		\g121_reg/NET0131 ,
		_w6951_
	);
	LUT2 #(
		.INIT('h8)
	) name5772 (
		_w5110_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h1)
	) name5773 (
		\g1496_reg/NET0131 ,
		\g1501_reg/NET0131 ,
		_w6953_
	);
	LUT2 #(
		.INIT('h8)
	) name5774 (
		_w5172_,
		_w6953_,
		_w6954_
	);
	LUT2 #(
		.INIT('h2)
	) name5775 (
		\g2950_reg/NET0131 ,
		\g51_pad ,
		_w6955_
	);
	LUT2 #(
		.INIT('h2)
	) name5776 (
		\g3080_reg/NET0131 ,
		\g3234_pad ,
		_w6956_
	);
	LUT2 #(
		.INIT('h1)
	) name5777 (
		_w2175_,
		_w3560_,
		_w6957_
	);
	LUT2 #(
		.INIT('h8)
	) name5778 (
		_w2175_,
		_w3560_,
		_w6958_
	);
	LUT2 #(
		.INIT('h1)
	) name5779 (
		_w6957_,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h8)
	) name5780 (
		_w3099_,
		_w6959_,
		_w6960_
	);
	LUT2 #(
		.INIT('h1)
	) name5781 (
		\g121_reg/NET0131 ,
		_w3075_,
		_w6961_
	);
	LUT2 #(
		.INIT('h1)
	) name5782 (
		_w3095_,
		_w6961_,
		_w6962_
	);
	LUT2 #(
		.INIT('h4)
	) name5783 (
		_w6960_,
		_w6962_,
		_w6963_
	);
	LUT2 #(
		.INIT('h2)
	) name5784 (
		\g2190_reg/NET0131 ,
		_w3331_,
		_w6964_
	);
	LUT2 #(
		.INIT('h2)
	) name5785 (
		_w1330_,
		_w3420_,
		_w6965_
	);
	LUT2 #(
		.INIT('h4)
	) name5786 (
		_w1330_,
		_w3420_,
		_w6966_
	);
	LUT2 #(
		.INIT('h1)
	) name5787 (
		_w6965_,
		_w6966_,
		_w6967_
	);
	LUT2 #(
		.INIT('h8)
	) name5788 (
		_w3336_,
		_w6967_,
		_w6968_
	);
	LUT2 #(
		.INIT('h1)
	) name5789 (
		_w6964_,
		_w6968_,
		_w6969_
	);
	LUT2 #(
		.INIT('h2)
	) name5790 (
		\g1088_reg/NET0131 ,
		_w3501_,
		_w6970_
	);
	LUT2 #(
		.INIT('h1)
	) name5791 (
		\g1088_reg/NET0131 ,
		\g246_reg/NET0131 ,
		_w6971_
	);
	LUT2 #(
		.INIT('h1)
	) name5792 (
		_w6970_,
		_w6971_,
		_w6972_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g101_reg/P0001  = \g101_reg/NET0131 ;
	assign \g105_reg/P0001  = \g105_reg/NET0131 ;
	assign \g109_reg/P0001  = \g109_reg/NET0131 ;
	assign \g1138_reg/P0001  = \g1138_reg/NET0131 ;
	assign \g113_reg/P0001  = \g113_reg/NET0131 ;
	assign \g1140_reg/P0001  = \g1140_reg/NET0131 ;
	assign \g117_reg/P0001  = \g117_reg/NET0131 ;
	assign \g121_reg/P0001  = \g121_reg/NET0131 ;
	assign \g125_reg/P0001  = \g125_reg/NET0131 ;
	assign \g1471_reg/P0001  = \g1471_reg/NET0131 ;
	assign \g1476_reg/P0001  = \g1476_reg/NET0131 ;
	assign \g1481_reg/P0001  = \g1481_reg/NET0131 ;
	assign \g1486_reg/P0001  = \g1486_reg/NET0131 ;
	assign \g1491_reg/P0001  = \g1491_reg/NET0131 ;
	assign \g1496_reg/P0001  = \g1496_reg/NET0131 ;
	assign \g1501_reg/P0001  = \g1501_reg/NET0131 ;
	assign \g1506_reg/P0001  = \g1506_reg/NET0131 ;
	assign \g16496_pad  = _w1181_ ;
	assign \g1660_reg/P0001  = \g1660_reg/NET0131 ;
	assign \g1662_reg/P0001  = \g1662_reg/NET0131 ;
	assign \g1664_reg/P0001  = \g1664_reg/NET0131 ;
	assign \g1666_reg/P0001  = \g1666_reg/NET0131 ;
	assign \g1668_reg/P0001  = \g1668_reg/NET0131 ;
	assign \g1670_reg/P0001  = \g1670_reg/NET0131 ;
	assign \g1672_reg/P0001  = \g1672_reg/NET0131 ;
	assign \g18/_0_  = _w1450_ ;
	assign \g1832_reg/P0001  = \g1832_reg/NET0131 ;
	assign \g1834_reg/P0001  = \g1834_reg/NET0131 ;
	assign \g2165_reg/P0001  = \g2165_reg/NET0131 ;
	assign \g2170_reg/P0001  = \g2170_reg/NET0131 ;
	assign \g2175_reg/P0001  = \g2175_reg/NET0131 ;
	assign \g2180_reg/P0001  = \g2180_reg/NET0131 ;
	assign \g2185_reg/P0001  = \g2185_reg/NET0131 ;
	assign \g2190_reg/P0001  = \g2190_reg/NET0131 ;
	assign \g2195_reg/P0001  = \g2195_reg/NET0131 ;
	assign \g2200_reg/P0001  = \g2200_reg/NET0131 ;
	assign \g2354_reg/P0001  = \g2354_reg/NET0131 ;
	assign \g2356_reg/P0001  = \g2356_reg/NET0131 ;
	assign \g2358_reg/P0001  = \g2358_reg/NET0131 ;
	assign \g2360_reg/P0001  = \g2360_reg/NET0131 ;
	assign \g2362_reg/P0001  = \g2362_reg/NET0131 ;
	assign \g2364_reg/P0001  = \g2364_reg/NET0131 ;
	assign \g2366_reg/P0001  = \g2366_reg/NET0131 ;
	assign \g2526_reg/P0001  = \g2526_reg/NET0131 ;
	assign \g2528_reg/P0001  = \g2528_reg/NET0131 ;
	assign \g25489_pad  = _w1461_ ;
	assign \g279_reg/P0001  = \g279_reg/NET0131 ;
	assign \g281_reg/P0001  = \g281_reg/NET0131 ;
	assign \g283_reg/P0001  = \g283_reg/NET0131 ;
	assign \g285_reg/P0001  = \g285_reg/NET0131 ;
	assign \g2879_reg/NET0131_syn_2  = \g2879_reg/NET0131 ;
	assign \g287_reg/P0001  = \g287_reg/NET0131 ;
	assign \g289_reg/P0001  = \g289_reg/NET0131 ;
	assign \g291_reg/P0001  = \g291_reg/NET0131 ;
	assign \g451_reg/P0001  = \g451_reg/NET0131 ;
	assign \g453_reg/P0001  = \g453_reg/NET0131 ;
	assign \g59421/_3_  = _w1466_ ;
	assign \g59425/_1_  = _w1469_ ;
	assign \g59435/_0_  = _w1493_ ;
	assign \g59436/_0_  = _w1497_ ;
	assign \g59441/_3_  = _w1500_ ;
	assign \g59442/_0_  = _w1524_ ;
	assign \g59445/_0_  = _w1527_ ;
	assign \g59453/_0_  = _w1710_ ;
	assign \g59462/_3_  = _w1713_ ;
	assign \g59466/_3_  = _w1716_ ;
	assign \g59467/_3_  = _w1719_ ;
	assign \g59468/_3_  = _w1722_ ;
	assign \g59469/_3_  = _w1725_ ;
	assign \g59470/_3_  = _w1728_ ;
	assign \g59471/_3_  = _w1731_ ;
	assign \g59472/_3_  = _w1734_ ;
	assign \g59473/_3_  = _w1737_ ;
	assign \g59489/_0_  = _w1900_ ;
	assign \g59498/_0_  = _w1919_ ;
	assign \g59499/_0_  = _w1925_ ;
	assign \g59500/_0_  = _w1932_ ;
	assign \g59502/_2_  = _w1940_ ;
	assign \g59503/_0_  = _w1946_ ;
	assign \g59505/_2_  = _w1952_ ;
	assign \g59507/_0_  = _w1959_ ;
	assign \g59508/_0_  = _w1966_ ;
	assign \g59533/_3_  = _w1969_ ;
	assign \g59534/_3_  = _w1972_ ;
	assign \g59535/_3_  = _w1975_ ;
	assign \g59536/_3_  = _w1978_ ;
	assign \g59537/_3_  = _w1981_ ;
	assign \g59538/_3_  = _w1984_ ;
	assign \g59539/_3_  = _w1987_ ;
	assign \g59540/_3_  = _w1990_ ;
	assign \g59548/_0_  = _w2009_ ;
	assign \g59550/_0_  = _w2277_ ;
	assign \g59551/_0_  = _w2280_ ;
	assign \g59552/_0_  = _w2283_ ;
	assign \g59554/_0_  = _w2557_ ;
	assign \g59555/_0_  = _w2560_ ;
	assign \g59556/_0_  = _w2563_ ;
	assign \g59557/_0_  = _w2566_ ;
	assign \g59558/_0_  = _w2569_ ;
	assign \g59559/_0_  = _w2843_ ;
	assign \g59560/_0_  = _w2846_ ;
	assign \g59561/_0_  = _w2849_ ;
	assign \g59639/_0_  = _w3012_ ;
	assign \g59694/_2_  = _w3029_ ;
	assign \g59695/_0_  = _w3037_ ;
	assign \g59697/_2_  = _w3043_ ;
	assign \g59698/_0_  = _w3049_ ;
	assign \g59699/_0_  = _w3056_ ;
	assign \g59700/_0_  = _w3062_ ;
	assign \g59705/_0_  = _w3115_ ;
	assign \g59706/_0_  = _w3118_ ;
	assign \g59707/_0_  = _w3121_ ;
	assign \g59708/_0_  = _w3168_ ;
	assign \g59709/_0_  = _w3171_ ;
	assign \g59710/_0_  = _w3174_ ;
	assign \g59711/_0_  = _w3187_ ;
	assign \g59712/_0_  = _w3190_ ;
	assign \g59713/_0_  = _w3193_ ;
	assign \g59714/_0_  = _w3206_ ;
	assign \g59715/_0_  = _w3209_ ;
	assign \g59716/_0_  = _w3212_ ;
	assign \g59717/_0_  = _w3243_ ;
	assign \g59718/_0_  = _w3246_ ;
	assign \g59719/_0_  = _w3249_ ;
	assign \g59720/_0_  = _w3298_ ;
	assign \g59721/_0_  = _w3350_ ;
	assign \g59722/_0_  = _w3353_ ;
	assign \g59723/_0_  = _w3356_ ;
	assign \g59724/_0_  = _w3359_ ;
	assign \g59725/_0_  = _w3372_ ;
	assign \g59726/_0_  = _w3375_ ;
	assign \g59727/_0_  = _w3378_ ;
	assign \g59728/_0_  = _w3381_ ;
	assign \g59729/_0_  = _w3395_ ;
	assign \g59730/_0_  = _w3398_ ;
	assign \g59731/_0_  = _w3408_ ;
	assign \g59732/_0_  = _w3411_ ;
	assign \g59733/_0_  = _w3441_ ;
	assign \g59734/_0_  = _w3444_ ;
	assign \g59735/_0_  = _w3447_ ;
	assign \g59736/_0_  = _w3450_ ;
	assign \g59737/_0_  = _w3453_ ;
	assign \g59738/_0_  = _w3466_ ;
	assign \g59739/_0_  = _w3469_ ;
	assign \g59740/_0_  = _w3472_ ;
	assign \g59741/_0_  = _w3486_ ;
	assign \g59742/_0_  = _w3489_ ;
	assign \g59743/_0_  = _w3504_ ;
	assign \g59744/_0_  = _w3507_ ;
	assign \g59745/_0_  = _w3510_ ;
	assign \g59747/_0_  = _w3539_ ;
	assign \g59748/_0_  = _w3542_ ;
	assign \g59749/_0_  = _w3545_ ;
	assign \g59750/_0_  = _w3578_ ;
	assign \g59751/_0_  = _w3581_ ;
	assign \g59752/_0_  = _w3584_ ;
	assign \g59753/_0_  = _w3591_ ;
	assign \g59754/_0_  = _w3598_ ;
	assign \g59755/_0_  = _w3608_ ;
	assign \g59756/_0_  = _w3611_ ;
	assign \g59757/_0_  = _w3614_ ;
	assign \g59758/_0_  = _w3624_ ;
	assign \g59759/_0_  = _w3627_ ;
	assign \g59760/_0_  = _w3630_ ;
	assign \g59761/_0_  = _w3640_ ;
	assign \g59762/_0_  = _w3643_ ;
	assign \g59763/_0_  = _w3646_ ;
	assign \g59764/_0_  = _w3656_ ;
	assign \g59765/_0_  = _w3659_ ;
	assign \g59766/_0_  = _w3662_ ;
	assign \g59915/_0_  = _w3830_ ;
	assign \g59952/_2_  = _w2005_ ;
	assign \g60046/_0_  = _w3840_ ;
	assign \g60048/_0_  = _w3847_ ;
	assign \g60049/_0_  = _w3854_ ;
	assign \g60051/_0_  = _w3861_ ;
	assign \g60063/_0_  = _w3880_ ;
	assign \g60103/_0_  = _w3886_ ;
	assign \g60104/_0_  = _w3893_ ;
	assign \g60105/_0_  = _w3909_ ;
	assign \g60107/_2_  = _w3918_ ;
	assign \g60108/_0_  = _w3924_ ;
	assign \g60109/_0_  = _w3931_ ;
	assign \g60110/_0_  = _w3937_ ;
	assign \g60112/_2_  = _w3943_ ;
	assign \g60119/_0_  = _w3949_ ;
	assign \g60120/_0_  = _w3956_ ;
	assign \g60121/_0_  = _w3963_ ;
	assign \g60122/_0_  = _w3968_ ;
	assign \g60123/_0_  = _w3973_ ;
	assign \g60124/_0_  = _w3979_ ;
	assign \g60126/_0_  = _w3984_ ;
	assign \g60127/_0_  = _w3993_ ;
	assign \g60128/_0_  = _w3999_ ;
	assign \g60129/_0_  = _w4005_ ;
	assign \g60130/_0_  = _w4013_ ;
	assign \g60135/_0_  = _w4022_ ;
	assign \g60136/_0_  = _w4028_ ;
	assign \g60137/_0_  = _w4034_ ;
	assign \g60138/_0_  = _w4040_ ;
	assign \g60139/_0_  = _w4046_ ;
	assign \g60143/_3_  = _w1547_ ;
	assign \g60144/_0_  = _w4053_ ;
	assign \g60145/_0_  = _w4060_ ;
	assign \g60339/_0_  = _w2001_ ;
	assign \g60404/_0_  = _w4064_ ;
	assign \g60427/_0_  = _w4068_ ;
	assign \g60428/_0_  = _w4072_ ;
	assign \g60429/_0_  = _w4076_ ;
	assign \g60434/_0_  = _w4093_ ;
	assign \g60435/_0_  = _w4099_ ;
	assign \g60437/_0_  = _w4107_ ;
	assign \g60438/_0_  = _w4113_ ;
	assign \g60439/_0_  = _w4120_ ;
	assign \g60440/_0_  = _w4126_ ;
	assign \g60441/_0_  = _w3876_ ;
	assign \g60448/_0_  = _w4281_ ;
	assign \g60451/_0_  = _w4429_ ;
	assign \g60452/_0_  = _w4432_ ;
	assign \g60453/_0_  = _w4435_ ;
	assign \g60459/_0_  = _w4442_ ;
	assign \g60460/_0_  = _w4449_ ;
	assign \g60523/_0_  = _w1542_ ;
	assign \g60534/_0_  = _w4458_ ;
	assign \g60535/_0_  = _w4461_ ;
	assign \g60536/_0_  = _w4464_ ;
	assign \g60585/_0_  = _w4467_ ;
	assign \g60586/_0_  = _w4469_ ;
	assign \g60587/_0_  = _w4472_ ;
	assign \g60588/_0_  = _w4475_ ;
	assign \g60591/_0_  = _w4527_ ;
	assign \g60592/_0_  = _w4531_ ;
	assign \g60599/_0_  = _w4583_ ;
	assign \g60601/_0_  = _w4587_ ;
	assign \g60602/_0_  = _w4591_ ;
	assign \g60603/_0_  = _w4643_ ;
	assign \g60604/_0_  = _w4695_ ;
	assign \g60605/_0_  = _w4699_ ;
	assign \g60606/_0_  = _w4703_ ;
	assign \g60607/_0_  = _w4707_ ;
	assign \g60608/_0_  = _w4711_ ;
	assign \g60609/_0_  = _w4715_ ;
	assign \g60613/_0_  = _w4859_ ;
	assign \g60614/_0_  = _w5003_ ;
	assign \g60615/_0_  = _w4278_ ;
	assign \g60694/_0_  = _w5006_ ;
	assign \g60708/_0_  = _w5011_ ;
	assign \g60709/_0_  = _w5017_ ;
	assign \g60710/_0_  = _w5022_ ;
	assign \g60785/_0_  = _w5026_ ;
	assign \g60787/_0_  = _w5028_ ;
	assign \g60788/_0_  = _w5030_ ;
	assign \g60799/_0_  = _w5033_ ;
	assign \g60801/_0_  = _w5034_ ;
	assign \g60802/_0_  = _w5035_ ;
	assign \g60803/_1__syn_2  = _w5038_ ;
	assign \g60805/_1__syn_2  = _w5039_ ;
	assign \g60806/_1__syn_2  = _w5040_ ;
	assign \g60808/_0_  = _w5042_ ;
	assign \g60810/_0_  = _w5043_ ;
	assign \g60811/_0_  = _w5044_ ;
	assign \g60825/_3_  = _w3872_ ;
	assign \g60896/_0_  = _w5059_ ;
	assign \g60980/_0_  = _w5090_ ;
	assign \g60981/_0_  = _w5121_ ;
	assign \g60985/_0_  = _w5152_ ;
	assign \g60986/_0_  = _w5183_ ;
	assign \g61012/_0_  = _w5184_ ;
	assign \g61013/_0_  = _w5185_ ;
	assign \g61015/_0_  = _w5186_ ;
	assign \g61017/_0_  = _w5187_ ;
	assign \g61122/_0_  = _w5195_ ;
	assign \g61123/_0_  = _w5203_ ;
	assign \g61124/_0_  = _w5211_ ;
	assign \g61125/_0_  = _w5219_ ;
	assign \g61222/_0_  = _w5220_ ;
	assign \g61223/_0_  = _w5221_ ;
	assign \g61224/_0_  = _w5222_ ;
	assign \g61225/_0_  = _w5223_ ;
	assign \g61228/_0_  = _w5224_ ;
	assign \g61229/_0_  = _w5225_ ;
	assign \g61230/_0_  = _w5226_ ;
	assign \g61231/_0_  = _w5227_ ;
	assign \g61281/_0_  = _w5230_ ;
	assign \g61293/_1_  = _w5232_ ;
	assign \g61307/_0__syn_2  = _w5233_ ;
	assign \g61309/_0__syn_2  = _w5234_ ;
	assign \g61310/_0__syn_2  = _w5235_ ;
	assign \g61311/_1_  = _w5236_ ;
	assign \g61312/_1_  = _w5237_ ;
	assign \g61313/_1_  = _w5238_ ;
	assign \g61324/_1_  = _w5239_ ;
	assign \g61325/_1_  = _w5240_ ;
	assign \g61326/_1_  = _w5241_ ;
	assign \g61328/_1_  = _w5242_ ;
	assign \g61329/_1_  = _w5243_ ;
	assign \g61330/_1_  = _w5244_ ;
	assign \g61332/_1_  = _w5293_ ;
	assign \g61333/_1_  = _w5338_ ;
	assign \g61334/_1_  = _w5383_ ;
	assign \g61335/_1_  = _w5428_ ;
	assign \g61336/_0_  = _w5445_ ;
	assign \g61338/_0_  = _w5462_ ;
	assign \g61339/_0_  = _w5465_ ;
	assign \g61340/_0_  = _w5468_ ;
	assign \g61377/_1_  = _w5490_ ;
	assign \g61378/_1_  = _w5491_ ;
	assign \g61379/_1_  = _w5492_ ;
	assign \g61388/_1_  = _w5526_ ;
	assign \g61391/_0_  = _w5541_ ;
	assign \g61394/_1_  = _w5542_ ;
	assign \g61395/_1_  = _w5543_ ;
	assign \g61396/_1_  = _w5565_ ;
	assign \g61398/_1_  = _w5566_ ;
	assign \g61399/_1_  = _w5567_ ;
	assign \g61421/_1_  = _w5601_ ;
	assign \g61422/_1_  = _w5602_ ;
	assign \g61423/_1_  = _w5603_ ;
	assign \g61524/_0_  = _w5630_ ;
	assign \g61525/_0_  = _w5634_ ;
	assign \g61526/_0_  = _w5638_ ;
	assign \g61527/_0_  = _w5663_ ;
	assign \g61528/_0_  = _w5667_ ;
	assign \g61529/_0_  = _w5671_ ;
	assign \g61530/_0_  = _w5705_ ;
	assign \g61531/_0_  = _w5709_ ;
	assign \g61532/_0_  = _w5713_ ;
	assign \g61533/_0_  = _w5723_ ;
	assign \g61534/_0_  = _w5726_ ;
	assign \g61535/_0_  = _w5729_ ;
	assign \g61536/_0_  = _w5750_ ;
	assign \g61537/_0_  = _w5754_ ;
	assign \g61538/_0_  = _w5758_ ;
	assign \g61539/_0_  = _w5761_ ;
	assign \g61540/_0_  = _w5781_ ;
	assign \g61541/_0_  = _w5785_ ;
	assign \g61542/_0_  = _w5789_ ;
	assign \g61543/_0_  = _w5798_ ;
	assign \g61544/_0_  = _w5831_ ;
	assign \g61545/_0_  = _w5834_ ;
	assign \g61546/_0_  = _w5837_ ;
	assign \g61547/_0_  = _w5841_ ;
	assign \g61548/_0_  = _w5845_ ;
	assign \g61549/_0_  = _w5855_ ;
	assign \g61550/_0_  = _w5858_ ;
	assign \g61551/_0_  = _w5861_ ;
	assign \g61552/_0_  = _w5877_ ;
	assign \g61553/_0_  = _w5897_ ;
	assign \g61554/_0_  = _w5930_ ;
	assign \g61555/_0_  = _w5934_ ;
	assign \g61556/_0_  = _w5938_ ;
	assign \g61557/_0_  = _w5946_ ;
	assign \g61558/_0_  = _w5949_ ;
	assign \g61559/_0_  = _w5952_ ;
	assign \g61560/_0_  = _w5956_ ;
	assign \g61561/_0_  = _w5960_ ;
	assign \g61562/_0_  = _w5970_ ;
	assign \g61563/_0_  = _w5973_ ;
	assign \g61564/_0_  = _w5976_ ;
	assign \g61565/_0_  = _w5979_ ;
	assign \g61566/_0_  = _w5982_ ;
	assign \g61620/_0_  = _w5986_ ;
	assign \g61621/_0_  = _w5990_ ;
	assign \g61622/_0_  = _w5994_ ;
	assign \g61623/_0_  = _w5998_ ;
	assign \g61753/_0_  = _w6000_ ;
	assign \g61764/_0_  = _w6002_ ;
	assign \g61786/_0_  = _w6004_ ;
	assign \g61795/_0_  = _w6006_ ;
	assign \g61801/_0_  = _w6016_ ;
	assign \g61803/_0_  = _w6018_ ;
	assign \g61808/_0_  = _w6020_ ;
	assign \g61848/_0_  = _w6023_ ;
	assign \g61850/_0_  = _w6026_ ;
	assign \g61851/_0_  = _w5442_ ;
	assign \g62097/_0_  = _w6030_ ;
	assign \g62102/_0_  = _w6034_ ;
	assign \g62115/_0_  = _w6037_ ;
	assign \g62119/_0_  = _w5485_ ;
	assign \g62130/_1_  = _w5710_ ;
	assign \g62131/_0_  = _w6040_ ;
	assign \g62132/_0_  = _w6051_ ;
	assign \g62139/_1_  = _w5751_ ;
	assign \g62140/_1_  = _w5653_ ;
	assign \g62141/_1_  = _w5664_ ;
	assign \g62144/_0_  = _w6056_ ;
	assign \g62145/_0_  = _w6059_ ;
	assign \g62146/_0_  = _w6062_ ;
	assign \g62147/_0_  = _w6065_ ;
	assign \g62150/_0_  = _w6068_ ;
	assign \g62151/_1_  = _w5674_ ;
	assign \g62152/_0_  = _w6071_ ;
	assign \g62153/_1_  = _w5706_ ;
	assign \g62156/_1_  = _w5668_ ;
	assign \g62157/_0_  = _w5520_ ;
	assign \g62159/_0_  = _w5560_ ;
	assign \g62161/_0_  = _w6076_ ;
	assign \g62187/_1_  = _w5772_ ;
	assign \g62190/_1_  = _w5782_ ;
	assign \g62191/_1_  = _w5740_ ;
	assign \g62192/_1_  = _w5786_ ;
	assign \g62194/_1_  = _w5800_ ;
	assign \g62195/_1_  = _w5838_ ;
	assign \g62196/_1_  = _w5842_ ;
	assign \g62203/_0_  = _w5595_ ;
	assign \g62204/_1_  = _w5755_ ;
	assign \g62207/_0__syn_2  = _w5888_ ;
	assign \g62208/_1_  = _w5899_ ;
	assign \g62209/_1_  = _w5931_ ;
	assign \g62210/_1_  = _w5935_ ;
	assign \g62211/_1_  = _w5953_ ;
	assign \g62212/_1_  = _w5957_ ;
	assign \g62217/_0_  = _w6079_ ;
	assign \g62286/_0_  = _w6096_ ;
	assign \g62287/_0_  = _w6098_ ;
	assign \g62288/_0_  = _w6101_ ;
	assign \g62289/_0_  = _w6104_ ;
	assign \g62290/_0_  = _w6106_ ;
	assign \g62291/_0_  = _w6108_ ;
	assign \g62292/_0_  = _w6110_ ;
	assign \g62435/_0_  = _w6113_ ;
	assign \g62436/_0_  = _w6116_ ;
	assign \g62439/_0_  = _w6119_ ;
	assign \g62456/_0_  = _w6122_ ;
	assign \g62486/_1_  = _w5605_ ;
	assign \g62492/_1_  = _w5631_ ;
	assign \g62494/_0_  = _w6125_ ;
	assign \g62495/_1_  = _w5635_ ;
	assign \g62497/_0_  = _w6128_ ;
	assign \g62537/_0_  = _w6132_ ;
	assign \g62544/_0_  = _w5652_ ;
	assign \g62546/_0_  = _w5739_ ;
	assign \g62547/_0_  = _w5771_ ;
	assign \g62549/_3_  = _w5887_ ;
	assign \g62552/_0_  = _w6133_ ;
	assign \g62554/_0_  = _w6137_ ;
	assign \g62555/_0_  = _w6138_ ;
	assign \g62556/_0_  = _w6142_ ;
	assign \g62558/_0_  = _w6146_ ;
	assign \g62559/_0_  = _w6147_ ;
	assign \g62561/_0_  = _w6151_ ;
	assign \g62562/_0_  = _w6152_ ;
	assign \g62566/_0_  = _w6155_ ;
	assign \g62567/_0_  = _w6158_ ;
	assign \g62568/_0_  = _w6160_ ;
	assign \g62569/_0_  = _w6163_ ;
	assign \g62570/_0_  = _w6165_ ;
	assign \g62571/_0_  = _w6168_ ;
	assign \g62572/_0_  = _w6171_ ;
	assign \g62573/_0_  = _w6174_ ;
	assign \g62574/_0_  = _w6177_ ;
	assign \g62575/_0_  = _w6180_ ;
	assign \g62576/_0_  = _w6183_ ;
	assign \g62577/_0_  = _w6186_ ;
	assign \g62578/_0_  = _w6189_ ;
	assign \g62579/_0_  = _w6192_ ;
	assign \g62580/_0_  = _w6195_ ;
	assign \g62581/_0_  = _w6198_ ;
	assign \g62582/_0_  = _w6201_ ;
	assign \g62583/_0_  = _w6204_ ;
	assign \g62584/_0_  = _w6207_ ;
	assign \g62585/_0_  = _w6210_ ;
	assign \g62586/_0_  = _w6213_ ;
	assign \g62587/_0_  = _w6216_ ;
	assign \g62588/_0_  = _w6219_ ;
	assign \g62589/_0_  = _w6222_ ;
	assign \g62590/_0_  = _w6225_ ;
	assign \g62591/_0_  = _w6228_ ;
	assign \g62592/_0_  = _w6231_ ;
	assign \g62593/_0_  = _w6234_ ;
	assign \g62594/_0_  = _w6237_ ;
	assign \g62595/_0_  = _w6240_ ;
	assign \g62596/_0_  = _w6243_ ;
	assign \g62597/_0_  = _w6246_ ;
	assign \g62602/_0_  = _w6249_ ;
	assign \g62607/_0_  = _w6252_ ;
	assign \g62608/_0_  = _w6255_ ;
	assign \g62609/_0_  = _w6258_ ;
	assign \g62619/_0_  = _w6261_ ;
	assign \g62620/_0_  = _w6264_ ;
	assign \g62621/_0_  = _w6267_ ;
	assign \g62622/_0_  = _w6270_ ;
	assign \g62623/_0_  = _w6273_ ;
	assign \g62624/_0_  = _w6276_ ;
	assign \g62626/_0_  = _w6279_ ;
	assign \g62627/_0_  = _w6282_ ;
	assign \g62628/_0_  = _w6285_ ;
	assign \g62629/_0_  = _w6288_ ;
	assign \g62630/_0_  = _w6291_ ;
	assign \g62631/_0_  = _w6294_ ;
	assign \g62632/_0_  = _w6297_ ;
	assign \g62633/_0_  = _w6300_ ;
	assign \g62634/_0_  = _w6303_ ;
	assign \g62635/_0_  = _w6306_ ;
	assign \g62636/_0_  = _w6309_ ;
	assign \g62637/_0_  = _w6312_ ;
	assign \g62638/_0_  = _w6315_ ;
	assign \g62639/_0_  = _w6318_ ;
	assign \g62640/_0_  = _w6321_ ;
	assign \g62641/_0_  = _w6324_ ;
	assign \g62642/_0_  = _w6327_ ;
	assign \g62643/_0_  = _w6330_ ;
	assign \g62644/_0_  = _w6333_ ;
	assign \g62645/_0_  = _w6336_ ;
	assign \g62646/_0_  = _w6339_ ;
	assign \g62647/_0_  = _w6342_ ;
	assign \g62648/_0_  = _w6345_ ;
	assign \g62649/_0_  = _w6348_ ;
	assign \g62650/_0_  = _w6351_ ;
	assign \g62651/_0_  = _w6354_ ;
	assign \g62652/_0_  = _w6357_ ;
	assign \g62653/_0_  = _w6360_ ;
	assign \g62654/_0_  = _w6363_ ;
	assign \g62655/_0_  = _w6366_ ;
	assign \g62656/_0_  = _w6369_ ;
	assign \g62657/_0_  = _w6372_ ;
	assign \g62658/_0_  = _w6375_ ;
	assign \g62659/_0_  = _w6378_ ;
	assign \g62660/_0_  = _w6381_ ;
	assign \g62661/_0_  = _w6383_ ;
	assign \g62674/_0_  = _w6386_ ;
	assign \g62682/_0_  = _w6389_ ;
	assign \g62683/_0_  = _w6391_ ;
	assign \g62689/_0_  = _w6394_ ;
	assign \g62690/_0_  = _w6397_ ;
	assign \g62691/_0_  = _w6400_ ;
	assign \g62694/_0_  = _w6403_ ;
	assign \g62695/_0_  = _w6406_ ;
	assign \g62696/_0_  = _w6409_ ;
	assign \g62698/_0_  = _w6412_ ;
	assign \g62699/_0_  = _w6415_ ;
	assign \g62700/_0_  = _w6418_ ;
	assign \g62723/_0_  = _w6421_ ;
	assign \g62724/_0_  = _w6424_ ;
	assign \g62725/_0_  = _w6427_ ;
	assign \g62726/_0_  = _w6430_ ;
	assign \g62727/_0_  = _w6433_ ;
	assign \g62728/_0_  = _w6436_ ;
	assign \g62735/_0_  = _w6439_ ;
	assign \g62736/_0_  = _w6442_ ;
	assign \g62737/_0_  = _w6445_ ;
	assign \g62738/_0_  = _w6448_ ;
	assign \g62739/_0_  = _w6451_ ;
	assign \g62740/_0_  = _w6454_ ;
	assign \g62754/_0_  = _w6457_ ;
	assign \g62762/_0_  = _w6460_ ;
	assign \g62763/_0_  = _w6463_ ;
	assign \g62764/_0_  = _w6466_ ;
	assign \g62780/_0_  = _w6469_ ;
	assign \g62781/_0_  = _w6472_ ;
	assign \g62785/_0_  = _w6475_ ;
	assign \g62786/_0_  = _w6478_ ;
	assign \g62787/_0_  = _w6481_ ;
	assign \g62791/_0_  = _w6484_ ;
	assign \g62792/_0_  = _w6487_ ;
	assign \g62794/_0_  = _w6490_ ;
	assign \g62804/_0_  = _w6492_ ;
	assign \g62806/_0_  = _w6494_ ;
	assign \g62807/_0_  = _w6496_ ;
	assign \g62811/_0_  = _w6498_ ;
	assign \g62968/_0_  = _w6501_ ;
	assign \g63005/_0_  = _w6504_ ;
	assign \g63041/_0_  = _w6506_ ;
	assign \g63116/_0_  = _w6510_ ;
	assign \g63157/_0_  = _w6514_ ;
	assign \g63164/_0_  = _w6516_ ;
	assign \g63170/_0_  = _w6520_ ;
	assign \g63189/_0_  = _w6522_ ;
	assign \g63202/_0_  = _w6525_ ;
	assign \g63206/_0_  = _w6527_ ;
	assign \g63207/_0_  = _w6538_ ;
	assign \g63265/_0_  = _w6541_ ;
	assign \g63266/_0_  = _w6544_ ;
	assign \g63269/_0_  = _w6547_ ;
	assign \g63271/_0_  = _w6550_ ;
	assign \g63272/_0_  = _w6553_ ;
	assign \g63273/_0_  = _w6556_ ;
	assign \g63274/_0_  = _w6559_ ;
	assign \g63275/_0_  = _w6562_ ;
	assign \g63276/_0_  = _w6565_ ;
	assign \g63277/_0_  = _w6568_ ;
	assign \g63278/_0_  = _w6571_ ;
	assign \g63280/_0_  = _w6574_ ;
	assign \g63281/_0_  = _w6577_ ;
	assign \g63282/_0_  = _w6580_ ;
	assign \g63283/_0_  = _w6583_ ;
	assign \g63284/_0_  = _w6586_ ;
	assign \g63285/_0_  = _w6589_ ;
	assign \g63286/_0_  = _w6592_ ;
	assign \g63287/_0_  = _w6595_ ;
	assign \g63288/_0_  = _w6598_ ;
	assign \g63289/_0_  = _w6601_ ;
	assign \g63290/_0_  = _w6604_ ;
	assign \g63292/_0_  = _w6607_ ;
	assign \g63293/_0_  = _w6610_ ;
	assign \g63294/_0_  = _w6613_ ;
	assign \g63295/_0_  = _w6616_ ;
	assign \g63296/_0_  = _w6619_ ;
	assign \g63297/_0_  = _w6622_ ;
	assign \g63298/_0_  = _w6625_ ;
	assign \g63299/_0_  = _w6628_ ;
	assign \g63302/_0_  = _w6631_ ;
	assign \g63303/_0_  = _w6634_ ;
	assign \g63304/_0_  = _w6637_ ;
	assign \g63305/_0_  = _w6640_ ;
	assign \g63306/_0_  = _w6643_ ;
	assign \g63307/_0_  = _w6646_ ;
	assign \g63308/_0_  = _w6649_ ;
	assign \g63309/_0_  = _w6652_ ;
	assign \g63310/_0_  = _w6655_ ;
	assign \g63311/_0_  = _w6658_ ;
	assign \g63312/_0_  = _w6661_ ;
	assign \g63313/_0_  = _w6664_ ;
	assign \g63314/_0_  = _w6667_ ;
	assign \g63315/_0_  = _w6670_ ;
	assign \g63316/_0_  = _w6673_ ;
	assign \g63317/_0_  = _w6676_ ;
	assign \g63318/_0_  = _w6679_ ;
	assign \g63319/_0_  = _w6682_ ;
	assign \g63320/_0_  = _w6685_ ;
	assign \g63321/_0_  = _w6688_ ;
	assign \g63322/_0_  = _w6691_ ;
	assign \g63323/_0_  = _w6694_ ;
	assign \g63324/_0_  = _w6697_ ;
	assign \g63325/_0_  = _w6700_ ;
	assign \g63326/_0_  = _w6703_ ;
	assign \g63327/_0_  = _w6706_ ;
	assign \g63328/_0_  = _w6709_ ;
	assign \g63329/_0_  = _w6712_ ;
	assign \g63330/_0_  = _w6715_ ;
	assign \g63331/_0_  = _w6718_ ;
	assign \g63339/_0_  = _w6721_ ;
	assign \g63505/_0_  = _w6724_ ;
	assign \g63525/_0_  = _w5264_ ;
	assign \g63543/_1_  = _w4465_ ;
	assign \g63602/_0_  = _w6727_ ;
	assign \g63653/_0_  = _w3320_ ;
	assign \g63663/_1_  = _w4473_ ;
	assign \g63677/_0_  = _w5343_ ;
	assign \g63694/_0_  = _w5399_ ;
	assign \g63729/_0_  = _w6730_ ;
	assign \g63766/_0_  = _w6733_ ;
	assign \g63771/_1_  = _w5023_ ;
	assign \g63773/_1_  = _w5029_ ;
	assign \g63784/_1_  = _w5027_ ;
	assign \g63964/_0_  = _w6758_ ;
	assign \g63965/_0_  = _w6782_ ;
	assign \g63966/_0_  = _w6785_ ;
	assign \g63967/_0_  = _w6788_ ;
	assign \g64257/_1_  = _w2551_ ;
	assign \g64266/_0_  = _w6791_ ;
	assign \g64275/_0_  = _w6794_ ;
	assign \g64400/_0_  = _w5036_ ;
	assign \g64416/_0_  = _w5309_ ;
	assign \g64470/_3_  = _w6799_ ;
	assign \g64473/_0_  = _w6804_ ;
	assign \g64474/_0_  = _w6809_ ;
	assign \g64475/_0_  = _w6814_ ;
	assign \g64479/_0_  = _w6826_ ;
	assign \g64480/_0_  = _w6830_ ;
	assign \g64481/_0_  = _w6834_ ;
	assign \g64483/_0_  = _w6839_ ;
	assign \g64484/_0_  = _w6844_ ;
	assign \g64485/_0_  = _w6847_ ;
	assign \g64486/_0_  = _w6850_ ;
	assign \g64493/_0_  = _w6855_ ;
	assign \g64494/_0_  = _w6860_ ;
	assign \g64495/_0_  = _w6865_ ;
	assign \g64496/_0_  = _w6870_ ;
	assign \g64505/_3_  = _w6873_ ;
	assign \g64507/_0_  = _w6878_ ;
	assign \g64508/_0_  = _w6883_ ;
	assign \g64510/_0_  = _w6888_ ;
	assign \g64511/_0_  = _w6893_ ;
	assign \g64544/_0_  = _w6896_ ;
	assign \g64545/_0_  = _w6899_ ;
	assign \g64546/_0_  = _w6902_ ;
	assign \g64639/_0_  = _w6905_ ;
	assign \g64641/_0_  = _w6908_ ;
	assign \g64642/_0_  = _w6911_ ;
	assign \g64645/_0_  = _w6914_ ;
	assign \g64650/_0_  = _w6917_ ;
	assign \g64737/_0_  = _w6920_ ;
	assign \g64738/_0_  = _w6923_ ;
	assign \g65066/_0_  = _w4993_ ;
	assign \g65070/_0_  = _w3754_ ;
	assign \g65090/_0_  = _w1826_ ;
	assign \g65102/_0_  = _w5076_ ;
	assign \g65102/_3_  = _w5076_ ;
	assign \g65126/_3_  = _w5478_ ;
	assign \g65147/_3_  = _w5514_ ;
	assign \g65163/_0_  = _w4849_ ;
	assign \g65176/_3_  = _w5553_ ;
	assign \g65178/_0_  = _w4370_ ;
	assign \g65182/_0_  = _w4835_ ;
	assign \g65190/_1_  = _w1745_ ;
	assign \g65191/_0_  = _w4268_ ;
	assign \g65196/_0_  = _w4224_ ;
	assign \g65268/_0_  = _w1643_ ;
	assign \g65275/_0_  = _w2929_ ;
	assign \g65290/_0_  = _w5138_ ;
	assign \g65290/_3_  = _w5138_ ;
	assign \g65291/_0_  = _w2938_ ;
	assign \g65292/_0_  = _w3673_ ;
	assign \g65298/_0_  = _w5107_ ;
	assign \g65298/_3_  = _w5107_ ;
	assign \g65314/_0_  = _w5169_ ;
	assign \g65314/_3_  = _w5169_ ;
	assign \g65319/_3_  = _w5589_ ;
	assign \g65335/_0_  = _w4947_ ;
	assign \g65342/_0_  = _w1633_ ;
	assign \g65348/_0_  = _w4416_ ;
	assign \g65422/_0_  = _w6926_ ;
	assign \g65465/_1_  = _w6827_ ;
	assign \g65469/_1_  = _w6831_ ;
	assign \g65478/_1_  = _w6821_ ;
	assign \g65507/_0_  = _w4136_ ;
	assign \g65548/_0_  = _w5085_ ;
	assign \g65699/_1_  = _w1223_ ;
	assign \g65713/_1_  = _w2610_ ;
	assign \g65835/_0_  = _w6927_ ;
	assign \g65860/_0_  = _w6820_ ;
	assign \g65863/_0_  = _w6928_ ;
	assign \g66094/_1_  = _w5116_ ;
	assign \g66102/_0_  = _w6931_ ;
	assign \g66107/_0_  = _w6934_ ;
	assign \g66130/_3_  = _w6937_ ;
	assign \g66131/_3_  = _w6940_ ;
	assign \g66228/_1_  = _w6099_ ;
	assign \g66348/_1_  = _w1466_ ;
	assign \g66543/_0_  = _w6942_ ;
	assign \g66549/_1_  = _w5178_ ;
	assign \g66640/_3_  = _w6945_ ;
	assign \g66641/_3_  = _w6948_ ;
	assign \g66950/_1_  = _w5045_ ;
	assign \g67111/_0_  = _w6949_ ;
	assign \g67219/_0_  = _w6950_ ;
	assign \g67263/_0_  = _w6952_ ;
	assign \g67909/_1_  = _w6102_ ;
	assign \g68049/_0_  = _w6954_ ;
	assign \g68220/_0_  = \g805_reg/NET0131 ;
	assign \g68413/_0_  = \g801_reg/NET0131 ;
	assign \g68511/_0_  = \g97_reg/NET0131 ;
	assign \g68536/_0_  = \g793_reg/NET0131 ;
	assign \g68543/_1_  = _w1462_ ;
	assign \g68554/_0_  = _w6955_ ;
	assign \g68559/_0_  = _w6956_ ;
	assign \g70915/_0_  = _w6963_ ;
	assign \g71108/_1_  = _w1537_ ;
	assign \g71115/_2_  = _w3665_ ;
	assign \g71244_dup/_0_  = _w2670_ ;
	assign \g71368/_0_  = _w6969_ ;
	assign \g71581/_0_  = _w6972_ ;
	assign \g71720/_0_  = _w1268_ ;
	assign \g785_reg/P0001  = \g785_reg/NET0131 ;
	assign \g789_reg/P0001  = \g789_reg/NET0131 ;
	assign \g797_reg/P0001  = \g797_reg/NET0131 ;
	assign \g809_reg/P0001  = \g809_reg/NET0131 ;
	assign \g813_reg/P0001  = \g813_reg/NET0131 ;
	assign \g966_reg/P0001  = \g966_reg/NET0131 ;
	assign \g968_reg/P0001  = \g968_reg/NET0131 ;
	assign \g970_reg/P0001  = \g970_reg/NET0131 ;
	assign \g972_reg/P0001  = \g972_reg/NET0131 ;
	assign \g974_reg/P0001  = \g974_reg/NET0131 ;
	assign \g976_reg/P0001  = \g976_reg/NET0131 ;
	assign \g978_reg/P0001  = \g978_reg/NET0131 ;
endmodule;