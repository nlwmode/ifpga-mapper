module top( \line1_pad  , \line2_pad  , \stato_reg[0]/NET0131  , \stato_reg[1]/NET0131  , \stato_reg[2]/NET0131  , \_al_n0  , \_al_n1  , \g220/_2_  , \g221/_0_  , \g222/_0_  , \g224/_0_  , \g44/_1_  );
  input \line1_pad  ;
  input \line2_pad  ;
  input \stato_reg[0]/NET0131  ;
  input \stato_reg[1]/NET0131  ;
  input \stato_reg[2]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g220/_2_  ;
  output \g221/_0_  ;
  output \g222/_0_  ;
  output \g224/_0_  ;
  output \g44/_1_  ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n6 = ~\stato_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n7 = ~\stato_reg[2]/NET0131  & ~n6 ;
  assign n8 = \stato_reg[0]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n9 = \stato_reg[2]/NET0131  & ~n8 ;
  assign n10 = ~n7 & ~n9 ;
  assign n11 = \line1_pad  & \line2_pad  ;
  assign n12 = ~\stato_reg[0]/NET0131  & ~n11 ;
  assign n13 = ~\line1_pad  & ~\line2_pad  ;
  assign n14 = \stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n15 = ~n13 & n14 ;
  assign n16 = ~n12 & n15 ;
  assign n17 = ~n10 & ~n16 ;
  assign n18 = ~\stato_reg[2]/NET0131  & n8 ;
  assign n19 = ~n11 & n18 ;
  assign n20 = ~\stato_reg[0]/NET0131  & n13 ;
  assign n21 = ~\stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n22 = n20 & n21 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = n17 & n23 ;
  assign n25 = ~n6 & ~n18 ;
  assign n26 = n11 & ~n25 ;
  assign n27 = \stato_reg[2]/NET0131  & ~n6 ;
  assign n28 = ~n13 & n27 ;
  assign n29 = ~n8 & ~n11 ;
  assign n30 = n7 & n29 ;
  assign n31 = ~n28 & ~n30 ;
  assign n32 = ~n26 & n31 ;
  assign n33 = ~n11 & ~n13 ;
  assign n34 = ~n27 & n33 ;
  assign n35 = n27 & ~n33 ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = n7 & ~n11 ;
  assign n38 = ~\stato_reg[0]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n39 = n13 & n38 ;
  assign n40 = ~n14 & ~n39 ;
  assign n41 = ~n37 & n40 ;
  assign n42 = \stato_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n43 = ~\stato_reg[2]/NET0131  & n42 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g220/_2_  = ~n24 ;
  assign \g221/_0_  = ~n32 ;
  assign \g222/_0_  = ~n36 ;
  assign \g224/_0_  = n41 ;
  assign \g44/_1_  = n43 ;
endmodule
