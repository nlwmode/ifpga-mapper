module top (\g108_reg/NET0131 , \g109_pad , \g1212_reg/NET0131 , \g1218_reg/NET0131 , \g1223_reg/NET0131 , \g1227_reg/NET0131 , \g1231_reg/NET0131 , \g1235_reg/NET0131 , \g1240_reg/NET0131 , \g1245_reg/NET0131 , \g1250_reg/NET0131 , \g1255_reg/NET0131 , \g1260_reg/NET0131 , \g1265_reg/NET0131 , \g1270_reg/NET0131 , \g1275_reg/NET0131 , \g1280_reg/NET0131 , \g1284_reg/NET0131 , \g1289_reg/NET0131 , \g1292_reg/NET0131 , \g1296_reg/NET0131 , \g1300_reg/NET0131 , \g1304_reg/NET0131 , \g1336_reg/NET0131 , \g1341_reg/NET0131 , \g1346_reg/NET0131 , \g1351_reg/NET0131 , \g1361_reg/NET0131 , \g1362_reg/NET0131 , \g1365_reg/NET0131 , \g1368_reg/NET0131 , \g1371_reg/NET0131 , \g1374_reg/NET0131 , \g1377_reg/NET0131 , \g1380_reg/NET0131 , \g1383_reg/NET0131 , \g1386_reg/NET0131 , \g1389_reg/NET0131 , \g1397_reg/NET0131 , \g1400_reg/NET0131 , \g1615_reg/NET0131 , \g1618_reg/NET0131 , \g1621_reg/NET0131 , \g1624_reg/NET0131 , \g1627_reg/NET0131 , \g1630_reg/NET0131 , \g1633_reg/NET0131 , \g1636_reg/NET0131 , \g1718_reg/NET0131 , \g186_reg/NET0131 , \g192_reg/NET0131 , \g197_reg/NET0131 , \g201_reg/NET0131 , \g207_reg/NET0131 , \g213_reg/NET0131 , \g219_reg/NET0131 , \g225_reg/NET0131 , \g231_reg/NET0131 , \g2355_pad , \g237_reg/NET0131 , \g243_reg/NET0131 , \g248_reg/NET0131 , \g3007_pad , \g305_reg/NET0131 , \g3069_pad , \g309_reg/NET0131 , \g312_reg/NET0131 , \g315_reg/NET0131 , \g318_reg/NET0131 , \g321_reg/NET0131 , \g324_reg/NET0131 , \g327_reg/NET0131 , \g330_reg/NET0131 , \g333_reg/NET0131 , \g369_reg/NET0131 , \g374_reg/NET0131 , \g378_reg/NET0131 , \g382_reg/NET0131 , \g386_reg/NET0131 , \g391_reg/NET0131 , \g396_reg/NET0131 , \g401_reg/NET0131 , \g406_reg/NET0131 , \g411_reg/NET0131 , \g416_reg/NET0131 , \g4173_pad , \g4174_pad , \g4175_pad , \g4176_pad , \g4177_pad , \g4178_pad , \g4179_pad , \g4180_pad , \g4181_pad , \g421_reg/NET0131 , \g426_reg/NET0131 , \g431_reg/NET0131 , \g435_reg/NET0131 , \g440_reg/NET0131 , \g444_reg/NET0131 , \g448_reg/NET0131 , \g452_reg/NET0131 , \g546_reg/NET0131 , \g549_reg/NET0131 , \g554_reg/NET0131 , \g557_reg/NET0131 , \g560_reg/NET0131 , \g563_reg/NET0131 , \g566_reg/NET0131 , \g569_reg/NET0131 , \g572_reg/NET0131 , \g575_reg/NET0131 , \g741_pad , \g742_pad , \g743_pad , \g744_pad , \g757_reg/NET0131 , \g876_reg/NET0131 , \g971_reg/NET0131 , \g976_reg/NET0131 , \g981_reg/NET0131 , \g986_reg/NET0131 , \g21280/_0_ , \g21281/_0_ , \g21282/_0_ , \g21307/_0_ , \g21322/_0_ , \g21333/_0_ , \g21334/_0_ , \g21338/_0_ , \g21350/_0_ , \g21355/_0_ , \g21356/_0_ , \g21357/_0_ , \g21358/_1_ , \g21359/_0_ , \g21370/_0_ , \g21371/_0_ , \g21378/_0_ , \g21379/_0_ , \g21380/_1_ , \g21381/_0_ , \g21390/_0_ , \g21394/_0_ , \g21396/_0_ , \g21397/_0_ , \g21398/_1_ , \g21412/_0_ , \g21413/_0_ , \g21419/_0_ , \g21420/_00_ , \g21421/_00_ , \g21424/_0_ , \g21425/_0_ , \g21426/_1_ , \g21437/_0_ , \g21444/_0_ , \g21450/_0_ , \g21455/_0_ , \g21457/_0_ , \g21458/_1_ , \g21459/_0_ , \g21470/_0_ , \g21486/_0_ , \g21487/_0_ , \g21495/_0_ , \g21498/_1_ , \g21499/_0_ , \g21500/_0_ , \g21502/_0_ , \g21503/_0_ , \g21508/_0_ , \g21509/_0_ , \g21510/_0_ , \g21511/_0_ , \g21515/_0_ , \g21520/_0_ , \g21523/_0_ , \g21524/_0_ , \g21525/_0_ , \g21538/_0_ , \g21544/_0_ , \g21550/_1_ , \g21562/_0_ , \g21563/_0_ , \g21584/_0_ , \g21591/_0_ , \g21593/_0_ , \g21601/_3_ , \g21603/_3_ , \g21605/_3_ , \g21607/_3_ , \g21609/_3_ , \g21611/_3_ , \g21613/_3_ , \g21615/_3_ , \g21617/_3_ , \g21619/_3_ , \g21621/_3_ , \g21623/_3_ , \g21625/_3_ , \g21627/_3_ , \g21640/_0_ , \g21641/_0_ , \g21642/_0_ , \g21693/_0_ , \g21694/_0_ , \g21735/_2_ , \g21745/_2_ , \g21796/_0_ , \g21799/_0_ , \g21803/_0_ , \g21812/_0_ , \g21814/_0_ , \g21816/_0_ , \g21828/_0_ , \g22203/_0_ , \g22260/_1_ , \g22317/_0_ , \g22339/_0_ , \g22392/_0_ , \g22395/_1_ , \g2601_pad , \g27_dup/_0_ , \g5816_pad );
	input \g108_reg/NET0131  ;
	input \g109_pad  ;
	input \g1212_reg/NET0131  ;
	input \g1218_reg/NET0131  ;
	input \g1223_reg/NET0131  ;
	input \g1227_reg/NET0131  ;
	input \g1231_reg/NET0131  ;
	input \g1235_reg/NET0131  ;
	input \g1240_reg/NET0131  ;
	input \g1245_reg/NET0131  ;
	input \g1250_reg/NET0131  ;
	input \g1255_reg/NET0131  ;
	input \g1260_reg/NET0131  ;
	input \g1265_reg/NET0131  ;
	input \g1270_reg/NET0131  ;
	input \g1275_reg/NET0131  ;
	input \g1280_reg/NET0131  ;
	input \g1284_reg/NET0131  ;
	input \g1289_reg/NET0131  ;
	input \g1292_reg/NET0131  ;
	input \g1296_reg/NET0131  ;
	input \g1300_reg/NET0131  ;
	input \g1304_reg/NET0131  ;
	input \g1336_reg/NET0131  ;
	input \g1341_reg/NET0131  ;
	input \g1346_reg/NET0131  ;
	input \g1351_reg/NET0131  ;
	input \g1361_reg/NET0131  ;
	input \g1362_reg/NET0131  ;
	input \g1365_reg/NET0131  ;
	input \g1368_reg/NET0131  ;
	input \g1371_reg/NET0131  ;
	input \g1374_reg/NET0131  ;
	input \g1377_reg/NET0131  ;
	input \g1380_reg/NET0131  ;
	input \g1383_reg/NET0131  ;
	input \g1386_reg/NET0131  ;
	input \g1389_reg/NET0131  ;
	input \g1397_reg/NET0131  ;
	input \g1400_reg/NET0131  ;
	input \g1615_reg/NET0131  ;
	input \g1618_reg/NET0131  ;
	input \g1621_reg/NET0131  ;
	input \g1624_reg/NET0131  ;
	input \g1627_reg/NET0131  ;
	input \g1630_reg/NET0131  ;
	input \g1633_reg/NET0131  ;
	input \g1636_reg/NET0131  ;
	input \g1718_reg/NET0131  ;
	input \g186_reg/NET0131  ;
	input \g192_reg/NET0131  ;
	input \g197_reg/NET0131  ;
	input \g201_reg/NET0131  ;
	input \g207_reg/NET0131  ;
	input \g213_reg/NET0131  ;
	input \g219_reg/NET0131  ;
	input \g225_reg/NET0131  ;
	input \g231_reg/NET0131  ;
	input \g2355_pad  ;
	input \g237_reg/NET0131  ;
	input \g243_reg/NET0131  ;
	input \g248_reg/NET0131  ;
	input \g3007_pad  ;
	input \g305_reg/NET0131  ;
	input \g3069_pad  ;
	input \g309_reg/NET0131  ;
	input \g312_reg/NET0131  ;
	input \g315_reg/NET0131  ;
	input \g318_reg/NET0131  ;
	input \g321_reg/NET0131  ;
	input \g324_reg/NET0131  ;
	input \g327_reg/NET0131  ;
	input \g330_reg/NET0131  ;
	input \g333_reg/NET0131  ;
	input \g369_reg/NET0131  ;
	input \g374_reg/NET0131  ;
	input \g378_reg/NET0131  ;
	input \g382_reg/NET0131  ;
	input \g386_reg/NET0131  ;
	input \g391_reg/NET0131  ;
	input \g396_reg/NET0131  ;
	input \g401_reg/NET0131  ;
	input \g406_reg/NET0131  ;
	input \g411_reg/NET0131  ;
	input \g416_reg/NET0131  ;
	input \g4173_pad  ;
	input \g4174_pad  ;
	input \g4175_pad  ;
	input \g4176_pad  ;
	input \g4177_pad  ;
	input \g4178_pad  ;
	input \g4179_pad  ;
	input \g4180_pad  ;
	input \g4181_pad  ;
	input \g421_reg/NET0131  ;
	input \g426_reg/NET0131  ;
	input \g431_reg/NET0131  ;
	input \g435_reg/NET0131  ;
	input \g440_reg/NET0131  ;
	input \g444_reg/NET0131  ;
	input \g448_reg/NET0131  ;
	input \g452_reg/NET0131  ;
	input \g546_reg/NET0131  ;
	input \g549_reg/NET0131  ;
	input \g554_reg/NET0131  ;
	input \g557_reg/NET0131  ;
	input \g560_reg/NET0131  ;
	input \g563_reg/NET0131  ;
	input \g566_reg/NET0131  ;
	input \g569_reg/NET0131  ;
	input \g572_reg/NET0131  ;
	input \g575_reg/NET0131  ;
	input \g741_pad  ;
	input \g742_pad  ;
	input \g743_pad  ;
	input \g744_pad  ;
	input \g757_reg/NET0131  ;
	input \g876_reg/NET0131  ;
	input \g971_reg/NET0131  ;
	input \g976_reg/NET0131  ;
	input \g981_reg/NET0131  ;
	input \g986_reg/NET0131  ;
	output \g21280/_0_  ;
	output \g21281/_0_  ;
	output \g21282/_0_  ;
	output \g21307/_0_  ;
	output \g21322/_0_  ;
	output \g21333/_0_  ;
	output \g21334/_0_  ;
	output \g21338/_0_  ;
	output \g21350/_0_  ;
	output \g21355/_0_  ;
	output \g21356/_0_  ;
	output \g21357/_0_  ;
	output \g21358/_1_  ;
	output \g21359/_0_  ;
	output \g21370/_0_  ;
	output \g21371/_0_  ;
	output \g21378/_0_  ;
	output \g21379/_0_  ;
	output \g21380/_1_  ;
	output \g21381/_0_  ;
	output \g21390/_0_  ;
	output \g21394/_0_  ;
	output \g21396/_0_  ;
	output \g21397/_0_  ;
	output \g21398/_1_  ;
	output \g21412/_0_  ;
	output \g21413/_0_  ;
	output \g21419/_0_  ;
	output \g21420/_00_  ;
	output \g21421/_00_  ;
	output \g21424/_0_  ;
	output \g21425/_0_  ;
	output \g21426/_1_  ;
	output \g21437/_0_  ;
	output \g21444/_0_  ;
	output \g21450/_0_  ;
	output \g21455/_0_  ;
	output \g21457/_0_  ;
	output \g21458/_1_  ;
	output \g21459/_0_  ;
	output \g21470/_0_  ;
	output \g21486/_0_  ;
	output \g21487/_0_  ;
	output \g21495/_0_  ;
	output \g21498/_1_  ;
	output \g21499/_0_  ;
	output \g21500/_0_  ;
	output \g21502/_0_  ;
	output \g21503/_0_  ;
	output \g21508/_0_  ;
	output \g21509/_0_  ;
	output \g21510/_0_  ;
	output \g21511/_0_  ;
	output \g21515/_0_  ;
	output \g21520/_0_  ;
	output \g21523/_0_  ;
	output \g21524/_0_  ;
	output \g21525/_0_  ;
	output \g21538/_0_  ;
	output \g21544/_0_  ;
	output \g21550/_1_  ;
	output \g21562/_0_  ;
	output \g21563/_0_  ;
	output \g21584/_0_  ;
	output \g21591/_0_  ;
	output \g21593/_0_  ;
	output \g21601/_3_  ;
	output \g21603/_3_  ;
	output \g21605/_3_  ;
	output \g21607/_3_  ;
	output \g21609/_3_  ;
	output \g21611/_3_  ;
	output \g21613/_3_  ;
	output \g21615/_3_  ;
	output \g21617/_3_  ;
	output \g21619/_3_  ;
	output \g21621/_3_  ;
	output \g21623/_3_  ;
	output \g21625/_3_  ;
	output \g21627/_3_  ;
	output \g21640/_0_  ;
	output \g21641/_0_  ;
	output \g21642/_0_  ;
	output \g21693/_0_  ;
	output \g21694/_0_  ;
	output \g21735/_2_  ;
	output \g21745/_2_  ;
	output \g21796/_0_  ;
	output \g21799/_0_  ;
	output \g21803/_0_  ;
	output \g21812/_0_  ;
	output \g21814/_0_  ;
	output \g21816/_0_  ;
	output \g21828/_0_  ;
	output \g22203/_0_  ;
	output \g22260/_1_  ;
	output \g22317/_0_  ;
	output \g22339/_0_  ;
	output \g22392/_0_  ;
	output \g22395/_1_  ;
	output \g2601_pad  ;
	output \g27_dup/_0_  ;
	output \g5816_pad  ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	LUT4 #(
		.INIT('h8000)
	) name0 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		\g378_reg/NET0131 ,
		\g382_reg/NET0131 ,
		_w124_
	);
	LUT4 #(
		.INIT('h0001)
	) name1 (
		\g396_reg/NET0131 ,
		\g401_reg/NET0131 ,
		\g406_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w125_
	);
	LUT4 #(
		.INIT('h0001)
	) name2 (
		\g386_reg/NET0131 ,
		\g391_reg/NET0131 ,
		\g431_reg/NET0131 ,
		\g435_reg/NET0131 ,
		_w126_
	);
	LUT3 #(
		.INIT('h01)
	) name3 (
		\g444_reg/NET0131 ,
		\g448_reg/NET0131 ,
		\g452_reg/NET0131 ,
		_w127_
	);
	LUT4 #(
		.INIT('h0001)
	) name4 (
		\g416_reg/NET0131 ,
		\g421_reg/NET0131 ,
		\g426_reg/NET0131 ,
		\g440_reg/NET0131 ,
		_w128_
	);
	LUT4 #(
		.INIT('h8000)
	) name5 (
		_w127_,
		_w128_,
		_w125_,
		_w126_,
		_w129_
	);
	LUT2 #(
		.INIT('h6)
	) name6 (
		\g431_reg/NET0131 ,
		\g435_reg/NET0131 ,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h6)
	) name8 (
		\g315_reg/NET0131 ,
		\g426_reg/NET0131 ,
		_w132_
	);
	LUT4 #(
		.INIT('h8241)
	) name9 (
		\g312_reg/NET0131 ,
		\g324_reg/NET0131 ,
		\g396_reg/NET0131 ,
		\g421_reg/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name11 (
		\g318_reg/NET0131 ,
		\g330_reg/NET0131 ,
		\g386_reg/NET0131 ,
		\g406_reg/NET0131 ,
		_w135_
	);
	LUT4 #(
		.INIT('haf23)
	) name12 (
		\g318_reg/NET0131 ,
		\g321_reg/NET0131 ,
		\g386_reg/NET0131 ,
		\g391_reg/NET0131 ,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w135_,
		_w136_,
		_w137_
	);
	LUT4 #(
		.INIT('h8caf)
	) name14 (
		\g321_reg/NET0131 ,
		\g333_reg/NET0131 ,
		\g391_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w138_
	);
	LUT4 #(
		.INIT('hf351)
	) name15 (
		\g309_reg/NET0131 ,
		\g330_reg/NET0131 ,
		\g406_reg/NET0131 ,
		\g416_reg/NET0131 ,
		_w139_
	);
	LUT2 #(
		.INIT('h6)
	) name16 (
		\g327_reg/NET0131 ,
		\g401_reg/NET0131 ,
		_w140_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name17 (
		\g309_reg/NET0131 ,
		\g333_reg/NET0131 ,
		\g411_reg/NET0131 ,
		\g416_reg/NET0131 ,
		_w141_
	);
	LUT4 #(
		.INIT('h4000)
	) name18 (
		_w140_,
		_w141_,
		_w138_,
		_w139_,
		_w142_
	);
	LUT3 #(
		.INIT('h80)
	) name19 (
		_w137_,
		_w134_,
		_w142_,
		_w143_
	);
	LUT4 #(
		.INIT('h84cc)
	) name20 (
		\g305_reg/NET0131 ,
		_w124_,
		_w131_,
		_w143_,
		_w144_
	);
	LUT4 #(
		.INIT('h0a02)
	) name21 (
		\g1212_reg/NET0131 ,
		\g3007_pad ,
		\g757_reg/NET0131 ,
		\g876_reg/NET0131 ,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\g109_pad ,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\g971_reg/NET0131 ,
		\g976_reg/NET0131 ,
		_w147_
	);
	LUT4 #(
		.INIT('h6c00)
	) name24 (
		\g971_reg/NET0131 ,
		\g976_reg/NET0131 ,
		_w144_,
		_w146_,
		_w148_
	);
	LUT3 #(
		.INIT('h80)
	) name25 (
		\g971_reg/NET0131 ,
		\g976_reg/NET0131 ,
		\g981_reg/NET0131 ,
		_w149_
	);
	LUT4 #(
		.INIT('h60a0)
	) name26 (
		\g981_reg/NET0131 ,
		_w144_,
		_w146_,
		_w147_,
		_w150_
	);
	LUT4 #(
		.INIT('h8000)
	) name27 (
		\g971_reg/NET0131 ,
		\g976_reg/NET0131 ,
		\g981_reg/NET0131 ,
		\g986_reg/NET0131 ,
		_w151_
	);
	LUT4 #(
		.INIT('h60a0)
	) name28 (
		\g986_reg/NET0131 ,
		_w144_,
		_w146_,
		_w149_,
		_w152_
	);
	LUT4 #(
		.INIT('h0001)
	) name29 (
		\g1362_reg/NET0131 ,
		\g1365_reg/NET0131 ,
		\g1368_reg/NET0131 ,
		\g1371_reg/NET0131 ,
		_w153_
	);
	LUT4 #(
		.INIT('h0001)
	) name30 (
		\g1386_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		\g197_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT4 #(
		.INIT('h0001)
	) name32 (
		\g1397_reg/NET0131 ,
		\g1400_reg/NET0131 ,
		\g186_reg/NET0131 ,
		\g192_reg/NET0131 ,
		_w156_
	);
	LUT4 #(
		.INIT('h0001)
	) name33 (
		\g1374_reg/NET0131 ,
		\g1377_reg/NET0131 ,
		\g1380_reg/NET0131 ,
		\g1383_reg/NET0131 ,
		_w157_
	);
	LUT4 #(
		.INIT('h0001)
	) name34 (
		\g231_reg/NET0131 ,
		\g237_reg/NET0131 ,
		\g243_reg/NET0131 ,
		\g248_reg/NET0131 ,
		_w158_
	);
	LUT4 #(
		.INIT('h0001)
	) name35 (
		\g207_reg/NET0131 ,
		\g213_reg/NET0131 ,
		\g219_reg/NET0131 ,
		\g225_reg/NET0131 ,
		_w159_
	);
	LUT4 #(
		.INIT('h8000)
	) name36 (
		_w158_,
		_w159_,
		_w156_,
		_w157_,
		_w160_
	);
	LUT4 #(
		.INIT('h9009)
	) name37 (
		\g1386_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		\g197_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w161_
	);
	LUT4 #(
		.INIT('h0660)
	) name38 (
		\g1386_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		\g197_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\g109_pad ,
		_w162_,
		_w163_
	);
	LUT4 #(
		.INIT('h8f00)
	) name40 (
		_w155_,
		_w160_,
		_w161_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\g213_reg/NET0131 ,
		\g2355_pad ,
		_w165_
	);
	LUT3 #(
		.INIT('hb8)
	) name42 (
		\g213_reg/NET0131 ,
		\g2355_pad ,
		\g557_reg/NET0131 ,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\g186_reg/NET0131 ,
		\g2355_pad ,
		_w167_
	);
	LUT3 #(
		.INIT('hb8)
	) name44 (
		\g186_reg/NET0131 ,
		\g2355_pad ,
		\g546_reg/NET0131 ,
		_w168_
	);
	LUT4 #(
		.INIT('h3022)
	) name45 (
		\g1615_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g213_reg/NET0131 ,
		\g2355_pad ,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\g219_reg/NET0131 ,
		\g2355_pad ,
		_w170_
	);
	LUT3 #(
		.INIT('hb8)
	) name47 (
		\g219_reg/NET0131 ,
		\g2355_pad ,
		\g560_reg/NET0131 ,
		_w171_
	);
	LUT4 #(
		.INIT('h3022)
	) name48 (
		\g1618_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g186_reg/NET0131 ,
		\g2355_pad ,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\g207_reg/NET0131 ,
		\g2355_pad ,
		_w173_
	);
	LUT3 #(
		.INIT('hb8)
	) name50 (
		\g207_reg/NET0131 ,
		\g2355_pad ,
		\g554_reg/NET0131 ,
		_w174_
	);
	LUT4 #(
		.INIT('h3022)
	) name51 (
		\g1621_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g219_reg/NET0131 ,
		\g2355_pad ,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\g109_pad ,
		\g186_reg/NET0131 ,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\g225_reg/NET0131 ,
		\g2355_pad ,
		_w177_
	);
	LUT3 #(
		.INIT('hb8)
	) name54 (
		\g225_reg/NET0131 ,
		\g2355_pad ,
		\g563_reg/NET0131 ,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\g109_pad ,
		\g1383_reg/NET0131 ,
		_w179_
	);
	LUT3 #(
		.INIT('hea)
	) name56 (
		\g1718_reg/NET0131 ,
		\g207_reg/NET0131 ,
		\g2355_pad ,
		_w180_
	);
	LUT4 #(
		.INIT('h3022)
	) name57 (
		\g1624_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g225_reg/NET0131 ,
		\g2355_pad ,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\g109_pad ,
		\g207_reg/NET0131 ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\g231_reg/NET0131 ,
		\g2355_pad ,
		_w183_
	);
	LUT3 #(
		.INIT('hb8)
	) name60 (
		\g231_reg/NET0131 ,
		\g2355_pad ,
		\g566_reg/NET0131 ,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\g109_pad ,
		\g1380_reg/NET0131 ,
		_w185_
	);
	LUT4 #(
		.INIT('h3022)
	) name62 (
		\g1627_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g231_reg/NET0131 ,
		\g2355_pad ,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\g2355_pad ,
		\g237_reg/NET0131 ,
		_w187_
	);
	LUT3 #(
		.INIT('hd8)
	) name64 (
		\g2355_pad ,
		\g237_reg/NET0131 ,
		\g569_reg/NET0131 ,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\g109_pad ,
		\g213_reg/NET0131 ,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\g4173_pad ,
		\g4174_pad ,
		_w190_
	);
	LUT3 #(
		.INIT('h80)
	) name67 (
		\g4173_pad ,
		\g4174_pad ,
		\g4175_pad ,
		_w191_
	);
	LUT4 #(
		.INIT('h8000)
	) name68 (
		\g4173_pad ,
		\g4174_pad ,
		\g4175_pad ,
		\g4176_pad ,
		_w192_
	);
	LUT3 #(
		.INIT('h80)
	) name69 (
		\g4177_pad ,
		\g4178_pad ,
		_w192_,
		_w193_
	);
	LUT4 #(
		.INIT('h8000)
	) name70 (
		\g4177_pad ,
		\g4178_pad ,
		\g4179_pad ,
		_w192_,
		_w194_
	);
	LUT4 #(
		.INIT('h1555)
	) name71 (
		\g1718_reg/NET0131 ,
		\g4180_pad ,
		\g4181_pad ,
		_w194_,
		_w195_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name72 (
		\g109_pad ,
		\g4180_pad ,
		\g4181_pad ,
		_w194_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\g109_pad ,
		\g1377_reg/NET0131 ,
		_w198_
	);
	LUT4 #(
		.INIT('h3202)
	) name75 (
		\g1630_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g2355_pad ,
		\g237_reg/NET0131 ,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\g1240_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		_w200_
	);
	LUT3 #(
		.INIT('h01)
	) name77 (
		\g1255_reg/NET0131 ,
		\g1260_reg/NET0131 ,
		\g1270_reg/NET0131 ,
		_w201_
	);
	LUT4 #(
		.INIT('h0001)
	) name78 (
		\g1235_reg/NET0131 ,
		\g1250_reg/NET0131 ,
		\g1265_reg/NET0131 ,
		\g1275_reg/NET0131 ,
		_w202_
	);
	LUT4 #(
		.INIT('h0001)
	) name79 (
		\g1292_reg/NET0131 ,
		\g1296_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w203_
	);
	LUT4 #(
		.INIT('h8000)
	) name80 (
		_w202_,
		_w200_,
		_w201_,
		_w203_,
		_w204_
	);
	LUT3 #(
		.INIT('h80)
	) name81 (
		_w202_,
		_w200_,
		_w201_,
		_w205_
	);
	LUT4 #(
		.INIT('h8900)
	) name82 (
		\g1280_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w207_
	);
	LUT3 #(
		.INIT('h80)
	) name84 (
		\g1218_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		\g1227_reg/NET0131 ,
		_w208_
	);
	LUT3 #(
		.INIT('h80)
	) name85 (
		\g1231_reg/NET0131 ,
		_w207_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w206_,
		_w209_,
		_w210_
	);
	LUT4 #(
		.INIT('h4044)
	) name87 (
		\g108_reg/NET0131 ,
		\g1212_reg/NET0131 ,
		\g1361_reg/NET0131 ,
		\g3069_pad ,
		_w211_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\g109_pad ,
		_w211_,
		_w212_
	);
	LUT4 #(
		.INIT('h8a00)
	) name89 (
		\g1346_reg/NET0131 ,
		_w206_,
		_w209_,
		_w212_,
		_w213_
	);
	LUT3 #(
		.INIT('h78)
	) name90 (
		\g1336_reg/NET0131 ,
		\g1341_reg/NET0131 ,
		\g1346_reg/NET0131 ,
		_w214_
	);
	LUT4 #(
		.INIT('h4000)
	) name91 (
		_w206_,
		_w209_,
		_w212_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('he)
	) name92 (
		_w213_,
		_w215_,
		_w216_
	);
	LUT4 #(
		.INIT('h8a00)
	) name93 (
		\g1351_reg/NET0131 ,
		_w206_,
		_w209_,
		_w212_,
		_w217_
	);
	LUT4 #(
		.INIT('h8000)
	) name94 (
		\g1336_reg/NET0131 ,
		\g1341_reg/NET0131 ,
		\g1346_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w218_
	);
	LUT4 #(
		.INIT('h7f80)
	) name95 (
		\g1336_reg/NET0131 ,
		\g1341_reg/NET0131 ,
		\g1346_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w219_
	);
	LUT4 #(
		.INIT('h4000)
	) name96 (
		_w206_,
		_w209_,
		_w212_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('he)
	) name97 (
		_w217_,
		_w220_,
		_w221_
	);
	LUT3 #(
		.INIT('hd8)
	) name98 (
		\g2355_pad ,
		\g243_reg/NET0131 ,
		\g572_reg/NET0131 ,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\g109_pad ,
		\g219_reg/NET0131 ,
		_w223_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\g109_pad ,
		\g1718_reg/NET0131 ,
		_w224_
	);
	LUT3 #(
		.INIT('h60)
	) name101 (
		\g4180_pad ,
		_w194_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\g109_pad ,
		\g1371_reg/NET0131 ,
		_w226_
	);
	LUT4 #(
		.INIT('hfece)
	) name103 (
		\g1633_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g2355_pad ,
		\g243_reg/NET0131 ,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\g109_pad ,
		\g225_reg/NET0131 ,
		_w228_
	);
	LUT3 #(
		.INIT('h60)
	) name105 (
		\g4179_pad ,
		_w193_,
		_w224_,
		_w229_
	);
	LUT3 #(
		.INIT('hd8)
	) name106 (
		\g2355_pad ,
		\g248_reg/NET0131 ,
		\g575_reg/NET0131 ,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\g109_pad ,
		\g1368_reg/NET0131 ,
		_w231_
	);
	LUT4 #(
		.INIT('hfece)
	) name108 (
		\g1636_reg/NET0131 ,
		\g1718_reg/NET0131 ,
		\g2355_pad ,
		\g248_reg/NET0131 ,
		_w232_
	);
	LUT4 #(
		.INIT('h6c00)
	) name109 (
		\g4177_pad ,
		\g4178_pad ,
		_w192_,
		_w224_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\g109_pad ,
		\g231_reg/NET0131 ,
		_w234_
	);
	LUT4 #(
		.INIT('h8000)
	) name111 (
		\g1218_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		\g1227_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		_w236_
	);
	LUT3 #(
		.INIT('h08)
	) name113 (
		\g1218_reg/NET0131 ,
		_w207_,
		_w235_,
		_w237_
	);
	LUT4 #(
		.INIT('ha060)
	) name114 (
		\g1218_reg/NET0131 ,
		_w207_,
		_w236_,
		_w235_,
		_w238_
	);
	LUT3 #(
		.INIT('h48)
	) name115 (
		\g1223_reg/NET0131 ,
		_w236_,
		_w237_,
		_w239_
	);
	LUT4 #(
		.INIT('h2a80)
	) name116 (
		\g109_pad ,
		\g1218_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		\g1227_reg/NET0131 ,
		_w240_
	);
	LUT3 #(
		.INIT('h20)
	) name117 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1227_reg/NET0131 ,
		_w241_
	);
	LUT4 #(
		.INIT('hfd20)
	) name118 (
		_w207_,
		_w235_,
		_w240_,
		_w241_,
		_w242_
	);
	LUT4 #(
		.INIT('hea00)
	) name119 (
		\g1231_reg/NET0131 ,
		_w207_,
		_w208_,
		_w236_,
		_w243_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name120 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		\g378_reg/NET0131 ,
		\g382_reg/NET0131 ,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		_w236_,
		_w244_,
		_w245_
	);
	LUT4 #(
		.INIT('h1999)
	) name122 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		\g378_reg/NET0131 ,
		\g382_reg/NET0131 ,
		_w246_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		_w236_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h0080)
	) name124 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		\g378_reg/NET0131 ,
		\g382_reg/NET0131 ,
		_w248_
	);
	LUT3 #(
		.INIT('h07)
	) name125 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		\g378_reg/NET0131 ,
		_w249_
	);
	LUT3 #(
		.INIT('h02)
	) name126 (
		_w236_,
		_w248_,
		_w249_,
		_w250_
	);
	LUT4 #(
		.INIT('h007f)
	) name127 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		\g378_reg/NET0131 ,
		\g382_reg/NET0131 ,
		_w251_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		_w236_,
		_w251_,
		_w252_
	);
	LUT4 #(
		.INIT('h80a0)
	) name129 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1275_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w253_
	);
	LUT4 #(
		.INIT('h7600)
	) name130 (
		\g1280_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		_w204_,
		_w209_,
		_w254_
	);
	LUT2 #(
		.INIT('he)
	) name131 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT3 #(
		.INIT('h60)
	) name132 (
		\g4177_pad ,
		_w192_,
		_w224_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\g109_pad ,
		\g1365_reg/NET0131 ,
		_w257_
	);
	LUT3 #(
		.INIT('hb8)
	) name134 (
		\g192_reg/NET0131 ,
		\g2355_pad ,
		\g549_reg/NET0131 ,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		\g201_reg/NET0131 ,
		\g2355_pad ,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\g109_pad ,
		\g237_reg/NET0131 ,
		_w260_
	);
	LUT3 #(
		.INIT('h60)
	) name137 (
		\g4176_pad ,
		_w191_,
		_w224_,
		_w261_
	);
	LUT3 #(
		.INIT('hea)
	) name138 (
		\g1718_reg/NET0131 ,
		\g192_reg/NET0131 ,
		\g2355_pad ,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\g109_pad ,
		\g1362_reg/NET0131 ,
		_w263_
	);
	LUT4 #(
		.INIT('h0220)
	) name140 (
		\g109_pad ,
		\g1718_reg/NET0131 ,
		\g4173_pad ,
		\g4174_pad ,
		_w264_
	);
	LUT3 #(
		.INIT('h40)
	) name141 (
		\g1212_reg/NET0131 ,
		\g1275_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w265_
	);
	LUT4 #(
		.INIT('h80a0)
	) name142 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1235_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w266_
	);
	LUT2 #(
		.INIT('he)
	) name143 (
		_w265_,
		_w266_,
		_w267_
	);
	LUT3 #(
		.INIT('h40)
	) name144 (
		\g1212_reg/NET0131 ,
		\g1235_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w268_
	);
	LUT4 #(
		.INIT('h80a0)
	) name145 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1240_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w269_
	);
	LUT2 #(
		.INIT('he)
	) name146 (
		_w268_,
		_w269_,
		_w270_
	);
	LUT3 #(
		.INIT('h40)
	) name147 (
		\g1212_reg/NET0131 ,
		\g1240_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w271_
	);
	LUT4 #(
		.INIT('h80a0)
	) name148 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w272_
	);
	LUT2 #(
		.INIT('he)
	) name149 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT3 #(
		.INIT('h40)
	) name150 (
		\g1212_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w274_
	);
	LUT4 #(
		.INIT('h80a0)
	) name151 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1250_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w275_
	);
	LUT2 #(
		.INIT('he)
	) name152 (
		_w274_,
		_w275_,
		_w276_
	);
	LUT3 #(
		.INIT('h40)
	) name153 (
		\g1212_reg/NET0131 ,
		\g1250_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w277_
	);
	LUT4 #(
		.INIT('h80a0)
	) name154 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1255_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w278_
	);
	LUT2 #(
		.INIT('he)
	) name155 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT3 #(
		.INIT('h40)
	) name156 (
		\g1212_reg/NET0131 ,
		\g1255_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w280_
	);
	LUT4 #(
		.INIT('h80a0)
	) name157 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1260_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w281_
	);
	LUT2 #(
		.INIT('he)
	) name158 (
		_w280_,
		_w281_,
		_w282_
	);
	LUT3 #(
		.INIT('h40)
	) name159 (
		\g1212_reg/NET0131 ,
		\g1260_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w283_
	);
	LUT4 #(
		.INIT('h80a0)
	) name160 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1265_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w284_
	);
	LUT2 #(
		.INIT('he)
	) name161 (
		_w283_,
		_w284_,
		_w285_
	);
	LUT3 #(
		.INIT('h40)
	) name162 (
		\g1212_reg/NET0131 ,
		\g1265_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w286_
	);
	LUT4 #(
		.INIT('h80a0)
	) name163 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1270_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w287_
	);
	LUT2 #(
		.INIT('he)
	) name164 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT3 #(
		.INIT('h40)
	) name165 (
		\g1212_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w289_
	);
	LUT4 #(
		.INIT('h80a0)
	) name166 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1280_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w290_
	);
	LUT2 #(
		.INIT('he)
	) name167 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT3 #(
		.INIT('h40)
	) name168 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1292_reg/NET0131 ,
		_w292_
	);
	LUT4 #(
		.INIT('h80a0)
	) name169 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w293_
	);
	LUT2 #(
		.INIT('he)
	) name170 (
		_w292_,
		_w293_,
		_w294_
	);
	LUT3 #(
		.INIT('h40)
	) name171 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1296_reg/NET0131 ,
		_w295_
	);
	LUT4 #(
		.INIT('h8a00)
	) name172 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1292_reg/NET0131 ,
		_w296_
	);
	LUT2 #(
		.INIT('he)
	) name173 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT3 #(
		.INIT('h40)
	) name174 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		_w298_
	);
	LUT4 #(
		.INIT('h8a00)
	) name175 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1296_reg/NET0131 ,
		_w299_
	);
	LUT2 #(
		.INIT('he)
	) name176 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT3 #(
		.INIT('h40)
	) name177 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w301_
	);
	LUT4 #(
		.INIT('h8a00)
	) name178 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		_w302_
	);
	LUT2 #(
		.INIT('he)
	) name179 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT3 #(
		.INIT('h40)
	) name180 (
		\g1212_reg/NET0131 ,
		\g1270_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w304_
	);
	LUT4 #(
		.INIT('h8a00)
	) name181 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w305_
	);
	LUT2 #(
		.INIT('he)
	) name182 (
		_w304_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		\g109_pad ,
		\g243_reg/NET0131 ,
		_w307_
	);
	LUT3 #(
		.INIT('h02)
	) name184 (
		\g109_pad ,
		\g1718_reg/NET0131 ,
		\g4173_pad ,
		_w308_
	);
	LUT3 #(
		.INIT('h60)
	) name185 (
		\g4175_pad ,
		_w190_,
		_w224_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		\g109_pad ,
		\g1400_reg/NET0131 ,
		_w310_
	);
	LUT2 #(
		.INIT('he)
	) name187 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w311_
	);
	LUT3 #(
		.INIT('h80)
	) name188 (
		\g109_pad ,
		\g741_pad ,
		\g742_pad ,
		_w312_
	);
	LUT3 #(
		.INIT('h80)
	) name189 (
		\g109_pad ,
		\g743_pad ,
		\g744_pad ,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\g109_pad ,
		\g1374_reg/NET0131 ,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		\g109_pad ,
		\g197_reg/NET0131 ,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\g109_pad ,
		\g201_reg/NET0131 ,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\g109_pad ,
		\g1389_reg/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\g109_pad ,
		\g1397_reg/NET0131 ,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\g109_pad ,
		\g192_reg/NET0131 ,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\g109_pad ,
		\g248_reg/NET0131 ,
		_w320_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name197 (
		\g1718_reg/NET0131 ,
		\g4180_pad ,
		\g4181_pad ,
		_w194_,
		_w321_
	);
	LUT3 #(
		.INIT('h60)
	) name198 (
		\g971_reg/NET0131 ,
		_w144_,
		_w146_,
		_w322_
	);
	LUT4 #(
		.INIT('h9a00)
	) name199 (
		\g1336_reg/NET0131 ,
		_w206_,
		_w209_,
		_w212_,
		_w323_
	);
	LUT4 #(
		.INIT('h8a00)
	) name200 (
		\g1341_reg/NET0131 ,
		_w206_,
		_w209_,
		_w212_,
		_w324_
	);
	LUT2 #(
		.INIT('h6)
	) name201 (
		\g1336_reg/NET0131 ,
		\g1341_reg/NET0131 ,
		_w325_
	);
	LUT4 #(
		.INIT('h4000)
	) name202 (
		_w206_,
		_w209_,
		_w212_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('he)
	) name203 (
		_w324_,
		_w326_,
		_w327_
	);
	LUT4 #(
		.INIT('heee2)
	) name204 (
		\g305_reg/NET0131 ,
		_w124_,
		_w129_,
		_w130_,
		_w328_
	);
	assign \g21280/_0_  = _w148_ ;
	assign \g21281/_0_  = _w150_ ;
	assign \g21282/_0_  = _w152_ ;
	assign \g21307/_0_  = _w164_ ;
	assign \g21322/_0_  = _w166_ ;
	assign \g21333/_0_  = _w168_ ;
	assign \g21334/_0_  = _w169_ ;
	assign \g21338/_0_  = _w171_ ;
	assign \g21350/_0_  = _w172_ ;
	assign \g21355/_0_  = _w174_ ;
	assign \g21356/_0_  = _w175_ ;
	assign \g21357/_0_  = _w176_ ;
	assign \g21358/_1_  = _w167_ ;
	assign \g21359/_0_  = _w178_ ;
	assign \g21370/_0_  = _w179_ ;
	assign \g21371/_0_  = _w180_ ;
	assign \g21378/_0_  = _w181_ ;
	assign \g21379/_0_  = _w182_ ;
	assign \g21380/_1_  = _w173_ ;
	assign \g21381/_0_  = _w184_ ;
	assign \g21390/_0_  = _w185_ ;
	assign \g21394/_0_  = _w186_ ;
	assign \g21396/_0_  = _w188_ ;
	assign \g21397/_0_  = _w189_ ;
	assign \g21398/_1_  = _w165_ ;
	assign \g21412/_0_  = _w197_ ;
	assign \g21413/_0_  = _w198_ ;
	assign \g21419/_0_  = _w199_ ;
	assign \g21420/_00_  = _w216_ ;
	assign \g21421/_00_  = _w221_ ;
	assign \g21424/_0_  = _w222_ ;
	assign \g21425/_0_  = _w223_ ;
	assign \g21426/_1_  = _w170_ ;
	assign \g21437/_0_  = _w225_ ;
	assign \g21444/_0_  = _w226_ ;
	assign \g21450/_0_  = _w227_ ;
	assign \g21455/_0_  = _w228_ ;
	assign \g21457/_0_  = _w229_ ;
	assign \g21458/_1_  = _w177_ ;
	assign \g21459/_0_  = _w230_ ;
	assign \g21470/_0_  = _w231_ ;
	assign \g21486/_0_  = _w232_ ;
	assign \g21487/_0_  = _w233_ ;
	assign \g21495/_0_  = _w234_ ;
	assign \g21498/_1_  = _w183_ ;
	assign \g21499/_0_  = _w238_ ;
	assign \g21500/_0_  = _w239_ ;
	assign \g21502/_0_  = _w242_ ;
	assign \g21503/_0_  = _w243_ ;
	assign \g21508/_0_  = _w245_ ;
	assign \g21509/_0_  = _w247_ ;
	assign \g21510/_0_  = _w250_ ;
	assign \g21511/_0_  = _w252_ ;
	assign \g21515/_0_  = _w255_ ;
	assign \g21520/_0_  = _w256_ ;
	assign \g21523/_0_  = _w257_ ;
	assign \g21524/_0_  = _w258_ ;
	assign \g21525/_0_  = _w259_ ;
	assign \g21538/_0_  = _w187_ ;
	assign \g21544/_0_  = _w260_ ;
	assign \g21550/_1_  = _w151_ ;
	assign \g21562/_0_  = _w261_ ;
	assign \g21563/_0_  = _w262_ ;
	assign \g21584/_0_  = _w218_ ;
	assign \g21591/_0_  = _w263_ ;
	assign \g21593/_0_  = _w264_ ;
	assign \g21601/_3_  = _w267_ ;
	assign \g21603/_3_  = _w270_ ;
	assign \g21605/_3_  = _w273_ ;
	assign \g21607/_3_  = _w276_ ;
	assign \g21609/_3_  = _w279_ ;
	assign \g21611/_3_  = _w282_ ;
	assign \g21613/_3_  = _w285_ ;
	assign \g21615/_3_  = _w288_ ;
	assign \g21617/_3_  = _w291_ ;
	assign \g21619/_3_  = _w294_ ;
	assign \g21621/_3_  = _w297_ ;
	assign \g21623/_3_  = _w300_ ;
	assign \g21625/_3_  = _w303_ ;
	assign \g21627/_3_  = _w306_ ;
	assign \g21640/_0_  = _w307_ ;
	assign \g21641/_0_  = _w308_ ;
	assign \g21642/_0_  = _w309_ ;
	assign \g21693/_0_  = _w310_ ;
	assign \g21694/_0_  = _w311_ ;
	assign \g21735/_2_  = _w312_ ;
	assign \g21745/_2_  = _w313_ ;
	assign \g21796/_0_  = _w314_ ;
	assign \g21799/_0_  = _w315_ ;
	assign \g21803/_0_  = _w316_ ;
	assign \g21812/_0_  = _w317_ ;
	assign \g21814/_0_  = _w318_ ;
	assign \g21816/_0_  = _w319_ ;
	assign \g21828/_0_  = _w320_ ;
	assign \g22203/_0_  = _w321_ ;
	assign \g22260/_1_  = _w144_ ;
	assign \g22317/_0_  = _w322_ ;
	assign \g22339/_0_  = _w323_ ;
	assign \g22392/_0_  = _w327_ ;
	assign \g22395/_1_  = _w210_ ;
	assign \g2601_pad  = 1'b0;
	assign \g27_dup/_0_  = _w328_ ;
	assign \g5816_pad  = 1'b1;
endmodule;