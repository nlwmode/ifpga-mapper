module top( \V10_0_pad  , \V11_0_pad  , \V12_0_pad  , \V13_0_pad  , \V14_0_pad  , \V15_0_pad  , \V16_0_pad  , \V17_0_pad  , \V18_0_pad  , \V22_2_pad  , \V22_3_pad  , \V22_4_pad  , \V22_5_pad  , \V27_0_pad  , \V27_3_pad  , \V29_0_pad  , \V7_1_pad  , \V7_2_pad  , \V7_3_pad  , \V7_4_pad  , \V7_5_pad  , \V7_6_pad  , \V7_7_pad  , \V8_0_pad  , \V9_0_pad  , \V27_1_pad  , \V27_2_pad  , \V27_4_pad  , \V28_0_pad  , \V30_0_pad  , \V32_0_pad  , \V33_0_pad  , \V34_0_pad  , \V35_0_pad  , \V36_0_pad  , \V37_0_pad  , \V38_0_pad  );
  input \V10_0_pad  ;
  input \V11_0_pad  ;
  input \V12_0_pad  ;
  input \V13_0_pad  ;
  input \V14_0_pad  ;
  input \V15_0_pad  ;
  input \V16_0_pad  ;
  input \V17_0_pad  ;
  input \V18_0_pad  ;
  input \V22_2_pad  ;
  input \V22_3_pad  ;
  input \V22_4_pad  ;
  input \V22_5_pad  ;
  input \V27_0_pad  ;
  input \V27_3_pad  ;
  input \V29_0_pad  ;
  input \V7_1_pad  ;
  input \V7_2_pad  ;
  input \V7_3_pad  ;
  input \V7_4_pad  ;
  input \V7_5_pad  ;
  input \V7_6_pad  ;
  input \V7_7_pad  ;
  input \V8_0_pad  ;
  input \V9_0_pad  ;
  output \V27_1_pad  ;
  output \V27_2_pad  ;
  output \V27_4_pad  ;
  output \V28_0_pad  ;
  output \V30_0_pad  ;
  output \V32_0_pad  ;
  output \V33_0_pad  ;
  output \V34_0_pad  ;
  output \V35_0_pad  ;
  output \V36_0_pad  ;
  output \V37_0_pad  ;
  output \V38_0_pad  ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n26 = ~\V7_5_pad  & ~\V7_6_pad  ;
  assign n27 = ~\V7_7_pad  & n26 ;
  assign n28 = ~\V7_1_pad  & ~\V7_2_pad  ;
  assign n29 = ~\V7_3_pad  & ~\V7_4_pad  ;
  assign n30 = n28 & n29 ;
  assign n31 = n27 & n30 ;
  assign n32 = \V29_0_pad  & \V8_0_pad  ;
  assign n33 = \V9_0_pad  & n32 ;
  assign n34 = n31 & n33 ;
  assign n35 = \V29_0_pad  & ~\V8_0_pad  ;
  assign n36 = ~\V9_0_pad  & n35 ;
  assign n37 = n31 & n36 ;
  assign n38 = ~\V27_0_pad  & \V29_0_pad  ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = ~n34 & n39 ;
  assign n41 = ~\V9_0_pad  & n32 ;
  assign n42 = n31 & n41 ;
  assign n43 = \V27_0_pad  & \V29_0_pad  ;
  assign n44 = ~n31 & n43 ;
  assign n45 = ~n42 & ~n44 ;
  assign n46 = ~\V22_2_pad  & ~\V27_3_pad  ;
  assign n47 = n31 & n35 ;
  assign n48 = ~\V10_0_pad  & ~n47 ;
  assign n49 = \V18_0_pad  & \V22_5_pad  ;
  assign n50 = \V11_0_pad  & \V22_5_pad  ;
  assign n51 = \V14_0_pad  & ~\V22_5_pad  ;
  assign n52 = \V22_3_pad  & n51 ;
  assign n53 = \V17_0_pad  & ~\V22_5_pad  ;
  assign n54 = \V22_3_pad  & n53 ;
  assign n55 = \V22_4_pad  & n51 ;
  assign n56 = \V22_4_pad  & n53 ;
  assign n57 = \V16_0_pad  & ~\V22_5_pad  ;
  assign n58 = ~\V12_0_pad  & ~\V13_0_pad  ;
  assign n59 = ~\V14_0_pad  & ~\V15_0_pad  ;
  assign n60 = n58 & n59 ;
  assign \V27_1_pad  = ~n40 ;
  assign \V27_2_pad  = ~n45 ;
  assign \V27_4_pad  = ~n46 ;
  assign \V28_0_pad  = ~n48 ;
  assign \V30_0_pad  = n49 ;
  assign \V32_0_pad  = n50 ;
  assign \V33_0_pad  = n52 ;
  assign \V34_0_pad  = n54 ;
  assign \V35_0_pad  = n55 ;
  assign \V36_0_pad  = n56 ;
  assign \V37_0_pad  = n57 ;
  assign \V38_0_pad  = ~n60 ;
endmodule
