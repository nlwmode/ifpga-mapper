module top( \dest_x[0]  , \dest_x[1]  , \dest_x[2]  , \dest_x[3]  , \dest_x[4]  , \dest_x[5]  , \dest_x[6]  , \dest_x[7]  , \dest_x[8]  , \dest_x[9]  , \dest_x[10]  , \dest_x[11]  , \dest_x[12]  , \dest_x[13]  , \dest_x[14]  , \dest_x[15]  , \dest_x[16]  , \dest_x[17]  , \dest_x[18]  , \dest_x[19]  , \dest_x[20]  , \dest_x[21]  , \dest_x[22]  , \dest_x[23]  , \dest_x[24]  , \dest_x[25]  , \dest_x[26]  , \dest_x[27]  , \dest_x[28]  , \dest_x[29]  , \dest_y[0]  , \dest_y[1]  , \dest_y[2]  , \dest_y[3]  , \dest_y[4]  , \dest_y[5]  , \dest_y[6]  , \dest_y[7]  , \dest_y[8]  , \dest_y[9]  , \dest_y[10]  , \dest_y[11]  , \dest_y[12]  , \dest_y[13]  , \dest_y[14]  , \dest_y[15]  , \dest_y[16]  , \dest_y[17]  , \dest_y[18]  , \dest_y[19]  , \dest_y[20]  , \dest_y[21]  , \dest_y[22]  , \dest_y[23]  , \dest_y[24]  , \dest_y[25]  , \dest_y[26]  , \dest_y[27]  , \dest_y[28]  , \dest_y[29]  , \outport[0]  , \outport[1]  , \outport[2]  , \outport[3]  , \outport[4]  , \outport[5]  , \outport[6]  , \outport[7]  , \outport[8]  , \outport[9]  , \outport[10]  , \outport[11]  , \outport[12]  , \outport[13]  , \outport[14]  , \outport[15]  , \outport[16]  , \outport[17]  , \outport[18]  , \outport[19]  , \outport[20]  , \outport[21]  , \outport[22]  , \outport[23]  , \outport[24]  , \outport[25]  , \outport[26]  , \outport[27]  , \outport[28]  , \outport[29]  );
  input \dest_x[0]  ;
  input \dest_x[1]  ;
  input \dest_x[2]  ;
  input \dest_x[3]  ;
  input \dest_x[4]  ;
  input \dest_x[5]  ;
  input \dest_x[6]  ;
  input \dest_x[7]  ;
  input \dest_x[8]  ;
  input \dest_x[9]  ;
  input \dest_x[10]  ;
  input \dest_x[11]  ;
  input \dest_x[12]  ;
  input \dest_x[13]  ;
  input \dest_x[14]  ;
  input \dest_x[15]  ;
  input \dest_x[16]  ;
  input \dest_x[17]  ;
  input \dest_x[18]  ;
  input \dest_x[19]  ;
  input \dest_x[20]  ;
  input \dest_x[21]  ;
  input \dest_x[22]  ;
  input \dest_x[23]  ;
  input \dest_x[24]  ;
  input \dest_x[25]  ;
  input \dest_x[26]  ;
  input \dest_x[27]  ;
  input \dest_x[28]  ;
  input \dest_x[29]  ;
  input \dest_y[0]  ;
  input \dest_y[1]  ;
  input \dest_y[2]  ;
  input \dest_y[3]  ;
  input \dest_y[4]  ;
  input \dest_y[5]  ;
  input \dest_y[6]  ;
  input \dest_y[7]  ;
  input \dest_y[8]  ;
  input \dest_y[9]  ;
  input \dest_y[10]  ;
  input \dest_y[11]  ;
  input \dest_y[12]  ;
  input \dest_y[13]  ;
  input \dest_y[14]  ;
  input \dest_y[15]  ;
  input \dest_y[16]  ;
  input \dest_y[17]  ;
  input \dest_y[18]  ;
  input \dest_y[19]  ;
  input \dest_y[20]  ;
  input \dest_y[21]  ;
  input \dest_y[22]  ;
  input \dest_y[23]  ;
  input \dest_y[24]  ;
  input \dest_y[25]  ;
  input \dest_y[26]  ;
  input \dest_y[27]  ;
  input \dest_y[28]  ;
  input \dest_y[29]  ;
  output \outport[0]  ;
  output \outport[1]  ;
  output \outport[2]  ;
  output \outport[3]  ;
  output \outport[4]  ;
  output \outport[5]  ;
  output \outport[6]  ;
  output \outport[7]  ;
  output \outport[8]  ;
  output \outport[9]  ;
  output \outport[10]  ;
  output \outport[11]  ;
  output \outport[12]  ;
  output \outport[13]  ;
  output \outport[14]  ;
  output \outport[15]  ;
  output \outport[16]  ;
  output \outport[17]  ;
  output \outport[18]  ;
  output \outport[19]  ;
  output \outport[20]  ;
  output \outport[21]  ;
  output \outport[22]  ;
  output \outport[23]  ;
  output \outport[24]  ;
  output \outport[25]  ;
  output \outport[26]  ;
  output \outport[27]  ;
  output \outport[28]  ;
  output \outport[29]  ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 ;
  assign n61 = \dest_x[22]  & ~\dest_x[23]  ;
  assign n62 = \dest_x[14]  & \dest_x[15]  ;
  assign n63 = ~\dest_x[16]  & ~\dest_x[18]  ;
  assign n64 = ~n62 & n63 ;
  assign n65 = ~\dest_x[9]  & ~\dest_x[10]  ;
  assign n66 = \dest_x[11]  & ~n65 ;
  assign n67 = ~\dest_x[12]  & ~\dest_x[13]  ;
  assign n68 = n63 & n67 ;
  assign n69 = ~n66 & n68 ;
  assign n70 = ~n64 & ~n69 ;
  assign n71 = ~\dest_x[17]  & ~\dest_x[18]  ;
  assign n72 = \dest_x[19]  & \dest_x[20]  ;
  assign n73 = ~n71 & n72 ;
  assign n74 = n70 & n73 ;
  assign n75 = ~\dest_x[21]  & ~n74 ;
  assign n76 = \dest_x[8]  & \dest_x[11]  ;
  assign n77 = \dest_x[6]  & \dest_x[7]  ;
  assign n78 = n76 & n77 ;
  assign n79 = \dest_x[4]  & \dest_x[5]  ;
  assign n80 = \dest_x[2]  & \dest_x[3]  ;
  assign n81 = n79 & n80 ;
  assign n82 = n78 & n81 ;
  assign n83 = \dest_x[17]  & ~\dest_x[18]  ;
  assign n84 = \dest_x[0]  & \dest_x[1]  ;
  assign n85 = n65 & n84 ;
  assign n86 = n83 & n85 ;
  assign n87 = n82 & n86 ;
  assign n88 = \dest_x[24]  & \dest_x[25]  ;
  assign n89 = \dest_x[20]  & ~\dest_x[21]  ;
  assign n90 = n88 & n89 ;
  assign n91 = \dest_x[19]  & ~\dest_x[26]  ;
  assign n92 = ~\dest_x[12]  & \dest_x[15]  ;
  assign n93 = n91 & n92 ;
  assign n94 = n90 & n93 ;
  assign n95 = \dest_x[27]  & \dest_x[28]  ;
  assign n96 = \dest_x[29]  & n95 ;
  assign n97 = n94 & n96 ;
  assign n98 = n87 & n97 ;
  assign n99 = ~\dest_x[16]  & ~n62 ;
  assign n100 = ~\dest_x[16]  & n67 ;
  assign n101 = ~n66 & n100 ;
  assign n102 = ~n99 & ~n101 ;
  assign n103 = \dest_x[14]  & ~n67 ;
  assign n104 = \dest_x[11]  & \dest_x[14]  ;
  assign n105 = ~n65 & n104 ;
  assign n106 = ~n103 & ~n105 ;
  assign n107 = \dest_x[11]  & \dest_x[13]  ;
  assign n108 = ~n65 & n107 ;
  assign n109 = \dest_x[12]  & \dest_x[13]  ;
  assign n110 = ~\dest_x[14]  & ~n109 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = n106 & ~n111 ;
  assign n113 = ~n102 & n112 ;
  assign n114 = n98 & n113 ;
  assign n115 = ~n75 & n114 ;
  assign n116 = n61 & n115 ;
  assign n117 = ~\dest_x[22]  & \dest_x[23]  ;
  assign n118 = ~\dest_x[21]  & n117 ;
  assign n119 = ~n74 & n118 ;
  assign n120 = n114 & n119 ;
  assign n121 = ~n116 & ~n120 ;
  assign n122 = \dest_x[23]  & n88 ;
  assign n123 = ~\dest_x[26]  & ~n122 ;
  assign n124 = ~\dest_x[21]  & ~\dest_x[22]  ;
  assign n125 = ~\dest_x[26]  & n124 ;
  assign n126 = ~n74 & n125 ;
  assign n127 = ~n123 & ~n126 ;
  assign n128 = n96 & n127 ;
  assign n129 = n121 & ~n128 ;
  assign n130 = ~n74 & n124 ;
  assign n131 = \dest_x[23]  & ~n130 ;
  assign n132 = \dest_x[22]  & ~n75 ;
  assign n133 = \dest_x[9]  & ~\dest_x[10]  ;
  assign n134 = ~\dest_x[7]  & n133 ;
  assign n135 = \dest_x[11]  & ~\dest_x[12]  ;
  assign n136 = ~\dest_x[8]  & ~\dest_x[13]  ;
  assign n137 = n135 & n136 ;
  assign n138 = n134 & n137 ;
  assign n139 = n90 & n138 ;
  assign n140 = ~\dest_x[1]  & ~\dest_x[2]  ;
  assign n141 = n83 & n140 ;
  assign n142 = ~\dest_x[5]  & ~\dest_x[6]  ;
  assign n143 = ~\dest_x[3]  & ~\dest_x[4]  ;
  assign n144 = n142 & n143 ;
  assign n145 = n141 & n144 ;
  assign n146 = n139 & n145 ;
  assign n147 = ~\dest_x[14]  & ~\dest_x[15]  ;
  assign n148 = ~\dest_x[12]  & n147 ;
  assign n149 = ~n66 & n148 ;
  assign n150 = \dest_x[16]  & ~n149 ;
  assign n151 = n102 & ~n150 ;
  assign n152 = n146 & n151 ;
  assign n153 = \dest_x[19]  & ~n71 ;
  assign n154 = n70 & n153 ;
  assign n155 = \dest_x[23]  & \dest_x[26]  ;
  assign n156 = n88 & n155 ;
  assign n157 = n154 & ~n156 ;
  assign n158 = n152 & n157 ;
  assign n159 = ~n132 & n158 ;
  assign n160 = n131 & n159 ;
  assign n161 = n128 & ~n160 ;
  assign n162 = ~n129 & ~n161 ;
  assign n163 = \dest_y[23]  & \dest_y[25]  ;
  assign n164 = \dest_y[24]  & n163 ;
  assign n165 = ~\dest_y[26]  & ~n164 ;
  assign n166 = \dest_y[14]  & \dest_y[15]  ;
  assign n167 = ~\dest_y[16]  & ~\dest_y[18]  ;
  assign n168 = ~n166 & n167 ;
  assign n169 = ~\dest_y[9]  & ~\dest_y[10]  ;
  assign n170 = \dest_y[11]  & ~n169 ;
  assign n171 = ~\dest_y[12]  & ~\dest_y[13]  ;
  assign n172 = n167 & n171 ;
  assign n173 = ~n170 & n172 ;
  assign n174 = ~n168 & ~n173 ;
  assign n175 = ~\dest_y[17]  & ~\dest_y[18]  ;
  assign n176 = \dest_y[19]  & \dest_y[20]  ;
  assign n177 = ~n175 & n176 ;
  assign n178 = n174 & n177 ;
  assign n179 = ~\dest_y[21]  & ~\dest_y[22]  ;
  assign n180 = ~\dest_y[26]  & n179 ;
  assign n181 = ~n178 & n180 ;
  assign n182 = ~n165 & ~n181 ;
  assign n183 = \dest_y[28]  & \dest_y[29]  ;
  assign n184 = \dest_y[27]  & n183 ;
  assign n185 = n182 & n184 ;
  assign n186 = \dest_x[0]  & ~n185 ;
  assign n187 = ~n129 & ~n186 ;
  assign n188 = ~n161 & ~n187 ;
  assign n189 = \dest_y[19]  & ~n175 ;
  assign n190 = n174 & n189 ;
  assign n191 = \dest_y[12]  & \dest_y[13]  ;
  assign n192 = \dest_y[11]  & \dest_y[13]  ;
  assign n193 = ~n169 & n192 ;
  assign n194 = ~n191 & ~n193 ;
  assign n195 = ~\dest_y[22]  & \dest_y[23]  ;
  assign n196 = ~\dest_y[18]  & \dest_y[19]  ;
  assign n197 = n195 & n196 ;
  assign n198 = \dest_y[15]  & ~\dest_y[16]  ;
  assign n199 = \dest_y[11]  & ~\dest_y[12]  ;
  assign n200 = n198 & n199 ;
  assign n201 = n197 & n200 ;
  assign n202 = n194 & n201 ;
  assign n203 = ~\dest_y[7]  & ~\dest_y[8]  ;
  assign n204 = ~\dest_y[5]  & ~\dest_y[6]  ;
  assign n205 = n203 & n204 ;
  assign n206 = ~\dest_y[3]  & ~\dest_y[4]  ;
  assign n207 = ~\dest_y[1]  & ~\dest_y[2]  ;
  assign n208 = n206 & n207 ;
  assign n209 = n205 & n208 ;
  assign n210 = \dest_y[9]  & ~\dest_y[10]  ;
  assign n211 = \dest_y[17]  & n210 ;
  assign n212 = n209 & n211 ;
  assign n213 = n202 & n212 ;
  assign n214 = \dest_y[14]  & ~n171 ;
  assign n215 = \dest_y[11]  & \dest_y[14]  ;
  assign n216 = ~n169 & n215 ;
  assign n217 = ~n214 & ~n216 ;
  assign n218 = ~\dest_y[20]  & \dest_y[21]  ;
  assign n219 = ~n217 & n218 ;
  assign n220 = n213 & n219 ;
  assign n221 = ~n190 & n220 ;
  assign n222 = \dest_y[20]  & ~n217 ;
  assign n223 = n213 & n222 ;
  assign n224 = ~\dest_y[21]  & n190 ;
  assign n225 = n223 & n224 ;
  assign n226 = ~n221 & ~n225 ;
  assign n227 = ~\dest_y[23]  & \dest_y[24]  ;
  assign n228 = \dest_y[24]  & n179 ;
  assign n229 = ~n178 & n228 ;
  assign n230 = ~n227 & ~n229 ;
  assign n231 = ~n178 & n179 ;
  assign n232 = \dest_y[23]  & ~\dest_y[24]  ;
  assign n233 = ~n231 & n232 ;
  assign n234 = n230 & ~n233 ;
  assign n235 = ~n226 & n234 ;
  assign n236 = \dest_y[26]  & n164 ;
  assign n237 = ~n231 & n236 ;
  assign n238 = ~\dest_x[0]  & ~\dest_y[0]  ;
  assign n239 = ~n237 & n238 ;
  assign n240 = n164 & ~n231 ;
  assign n241 = \dest_y[23]  & \dest_y[24]  ;
  assign n242 = ~\dest_y[25]  & ~n241 ;
  assign n243 = ~\dest_y[25]  & n179 ;
  assign n244 = ~n178 & n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = ~n240 & n245 ;
  assign n247 = n239 & ~n246 ;
  assign n248 = n235 & n247 ;
  assign n249 = n185 & ~n248 ;
  assign n250 = ~\dest_y[27]  & ~n237 ;
  assign n251 = ~n231 & n241 ;
  assign n252 = ~\dest_y[20]  & ~n190 ;
  assign n253 = ~n251 & ~n252 ;
  assign n254 = ~\dest_y[23]  & ~\dest_y[24]  ;
  assign n255 = ~\dest_y[24]  & n179 ;
  assign n256 = ~n178 & n255 ;
  assign n257 = ~n254 & ~n256 ;
  assign n258 = ~\dest_y[17]  & n217 ;
  assign n259 = n169 & n183 ;
  assign n260 = \dest_y[14]  & ~\dest_y[21]  ;
  assign n261 = \dest_y[8]  & ~\dest_y[13]  ;
  assign n262 = n260 & n261 ;
  assign n263 = \dest_y[6]  & \dest_y[7]  ;
  assign n264 = \dest_y[4]  & \dest_y[5]  ;
  assign n265 = n263 & n264 ;
  assign n266 = n262 & n265 ;
  assign n267 = n259 & n266 ;
  assign n268 = \dest_y[2]  & \dest_y[3]  ;
  assign n269 = \dest_y[0]  & \dest_y[1]  ;
  assign n270 = n268 & n269 ;
  assign n271 = n201 & n270 ;
  assign n272 = n267 & n271 ;
  assign n273 = ~n258 & n272 ;
  assign n274 = \dest_y[17]  & ~n217 ;
  assign n275 = ~n178 & ~n274 ;
  assign n276 = n273 & n275 ;
  assign n277 = n257 & n276 ;
  assign n278 = n253 & n277 ;
  assign n279 = \dest_y[27]  & n182 ;
  assign n280 = n246 & ~n279 ;
  assign n281 = n278 & n280 ;
  assign n282 = ~n250 & n281 ;
  assign n283 = ~n161 & ~n282 ;
  assign n284 = ~n249 & n283 ;
  assign n285 = ~n188 & ~n284 ;
  assign n286 = \dest_x[0]  & \dest_y[0]  ;
  assign n287 = ~n237 & ~n286 ;
  assign n288 = ~n246 & n287 ;
  assign n289 = n235 & n288 ;
  assign n290 = n185 & ~n289 ;
  assign n291 = n162 & n290 ;
  assign \outport[0]  = ~n162 ;
  assign \outport[1]  = ~n285 ;
  assign \outport[2]  = n291 ;
  assign \outport[3]  = 1'b0 ;
  assign \outport[4]  = 1'b0 ;
  assign \outport[5]  = 1'b0 ;
  assign \outport[6]  = 1'b0 ;
  assign \outport[7]  = 1'b0 ;
  assign \outport[8]  = 1'b0 ;
  assign \outport[9]  = 1'b0 ;
  assign \outport[10]  = 1'b0 ;
  assign \outport[11]  = 1'b0 ;
  assign \outport[12]  = 1'b0 ;
  assign \outport[13]  = 1'b0 ;
  assign \outport[14]  = 1'b0 ;
  assign \outport[15]  = 1'b0 ;
  assign \outport[16]  = 1'b0 ;
  assign \outport[17]  = 1'b0 ;
  assign \outport[18]  = 1'b0 ;
  assign \outport[19]  = 1'b0 ;
  assign \outport[20]  = 1'b0 ;
  assign \outport[21]  = 1'b0 ;
  assign \outport[22]  = 1'b0 ;
  assign \outport[23]  = 1'b0 ;
  assign \outport[24]  = 1'b0 ;
  assign \outport[25]  = 1'b0 ;
  assign \outport[26]  = 1'b0 ;
  assign \outport[27]  = 1'b0 ;
  assign \outport[28]  = 1'b0 ;
  assign \outport[29]  = 1'b0 ;
endmodule
