module top (\n1035gat_reg/NET0131 , \n1045gat_reg/NET0131 , \n1068gat_reg/NET0131 , \n1072gat_reg/NET0131 , \n1080gat_reg/NET0131 , \n1121gat_reg/NET0131 , \n1135gat_reg/NET0131 , \n1148gat_reg/NET0131 , \n1197gat_reg/NET0131 , \n1226gat_reg/NET0131 , \n1241gat_reg/NET0131 , \n1282gat_reg/NET0131 , \n1294gat_reg/NET0131 , \n1312gat_reg/NET0131 , \n1316gat_reg/NET0131 , \n1332gat_reg/NET0131 , \n1336gat_reg/NET0131 , \n1340gat_reg/NET0131 , \n1363gat_reg/NET0131 , \n1389gat_reg/NET0131 , \n1394gat_reg/NET0131 , \n1433gat_reg/NET0131 , \n1456gat_reg/NET0131 , \n1462gat_reg/NET0131 , \n148gat_reg/NET0131 , \n1496gat_reg/NET0131 , \n1508gat_reg/NET0131 , \n1525gat_reg/NET0131 , \n152gat_reg/NET0131 , \n156gat_reg/NET0131 , \n1588gat_reg/NET0131 , \n1596gat_reg/NET0131 , \n160gat_reg/NET0131 , \n1675gat_reg/NET0131 , \n1678gat_reg/NET0131 , \n1740gat_reg/NET0131 , \n1748gat_reg/NET0131 , \n1763gat_reg/NET0131 , \n1767gat_reg/NET0131 , \n1771gat_reg/NET0131 , \n1775gat_reg/NET0131 , \n1807gat_reg/NET0131 , \n1821gat_reg/NET0131 , \n1829gat_reg/NET0131 , \n1834gat_reg/NET0131 , \n1850gat_reg/NET0131 , \n1871gat_reg/NET0131 , \n1880gat_reg/NET0131 , \n1899gat_reg/NET0131 , \n1975gat_reg/NET0131 , \n2021gat_reg/NET0131 , \n2025gat_reg/NET0131 , \n2029gat_reg/NET0131 , \n2033gat_reg/NET0131 , \n2037gat_reg/NET0131 , \n2040gat_reg/NET0131 , \n2044gat_reg/NET0131 , \n2061gat_reg/NET0131 , \n2084gat_reg/NET0131 , \n2091gat_reg/NET0131 , \n2095gat_reg/NET0131 , \n2099gat_reg/NET0131 , \n2102gat_reg/NET0131 , \n2110gat_reg/NET0131 , \n2117gat_reg/NET0131 , \n2121gat_reg/NET0131 , \n2125gat_reg/NET0131 , \n2135gat_reg/NET0131 , \n2139gat_reg/NET0131 , \n2143gat_reg/NET0131 , \n2155gat_reg/NET0131 , \n2169gat_reg/NET0131 , \n2176gat_reg/NET0131 , \n2179gat_reg/NET0131 , \n2182gat_reg/NET0131 , \n2190gat_reg/NET0131 , \n2203gat_reg/NET0131 , \n2207gat_reg/NET0131 , \n2262gat_reg/NET0131 , \n2266gat_reg/NET0131 , \n2270gat_reg/NET0131 , \n2319gat_reg/NET0131 , \n2339gat_reg/NET0131 , \n2343gat_reg/NET0131 , \n2347gat_reg/NET0131 , \n2390gat_reg/NET0131 , \n2394gat_reg/NET0131 , \n2399gat_reg/NET0131 , \n2403gat_reg/NET0131 , \n2407gat_reg/NET0131 , \n2440gat_reg/NET0131 , \n2446gat_reg/NET0131 , \n2450gat_reg/NET0131 , \n2454gat_reg/NET0131 , \n2458gat_reg/NET0131 , \n2464gat_reg/NET0131 , \n2468gat_reg/NET0131 , \n2472gat_reg/NET0131 , \n2476gat_reg/NET0131 , \n2490gat_reg/NET0131 , \n2495gat_reg/NET0131 , \n2502gat_reg/NET0131 , \n2506gat_reg/NET0131 , \n2510gat_reg/NET0131 , \n2514gat_reg/NET0131 , \n2518gat_reg/NET0131 , \n2526gat_reg/NET0131 , \n2543gat_reg/NET0131 , \n2562gat_reg/NET0131 , \n256gat_reg/NET0131 , \n2588gat_reg/NET0131 , \n2592gat_reg/NET0131 , \n2599gat_reg/NET0131 , \n2622gat_reg/NET0131 , \n2626gat_reg/NET0131 , \n2630gat_reg/NET0131 , \n2634gat_reg/NET0131 , \n2640gat_reg/NET0131 , \n2644gat_reg/NET0131 , \n2658gat_reg/NET0131 , \n271gat_reg/NET0131 , \n3065gat_pad , \n3066gat_pad , \n3067gat_pad , \n3068gat_pad , \n3069gat_pad , \n3070gat_pad , \n3071gat_pad , \n3072gat_pad , \n3073gat_pad , \n3074gat_pad , \n3075gat_pad , \n3076gat_pad , \n3077gat_pad , \n3078gat_pad , \n3079gat_pad , \n3080gat_pad , \n3081gat_pad , \n3082gat_pad , \n3083gat_pad , \n3084gat_pad , \n3085gat_pad , \n3086gat_pad , \n3087gat_pad , \n3088gat_pad , \n3089gat_pad , \n3090gat_pad , \n3091gat_pad , \n3092gat_pad , \n3093gat_pad , \n3094gat_pad , \n3095gat_pad , \n3097gat_pad , \n3098gat_pad , \n3099gat_pad , \n3100gat_pad , \n314gat_reg/NET0131 , \n318gat_reg/NET0131 , \n322gat_reg/NET0131 , \n327gat_reg/NET0131 , \n331gat_reg/NET0131 , \n337gat_reg/NET0131 , \n341gat_reg/NET0131 , \n366gat_reg/NET0131 , \n384gat_reg/NET0131 , \n388gat_reg/NET0131 , \n398gat_reg/NET0131 , \n402gat_reg/NET0131 , \n463gat_reg/NET0131 , \n470gat_reg/NET0131 , \n553gat_reg/NET0131 , \n561gat_reg/NET0131 , \n580gat_reg/NET0131 , \n584gat_reg/NET0131 , \n614gat_reg/NET0131 , \n659gat_reg/NET0131 , \n667gat_reg/NET0131 , \n673gat_reg/NET0131 , \n680gat_reg/NET0131 , \n684gat_reg/NET0131 , \n699gat_reg/NET0131 , \n707gat_reg/NET0131 , \n777gat_reg/NET0131 , \n816gat_reg/NET0131 , \n820gat_reg/NET0131 , \n824gat_reg/NET0131 , \n830gat_reg/NET0131 , \n834gat_reg/NET0131 , \n838gat_reg/NET0131 , \n842gat_reg/NET0131 , \n846gat_reg/NET0131 , \n861gat_reg/NET0131 , \n865gat_reg/NET0131 , \n883gat_reg/NET0131 , \n919gat_reg/NET0131 , \n931gat_reg/NET0131 , \n957gat_reg/NET0131 , \_al_n0 , \g17_dup/_0_ , \g6952/_2_ , \g6953/_2_ , \g6961/_0_ , \g7076/_0_ , \g7077/_0_ , \g7079/_0_ , \g7081/_0_ , \g7082/_0_ , \g7083/_0_ , \g7146/_0_ , \g7147/_0_ , \g7148/_0_ , \g7149/_0_ , \g7150/_0_ , \g7151/_0_ , \g7152/_0_ , \g7153/_0_ , \g7154/_0_ , \g7156/_2_ , \g7161/_2_ , \g7165/_2_ , \g7174/_0_ , \g7180/_00_ , \g7182/_3_ , \g7191/_0_ , \g7204/_0_ , \g7209/_3_ , \g7220/_0_ , \g7229/_0_ , \g7233/_0_ , \g7234/_0_ , \g7235/_0_ , \g7236/_0_ , \g7237/_0_ , \g7238/_0_ , \g7241/_3_ , \g7264/_0_ , \g7265/_0_ , \g7266/_0_ , \g7267/_0_ , \g7268/_0_ , \g7301/_0_ , \g7326/_3_ , \g7350/_2_ , \g7352/_0_ , \g7356/_0_ , \g7359/_0_ , \g7389/_3_ , \g7417/_0_ , \g7418/_0_ , \g7419/_0_ , \g7444/_0_ , \g7445/_0_ , \g7449/_3_ , \g7451/_3_ , \g7454/_0_ , \g7467/_3_ , \g7476/_0_ , \g7480/_0_ , \g7494/_0_ , \g7509/_0_ , \g7514/_0_ , \g7517/_3_ , \g7524/_0_ , \g7558/_0_ , \g7560/_0_ , \g7561/_0_ , \g7563/_0_ , \g7567/_0_ , \g7572/_0_ , \g7579/_0_ , \g7605/_0_ , \g7625/_0_ , \g7627/_0_ , \g7671/_0_ , \g7675/_0_ , \g7689/_0_ , \g7697/_0_ , \g7743/_1_ , \g7764/_1_ , \g7769/_0_ , \g7771/_2_ , \g7779/_0_ , \g7852/_0_ , \g7873/_0_ , \g7884/_3_ , \g7889/_0_ , \g7902/_1_ , \g7992/_3_ , \g7994/_3_ , \g7996/_3_ , \g7998/_3_ , \g8000/_3_ , \g8002/_3_ , \g8004/_3_ , \g8006/_3_ , \g8008/_3_ , \g8150/_0_ , \g8151/_0_ , \g8157/_0_ , \g8163/_0_ , \g8172/_0_ , \g8197/_0_ , \g8211/_0_ , \g8223/_0_ , \g8237/_0_ , \g8251/_0_ , \g8261/_0_ , \g8272/_0_ , \g8287/_0_ , \g8647/_0_ , \g8671/_0_ , \g8672/_0_ , \g8735/_0_ , \g8766/_0_ , \g8811/_0_ , \g8821/_0_ , \g8856/_0_ , \g8858/_3_ , \g8868/_0_ , \g8880/_2_ , \g8886/_0_ , \g8900/_0_ , \g8932/_0_ , \g8991/_3_ , \g9014/_3_ , \g9074/_0_ , \g9091/_0_ , \g9105/_0_ , \g9107/_1_ , \g9111/_0_ , \n1332gat_reg/P0001 , \n1363gat_reg/P0001 , \n1394gat_reg/P0001 , \n1433gat_reg/P0001 , \n1775gat_reg/P0001 , \n2025gat_reg/P0001 , \n2029gat_reg/P0001 , \n2033gat_reg/P0001 , \n2044gat_reg/P0001 , \n2121gat_reg/P0001 , \n2125gat_reg/P0001 , \n2458gat_reg/P0001 , \n2472gat_reg/P0001 , \n2592gat_reg/P0001 , \n3104gat_pad , \n3105gat_pad , \n3106gat_pad , \n3107gat_pad , \n3108gat_pad , \n3109gat_pad , \n3110gat_pad , \n3111gat_pad , \n3112gat_pad , \n3113gat_pad , \n3114gat_pad , \n3116gat_pad , \n3117gat_pad , \n3118gat_pad , \n3119gat_pad , \n3120gat_pad , \n3121gat_pad , \n3122gat_pad , \n3123gat_pad , \n3124gat_pad , \n3125gat_pad , \n3126gat_pad , \n3127gat_pad , \n3128gat_pad , \n3130gat_pad , \n3131gat_pad , \n3132gat_pad , \n3133gat_pad , \n3134gat_pad , \n3135gat_pad , \n3136gat_pad , \n3137gat_pad , \n3138gat_pad , \n3140gat_pad , \n3142gat_pad , \n3143gat_pad , \n3144gat_pad , \n3145gat_pad , \n3146gat_pad , \n3147gat_pad , \n3148gat_pad , \n3149gat_pad , \n3150gat_pad , \n3151gat_pad , \n684gat_reg/P0001 , \n824gat_reg/P0001 , \n883gat_reg/P0001 );
	input \n1035gat_reg/NET0131  ;
	input \n1045gat_reg/NET0131  ;
	input \n1068gat_reg/NET0131  ;
	input \n1072gat_reg/NET0131  ;
	input \n1080gat_reg/NET0131  ;
	input \n1121gat_reg/NET0131  ;
	input \n1135gat_reg/NET0131  ;
	input \n1148gat_reg/NET0131  ;
	input \n1197gat_reg/NET0131  ;
	input \n1226gat_reg/NET0131  ;
	input \n1241gat_reg/NET0131  ;
	input \n1282gat_reg/NET0131  ;
	input \n1294gat_reg/NET0131  ;
	input \n1312gat_reg/NET0131  ;
	input \n1316gat_reg/NET0131  ;
	input \n1332gat_reg/NET0131  ;
	input \n1336gat_reg/NET0131  ;
	input \n1340gat_reg/NET0131  ;
	input \n1363gat_reg/NET0131  ;
	input \n1389gat_reg/NET0131  ;
	input \n1394gat_reg/NET0131  ;
	input \n1433gat_reg/NET0131  ;
	input \n1456gat_reg/NET0131  ;
	input \n1462gat_reg/NET0131  ;
	input \n148gat_reg/NET0131  ;
	input \n1496gat_reg/NET0131  ;
	input \n1508gat_reg/NET0131  ;
	input \n1525gat_reg/NET0131  ;
	input \n152gat_reg/NET0131  ;
	input \n156gat_reg/NET0131  ;
	input \n1588gat_reg/NET0131  ;
	input \n1596gat_reg/NET0131  ;
	input \n160gat_reg/NET0131  ;
	input \n1675gat_reg/NET0131  ;
	input \n1678gat_reg/NET0131  ;
	input \n1740gat_reg/NET0131  ;
	input \n1748gat_reg/NET0131  ;
	input \n1763gat_reg/NET0131  ;
	input \n1767gat_reg/NET0131  ;
	input \n1771gat_reg/NET0131  ;
	input \n1775gat_reg/NET0131  ;
	input \n1807gat_reg/NET0131  ;
	input \n1821gat_reg/NET0131  ;
	input \n1829gat_reg/NET0131  ;
	input \n1834gat_reg/NET0131  ;
	input \n1850gat_reg/NET0131  ;
	input \n1871gat_reg/NET0131  ;
	input \n1880gat_reg/NET0131  ;
	input \n1899gat_reg/NET0131  ;
	input \n1975gat_reg/NET0131  ;
	input \n2021gat_reg/NET0131  ;
	input \n2025gat_reg/NET0131  ;
	input \n2029gat_reg/NET0131  ;
	input \n2033gat_reg/NET0131  ;
	input \n2037gat_reg/NET0131  ;
	input \n2040gat_reg/NET0131  ;
	input \n2044gat_reg/NET0131  ;
	input \n2061gat_reg/NET0131  ;
	input \n2084gat_reg/NET0131  ;
	input \n2091gat_reg/NET0131  ;
	input \n2095gat_reg/NET0131  ;
	input \n2099gat_reg/NET0131  ;
	input \n2102gat_reg/NET0131  ;
	input \n2110gat_reg/NET0131  ;
	input \n2117gat_reg/NET0131  ;
	input \n2121gat_reg/NET0131  ;
	input \n2125gat_reg/NET0131  ;
	input \n2135gat_reg/NET0131  ;
	input \n2139gat_reg/NET0131  ;
	input \n2143gat_reg/NET0131  ;
	input \n2155gat_reg/NET0131  ;
	input \n2169gat_reg/NET0131  ;
	input \n2176gat_reg/NET0131  ;
	input \n2179gat_reg/NET0131  ;
	input \n2182gat_reg/NET0131  ;
	input \n2190gat_reg/NET0131  ;
	input \n2203gat_reg/NET0131  ;
	input \n2207gat_reg/NET0131  ;
	input \n2262gat_reg/NET0131  ;
	input \n2266gat_reg/NET0131  ;
	input \n2270gat_reg/NET0131  ;
	input \n2319gat_reg/NET0131  ;
	input \n2339gat_reg/NET0131  ;
	input \n2343gat_reg/NET0131  ;
	input \n2347gat_reg/NET0131  ;
	input \n2390gat_reg/NET0131  ;
	input \n2394gat_reg/NET0131  ;
	input \n2399gat_reg/NET0131  ;
	input \n2403gat_reg/NET0131  ;
	input \n2407gat_reg/NET0131  ;
	input \n2440gat_reg/NET0131  ;
	input \n2446gat_reg/NET0131  ;
	input \n2450gat_reg/NET0131  ;
	input \n2454gat_reg/NET0131  ;
	input \n2458gat_reg/NET0131  ;
	input \n2464gat_reg/NET0131  ;
	input \n2468gat_reg/NET0131  ;
	input \n2472gat_reg/NET0131  ;
	input \n2476gat_reg/NET0131  ;
	input \n2490gat_reg/NET0131  ;
	input \n2495gat_reg/NET0131  ;
	input \n2502gat_reg/NET0131  ;
	input \n2506gat_reg/NET0131  ;
	input \n2510gat_reg/NET0131  ;
	input \n2514gat_reg/NET0131  ;
	input \n2518gat_reg/NET0131  ;
	input \n2526gat_reg/NET0131  ;
	input \n2543gat_reg/NET0131  ;
	input \n2562gat_reg/NET0131  ;
	input \n256gat_reg/NET0131  ;
	input \n2588gat_reg/NET0131  ;
	input \n2592gat_reg/NET0131  ;
	input \n2599gat_reg/NET0131  ;
	input \n2622gat_reg/NET0131  ;
	input \n2626gat_reg/NET0131  ;
	input \n2630gat_reg/NET0131  ;
	input \n2634gat_reg/NET0131  ;
	input \n2640gat_reg/NET0131  ;
	input \n2644gat_reg/NET0131  ;
	input \n2658gat_reg/NET0131  ;
	input \n271gat_reg/NET0131  ;
	input \n3065gat_pad  ;
	input \n3066gat_pad  ;
	input \n3067gat_pad  ;
	input \n3068gat_pad  ;
	input \n3069gat_pad  ;
	input \n3070gat_pad  ;
	input \n3071gat_pad  ;
	input \n3072gat_pad  ;
	input \n3073gat_pad  ;
	input \n3074gat_pad  ;
	input \n3075gat_pad  ;
	input \n3076gat_pad  ;
	input \n3077gat_pad  ;
	input \n3078gat_pad  ;
	input \n3079gat_pad  ;
	input \n3080gat_pad  ;
	input \n3081gat_pad  ;
	input \n3082gat_pad  ;
	input \n3083gat_pad  ;
	input \n3084gat_pad  ;
	input \n3085gat_pad  ;
	input \n3086gat_pad  ;
	input \n3087gat_pad  ;
	input \n3088gat_pad  ;
	input \n3089gat_pad  ;
	input \n3090gat_pad  ;
	input \n3091gat_pad  ;
	input \n3092gat_pad  ;
	input \n3093gat_pad  ;
	input \n3094gat_pad  ;
	input \n3095gat_pad  ;
	input \n3097gat_pad  ;
	input \n3098gat_pad  ;
	input \n3099gat_pad  ;
	input \n3100gat_pad  ;
	input \n314gat_reg/NET0131  ;
	input \n318gat_reg/NET0131  ;
	input \n322gat_reg/NET0131  ;
	input \n327gat_reg/NET0131  ;
	input \n331gat_reg/NET0131  ;
	input \n337gat_reg/NET0131  ;
	input \n341gat_reg/NET0131  ;
	input \n366gat_reg/NET0131  ;
	input \n384gat_reg/NET0131  ;
	input \n388gat_reg/NET0131  ;
	input \n398gat_reg/NET0131  ;
	input \n402gat_reg/NET0131  ;
	input \n463gat_reg/NET0131  ;
	input \n470gat_reg/NET0131  ;
	input \n553gat_reg/NET0131  ;
	input \n561gat_reg/NET0131  ;
	input \n580gat_reg/NET0131  ;
	input \n584gat_reg/NET0131  ;
	input \n614gat_reg/NET0131  ;
	input \n659gat_reg/NET0131  ;
	input \n667gat_reg/NET0131  ;
	input \n673gat_reg/NET0131  ;
	input \n680gat_reg/NET0131  ;
	input \n684gat_reg/NET0131  ;
	input \n699gat_reg/NET0131  ;
	input \n707gat_reg/NET0131  ;
	input \n777gat_reg/NET0131  ;
	input \n816gat_reg/NET0131  ;
	input \n820gat_reg/NET0131  ;
	input \n824gat_reg/NET0131  ;
	input \n830gat_reg/NET0131  ;
	input \n834gat_reg/NET0131  ;
	input \n838gat_reg/NET0131  ;
	input \n842gat_reg/NET0131  ;
	input \n846gat_reg/NET0131  ;
	input \n861gat_reg/NET0131  ;
	input \n865gat_reg/NET0131  ;
	input \n883gat_reg/NET0131  ;
	input \n919gat_reg/NET0131  ;
	input \n931gat_reg/NET0131  ;
	input \n957gat_reg/NET0131  ;
	output \_al_n0  ;
	output \g17_dup/_0_  ;
	output \g6952/_2_  ;
	output \g6953/_2_  ;
	output \g6961/_0_  ;
	output \g7076/_0_  ;
	output \g7077/_0_  ;
	output \g7079/_0_  ;
	output \g7081/_0_  ;
	output \g7082/_0_  ;
	output \g7083/_0_  ;
	output \g7146/_0_  ;
	output \g7147/_0_  ;
	output \g7148/_0_  ;
	output \g7149/_0_  ;
	output \g7150/_0_  ;
	output \g7151/_0_  ;
	output \g7152/_0_  ;
	output \g7153/_0_  ;
	output \g7154/_0_  ;
	output \g7156/_2_  ;
	output \g7161/_2_  ;
	output \g7165/_2_  ;
	output \g7174/_0_  ;
	output \g7180/_00_  ;
	output \g7182/_3_  ;
	output \g7191/_0_  ;
	output \g7204/_0_  ;
	output \g7209/_3_  ;
	output \g7220/_0_  ;
	output \g7229/_0_  ;
	output \g7233/_0_  ;
	output \g7234/_0_  ;
	output \g7235/_0_  ;
	output \g7236/_0_  ;
	output \g7237/_0_  ;
	output \g7238/_0_  ;
	output \g7241/_3_  ;
	output \g7264/_0_  ;
	output \g7265/_0_  ;
	output \g7266/_0_  ;
	output \g7267/_0_  ;
	output \g7268/_0_  ;
	output \g7301/_0_  ;
	output \g7326/_3_  ;
	output \g7350/_2_  ;
	output \g7352/_0_  ;
	output \g7356/_0_  ;
	output \g7359/_0_  ;
	output \g7389/_3_  ;
	output \g7417/_0_  ;
	output \g7418/_0_  ;
	output \g7419/_0_  ;
	output \g7444/_0_  ;
	output \g7445/_0_  ;
	output \g7449/_3_  ;
	output \g7451/_3_  ;
	output \g7454/_0_  ;
	output \g7467/_3_  ;
	output \g7476/_0_  ;
	output \g7480/_0_  ;
	output \g7494/_0_  ;
	output \g7509/_0_  ;
	output \g7514/_0_  ;
	output \g7517/_3_  ;
	output \g7524/_0_  ;
	output \g7558/_0_  ;
	output \g7560/_0_  ;
	output \g7561/_0_  ;
	output \g7563/_0_  ;
	output \g7567/_0_  ;
	output \g7572/_0_  ;
	output \g7579/_0_  ;
	output \g7605/_0_  ;
	output \g7625/_0_  ;
	output \g7627/_0_  ;
	output \g7671/_0_  ;
	output \g7675/_0_  ;
	output \g7689/_0_  ;
	output \g7697/_0_  ;
	output \g7743/_1_  ;
	output \g7764/_1_  ;
	output \g7769/_0_  ;
	output \g7771/_2_  ;
	output \g7779/_0_  ;
	output \g7852/_0_  ;
	output \g7873/_0_  ;
	output \g7884/_3_  ;
	output \g7889/_0_  ;
	output \g7902/_1_  ;
	output \g7992/_3_  ;
	output \g7994/_3_  ;
	output \g7996/_3_  ;
	output \g7998/_3_  ;
	output \g8000/_3_  ;
	output \g8002/_3_  ;
	output \g8004/_3_  ;
	output \g8006/_3_  ;
	output \g8008/_3_  ;
	output \g8150/_0_  ;
	output \g8151/_0_  ;
	output \g8157/_0_  ;
	output \g8163/_0_  ;
	output \g8172/_0_  ;
	output \g8197/_0_  ;
	output \g8211/_0_  ;
	output \g8223/_0_  ;
	output \g8237/_0_  ;
	output \g8251/_0_  ;
	output \g8261/_0_  ;
	output \g8272/_0_  ;
	output \g8287/_0_  ;
	output \g8647/_0_  ;
	output \g8671/_0_  ;
	output \g8672/_0_  ;
	output \g8735/_0_  ;
	output \g8766/_0_  ;
	output \g8811/_0_  ;
	output \g8821/_0_  ;
	output \g8856/_0_  ;
	output \g8858/_3_  ;
	output \g8868/_0_  ;
	output \g8880/_2_  ;
	output \g8886/_0_  ;
	output \g8900/_0_  ;
	output \g8932/_0_  ;
	output \g8991/_3_  ;
	output \g9014/_3_  ;
	output \g9074/_0_  ;
	output \g9091/_0_  ;
	output \g9105/_0_  ;
	output \g9107/_1_  ;
	output \g9111/_0_  ;
	output \n1332gat_reg/P0001  ;
	output \n1363gat_reg/P0001  ;
	output \n1394gat_reg/P0001  ;
	output \n1433gat_reg/P0001  ;
	output \n1775gat_reg/P0001  ;
	output \n2025gat_reg/P0001  ;
	output \n2029gat_reg/P0001  ;
	output \n2033gat_reg/P0001  ;
	output \n2044gat_reg/P0001  ;
	output \n2121gat_reg/P0001  ;
	output \n2125gat_reg/P0001  ;
	output \n2458gat_reg/P0001  ;
	output \n2472gat_reg/P0001  ;
	output \n2592gat_reg/P0001  ;
	output \n3104gat_pad  ;
	output \n3105gat_pad  ;
	output \n3106gat_pad  ;
	output \n3107gat_pad  ;
	output \n3108gat_pad  ;
	output \n3109gat_pad  ;
	output \n3110gat_pad  ;
	output \n3111gat_pad  ;
	output \n3112gat_pad  ;
	output \n3113gat_pad  ;
	output \n3114gat_pad  ;
	output \n3116gat_pad  ;
	output \n3117gat_pad  ;
	output \n3118gat_pad  ;
	output \n3119gat_pad  ;
	output \n3120gat_pad  ;
	output \n3121gat_pad  ;
	output \n3122gat_pad  ;
	output \n3123gat_pad  ;
	output \n3124gat_pad  ;
	output \n3125gat_pad  ;
	output \n3126gat_pad  ;
	output \n3127gat_pad  ;
	output \n3128gat_pad  ;
	output \n3130gat_pad  ;
	output \n3131gat_pad  ;
	output \n3132gat_pad  ;
	output \n3133gat_pad  ;
	output \n3134gat_pad  ;
	output \n3135gat_pad  ;
	output \n3136gat_pad  ;
	output \n3137gat_pad  ;
	output \n3138gat_pad  ;
	output \n3140gat_pad  ;
	output \n3142gat_pad  ;
	output \n3143gat_pad  ;
	output \n3144gat_pad  ;
	output \n3145gat_pad  ;
	output \n3146gat_pad  ;
	output \n3147gat_pad  ;
	output \n3148gat_pad  ;
	output \n3149gat_pad  ;
	output \n3150gat_pad  ;
	output \n3151gat_pad  ;
	output \n684gat_reg/P0001  ;
	output \n824gat_reg/P0001  ;
	output \n883gat_reg/P0001  ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\n2454gat_reg/NET0131 ,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\n846gat_reg/NET0131 ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\n3088gat_pad ,
		\n3095gat_pad ,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\n3087gat_pad ,
		\n3093gat_pad ,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\n3087gat_pad ,
		\n3095gat_pad ,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\n3086gat_pad ,
		\n3093gat_pad ,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		_w203_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\n3086gat_pad ,
		\n3095gat_pad ,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\n3085gat_pad ,
		\n3093gat_pad ,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w208_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\n673gat_reg/NET0131 ,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w207_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		_w207_,
		_w210_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\n659gat_reg/NET0131 ,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\n659gat_reg/NET0131 ,
		_w216_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\n553gat_reg/NET0131 ,
		\n777gat_reg/NET0131 ,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\n553gat_reg/NET0131 ,
		\n777gat_reg/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w220_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\n314gat_reg/NET0131 ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\n314gat_reg/NET0131 ,
		_w222_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\n366gat_reg/NET0131 ,
		\n561gat_reg/NET0131 ,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\n366gat_reg/NET0131 ,
		\n561gat_reg/NET0131 ,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		_w225_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w225_,
		_w228_,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w229_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w219_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w219_,
		_w231_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w213_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\n820gat_reg/NET0131 ,
		_w203_,
		_w236_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		_w206_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w203_,
		_w206_,
		_w238_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\n842gat_reg/NET0131 ,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w237_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w210_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w210_,
		_w238_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		\n1241gat_reg/NET0131 ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w212_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w241_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w235_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\n3083gat_pad ,
		\n3084gat_pad ,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\n3093gat_pad ,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w247_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		\n3088gat_pad ,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\n3085gat_pad ,
		_w248_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\n3095gat_pad ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\n3086gat_pad ,
		\n3087gat_pad ,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w201_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w253_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w251_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w246_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\n3086gat_pad ,
		\n3087gat_pad ,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\n3095gat_pad ,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w253_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w209_,
		_w254_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\n3088gat_pad ,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w250_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w261_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\n1045gat_reg/NET0131 ,
		\n1072gat_reg/NET0131 ,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		\n1045gat_reg/NET0131 ,
		\n1072gat_reg/NET0131 ,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\n1035gat_reg/NET0131 ,
		\n1121gat_reg/NET0131 ,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\n1035gat_reg/NET0131 ,
		\n1121gat_reg/NET0131 ,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\n1282gat_reg/NET0131 ,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\n1282gat_reg/NET0131 ,
		_w271_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\n1135gat_reg/NET0131 ,
		\n931gat_reg/NET0131 ,
		_w275_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\n1135gat_reg/NET0131 ,
		\n931gat_reg/NET0131 ,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\n1226gat_reg/NET0131 ,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\n1226gat_reg/NET0131 ,
		_w277_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		_w274_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w274_,
		_w280_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w268_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w268_,
		_w283_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w213_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w203_,
		_w206_,
		_w288_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w210_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\n830gat_reg/NET0131 ,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		\n842gat_reg/NET0131 ,
		_w242_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w287_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w265_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w258_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\n2464gat_reg/NET0131 ,
		\n2468gat_reg/NET0131 ,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\n2476gat_reg/NET0131 ,
		\n2518gat_reg/NET0131 ,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\n2526gat_reg/NET0131 ,
		\n2599gat_reg/NET0131 ,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\n3090gat_pad ,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w296_,
		_w297_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\n667gat_reg/NET0131 ,
		_w234_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\n667gat_reg/NET0131 ,
		_w234_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\n3069gat_pad ,
		\n3093gat_pad ,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\n3078gat_pad ,
		\n3095gat_pad ,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		\n2562gat_reg/NET0131 ,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w308_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\n2490gat_reg/NET0131 ,
		\n2543gat_reg/NET0131 ,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\n2630gat_reg/NET0131 ,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\n2155gat_reg/NET0131 ,
		\n2622gat_reg/NET0131 ,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		\n2626gat_reg/NET0131 ,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w313_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\n2543gat_reg/NET0131 ,
		\n2630gat_reg/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		\n2622gat_reg/NET0131 ,
		\n2626gat_reg/NET0131 ,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\n2155gat_reg/NET0131 ,
		\n2490gat_reg/NET0131 ,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w317_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w318_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w316_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\n2454gat_reg/NET0131 ,
		_w323_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w327_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		\n2454gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		\n919gat_reg/NET0131 ,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w327_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w200_,
		_w326_,
		_w331_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\n2562gat_reg/NET0131 ,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w308_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\n2207gat_reg/NET0131 ,
		_w311_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w335_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w322_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		_w332_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		_w307_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\n3070gat_pad ,
		\n3093gat_pad ,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\n3079gat_pad ,
		\n3095gat_pad ,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w341_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		_w339_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\n3072gat_pad ,
		\n3093gat_pad ,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\n3081gat_pad ,
		\n3095gat_pad ,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w345_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w339_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\n3071gat_pad ,
		\n3093gat_pad ,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\n3080gat_pad ,
		\n3095gat_pad ,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w349_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w339_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\n3065gat_pad ,
		\n3093gat_pad ,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\n3074gat_pad ,
		\n3095gat_pad ,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w353_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w339_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\n3073gat_pad ,
		\n3093gat_pad ,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\n3082gat_pad ,
		\n3095gat_pad ,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w357_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w339_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\n1871gat_reg/NET0131 ,
		_w252_,
		_w361_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w204_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\n3094gat_pad ,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		_w208_,
		_w361_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		\n3088gat_pad ,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w363_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\n1871gat_reg/NET0131 ,
		_w249_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\n3088gat_pad ,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\n3087gat_pad ,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\n3091gat_pad ,
		\n3092gat_pad ,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\n3085gat_pad ,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\n3086gat_pad ,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w369_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w366_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		\n3068gat_pad ,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w339_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name179 (
		\n3065gat_pad ,
		_w374_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w339_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\n3069gat_pad ,
		_w374_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w339_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		\n3066gat_pad ,
		_w374_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w339_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\n3067gat_pad ,
		_w374_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w339_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		\n3070gat_pad ,
		_w374_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w339_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\n3073gat_pad ,
		_w374_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w339_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\n3072gat_pad ,
		_w374_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w339_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\n3071gat_pad ,
		_w374_,
		_w391_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w339_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		\n1312gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		_w393_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\n1880gat_reg/NET0131 ,
		\n2021gat_reg/NET0131 ,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\n1880gat_reg/NET0131 ,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		\n2347gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		\n2407gat_reg/NET0131 ,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\n2403gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\n2403gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w400_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h2)
	) name205 (
		\n2347gat_reg/NET0131 ,
		\n2407gat_reg/NET0131 ,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\n398gat_reg/NET0131 ,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w402_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		_w324_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w399_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w397_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w409_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w412_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\n846gat_reg/NET0131 ,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name217 (
		\n846gat_reg/NET0131 ,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		\n919gat_reg/NET0131 ,
		_w413_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		_w415_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w411_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		_w405_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w408_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		\n2102gat_reg/NET0131 ,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\n1850gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		\n2139gat_reg/NET0131 ,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w423_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w422_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w428_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		\n2061gat_reg/NET0131 ,
		_w422_,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		\n1850gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w428_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w429_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w427_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w396_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		_w420_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w394_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		\n2502gat_reg/NET0131 ,
		\n2506gat_reg/NET0131 ,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		\n2510gat_reg/NET0131 ,
		\n2588gat_reg/NET0131 ,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		\n2658gat_reg/NET0131 ,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w437_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\n3100gat_pad ,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w393_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w436_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w399_,
		_w410_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w432_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		_w435_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\n2622gat_reg/NET0131 ,
		\n2626gat_reg/NET0131 ,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w318_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\n2543gat_reg/NET0131 ,
		\n2630gat_reg/NET0131 ,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w317_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		\n2490gat_reg/NET0131 ,
		\n2634gat_reg/NET0131 ,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\n2490gat_reg/NET0131 ,
		\n2634gat_reg/NET0131 ,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w451_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w450_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w450_,
		_w453_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w454_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w448_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w448_,
		_w456_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w457_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		_w426_,
		_w435_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w461_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		\n2135gat_reg/NET0131 ,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		\n2179gat_reg/NET0131 ,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		\n2182gat_reg/NET0131 ,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		\n2143gat_reg/NET0131 ,
		_w425_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\n1850gat_reg/NET0131 ,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\n1740gat_reg/NET0131 ,
		_w422_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h4)
	) name271 (
		\n1740gat_reg/NET0131 ,
		_w432_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		\n1496gat_reg/NET0131 ,
		\n2091gat_reg/NET0131 ,
		_w470_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		_w427_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h4)
	) name274 (
		\n2061gat_reg/NET0131 ,
		_w423_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w428_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w422_,
		_w470_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w468_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w469_,
		_w471_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w476_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w410_,
		_w422_,
		_w479_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w414_,
		_w422_,
		_w480_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		_w399_,
		_w479_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w480_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h4)
	) name285 (
		_w464_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w478_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\n2562gat_reg/NET0131 ,
		_w309_,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w313_,
		_w447_,
		_w486_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w487_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w485_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w486_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		\n2135gat_reg/NET0131 ,
		_w461_,
		_w490_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w462_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		\n2099gat_reg/NET0131 ,
		_w394_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		\n2037gat_reg/NET0131 ,
		\n2095gat_reg/NET0131 ,
		_w493_
	);
	LUT2 #(
		.INIT('h4)
	) name296 (
		_w492_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w441_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		_w491_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w497_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\n2266gat_reg/NET0131 ,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		\n2266gat_reg/NET0131 ,
		_w497_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w495_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		\n699gat_reg/NET0131 ,
		\n824gat_reg/NET0131 ,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		\n699gat_reg/NET0131 ,
		\n824gat_reg/NET0131 ,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		\n680gat_reg/NET0131 ,
		\n883gat_reg/NET0131 ,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		\n680gat_reg/NET0131 ,
		\n883gat_reg/NET0131 ,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w505_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		_w504_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		_w504_,
		_w507_,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w508_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		\n580gat_reg/NET0131 ,
		\n820gat_reg/NET0131 ,
		_w511_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\n580gat_reg/NET0131 ,
		\n820gat_reg/NET0131 ,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w511_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		\n584gat_reg/NET0131 ,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		\n584gat_reg/NET0131 ,
		_w513_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		\n684gat_reg/NET0131 ,
		\n816gat_reg/NET0131 ,
		_w517_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		\n684gat_reg/NET0131 ,
		\n816gat_reg/NET0131 ,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w517_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		_w516_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		_w516_,
		_w519_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w520_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w510_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w510_,
		_w522_,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w523_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		\n2390gat_reg/NET0131 ,
		\n2495gat_reg/NET0131 ,
		_w526_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\n2390gat_reg/NET0131 ,
		\n2495gat_reg/NET0131 ,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w526_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		\n2270gat_reg/NET0131 ,
		\n2339gat_reg/NET0131 ,
		_w529_
	);
	LUT2 #(
		.INIT('h4)
	) name332 (
		\n2270gat_reg/NET0131 ,
		\n2339gat_reg/NET0131 ,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w529_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w528_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w528_,
		_w531_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w532_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		_w495_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w478_,
		_w495_,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w537_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h2)
	) name342 (
		\n2143gat_reg/NET0131 ,
		_w425_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w465_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		_w538_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		\n2061gat_reg/NET0131 ,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\n2061gat_reg/NET0131 ,
		_w543_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w544_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		_w538_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		\n1850gat_reg/NET0131 ,
		_w465_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w466_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w538_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w424_,
		_w428_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w465_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		\n1975gat_reg/NET0131 ,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h2)
	) name356 (
		\n1975gat_reg/NET0131 ,
		_w552_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w553_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		_w538_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\n614gat_reg/NET0131 ,
		\n838gat_reg/NET0131 ,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		\n614gat_reg/NET0131 ,
		\n838gat_reg/NET0131 ,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w324_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w198_,
		_w323_,
		_w562_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w561_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w561_,
		_w562_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w563_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		\n707gat_reg/NET0131 ,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		\n707gat_reg/NET0131 ,
		_w565_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w566_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		\n830gat_reg/NET0131 ,
		\n834gat_reg/NET0131 ,
		_w569_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		\n830gat_reg/NET0131 ,
		\n834gat_reg/NET0131 ,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		_w568_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		_w568_,
		_w571_,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w572_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		_w559_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		_w559_,
		_w574_,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w482_,
		_w495_,
		_w578_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		\n2403gat_reg/NET0131 ,
		_w412_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		\n2347gat_reg/NET0131 ,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		\n2347gat_reg/NET0131 ,
		_w579_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		_w578_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		\n2347gat_reg/NET0131 ,
		\n2407gat_reg/NET0131 ,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w403_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w580_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w580_,
		_w585_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		_w578_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		\n2347gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name393 (
		\n2440gat_reg/NET0131 ,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w414_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		\n2644gat_reg/NET0131 ,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\n2644gat_reg/NET0131 ,
		_w592_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w578_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		\n2403gat_reg/NET0131 ,
		_w412_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w579_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w578_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w397_,
		_w578_,
		_w600_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		\n2403gat_reg/NET0131 ,
		_w584_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		_w410_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w433_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		\n1850gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w428_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w429_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		\n2454gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w327_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		_w332_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		\n1316gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		_w610_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		\n2040gat_reg/NET0131 ,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		\n1294gat_reg/NET0131 ,
		\n673gat_reg/NET0131 ,
		_w612_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		\n1294gat_reg/NET0131 ,
		\n673gat_reg/NET0131 ,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w612_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		\n1068gat_reg/NET0131 ,
		\n861gat_reg/NET0131 ,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		\n1068gat_reg/NET0131 ,
		\n861gat_reg/NET0131 ,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w615_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h2)
	) name420 (
		_w614_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w614_,
		_w617_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		\n1148gat_reg/NET0131 ,
		\n865gat_reg/NET0131 ,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\n1148gat_reg/NET0131 ,
		\n865gat_reg/NET0131 ,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w621_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\n1080gat_reg/NET0131 ,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\n1080gat_reg/NET0131 ,
		_w623_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w624_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		\n1241gat_reg/NET0131 ,
		\n957gat_reg/NET0131 ,
		_w627_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		\n1241gat_reg/NET0131 ,
		\n957gat_reg/NET0131 ,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w627_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		_w626_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name433 (
		_w626_,
		_w629_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w630_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		_w620_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w620_,
		_w632_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name438 (
		_w199_,
		_w409_,
		_w636_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		\n1821gat_reg/NET0131 ,
		\n1829gat_reg/NET0131 ,
		_w637_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\n2446gat_reg/NET0131 ,
		\n2450gat_reg/NET0131 ,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\n3100gat_pad ,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		\n2472gat_reg/NET0131 ,
		_w637_,
		_w640_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w636_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		\n2454gat_reg/NET0131 ,
		\n271gat_reg/NET0131 ,
		_w643_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		_w641_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w199_,
		_w560_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w641_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		\n3094gat_pad ,
		_w362_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\n3088gat_pad ,
		_w364_,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w647_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		\n3080gat_pad ,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		\n3088gat_pad ,
		_w367_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		\n3086gat_pad ,
		_w371_,
		_w652_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		\n3087gat_pad ,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w651_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		\n3071gat_pad ,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w649_,
		_w654_,
		_w656_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w199_,
		_w324_,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		\n388gat_reg/NET0131 ,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		\n331gat_reg/NET0131 ,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		\n331gat_reg/NET0131 ,
		_w658_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w659_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w656_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w650_,
		_w655_,
		_w663_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w662_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w368_,
		_w653_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w649_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		_w198_,
		_w329_,
		_w667_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		\n156gat_reg/NET0131 ,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		\n152gat_reg/NET0131 ,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		\n256gat_reg/NET0131 ,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		\n148gat_reg/NET0131 ,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		\n148gat_reg/NET0131 ,
		_w670_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w671_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h2)
	) name476 (
		_w666_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		\n3065gat_pad ,
		_w666_,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w674_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		\n152gat_reg/NET0131 ,
		\n256gat_reg/NET0131 ,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		\n156gat_reg/NET0131 ,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		_w667_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		\n470gat_reg/NET0131 ,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		\n470gat_reg/NET0131 ,
		_w679_,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w680_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h2)
	) name485 (
		_w666_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		\n3073gat_pad ,
		_w666_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w683_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		\n3083gat_pad ,
		\n3088gat_pad ,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\n3083gat_pad ,
		\n3088gat_pad ,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w686_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		\n3084gat_pad ,
		\n3085gat_pad ,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		\n3084gat_pad ,
		\n3085gat_pad ,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		\n3089gat_pad ,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		\n3089gat_pad ,
		_w691_,
		_w693_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w692_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w254_,
		_w259_,
		_w695_
	);
	LUT2 #(
		.INIT('h2)
	) name498 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		_w694_,
		_w695_,
		_w697_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w696_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w688_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w688_,
		_w698_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w699_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		\n256gat_reg/NET0131 ,
		_w669_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w670_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		_w666_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h2)
	) name507 (
		\n3066gat_pad ,
		_w666_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w704_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		\n3079gat_pad ,
		_w649_,
		_w707_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\n3070gat_pad ,
		_w654_,
		_w708_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\n327gat_reg/NET0131 ,
		_w659_,
		_w709_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		\n327gat_reg/NET0131 ,
		_w659_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		_w709_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		_w656_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w707_,
		_w708_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		\n152gat_reg/NET0131 ,
		_w668_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w669_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		_w666_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		\n3067gat_pad ,
		_w666_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w717_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w326_,
		_w608_,
		_w720_
	);
	LUT2 #(
		.INIT('h4)
	) name523 (
		_w330_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w199_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\n156gat_reg/NET0131 ,
		_w667_,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w668_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		_w666_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h2)
	) name528 (
		\n3068gat_pad ,
		_w666_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w725_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h8)
	) name530 (
		\n3067gat_pad ,
		_w654_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		\n3076gat_pad ,
		_w649_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w728_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		\n3068gat_pad ,
		_w654_,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		\n3077gat_pad ,
		_w649_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w731_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name536 (
		\n3065gat_pad ,
		_w654_,
		_w734_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		\n3074gat_pad ,
		_w649_,
		_w735_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w734_,
		_w735_,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		\n3066gat_pad ,
		_w654_,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		\n3075gat_pad ,
		_w649_,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w737_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		\n2562gat_reg/NET0131 ,
		\n2640gat_reg/NET0131 ,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		\n2562gat_reg/NET0131 ,
		\n2640gat_reg/NET0131 ,
		_w741_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w740_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name545 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		_w743_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w333_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w745_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w308_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		_w744_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		_w744_,
		_w746_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w747_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w742_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w742_,
		_w749_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h2)
	) name555 (
		\n2117gat_reg/NET0131 ,
		\n2125gat_reg/NET0131 ,
		_w753_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w639_,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		_w363_,
		_w648_,
		_w755_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		\n3087gat_pad ,
		_w372_,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w651_,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w755_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		\n2319gat_reg/NET0131 ,
		\n3099gat_pad ,
		_w759_
	);
	LUT2 #(
		.INIT('h8)
	) name562 (
		_w414_,
		_w601_,
		_w760_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		_w466_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name564 (
		\n2061gat_reg/NET0131 ,
		_w423_,
		_w762_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		_w428_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name566 (
		\n2403gat_reg/NET0131 ,
		_w397_,
		_w764_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w403_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w763_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		_w426_,
		_w760_,
		_w767_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		_w472_,
		_w537_,
		_w768_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		_w602_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		_w423_,
		_w544_,
		_w770_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w602_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		\n1312gat_reg/NET0131 ,
		_w763_,
		_w772_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w773_
	);
	LUT2 #(
		.INIT('h8)
	) name576 (
		_w762_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		_w324_,
		_w327_,
		_w775_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		\n3066gat_pad ,
		\n3093gat_pad ,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name579 (
		\n3075gat_pad ,
		\n3095gat_pad ,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w776_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		\n3068gat_pad ,
		\n3093gat_pad ,
		_w779_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\n3077gat_pad ,
		\n3095gat_pad ,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w779_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\n3067gat_pad ,
		\n3093gat_pad ,
		_w782_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\n3076gat_pad ,
		\n3095gat_pad ,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w782_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		\n337gat_reg/NET0131 ,
		\n341gat_reg/NET0131 ,
		_w785_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		\n337gat_reg/NET0131 ,
		\n341gat_reg/NET0131 ,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\n160gat_reg/NET0131 ,
		_w565_,
		_w788_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		\n160gat_reg/NET0131 ,
		_w565_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		\n271gat_reg/NET0131 ,
		\n842gat_reg/NET0131 ,
		_w791_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\n271gat_reg/NET0131 ,
		\n842gat_reg/NET0131 ,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w791_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		_w790_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		_w790_,
		_w793_,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		_w794_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w787_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w787_,
		_w796_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		_w797_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		_w339_,
		_w784_,
		_w800_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		_w339_,
		_w781_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		\n3078gat_pad ,
		_w649_,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		\n3069gat_pad ,
		_w654_,
		_w803_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		\n384gat_reg/NET0131 ,
		_w710_,
		_w804_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		\n384gat_reg/NET0131 ,
		_w710_,
		_w805_
	);
	LUT2 #(
		.INIT('h2)
	) name608 (
		_w656_,
		_w804_,
		_w806_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w805_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		_w802_,
		_w803_,
		_w808_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		_w807_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		\n3082gat_pad ,
		_w649_,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name613 (
		\n3073gat_pad ,
		_w654_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name614 (
		\n327gat_reg/NET0131 ,
		\n331gat_reg/NET0131 ,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		\n388gat_reg/NET0131 ,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		_w657_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		\n463gat_reg/NET0131 ,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h2)
	) name618 (
		\n463gat_reg/NET0131 ,
		_w814_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w815_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w656_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w810_,
		_w811_,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h4)
	) name623 (
		_w339_,
		_w778_,
		_w821_
	);
	LUT2 #(
		.INIT('h8)
	) name624 (
		\n3081gat_pad ,
		_w649_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		\n3072gat_pad ,
		_w654_,
		_w823_
	);
	LUT2 #(
		.INIT('h2)
	) name626 (
		\n388gat_reg/NET0131 ,
		_w657_,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		_w658_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h8)
	) name628 (
		_w656_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w822_,
		_w823_,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		_w826_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		\n1312gat_reg/NET0131 ,
		\n2169gat_reg/NET0131 ,
		_w829_
	);
	LUT2 #(
		.INIT('h4)
	) name632 (
		_w441_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		_w435_,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		\n1197gat_reg/NET0131 ,
		_w286_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		\n1197gat_reg/NET0131 ,
		_w286_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w832_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		\n3086gat_pad ,
		_w201_,
		_w835_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		_w363_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		_w837_
	);
	LUT2 #(
		.INIT('h8)
	) name640 (
		_w369_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		_w370_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		_w549_,
		_w836_,
		_w840_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		_w839_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		_w365_,
		_w647_,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		_w369_,
		_w652_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		_w541_,
		_w842_,
		_w844_
	);
	LUT2 #(
		.INIT('h4)
	) name647 (
		_w843_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		\n1771gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		_w846_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		\n1871gat_reg/NET0131 ,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		\n1035gat_reg/NET0131 ,
		_w588_,
		_w848_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		\n1072gat_reg/NET0131 ,
		_w582_,
		_w849_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		\n1121gat_reg/NET0131 ,
		_w598_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		\n931gat_reg/NET0131 ,
		_w397_,
		_w851_
	);
	LUT2 #(
		.INIT('h2)
	) name654 (
		\n1135gat_reg/NET0131 ,
		_w491_,
		_w852_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		\n1282gat_reg/NET0131 ,
		_w535_,
		_w853_
	);
	LUT2 #(
		.INIT('h4)
	) name656 (
		\n659gat_reg/NET0131 ,
		_w213_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name657 (
		\n1068gat_reg/NET0131 ,
		_w242_,
		_w855_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w210_,
		_w238_,
		_w856_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		\n271gat_reg/NET0131 ,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h4)
	) name660 (
		\n680gat_reg/NET0131 ,
		_w289_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w854_,
		_w855_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w857_,
		_w858_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name663 (
		_w859_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w261_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h2)
	) name665 (
		_w701_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		\n580gat_reg/NET0131 ,
		_w289_,
		_w864_
	);
	LUT2 #(
		.INIT('h4)
	) name667 (
		\n337gat_reg/NET0131 ,
		_w856_,
		_w865_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		\n777gat_reg/NET0131 ,
		_w213_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		\n861gat_reg/NET0131 ,
		_w242_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w864_,
		_w865_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w866_,
		_w867_,
		_w869_
	);
	LUT2 #(
		.INIT('h8)
	) name672 (
		_w868_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h2)
	) name673 (
		_w261_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		_w799_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		\n816gat_reg/NET0131 ,
		_w289_,
		_w873_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		\n160gat_reg/NET0131 ,
		_w856_,
		_w874_
	);
	LUT2 #(
		.INIT('h4)
	) name677 (
		\n553gat_reg/NET0131 ,
		_w213_,
		_w875_
	);
	LUT2 #(
		.INIT('h4)
	) name678 (
		\n957gat_reg/NET0131 ,
		_w242_,
		_w876_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w873_,
		_w874_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		_w875_,
		_w876_,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		_w877_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h2)
	) name682 (
		_w261_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		_w635_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h4)
	) name684 (
		\n322gat_reg/NET0131 ,
		_w213_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name685 (
		\n865gat_reg/NET0131 ,
		_w242_,
		_w883_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		\n341gat_reg/NET0131 ,
		_w856_,
		_w884_
	);
	LUT2 #(
		.INIT('h4)
	) name687 (
		\n584gat_reg/NET0131 ,
		_w289_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		_w882_,
		_w883_,
		_w886_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w884_,
		_w885_,
		_w887_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w886_,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		_w261_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h2)
	) name692 (
		_w799_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h4)
	) name693 (
		\n699gat_reg/NET0131 ,
		_w289_,
		_w891_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		\n398gat_reg/NET0131 ,
		_w856_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		\n314gat_reg/NET0131 ,
		_w213_,
		_w893_
	);
	LUT2 #(
		.INIT('h4)
	) name696 (
		\n1148gat_reg/NET0131 ,
		_w242_,
		_w894_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w891_,
		_w892_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w893_,
		_w894_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		_w261_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h2)
	) name701 (
		_w525_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		\n684gat_reg/NET0131 ,
		_w289_,
		_w900_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		\n402gat_reg/NET0131 ,
		_w856_,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name704 (
		\n318gat_reg/NET0131 ,
		_w213_,
		_w902_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		\n1080gat_reg/NET0131 ,
		_w242_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		_w900_,
		_w901_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w902_,
		_w903_,
		_w905_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w904_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		_w261_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h2)
	) name710 (
		_w577_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		\n561gat_reg/NET0131 ,
		_w213_,
		_w909_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		\n1294gat_reg/NET0131 ,
		_w242_,
		_w910_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		\n846gat_reg/NET0131 ,
		_w856_,
		_w911_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		\n824gat_reg/NET0131 ,
		_w289_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w909_,
		_w910_,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		_w911_,
		_w912_,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		_w913_,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		_w261_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		_w304_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		\n883gat_reg/NET0131 ,
		_w289_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name721 (
		\n366gat_reg/NET0131 ,
		_w213_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		\n919gat_reg/NET0131 ,
		_w203_,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w210_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		_w206_,
		_w211_,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w921_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w918_,
		_w919_,
		_w924_
	);
	LUT2 #(
		.INIT('h4)
	) name727 (
		_w923_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		_w261_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		_w834_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h4)
	) name730 (
		_w246_,
		_w261_,
		_w928_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		_w534_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w257_,
		_w861_,
		_w930_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		\n1035gat_reg/NET0131 ,
		_w213_,
		_w931_
	);
	LUT2 #(
		.INIT('h4)
	) name734 (
		\n834gat_reg/NET0131 ,
		_w289_,
		_w932_
	);
	LUT2 #(
		.INIT('h4)
	) name735 (
		\n271gat_reg/NET0131 ,
		_w242_,
		_w933_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w931_,
		_w932_,
		_w934_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		_w933_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		_w265_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w930_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		_w257_,
		_w870_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name741 (
		\n838gat_reg/NET0131 ,
		_w289_,
		_w939_
	);
	LUT2 #(
		.INIT('h4)
	) name742 (
		\n1072gat_reg/NET0131 ,
		_w213_,
		_w940_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		\n337gat_reg/NET0131 ,
		_w242_,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w939_,
		_w940_,
		_w942_
	);
	LUT2 #(
		.INIT('h4)
	) name745 (
		_w941_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		_w265_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w938_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w257_,
		_w879_,
		_w946_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		\n707gat_reg/NET0131 ,
		_w289_,
		_w947_
	);
	LUT2 #(
		.INIT('h4)
	) name750 (
		\n1121gat_reg/NET0131 ,
		_w213_,
		_w948_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		\n160gat_reg/NET0131 ,
		_w242_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w947_,
		_w948_,
		_w950_
	);
	LUT2 #(
		.INIT('h4)
	) name753 (
		_w949_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w265_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w946_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		_w257_,
		_w888_,
		_w954_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		\n614gat_reg/NET0131 ,
		_w289_,
		_w955_
	);
	LUT2 #(
		.INIT('h4)
	) name758 (
		\n931gat_reg/NET0131 ,
		_w213_,
		_w956_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		\n341gat_reg/NET0131 ,
		_w242_,
		_w957_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w955_,
		_w956_,
		_w958_
	);
	LUT2 #(
		.INIT('h4)
	) name761 (
		_w957_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w265_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w954_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		\n1045gat_reg/NET0131 ,
		_w213_,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w242_,
		_w289_,
		_w963_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		\n398gat_reg/NET0131 ,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w962_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w265_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w257_,
		_w897_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w966_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		\n1135gat_reg/NET0131 ,
		_w213_,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		\n402gat_reg/NET0131 ,
		_w963_,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w969_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w265_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w257_,
		_w906_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w972_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		\n1282gat_reg/NET0131 ,
		_w213_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		\n846gat_reg/NET0131 ,
		_w963_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		_w975_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w265_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w257_,
		_w915_,
		_w979_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w978_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		\n1226gat_reg/NET0131 ,
		_w213_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		\n919gat_reg/NET0131 ,
		_w963_,
		_w982_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w981_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		_w265_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		_w257_,
		_w925_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		_w984_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		_w200_,
		_w311_,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		_w486_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		\n1340gat_reg/NET0131 ,
		_w609_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w335_,
		_w422_,
		_w990_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w989_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		\n1462gat_reg/NET0131 ,
		_w422_,
		_w992_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		\n1394gat_reg/NET0131 ,
		_w396_,
		_w993_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		_w992_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w991_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		\n1508gat_reg/NET0131 ,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		\n1829gat_reg/NET0131 ,
		\n3097gat_pad ,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		_w394_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h2)
	) name801 (
		\n1821gat_reg/NET0131 ,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		\n1775gat_reg/NET0131 ,
		\n1871gat_reg/NET0131 ,
		_w1000_
	);
	LUT2 #(
		.INIT('h4)
	) name803 (
		\n3098gat_pad ,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		_w999_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		\n1394gat_reg/NET0131 ,
		_w608_,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		\n1596gat_reg/NET0131 ,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		_w422_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		\n1678gat_reg/NET0131 ,
		_w992_,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name809 (
		_w1005_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h4)
	) name810 (
		\n1394gat_reg/NET0131 ,
		_w422_,
		_w1008_
	);
	LUT2 #(
		.INIT('h4)
	) name811 (
		_w332_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		\n1525gat_reg/NET0131 ,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		\n1588gat_reg/NET0131 ,
		\n1596gat_reg/NET0131 ,
		_w1011_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		_w422_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w1002_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h4)
	) name816 (
		_w1007_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		_w1010_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		_w996_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		\n1340gat_reg/NET0131 ,
		\n1807gat_reg/NET0131 ,
		_w1017_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		_w396_,
		_w989_,
		_w1018_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		\n1456gat_reg/NET0131 ,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w1017_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w422_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		\n1675gat_reg/NET0131 ,
		_w1009_,
		_w1022_
	);
	LUT2 #(
		.INIT('h2)
	) name825 (
		\n1336gat_reg/NET0131 ,
		_w332_,
		_w1023_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		_w396_,
		_w608_,
		_w1024_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h4)
	) name828 (
		\n1748gat_reg/NET0131 ,
		_w422_,
		_w1026_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		_w1025_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w1022_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name831 (
		_w1021_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		\n1080gat_reg/NET0131 ,
		_w396_,
		_w1030_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\n684gat_reg/NET0131 ,
		_w396_,
		_w1031_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		_w1032_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		\n2562gat_reg/NET0131 ,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h8)
	) name836 (
		_w745_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		_w1030_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h4)
	) name838 (
		_w1031_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		\n1148gat_reg/NET0131 ,
		_w396_,
		_w1037_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		\n699gat_reg/NET0131 ,
		_w396_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		\n2562gat_reg/NET0131 ,
		_w1032_,
		_w1039_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		_w745_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		_w1037_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h4)
	) name844 (
		_w1038_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		_w310_,
		_w720_,
		_w1043_
	);
	LUT2 #(
		.INIT('h2)
	) name846 (
		\n2084gat_reg/NET0131 ,
		_w326_,
		_w1044_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w485_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		\n2562gat_reg/NET0131 ,
		_w743_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		\n816gat_reg/NET0131 ,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h4)
	) name850 (
		\n680gat_reg/NET0131 ,
		_w334_,
		_w1048_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		\n2562gat_reg/NET0131 ,
		_w743_,
		_w1049_
	);
	LUT2 #(
		.INIT('h4)
	) name852 (
		\n584gat_reg/NET0131 ,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h4)
	) name853 (
		\n2562gat_reg/NET0131 ,
		_w333_,
		_w1051_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		\n580gat_reg/NET0131 ,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		_w1047_,
		_w1048_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w1050_,
		_w1052_,
		_w1054_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		_w1053_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w396_,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h4)
	) name859 (
		\n1068gat_reg/NET0131 ,
		_w334_,
		_w1057_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		\n865gat_reg/NET0131 ,
		_w1049_,
		_w1058_
	);
	LUT2 #(
		.INIT('h4)
	) name861 (
		\n861gat_reg/NET0131 ,
		_w1051_,
		_w1059_
	);
	LUT2 #(
		.INIT('h4)
	) name862 (
		\n957gat_reg/NET0131 ,
		_w1046_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name863 (
		_w1057_,
		_w1058_,
		_w1061_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w1059_,
		_w1060_,
		_w1062_
	);
	LUT2 #(
		.INIT('h8)
	) name865 (
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		_w396_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		_w1043_,
		_w1045_,
		_w1065_
	);
	LUT2 #(
		.INIT('h4)
	) name868 (
		_w1056_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w1064_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h2)
	) name870 (
		_w745_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h8)
	) name871 (
		\n824gat_reg/NET0131 ,
		_w396_,
		_w1069_
	);
	LUT2 #(
		.INIT('h2)
	) name872 (
		\n1294gat_reg/NET0131 ,
		_w396_,
		_w1070_
	);
	LUT2 #(
		.INIT('h2)
	) name873 (
		_w485_,
		_w1069_,
		_w1071_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		_w1070_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		\n883gat_reg/NET0131 ,
		_w396_,
		_w1073_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		\n673gat_reg/NET0131 ,
		_w396_,
		_w1074_
	);
	LUT2 #(
		.INIT('h2)
	) name877 (
		_w310_,
		_w1073_,
		_w1075_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		_w1074_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		\n337gat_reg/NET0131 ,
		_w1051_,
		_w1077_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		\n271gat_reg/NET0131 ,
		_w334_,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name881 (
		\n341gat_reg/NET0131 ,
		_w1049_,
		_w1079_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		\n160gat_reg/NET0131 ,
		_w1046_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w396_,
		_w1077_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1078_,
		_w1079_,
		_w1082_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		_w1080_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name886 (
		_w1081_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		\n614gat_reg/NET0131 ,
		_w1049_,
		_w1085_
	);
	LUT2 #(
		.INIT('h4)
	) name888 (
		\n834gat_reg/NET0131 ,
		_w334_,
		_w1086_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		\n707gat_reg/NET0131 ,
		_w1046_,
		_w1087_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		\n838gat_reg/NET0131 ,
		_w1051_,
		_w1088_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		_w396_,
		_w1085_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1086_,
		_w1087_,
		_w1090_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		_w1088_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w1089_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1084_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w1072_,
		_w1076_,
		_w1094_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w1093_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h4)
	) name898 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name900 (
		_w1036_,
		_w1042_,
		_w1098_
	);
	LUT2 #(
		.INIT('h4)
	) name901 (
		_w1068_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		_w1097_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		\n1389gat_reg/NET0131 ,
		_w1100_,
		_w1101_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		\n1508gat_reg/NET0131 ,
		_w422_,
		_w1102_
	);
	LUT2 #(
		.INIT('h8)
	) name905 (
		\n1678gat_reg/NET0131 ,
		_w422_,
		_w1103_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		\n1394gat_reg/NET0131 ,
		_w396_,
		_w1104_
	);
	LUT2 #(
		.INIT('h4)
	) name907 (
		_w1102_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h4)
	) name908 (
		_w1103_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name909 (
		\n1871gat_reg/NET0131 ,
		\n2592gat_reg/NET0131 ,
		_w1107_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		\n673gat_reg/NET0131 ,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h4)
	) name911 (
		\n322gat_reg/NET0131 ,
		_w1051_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name912 (
		\n314gat_reg/NET0131 ,
		_w1046_,
		_w1110_
	);
	LUT2 #(
		.INIT('h4)
	) name913 (
		\n366gat_reg/NET0131 ,
		_w1033_,
		_w1111_
	);
	LUT2 #(
		.INIT('h4)
	) name914 (
		\n553gat_reg/NET0131 ,
		_w334_,
		_w1112_
	);
	LUT2 #(
		.INIT('h4)
	) name915 (
		\n561gat_reg/NET0131 ,
		_w1039_,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name916 (
		\n659gat_reg/NET0131 ,
		_w485_,
		_w1114_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		\n777gat_reg/NET0131 ,
		_w310_,
		_w1115_
	);
	LUT2 #(
		.INIT('h4)
	) name918 (
		\n318gat_reg/NET0131 ,
		_w1049_,
		_w1116_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w1109_,
		_w1110_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1111_,
		_w1112_,
		_w1118_
	);
	LUT2 #(
		.INIT('h1)
	) name921 (
		_w1113_,
		_w1114_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w1115_,
		_w1116_,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name923 (
		_w1119_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		_w1117_,
		_w1118_,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name925 (
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h2)
	) name926 (
		_w487_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		\n919gat_reg/NET0131 ,
		_w234_,
		_w1125_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		\n919gat_reg/NET0131 ,
		_w234_,
		_w1126_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		_w308_,
		_w485_,
		_w1127_
	);
	LUT2 #(
		.INIT('h4)
	) name930 (
		_w1125_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w1126_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1124_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		_w608_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name934 (
		_w1106_,
		_w1108_,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		_w1101_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h4)
	) name936 (
		_w1131_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		_w459_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h4)
	) name938 (
		_w752_,
		_w1134_,
		_w1136_
	);
	LUT2 #(
		.INIT('h8)
	) name939 (
		\n2514gat_reg/NET0131 ,
		_w846_,
		_w1137_
	);
	LUT2 #(
		.INIT('h2)
	) name940 (
		_w609_,
		_w1137_,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		\n1871gat_reg/NET0131 ,
		_w1137_,
		_w1139_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		\n2033gat_reg/NET0131 ,
		\n2110gat_reg/NET0131 ,
		_w1140_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		\n2169gat_reg/NET0131 ,
		\n2176gat_reg/NET0131 ,
		_w1141_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		_w1140_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		_w493_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		_w1139_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		\n2454gat_reg/NET0131 ,
		\n337gat_reg/NET0131 ,
		_w1145_
	);
	LUT2 #(
		.INIT('h2)
	) name948 (
		_w546_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name949 (
		_w362_,
		_w835_,
		_w1147_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		_w537_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w838_,
		_w1148_,
		_w1149_
	);
	assign \_al_n0  = 1'b0;
	assign \g17_dup/_0_  = _w200_ ;
	assign \g6952/_2_  = _w295_ ;
	assign \g6953/_2_  = _w301_ ;
	assign \g6961/_0_  = _w304_ ;
	assign \g7076/_0_  = _w340_ ;
	assign \g7077/_0_  = _w344_ ;
	assign \g7079/_0_  = _w348_ ;
	assign \g7081/_0_  = _w352_ ;
	assign \g7082/_0_  = _w356_ ;
	assign \g7083/_0_  = _w360_ ;
	assign \g7146/_0_  = _w376_ ;
	assign \g7147/_0_  = _w378_ ;
	assign \g7148/_0_  = _w380_ ;
	assign \g7149/_0_  = _w382_ ;
	assign \g7150/_0_  = _w384_ ;
	assign \g7151/_0_  = _w386_ ;
	assign \g7152/_0_  = _w388_ ;
	assign \g7153/_0_  = _w390_ ;
	assign \g7154/_0_  = _w392_ ;
	assign \g7156/_2_  = _w443_ ;
	assign \g7161/_2_  = _w446_ ;
	assign \g7165/_2_  = _w459_ ;
	assign \g7174/_0_  = _w460_ ;
	assign \g7180/_00_  = _w484_ ;
	assign \g7182/_3_  = _w489_ ;
	assign \g7191/_0_  = _w496_ ;
	assign \g7204/_0_  = _w501_ ;
	assign \g7209/_3_  = _w525_ ;
	assign \g7220/_0_  = \n2543gat_reg/NET0131 ;
	assign \g7229/_0_  = _w534_ ;
	assign \g7233/_0_  = _w536_ ;
	assign \g7234/_0_  = _w539_ ;
	assign \g7235/_0_  = _w542_ ;
	assign \g7236/_0_  = _w547_ ;
	assign \g7237/_0_  = _w550_ ;
	assign \g7238/_0_  = _w556_ ;
	assign \g7241/_3_  = _w577_ ;
	assign \g7264/_0_  = _w583_ ;
	assign \g7265/_0_  = _w589_ ;
	assign \g7266/_0_  = _w596_ ;
	assign \g7267/_0_  = _w599_ ;
	assign \g7268/_0_  = _w600_ ;
	assign \g7301/_0_  = _w603_ ;
	assign \g7326/_3_  = _w606_ ;
	assign \g7350/_2_  = _w609_ ;
	assign \g7352/_0_  = \n838gat_reg/NET0131 ;
	assign \g7356/_0_  = _w611_ ;
	assign \g7359/_0_  = _w440_ ;
	assign \g7389/_3_  = _w635_ ;
	assign \g7417/_0_  = _w642_ ;
	assign \g7418/_0_  = _w644_ ;
	assign \g7419/_0_  = _w646_ ;
	assign \g7444/_0_  = _w664_ ;
	assign \g7445/_0_  = _w676_ ;
	assign \g7449/_3_  = _w685_ ;
	assign \g7451/_3_  = _w701_ ;
	assign \g7454/_0_  = \n707gat_reg/NET0131 ;
	assign \g7467/_3_  = _w706_ ;
	assign \g7476/_0_  = \n614gat_reg/NET0131 ;
	assign \g7480/_0_  = _w714_ ;
	assign \g7494/_0_  = _w719_ ;
	assign \g7509/_0_  = \n2176gat_reg/NET0131 ;
	assign \g7514/_0_  = _w722_ ;
	assign \g7517/_3_  = _w727_ ;
	assign \g7524/_0_  = \n2095gat_reg/NET0131 ;
	assign \g7558/_0_  = _w730_ ;
	assign \g7560/_0_  = _w733_ ;
	assign \g7561/_0_  = _w736_ ;
	assign \g7563/_0_  = _w739_ ;
	assign \g7567/_0_  = _w752_ ;
	assign \g7572/_0_  = \n1821gat_reg/NET0131 ;
	assign \g7579/_0_  = _w754_ ;
	assign \g7605/_0_  = _w758_ ;
	assign \g7625/_0_  = _w759_ ;
	assign \g7627/_0_  = _w721_ ;
	assign \g7671/_0_  = _w761_ ;
	assign \g7675/_0_  = _w766_ ;
	assign \g7689/_0_  = _w767_ ;
	assign \g7697/_0_  = _w769_ ;
	assign \g7743/_1_  = _w636_ ;
	assign \g7764/_1_  = _w645_ ;
	assign \g7769/_0_  = _w771_ ;
	assign \g7771/_2_  = _w768_ ;
	assign \g7779/_0_  = _w772_ ;
	assign \g7852/_0_  = _w774_ ;
	assign \g7873/_0_  = _w775_ ;
	assign \g7884/_3_  = _w473_ ;
	assign \g7889/_0_  = \n2110gat_reg/NET0131 ;
	assign \g7902/_1_  = _w643_ ;
	assign \g7992/_3_  = _w778_ ;
	assign \g7994/_3_  = _w343_ ;
	assign \g7996/_3_  = _w351_ ;
	assign \g7998/_3_  = _w781_ ;
	assign \g8000/_3_  = _w784_ ;
	assign \g8002/_3_  = _w307_ ;
	assign \g8004/_3_  = _w359_ ;
	assign \g8006/_3_  = _w355_ ;
	assign \g8008/_3_  = _w347_ ;
	assign \g8150/_0_  = \n2626gat_reg/NET0131 ;
	assign \g8151/_0_  = \n2495gat_reg/NET0131 ;
	assign \g8157/_0_  = \n2037gat_reg/NET0131 ;
	assign \g8163/_0_  = \n830gat_reg/NET0131 ;
	assign \g8172/_0_  = \n2490gat_reg/NET0131 ;
	assign \g8197/_0_  = \n834gat_reg/NET0131 ;
	assign \g8211/_0_  = \n2562gat_reg/NET0131 ;
	assign \g8223/_0_  = \n2634gat_reg/NET0131 ;
	assign \g8237/_0_  = \n2203gat_reg/NET0131 ;
	assign \g8251/_0_  = \n2640gat_reg/NET0131 ;
	assign \g8261/_0_  = \n820gat_reg/NET0131 ;
	assign \g8272/_0_  = \n1316gat_reg/NET0131 ;
	assign \g8287/_0_  = \n699gat_reg/NET0131 ;
	assign \g8647/_0_  = \n2207gat_reg/NET0131 ;
	assign \g8671/_0_  = \n2343gat_reg/NET0131 ;
	assign \g8672/_0_  = \n2399gat_reg/NET0131 ;
	assign \g8735/_0_  = _w799_ ;
	assign \g8766/_0_  = _w800_ ;
	assign \g8811/_0_  = _w801_ ;
	assign \g8821/_0_  = _w809_ ;
	assign \g8856/_0_  = _w578_ ;
	assign \g8858/_3_  = _w495_ ;
	assign \g8868/_0_  = _w422_ ;
	assign \g8880/_2_  = _w538_ ;
	assign \g8886/_0_  = _w820_ ;
	assign \g8900/_0_  = _w821_ ;
	assign \g8932/_0_  = _w828_ ;
	assign \g8991/_3_  = _w436_ ;
	assign \g9014/_3_  = _w831_ ;
	assign \g9074/_0_  = _w466_ ;
	assign \g9091/_0_  = \n2622gat_reg/NET0131 ;
	assign \g9105/_0_  = \n2630gat_reg/NET0131 ;
	assign \g9107/_1_  = _w332_ ;
	assign \g9111/_0_  = _w834_ ;
	assign \n1332gat_reg/P0001  = \n1332gat_reg/NET0131 ;
	assign \n1363gat_reg/P0001  = \n1363gat_reg/NET0131 ;
	assign \n1394gat_reg/P0001  = \n1394gat_reg/NET0131 ;
	assign \n1433gat_reg/P0001  = \n1433gat_reg/NET0131 ;
	assign \n1775gat_reg/P0001  = \n1775gat_reg/NET0131 ;
	assign \n2025gat_reg/P0001  = \n2025gat_reg/NET0131 ;
	assign \n2029gat_reg/P0001  = \n2029gat_reg/NET0131 ;
	assign \n2033gat_reg/P0001  = \n2033gat_reg/NET0131 ;
	assign \n2044gat_reg/P0001  = \n2044gat_reg/NET0131 ;
	assign \n2121gat_reg/P0001  = \n2121gat_reg/NET0131 ;
	assign \n2125gat_reg/P0001  = \n2125gat_reg/NET0131 ;
	assign \n2458gat_reg/P0001  = \n2458gat_reg/NET0131 ;
	assign \n2472gat_reg/P0001  = \n2472gat_reg/NET0131 ;
	assign \n2592gat_reg/P0001  = \n2592gat_reg/NET0131 ;
	assign \n3104gat_pad  = _w841_ ;
	assign \n3105gat_pad  = _w845_ ;
	assign \n3106gat_pad  = \n1871gat_reg/NET0131 ;
	assign \n3107gat_pad  = _w847_ ;
	assign \n3108gat_pad  = _w848_ ;
	assign \n3109gat_pad  = _w849_ ;
	assign \n3110gat_pad  = _w850_ ;
	assign \n3111gat_pad  = _w851_ ;
	assign \n3112gat_pad  = 1'b0;
	assign \n3113gat_pad  = _w852_ ;
	assign \n3114gat_pad  = _w853_ ;
	assign \n3116gat_pad  = _w286_ ;
	assign \n3117gat_pad  = _w863_ ;
	assign \n3118gat_pad  = _w872_ ;
	assign \n3119gat_pad  = _w881_ ;
	assign \n3120gat_pad  = _w890_ ;
	assign \n3121gat_pad  = _w899_ ;
	assign \n3122gat_pad  = _w908_ ;
	assign \n3123gat_pad  = _w917_ ;
	assign \n3124gat_pad  = _w927_ ;
	assign \n3125gat_pad  = _w929_ ;
	assign \n3126gat_pad  = \n2339gat_reg/NET0131 ;
	assign \n3127gat_pad  = \n2270gat_reg/NET0131 ;
	assign \n3128gat_pad  = \n2390gat_reg/NET0131 ;
	assign \n3130gat_pad  = _w937_ ;
	assign \n3131gat_pad  = _w945_ ;
	assign \n3132gat_pad  = _w953_ ;
	assign \n3133gat_pad  = _w961_ ;
	assign \n3134gat_pad  = _w968_ ;
	assign \n3135gat_pad  = _w974_ ;
	assign \n3136gat_pad  = _w980_ ;
	assign \n3137gat_pad  = _w986_ ;
	assign \n3138gat_pad  = _w988_ ;
	assign \n3140gat_pad  = _w1016_ ;
	assign \n3142gat_pad  = _w1029_ ;
	assign \n3143gat_pad  = _w1135_ ;
	assign \n3144gat_pad  = _w1136_ ;
	assign \n3145gat_pad  = _w1138_ ;
	assign \n3146gat_pad  = _w1144_ ;
	assign \n3147gat_pad  = _w638_ ;
	assign \n3148gat_pad  = \n2450gat_reg/NET0131 ;
	assign \n3149gat_pad  = _w396_ ;
	assign \n3150gat_pad  = _w1146_ ;
	assign \n3151gat_pad  = _w1149_ ;
	assign \n684gat_reg/P0001  = \n684gat_reg/NET0131 ;
	assign \n824gat_reg/P0001  = \n824gat_reg/NET0131 ;
	assign \n883gat_reg/P0001  = \n883gat_reg/NET0131 ;
endmodule;