module top( \G0_pad  , \G10_pad  , \G11_pad  , \G12_pad  , \G13_pad  , \G1_pad  , \G29_reg/NET0131  , \G2_pad  , \G30_reg/NET0131  , \G31_reg/NET0131  , \G32_reg/NET0131  , \G33_reg/NET0131  , \G34_reg/NET0131  , \G35_reg/NET0131  , \G36_reg/NET0131  , \G37_reg/NET0131  , \G38_reg/NET0131  , \G39_reg/NET0131  , \G3_pad  , \G40_reg/NET0131  , \G41_reg/NET0131  , \G42_reg/NET0131  , \G43_reg/NET0131  , \G44_reg/NET0131  , \G46_reg/NET0131  , \G4_pad  , \G5_pad  , \G6_pad  , \G7_pad  , \G8_pad  , \G9_pad  , \G530_pad  , \G532_pad  , \G542_pad  , \G546_pad  , \G547_pad  , \G548_pad  , \G549_pad  , \G550_pad  , \G551_pad  , \G552_pad  , \_al_n0  , \_al_n1  , \g1594/_3_  , \g1613/_0_  , \g1618/_0_  , \g1620/_2_  , \g1692/_0_  , \g1727/_0_  , \g1740/_0_  , \g1742/_0_  , \g1760/_0_  , \g1769/_3_  , \g1771/_0_  , \g1780/_0_  , \g1799/_0_  , \g1867/_0_  , \g1873/_0_  , \g1900/_0_  , \g1930/_0_  , \g1936/_0_  , \g2340/_2_  , \g2396/_1_  , \g2408/_0_  );
  input \G0_pad  ;
  input \G10_pad  ;
  input \G11_pad  ;
  input \G12_pad  ;
  input \G13_pad  ;
  input \G1_pad  ;
  input \G29_reg/NET0131  ;
  input \G2_pad  ;
  input \G30_reg/NET0131  ;
  input \G31_reg/NET0131  ;
  input \G32_reg/NET0131  ;
  input \G33_reg/NET0131  ;
  input \G34_reg/NET0131  ;
  input \G35_reg/NET0131  ;
  input \G36_reg/NET0131  ;
  input \G37_reg/NET0131  ;
  input \G38_reg/NET0131  ;
  input \G39_reg/NET0131  ;
  input \G3_pad  ;
  input \G40_reg/NET0131  ;
  input \G41_reg/NET0131  ;
  input \G42_reg/NET0131  ;
  input \G43_reg/NET0131  ;
  input \G44_reg/NET0131  ;
  input \G46_reg/NET0131  ;
  input \G4_pad  ;
  input \G5_pad  ;
  input \G6_pad  ;
  input \G7_pad  ;
  input \G8_pad  ;
  input \G9_pad  ;
  output \G530_pad  ;
  output \G532_pad  ;
  output \G542_pad  ;
  output \G546_pad  ;
  output \G547_pad  ;
  output \G548_pad  ;
  output \G549_pad  ;
  output \G550_pad  ;
  output \G551_pad  ;
  output \G552_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1594/_3_  ;
  output \g1613/_0_  ;
  output \g1618/_0_  ;
  output \g1620/_2_  ;
  output \g1692/_0_  ;
  output \g1727/_0_  ;
  output \g1740/_0_  ;
  output \g1742/_0_  ;
  output \g1760/_0_  ;
  output \g1769/_3_  ;
  output \g1771/_0_  ;
  output \g1780/_0_  ;
  output \g1799/_0_  ;
  output \g1867/_0_  ;
  output \g1873/_0_  ;
  output \g1900/_0_  ;
  output \g1930/_0_  ;
  output \g1936/_0_  ;
  output \g2340/_2_  ;
  output \g2396/_1_  ;
  output \g2408/_0_  ;
  wire n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 ;
  assign n32 = \G3_pad  & ~\G4_pad  ;
  assign n33 = \G11_pad  & ~\G5_pad  ;
  assign n34 = \G35_reg/NET0131  & n33 ;
  assign n35 = n32 & n34 ;
  assign n36 = \G2_pad  & n35 ;
  assign n37 = ~\G7_pad  & ~\G8_pad  ;
  assign n38 = ~\G10_pad  & ~\G11_pad  ;
  assign n39 = n37 & n38 ;
  assign n40 = \G9_pad  & n39 ;
  assign n41 = \G10_pad  & \G7_pad  ;
  assign n42 = \G11_pad  & \G9_pad  ;
  assign n43 = \G8_pad  & n42 ;
  assign n44 = n41 & n43 ;
  assign n45 = ~n40 & ~n44 ;
  assign n46 = \G4_pad  & \G6_pad  ;
  assign n47 = \G3_pad  & \G5_pad  ;
  assign n48 = n46 & n47 ;
  assign n49 = \G2_pad  & n48 ;
  assign n50 = ~n45 & n49 ;
  assign n51 = ~n36 & ~n50 ;
  assign n52 = ~\G10_pad  & \G7_pad  ;
  assign n53 = \G10_pad  & \G9_pad  ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = \G7_pad  & ~\G8_pad  ;
  assign n56 = \G8_pad  & \G9_pad  ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = ~n54 & n57 ;
  assign n59 = \G11_pad  & \G5_pad  ;
  assign n60 = n46 & n59 ;
  assign n61 = ~\G3_pad  & n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = \G36_reg/NET0131  & ~\G3_pad  ;
  assign n64 = ~\G6_pad  & n63 ;
  assign n65 = ~n62 & ~n64 ;
  assign n66 = ~\G7_pad  & \G8_pad  ;
  assign n67 = ~\G10_pad  & \G9_pad  ;
  assign n68 = n66 & n67 ;
  assign n69 = ~n58 & ~n68 ;
  assign n70 = \G3_pad  & \G4_pad  ;
  assign n71 = \G6_pad  & n70 ;
  assign n72 = n33 & n71 ;
  assign n73 = ~n69 & n72 ;
  assign n74 = n65 & ~n73 ;
  assign n75 = ~\G2_pad  & ~n74 ;
  assign n76 = n51 & ~n75 ;
  assign n77 = n41 & ~n43 ;
  assign n78 = \G7_pad  & n67 ;
  assign n79 = \G30_reg/NET0131  & n66 ;
  assign n80 = ~n78 & ~n79 ;
  assign n81 = ~n77 & n80 ;
  assign n82 = \G32_reg/NET0131  & ~n81 ;
  assign n83 = ~\G13_pad  & ~n82 ;
  assign n84 = ~\G12_pad  & ~n65 ;
  assign n85 = n83 & n84 ;
  assign n86 = ~n76 & n85 ;
  assign n87 = \G11_pad  & \G8_pad  ;
  assign n88 = ~n38 & ~n87 ;
  assign n89 = ~\G6_pad  & \G7_pad  ;
  assign n90 = \G30_reg/NET0131  & n89 ;
  assign n91 = \G31_reg/NET0131  & \G8_pad  ;
  assign n92 = ~n67 & ~n91 ;
  assign n93 = ~n90 & n92 ;
  assign n94 = ~n88 & n93 ;
  assign n95 = ~\G31_reg/NET0131  & n56 ;
  assign n96 = ~\G8_pad  & n53 ;
  assign n97 = ~n95 & ~n96 ;
  assign n98 = ~\G11_pad  & ~\G7_pad  ;
  assign n99 = ~n97 & n98 ;
  assign n100 = ~n94 & ~n99 ;
  assign n101 = \G0_pad  & \G3_pad  ;
  assign n102 = ~\G3_pad  & \G5_pad  ;
  assign n103 = ~\G4_pad  & ~n102 ;
  assign n104 = ~n101 & n103 ;
  assign n105 = \G46_reg/NET0131  & ~n104 ;
  assign n106 = \G12_pad  & ~\G13_pad  ;
  assign n107 = ~\G30_reg/NET0131  & ~\G6_pad  ;
  assign n108 = \G11_pad  & n107 ;
  assign n109 = \G11_pad  & ~\G9_pad  ;
  assign n110 = n37 & n109 ;
  assign n111 = ~n108 & ~n110 ;
  assign n112 = n106 & n111 ;
  assign n113 = n105 & n112 ;
  assign n114 = n100 & n113 ;
  assign n115 = \G0_pad  & ~n32 ;
  assign n116 = \G1_pad  & ~n115 ;
  assign n117 = \G4_pad  & ~n47 ;
  assign n118 = ~\G1_pad  & \G5_pad  ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = ~n116 & n119 ;
  assign n121 = ~\G0_pad  & ~\G1_pad  ;
  assign n122 = \G2_pad  & ~n121 ;
  assign n123 = ~n120 & n122 ;
  assign n124 = n114 & n123 ;
  assign n125 = ~n86 & ~n124 ;
  assign n126 = \G1_pad  & \G3_pad  ;
  assign n127 = \G5_pad  & n126 ;
  assign n128 = \G2_pad  & n46 ;
  assign n129 = n127 & n128 ;
  assign n130 = ~n45 & n129 ;
  assign n131 = \G13_pad  & n130 ;
  assign n132 = ~\G1_pad  & \G3_pad  ;
  assign n133 = n46 & n132 ;
  assign n134 = ~\G4_pad  & \G6_pad  ;
  assign n135 = n126 & n134 ;
  assign n136 = ~n133 & ~n135 ;
  assign n137 = ~\G9_pad  & n52 ;
  assign n138 = n87 & n137 ;
  assign n139 = \G11_pad  & ~\G7_pad  ;
  assign n140 = n96 & n139 ;
  assign n141 = ~n138 & ~n140 ;
  assign n142 = ~n136 & ~n141 ;
  assign n143 = n67 & n87 ;
  assign n144 = ~\G7_pad  & n133 ;
  assign n145 = n143 & n144 ;
  assign n146 = ~\G8_pad  & n52 ;
  assign n147 = ~\G4_pad  & ~\G6_pad  ;
  assign n148 = n132 & n147 ;
  assign n149 = n109 & n148 ;
  assign n150 = n146 & n149 ;
  assign n151 = ~n145 & ~n150 ;
  assign n152 = ~n142 & n151 ;
  assign n153 = \G2_pad  & ~\G5_pad  ;
  assign n154 = \G13_pad  & n153 ;
  assign n155 = ~n152 & n154 ;
  assign n156 = ~n131 & ~n155 ;
  assign n157 = ~n71 & n156 ;
  assign n158 = \G10_pad  & ~\G8_pad  ;
  assign n159 = n42 & n158 ;
  assign n160 = ~n156 & n159 ;
  assign n161 = n83 & n159 ;
  assign n162 = ~n76 & n161 ;
  assign n163 = ~n160 & ~n162 ;
  assign n164 = ~n157 & ~n163 ;
  assign n165 = \G5_pad  & \G9_pad  ;
  assign n166 = n39 & n165 ;
  assign n167 = \G6_pad  & n166 ;
  assign n168 = n58 & n134 ;
  assign n169 = ~n167 & ~n168 ;
  assign n170 = ~n156 & ~n169 ;
  assign n171 = n83 & ~n169 ;
  assign n172 = ~n76 & n171 ;
  assign n173 = ~n170 & ~n172 ;
  assign n174 = ~\G5_pad  & ~n134 ;
  assign n175 = ~\G1_pad  & \G2_pad  ;
  assign n176 = ~n174 & n175 ;
  assign n177 = ~n81 & n176 ;
  assign n178 = ~n46 & n47 ;
  assign n179 = ~\G2_pad  & \G3_pad  ;
  assign n180 = \G6_pad  & n179 ;
  assign n181 = ~n178 & ~n180 ;
  assign n182 = \G4_pad  & ~\G5_pad  ;
  assign n183 = ~\G3_pad  & n182 ;
  assign n184 = n181 & ~n183 ;
  assign n185 = \G2_pad  & ~\G3_pad  ;
  assign n186 = \G6_pad  & n185 ;
  assign n187 = n46 & ~n47 ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = \G2_pad  & \G4_pad  ;
  assign n190 = ~\G4_pad  & \G5_pad  ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = ~\G6_pad  & ~n191 ;
  assign n193 = n188 & ~n192 ;
  assign n194 = n184 & n193 ;
  assign n195 = \G1_pad  & ~n81 ;
  assign n196 = ~n194 & n195 ;
  assign n197 = ~n177 & ~n196 ;
  assign n198 = \G13_pad  & ~\G43_reg/NET0131  ;
  assign n199 = ~n197 & n198 ;
  assign n200 = n60 & n137 ;
  assign n201 = ~n147 & ~n200 ;
  assign n202 = ~\G3_pad  & ~n201 ;
  assign n203 = n83 & n202 ;
  assign n204 = ~n76 & n203 ;
  assign n205 = ~n199 & ~n204 ;
  assign n206 = n173 & n205 ;
  assign n207 = ~n164 & n206 ;
  assign n208 = ~\G12_pad  & ~n207 ;
  assign n209 = \G5_pad  & n179 ;
  assign n210 = \G4_pad  & n209 ;
  assign n211 = ~\G3_pad  & ~\G5_pad  ;
  assign n212 = ~\G2_pad  & ~n211 ;
  assign n213 = \G4_pad  & ~n126 ;
  assign n214 = ~n212 & n213 ;
  assign n215 = ~n210 & ~n214 ;
  assign n216 = \G1_pad  & ~n70 ;
  assign n217 = ~n185 & n216 ;
  assign n218 = n215 & ~n217 ;
  assign n219 = \G0_pad  & ~n218 ;
  assign n220 = n114 & n219 ;
  assign n221 = ~n208 & ~n220 ;
  assign n222 = \G34_reg/NET0131  & \G8_pad  ;
  assign n223 = n78 & n222 ;
  assign n224 = \G6_pad  & n78 ;
  assign n225 = n114 & n224 ;
  assign n226 = ~n223 & ~n225 ;
  assign n227 = \G34_reg/NET0131  & ~n56 ;
  assign n228 = n41 & n227 ;
  assign n229 = ~\G10_pad  & ~n55 ;
  assign n230 = ~\G9_pad  & ~n229 ;
  assign n231 = \G10_pad  & \G8_pad  ;
  assign n232 = \G7_pad  & \G9_pad  ;
  assign n233 = n231 & ~n232 ;
  assign n234 = ~n159 & ~n233 ;
  assign n235 = ~n230 & n234 ;
  assign n236 = \G6_pad  & ~n235 ;
  assign n237 = n114 & n236 ;
  assign n238 = ~n228 & ~n237 ;
  assign n239 = n226 & n238 ;
  assign n240 = n53 & n89 ;
  assign n241 = \G10_pad  & ~\G9_pad  ;
  assign n242 = ~n38 & n66 ;
  assign n243 = ~n241 & n242 ;
  assign n244 = ~\G8_pad  & n42 ;
  assign n245 = ~n66 & n67 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = ~n243 & n246 ;
  assign n248 = \G6_pad  & ~n247 ;
  assign n249 = ~n240 & ~n248 ;
  assign n250 = n114 & ~n249 ;
  assign n251 = ~\G7_pad  & ~n231 ;
  assign n252 = \G8_pad  & n41 ;
  assign n253 = \G34_reg/NET0131  & \G9_pad  ;
  assign n254 = ~n252 & n253 ;
  assign n255 = ~n251 & n254 ;
  assign n256 = ~n250 & ~n255 ;
  assign n257 = ~\G42_reg/NET0131  & n114 ;
  assign n258 = ~\G10_pad  & ~\G7_pad  ;
  assign n259 = \G9_pad  & n258 ;
  assign n260 = ~n37 & ~n259 ;
  assign n261 = n231 & n232 ;
  assign n262 = ~n137 & ~n261 ;
  assign n263 = n260 & n262 ;
  assign n264 = \G11_pad  & \G34_reg/NET0131  ;
  assign n265 = n263 & n264 ;
  assign n266 = ~n257 & ~n265 ;
  assign n267 = ~\G12_pad  & \G13_pad  ;
  assign n268 = n46 & n102 ;
  assign n269 = ~n209 & ~n268 ;
  assign n270 = ~n32 & n153 ;
  assign n271 = ~n190 & ~n270 ;
  assign n272 = n269 & n271 ;
  assign n273 = \G1_pad  & ~n272 ;
  assign n274 = n267 & n273 ;
  assign n275 = ~n197 & n274 ;
  assign n276 = \G1_pad  & \G4_pad  ;
  assign n277 = ~n101 & n276 ;
  assign n278 = n114 & n277 ;
  assign n279 = ~\G13_pad  & ~\G33_reg/NET0131  ;
  assign n280 = \G3_pad  & n279 ;
  assign n281 = ~\G12_pad  & \G32_reg/NET0131  ;
  assign n282 = ~\G13_pad  & n281 ;
  assign n283 = ~n81 & n282 ;
  assign n284 = \G2_pad  & \G5_pad  ;
  assign n285 = ~n70 & n284 ;
  assign n286 = n283 & n285 ;
  assign n287 = ~n280 & ~n286 ;
  assign n288 = ~n278 & n287 ;
  assign n289 = ~n275 & n288 ;
  assign n290 = ~n276 & n284 ;
  assign n291 = n153 & n276 ;
  assign n292 = ~n290 & ~n291 ;
  assign n293 = n267 & ~n292 ;
  assign n294 = ~n197 & n293 ;
  assign n295 = ~\G0_pad  & \G3_pad  ;
  assign n296 = n276 & n295 ;
  assign n297 = \G0_pad  & ~\G29_reg/NET0131  ;
  assign n298 = ~n296 & ~n297 ;
  assign n299 = n114 & ~n298 ;
  assign n300 = n47 & ~n189 ;
  assign n301 = n283 & n300 ;
  assign n302 = ~n280 & ~n301 ;
  assign n303 = ~n299 & n302 ;
  assign n304 = ~n294 & n303 ;
  assign n305 = ~\G3_pad  & n46 ;
  assign n306 = \G1_pad  & ~n182 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = ~\G5_pad  & \G6_pad  ;
  assign n309 = n179 & n308 ;
  assign n310 = ~\G2_pad  & n70 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = n307 & n311 ;
  assign n313 = ~\G1_pad  & ~n189 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = n267 & n314 ;
  assign n316 = ~n197 & n315 ;
  assign n317 = \G39_reg/NET0131  & \G4_pad  ;
  assign n318 = n283 & n317 ;
  assign n319 = ~\G0_pad  & n276 ;
  assign n320 = n101 & ~n276 ;
  assign n321 = ~n319 & ~n320 ;
  assign n322 = \G5_pad  & ~n321 ;
  assign n323 = \G0_pad  & \G2_pad  ;
  assign n324 = \G1_pad  & ~n323 ;
  assign n325 = \G0_pad  & n189 ;
  assign n326 = ~n324 & ~n325 ;
  assign n327 = n102 & ~n326 ;
  assign n328 = ~n322 & ~n327 ;
  assign n329 = n114 & ~n328 ;
  assign n330 = ~n318 & ~n329 ;
  assign n331 = ~n316 & n330 ;
  assign n332 = ~\G40_reg/NET0131  & n114 ;
  assign n333 = ~\G6_pad  & ~n332 ;
  assign n334 = \G4_pad  & ~n284 ;
  assign n335 = \G2_pad  & ~n276 ;
  assign n336 = ~n47 & ~n335 ;
  assign n337 = ~n334 & n336 ;
  assign n338 = n267 & ~n337 ;
  assign n339 = ~n197 & n338 ;
  assign n340 = \G2_pad  & n190 ;
  assign n341 = ~n47 & n189 ;
  assign n342 = ~n340 & ~n341 ;
  assign n343 = n179 & ~n182 ;
  assign n344 = n342 & ~n343 ;
  assign n345 = n283 & ~n344 ;
  assign n346 = ~n332 & ~n345 ;
  assign n347 = ~n339 & n346 ;
  assign n348 = ~n333 & ~n347 ;
  assign n349 = n139 & n158 ;
  assign n350 = \G6_pad  & ~\G9_pad  ;
  assign n351 = ~\G0_pad  & ~\G4_pad  ;
  assign n352 = n211 & n351 ;
  assign n353 = n350 & n352 ;
  assign n354 = n349 & n353 ;
  assign n355 = n52 & n351 ;
  assign n356 = \G37_reg/NET0131  & n47 ;
  assign n357 = n87 & n356 ;
  assign n358 = n355 & n357 ;
  assign n359 = \G0_pad  & n48 ;
  assign n360 = n44 & n359 ;
  assign n361 = ~n358 & ~n360 ;
  assign n362 = ~n354 & n361 ;
  assign n363 = \G1_pad  & \G2_pad  ;
  assign n364 = ~n362 & n363 ;
  assign n365 = n105 & n111 ;
  assign n366 = n100 & n365 ;
  assign n367 = n106 & n127 ;
  assign n368 = ~n366 & n367 ;
  assign n369 = n364 & n368 ;
  assign n370 = \G38_reg/NET0131  & n350 ;
  assign n371 = ~n41 & ~n370 ;
  assign n372 = n369 & ~n371 ;
  assign n373 = \G12_pad  & ~n372 ;
  assign n374 = n52 & n350 ;
  assign n375 = ~n47 & ~n374 ;
  assign n376 = \G8_pad  & ~n375 ;
  assign n377 = ~n156 & n376 ;
  assign n378 = n83 & n376 ;
  assign n379 = ~n76 & n378 ;
  assign n380 = ~n377 & ~n379 ;
  assign n381 = n58 & n71 ;
  assign n382 = ~n156 & n381 ;
  assign n383 = ~n372 & ~n382 ;
  assign n384 = n380 & n383 ;
  assign n385 = ~n373 & ~n384 ;
  assign n386 = \G2_pad  & n385 ;
  assign n387 = ~\G12_pad  & n83 ;
  assign n388 = n53 & n60 ;
  assign n389 = ~\G5_pad  & n38 ;
  assign n390 = n147 & n389 ;
  assign n391 = ~n388 & ~n390 ;
  assign n392 = n37 & ~n391 ;
  assign n393 = ~\G6_pad  & n182 ;
  assign n394 = n44 & n393 ;
  assign n395 = ~n381 & ~n394 ;
  assign n396 = ~n392 & n395 ;
  assign n397 = n387 & ~n396 ;
  assign n398 = ~n76 & n397 ;
  assign n399 = ~n386 & ~n398 ;
  assign n400 = \G2_pad  & n182 ;
  assign n401 = n281 & n400 ;
  assign n402 = ~n81 & n401 ;
  assign n403 = \G0_pad  & \G12_pad  ;
  assign n404 = \G1_pad  & ~\G4_pad  ;
  assign n405 = n403 & n404 ;
  assign n406 = n111 & n405 ;
  assign n407 = n105 & n406 ;
  assign n408 = n100 & n407 ;
  assign n409 = ~n402 & ~n408 ;
  assign n410 = ~n152 & n153 ;
  assign n411 = ~n130 & ~n410 ;
  assign n412 = n197 & n267 ;
  assign n413 = ~n411 & n412 ;
  assign n414 = ~n76 & n387 ;
  assign n415 = n106 & ~n366 ;
  assign n416 = n364 & n415 ;
  assign n417 = ~n414 & ~n416 ;
  assign n418 = ~n413 & n417 ;
  assign n419 = n411 & n412 ;
  assign n420 = ~n364 & n415 ;
  assign n421 = ~\G12_pad  & ~\G13_pad  ;
  assign n422 = ~n82 & n421 ;
  assign n423 = n51 & n422 ;
  assign n424 = ~n75 & n423 ;
  assign n425 = ~n420 & ~n424 ;
  assign n426 = ~n419 & n425 ;
  assign n427 = ~\G2_pad  & ~\G3_pad  ;
  assign n428 = ~n182 & n427 ;
  assign n429 = n179 & n182 ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = \G0_pad  & n430 ;
  assign n432 = ~\G1_pad  & ~n431 ;
  assign n433 = \G2_pad  & ~n118 ;
  assign n434 = ~n117 & n433 ;
  assign n435 = ~n116 & n434 ;
  assign n436 = ~\G10_pad  & ~\G30_reg/NET0131  ;
  assign n437 = \G7_pad  & ~n436 ;
  assign n438 = ~\G6_pad  & ~n437 ;
  assign n439 = ~n435 & ~n438 ;
  assign n440 = ~n432 & n439 ;
  assign n441 = \G6_pad  & \G9_pad  ;
  assign n442 = ~\G11_pad  & \G7_pad  ;
  assign n443 = n441 & n442 ;
  assign n444 = ~n90 & ~n443 ;
  assign n445 = \G8_pad  & ~n444 ;
  assign n446 = ~n91 & ~n143 ;
  assign n447 = \G6_pad  & ~n446 ;
  assign n448 = ~n445 & ~n447 ;
  assign n449 = ~\G9_pad  & n55 ;
  assign n450 = n231 & n350 ;
  assign n451 = ~n449 & ~n450 ;
  assign n452 = ~n67 & n89 ;
  assign n453 = ~n41 & n441 ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = n451 & n454 ;
  assign n456 = \G11_pad  & ~n455 ;
  assign n457 = ~\G6_pad  & n189 ;
  assign n458 = ~\G5_pad  & n46 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = n126 & ~n459 ;
  assign n461 = \G1_pad  & ~n181 ;
  assign n462 = \G3_pad  & n175 ;
  assign n463 = ~n174 & n462 ;
  assign n464 = ~n461 & ~n463 ;
  assign n465 = ~n460 & n464 ;
  assign n466 = n37 & n53 ;
  assign n467 = n60 & n466 ;
  assign n468 = ~\G4_pad  & n41 ;
  assign n469 = n43 & n468 ;
  assign n470 = ~\G9_pad  & n39 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = ~\G5_pad  & ~\G6_pad  ;
  assign n473 = ~n471 & n472 ;
  assign n474 = ~n467 & ~n473 ;
  assign n475 = \G6_pad  & n58 ;
  assign n476 = ~\G6_pad  & ~\G9_pad  ;
  assign n477 = n146 & n476 ;
  assign n478 = ~n475 & ~n477 ;
  assign n479 = ~\G5_pad  & n39 ;
  assign n480 = ~\G5_pad  & n41 ;
  assign n481 = n43 & n480 ;
  assign n482 = ~n479 & ~n481 ;
  assign n483 = ~n71 & n284 ;
  assign n484 = ~n174 & n179 ;
  assign n485 = ~n400 & ~n484 ;
  assign n486 = ~n483 & n485 ;
  assign n487 = ~n70 & ~n190 ;
  assign n488 = n175 & ~n487 ;
  assign n489 = ~n343 & ~n488 ;
  assign n490 = \G2_pad  & ~n47 ;
  assign n491 = ~n209 & ~n490 ;
  assign n492 = \G10_pad  & ~n42 ;
  assign n493 = ~n139 & ~n492 ;
  assign n494 = ~\G10_pad  & ~n109 ;
  assign n495 = ~n441 & ~n476 ;
  assign n496 = n41 & ~n441 ;
  assign n497 = n114 & n496 ;
  assign n498 = \G34_reg/NET0131  & n233 ;
  assign n499 = ~n497 & ~n498 ;
  assign n500 = n226 & n499 ;
  assign n501 = ~\G4_pad  & n58 ;
  assign n502 = ~n156 & n501 ;
  assign n503 = n83 & n501 ;
  assign n504 = ~n76 & n503 ;
  assign n505 = ~n502 & ~n504 ;
  assign n506 = ~\G7_pad  & ~\G9_pad  ;
  assign n507 = ~\G10_pad  & ~n506 ;
  assign n508 = n182 & n507 ;
  assign n509 = ~n156 & n508 ;
  assign n510 = n505 & ~n509 ;
  assign n511 = ~\G12_pad  & \G6_pad  ;
  assign n512 = ~n510 & n511 ;
  assign n513 = ~\G3_pad  & ~\G44_reg/NET0131  ;
  assign n514 = n72 & n507 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = ~\G12_pad  & ~n515 ;
  assign n517 = n83 & n516 ;
  assign n518 = ~n76 & n517 ;
  assign n519 = \G37_reg/NET0131  & \G38_reg/NET0131  ;
  assign n520 = n369 & n519 ;
  assign n521 = ~n518 & ~n520 ;
  assign n522 = ~n512 & n521 ;
  assign n523 = ~n197 & n267 ;
  assign n524 = ~n283 & ~n523 ;
  assign \G530_pad  = ~n125 ;
  assign \G532_pad  = ~n221 ;
  assign \G542_pad  = ~n239 ;
  assign \G546_pad  = ~\G41_reg/NET0131  ;
  assign \G547_pad  = ~n256 ;
  assign \G548_pad  = ~n266 ;
  assign \G549_pad  = ~n289 ;
  assign \G550_pad  = ~n304 ;
  assign \G551_pad  = ~n331 ;
  assign \G552_pad  = n348 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1594/_3_  = ~n399 ;
  assign \g1613/_0_  = n409 ;
  assign \g1618/_0_  = ~n418 ;
  assign \g1620/_2_  = ~n426 ;
  assign \g1692/_0_  = n440 ;
  assign \g1727/_0_  = n448 ;
  assign \g1740/_0_  = ~n456 ;
  assign \g1742/_0_  = n465 ;
  assign \g1760/_0_  = n474 ;
  assign \g1769/_3_  = ~n478 ;
  assign \g1771/_0_  = ~n482 ;
  assign \g1780/_0_  = ~n486 ;
  assign \g1799/_0_  = n489 ;
  assign \g1867/_0_  = ~n491 ;
  assign \g1873/_0_  = ~n493 ;
  assign \g1900/_0_  = n355 ;
  assign \g1930/_0_  = ~n494 ;
  assign \g1936/_0_  = n495 ;
  assign \g2340/_2_  = n500 ;
  assign \g2396/_1_  = ~n522 ;
  assign \g2408/_0_  = ~n524 ;
endmodule
