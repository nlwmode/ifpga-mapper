module top( \a0_pad  , \a1_pad  , \a2_pad  , \a3_pad  , \a4_pad  , \b0_pad  , \b1_pad  , \b2_pad  , \b3_pad  , \b4_pad  , \b5_pad  , b_pad , \c0_pad  , \c1_pad  , \c2_pad  , \c3_pad  , \c4_pad  , \c5_pad  , c_pad , \d0_pad  , \d1_pad  , \d2_pad  , \d3_pad  , \d4_pad  , \d5_pad  , d_pad , \e0_pad  , \e2_pad  , \e3_pad  , \e4_pad  , \e5_pad  , e_pad , \f0_pad  , \f1_pad  , \f2_pad  , \f3_pad  , \f4_pad  , \f5_pad  , f_pad , \g0_pad  , \g1_pad  , \g2_pad  , \g3_pad  , \g4_pad  , g_pad , \h0_pad  , \h1_pad  , \h2_pad  , \h3_pad  , \h4_pad  , \h5_pad  , h_pad , \i0_pad  , \i10_pad  , \i1_pad  , \i2_pad  , \i3_pad  , \i4_pad  , \i5_pad  , i_pad , \j0_pad  , \j2_pad  , \j3_pad  , \j4_pad  , \j5_pad  , j_pad , \k0_pad  , \k1_pad  , \k2_pad  , \k3_pad  , \k4_pad  , \k5_pad  , k_pad , \l0_pad  , \l1_pad  , \l2_pad  , \l3_pad  , \l4_pad  , \l5_pad  , \l6_pad  , l_pad , \m0_pad  , \m1_pad  , \m2_pad  , \m3_pad  , \m4_pad  , \m5_pad  , \m6_pad  , m_pad , \n0_pad  , \n1_pad  , \n2_pad  , \n3_pad  , \n4_pad  , \n5_pad  , n_pad , \o0_pad  , \o1_pad  , \o2_pad  , \o3_pad  , \o4_pad  , \o5_pad  , o_pad , \p0_pad  , \p10_pad  , \p1_pad  , \p2_pad  , \p3_pad  , \p4_pad  , \p5_pad  , p_pad , \q0_pad  , \q1_pad  , \q2_pad  , \q3_pad  , \q4_pad  , \q5_pad  , q_pad , \r0_pad  , \r1_pad  , \r2_pad  , \r3_pad  , \r4_pad  , \r5_pad  , \r6_pad  , r_pad , \s0_pad  , \s1_pad  , \s2_pad  , \s3_pad  , \s4_pad  , s_pad , \t0_pad  , \t1_pad  , \t2_pad  , \t3_pad  , \t4_pad  , t_pad , \u0_pad  , \u1_pad  , \u2_pad  , \u3_pad  , \u4_pad  , u_pad , \v0_pad  , \v1_pad  , \v2_pad  , \v3_pad  , \v4_pad  , v_pad , \w0_pad  , \w1_pad  , \w2_pad  , \w3_pad  , \w4_pad  , w_pad , \x0_pad  , \x1_pad  , \x2_pad  , \x3_pad  , \x4_pad  , \y0_pad  , \y1_pad  , \y2_pad  , \y3_pad  , \y4_pad  , \z0_pad  , \z1_pad  , \z2_pad  , \z3_pad  , \z4_pad  , z_pad , \a10_pad  , \a6_pad  , \a7_pad  , \a8_pad  , \a9_pad  , \b10_pad  , \b6_pad  , \b7_pad  , \b8_pad  , \b9_pad  , \c10_pad  , \c53  , \c6_pad  , \c7_pad  , \c8_pad  , \c9_pad  , \d10_pad  , \d6_pad  , \d7_pad  , \d8_pad  , \d9_pad  , \e10_pad  , \e6_pad  , \e7_pad  , \e8_pad  , \e9_pad  , \f10_pad  , \f22  , \f6_pad  , \f7_pad  , \f8_pad  , \f9_pad  , \g10_pad  , \g6_pad  , \g7_pad  , \g8_pad  , \g9_pad  , \h6_pad  , \h7_pad  , \h8_pad  , \h9_pad  , \i6_pad  , \i7_pad  , \i8_pad  , \i9_pad  , \j10_pad  , \j6_pad  , \j7_pad  , \j8_pad  , \j9_pad  , \k10_pad  , \k53  , \k6_pad  , \k7_pad  , \k8_pad  , \k9_pad  , \l10_pad  , \l7_pad  , \l8_pad  , \l9_pad  , \m10_pad  , \m7_pad  , \m8_pad  , \m9_pad  , \n10_pad  , \n6_pad  , \n7_pad  , \n8_pad  , \n9_pad  , \o10_pad  , \o6_pad  , \o7_pad  , \o8_pad  , \o9_pad  , \p6_pad  , \p7_pad  , \p8_pad  , \p9_pad  , \q10_pad  , \q6_pad  , \q7_pad  , \q8_pad  , \q9_pad  , \r10_pad  , \r7_pad  , \r8_pad  , \r9_pad  , \s5_pad  , \s7_pad  , \s8_pad  , \s9_pad  , \t10_pad  , \t5_pad  , \t6_pad  , \t7_pad  , \t8_pad  , \t9_pad  , \u5_pad  , \u7_pad  , \u8_pad  , \u9_pad  , \v10_pad  , \v5_pad  , \v6_pad  , \v7_pad  , \v8_pad  , \v9_pad  , \w10_pad  , \w5_pad  , \w6_pad  , \w7_pad  , \w8_pad  , \w9_pad  , \x10_pad  , \x21  , \x5_pad  , \x6_pad  , \x7_pad  , \x8_pad  , \x9_pad  , \y10_pad  , \y5_pad  , \y6_pad  , \y7_pad  , \y8_pad  , \y9_pad  , \z5_pad  , \z6_pad  , \z7_pad  , \z8_pad  , \z9_pad  );
  input \a0_pad  ;
  input \a1_pad  ;
  input \a2_pad  ;
  input \a3_pad  ;
  input \a4_pad  ;
  input \b0_pad  ;
  input \b1_pad  ;
  input \b2_pad  ;
  input \b3_pad  ;
  input \b4_pad  ;
  input \b5_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input \c1_pad  ;
  input \c2_pad  ;
  input \c3_pad  ;
  input \c4_pad  ;
  input \c5_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input \d1_pad  ;
  input \d2_pad  ;
  input \d3_pad  ;
  input \d4_pad  ;
  input \d5_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input \e2_pad  ;
  input \e3_pad  ;
  input \e4_pad  ;
  input \e5_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input \f1_pad  ;
  input \f2_pad  ;
  input \f3_pad  ;
  input \f4_pad  ;
  input \f5_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input \g1_pad  ;
  input \g2_pad  ;
  input \g3_pad  ;
  input \g4_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input \h1_pad  ;
  input \h2_pad  ;
  input \h3_pad  ;
  input \h4_pad  ;
  input \h5_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input \i10_pad  ;
  input \i1_pad  ;
  input \i2_pad  ;
  input \i3_pad  ;
  input \i4_pad  ;
  input \i5_pad  ;
  input i_pad ;
  input \j0_pad  ;
  input \j2_pad  ;
  input \j3_pad  ;
  input \j4_pad  ;
  input \j5_pad  ;
  input j_pad ;
  input \k0_pad  ;
  input \k1_pad  ;
  input \k2_pad  ;
  input \k3_pad  ;
  input \k4_pad  ;
  input \k5_pad  ;
  input k_pad ;
  input \l0_pad  ;
  input \l1_pad  ;
  input \l2_pad  ;
  input \l3_pad  ;
  input \l4_pad  ;
  input \l5_pad  ;
  input \l6_pad  ;
  input l_pad ;
  input \m0_pad  ;
  input \m1_pad  ;
  input \m2_pad  ;
  input \m3_pad  ;
  input \m4_pad  ;
  input \m5_pad  ;
  input \m6_pad  ;
  input m_pad ;
  input \n0_pad  ;
  input \n1_pad  ;
  input \n2_pad  ;
  input \n3_pad  ;
  input \n4_pad  ;
  input \n5_pad  ;
  input n_pad ;
  input \o0_pad  ;
  input \o1_pad  ;
  input \o2_pad  ;
  input \o3_pad  ;
  input \o4_pad  ;
  input \o5_pad  ;
  input o_pad ;
  input \p0_pad  ;
  input \p10_pad  ;
  input \p1_pad  ;
  input \p2_pad  ;
  input \p3_pad  ;
  input \p4_pad  ;
  input \p5_pad  ;
  input p_pad ;
  input \q0_pad  ;
  input \q1_pad  ;
  input \q2_pad  ;
  input \q3_pad  ;
  input \q4_pad  ;
  input \q5_pad  ;
  input q_pad ;
  input \r0_pad  ;
  input \r1_pad  ;
  input \r2_pad  ;
  input \r3_pad  ;
  input \r4_pad  ;
  input \r5_pad  ;
  input \r6_pad  ;
  input r_pad ;
  input \s0_pad  ;
  input \s1_pad  ;
  input \s2_pad  ;
  input \s3_pad  ;
  input \s4_pad  ;
  input s_pad ;
  input \t0_pad  ;
  input \t1_pad  ;
  input \t2_pad  ;
  input \t3_pad  ;
  input \t4_pad  ;
  input t_pad ;
  input \u0_pad  ;
  input \u1_pad  ;
  input \u2_pad  ;
  input \u3_pad  ;
  input \u4_pad  ;
  input u_pad ;
  input \v0_pad  ;
  input \v1_pad  ;
  input \v2_pad  ;
  input \v3_pad  ;
  input \v4_pad  ;
  input v_pad ;
  input \w0_pad  ;
  input \w1_pad  ;
  input \w2_pad  ;
  input \w3_pad  ;
  input \w4_pad  ;
  input w_pad ;
  input \x0_pad  ;
  input \x1_pad  ;
  input \x2_pad  ;
  input \x3_pad  ;
  input \x4_pad  ;
  input \y0_pad  ;
  input \y1_pad  ;
  input \y2_pad  ;
  input \y3_pad  ;
  input \y4_pad  ;
  input \z0_pad  ;
  input \z1_pad  ;
  input \z2_pad  ;
  input \z3_pad  ;
  input \z4_pad  ;
  input z_pad ;
  output \a10_pad  ;
  output \a6_pad  ;
  output \a7_pad  ;
  output \a8_pad  ;
  output \a9_pad  ;
  output \b10_pad  ;
  output \b6_pad  ;
  output \b7_pad  ;
  output \b8_pad  ;
  output \b9_pad  ;
  output \c10_pad  ;
  output \c53  ;
  output \c6_pad  ;
  output \c7_pad  ;
  output \c8_pad  ;
  output \c9_pad  ;
  output \d10_pad  ;
  output \d6_pad  ;
  output \d7_pad  ;
  output \d8_pad  ;
  output \d9_pad  ;
  output \e10_pad  ;
  output \e6_pad  ;
  output \e7_pad  ;
  output \e8_pad  ;
  output \e9_pad  ;
  output \f10_pad  ;
  output \f22  ;
  output \f6_pad  ;
  output \f7_pad  ;
  output \f8_pad  ;
  output \f9_pad  ;
  output \g10_pad  ;
  output \g6_pad  ;
  output \g7_pad  ;
  output \g8_pad  ;
  output \g9_pad  ;
  output \h6_pad  ;
  output \h7_pad  ;
  output \h8_pad  ;
  output \h9_pad  ;
  output \i6_pad  ;
  output \i7_pad  ;
  output \i8_pad  ;
  output \i9_pad  ;
  output \j10_pad  ;
  output \j6_pad  ;
  output \j7_pad  ;
  output \j8_pad  ;
  output \j9_pad  ;
  output \k10_pad  ;
  output \k53  ;
  output \k6_pad  ;
  output \k7_pad  ;
  output \k8_pad  ;
  output \k9_pad  ;
  output \l10_pad  ;
  output \l7_pad  ;
  output \l8_pad  ;
  output \l9_pad  ;
  output \m10_pad  ;
  output \m7_pad  ;
  output \m8_pad  ;
  output \m9_pad  ;
  output \n10_pad  ;
  output \n6_pad  ;
  output \n7_pad  ;
  output \n8_pad  ;
  output \n9_pad  ;
  output \o10_pad  ;
  output \o6_pad  ;
  output \o7_pad  ;
  output \o8_pad  ;
  output \o9_pad  ;
  output \p6_pad  ;
  output \p7_pad  ;
  output \p8_pad  ;
  output \p9_pad  ;
  output \q10_pad  ;
  output \q6_pad  ;
  output \q7_pad  ;
  output \q8_pad  ;
  output \q9_pad  ;
  output \r10_pad  ;
  output \r7_pad  ;
  output \r8_pad  ;
  output \r9_pad  ;
  output \s5_pad  ;
  output \s7_pad  ;
  output \s8_pad  ;
  output \s9_pad  ;
  output \t10_pad  ;
  output \t5_pad  ;
  output \t6_pad  ;
  output \t7_pad  ;
  output \t8_pad  ;
  output \t9_pad  ;
  output \u5_pad  ;
  output \u7_pad  ;
  output \u8_pad  ;
  output \u9_pad  ;
  output \v10_pad  ;
  output \v5_pad  ;
  output \v6_pad  ;
  output \v7_pad  ;
  output \v8_pad  ;
  output \v9_pad  ;
  output \w10_pad  ;
  output \w5_pad  ;
  output \w6_pad  ;
  output \w7_pad  ;
  output \w8_pad  ;
  output \w9_pad  ;
  output \x10_pad  ;
  output \x21  ;
  output \x5_pad  ;
  output \x6_pad  ;
  output \x7_pad  ;
  output \x8_pad  ;
  output \x9_pad  ;
  output \y10_pad  ;
  output \y5_pad  ;
  output \y6_pad  ;
  output \y7_pad  ;
  output \y8_pad  ;
  output \y9_pad  ;
  output \z5_pad  ;
  output \z6_pad  ;
  output \z7_pad  ;
  output \z8_pad  ;
  output \z9_pad  ;
  wire n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 ;
  assign n173 = ~\n5_pad  & ~z_pad ;
  assign n174 = \l5_pad  & \m5_pad  ;
  assign n175 = n173 & n174 ;
  assign n176 = \r5_pad  & n175 ;
  assign n182 = ~\i5_pad  & \o5_pad  ;
  assign n183 = \p10_pad  & n182 ;
  assign n184 = ~\d5_pad  & ~\e5_pad  ;
  assign n185 = ~\b5_pad  & \i10_pad  ;
  assign n186 = n184 & n185 ;
  assign n187 = ~n183 & n186 ;
  assign n188 = ~\e5_pad  & ~n187 ;
  assign n189 = ~\c5_pad  & n188 ;
  assign n190 = n184 & ~n185 ;
  assign n191 = n183 & n190 ;
  assign n192 = ~\d5_pad  & ~n191 ;
  assign n193 = n189 & n192 ;
  assign n199 = ~n176 & n193 ;
  assign n200 = \r4_pad  & ~n199 ;
  assign n201 = \s4_pad  & n200 ;
  assign n203 = ~\t4_pad  & ~n201 ;
  assign n177 = \r4_pad  & n176 ;
  assign n178 = \l5_pad  & ~\m5_pad  ;
  assign n179 = \n5_pad  & ~z_pad ;
  assign n180 = n178 & n179 ;
  assign n181 = ~z_pad & ~n180 ;
  assign n194 = ~\l5_pad  & ~\m5_pad  ;
  assign n195 = ~\n5_pad  & n194 ;
  assign n196 = n193 & n195 ;
  assign n197 = n181 & ~n196 ;
  assign n198 = ~n177 & n197 ;
  assign n202 = \t4_pad  & n201 ;
  assign n204 = n198 & ~n202 ;
  assign n205 = ~n203 & n204 ;
  assign n216 = \m4_pad  & \q0_pad  ;
  assign n214 = \n0_pad  & \p5_pad  ;
  assign n215 = \f3_pad  & \m0_pad  ;
  assign n221 = ~n214 & ~n215 ;
  assign n222 = ~n216 & n221 ;
  assign n210 = \m5_pad  & \p0_pad  ;
  assign n211 = \h4_pad  & \r0_pad  ;
  assign n219 = ~n210 & ~n211 ;
  assign n212 = \k0_pad  & \q3_pad  ;
  assign n213 = \l0_pad  & \m3_pad  ;
  assign n220 = ~n212 & ~n213 ;
  assign n223 = n219 & n220 ;
  assign n206 = \o0_pad  & \r5_pad  ;
  assign n207 = \r4_pad  & \u0_pad  ;
  assign n217 = ~n206 & ~n207 ;
  assign n208 = \t0_pad  & \w4_pad  ;
  assign n209 = \d4_pad  & \s0_pad  ;
  assign n218 = ~n208 & ~n209 ;
  assign n224 = n217 & n218 ;
  assign n225 = n223 & n224 ;
  assign n226 = n222 & n225 ;
  assign n244 = ~\k1_pad  & \o1_pad  ;
  assign n245 = \r6_pad  & n244 ;
  assign n246 = ~\h1_pad  & ~\i1_pad  ;
  assign n247 = ~\f1_pad  & \m6_pad  ;
  assign n248 = n246 & n247 ;
  assign n249 = ~n245 & n248 ;
  assign n250 = ~\i1_pad  & ~n249 ;
  assign n251 = ~\g1_pad  & n250 ;
  assign n252 = ~i_pad & n251 ;
  assign n253 = \s1_pad  & n252 ;
  assign n254 = ~\s1_pad  & ~n252 ;
  assign n230 = ~\a1_pad  & ~\b1_pad  ;
  assign n231 = ~\c1_pad  & n230 ;
  assign n256 = \r1_pad  & n231 ;
  assign n257 = ~\q1_pad  & ~n256 ;
  assign n258 = ~\z0_pad  & ~n257 ;
  assign n259 = ~\p1_pad  & ~n258 ;
  assign n237 = ~\l1_pad  & ~\m1_pad  ;
  assign n238 = ~\n1_pad  & n237 ;
  assign n239 = ~b_pad & ~n238 ;
  assign n255 = ~\v0_pad  & ~n239 ;
  assign n232 = ~\x0_pad  & ~\y0_pad  ;
  assign n260 = \w0_pad  & n232 ;
  assign n261 = n255 & n260 ;
  assign n262 = ~n259 & n261 ;
  assign n263 = ~h_pad & ~n262 ;
  assign n264 = ~n254 & ~n263 ;
  assign n265 = ~n253 & n264 ;
  assign n267 = ~\t1_pad  & n265 ;
  assign n227 = ~b_pad & \l1_pad  ;
  assign n228 = ~\m1_pad  & n227 ;
  assign n229 = ~\n1_pad  & n228 ;
  assign n233 = ~\d1_pad  & ~\w0_pad  ;
  assign n234 = ~\z0_pad  & n233 ;
  assign n235 = n232 & n234 ;
  assign n236 = n231 & n235 ;
  assign n240 = \v0_pad  & ~n239 ;
  assign n241 = n236 & n240 ;
  assign n242 = ~n229 & ~n241 ;
  assign n266 = \t1_pad  & ~n265 ;
  assign n268 = n242 & ~n266 ;
  assign n269 = ~n267 & n268 ;
  assign n243 = ~\x2_pad  & ~n242 ;
  assign n270 = ~b_pad & ~n243 ;
  assign n271 = ~n269 & n270 ;
  assign n272 = ~n239 & ~n251 ;
  assign n273 = ~g_pad & ~n272 ;
  assign n274 = ~b_pad & \m1_pad  ;
  assign n275 = ~\n1_pad  & n274 ;
  assign n276 = ~\l1_pad  & n275 ;
  assign n277 = ~b_pad & ~n276 ;
  assign n278 = ~n273 & ~n277 ;
  assign n296 = n246 & ~n247 ;
  assign n297 = n245 & n296 ;
  assign n298 = ~\h1_pad  & ~n297 ;
  assign n299 = n251 & n298 ;
  assign n300 = n236 & n255 ;
  assign n301 = ~n299 & n300 ;
  assign n279 = \l1_pad  & n275 ;
  assign n294 = \r1_pad  & ~\v0_pad  ;
  assign n295 = n279 & ~n294 ;
  assign n302 = ~f_pad & ~n295 ;
  assign n303 = ~n301 & n302 ;
  assign n280 = ~j_pad & \q1_pad  ;
  assign n281 = n279 & n280 ;
  assign n282 = \q2_pad  & \r2_pad  ;
  assign n283 = ~n281 & ~n282 ;
  assign n284 = \s2_pad  & ~n283 ;
  assign n285 = ~j_pad & \p1_pad  ;
  assign n286 = n279 & n285 ;
  assign n287 = ~n284 & ~n286 ;
  assign n288 = ~n273 & n287 ;
  assign n289 = ~\q2_pad  & ~\r2_pad  ;
  assign n290 = ~n281 & ~n289 ;
  assign n291 = ~\s2_pad  & ~n290 ;
  assign n292 = ~n286 & ~n291 ;
  assign n293 = n273 & n292 ;
  assign n304 = ~n288 & ~n293 ;
  assign n305 = ~n303 & n304 ;
  assign n307 = \t2_pad  & n305 ;
  assign n306 = ~\t2_pad  & ~n305 ;
  assign n308 = n277 & ~n306 ;
  assign n309 = ~n307 & n308 ;
  assign n310 = ~n278 & ~n309 ;
  assign n311 = ~z_pad & ~n195 ;
  assign n312 = ~n189 & ~n311 ;
  assign n313 = ~\e0_pad  & ~n312 ;
  assign n314 = ~\l5_pad  & \m5_pad  ;
  assign n315 = n173 & n314 ;
  assign n316 = ~z_pad & ~n315 ;
  assign n317 = ~n313 & ~n316 ;
  assign n318 = ~\f3_pad  & ~\g3_pad  ;
  assign n319 = ~\h0_pad  & \q5_pad  ;
  assign n320 = n175 & n319 ;
  assign n321 = ~n318 & ~n320 ;
  assign n322 = ~\h3_pad  & ~n321 ;
  assign n323 = ~\h0_pad  & \p5_pad  ;
  assign n324 = n175 & n323 ;
  assign n325 = ~n322 & ~n324 ;
  assign n326 = ~\i3_pad  & ~n325 ;
  assign n327 = ~\h0_pad  & ~n326 ;
  assign n328 = \j3_pad  & ~n327 ;
  assign n329 = ~\p3_pad  & n328 ;
  assign n330 = ~\h0_pad  & ~n329 ;
  assign n331 = ~\q3_pad  & ~n330 ;
  assign n332 = ~\r3_pad  & n331 ;
  assign n333 = n313 & ~n332 ;
  assign n334 = \q3_pad  & \r3_pad  ;
  assign n335 = ~n313 & ~n334 ;
  assign n339 = ~\t4_pad  & ~\u4_pad  ;
  assign n340 = ~\v4_pad  & ~\w4_pad  ;
  assign n341 = ~\x4_pad  & ~\y4_pad  ;
  assign n342 = n340 & n341 ;
  assign n343 = n339 & n342 ;
  assign n344 = ~\s4_pad  & ~\z4_pad  ;
  assign n345 = ~n311 & n344 ;
  assign n346 = n343 & n345 ;
  assign n347 = ~\r4_pad  & n346 ;
  assign n348 = ~n193 & n347 ;
  assign n336 = ~\j5_pad  & \k5_pad  ;
  assign n337 = ~\r4_pad  & \r5_pad  ;
  assign n338 = n336 & ~n337 ;
  assign n349 = ~\d0_pad  & ~n338 ;
  assign n350 = ~n348 & n349 ;
  assign n351 = \f3_pad  & \g3_pad  ;
  assign n352 = ~n320 & ~n351 ;
  assign n353 = \h3_pad  & ~n352 ;
  assign n354 = ~n324 & ~n353 ;
  assign n355 = \i3_pad  & ~n354 ;
  assign n356 = ~\h0_pad  & ~n355 ;
  assign n357 = \k3_pad  & ~n356 ;
  assign n358 = \p3_pad  & n357 ;
  assign n359 = ~\h0_pad  & ~n313 ;
  assign n360 = ~n358 & n359 ;
  assign n361 = ~n350 & ~n360 ;
  assign n362 = ~n335 & n361 ;
  assign n363 = ~n333 & n362 ;
  assign n364 = ~\s3_pad  & ~n313 ;
  assign n365 = \s3_pad  & n313 ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = n363 & n366 ;
  assign n369 = \t3_pad  & n367 ;
  assign n368 = ~\t3_pad  & ~n367 ;
  assign n370 = n316 & ~n368 ;
  assign n371 = ~n369 & n370 ;
  assign n372 = ~n317 & ~n371 ;
  assign n374 = ~\u4_pad  & ~n202 ;
  assign n373 = \u4_pad  & n202 ;
  assign n375 = n198 & ~n373 ;
  assign n376 = ~n374 & n375 ;
  assign n393 = \s0_pad  & n350 ;
  assign n394 = ~\j0_pad  & \q5_pad  ;
  assign n395 = \d4_pad  & \e4_pad  ;
  assign n396 = \f4_pad  & n395 ;
  assign n397 = ~n394 & ~n396 ;
  assign n398 = \i4_pad  & ~n397 ;
  assign n399 = ~\j0_pad  & ~\p5_pad  ;
  assign n400 = ~n398 & n399 ;
  assign n401 = \g4_pad  & ~n400 ;
  assign n402 = \p4_pad  & n401 ;
  assign n403 = \q0_pad  & n402 ;
  assign n380 = \p3_pad  & \s3_pad  ;
  assign n381 = \t3_pad  & n380 ;
  assign n382 = n334 & n381 ;
  assign n383 = \m0_pad  & n382 ;
  assign n377 = \n5_pad  & \p0_pad  ;
  assign n378 = \l0_pad  & \l3_pad  ;
  assign n406 = ~n377 & ~n378 ;
  assign n379 = \g4_pad  & \r0_pad  ;
  assign n391 = \l5_pad  & \u0_pad  ;
  assign n407 = ~n379 & ~n391 ;
  assign n404 = \t0_pad  & \v4_pad  ;
  assign n405 = \n0_pad  & \q5_pad  ;
  assign n408 = ~n404 & ~n405 ;
  assign n409 = n407 & n408 ;
  assign n410 = n406 & n409 ;
  assign n411 = ~n383 & n410 ;
  assign n386 = ~\r3_pad  & ~\s3_pad  ;
  assign n387 = ~\t3_pad  & n386 ;
  assign n384 = \n3_pad  & ~\o3_pad  ;
  assign n385 = ~\p3_pad  & ~\q3_pad  ;
  assign n388 = n384 & n385 ;
  assign n389 = n387 & n388 ;
  assign n390 = \k0_pad  & n389 ;
  assign n392 = \o0_pad  & ~n316 ;
  assign n412 = ~n390 & ~n392 ;
  assign n413 = n411 & n412 ;
  assign n414 = ~n403 & n413 ;
  assign n415 = ~n393 & n414 ;
  assign n417 = ~\s1_pad  & ~\t1_pad  ;
  assign n418 = \t1_pad  & ~n252 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = n264 & ~n419 ;
  assign n422 = ~\u1_pad  & n420 ;
  assign n421 = \u1_pad  & ~n420 ;
  assign n423 = n242 & ~n421 ;
  assign n424 = ~n422 & n423 ;
  assign n416 = ~\y2_pad  & ~n242 ;
  assign n425 = ~b_pad & ~n416 ;
  assign n426 = ~n424 & n425 ;
  assign n427 = ~\w2_pad  & ~\x2_pad  ;
  assign n428 = ~\y2_pad  & ~\z2_pad  ;
  assign n429 = n427 & n428 ;
  assign n430 = n277 & ~n429 ;
  assign n431 = ~n278 & ~n430 ;
  assign n432 = \r4_pad  & n346 ;
  assign n433 = n173 & n178 ;
  assign n434 = ~n432 & ~n433 ;
  assign n437 = \r5_pad  & n343 ;
  assign n436 = \q5_pad  & ~\v4_pad  ;
  assign n438 = ~\p5_pad  & ~n436 ;
  assign n439 = ~n437 & n438 ;
  assign n440 = ~\r4_pad  & \s4_pad  ;
  assign n441 = n339 & n440 ;
  assign n442 = ~n311 & n441 ;
  assign n443 = ~n439 & n442 ;
  assign n444 = ~\f0_pad  & ~n443 ;
  assign n445 = \u3_pad  & ~n444 ;
  assign n446 = ~\u3_pad  & n444 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = n434 & ~n447 ;
  assign n435 = ~\l3_pad  & ~n434 ;
  assign n449 = ~z_pad & ~n435 ;
  assign n450 = ~n448 & n449 ;
  assign n452 = \v4_pad  & n373 ;
  assign n451 = ~\v4_pad  & ~n373 ;
  assign n453 = n198 & ~n451 ;
  assign n454 = ~n452 & n453 ;
  assign n455 = n179 & n194 ;
  assign n456 = n175 & n389 ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = n175 & n185 ;
  assign n459 = n382 & n458 ;
  assign n460 = n174 & n179 ;
  assign n461 = ~n433 & ~n460 ;
  assign n462 = ~n459 & n461 ;
  assign n463 = n457 & n462 ;
  assign n468 = \r1_pad  & n279 ;
  assign n469 = n299 & ~n468 ;
  assign n471 = ~\v0_pad  & n469 ;
  assign n464 = \n1_pad  & n228 ;
  assign n465 = ~b_pad & ~n464 ;
  assign n466 = n238 & n299 ;
  assign n467 = n465 & ~n466 ;
  assign n470 = \v0_pad  & ~n469 ;
  assign n472 = n467 & ~n470 ;
  assign n473 = ~n471 & n472 ;
  assign n475 = \s1_pad  & \t1_pad  ;
  assign n476 = \u1_pad  & n475 ;
  assign n477 = ~k_pad & ~n476 ;
  assign n478 = ~n252 & n477 ;
  assign n479 = ~\u1_pad  & n417 ;
  assign n480 = ~k_pad & ~n479 ;
  assign n481 = n252 & n480 ;
  assign n482 = ~n478 & ~n481 ;
  assign n483 = ~n263 & n482 ;
  assign n485 = \v1_pad  & n483 ;
  assign n484 = ~\v1_pad  & ~n483 ;
  assign n486 = n242 & ~n484 ;
  assign n487 = ~n485 & n486 ;
  assign n474 = \z2_pad  & ~n242 ;
  assign n488 = ~b_pad & ~n474 ;
  assign n489 = ~n487 & n488 ;
  assign n490 = \w2_pad  & \x2_pad  ;
  assign n491 = \y2_pad  & \z2_pad  ;
  assign n492 = n490 & n491 ;
  assign n493 = n277 & n492 ;
  assign n495 = ~\g0_pad  & n189 ;
  assign n496 = \u3_pad  & n495 ;
  assign n497 = ~\u3_pad  & ~n495 ;
  assign n498 = ~n444 & ~n497 ;
  assign n499 = ~n496 & n498 ;
  assign n501 = ~\v3_pad  & n499 ;
  assign n500 = \v3_pad  & ~n499 ;
  assign n502 = n434 & ~n500 ;
  assign n503 = ~n501 & n502 ;
  assign n494 = ~\m3_pad  & ~n434 ;
  assign n504 = ~z_pad & ~n494 ;
  assign n505 = ~n503 & n504 ;
  assign n507 = \w4_pad  & n452 ;
  assign n506 = ~\w4_pad  & ~n452 ;
  assign n508 = n198 & ~n506 ;
  assign n509 = ~n507 & n508 ;
  assign n513 = \w0_pad  & n470 ;
  assign n510 = \v0_pad  & n468 ;
  assign n511 = n467 & ~n510 ;
  assign n512 = ~\w0_pad  & ~n470 ;
  assign n514 = n511 & ~n512 ;
  assign n515 = ~n513 & n514 ;
  assign n517 = ~\v1_pad  & ~n480 ;
  assign n518 = n252 & ~n517 ;
  assign n519 = \v1_pad  & ~n477 ;
  assign n520 = ~n252 & ~n519 ;
  assign n521 = ~n518 & ~n520 ;
  assign n522 = ~n263 & n521 ;
  assign n524 = \w1_pad  & n522 ;
  assign n523 = ~\w1_pad  & ~n522 ;
  assign n525 = n242 & ~n523 ;
  assign n526 = ~n524 & n525 ;
  assign n516 = \a3_pad  & ~n242 ;
  assign n527 = ~b_pad & ~n516 ;
  assign n528 = ~n526 & n527 ;
  assign n529 = ~\t2_pad  & ~n292 ;
  assign n530 = ~j_pad & ~n529 ;
  assign n531 = n273 & ~n530 ;
  assign n532 = \t2_pad  & ~n287 ;
  assign n533 = ~j_pad & ~n532 ;
  assign n534 = ~n273 & ~n533 ;
  assign n535 = ~n531 & ~n534 ;
  assign n536 = ~n303 & ~n535 ;
  assign n538 = ~\w2_pad  & ~n536 ;
  assign n537 = \w2_pad  & n536 ;
  assign n539 = n277 & ~n537 ;
  assign n540 = ~n538 & n539 ;
  assign n542 = ~\u3_pad  & ~\v3_pad  ;
  assign n543 = \v3_pad  & ~n495 ;
  assign n544 = ~n542 & ~n543 ;
  assign n545 = n498 & ~n544 ;
  assign n547 = ~\w3_pad  & n545 ;
  assign n546 = \w3_pad  & ~n545 ;
  assign n548 = n434 & ~n546 ;
  assign n549 = ~n547 & n548 ;
  assign n541 = ~\n3_pad  & ~n434 ;
  assign n550 = ~z_pad & ~n541 ;
  assign n551 = ~n549 & n550 ;
  assign n554 = ~\x4_pad  & ~n507 ;
  assign n552 = \w4_pad  & \x4_pad  ;
  assign n553 = n452 & n552 ;
  assign n555 = n198 & ~n553 ;
  assign n556 = ~n554 & n555 ;
  assign n558 = \x0_pad  & n513 ;
  assign n557 = ~\x0_pad  & ~n513 ;
  assign n559 = n511 & ~n557 ;
  assign n560 = ~n558 & n559 ;
  assign n562 = ~\w1_pad  & n517 ;
  assign n563 = n252 & ~n562 ;
  assign n564 = \w1_pad  & n519 ;
  assign n565 = ~n252 & ~n564 ;
  assign n566 = ~n563 & ~n565 ;
  assign n567 = ~n263 & n566 ;
  assign n569 = \x1_pad  & n567 ;
  assign n568 = ~\x1_pad  & ~n567 ;
  assign n570 = n242 & ~n568 ;
  assign n571 = ~n569 & n570 ;
  assign n561 = \b3_pad  & ~n242 ;
  assign n572 = ~b_pad & ~n561 ;
  assign n573 = ~n571 & n572 ;
  assign n575 = ~\w2_pad  & ~n531 ;
  assign n574 = \w2_pad  & ~n534 ;
  assign n576 = ~n303 & ~n574 ;
  assign n577 = ~n575 & n576 ;
  assign n579 = ~\x2_pad  & ~n577 ;
  assign n578 = \x2_pad  & n577 ;
  assign n580 = n277 & ~n578 ;
  assign n581 = ~n579 & n580 ;
  assign n583 = ~\w3_pad  & n542 ;
  assign n584 = ~\i0_pad  & n495 ;
  assign n585 = ~n583 & n584 ;
  assign n586 = \u3_pad  & \v3_pad  ;
  assign n587 = \w3_pad  & n586 ;
  assign n588 = ~\i0_pad  & ~n587 ;
  assign n589 = ~n495 & n588 ;
  assign n590 = ~n444 & ~n589 ;
  assign n591 = ~n585 & n590 ;
  assign n593 = \x3_pad  & n591 ;
  assign n592 = ~\x3_pad  & ~n591 ;
  assign n594 = n434 & ~n592 ;
  assign n595 = ~n593 & n594 ;
  assign n582 = \o3_pad  & ~n434 ;
  assign n596 = ~z_pad & ~n582 ;
  assign n597 = ~n595 & n596 ;
  assign n599 = \y4_pad  & n553 ;
  assign n598 = ~\y4_pad  & ~n553 ;
  assign n600 = n198 & ~n598 ;
  assign n601 = ~n599 & n600 ;
  assign n603 = \c3_pad  & \d3_pad  ;
  assign n604 = \e3_pad  & n603 ;
  assign n605 = n247 & n604 ;
  assign n606 = n279 & ~n605 ;
  assign n602 = n247 & n276 ;
  assign n607 = ~n229 & ~n602 ;
  assign n608 = ~n606 & n607 ;
  assign n610 = \y0_pad  & n558 ;
  assign n609 = ~\y0_pad  & ~n558 ;
  assign n611 = n511 & ~n609 ;
  assign n612 = ~n610 & n611 ;
  assign n617 = \x1_pad  & n564 ;
  assign n618 = ~k_pad & ~n617 ;
  assign n619 = ~n252 & n618 ;
  assign n614 = ~\x1_pad  & n562 ;
  assign n615 = ~k_pad & ~n614 ;
  assign n616 = n252 & n615 ;
  assign n620 = ~n263 & ~n616 ;
  assign n621 = ~n619 & n620 ;
  assign n623 = ~\y1_pad  & n621 ;
  assign n622 = \y1_pad  & ~n621 ;
  assign n624 = n242 & ~n622 ;
  assign n625 = ~n623 & n624 ;
  assign n613 = ~\c3_pad  & ~n242 ;
  assign n626 = ~b_pad & ~n613 ;
  assign n627 = ~n625 & n626 ;
  assign n628 = n427 & n531 ;
  assign n629 = n490 & n534 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = ~n303 & ~n630 ;
  assign n633 = ~\y2_pad  & ~n631 ;
  assign n632 = \y2_pad  & n631 ;
  assign n634 = n277 & ~n632 ;
  assign n635 = ~n633 & n634 ;
  assign n640 = \x3_pad  & ~n588 ;
  assign n641 = ~n495 & ~n640 ;
  assign n637 = ~\i0_pad  & ~n583 ;
  assign n638 = ~\x3_pad  & ~n637 ;
  assign n639 = n495 & ~n638 ;
  assign n642 = ~n444 & ~n639 ;
  assign n643 = ~n641 & n642 ;
  assign n645 = \y3_pad  & n643 ;
  assign n644 = ~\y3_pad  & ~n643 ;
  assign n646 = n434 & ~n644 ;
  assign n647 = ~n645 & n646 ;
  assign n636 = \p3_pad  & ~n434 ;
  assign n648 = ~z_pad & ~n636 ;
  assign n649 = ~n647 & n648 ;
  assign n651 = \z4_pad  & n599 ;
  assign n650 = ~\z4_pad  & ~n599 ;
  assign n652 = n198 & ~n650 ;
  assign n653 = ~n651 & n652 ;
  assign n656 = ~\z0_pad  & ~n610 ;
  assign n654 = \y0_pad  & \z0_pad  ;
  assign n655 = n558 & n654 ;
  assign n657 = n511 & ~n655 ;
  assign n658 = ~n656 & n657 ;
  assign n660 = \y1_pad  & ~n252 ;
  assign n661 = ~n618 & n660 ;
  assign n662 = ~\y1_pad  & n252 ;
  assign n663 = ~n615 & n662 ;
  assign n664 = ~n661 & ~n663 ;
  assign n665 = ~n263 & ~n664 ;
  assign n667 = \z1_pad  & n665 ;
  assign n666 = ~\z1_pad  & ~n665 ;
  assign n668 = n242 & ~n666 ;
  assign n669 = ~n667 & n668 ;
  assign n659 = \d3_pad  & ~n242 ;
  assign n670 = ~b_pad & ~n659 ;
  assign n671 = ~n669 & n670 ;
  assign n673 = \y2_pad  & ~n629 ;
  assign n672 = ~\y2_pad  & ~n628 ;
  assign n674 = ~n303 & ~n672 ;
  assign n675 = ~n673 & n674 ;
  assign n677 = \z2_pad  & n675 ;
  assign n676 = ~\z2_pad  & ~n675 ;
  assign n678 = n277 & ~n676 ;
  assign n679 = ~n677 & n678 ;
  assign n680 = ~n278 & ~n679 ;
  assign n684 = \y3_pad  & n640 ;
  assign n685 = ~n495 & ~n684 ;
  assign n682 = ~\y3_pad  & n638 ;
  assign n683 = n495 & ~n682 ;
  assign n686 = ~n444 & ~n683 ;
  assign n687 = ~n685 & n686 ;
  assign n689 = \z3_pad  & n687 ;
  assign n688 = ~\z3_pad  & ~n687 ;
  assign n690 = n434 & ~n688 ;
  assign n691 = ~n689 & n690 ;
  assign n681 = \q3_pad  & ~n434 ;
  assign n692 = ~z_pad & ~n681 ;
  assign n693 = ~n691 & n692 ;
  assign n695 = \a1_pad  & n655 ;
  assign n694 = ~\a1_pad  & ~n655 ;
  assign n696 = n511 & ~n694 ;
  assign n697 = ~n695 & n696 ;
  assign n700 = \z1_pad  & ~n661 ;
  assign n699 = ~\z1_pad  & ~n663 ;
  assign n701 = ~n263 & ~n699 ;
  assign n702 = ~n700 & n701 ;
  assign n704 = \a2_pad  & n702 ;
  assign n703 = ~\a2_pad  & ~n702 ;
  assign n705 = n242 & ~n703 ;
  assign n706 = ~n704 & n705 ;
  assign n698 = \e3_pad  & ~n242 ;
  assign n707 = ~b_pad & ~n698 ;
  assign n708 = ~n706 & n707 ;
  assign n711 = \v2_pad  & ~n533 ;
  assign n712 = ~n273 & ~n711 ;
  assign n709 = \u2_pad  & ~n530 ;
  assign n710 = n273 & ~n709 ;
  assign n713 = ~n303 & ~n710 ;
  assign n714 = ~n712 & n713 ;
  assign n716 = \a3_pad  & n714 ;
  assign n715 = ~\a3_pad  & ~n714 ;
  assign n717 = n277 & ~n715 ;
  assign n718 = ~n716 & n717 ;
  assign n719 = ~n278 & ~n718 ;
  assign n723 = \z3_pad  & n684 ;
  assign n724 = ~\i0_pad  & ~n495 ;
  assign n725 = ~n723 & n724 ;
  assign n721 = ~\z3_pad  & n682 ;
  assign n722 = n584 & ~n721 ;
  assign n726 = ~n444 & ~n722 ;
  assign n727 = ~n725 & n726 ;
  assign n728 = ~\a4_pad  & ~n727 ;
  assign n729 = \a4_pad  & n727 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = n434 & ~n730 ;
  assign n720 = ~\r3_pad  & ~n434 ;
  assign n732 = ~z_pad & ~n720 ;
  assign n733 = ~n731 & n732 ;
  assign n735 = \b1_pad  & n695 ;
  assign n734 = ~\b1_pad  & ~n695 ;
  assign n736 = n511 & ~n734 ;
  assign n737 = ~n735 & n736 ;
  assign n738 = \b2_pad  & ~b_pad ;
  assign n739 = ~\a3_pad  & n709 ;
  assign n740 = ~j_pad & ~n739 ;
  assign n741 = n273 & n740 ;
  assign n742 = \a3_pad  & n711 ;
  assign n743 = ~j_pad & ~n273 ;
  assign n744 = ~n742 & n743 ;
  assign n745 = ~n303 & ~n744 ;
  assign n746 = ~n741 & n745 ;
  assign n748 = \b3_pad  & n746 ;
  assign n747 = ~\b3_pad  & ~n746 ;
  assign n749 = n277 & ~n747 ;
  assign n750 = ~n748 & n749 ;
  assign n751 = ~n278 & ~n750 ;
  assign n753 = ~\a4_pad  & ~n495 ;
  assign n754 = \a4_pad  & n495 ;
  assign n755 = ~n753 & ~n754 ;
  assign n756 = n727 & n755 ;
  assign n757 = \b4_pad  & ~n756 ;
  assign n758 = ~\b4_pad  & n756 ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = n434 & ~n759 ;
  assign n752 = \s3_pad  & ~n434 ;
  assign n761 = ~z_pad & ~n752 ;
  assign n762 = ~n760 & n761 ;
  assign n764 = \c1_pad  & n735 ;
  assign n763 = ~\c1_pad  & ~n735 ;
  assign n765 = n511 & ~n763 ;
  assign n766 = ~n764 & n765 ;
  assign n767 = ~\b2_pad  & ~\c2_pad  ;
  assign n768 = \b2_pad  & \c2_pad  ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = ~b_pad & ~n769 ;
  assign n771 = ~\b3_pad  & ~n740 ;
  assign n772 = n273 & ~n771 ;
  assign n773 = ~\b3_pad  & ~n273 ;
  assign n774 = n745 & ~n773 ;
  assign n775 = ~n772 & n774 ;
  assign n777 = \c3_pad  & n775 ;
  assign n776 = ~\c3_pad  & ~n775 ;
  assign n778 = n277 & ~n776 ;
  assign n779 = ~n777 & n778 ;
  assign n781 = ~\b4_pad  & ~n495 ;
  assign n782 = \b4_pad  & n495 ;
  assign n783 = ~n781 & ~n782 ;
  assign n784 = n756 & n783 ;
  assign n786 = \c4_pad  & n784 ;
  assign n785 = ~\c4_pad  & ~n784 ;
  assign n787 = n434 & ~n785 ;
  assign n788 = ~n786 & n787 ;
  assign n780 = \t3_pad  & ~n434 ;
  assign n789 = ~z_pad & ~n780 ;
  assign n790 = ~n788 & n789 ;
  assign n791 = \d5_pad  & ~n185 ;
  assign n792 = n181 & n791 ;
  assign n793 = ~n191 & ~n792 ;
  assign n795 = n175 & ~n459 ;
  assign n794 = n185 & n315 ;
  assign n796 = ~n433 & ~n794 ;
  assign n797 = ~n795 & n796 ;
  assign n799 = \d1_pad  & n764 ;
  assign n798 = ~\d1_pad  & ~n764 ;
  assign n800 = n511 & ~n798 ;
  assign n801 = ~n799 & n800 ;
  assign n802 = \d2_pad  & n768 ;
  assign n803 = ~\d2_pad  & ~n768 ;
  assign n804 = ~n802 & ~n803 ;
  assign n805 = ~b_pad & ~n804 ;
  assign n806 = ~\c3_pad  & ~n273 ;
  assign n807 = \c3_pad  & n273 ;
  assign n808 = ~n806 & ~n807 ;
  assign n809 = n775 & n808 ;
  assign n811 = \d3_pad  & n809 ;
  assign n810 = ~\d3_pad  & ~n809 ;
  assign n812 = n277 & ~n810 ;
  assign n813 = ~n811 & n812 ;
  assign n814 = ~n278 & ~n813 ;
  assign n815 = \d4_pad  & ~z_pad ;
  assign n816 = \e5_pad  & ~n183 ;
  assign n817 = n181 & n816 ;
  assign n818 = ~n187 & ~n817 ;
  assign n819 = ~l_pad & \q1_pad  ;
  assign n820 = ~n802 & ~n819 ;
  assign n821 = \g2_pad  & ~n820 ;
  assign n822 = ~l_pad & ~\p1_pad  ;
  assign n823 = ~n821 & n822 ;
  assign n824 = \e2_pad  & ~n823 ;
  assign n825 = \n2_pad  & n824 ;
  assign n826 = ~n464 & ~n825 ;
  assign n828 = ~\e2_pad  & n823 ;
  assign n829 = ~n824 & ~n828 ;
  assign n830 = n826 & n829 ;
  assign n827 = \s1_pad  & ~n826 ;
  assign n831 = ~b_pad & ~n827 ;
  assign n832 = ~n830 & n831 ;
  assign n833 = ~\c3_pad  & ~\d3_pad  ;
  assign n834 = n771 & n833 ;
  assign n835 = n273 & ~n834 ;
  assign n836 = ~n273 & ~n603 ;
  assign n837 = n774 & ~n836 ;
  assign n838 = ~n835 & n837 ;
  assign n840 = \e3_pad  & n838 ;
  assign n839 = ~\e3_pad  & ~n838 ;
  assign n841 = n277 & ~n839 ;
  assign n842 = ~n840 & n841 ;
  assign n843 = ~n278 & ~n842 ;
  assign n844 = ~\d4_pad  & ~\e4_pad  ;
  assign n845 = ~n395 & ~n844 ;
  assign n846 = ~z_pad & ~n845 ;
  assign n848 = ~\h5_pad  & n402 ;
  assign n847 = \h5_pad  & ~n402 ;
  assign n849 = ~n178 & ~n847 ;
  assign n850 = ~n848 & n849 ;
  assign n851 = ~z_pad & ~n850 ;
  assign n852 = ~\h5_pad  & n851 ;
  assign n853 = ~\p10_pad  & n852 ;
  assign n854 = ~\f5_pad  & ~n853 ;
  assign n855 = \f5_pad  & n852 ;
  assign n856 = ~n178 & ~n855 ;
  assign n857 = ~n854 & n856 ;
  assign n858 = ~z_pad & ~n857 ;
  assign n860 = \f2_pad  & n824 ;
  assign n861 = ~\f2_pad  & ~n824 ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = n826 & n862 ;
  assign n859 = \t1_pad  & ~n826 ;
  assign n864 = ~b_pad & ~n859 ;
  assign n865 = ~n863 & n864 ;
  assign n867 = ~\f3_pad  & n350 ;
  assign n866 = \f3_pad  & ~n350 ;
  assign n868 = n316 & ~n866 ;
  assign n869 = ~n867 & n868 ;
  assign n870 = ~\f4_pad  & ~n395 ;
  assign n871 = ~n396 & ~n870 ;
  assign n872 = ~z_pad & ~n871 ;
  assign n873 = \p10_pad  & ~n852 ;
  assign n874 = n856 & ~n873 ;
  assign n875 = ~z_pad & ~n874 ;
  assign n876 = ~\g2_pad  & n820 ;
  assign n877 = ~n821 & ~n876 ;
  assign n878 = ~b_pad & ~n877 ;
  assign n880 = \f3_pad  & n313 ;
  assign n879 = ~\f3_pad  & ~n313 ;
  assign n881 = ~n350 & ~n879 ;
  assign n882 = ~n880 & n881 ;
  assign n884 = ~\g3_pad  & ~n882 ;
  assign n883 = \g3_pad  & n882 ;
  assign n885 = n316 & ~n883 ;
  assign n886 = ~n884 & n885 ;
  assign n887 = ~n180 & ~n402 ;
  assign n889 = ~\g4_pad  & n400 ;
  assign n890 = ~n401 & ~n889 ;
  assign n891 = n887 & n890 ;
  assign n888 = \u3_pad  & ~n887 ;
  assign n892 = ~z_pad & ~n888 ;
  assign n893 = ~n891 & n892 ;
  assign n894 = \h1_pad  & ~n247 ;
  assign n895 = n465 & n894 ;
  assign n896 = ~n297 & ~n895 ;
  assign n897 = ~\h2_pad  & ~n860 ;
  assign n898 = \f2_pad  & \h2_pad  ;
  assign n899 = n824 & n898 ;
  assign n900 = n826 & ~n899 ;
  assign n901 = ~n897 & n900 ;
  assign n902 = \u1_pad  & ~n826 ;
  assign n903 = ~b_pad & ~n902 ;
  assign n904 = ~n901 & n903 ;
  assign n906 = ~n313 & n352 ;
  assign n905 = n313 & n321 ;
  assign n907 = ~n350 & ~n905 ;
  assign n908 = ~n906 & n907 ;
  assign n910 = ~\h3_pad  & ~n908 ;
  assign n909 = \h3_pad  & n908 ;
  assign n911 = n316 & ~n909 ;
  assign n912 = ~n910 & n911 ;
  assign n914 = \h4_pad  & n401 ;
  assign n915 = ~\h4_pad  & ~n401 ;
  assign n916 = ~n914 & ~n915 ;
  assign n917 = n887 & n916 ;
  assign n913 = \v3_pad  & ~n887 ;
  assign n918 = ~z_pad & ~n913 ;
  assign n919 = ~n917 & n918 ;
  assign n920 = \i1_pad  & ~n245 ;
  assign n921 = n465 & n920 ;
  assign n922 = ~n249 & ~n921 ;
  assign n925 = ~\i2_pad  & ~n899 ;
  assign n924 = \i2_pad  & n899 ;
  assign n926 = n826 & ~n924 ;
  assign n927 = ~n925 & n926 ;
  assign n923 = \v1_pad  & ~n826 ;
  assign n928 = ~b_pad & ~n923 ;
  assign n929 = ~n927 & n928 ;
  assign n931 = ~n313 & n354 ;
  assign n930 = n313 & n325 ;
  assign n932 = ~n350 & ~n930 ;
  assign n933 = ~n931 & n932 ;
  assign n935 = \i3_pad  & n933 ;
  assign n934 = ~\i3_pad  & ~n933 ;
  assign n936 = n316 & ~n934 ;
  assign n937 = ~n935 & n936 ;
  assign n938 = ~n317 & ~n937 ;
  assign n939 = ~\i4_pad  & n397 ;
  assign n940 = ~n398 & ~n939 ;
  assign n941 = ~z_pad & ~n940 ;
  assign n944 = \j5_pad  & n175 ;
  assign n942 = ~z_pad & ~n336 ;
  assign n943 = ~\j5_pad  & ~n175 ;
  assign n945 = n942 & ~n943 ;
  assign n946 = ~n944 & n945 ;
  assign n948 = ~\r6_pad  & ~n825 ;
  assign n947 = \r6_pad  & n825 ;
  assign n949 = ~b_pad & ~n947 ;
  assign n950 = ~n948 & n949 ;
  assign n951 = ~n228 & ~n950 ;
  assign n953 = ~\j2_pad  & ~n924 ;
  assign n954 = \i2_pad  & \j2_pad  ;
  assign n955 = n898 & n954 ;
  assign n956 = n824 & n955 ;
  assign n957 = n826 & ~n956 ;
  assign n958 = ~n953 & n957 ;
  assign n952 = \w1_pad  & ~n826 ;
  assign n959 = ~b_pad & ~n952 ;
  assign n960 = ~n958 & n959 ;
  assign n961 = ~\l3_pad  & ~\m3_pad  ;
  assign n962 = ~\n3_pad  & ~\o3_pad  ;
  assign n963 = n961 & n962 ;
  assign n964 = n316 & ~n963 ;
  assign n965 = ~n317 & ~n964 ;
  assign n966 = ~\j4_pad  & ~n914 ;
  assign n967 = \h4_pad  & \j4_pad  ;
  assign n968 = n401 & n967 ;
  assign n969 = n887 & ~n968 ;
  assign n970 = ~n966 & n969 ;
  assign n971 = \w3_pad  & ~n887 ;
  assign n972 = ~z_pad & ~n971 ;
  assign n973 = ~n970 & n972 ;
  assign n975 = \k5_pad  & n944 ;
  assign n974 = ~\k5_pad  & ~n944 ;
  assign n976 = n942 & ~n974 ;
  assign n977 = ~n975 & n976 ;
  assign n979 = ~l_pad & ~n956 ;
  assign n981 = ~\k2_pad  & n979 ;
  assign n980 = \k2_pad  & ~n979 ;
  assign n982 = n826 & ~n980 ;
  assign n983 = ~n981 & n982 ;
  assign n978 = \x1_pad  & ~n826 ;
  assign n984 = ~b_pad & ~n978 ;
  assign n985 = ~n983 & n984 ;
  assign n986 = \l3_pad  & \m3_pad  ;
  assign n987 = \n3_pad  & \o3_pad  ;
  assign n988 = n986 & n987 ;
  assign n989 = n316 & n988 ;
  assign n992 = ~\k4_pad  & ~n968 ;
  assign n991 = \k4_pad  & n968 ;
  assign n993 = n887 & ~n991 ;
  assign n994 = ~n992 & n993 ;
  assign n990 = \x3_pad  & ~n887 ;
  assign n995 = ~z_pad & ~n990 ;
  assign n996 = ~n994 & n995 ;
  assign n1007 = \o2_pad  & s_pad ;
  assign n1005 = r_pad & \u1_pad  ;
  assign n1006 = o_pad & \t2_pad  ;
  assign n1012 = ~n1005 & ~n1006 ;
  assign n1013 = ~n1007 & n1012 ;
  assign n1001 = q_pad & \x1_pad  ;
  assign n1002 = \j2_pad  & t_pad ;
  assign n1010 = ~n1001 & ~n1002 ;
  assign n1003 = \a3_pad  & n_pad ;
  assign n1004 = \e3_pad  & m_pad ;
  assign n1011 = ~n1003 & ~n1004 ;
  assign n1014 = n1010 & n1011 ;
  assign n997 = \a2_pad  & p_pad ;
  assign n998 = w_pad & \y0_pad  ;
  assign n1008 = ~n997 & ~n998 ;
  assign n999 = \d1_pad  & v_pad ;
  assign n1000 = \g2_pad  & u_pad ;
  assign n1009 = ~n999 & ~n1000 ;
  assign n1015 = n1008 & n1009 ;
  assign n1016 = n1014 & n1015 ;
  assign n1017 = n1013 & n1016 ;
  assign n1020 = \l2_pad  & n980 ;
  assign n1019 = ~\l2_pad  & ~n980 ;
  assign n1021 = n826 & ~n1019 ;
  assign n1022 = ~n1020 & n1021 ;
  assign n1018 = \y1_pad  & ~n826 ;
  assign n1023 = ~b_pad & ~n1018 ;
  assign n1024 = ~n1022 & n1023 ;
  assign n1026 = n313 & n327 ;
  assign n1025 = ~n313 & n356 ;
  assign n1027 = ~n350 & ~n1025 ;
  assign n1028 = ~n1026 & n1027 ;
  assign n1030 = \l3_pad  & n1028 ;
  assign n1029 = ~\l3_pad  & ~n1028 ;
  assign n1031 = n316 & ~n1029 ;
  assign n1032 = ~n1030 & n1031 ;
  assign n1034 = ~\l4_pad  & ~n991 ;
  assign n1035 = \k4_pad  & \l4_pad  ;
  assign n1036 = n967 & n1035 ;
  assign n1037 = n401 & n1036 ;
  assign n1038 = n887 & ~n1037 ;
  assign n1039 = ~n1034 & n1038 ;
  assign n1033 = \y3_pad  & ~n887 ;
  assign n1040 = ~z_pad & ~n1033 ;
  assign n1041 = ~n1039 & n1040 ;
  assign n1042 = \r5_pad  & ~n599 ;
  assign n1043 = \z4_pad  & ~n1042 ;
  assign n1044 = ~\a0_pad  & ~n1043 ;
  assign n1045 = n195 & ~n1044 ;
  assign n1047 = n175 & ~n185 ;
  assign n1048 = ~n389 & n1047 ;
  assign n1046 = \m5_pad  & \n5_pad  ;
  assign n1049 = ~n315 & ~n1046 ;
  assign n1050 = ~n1048 & n1049 ;
  assign n1051 = n457 & n1050 ;
  assign n1052 = ~n1045 & n1051 ;
  assign n1053 = ~z_pad & ~n1052 ;
  assign n1064 = \m2_pad  & s_pad ;
  assign n1062 = q_pad & \w1_pad  ;
  assign n1063 = o_pad & \s2_pad  ;
  assign n1069 = ~n1062 & ~n1063 ;
  assign n1070 = ~n1064 & n1069 ;
  assign n1058 = r_pad & \t1_pad  ;
  assign n1059 = \i2_pad  & t_pad ;
  assign n1067 = ~n1058 & ~n1059 ;
  assign n1060 = n_pad & \z2_pad  ;
  assign n1061 = \d3_pad  & m_pad ;
  assign n1068 = ~n1060 & ~n1061 ;
  assign n1071 = n1067 & n1068 ;
  assign n1054 = p_pad & \z1_pad  ;
  assign n1055 = w_pad & \x0_pad  ;
  assign n1065 = ~n1054 & ~n1055 ;
  assign n1056 = \c1_pad  & v_pad ;
  assign n1057 = \d2_pad  & u_pad ;
  assign n1066 = ~n1056 & ~n1057 ;
  assign n1072 = n1065 & n1066 ;
  assign n1073 = n1071 & n1072 ;
  assign n1074 = n1070 & n1073 ;
  assign n1075 = \r1_pad  & ~n764 ;
  assign n1076 = \d1_pad  & ~n1075 ;
  assign n1077 = ~c_pad & ~n1076 ;
  assign n1078 = n238 & ~n1077 ;
  assign n1081 = ~\e3_pad  & \y2_pad  ;
  assign n1082 = ~\z2_pad  & n1081 ;
  assign n1080 = ~\a3_pad  & ~\b3_pad  ;
  assign n1083 = n833 & n1080 ;
  assign n1084 = n1082 & n1083 ;
  assign n1089 = ~n247 & n279 ;
  assign n1090 = ~n1084 & n1089 ;
  assign n1085 = n279 & n1084 ;
  assign n1086 = ~b_pad & \n1_pad  ;
  assign n1087 = n237 & n1086 ;
  assign n1088 = ~n1085 & ~n1087 ;
  assign n1079 = \m1_pad  & \n1_pad  ;
  assign n1091 = ~n276 & ~n1079 ;
  assign n1092 = n1088 & n1091 ;
  assign n1093 = ~n1090 & n1092 ;
  assign n1094 = ~n1078 & n1093 ;
  assign n1095 = ~b_pad & ~n1094 ;
  assign n1098 = \m2_pad  & n1020 ;
  assign n1097 = ~\m2_pad  & ~n1020 ;
  assign n1099 = n826 & ~n1097 ;
  assign n1100 = ~n1098 & n1099 ;
  assign n1096 = \z1_pad  & ~n826 ;
  assign n1101 = ~b_pad & ~n1096 ;
  assign n1102 = ~n1100 & n1101 ;
  assign n1103 = ~\l3_pad  & ~n313 ;
  assign n1104 = \l3_pad  & n313 ;
  assign n1105 = ~n1103 & ~n1104 ;
  assign n1106 = n1028 & n1105 ;
  assign n1108 = \m3_pad  & n1106 ;
  assign n1107 = ~\m3_pad  & ~n1106 ;
  assign n1109 = n316 & ~n1107 ;
  assign n1110 = ~n1108 & n1109 ;
  assign n1112 = ~\j0_pad  & ~n1037 ;
  assign n1114 = ~\m4_pad  & n1112 ;
  assign n1113 = \m4_pad  & ~n1112 ;
  assign n1115 = n887 & ~n1113 ;
  assign n1116 = ~n1114 & n1115 ;
  assign n1111 = \z3_pad  & ~n887 ;
  assign n1117 = ~z_pad & ~n1111 ;
  assign n1118 = ~n1116 & n1117 ;
  assign n1129 = \l2_pad  & s_pad ;
  assign n1127 = q_pad & \v1_pad  ;
  assign n1128 = o_pad & \r2_pad  ;
  assign n1134 = ~n1127 & ~n1128 ;
  assign n1135 = ~n1129 & n1134 ;
  assign n1123 = r_pad & \s1_pad  ;
  assign n1124 = \h2_pad  & t_pad ;
  assign n1132 = ~n1123 & ~n1124 ;
  assign n1125 = n_pad & \y2_pad  ;
  assign n1126 = \c3_pad  & m_pad ;
  assign n1133 = ~n1125 & ~n1126 ;
  assign n1136 = n1132 & n1133 ;
  assign n1119 = p_pad & \y1_pad  ;
  assign n1120 = \w0_pad  & w_pad ;
  assign n1130 = ~n1119 & ~n1120 ;
  assign n1121 = \b1_pad  & v_pad ;
  assign n1122 = \c2_pad  & u_pad ;
  assign n1131 = ~n1121 & ~n1122 ;
  assign n1137 = n1130 & n1131 ;
  assign n1138 = n1136 & n1137 ;
  assign n1139 = n1135 & n1138 ;
  assign n1140 = ~b_pad & ~n826 ;
  assign n1141 = \k2_pad  & \l2_pad  ;
  assign n1142 = \m2_pad  & \o2_pad  ;
  assign n1143 = n1141 & n1142 ;
  assign n1144 = n955 & n1143 ;
  assign n1145 = ~n1140 & n1144 ;
  assign n1146 = ~\m3_pad  & ~n313 ;
  assign n1147 = \m3_pad  & n313 ;
  assign n1148 = ~n1146 & ~n1147 ;
  assign n1149 = n1106 & n1148 ;
  assign n1151 = \n3_pad  & n1149 ;
  assign n1150 = ~\n3_pad  & ~n1149 ;
  assign n1152 = n316 & ~n1150 ;
  assign n1153 = ~n1151 & n1152 ;
  assign n1156 = \n4_pad  & n1113 ;
  assign n1155 = ~\n4_pad  & ~n1113 ;
  assign n1157 = n887 & ~n1155 ;
  assign n1158 = ~n1156 & n1157 ;
  assign n1154 = \a4_pad  & ~n887 ;
  assign n1159 = ~z_pad & ~n1154 ;
  assign n1160 = ~n1158 & n1159 ;
  assign n1171 = \k2_pad  & s_pad ;
  assign n1169 = \m1_pad  & r_pad ;
  assign n1170 = o_pad & \q2_pad  ;
  assign n1176 = ~n1169 & ~n1170 ;
  assign n1177 = ~n1171 & n1176 ;
  assign n1165 = q_pad & \r1_pad  ;
  assign n1166 = \f2_pad  & t_pad ;
  assign n1174 = ~n1165 & ~n1166 ;
  assign n1167 = n_pad & \x2_pad  ;
  assign n1168 = \b3_pad  & m_pad ;
  assign n1175 = ~n1167 & ~n1168 ;
  assign n1178 = n1174 & n1175 ;
  assign n1161 = \p1_pad  & p_pad ;
  assign n1162 = \v0_pad  & w_pad ;
  assign n1172 = ~n1161 & ~n1162 ;
  assign n1163 = \a1_pad  & v_pad ;
  assign n1164 = \b2_pad  & u_pad ;
  assign n1173 = ~n1163 & ~n1164 ;
  assign n1179 = n1172 & n1173 ;
  assign n1180 = n1178 & n1179 ;
  assign n1181 = n1177 & n1180 ;
  assign n1184 = ~\o2_pad  & ~n1098 ;
  assign n1183 = ~n979 & n1143 ;
  assign n1185 = n826 & ~n1183 ;
  assign n1186 = ~n1184 & n1185 ;
  assign n1182 = \a2_pad  & ~n826 ;
  assign n1187 = ~b_pad & ~n1182 ;
  assign n1188 = ~n1186 & n1187 ;
  assign n1189 = ~\n3_pad  & ~n313 ;
  assign n1190 = \n3_pad  & n313 ;
  assign n1191 = ~n1189 & ~n1190 ;
  assign n1192 = n1149 & n1191 ;
  assign n1194 = \o3_pad  & n1192 ;
  assign n1193 = ~\o3_pad  & ~n1192 ;
  assign n1195 = n316 & ~n1193 ;
  assign n1196 = ~n1194 & n1195 ;
  assign n1197 = ~n317 & ~n1196 ;
  assign n1200 = \o4_pad  & n1156 ;
  assign n1199 = ~\o4_pad  & ~n1156 ;
  assign n1201 = n887 & ~n1199 ;
  assign n1202 = ~n1200 & n1201 ;
  assign n1198 = \b4_pad  & ~n887 ;
  assign n1203 = ~z_pad & ~n1198 ;
  assign n1204 = ~n1202 & n1203 ;
  assign n1207 = ~\b0_pad  & ~n455 ;
  assign n1205 = ~\c0_pad  & ~n460 ;
  assign n1216 = \p5_pad  & n1205 ;
  assign n1217 = n1207 & n1216 ;
  assign n1210 = ~\p5_pad  & ~\q5_pad  ;
  assign n1211 = ~\r5_pad  & ~n1210 ;
  assign n1212 = \r5_pad  & n1210 ;
  assign n1213 = ~n1211 & ~n1212 ;
  assign n1209 = \p5_pad  & \q5_pad  ;
  assign n1214 = ~z_pad & ~n1209 ;
  assign n1215 = ~n1213 & n1214 ;
  assign n1206 = \r5_pad  & ~n1205 ;
  assign n1208 = \q5_pad  & ~n1207 ;
  assign n1218 = ~n1206 & ~n1208 ;
  assign n1219 = n1215 & n1218 ;
  assign n1220 = ~n1217 & n1219 ;
  assign n1228 = u_pad & n303 ;
  assign n1229 = s_pad & n825 ;
  assign n1226 = q_pad & ~n277 ;
  assign n1230 = m_pad & n1084 ;
  assign n1231 = o_pad & n604 ;
  assign n1221 = p_pad & \q1_pad  ;
  assign n1222 = \e2_pad  & t_pad ;
  assign n1232 = ~n1221 & ~n1222 ;
  assign n1223 = \l1_pad  & w_pad ;
  assign n1224 = v_pad & \z0_pad  ;
  assign n1233 = ~n1223 & ~n1224 ;
  assign n1225 = n_pad & \w2_pad  ;
  assign n1227 = \n1_pad  & r_pad ;
  assign n1234 = ~n1225 & ~n1227 ;
  assign n1235 = n1233 & n1234 ;
  assign n1236 = n1232 & n1235 ;
  assign n1237 = ~n1231 & n1236 ;
  assign n1238 = ~n1230 & n1237 ;
  assign n1239 = ~n1226 & n1238 ;
  assign n1240 = ~n1229 & n1239 ;
  assign n1241 = ~n1228 & n1240 ;
  assign n1245 = ~d_pad & ~n1087 ;
  assign n1242 = n227 & n1079 ;
  assign n1243 = ~e_pad & ~n1242 ;
  assign n1254 = \p1_pad  & n1243 ;
  assign n1255 = n1245 & n1254 ;
  assign n1248 = ~\p1_pad  & ~\q1_pad  ;
  assign n1249 = ~\r1_pad  & ~n1248 ;
  assign n1250 = \r1_pad  & n1248 ;
  assign n1251 = ~n1249 & ~n1250 ;
  assign n1247 = \p1_pad  & \q1_pad  ;
  assign n1252 = ~b_pad & ~n1247 ;
  assign n1253 = ~n1251 & n1252 ;
  assign n1244 = \r1_pad  & ~n1243 ;
  assign n1246 = \q1_pad  & ~n1245 ;
  assign n1256 = ~n1244 & ~n1246 ;
  assign n1257 = n1253 & n1256 ;
  assign n1258 = ~n1255 & n1257 ;
  assign n1259 = \p2_pad  & ~n947 ;
  assign n1260 = ~\l6_pad  & n947 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1263 = n313 & ~n328 ;
  assign n1262 = ~n313 & ~n357 ;
  assign n1264 = ~n350 & ~n1262 ;
  assign n1265 = ~n1263 & n1264 ;
  assign n1267 = \p3_pad  & n1265 ;
  assign n1266 = ~\p3_pad  & ~n1265 ;
  assign n1268 = n316 & ~n1266 ;
  assign n1269 = ~n1267 & n1268 ;
  assign n1270 = ~n317 & ~n1269 ;
  assign n1271 = ~z_pad & ~n887 ;
  assign n1272 = \m4_pad  & \n4_pad  ;
  assign n1273 = \o4_pad  & \q4_pad  ;
  assign n1274 = n1272 & n1273 ;
  assign n1275 = n1036 & n1274 ;
  assign n1276 = ~n1271 & n1275 ;
  assign n1279 = \q5_pad  & n1205 ;
  assign n1280 = n1207 & n1279 ;
  assign n1277 = \r5_pad  & ~n1207 ;
  assign n1278 = \p5_pad  & ~n1205 ;
  assign n1281 = ~n1277 & ~n1278 ;
  assign n1282 = ~n1280 & n1281 ;
  assign n1283 = n1215 & ~n1282 ;
  assign n1284 = n279 & n605 ;
  assign n1285 = ~n229 & ~n1242 ;
  assign n1286 = ~n1284 & n1285 ;
  assign n1287 = n1088 & n1286 ;
  assign n1298 = \q0_pad  & \q4_pad  ;
  assign n1296 = \p0_pad  & \w3_pad  ;
  assign n1297 = \i3_pad  & \m0_pad  ;
  assign n1303 = ~n1296 & ~n1297 ;
  assign n1304 = ~n1298 & n1303 ;
  assign n1292 = \o0_pad  & \z3_pad  ;
  assign n1293 = \l4_pad  & \r0_pad  ;
  assign n1301 = ~n1292 & ~n1293 ;
  assign n1294 = \k0_pad  & \t3_pad  ;
  assign n1295 = \l0_pad  & \p3_pad  ;
  assign n1302 = ~n1294 & ~n1295 ;
  assign n1305 = n1301 & n1302 ;
  assign n1288 = \c4_pad  & \n0_pad  ;
  assign n1289 = \u0_pad  & \u4_pad  ;
  assign n1299 = ~n1288 & ~n1289 ;
  assign n1290 = \t0_pad  & \z4_pad  ;
  assign n1291 = \i4_pad  & \s0_pad  ;
  assign n1300 = ~n1290 & ~n1291 ;
  assign n1306 = n1299 & n1300 ;
  assign n1307 = n1305 & n1306 ;
  assign n1308 = n1304 & n1307 ;
  assign n1311 = \q1_pad  & n1243 ;
  assign n1312 = n1245 & n1311 ;
  assign n1309 = \r1_pad  & ~n1245 ;
  assign n1310 = \p1_pad  & ~n1243 ;
  assign n1313 = ~n1309 & ~n1310 ;
  assign n1314 = ~n1312 & n1313 ;
  assign n1315 = n1253 & ~n1314 ;
  assign n1317 = ~\q2_pad  & n303 ;
  assign n1316 = \q2_pad  & ~n303 ;
  assign n1318 = n277 & ~n1316 ;
  assign n1319 = ~n1317 & n1318 ;
  assign n1320 = n313 & n330 ;
  assign n1321 = n361 & ~n1320 ;
  assign n1323 = \q3_pad  & n1321 ;
  assign n1322 = ~\q3_pad  & ~n1321 ;
  assign n1324 = n316 & ~n1322 ;
  assign n1325 = ~n1323 & n1324 ;
  assign n1326 = ~n317 & ~n1325 ;
  assign n1329 = ~\q4_pad  & ~n1200 ;
  assign n1328 = ~n1112 & n1274 ;
  assign n1330 = n887 & ~n1328 ;
  assign n1331 = ~n1329 & n1330 ;
  assign n1327 = \c4_pad  & ~n887 ;
  assign n1332 = ~z_pad & ~n1327 ;
  assign n1333 = ~n1331 & n1332 ;
  assign n1336 = \r5_pad  & n1205 ;
  assign n1337 = n1207 & n1336 ;
  assign n1334 = \p5_pad  & ~n1207 ;
  assign n1335 = \q5_pad  & ~n1205 ;
  assign n1338 = ~n1334 & ~n1335 ;
  assign n1339 = ~n1337 & n1338 ;
  assign n1340 = n1215 & ~n1339 ;
  assign n1351 = \o4_pad  & \q0_pad  ;
  assign n1349 = \p0_pad  & \v3_pad  ;
  assign n1350 = \h3_pad  & \m0_pad  ;
  assign n1356 = ~n1349 & ~n1350 ;
  assign n1357 = ~n1351 & n1356 ;
  assign n1345 = \o0_pad  & \y3_pad  ;
  assign n1346 = \k4_pad  & \r0_pad  ;
  assign n1354 = ~n1345 & ~n1346 ;
  assign n1347 = \k0_pad  & \s3_pad  ;
  assign n1348 = \l0_pad  & \o3_pad  ;
  assign n1355 = ~n1347 & ~n1348 ;
  assign n1358 = n1354 & n1355 ;
  assign n1341 = \b4_pad  & \n0_pad  ;
  assign n1342 = \t4_pad  & \u0_pad  ;
  assign n1352 = ~n1341 & ~n1342 ;
  assign n1343 = \t0_pad  & \y4_pad  ;
  assign n1344 = \f4_pad  & \s0_pad  ;
  assign n1353 = ~n1343 & ~n1344 ;
  assign n1359 = n1352 & n1353 ;
  assign n1360 = n1358 & n1359 ;
  assign n1361 = n1357 & n1360 ;
  assign n1364 = \r1_pad  & n1243 ;
  assign n1365 = n1245 & n1364 ;
  assign n1362 = \p1_pad  & ~n1245 ;
  assign n1363 = \q1_pad  & ~n1243 ;
  assign n1366 = ~n1362 & ~n1363 ;
  assign n1367 = ~n1365 & n1366 ;
  assign n1368 = n1253 & ~n1367 ;
  assign n1370 = \q2_pad  & n273 ;
  assign n1369 = ~\q2_pad  & ~n273 ;
  assign n1371 = ~n303 & ~n1369 ;
  assign n1372 = ~n1370 & n1371 ;
  assign n1374 = ~\r2_pad  & ~n1372 ;
  assign n1373 = \r2_pad  & n1372 ;
  assign n1375 = n277 & ~n1373 ;
  assign n1376 = ~n1374 & n1375 ;
  assign n1378 = n313 & ~n331 ;
  assign n1377 = ~\q3_pad  & ~n313 ;
  assign n1379 = n361 & ~n1377 ;
  assign n1380 = ~n1378 & n1379 ;
  assign n1382 = ~\r3_pad  & ~n1380 ;
  assign n1381 = \r3_pad  & n1380 ;
  assign n1383 = n316 & ~n1381 ;
  assign n1384 = ~n1382 & n1383 ;
  assign n1385 = ~\r4_pad  & n199 ;
  assign n1386 = n197 & ~n200 ;
  assign n1387 = ~n1385 & n1386 ;
  assign n1398 = \n4_pad  & \q0_pad  ;
  assign n1396 = \p0_pad  & \u3_pad  ;
  assign n1397 = \g3_pad  & \m0_pad  ;
  assign n1403 = ~n1396 & ~n1397 ;
  assign n1404 = ~n1398 & n1403 ;
  assign n1392 = \o0_pad  & \x3_pad  ;
  assign n1393 = \j4_pad  & \r0_pad  ;
  assign n1401 = ~n1392 & ~n1393 ;
  assign n1394 = \k0_pad  & \r3_pad  ;
  assign n1395 = \l0_pad  & \n3_pad  ;
  assign n1402 = ~n1394 & ~n1395 ;
  assign n1405 = n1401 & n1402 ;
  assign n1388 = \a4_pad  & \n0_pad  ;
  assign n1389 = \s4_pad  & \u0_pad  ;
  assign n1399 = ~n1388 & ~n1389 ;
  assign n1390 = \t0_pad  & \x4_pad  ;
  assign n1391 = \e4_pad  & \s0_pad  ;
  assign n1400 = ~n1390 & ~n1391 ;
  assign n1406 = n1399 & n1400 ;
  assign n1407 = n1405 & n1406 ;
  assign n1408 = n1404 & n1407 ;
  assign n1410 = \s1_pad  & ~n263 ;
  assign n1411 = ~\s1_pad  & n263 ;
  assign n1412 = ~n1410 & ~n1411 ;
  assign n1413 = n242 & ~n1412 ;
  assign n1409 = ~\w2_pad  & ~n242 ;
  assign n1414 = ~b_pad & ~n1409 ;
  assign n1415 = ~n1413 & n1414 ;
  assign n1417 = ~n273 & n283 ;
  assign n1416 = n273 & n290 ;
  assign n1418 = ~n303 & ~n1416 ;
  assign n1419 = ~n1417 & n1418 ;
  assign n1421 = ~\s2_pad  & ~n1419 ;
  assign n1420 = \s2_pad  & n1419 ;
  assign n1422 = n277 & ~n1420 ;
  assign n1423 = ~n1421 & n1422 ;
  assign n1425 = ~\s3_pad  & ~n363 ;
  assign n1424 = \s3_pad  & n363 ;
  assign n1426 = n316 & ~n1424 ;
  assign n1427 = ~n1425 & n1426 ;
  assign n1428 = ~n317 & ~n1427 ;
  assign n1429 = ~\s4_pad  & ~n200 ;
  assign n1430 = n198 & ~n201 ;
  assign n1431 = ~n1429 & n1430 ;
  assign \a10_pad  = n205 ;
  assign \a6_pad  = ~n226 ;
  assign \a7_pad  = n271 ;
  assign \a8_pad  = ~n310 ;
  assign \a9_pad  = ~n372 ;
  assign \b10_pad  = n376 ;
  assign \b6_pad  = ~n415 ;
  assign \b7_pad  = n426 ;
  assign \b8_pad  = n431 ;
  assign \b9_pad  = n450 ;
  assign \c10_pad  = n454 ;
  assign \c53  = ~n463 ;
  assign \c6_pad  = n473 ;
  assign \c7_pad  = ~n489 ;
  assign \c8_pad  = n493 ;
  assign \c9_pad  = n505 ;
  assign \d10_pad  = n509 ;
  assign \d6_pad  = n515 ;
  assign \d7_pad  = ~n528 ;
  assign \d8_pad  = n540 ;
  assign \d9_pad  = n551 ;
  assign \e10_pad  = n556 ;
  assign \e6_pad  = n560 ;
  assign \e7_pad  = ~n573 ;
  assign \e8_pad  = n581 ;
  assign \e9_pad  = ~n597 ;
  assign \f10_pad  = n601 ;
  assign \f22  = ~n608 ;
  assign \f6_pad  = n612 ;
  assign \f7_pad  = n627 ;
  assign \f8_pad  = n635 ;
  assign \f9_pad  = ~n649 ;
  assign \g10_pad  = n653 ;
  assign \g6_pad  = n658 ;
  assign \g7_pad  = ~n671 ;
  assign \g8_pad  = ~n680 ;
  assign \g9_pad  = ~n693 ;
  assign \h6_pad  = n697 ;
  assign \h7_pad  = ~n708 ;
  assign \h8_pad  = ~n719 ;
  assign \h9_pad  = n733 ;
  assign \i6_pad  = n737 ;
  assign \i7_pad  = ~n738 ;
  assign \i8_pad  = ~n751 ;
  assign \i9_pad  = ~n762 ;
  assign \j10_pad  = ~n188 ;
  assign \j6_pad  = n766 ;
  assign \j7_pad  = ~n770 ;
  assign \j8_pad  = n779 ;
  assign \j9_pad  = ~n790 ;
  assign \k10_pad  = ~n793 ;
  assign \k53  = ~n797 ;
  assign \k6_pad  = n801 ;
  assign \k7_pad  = ~n805 ;
  assign \k8_pad  = ~n814 ;
  assign \k9_pad  = ~n815 ;
  assign \l10_pad  = ~n818 ;
  assign \l7_pad  = ~n832 ;
  assign \l8_pad  = ~n843 ;
  assign \l9_pad  = ~n846 ;
  assign \m10_pad  = ~n858 ;
  assign \m7_pad  = ~n865 ;
  assign \m8_pad  = n869 ;
  assign \m9_pad  = ~n872 ;
  assign \n10_pad  = n875 ;
  assign \n6_pad  = ~n250 ;
  assign \n7_pad  = ~n878 ;
  assign \n8_pad  = n886 ;
  assign \n9_pad  = ~n893 ;
  assign \o10_pad  = n851 ;
  assign \o6_pad  = ~n896 ;
  assign \o7_pad  = ~n904 ;
  assign \o8_pad  = n912 ;
  assign \o9_pad  = ~n919 ;
  assign \p6_pad  = ~n922 ;
  assign \p7_pad  = ~n929 ;
  assign \p8_pad  = ~n938 ;
  assign \p9_pad  = ~n941 ;
  assign \q10_pad  = n946 ;
  assign \q6_pad  = ~n951 ;
  assign \q7_pad  = ~n960 ;
  assign \q8_pad  = n965 ;
  assign \q9_pad  = ~n973 ;
  assign \r10_pad  = n977 ;
  assign \r7_pad  = ~n985 ;
  assign \r8_pad  = n989 ;
  assign \r9_pad  = ~n996 ;
  assign \s5_pad  = ~n1017 ;
  assign \s7_pad  = ~n1024 ;
  assign \s8_pad  = n1032 ;
  assign \s9_pad  = ~n1041 ;
  assign \t10_pad  = n1053 ;
  assign \t5_pad  = ~n1074 ;
  assign \t6_pad  = n1095 ;
  assign \t7_pad  = ~n1102 ;
  assign \t8_pad  = n1110 ;
  assign \t9_pad  = ~n1118 ;
  assign \u5_pad  = ~n1139 ;
  assign \u7_pad  = n1145 ;
  assign \u8_pad  = n1153 ;
  assign \u9_pad  = ~n1160 ;
  assign \v10_pad  = ~n311 ;
  assign \v5_pad  = ~n1181 ;
  assign \v6_pad  = ~n239 ;
  assign \v7_pad  = ~n1188 ;
  assign \v8_pad  = ~n1197 ;
  assign \v9_pad  = ~n1204 ;
  assign \w10_pad  = ~n1220 ;
  assign \w5_pad  = ~n1241 ;
  assign \w6_pad  = ~n1258 ;
  assign \w7_pad  = ~n1261 ;
  assign \w8_pad  = ~n1270 ;
  assign \w9_pad  = n1276 ;
  assign \x10_pad  = n1283 ;
  assign \x21  = ~n1287 ;
  assign \x5_pad  = ~n1308 ;
  assign \x6_pad  = n1315 ;
  assign \x7_pad  = n1319 ;
  assign \x8_pad  = ~n1326 ;
  assign \x9_pad  = ~n1333 ;
  assign \y10_pad  = n1340 ;
  assign \y5_pad  = ~n1361 ;
  assign \y6_pad  = n1368 ;
  assign \y7_pad  = n1376 ;
  assign \y8_pad  = n1384 ;
  assign \y9_pad  = n1387 ;
  assign \z5_pad  = ~n1408 ;
  assign \z6_pad  = n1415 ;
  assign \z7_pad  = n1423 ;
  assign \z8_pad  = ~n1428 ;
  assign \z9_pad  = n1431 ;
endmodule
