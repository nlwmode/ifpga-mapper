module top (\101(0)_pad , \104(1)_pad , \107(2)_pad , \110(3)_pad , \113(4)_pad , \116(5)_pad , \119(6)_pad , \122(7)_pad , \125(8)_pad , \128(9)_pad , \131(10)_pad , \134(11)_pad , \137(12)_pad , \140(13)_pad , \143(14)_pad , \146(15)_pad , \210(16)_pad , \214(17)_pad , \217(18)_pad , \221(19)_pad , \224(20)_pad , \227(21)_pad , \234(22)_pad , \237(23)_pad , \469(24)_pad , \472(25)_pad , \475(26)_pad , \478(27)_pad , \898(28)_pad , \900(29)_pad , \902(30)_pad , \952(31)_pad , \953(32)_pad , \12(862)_pad , \15(861)_pad , \18(860)_pad , \21(859)_pad , \24(858)_pad , \27(857)_pad , \3(865)_pad , \30(856)_pad , \33(855)_pad , \36(854)_pad , \39(853)_pad , \42(852)_pad , \45(851)_pad , \48(850)_pad , \51(899)_pad , \54(900)_pad , \57(912)_pad , \6(864)_pad , \60(901)_pad , \63(902)_pad , \66(903)_pad , \69(908)_pad , \72(909)_pad , \75(866)_pad , \9(863)_pad );
	input \101(0)_pad  ;
	input \104(1)_pad  ;
	input \107(2)_pad  ;
	input \110(3)_pad  ;
	input \113(4)_pad  ;
	input \116(5)_pad  ;
	input \119(6)_pad  ;
	input \122(7)_pad  ;
	input \125(8)_pad  ;
	input \128(9)_pad  ;
	input \131(10)_pad  ;
	input \134(11)_pad  ;
	input \137(12)_pad  ;
	input \140(13)_pad  ;
	input \143(14)_pad  ;
	input \146(15)_pad  ;
	input \210(16)_pad  ;
	input \214(17)_pad  ;
	input \217(18)_pad  ;
	input \221(19)_pad  ;
	input \224(20)_pad  ;
	input \227(21)_pad  ;
	input \234(22)_pad  ;
	input \237(23)_pad  ;
	input \469(24)_pad  ;
	input \472(25)_pad  ;
	input \475(26)_pad  ;
	input \478(27)_pad  ;
	input \898(28)_pad  ;
	input \900(29)_pad  ;
	input \902(30)_pad  ;
	input \952(31)_pad  ;
	input \953(32)_pad  ;
	output \12(862)_pad  ;
	output \15(861)_pad  ;
	output \18(860)_pad  ;
	output \21(859)_pad  ;
	output \24(858)_pad  ;
	output \27(857)_pad  ;
	output \3(865)_pad  ;
	output \30(856)_pad  ;
	output \33(855)_pad  ;
	output \36(854)_pad  ;
	output \39(853)_pad  ;
	output \42(852)_pad  ;
	output \45(851)_pad  ;
	output \48(850)_pad  ;
	output \51(899)_pad  ;
	output \54(900)_pad  ;
	output \57(912)_pad  ;
	output \6(864)_pad  ;
	output \60(901)_pad  ;
	output \63(902)_pad  ;
	output \66(903)_pad  ;
	output \69(908)_pad  ;
	output \72(909)_pad  ;
	output \75(866)_pad  ;
	output \9(863)_pad  ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	LUT3 #(
		.INIT('h69)
	) name0 (
		\128(9)_pad ,
		\143(14)_pad ,
		\146(15)_pad ,
		_w35_
	);
	LUT3 #(
		.INIT('h96)
	) name1 (
		\131(10)_pad ,
		\134(11)_pad ,
		\137(12)_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\227(21)_pad ,
		\953(32)_pad ,
		_w37_
	);
	LUT3 #(
		.INIT('h96)
	) name3 (
		_w35_,
		_w36_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h6)
	) name4 (
		\104(1)_pad ,
		\107(2)_pad ,
		_w39_
	);
	LUT3 #(
		.INIT('h69)
	) name5 (
		\101(0)_pad ,
		\110(3)_pad ,
		\140(13)_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h9)
	) name6 (
		_w39_,
		_w40_,
		_w41_
	);
	LUT4 #(
		.INIT('h4554)
	) name7 (
		\469(24)_pad ,
		\902(30)_pad ,
		_w38_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\469(24)_pad ,
		\902(30)_pad ,
		_w43_
	);
	LUT3 #(
		.INIT('h60)
	) name9 (
		_w39_,
		_w40_,
		_w43_,
		_w44_
	);
	LUT3 #(
		.INIT('h90)
	) name10 (
		_w39_,
		_w40_,
		_w43_,
		_w45_
	);
	LUT3 #(
		.INIT('ha2)
	) name11 (
		\221(19)_pad ,
		\234(22)_pad ,
		\902(30)_pad ,
		_w46_
	);
	LUT4 #(
		.INIT('h001b)
	) name12 (
		_w38_,
		_w44_,
		_w45_,
		_w46_,
		_w47_
	);
	LUT4 #(
		.INIT('h9669)
	) name13 (
		\101(0)_pad ,
		\113(4)_pad ,
		\116(5)_pad ,
		\119(6)_pad ,
		_w48_
	);
	LUT4 #(
		.INIT('h6996)
	) name14 (
		\104(1)_pad ,
		\107(2)_pad ,
		\110(3)_pad ,
		\122(7)_pad ,
		_w49_
	);
	LUT3 #(
		.INIT('h59)
	) name15 (
		\125(8)_pad ,
		\224(20)_pad ,
		\953(32)_pad ,
		_w50_
	);
	LUT4 #(
		.INIT('h9669)
	) name16 (
		_w35_,
		_w48_,
		_w49_,
		_w50_,
		_w51_
	);
	LUT3 #(
		.INIT('ha8)
	) name17 (
		\210(16)_pad ,
		\237(23)_pad ,
		\902(30)_pad ,
		_w52_
	);
	LUT3 #(
		.INIT('ha8)
	) name18 (
		\214(17)_pad ,
		\237(23)_pad ,
		\902(30)_pad ,
		_w53_
	);
	LUT4 #(
		.INIT('hff4b)
	) name19 (
		\902(30)_pad ,
		_w51_,
		_w52_,
		_w53_,
		_w54_
	);
	LUT3 #(
		.INIT('h04)
	) name20 (
		_w42_,
		_w47_,
		_w54_,
		_w55_
	);
	LUT3 #(
		.INIT('h02)
	) name21 (
		\210(16)_pad ,
		\237(23)_pad ,
		\953(32)_pad ,
		_w56_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name22 (
		\210(16)_pad ,
		\237(23)_pad ,
		\902(30)_pad ,
		\953(32)_pad ,
		_w57_
	);
	LUT4 #(
		.INIT('h69ff)
	) name23 (
		_w35_,
		_w36_,
		_w48_,
		_w57_,
		_w58_
	);
	LUT4 #(
		.INIT('h0002)
	) name24 (
		\210(16)_pad ,
		\237(23)_pad ,
		\902(30)_pad ,
		\953(32)_pad ,
		_w59_
	);
	LUT4 #(
		.INIT('h96ff)
	) name25 (
		_w35_,
		_w36_,
		_w48_,
		_w59_,
		_w60_
	);
	LUT3 #(
		.INIT('h6a)
	) name26 (
		\472(25)_pad ,
		_w58_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h6)
	) name27 (
		\125(8)_pad ,
		\140(13)_pad ,
		_w62_
	);
	LUT3 #(
		.INIT('h96)
	) name28 (
		\125(8)_pad ,
		\140(13)_pad ,
		\146(15)_pad ,
		_w63_
	);
	LUT2 #(
		.INIT('h6)
	) name29 (
		\119(6)_pad ,
		\128(9)_pad ,
		_w64_
	);
	LUT2 #(
		.INIT('h9)
	) name30 (
		\110(3)_pad ,
		\137(12)_pad ,
		_w65_
	);
	LUT3 #(
		.INIT('h08)
	) name31 (
		\221(19)_pad ,
		\234(22)_pad ,
		\953(32)_pad ,
		_w66_
	);
	LUT4 #(
		.INIT('h6996)
	) name32 (
		_w63_,
		_w64_,
		_w65_,
		_w66_,
		_w67_
	);
	LUT3 #(
		.INIT('ha2)
	) name33 (
		\217(18)_pad ,
		\234(22)_pad ,
		\902(30)_pad ,
		_w68_
	);
	LUT3 #(
		.INIT('h1e)
	) name34 (
		\902(30)_pad ,
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w61_,
		_w69_,
		_w70_
	);
	LUT4 #(
		.INIT('h9669)
	) name36 (
		\122(7)_pad ,
		\125(8)_pad ,
		\140(13)_pad ,
		\146(15)_pad ,
		_w71_
	);
	LUT3 #(
		.INIT('h02)
	) name37 (
		\214(17)_pad ,
		\237(23)_pad ,
		\953(32)_pad ,
		_w72_
	);
	LUT2 #(
		.INIT('h6)
	) name38 (
		\104(1)_pad ,
		\113(4)_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h9)
	) name39 (
		\131(10)_pad ,
		\143(14)_pad ,
		_w74_
	);
	LUT3 #(
		.INIT('h06)
	) name40 (
		\131(10)_pad ,
		\143(14)_pad ,
		\902(30)_pad ,
		_w75_
	);
	LUT4 #(
		.INIT('h1400)
	) name41 (
		_w71_,
		_w72_,
		_w73_,
		_w75_,
		_w76_
	);
	LUT3 #(
		.INIT('h09)
	) name42 (
		\131(10)_pad ,
		\143(14)_pad ,
		\902(30)_pad ,
		_w77_
	);
	LUT4 #(
		.INIT('h4100)
	) name43 (
		_w71_,
		_w72_,
		_w73_,
		_w77_,
		_w78_
	);
	LUT4 #(
		.INIT('h2800)
	) name44 (
		_w71_,
		_w72_,
		_w73_,
		_w77_,
		_w79_
	);
	LUT4 #(
		.INIT('h8200)
	) name45 (
		_w71_,
		_w72_,
		_w73_,
		_w75_,
		_w80_
	);
	LUT4 #(
		.INIT('h0001)
	) name46 (
		_w76_,
		_w78_,
		_w79_,
		_w80_,
		_w81_
	);
	LUT3 #(
		.INIT('h08)
	) name47 (
		\217(18)_pad ,
		\234(22)_pad ,
		\953(32)_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h6)
	) name48 (
		\134(11)_pad ,
		\143(14)_pad ,
		_w83_
	);
	LUT4 #(
		.INIT('h6996)
	) name49 (
		\107(2)_pad ,
		\116(5)_pad ,
		\122(7)_pad ,
		\128(9)_pad ,
		_w84_
	);
	LUT3 #(
		.INIT('h69)
	) name50 (
		_w82_,
		_w83_,
		_w84_,
		_w85_
	);
	LUT3 #(
		.INIT('ha9)
	) name51 (
		\478(27)_pad ,
		\902(30)_pad ,
		_w85_,
		_w86_
	);
	LUT4 #(
		.INIT('h7000)
	) name52 (
		\234(22)_pad ,
		\237(23)_pad ,
		\902(30)_pad ,
		\953(32)_pad ,
		_w87_
	);
	LUT4 #(
		.INIT('h0070)
	) name53 (
		\234(22)_pad ,
		\237(23)_pad ,
		\952(31)_pad ,
		\953(32)_pad ,
		_w88_
	);
	LUT3 #(
		.INIT('h0b)
	) name54 (
		\898(28)_pad ,
		_w87_,
		_w88_,
		_w89_
	);
	LUT4 #(
		.INIT('h0056)
	) name55 (
		\478(27)_pad ,
		\902(30)_pad ,
		_w85_,
		_w89_,
		_w90_
	);
	LUT3 #(
		.INIT('h60)
	) name56 (
		\475(26)_pad ,
		_w81_,
		_w90_,
		_w91_
	);
	LUT3 #(
		.INIT('h80)
	) name57 (
		_w55_,
		_w70_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name58 (
		\110(3)_pad ,
		_w55_,
		_w70_,
		_w91_,
		_w93_
	);
	LUT4 #(
		.INIT('h0010)
	) name59 (
		\110(3)_pad ,
		_w42_,
		_w47_,
		_w54_,
		_w94_
	);
	LUT3 #(
		.INIT('h80)
	) name60 (
		_w70_,
		_w91_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('he)
	) name61 (
		_w93_,
		_w95_,
		_w96_
	);
	LUT4 #(
		.INIT('h050d)
	) name62 (
		\221(19)_pad ,
		\234(22)_pad ,
		\469(24)_pad ,
		\902(30)_pad ,
		_w97_
	);
	LUT4 #(
		.INIT('hbe00)
	) name63 (
		\902(30)_pad ,
		_w38_,
		_w41_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h50d0)
	) name64 (
		\221(19)_pad ,
		\234(22)_pad ,
		\469(24)_pad ,
		\902(30)_pad ,
		_w99_
	);
	LUT4 #(
		.INIT('h4100)
	) name65 (
		\902(30)_pad ,
		_w38_,
		_w41_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w98_,
		_w100_,
		_w101_
	);
	LUT3 #(
		.INIT('h54)
	) name67 (
		_w54_,
		_w98_,
		_w100_,
		_w102_
	);
	LUT3 #(
		.INIT('h90)
	) name68 (
		\475(26)_pad ,
		_w81_,
		_w90_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w61_,
		_w69_,
		_w104_
	);
	LUT3 #(
		.INIT('h80)
	) name70 (
		_w102_,
		_w103_,
		_w104_,
		_w105_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name71 (
		\113(4)_pad ,
		_w102_,
		_w103_,
		_w104_,
		_w106_
	);
	LUT4 #(
		.INIT('h00a9)
	) name72 (
		\478(27)_pad ,
		\902(30)_pad ,
		_w85_,
		_w89_,
		_w107_
	);
	LUT3 #(
		.INIT('h60)
	) name73 (
		\475(26)_pad ,
		_w81_,
		_w107_,
		_w108_
	);
	LUT3 #(
		.INIT('h80)
	) name74 (
		_w102_,
		_w104_,
		_w108_,
		_w109_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name75 (
		\116(5)_pad ,
		_w102_,
		_w104_,
		_w108_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w61_,
		_w69_,
		_w111_
	);
	LUT3 #(
		.INIT('h80)
	) name77 (
		_w91_,
		_w102_,
		_w111_,
		_w112_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name78 (
		\119(6)_pad ,
		_w91_,
		_w102_,
		_w111_,
		_w113_
	);
	LUT4 #(
		.INIT('h1110)
	) name79 (
		\119(6)_pad ,
		_w54_,
		_w98_,
		_w100_,
		_w114_
	);
	LUT3 #(
		.INIT('h80)
	) name80 (
		_w91_,
		_w111_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('he)
	) name81 (
		_w113_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w61_,
		_w69_,
		_w117_
	);
	LUT3 #(
		.INIT('h90)
	) name83 (
		\475(26)_pad ,
		_w81_,
		_w107_,
		_w118_
	);
	LUT3 #(
		.INIT('h80)
	) name84 (
		_w102_,
		_w117_,
		_w118_,
		_w119_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name85 (
		\122(7)_pad ,
		_w102_,
		_w117_,
		_w118_,
		_w120_
	);
	LUT4 #(
		.INIT('h1110)
	) name86 (
		\122(7)_pad ,
		_w54_,
		_w98_,
		_w100_,
		_w121_
	);
	LUT3 #(
		.INIT('h80)
	) name87 (
		_w117_,
		_w118_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('he)
	) name88 (
		_w120_,
		_w122_,
		_w123_
	);
	LUT3 #(
		.INIT('h0b)
	) name89 (
		\900(29)_pad ,
		_w87_,
		_w88_,
		_w124_
	);
	LUT4 #(
		.INIT('h0056)
	) name90 (
		\478(27)_pad ,
		\902(30)_pad ,
		_w85_,
		_w124_,
		_w125_
	);
	LUT3 #(
		.INIT('h90)
	) name91 (
		\475(26)_pad ,
		_w81_,
		_w125_,
		_w126_
	);
	LUT3 #(
		.INIT('h80)
	) name92 (
		_w70_,
		_w102_,
		_w126_,
		_w127_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name93 (
		\125(8)_pad ,
		_w70_,
		_w102_,
		_w126_,
		_w128_
	);
	LUT4 #(
		.INIT('h1110)
	) name94 (
		\125(8)_pad ,
		_w54_,
		_w98_,
		_w100_,
		_w129_
	);
	LUT3 #(
		.INIT('h80)
	) name95 (
		_w70_,
		_w126_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('he)
	) name96 (
		_w128_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h80)
	) name97 (
		_w55_,
		_w91_,
		_w104_,
		_w132_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name98 (
		\101(0)_pad ,
		_w55_,
		_w91_,
		_w104_,
		_w133_
	);
	LUT4 #(
		.INIT('h00a9)
	) name99 (
		\478(27)_pad ,
		\902(30)_pad ,
		_w85_,
		_w124_,
		_w134_
	);
	LUT3 #(
		.INIT('h60)
	) name100 (
		\475(26)_pad ,
		_w81_,
		_w134_,
		_w135_
	);
	LUT3 #(
		.INIT('h80)
	) name101 (
		_w55_,
		_w111_,
		_w135_,
		_w136_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name102 (
		\128(9)_pad ,
		_w55_,
		_w111_,
		_w135_,
		_w137_
	);
	LUT4 #(
		.INIT('h004b)
	) name103 (
		\902(30)_pad ,
		_w51_,
		_w52_,
		_w53_,
		_w138_
	);
	LUT3 #(
		.INIT('h40)
	) name104 (
		_w42_,
		_w47_,
		_w138_,
		_w139_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name105 (
		\131(10)_pad ,
		_w104_,
		_w126_,
		_w139_,
		_w140_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name106 (
		\134(11)_pad ,
		_w104_,
		_w135_,
		_w139_,
		_w141_
	);
	LUT3 #(
		.INIT('h60)
	) name107 (
		\475(26)_pad ,
		_w81_,
		_w125_,
		_w142_
	);
	LUT3 #(
		.INIT('h80)
	) name108 (
		_w111_,
		_w139_,
		_w142_,
		_w143_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name109 (
		\137(12)_pad ,
		_w111_,
		_w139_,
		_w142_,
		_w144_
	);
	LUT4 #(
		.INIT('h1000)
	) name110 (
		\137(12)_pad ,
		_w42_,
		_w47_,
		_w138_,
		_w145_
	);
	LUT3 #(
		.INIT('h80)
	) name111 (
		_w111_,
		_w142_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('he)
	) name112 (
		_w144_,
		_w146_,
		_w147_
	);
	LUT3 #(
		.INIT('h80)
	) name113 (
		_w70_,
		_w126_,
		_w139_,
		_w148_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name114 (
		\140(13)_pad ,
		_w70_,
		_w126_,
		_w139_,
		_w149_
	);
	LUT3 #(
		.INIT('h90)
	) name115 (
		\475(26)_pad ,
		_w81_,
		_w134_,
		_w150_
	);
	LUT3 #(
		.INIT('h80)
	) name116 (
		_w55_,
		_w104_,
		_w150_,
		_w151_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name117 (
		\143(14)_pad ,
		_w55_,
		_w104_,
		_w150_,
		_w152_
	);
	LUT3 #(
		.INIT('h80)
	) name118 (
		_w55_,
		_w111_,
		_w126_,
		_w153_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name119 (
		\146(15)_pad ,
		_w55_,
		_w111_,
		_w126_,
		_w154_
	);
	LUT4 #(
		.INIT('h0001)
	) name120 (
		_w143_,
		_w148_,
		_w151_,
		_w153_,
		_w155_
	);
	LUT4 #(
		.INIT('h57ff)
	) name121 (
		_w104_,
		_w126_,
		_w135_,
		_w139_,
		_w156_
	);
	LUT3 #(
		.INIT('h10)
	) name122 (
		_w127_,
		_w136_,
		_w156_,
		_w157_
	);
	LUT4 #(
		.INIT('h57ff)
	) name123 (
		_w55_,
		_w103_,
		_w108_,
		_w117_,
		_w158_
	);
	LUT3 #(
		.INIT('h10)
	) name124 (
		_w119_,
		_w132_,
		_w158_,
		_w159_
	);
	LUT4 #(
		.INIT('h0001)
	) name125 (
		_w92_,
		_w105_,
		_w109_,
		_w112_,
		_w160_
	);
	LUT4 #(
		.INIT('h8000)
	) name126 (
		_w155_,
		_w157_,
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\210(16)_pad ,
		\902(30)_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		\952(31)_pad ,
		\953(32)_pad ,
		_w163_
	);
	LUT4 #(
		.INIT('h009a)
	) name129 (
		_w51_,
		_w161_,
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h6)
	) name130 (
		_w38_,
		_w41_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\469(24)_pad ,
		\902(30)_pad ,
		_w166_
	);
	LUT4 #(
		.INIT('h1203)
	) name132 (
		_w161_,
		_w163_,
		_w165_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('h9669)
	) name133 (
		_w35_,
		_w36_,
		_w48_,
		_w56_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\472(25)_pad ,
		\902(30)_pad ,
		_w169_
	);
	LUT4 #(
		.INIT('h1203)
	) name135 (
		_w161_,
		_w163_,
		_w168_,
		_w169_,
		_w170_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name136 (
		\104(1)_pad ,
		_w55_,
		_w103_,
		_w117_,
		_w171_
	);
	LUT4 #(
		.INIT('h9669)
	) name137 (
		_w71_,
		_w72_,
		_w73_,
		_w74_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\475(26)_pad ,
		\902(30)_pad ,
		_w173_
	);
	LUT4 #(
		.INIT('h1203)
	) name139 (
		_w161_,
		_w163_,
		_w172_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\478(27)_pad ,
		\902(30)_pad ,
		_w175_
	);
	LUT4 #(
		.INIT('h0605)
	) name141 (
		_w85_,
		_w161_,
		_w163_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\217(18)_pad ,
		\902(30)_pad ,
		_w177_
	);
	LUT4 #(
		.INIT('h0605)
	) name143 (
		_w67_,
		_w161_,
		_w163_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		\224(20)_pad ,
		\953(32)_pad ,
		_w179_
	);
	LUT3 #(
		.INIT('h06)
	) name145 (
		_w48_,
		_w49_,
		_w179_,
		_w180_
	);
	LUT4 #(
		.INIT('hea00)
	) name146 (
		\953(32)_pad ,
		_w159_,
		_w160_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		\898(28)_pad ,
		\953(32)_pad ,
		_w182_
	);
	LUT3 #(
		.INIT('h90)
	) name148 (
		_w48_,
		_w49_,
		_w179_,
		_w183_
	);
	LUT3 #(
		.INIT('h41)
	) name149 (
		\953(32)_pad ,
		_w48_,
		_w49_,
		_w184_
	);
	LUT4 #(
		.INIT('h080f)
	) name150 (
		_w159_,
		_w160_,
		_w183_,
		_w184_,
		_w185_
	);
	LUT3 #(
		.INIT('hef)
	) name151 (
		_w181_,
		_w182_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		\227(21)_pad ,
		\953(32)_pad ,
		_w187_
	);
	LUT4 #(
		.INIT('h0096)
	) name153 (
		_w35_,
		_w36_,
		_w62_,
		_w187_,
		_w188_
	);
	LUT4 #(
		.INIT('hea00)
	) name154 (
		\953(32)_pad ,
		_w155_,
		_w157_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		\900(29)_pad ,
		\953(32)_pad ,
		_w190_
	);
	LUT4 #(
		.INIT('h0096)
	) name156 (
		_w35_,
		_w36_,
		_w62_,
		_w190_,
		_w191_
	);
	LUT3 #(
		.INIT('h8f)
	) name157 (
		\227(21)_pad ,
		\900(29)_pad ,
		\953(32)_pad ,
		_w192_
	);
	LUT4 #(
		.INIT('hea00)
	) name158 (
		\953(32)_pad ,
		_w155_,
		_w157_,
		_w192_,
		_w193_
	);
	LUT3 #(
		.INIT('hab)
	) name159 (
		_w189_,
		_w191_,
		_w193_,
		_w194_
	);
	LUT3 #(
		.INIT('h06)
	) name160 (
		\475(26)_pad ,
		_w81_,
		_w86_,
		_w195_
	);
	LUT4 #(
		.INIT('h0600)
	) name161 (
		\475(26)_pad ,
		_w81_,
		_w86_,
		_w138_,
		_w196_
	);
	LUT4 #(
		.INIT('h4555)
	) name162 (
		\953(32)_pad ,
		_w101_,
		_w117_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		\952(31)_pad ,
		_w197_,
		_w198_
	);
	LUT3 #(
		.INIT('h10)
	) name164 (
		_w98_,
		_w100_,
		_w138_,
		_w199_
	);
	LUT4 #(
		.INIT('h1b00)
	) name165 (
		_w38_,
		_w44_,
		_w45_,
		_w46_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		_w42_,
		_w200_,
		_w201_
	);
	LUT4 #(
		.INIT('h7737)
	) name167 (
		_w102_,
		_w195_,
		_w199_,
		_w201_,
		_w202_
	);
	LUT4 #(
		.INIT('h2112)
	) name168 (
		\475(26)_pad ,
		_w53_,
		_w81_,
		_w86_,
		_w203_
	);
	LUT3 #(
		.INIT('h4b)
	) name169 (
		\902(30)_pad ,
		_w51_,
		_w52_,
		_w204_
	);
	LUT4 #(
		.INIT('ha090)
	) name170 (
		\478(27)_pad ,
		\902(30)_pad ,
		_w53_,
		_w85_,
		_w205_
	);
	LUT4 #(
		.INIT('h007b)
	) name171 (
		\475(26)_pad ,
		_w53_,
		_w81_,
		_w205_,
		_w206_
	);
	LUT4 #(
		.INIT('h1000)
	) name172 (
		_w101_,
		_w203_,
		_w204_,
		_w206_,
		_w207_
	);
	LUT3 #(
		.INIT('he0)
	) name173 (
		_w61_,
		_w69_,
		_w88_,
		_w208_
	);
	LUT4 #(
		.INIT('hdc00)
	) name174 (
		_w101_,
		_w117_,
		_w196_,
		_w208_,
		_w209_
	);
	LUT4 #(
		.INIT('hf700)
	) name175 (
		_w117_,
		_w202_,
		_w207_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		_w197_,
		_w210_,
		_w211_
	);
	LUT3 #(
		.INIT('h13)
	) name177 (
		_w161_,
		_w198_,
		_w211_,
		_w212_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name178 (
		\107(2)_pad ,
		_w55_,
		_w108_,
		_w117_,
		_w213_
	);
	assign \12(862)_pad  = _w96_ ;
	assign \15(861)_pad  = _w106_ ;
	assign \18(860)_pad  = _w110_ ;
	assign \21(859)_pad  = _w116_ ;
	assign \24(858)_pad  = _w123_ ;
	assign \27(857)_pad  = _w131_ ;
	assign \3(865)_pad  = _w133_ ;
	assign \30(856)_pad  = _w137_ ;
	assign \33(855)_pad  = _w140_ ;
	assign \36(854)_pad  = _w141_ ;
	assign \39(853)_pad  = _w147_ ;
	assign \42(852)_pad  = _w149_ ;
	assign \45(851)_pad  = _w152_ ;
	assign \48(850)_pad  = _w154_ ;
	assign \51(899)_pad  = _w164_ ;
	assign \54(900)_pad  = _w167_ ;
	assign \57(912)_pad  = _w170_ ;
	assign \6(864)_pad  = _w171_ ;
	assign \60(901)_pad  = _w174_ ;
	assign \63(902)_pad  = _w176_ ;
	assign \66(903)_pad  = _w178_ ;
	assign \69(908)_pad  = _w186_ ;
	assign \72(909)_pad  = _w194_ ;
	assign \75(866)_pad  = _w212_ ;
	assign \9(863)_pad  = _w213_ ;
endmodule;