module top( \B_reg/NET0131  , \IR_reg[0]/NET0131  , \IR_reg[10]/NET0131  , \IR_reg[11]/NET0131  , \IR_reg[12]/NET0131  , \IR_reg[13]/NET0131  , \IR_reg[14]/NET0131  , \IR_reg[15]/NET0131  , \IR_reg[16]/NET0131  , \IR_reg[17]/NET0131  , \IR_reg[18]/NET0131  , \IR_reg[19]/NET0131  , \IR_reg[1]/NET0131  , \IR_reg[20]/NET0131  , \IR_reg[21]/NET0131  , \IR_reg[22]/NET0131  , \IR_reg[23]/NET0131  , \IR_reg[24]/NET0131  , \IR_reg[25]/NET0131  , \IR_reg[26]/NET0131  , \IR_reg[27]/NET0131  , \IR_reg[28]/NET0131  , \IR_reg[29]/NET0131  , \IR_reg[2]/NET0131  , \IR_reg[30]/NET0131  , \IR_reg[31]/NET0131  , \IR_reg[3]/NET0131  , \IR_reg[4]/NET0131  , \IR_reg[5]/NET0131  , \IR_reg[6]/NET0131  , \IR_reg[7]/NET0131  , \IR_reg[8]/NET0131  , \IR_reg[9]/NET0131  , \addr[0]_pad  , \addr[10]_pad  , \addr[11]_pad  , \addr[12]_pad  , \addr[13]_pad  , \addr[14]_pad  , \addr[15]_pad  , \addr[16]_pad  , \addr[17]_pad  , \addr[18]_pad  , \addr[19]_pad  , \addr[1]_pad  , \addr[2]_pad  , \addr[3]_pad  , \addr[4]_pad  , \addr[5]_pad  , \addr[6]_pad  , \addr[7]_pad  , \addr[8]_pad  , \addr[9]_pad  , \d_reg[0]/NET0131  , \d_reg[1]/NET0131  , \datai[0]_pad  , \datai[10]_pad  , \datai[11]_pad  , \datai[12]_pad  , \datai[13]_pad  , \datai[14]_pad  , \datai[15]_pad  , \datai[16]_pad  , \datai[17]_pad  , \datai[18]_pad  , \datai[19]_pad  , \datai[1]_pad  , \datai[20]_pad  , \datai[21]_pad  , \datai[22]_pad  , \datai[23]_pad  , \datai[24]_pad  , \datai[25]_pad  , \datai[26]_pad  , \datai[27]_pad  , \datai[28]_pad  , \datai[29]_pad  , \datai[2]_pad  , \datai[30]_pad  , \datai[31]_pad  , \datai[3]_pad  , \datai[4]_pad  , \datai[5]_pad  , \datai[6]_pad  , \datai[7]_pad  , \datai[8]_pad  , \datai[9]_pad  , \datao[15]_pad  , \datao[28]_pad  , \datao[8]_pad  , \reg0_reg[0]/NET0131  , \reg0_reg[10]/NET0131  , \reg0_reg[11]/NET0131  , \reg0_reg[12]/NET0131  , \reg0_reg[13]/NET0131  , \reg0_reg[14]/NET0131  , \reg0_reg[15]/NET0131  , \reg0_reg[16]/NET0131  , \reg0_reg[17]/NET0131  , \reg0_reg[18]/NET0131  , \reg0_reg[19]/NET0131  , \reg0_reg[1]/NET0131  , \reg0_reg[20]/NET0131  , \reg0_reg[21]/NET0131  , \reg0_reg[22]/NET0131  , \reg0_reg[23]/NET0131  , \reg0_reg[24]/NET0131  , \reg0_reg[25]/NET0131  , \reg0_reg[26]/NET0131  , \reg0_reg[27]/NET0131  , \reg0_reg[28]/NET0131  , \reg0_reg[29]/NET0131  , \reg0_reg[2]/NET0131  , \reg0_reg[30]/NET0131  , \reg0_reg[31]/NET0131  , \reg0_reg[3]/NET0131  , \reg0_reg[4]/NET0131  , \reg0_reg[5]/NET0131  , \reg0_reg[6]/NET0131  , \reg0_reg[7]/NET0131  , \reg0_reg[8]/NET0131  , \reg0_reg[9]/NET0131  , \reg1_reg[0]/NET0131  , \reg1_reg[10]/NET0131  , \reg1_reg[11]/NET0131  , \reg1_reg[12]/NET0131  , \reg1_reg[13]/NET0131  , \reg1_reg[14]/NET0131  , \reg1_reg[15]/NET0131  , \reg1_reg[16]/NET0131  , \reg1_reg[17]/NET0131  , \reg1_reg[18]/NET0131  , \reg1_reg[19]/NET0131  , \reg1_reg[1]/NET0131  , \reg1_reg[20]/NET0131  , \reg1_reg[21]/NET0131  , \reg1_reg[22]/NET0131  , \reg1_reg[23]/NET0131  , \reg1_reg[24]/NET0131  , \reg1_reg[25]/NET0131  , \reg1_reg[26]/NET0131  , \reg1_reg[27]/NET0131  , \reg1_reg[28]/NET0131  , \reg1_reg[29]/NET0131  , \reg1_reg[2]/NET0131  , \reg1_reg[30]/NET0131  , \reg1_reg[31]/NET0131  , \reg1_reg[3]/NET0131  , \reg1_reg[4]/NET0131  , \reg1_reg[5]/NET0131  , \reg1_reg[6]/NET0131  , \reg1_reg[7]/NET0131  , \reg1_reg[8]/NET0131  , \reg1_reg[9]/NET0131  , \reg2_reg[0]/NET0131  , \reg2_reg[10]/NET0131  , \reg2_reg[11]/NET0131  , \reg2_reg[12]/NET0131  , \reg2_reg[13]/NET0131  , \reg2_reg[14]/NET0131  , \reg2_reg[15]/NET0131  , \reg2_reg[16]/NET0131  , \reg2_reg[17]/NET0131  , \reg2_reg[18]/NET0131  , \reg2_reg[19]/NET0131  , \reg2_reg[1]/NET0131  , \reg2_reg[20]/NET0131  , \reg2_reg[21]/NET0131  , \reg2_reg[22]/NET0131  , \reg2_reg[23]/NET0131  , \reg2_reg[24]/NET0131  , \reg2_reg[25]/NET0131  , \reg2_reg[26]/NET0131  , \reg2_reg[27]/NET0131  , \reg2_reg[28]/NET0131  , \reg2_reg[29]/NET0131  , \reg2_reg[2]/NET0131  , \reg2_reg[30]/NET0131  , \reg2_reg[31]/NET0131  , \reg2_reg[3]/NET0131  , \reg2_reg[4]/NET0131  , \reg2_reg[5]/NET0131  , \reg2_reg[6]/NET0131  , \reg2_reg[7]/NET0131  , \reg2_reg[8]/NET0131  , \reg2_reg[9]/NET0131  , \reg3_reg[0]/NET0131  , \reg3_reg[10]/NET0131  , \reg3_reg[11]/NET0131  , \reg3_reg[12]/NET0131  , \reg3_reg[13]/NET0131  , \reg3_reg[14]/NET0131  , \reg3_reg[15]/NET0131  , \reg3_reg[16]/NET0131  , \reg3_reg[17]/NET0131  , \reg3_reg[18]/NET0131  , \reg3_reg[19]/NET0131  , \reg3_reg[1]/NET0131  , \reg3_reg[20]/NET0131  , \reg3_reg[21]/NET0131  , \reg3_reg[22]/NET0131  , \reg3_reg[23]/NET0131  , \reg3_reg[24]/NET0131  , \reg3_reg[25]/NET0131  , \reg3_reg[26]/NET0131  , \reg3_reg[27]/NET0131  , \reg3_reg[28]/NET0131  , \reg3_reg[2]/NET0131  , \reg3_reg[3]/NET0131  , \reg3_reg[4]/NET0131  , \reg3_reg[5]/NET0131  , \reg3_reg[6]/NET0131  , \reg3_reg[7]/NET0131  , \reg3_reg[8]/NET0131  , \reg3_reg[9]/NET0131  , \state_reg[0]/NET0131  , \_al_n0  , \_al_n1  , \g22/_0_  , \g32_dup/_0_  , \g35904/_0_  , \g35905/_0_  , \g35906/_0_  , \g35907/_0_  , \g35908/_0_  , \g35909/_0_  , \g35910/_0_  , \g35911/_0_  , \g35932/_0_  , \g35955/_0_  , \g35956/_0_  , \g35957/_0_  , \g35962/_0_  , \g35967/_0_  , \g35968/_0_  , \g35971/_0_  , \g35972/_0_  , \g35973/_0_  , \g35974/_0_  , \g35975/_0_  , \g35976/_0_  , \g35977/_0_  , \g35978/_0_  , \g36015/_0_  , \g36016/_0_  , \g36018/_0_  , \g36022/_0_  , \g36023/_0_  , \g36025/_0_  , \g36029/_0_  , \g36030/_0_  , \g36031/_0_  , \g36032/_0_  , \g36033/_0_  , \g36034/_0_  , \g36035/_0_  , \g36036/_0_  , \g36038/_0_  , \g36039/_0_  , \g36040/_0_  , \g36041/_0_  , \g36073/_0_  , \g36087/_0_  , \g36091/_0_  , \g36092/_0_  , \g36093/_0_  , \g36094/_0_  , \g36096/_0_  , \g36097/_0_  , \g36098/_0_  , \g36099/_0_  , \g36100/_0_  , \g36101/_0_  , \g36102/_0_  , \g36103/_0_  , \g36104/_0_  , \g36105/_0_  , \g36106/_0_  , \g36107/_0_  , \g36108/_0_  , \g36109/_0_  , \g36110/_0_  , \g36111/_0_  , \g36112/_0_  , \g36113/_0_  , \g36165/_0_  , \g36169/_0_  , \g36170/_0_  , \g36171/_0_  , \g36172/_0_  , \g36198/_0_  , \g36199/_0_  , \g36200/_0_  , \g36201/_0_  , \g36202/_0_  , \g36203/_0_  , \g36205/_0_  , \g36206/_0_  , \g36207/_0_  , \g36208/_0_  , \g36209/_0_  , \g36240/_0_  , \g36281/_0_  , \g36282/_0_  , \g36283/_0_  , \g36284/_0_  , \g36285/_0_  , \g36286/_0_  , \g36287/_0_  , \g36288/_0_  , \g36289/_0_  , \g36290/_0_  , \g36291/_0_  , \g36292/_0_  , \g36293/_0_  , \g36294/_0_  , \g36295/_0_  , \g36296/_0_  , \g36297/_0_  , \g36298/_0_  , \g36330/_0_  , \g36385/_0_  , \g36390/_0_  , \g36391/_0_  , \g36392/_0_  , \g36393/_0_  , \g36394/_0_  , \g36470/_0_  , \g36471/_0_  , \g36472/_0_  , \g36473/_0_  , \g36474/_0_  , \g36475/_0_  , \g38/_0_  , \g38399/_0_  , \g38400/_0_  , \g39639/_0_  , \g39641/_0_  , \g39644/_0_  , \g39647/_0_  , \g39648/_0_  , \g39650/_0_  , \g39654/_0_  , \g39658/_0_  , \g39660/_0_  , \g39662/_0_  , \g39663/_0_  , \g39665/_0_  , \g39666/_0_  , \g39667/_0_  , \g39730/_0_  , \g39796/_0_  , \g39930/_0_  , \g39931/_0_  , \g39932/_0_  , \g40045/_0_  , \g40150/u3_syn_4  , \g40608/_0_  , \g41017/u3_syn_4  , \g42159/_0_  , \g42169/_0_  , \g42174/_0_  , \g42483/_0_  , \g42736/_0_  , \g42746/_0_  , \g42755/_0_  , \g42767/_0_  , \g42776/_0_  , \g42871_dup/_1_  , \g42908/_0_  , \g42938/_0_  , \g42969/_0_  , \g43022/_0_  , \g44035/_1__syn_2  , \g44227/_3_  , \g44260/_3_  , \g44261/_3_  , \g44262/_3_  , \g44311/_3_  , \g44378/_3_  , \g44379/_3_  , \g44383/_3_  , \g44384/_3_  , \g44385/_3_  , \g44386/_3_  , \g44390/_3_  , \g44391/_3_  , \g44492/_3_  , \g44493/_3_  , \g44494/_3_  , \g44495/_3_  , \g44496/_3_  , \g44497/_3_  , \g44498/_3_  , \g44499/_3_  , \g44575/_3_  , \g44589/_3_  , \g44596/_3_  , \g44615/_3_  , \g44795/_3_  , \g44803/_3_  , \g44804/_3_  , \g44888/_3_  , \g44889/_3_  , \g45004/_3_  , \g46129/_0_  , \g46133/_0_  , \g46265/_2_  , \g46313/_0_  , \g46372/_0_  , \g46377/_0_  , \g46399/_0_  , \g46405/_0_  , \g46427/_0_  , \g46461/_0_  , \g46526/_0_  , \g46576/_0_  , \g46608/_0_  , \g46697/_0_  , \g46778/_0_  , \g47007/_0_  , \g47023/_0_  , \g47077/_1_  , \g47097/_0_  , \g47109/_1_  , \g47142_dup/_1_  , \g47256/_0_  , \g47328/_0_  , \g47373/_0_  , \g47465/_0_  , \g47518/_0_  , \g47556/_1_  , \g56/_0_  , \state_reg[0]/NET0131_syn_2  );
  input \B_reg/NET0131  ;
  input \IR_reg[0]/NET0131  ;
  input \IR_reg[10]/NET0131  ;
  input \IR_reg[11]/NET0131  ;
  input \IR_reg[12]/NET0131  ;
  input \IR_reg[13]/NET0131  ;
  input \IR_reg[14]/NET0131  ;
  input \IR_reg[15]/NET0131  ;
  input \IR_reg[16]/NET0131  ;
  input \IR_reg[17]/NET0131  ;
  input \IR_reg[18]/NET0131  ;
  input \IR_reg[19]/NET0131  ;
  input \IR_reg[1]/NET0131  ;
  input \IR_reg[20]/NET0131  ;
  input \IR_reg[21]/NET0131  ;
  input \IR_reg[22]/NET0131  ;
  input \IR_reg[23]/NET0131  ;
  input \IR_reg[24]/NET0131  ;
  input \IR_reg[25]/NET0131  ;
  input \IR_reg[26]/NET0131  ;
  input \IR_reg[27]/NET0131  ;
  input \IR_reg[28]/NET0131  ;
  input \IR_reg[29]/NET0131  ;
  input \IR_reg[2]/NET0131  ;
  input \IR_reg[30]/NET0131  ;
  input \IR_reg[31]/NET0131  ;
  input \IR_reg[3]/NET0131  ;
  input \IR_reg[4]/NET0131  ;
  input \IR_reg[5]/NET0131  ;
  input \IR_reg[6]/NET0131  ;
  input \IR_reg[7]/NET0131  ;
  input \IR_reg[8]/NET0131  ;
  input \IR_reg[9]/NET0131  ;
  input \addr[0]_pad  ;
  input \addr[10]_pad  ;
  input \addr[11]_pad  ;
  input \addr[12]_pad  ;
  input \addr[13]_pad  ;
  input \addr[14]_pad  ;
  input \addr[15]_pad  ;
  input \addr[16]_pad  ;
  input \addr[17]_pad  ;
  input \addr[18]_pad  ;
  input \addr[19]_pad  ;
  input \addr[1]_pad  ;
  input \addr[2]_pad  ;
  input \addr[3]_pad  ;
  input \addr[4]_pad  ;
  input \addr[5]_pad  ;
  input \addr[6]_pad  ;
  input \addr[7]_pad  ;
  input \addr[8]_pad  ;
  input \addr[9]_pad  ;
  input \d_reg[0]/NET0131  ;
  input \d_reg[1]/NET0131  ;
  input \datai[0]_pad  ;
  input \datai[10]_pad  ;
  input \datai[11]_pad  ;
  input \datai[12]_pad  ;
  input \datai[13]_pad  ;
  input \datai[14]_pad  ;
  input \datai[15]_pad  ;
  input \datai[16]_pad  ;
  input \datai[17]_pad  ;
  input \datai[18]_pad  ;
  input \datai[19]_pad  ;
  input \datai[1]_pad  ;
  input \datai[20]_pad  ;
  input \datai[21]_pad  ;
  input \datai[22]_pad  ;
  input \datai[23]_pad  ;
  input \datai[24]_pad  ;
  input \datai[25]_pad  ;
  input \datai[26]_pad  ;
  input \datai[27]_pad  ;
  input \datai[28]_pad  ;
  input \datai[29]_pad  ;
  input \datai[2]_pad  ;
  input \datai[30]_pad  ;
  input \datai[31]_pad  ;
  input \datai[3]_pad  ;
  input \datai[4]_pad  ;
  input \datai[5]_pad  ;
  input \datai[6]_pad  ;
  input \datai[7]_pad  ;
  input \datai[8]_pad  ;
  input \datai[9]_pad  ;
  input \datao[15]_pad  ;
  input \datao[28]_pad  ;
  input \datao[8]_pad  ;
  input \reg0_reg[0]/NET0131  ;
  input \reg0_reg[10]/NET0131  ;
  input \reg0_reg[11]/NET0131  ;
  input \reg0_reg[12]/NET0131  ;
  input \reg0_reg[13]/NET0131  ;
  input \reg0_reg[14]/NET0131  ;
  input \reg0_reg[15]/NET0131  ;
  input \reg0_reg[16]/NET0131  ;
  input \reg0_reg[17]/NET0131  ;
  input \reg0_reg[18]/NET0131  ;
  input \reg0_reg[19]/NET0131  ;
  input \reg0_reg[1]/NET0131  ;
  input \reg0_reg[20]/NET0131  ;
  input \reg0_reg[21]/NET0131  ;
  input \reg0_reg[22]/NET0131  ;
  input \reg0_reg[23]/NET0131  ;
  input \reg0_reg[24]/NET0131  ;
  input \reg0_reg[25]/NET0131  ;
  input \reg0_reg[26]/NET0131  ;
  input \reg0_reg[27]/NET0131  ;
  input \reg0_reg[28]/NET0131  ;
  input \reg0_reg[29]/NET0131  ;
  input \reg0_reg[2]/NET0131  ;
  input \reg0_reg[30]/NET0131  ;
  input \reg0_reg[31]/NET0131  ;
  input \reg0_reg[3]/NET0131  ;
  input \reg0_reg[4]/NET0131  ;
  input \reg0_reg[5]/NET0131  ;
  input \reg0_reg[6]/NET0131  ;
  input \reg0_reg[7]/NET0131  ;
  input \reg0_reg[8]/NET0131  ;
  input \reg0_reg[9]/NET0131  ;
  input \reg1_reg[0]/NET0131  ;
  input \reg1_reg[10]/NET0131  ;
  input \reg1_reg[11]/NET0131  ;
  input \reg1_reg[12]/NET0131  ;
  input \reg1_reg[13]/NET0131  ;
  input \reg1_reg[14]/NET0131  ;
  input \reg1_reg[15]/NET0131  ;
  input \reg1_reg[16]/NET0131  ;
  input \reg1_reg[17]/NET0131  ;
  input \reg1_reg[18]/NET0131  ;
  input \reg1_reg[19]/NET0131  ;
  input \reg1_reg[1]/NET0131  ;
  input \reg1_reg[20]/NET0131  ;
  input \reg1_reg[21]/NET0131  ;
  input \reg1_reg[22]/NET0131  ;
  input \reg1_reg[23]/NET0131  ;
  input \reg1_reg[24]/NET0131  ;
  input \reg1_reg[25]/NET0131  ;
  input \reg1_reg[26]/NET0131  ;
  input \reg1_reg[27]/NET0131  ;
  input \reg1_reg[28]/NET0131  ;
  input \reg1_reg[29]/NET0131  ;
  input \reg1_reg[2]/NET0131  ;
  input \reg1_reg[30]/NET0131  ;
  input \reg1_reg[31]/NET0131  ;
  input \reg1_reg[3]/NET0131  ;
  input \reg1_reg[4]/NET0131  ;
  input \reg1_reg[5]/NET0131  ;
  input \reg1_reg[6]/NET0131  ;
  input \reg1_reg[7]/NET0131  ;
  input \reg1_reg[8]/NET0131  ;
  input \reg1_reg[9]/NET0131  ;
  input \reg2_reg[0]/NET0131  ;
  input \reg2_reg[10]/NET0131  ;
  input \reg2_reg[11]/NET0131  ;
  input \reg2_reg[12]/NET0131  ;
  input \reg2_reg[13]/NET0131  ;
  input \reg2_reg[14]/NET0131  ;
  input \reg2_reg[15]/NET0131  ;
  input \reg2_reg[16]/NET0131  ;
  input \reg2_reg[17]/NET0131  ;
  input \reg2_reg[18]/NET0131  ;
  input \reg2_reg[19]/NET0131  ;
  input \reg2_reg[1]/NET0131  ;
  input \reg2_reg[20]/NET0131  ;
  input \reg2_reg[21]/NET0131  ;
  input \reg2_reg[22]/NET0131  ;
  input \reg2_reg[23]/NET0131  ;
  input \reg2_reg[24]/NET0131  ;
  input \reg2_reg[25]/NET0131  ;
  input \reg2_reg[26]/NET0131  ;
  input \reg2_reg[27]/NET0131  ;
  input \reg2_reg[28]/NET0131  ;
  input \reg2_reg[29]/NET0131  ;
  input \reg2_reg[2]/NET0131  ;
  input \reg2_reg[30]/NET0131  ;
  input \reg2_reg[31]/NET0131  ;
  input \reg2_reg[3]/NET0131  ;
  input \reg2_reg[4]/NET0131  ;
  input \reg2_reg[5]/NET0131  ;
  input \reg2_reg[6]/NET0131  ;
  input \reg2_reg[7]/NET0131  ;
  input \reg2_reg[8]/NET0131  ;
  input \reg2_reg[9]/NET0131  ;
  input \reg3_reg[0]/NET0131  ;
  input \reg3_reg[10]/NET0131  ;
  input \reg3_reg[11]/NET0131  ;
  input \reg3_reg[12]/NET0131  ;
  input \reg3_reg[13]/NET0131  ;
  input \reg3_reg[14]/NET0131  ;
  input \reg3_reg[15]/NET0131  ;
  input \reg3_reg[16]/NET0131  ;
  input \reg3_reg[17]/NET0131  ;
  input \reg3_reg[18]/NET0131  ;
  input \reg3_reg[19]/NET0131  ;
  input \reg3_reg[1]/NET0131  ;
  input \reg3_reg[20]/NET0131  ;
  input \reg3_reg[21]/NET0131  ;
  input \reg3_reg[22]/NET0131  ;
  input \reg3_reg[23]/NET0131  ;
  input \reg3_reg[24]/NET0131  ;
  input \reg3_reg[25]/NET0131  ;
  input \reg3_reg[26]/NET0131  ;
  input \reg3_reg[27]/NET0131  ;
  input \reg3_reg[28]/NET0131  ;
  input \reg3_reg[2]/NET0131  ;
  input \reg3_reg[3]/NET0131  ;
  input \reg3_reg[4]/NET0131  ;
  input \reg3_reg[5]/NET0131  ;
  input \reg3_reg[6]/NET0131  ;
  input \reg3_reg[7]/NET0131  ;
  input \reg3_reg[8]/NET0131  ;
  input \reg3_reg[9]/NET0131  ;
  input \state_reg[0]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g22/_0_  ;
  output \g32_dup/_0_  ;
  output \g35904/_0_  ;
  output \g35905/_0_  ;
  output \g35906/_0_  ;
  output \g35907/_0_  ;
  output \g35908/_0_  ;
  output \g35909/_0_  ;
  output \g35910/_0_  ;
  output \g35911/_0_  ;
  output \g35932/_0_  ;
  output \g35955/_0_  ;
  output \g35956/_0_  ;
  output \g35957/_0_  ;
  output \g35962/_0_  ;
  output \g35967/_0_  ;
  output \g35968/_0_  ;
  output \g35971/_0_  ;
  output \g35972/_0_  ;
  output \g35973/_0_  ;
  output \g35974/_0_  ;
  output \g35975/_0_  ;
  output \g35976/_0_  ;
  output \g35977/_0_  ;
  output \g35978/_0_  ;
  output \g36015/_0_  ;
  output \g36016/_0_  ;
  output \g36018/_0_  ;
  output \g36022/_0_  ;
  output \g36023/_0_  ;
  output \g36025/_0_  ;
  output \g36029/_0_  ;
  output \g36030/_0_  ;
  output \g36031/_0_  ;
  output \g36032/_0_  ;
  output \g36033/_0_  ;
  output \g36034/_0_  ;
  output \g36035/_0_  ;
  output \g36036/_0_  ;
  output \g36038/_0_  ;
  output \g36039/_0_  ;
  output \g36040/_0_  ;
  output \g36041/_0_  ;
  output \g36073/_0_  ;
  output \g36087/_0_  ;
  output \g36091/_0_  ;
  output \g36092/_0_  ;
  output \g36093/_0_  ;
  output \g36094/_0_  ;
  output \g36096/_0_  ;
  output \g36097/_0_  ;
  output \g36098/_0_  ;
  output \g36099/_0_  ;
  output \g36100/_0_  ;
  output \g36101/_0_  ;
  output \g36102/_0_  ;
  output \g36103/_0_  ;
  output \g36104/_0_  ;
  output \g36105/_0_  ;
  output \g36106/_0_  ;
  output \g36107/_0_  ;
  output \g36108/_0_  ;
  output \g36109/_0_  ;
  output \g36110/_0_  ;
  output \g36111/_0_  ;
  output \g36112/_0_  ;
  output \g36113/_0_  ;
  output \g36165/_0_  ;
  output \g36169/_0_  ;
  output \g36170/_0_  ;
  output \g36171/_0_  ;
  output \g36172/_0_  ;
  output \g36198/_0_  ;
  output \g36199/_0_  ;
  output \g36200/_0_  ;
  output \g36201/_0_  ;
  output \g36202/_0_  ;
  output \g36203/_0_  ;
  output \g36205/_0_  ;
  output \g36206/_0_  ;
  output \g36207/_0_  ;
  output \g36208/_0_  ;
  output \g36209/_0_  ;
  output \g36240/_0_  ;
  output \g36281/_0_  ;
  output \g36282/_0_  ;
  output \g36283/_0_  ;
  output \g36284/_0_  ;
  output \g36285/_0_  ;
  output \g36286/_0_  ;
  output \g36287/_0_  ;
  output \g36288/_0_  ;
  output \g36289/_0_  ;
  output \g36290/_0_  ;
  output \g36291/_0_  ;
  output \g36292/_0_  ;
  output \g36293/_0_  ;
  output \g36294/_0_  ;
  output \g36295/_0_  ;
  output \g36296/_0_  ;
  output \g36297/_0_  ;
  output \g36298/_0_  ;
  output \g36330/_0_  ;
  output \g36385/_0_  ;
  output \g36390/_0_  ;
  output \g36391/_0_  ;
  output \g36392/_0_  ;
  output \g36393/_0_  ;
  output \g36394/_0_  ;
  output \g36470/_0_  ;
  output \g36471/_0_  ;
  output \g36472/_0_  ;
  output \g36473/_0_  ;
  output \g36474/_0_  ;
  output \g36475/_0_  ;
  output \g38/_0_  ;
  output \g38399/_0_  ;
  output \g38400/_0_  ;
  output \g39639/_0_  ;
  output \g39641/_0_  ;
  output \g39644/_0_  ;
  output \g39647/_0_  ;
  output \g39648/_0_  ;
  output \g39650/_0_  ;
  output \g39654/_0_  ;
  output \g39658/_0_  ;
  output \g39660/_0_  ;
  output \g39662/_0_  ;
  output \g39663/_0_  ;
  output \g39665/_0_  ;
  output \g39666/_0_  ;
  output \g39667/_0_  ;
  output \g39730/_0_  ;
  output \g39796/_0_  ;
  output \g39930/_0_  ;
  output \g39931/_0_  ;
  output \g39932/_0_  ;
  output \g40045/_0_  ;
  output \g40150/u3_syn_4  ;
  output \g40608/_0_  ;
  output \g41017/u3_syn_4  ;
  output \g42159/_0_  ;
  output \g42169/_0_  ;
  output \g42174/_0_  ;
  output \g42483/_0_  ;
  output \g42736/_0_  ;
  output \g42746/_0_  ;
  output \g42755/_0_  ;
  output \g42767/_0_  ;
  output \g42776/_0_  ;
  output \g42871_dup/_1_  ;
  output \g42908/_0_  ;
  output \g42938/_0_  ;
  output \g42969/_0_  ;
  output \g43022/_0_  ;
  output \g44035/_1__syn_2  ;
  output \g44227/_3_  ;
  output \g44260/_3_  ;
  output \g44261/_3_  ;
  output \g44262/_3_  ;
  output \g44311/_3_  ;
  output \g44378/_3_  ;
  output \g44379/_3_  ;
  output \g44383/_3_  ;
  output \g44384/_3_  ;
  output \g44385/_3_  ;
  output \g44386/_3_  ;
  output \g44390/_3_  ;
  output \g44391/_3_  ;
  output \g44492/_3_  ;
  output \g44493/_3_  ;
  output \g44494/_3_  ;
  output \g44495/_3_  ;
  output \g44496/_3_  ;
  output \g44497/_3_  ;
  output \g44498/_3_  ;
  output \g44499/_3_  ;
  output \g44575/_3_  ;
  output \g44589/_3_  ;
  output \g44596/_3_  ;
  output \g44615/_3_  ;
  output \g44795/_3_  ;
  output \g44803/_3_  ;
  output \g44804/_3_  ;
  output \g44888/_3_  ;
  output \g44889/_3_  ;
  output \g45004/_3_  ;
  output \g46129/_0_  ;
  output \g46133/_0_  ;
  output \g46265/_2_  ;
  output \g46313/_0_  ;
  output \g46372/_0_  ;
  output \g46377/_0_  ;
  output \g46399/_0_  ;
  output \g46405/_0_  ;
  output \g46427/_0_  ;
  output \g46461/_0_  ;
  output \g46526/_0_  ;
  output \g46576/_0_  ;
  output \g46608/_0_  ;
  output \g46697/_0_  ;
  output \g46778/_0_  ;
  output \g47007/_0_  ;
  output \g47023/_0_  ;
  output \g47077/_1_  ;
  output \g47097/_0_  ;
  output \g47109/_1_  ;
  output \g47142_dup/_1_  ;
  output \g47256/_0_  ;
  output \g47328/_0_  ;
  output \g47373/_0_  ;
  output \g47465/_0_  ;
  output \g47518/_0_  ;
  output \g47556/_1_  ;
  output \g56/_0_  ;
  output \state_reg[0]/NET0131_syn_2  ;
  wire n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 ;
  assign n218 = \reg3_reg[3]/NET0131  & \reg3_reg[4]/NET0131  ;
  assign n219 = \reg3_reg[5]/NET0131  & n218 ;
  assign n220 = \reg3_reg[6]/NET0131  & n219 ;
  assign n221 = \reg3_reg[7]/NET0131  & n220 ;
  assign n222 = \reg3_reg[8]/NET0131  & n221 ;
  assign n223 = \reg3_reg[9]/NET0131  & n222 ;
  assign n224 = \reg3_reg[10]/NET0131  & n223 ;
  assign n225 = \reg3_reg[11]/NET0131  & n224 ;
  assign n226 = \reg3_reg[12]/NET0131  & n225 ;
  assign n227 = \reg3_reg[13]/NET0131  & \reg3_reg[14]/NET0131  ;
  assign n228 = \reg3_reg[15]/NET0131  & \reg3_reg[16]/NET0131  ;
  assign n229 = n227 & n228 ;
  assign n230 = n226 & n229 ;
  assign n231 = ~\reg3_reg[17]/NET0131  & ~n230 ;
  assign n232 = \reg3_reg[17]/NET0131  & n230 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = ~\IR_reg[20]/NET0131  & ~\IR_reg[21]/NET0131  ;
  assign n235 = ~\IR_reg[14]/NET0131  & ~\IR_reg[15]/NET0131  ;
  assign n236 = ~\IR_reg[0]/NET0131  & ~\IR_reg[1]/NET0131  ;
  assign n237 = ~\IR_reg[2]/NET0131  & ~\IR_reg[3]/NET0131  ;
  assign n238 = n236 & n237 ;
  assign n239 = ~\IR_reg[4]/NET0131  & n238 ;
  assign n240 = ~\IR_reg[5]/NET0131  & ~\IR_reg[6]/NET0131  ;
  assign n241 = ~\IR_reg[7]/NET0131  & n240 ;
  assign n242 = n239 & n241 ;
  assign n243 = ~\IR_reg[10]/NET0131  & ~\IR_reg[9]/NET0131  ;
  assign n244 = ~\IR_reg[11]/NET0131  & ~\IR_reg[8]/NET0131  ;
  assign n245 = n243 & n244 ;
  assign n246 = ~\IR_reg[12]/NET0131  & n245 ;
  assign n247 = ~\IR_reg[13]/NET0131  & n246 ;
  assign n248 = n242 & n247 ;
  assign n249 = n235 & n248 ;
  assign n250 = ~\IR_reg[16]/NET0131  & ~\IR_reg[17]/NET0131  ;
  assign n251 = ~\IR_reg[18]/NET0131  & n250 ;
  assign n252 = ~\IR_reg[19]/NET0131  & n251 ;
  assign n253 = n249 & n252 ;
  assign n254 = n234 & n253 ;
  assign n255 = ~\IR_reg[22]/NET0131  & n254 ;
  assign n256 = \IR_reg[31]/NET0131  & ~n255 ;
  assign n257 = ~\IR_reg[23]/NET0131  & ~n256 ;
  assign n258 = \IR_reg[23]/NET0131  & n256 ;
  assign n259 = ~n257 & ~n258 ;
  assign n282 = \IR_reg[31]/NET0131  & ~n249 ;
  assign n262 = ~\IR_reg[22]/NET0131  & ~\IR_reg[23]/NET0131  ;
  assign n263 = n234 & n262 ;
  assign n264 = n252 & n263 ;
  assign n283 = \IR_reg[31]/NET0131  & ~n264 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = \IR_reg[24]/NET0131  & ~n284 ;
  assign n286 = ~\IR_reg[24]/NET0131  & n284 ;
  assign n287 = ~n285 & ~n286 ;
  assign n265 = ~\IR_reg[24]/NET0131  & ~\IR_reg[25]/NET0131  ;
  assign n266 = n235 & n265 ;
  assign n267 = n264 & n266 ;
  assign n268 = n248 & n267 ;
  assign n269 = \IR_reg[31]/NET0131  & ~n268 ;
  assign n270 = \IR_reg[26]/NET0131  & ~n269 ;
  assign n271 = ~\IR_reg[26]/NET0131  & n269 ;
  assign n272 = ~n270 & ~n271 ;
  assign n273 = n242 & n246 ;
  assign n274 = ~\IR_reg[13]/NET0131  & ~\IR_reg[24]/NET0131  ;
  assign n275 = n235 & n274 ;
  assign n276 = n264 & n275 ;
  assign n277 = n273 & n276 ;
  assign n278 = \IR_reg[31]/NET0131  & ~n277 ;
  assign n279 = \IR_reg[25]/NET0131  & ~n278 ;
  assign n280 = ~\IR_reg[25]/NET0131  & n278 ;
  assign n281 = ~n279 & ~n280 ;
  assign n288 = ~n272 & ~n281 ;
  assign n289 = n287 & n288 ;
  assign n290 = ~n259 & n289 ;
  assign n291 = n233 & n290 ;
  assign n292 = ~n259 & ~n289 ;
  assign n293 = \B_reg/NET0131  & ~n287 ;
  assign n294 = n281 & n293 ;
  assign n295 = ~\d_reg[0]/NET0131  & ~n294 ;
  assign n296 = ~n272 & ~n295 ;
  assign n297 = ~\B_reg/NET0131  & n281 ;
  assign n298 = ~n272 & ~n297 ;
  assign n299 = n287 & ~n298 ;
  assign n300 = ~n296 & ~n299 ;
  assign n301 = n272 & n281 ;
  assign n302 = ~\B_reg/NET0131  & n287 ;
  assign n303 = ~n293 & ~n302 ;
  assign n304 = n281 & ~n303 ;
  assign n305 = ~\d_reg[1]/NET0131  & ~n272 ;
  assign n306 = ~n304 & n305 ;
  assign n307 = ~n301 & ~n306 ;
  assign n308 = ~n300 & n307 ;
  assign n358 = n233 & ~n308 ;
  assign n334 = ~\IR_reg[26]/NET0131  & ~\IR_reg[27]/NET0131  ;
  assign n335 = n265 & n334 ;
  assign n336 = n264 & n335 ;
  assign n337 = \IR_reg[31]/NET0131  & ~n336 ;
  assign n338 = ~n282 & ~n337 ;
  assign n339 = \IR_reg[28]/NET0131  & ~n338 ;
  assign n340 = ~\IR_reg[28]/NET0131  & n338 ;
  assign n341 = ~n339 & ~n340 ;
  assign n359 = ~\IR_reg[28]/NET0131  & n334 ;
  assign n360 = ~\IR_reg[25]/NET0131  & n359 ;
  assign n361 = n277 & n360 ;
  assign n362 = \IR_reg[31]/NET0131  & ~n361 ;
  assign n363 = \IR_reg[29]/NET0131  & n362 ;
  assign n364 = ~\IR_reg[29]/NET0131  & ~n362 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = ~\IR_reg[29]/NET0131  & n359 ;
  assign n367 = \IR_reg[31]/NET0131  & ~n366 ;
  assign n368 = ~n269 & ~n367 ;
  assign n369 = \IR_reg[30]/NET0131  & ~n368 ;
  assign n370 = ~\IR_reg[30]/NET0131  & n368 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = ~n365 & n371 ;
  assign n373 = \reg2_reg[2]/NET0131  & n372 ;
  assign n374 = n365 & ~n371 ;
  assign n375 = \reg1_reg[2]/NET0131  & n374 ;
  assign n380 = ~n373 & ~n375 ;
  assign n376 = ~n365 & ~n371 ;
  assign n377 = \reg0_reg[2]/NET0131  & n376 ;
  assign n378 = n365 & n371 ;
  assign n379 = \reg3_reg[2]/NET0131  & n378 ;
  assign n381 = ~n377 & ~n379 ;
  assign n382 = n380 & n381 ;
  assign n383 = \reg1_reg[1]/NET0131  & n374 ;
  assign n384 = \reg0_reg[1]/NET0131  & n376 ;
  assign n387 = ~n383 & ~n384 ;
  assign n385 = \reg2_reg[1]/NET0131  & n372 ;
  assign n386 = \reg3_reg[1]/NET0131  & n378 ;
  assign n388 = ~n385 & ~n386 ;
  assign n389 = n387 & n388 ;
  assign n390 = \reg1_reg[0]/NET0131  & n374 ;
  assign n391 = \reg0_reg[0]/NET0131  & n376 ;
  assign n394 = ~n390 & ~n391 ;
  assign n392 = \reg3_reg[0]/NET0131  & n378 ;
  assign n393 = \reg2_reg[0]/NET0131  & n372 ;
  assign n395 = ~n392 & ~n393 ;
  assign n396 = n394 & n395 ;
  assign n397 = \reg3_reg[17]/NET0131  & \reg3_reg[18]/NET0131  ;
  assign n398 = n230 & n397 ;
  assign n399 = \reg3_reg[19]/NET0131  & \reg3_reg[20]/NET0131  ;
  assign n400 = \reg3_reg[21]/NET0131  & n399 ;
  assign n401 = \reg3_reg[22]/NET0131  & n400 ;
  assign n402 = \reg3_reg[23]/NET0131  & n401 ;
  assign n403 = \reg3_reg[24]/NET0131  & n402 ;
  assign n404 = n398 & n403 ;
  assign n405 = \reg3_reg[25]/NET0131  & \reg3_reg[26]/NET0131  ;
  assign n406 = \reg3_reg[27]/NET0131  & \reg3_reg[28]/NET0131  ;
  assign n407 = n405 & n406 ;
  assign n408 = n404 & n407 ;
  assign n409 = n378 & n408 ;
  assign n412 = \reg0_reg[31]/NET0131  & n376 ;
  assign n410 = \reg1_reg[31]/NET0131  & n374 ;
  assign n411 = \reg2_reg[31]/NET0131  & n372 ;
  assign n413 = ~n410 & ~n411 ;
  assign n414 = ~n412 & n413 ;
  assign n415 = ~n409 & n414 ;
  assign n416 = ~n396 & ~n415 ;
  assign n417 = ~n389 & n416 ;
  assign n418 = ~n382 & n417 ;
  assign n419 = ~\reg3_reg[3]/NET0131  & n378 ;
  assign n420 = \reg2_reg[3]/NET0131  & n372 ;
  assign n423 = ~n419 & ~n420 ;
  assign n421 = \reg1_reg[3]/NET0131  & n374 ;
  assign n422 = \reg0_reg[3]/NET0131  & n376 ;
  assign n424 = ~n421 & ~n422 ;
  assign n425 = n423 & n424 ;
  assign n426 = ~\reg3_reg[3]/NET0131  & ~\reg3_reg[4]/NET0131  ;
  assign n427 = ~n218 & ~n426 ;
  assign n428 = n378 & n427 ;
  assign n429 = \reg1_reg[4]/NET0131  & n374 ;
  assign n432 = ~n428 & ~n429 ;
  assign n430 = \reg2_reg[4]/NET0131  & n372 ;
  assign n431 = \reg0_reg[4]/NET0131  & n376 ;
  assign n433 = ~n430 & ~n431 ;
  assign n434 = n432 & n433 ;
  assign n435 = ~n425 & ~n434 ;
  assign n436 = n418 & n435 ;
  assign n437 = \reg1_reg[6]/NET0131  & n374 ;
  assign n438 = \reg0_reg[6]/NET0131  & n376 ;
  assign n443 = ~n437 & ~n438 ;
  assign n439 = \reg2_reg[6]/NET0131  & n372 ;
  assign n440 = ~\reg3_reg[6]/NET0131  & ~n219 ;
  assign n441 = ~n220 & ~n440 ;
  assign n442 = n378 & n441 ;
  assign n444 = ~n439 & ~n442 ;
  assign n445 = n443 & n444 ;
  assign n446 = ~\reg3_reg[5]/NET0131  & ~n218 ;
  assign n447 = ~n219 & ~n446 ;
  assign n448 = n378 & n447 ;
  assign n449 = \reg1_reg[5]/NET0131  & n374 ;
  assign n452 = ~n448 & ~n449 ;
  assign n450 = \reg0_reg[5]/NET0131  & n376 ;
  assign n451 = \reg2_reg[5]/NET0131  & n372 ;
  assign n453 = ~n450 & ~n451 ;
  assign n454 = n452 & n453 ;
  assign n455 = ~n445 & ~n454 ;
  assign n456 = n436 & n455 ;
  assign n475 = \reg1_reg[7]/NET0131  & n374 ;
  assign n476 = \reg0_reg[7]/NET0131  & n376 ;
  assign n481 = ~n475 & ~n476 ;
  assign n477 = \reg2_reg[7]/NET0131  & n372 ;
  assign n478 = ~\reg3_reg[7]/NET0131  & ~n220 ;
  assign n479 = ~n221 & ~n478 ;
  assign n480 = n378 & n479 ;
  assign n482 = ~n477 & ~n480 ;
  assign n483 = n481 & n482 ;
  assign n457 = \reg0_reg[8]/NET0131  & n376 ;
  assign n458 = \reg1_reg[8]/NET0131  & n374 ;
  assign n463 = ~n457 & ~n458 ;
  assign n459 = ~\reg3_reg[8]/NET0131  & ~n221 ;
  assign n460 = ~n222 & ~n459 ;
  assign n461 = n378 & n460 ;
  assign n462 = \reg2_reg[8]/NET0131  & n372 ;
  assign n464 = ~n461 & ~n462 ;
  assign n465 = n463 & n464 ;
  assign n466 = \reg1_reg[9]/NET0131  & n374 ;
  assign n467 = \reg0_reg[9]/NET0131  & n376 ;
  assign n472 = ~n466 & ~n467 ;
  assign n468 = ~\reg3_reg[9]/NET0131  & ~n222 ;
  assign n469 = ~n223 & ~n468 ;
  assign n470 = n378 & n469 ;
  assign n471 = \reg2_reg[9]/NET0131  & n372 ;
  assign n473 = ~n470 & ~n471 ;
  assign n474 = n472 & n473 ;
  assign n484 = ~n465 & ~n474 ;
  assign n485 = ~n483 & n484 ;
  assign n486 = n456 & n485 ;
  assign n487 = ~\reg3_reg[12]/NET0131  & ~n225 ;
  assign n488 = ~n226 & ~n487 ;
  assign n489 = n378 & n488 ;
  assign n490 = \reg2_reg[12]/NET0131  & n372 ;
  assign n493 = ~n489 & ~n490 ;
  assign n491 = \reg0_reg[12]/NET0131  & n376 ;
  assign n492 = \reg1_reg[12]/NET0131  & n374 ;
  assign n494 = ~n491 & ~n492 ;
  assign n495 = n493 & n494 ;
  assign n496 = \reg0_reg[11]/NET0131  & n376 ;
  assign n497 = \reg1_reg[11]/NET0131  & n374 ;
  assign n502 = ~n496 & ~n497 ;
  assign n498 = \reg2_reg[11]/NET0131  & n372 ;
  assign n499 = ~\reg3_reg[11]/NET0131  & ~n224 ;
  assign n500 = ~n225 & ~n499 ;
  assign n501 = n378 & n500 ;
  assign n503 = ~n498 & ~n501 ;
  assign n504 = n502 & n503 ;
  assign n505 = \reg2_reg[10]/NET0131  & n372 ;
  assign n506 = \reg1_reg[10]/NET0131  & n374 ;
  assign n511 = ~n505 & ~n506 ;
  assign n507 = ~\reg3_reg[10]/NET0131  & ~n223 ;
  assign n508 = ~n224 & ~n507 ;
  assign n509 = n378 & n508 ;
  assign n510 = \reg0_reg[10]/NET0131  & n376 ;
  assign n512 = ~n509 & ~n510 ;
  assign n513 = n511 & n512 ;
  assign n514 = ~n504 & ~n513 ;
  assign n515 = ~n495 & n514 ;
  assign n516 = n486 & n515 ;
  assign n517 = \reg3_reg[13]/NET0131  & n226 ;
  assign n530 = \reg3_reg[14]/NET0131  & n517 ;
  assign n531 = \reg3_reg[15]/NET0131  & n530 ;
  assign n550 = ~\reg3_reg[16]/NET0131  & ~n531 ;
  assign n551 = ~n230 & ~n550 ;
  assign n552 = n378 & n551 ;
  assign n549 = \reg0_reg[16]/NET0131  & n376 ;
  assign n547 = \reg2_reg[16]/NET0131  & n372 ;
  assign n548 = \reg1_reg[16]/NET0131  & n374 ;
  assign n553 = ~n547 & ~n548 ;
  assign n554 = ~n549 & n553 ;
  assign n555 = ~n552 & n554 ;
  assign n541 = ~\reg3_reg[14]/NET0131  & ~n517 ;
  assign n542 = ~n530 & ~n541 ;
  assign n543 = n378 & n542 ;
  assign n540 = \reg2_reg[14]/NET0131  & n372 ;
  assign n538 = \reg0_reg[14]/NET0131  & n376 ;
  assign n539 = \reg1_reg[14]/NET0131  & n374 ;
  assign n544 = ~n538 & ~n539 ;
  assign n545 = ~n540 & n544 ;
  assign n546 = ~n543 & n545 ;
  assign n518 = ~\reg3_reg[13]/NET0131  & ~n226 ;
  assign n519 = ~n517 & ~n518 ;
  assign n520 = n378 & n519 ;
  assign n521 = \reg1_reg[13]/NET0131  & n374 ;
  assign n524 = ~n520 & ~n521 ;
  assign n522 = \reg2_reg[13]/NET0131  & n372 ;
  assign n523 = \reg0_reg[13]/NET0131  & n376 ;
  assign n525 = ~n522 & ~n523 ;
  assign n526 = n524 & n525 ;
  assign n532 = ~\reg3_reg[15]/NET0131  & ~n530 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = n378 & n533 ;
  assign n529 = \reg2_reg[15]/NET0131  & n372 ;
  assign n527 = \reg0_reg[15]/NET0131  & n376 ;
  assign n528 = \reg1_reg[15]/NET0131  & n374 ;
  assign n535 = ~n527 & ~n528 ;
  assign n536 = ~n529 & n535 ;
  assign n537 = ~n534 & n536 ;
  assign n556 = ~n526 & ~n537 ;
  assign n557 = ~n546 & n556 ;
  assign n558 = ~n555 & n557 ;
  assign n559 = n516 & n558 ;
  assign n563 = n233 & n378 ;
  assign n562 = \reg0_reg[17]/NET0131  & n376 ;
  assign n560 = \reg1_reg[17]/NET0131  & n374 ;
  assign n561 = \reg2_reg[17]/NET0131  & n372 ;
  assign n564 = ~n560 & ~n561 ;
  assign n565 = ~n562 & n564 ;
  assign n566 = ~n563 & n565 ;
  assign n567 = n559 & ~n566 ;
  assign n571 = ~\reg3_reg[18]/NET0131  & ~n232 ;
  assign n572 = ~n398 & ~n571 ;
  assign n573 = n378 & n572 ;
  assign n570 = \reg2_reg[18]/NET0131  & n372 ;
  assign n568 = \reg1_reg[18]/NET0131  & n374 ;
  assign n569 = \reg0_reg[18]/NET0131  & n376 ;
  assign n574 = ~n568 & ~n569 ;
  assign n575 = ~n570 & n574 ;
  assign n576 = ~n573 & n575 ;
  assign n577 = ~n567 & n576 ;
  assign n578 = ~n566 & ~n576 ;
  assign n579 = n559 & n578 ;
  assign n580 = ~n577 & ~n579 ;
  assign n581 = ~n341 & ~n580 ;
  assign n582 = n341 & n555 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n308 & n583 ;
  assign n585 = ~n358 & ~n584 ;
  assign n313 = \IR_reg[31]/NET0131  & ~n253 ;
  assign n314 = \IR_reg[20]/NET0131  & \IR_reg[31]/NET0131  ;
  assign n315 = ~n313 & ~n314 ;
  assign n316 = \IR_reg[21]/NET0131  & ~n315 ;
  assign n317 = ~\IR_reg[21]/NET0131  & n315 ;
  assign n318 = ~n316 & ~n317 ;
  assign n320 = ~\IR_reg[20]/NET0131  & ~n313 ;
  assign n321 = ~n253 & n314 ;
  assign n322 = ~n320 & ~n321 ;
  assign n586 = n318 & ~n322 ;
  assign n309 = \IR_reg[22]/NET0131  & ~\IR_reg[31]/NET0131  ;
  assign n310 = \IR_reg[22]/NET0131  & ~n254 ;
  assign n311 = n256 & ~n310 ;
  assign n312 = ~n309 & ~n311 ;
  assign n323 = \IR_reg[31]/NET0131  & ~n251 ;
  assign n324 = ~n282 & ~n323 ;
  assign n325 = \IR_reg[19]/NET0131  & ~n324 ;
  assign n326 = ~\IR_reg[19]/NET0131  & n324 ;
  assign n327 = ~n325 & ~n326 ;
  assign n587 = ~n312 & ~n327 ;
  assign n588 = n586 & n587 ;
  assign n589 = ~n585 & n588 ;
  assign n342 = ~\IR_reg[25]/NET0131  & ~\IR_reg[26]/NET0131  ;
  assign n343 = \IR_reg[31]/NET0131  & ~n342 ;
  assign n344 = ~n278 & ~n343 ;
  assign n345 = \IR_reg[27]/NET0131  & ~n344 ;
  assign n346 = ~\IR_reg[27]/NET0131  & n344 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n341 & ~n347 ;
  assign n349 = \IR_reg[16]/NET0131  & \IR_reg[31]/NET0131  ;
  assign n350 = ~n282 & ~n349 ;
  assign n351 = \IR_reg[17]/NET0131  & ~n350 ;
  assign n352 = ~\IR_reg[17]/NET0131  & n350 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = n348 & ~n353 ;
  assign n355 = ~\datai[17]_pad  & ~n348 ;
  assign n356 = ~n354 & ~n355 ;
  assign n590 = ~n356 & n566 ;
  assign n591 = n356 & ~n566 ;
  assign n592 = ~n590 & ~n591 ;
  assign n593 = ~\IR_reg[8]/NET0131  & n242 ;
  assign n594 = \IR_reg[31]/NET0131  & ~n593 ;
  assign n595 = \IR_reg[31]/NET0131  & ~n243 ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = \IR_reg[11]/NET0131  & ~n596 ;
  assign n598 = ~\IR_reg[11]/NET0131  & n596 ;
  assign n599 = ~n597 & ~n598 ;
  assign n600 = n348 & n599 ;
  assign n601 = \datai[11]_pad  & ~n348 ;
  assign n602 = ~n600 & ~n601 ;
  assign n603 = n504 & ~n602 ;
  assign n604 = \IR_reg[31]/NET0131  & ~n242 ;
  assign n605 = \IR_reg[31]/NET0131  & ~n245 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = \IR_reg[12]/NET0131  & ~n606 ;
  assign n608 = ~\IR_reg[12]/NET0131  & n606 ;
  assign n609 = ~n607 & ~n608 ;
  assign n610 = n348 & n609 ;
  assign n611 = \datai[12]_pad  & ~n348 ;
  assign n612 = ~n610 & ~n611 ;
  assign n613 = n495 & ~n612 ;
  assign n614 = ~n603 & ~n613 ;
  assign n615 = \IR_reg[31]/NET0131  & \IR_reg[9]/NET0131  ;
  assign n616 = ~n594 & ~n615 ;
  assign n617 = \IR_reg[10]/NET0131  & ~n616 ;
  assign n618 = ~\IR_reg[10]/NET0131  & n616 ;
  assign n619 = ~n617 & ~n618 ;
  assign n620 = n348 & n619 ;
  assign n621 = \datai[10]_pad  & ~n348 ;
  assign n622 = ~n620 & ~n621 ;
  assign n623 = n513 & ~n622 ;
  assign n624 = ~n513 & n622 ;
  assign n625 = \IR_reg[9]/NET0131  & ~n594 ;
  assign n626 = ~\IR_reg[9]/NET0131  & n594 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = n348 & ~n627 ;
  assign n629 = \datai[9]_pad  & ~n348 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = ~n474 & n630 ;
  assign n632 = ~n624 & ~n631 ;
  assign n633 = ~n623 & ~n632 ;
  assign n634 = n614 & n633 ;
  assign n635 = ~n495 & n612 ;
  assign n636 = ~n504 & n602 ;
  assign n637 = ~n635 & ~n636 ;
  assign n638 = ~n613 & ~n637 ;
  assign n639 = ~n634 & ~n638 ;
  assign n640 = \IR_reg[31]/NET0131  & ~n248 ;
  assign n641 = \IR_reg[14]/NET0131  & ~n640 ;
  assign n642 = ~\IR_reg[14]/NET0131  & n640 ;
  assign n643 = ~n641 & ~n642 ;
  assign n644 = n348 & ~n643 ;
  assign n645 = \datai[14]_pad  & ~n348 ;
  assign n646 = ~n644 & ~n645 ;
  assign n647 = n546 & ~n646 ;
  assign n648 = \IR_reg[31]/NET0131  & ~n273 ;
  assign n649 = \IR_reg[13]/NET0131  & n648 ;
  assign n650 = ~\IR_reg[13]/NET0131  & ~n648 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = n348 & n651 ;
  assign n653 = \datai[13]_pad  & ~n348 ;
  assign n654 = ~n652 & ~n653 ;
  assign n655 = n526 & ~n654 ;
  assign n656 = ~n647 & ~n655 ;
  assign n657 = \datai[16]_pad  & ~n348 ;
  assign n658 = ~\IR_reg[16]/NET0131  & ~n282 ;
  assign n659 = ~n249 & n349 ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = n348 & n660 ;
  assign n662 = ~n657 & ~n661 ;
  assign n663 = n555 & ~n662 ;
  assign n664 = \IR_reg[14]/NET0131  & \IR_reg[31]/NET0131  ;
  assign n665 = ~n640 & ~n664 ;
  assign n666 = \IR_reg[15]/NET0131  & ~n665 ;
  assign n667 = ~\IR_reg[15]/NET0131  & n665 ;
  assign n668 = ~n666 & ~n667 ;
  assign n669 = n348 & ~n668 ;
  assign n670 = ~\datai[15]_pad  & ~n348 ;
  assign n671 = ~n669 & ~n670 ;
  assign n672 = n537 & n671 ;
  assign n673 = ~n663 & ~n672 ;
  assign n674 = n656 & n673 ;
  assign n675 = ~n639 & n674 ;
  assign n676 = ~n546 & n646 ;
  assign n677 = ~n526 & n654 ;
  assign n678 = ~n676 & ~n677 ;
  assign n679 = ~n647 & ~n678 ;
  assign n680 = n673 & n679 ;
  assign n681 = ~n555 & n662 ;
  assign n682 = ~n537 & ~n671 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = ~n663 & ~n683 ;
  assign n685 = ~n680 & ~n684 ;
  assign n686 = ~n675 & n685 ;
  assign n687 = n474 & ~n630 ;
  assign n688 = ~n623 & ~n687 ;
  assign n689 = n614 & n688 ;
  assign n690 = \IR_reg[31]/NET0131  & ~n239 ;
  assign n691 = \IR_reg[31]/NET0131  & ~n240 ;
  assign n692 = ~n690 & ~n691 ;
  assign n693 = \IR_reg[7]/NET0131  & ~n692 ;
  assign n694 = ~\IR_reg[7]/NET0131  & n692 ;
  assign n695 = ~n693 & ~n694 ;
  assign n696 = n348 & n695 ;
  assign n697 = \datai[7]_pad  & ~n348 ;
  assign n698 = ~n696 & ~n697 ;
  assign n699 = n483 & ~n698 ;
  assign n700 = ~\IR_reg[8]/NET0131  & ~n604 ;
  assign n701 = \IR_reg[8]/NET0131  & n604 ;
  assign n702 = ~n700 & ~n701 ;
  assign n703 = n348 & n702 ;
  assign n704 = \datai[8]_pad  & ~n348 ;
  assign n705 = ~n703 & ~n704 ;
  assign n706 = n465 & ~n705 ;
  assign n707 = ~n699 & ~n706 ;
  assign n708 = \IR_reg[31]/NET0131  & \IR_reg[5]/NET0131  ;
  assign n709 = ~n690 & ~n708 ;
  assign n710 = \IR_reg[6]/NET0131  & ~n709 ;
  assign n711 = ~\IR_reg[6]/NET0131  & n709 ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = n348 & n712 ;
  assign n714 = \datai[6]_pad  & ~n348 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = n445 & ~n715 ;
  assign n717 = ~n445 & n715 ;
  assign n718 = \datai[5]_pad  & ~n348 ;
  assign n719 = ~\IR_reg[5]/NET0131  & ~n690 ;
  assign n720 = ~n239 & n708 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = n348 & n721 ;
  assign n723 = ~n718 & ~n722 ;
  assign n724 = ~n454 & n723 ;
  assign n725 = ~n717 & ~n724 ;
  assign n726 = ~n716 & ~n725 ;
  assign n727 = n707 & n726 ;
  assign n728 = ~n465 & n705 ;
  assign n729 = ~n483 & n698 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~n706 & ~n730 ;
  assign n732 = ~n727 & ~n731 ;
  assign n733 = \IR_reg[31]/NET0131  & ~n238 ;
  assign n734 = \IR_reg[4]/NET0131  & ~n733 ;
  assign n735 = ~\IR_reg[4]/NET0131  & n733 ;
  assign n736 = ~n734 & ~n735 ;
  assign n737 = n348 & ~n736 ;
  assign n738 = \datai[4]_pad  & ~n348 ;
  assign n739 = ~n737 & ~n738 ;
  assign n740 = n434 & ~n739 ;
  assign n741 = \IR_reg[0]/NET0131  & \IR_reg[31]/NET0131  ;
  assign n742 = ~\IR_reg[1]/NET0131  & ~n741 ;
  assign n743 = \IR_reg[1]/NET0131  & n741 ;
  assign n744 = ~n742 & ~n743 ;
  assign n745 = n348 & n744 ;
  assign n746 = \datai[1]_pad  & ~n348 ;
  assign n747 = ~n745 & ~n746 ;
  assign n748 = n389 & ~n747 ;
  assign n749 = \datai[0]_pad  & ~n348 ;
  assign n750 = \IR_reg[0]/NET0131  & n348 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = n396 & ~n751 ;
  assign n753 = ~n748 & ~n752 ;
  assign n754 = ~n389 & n747 ;
  assign n755 = \datai[2]_pad  & ~n348 ;
  assign n756 = \IR_reg[31]/NET0131  & ~n236 ;
  assign n757 = \IR_reg[2]/NET0131  & ~n756 ;
  assign n758 = ~\IR_reg[2]/NET0131  & n756 ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = n348 & ~n759 ;
  assign n761 = ~n755 & ~n760 ;
  assign n762 = ~n382 & n761 ;
  assign n763 = ~n754 & ~n762 ;
  assign n764 = ~n753 & n763 ;
  assign n765 = \IR_reg[2]/NET0131  & \IR_reg[31]/NET0131  ;
  assign n766 = ~n756 & ~n765 ;
  assign n767 = \IR_reg[3]/NET0131  & ~n766 ;
  assign n768 = ~\IR_reg[3]/NET0131  & n766 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = n348 & n769 ;
  assign n771 = \datai[3]_pad  & ~n348 ;
  assign n772 = ~n770 & ~n771 ;
  assign n773 = n425 & ~n772 ;
  assign n774 = n382 & ~n761 ;
  assign n775 = ~n773 & ~n774 ;
  assign n776 = ~n764 & n775 ;
  assign n777 = ~n425 & n772 ;
  assign n778 = ~n434 & n739 ;
  assign n779 = ~n777 & ~n778 ;
  assign n780 = ~n776 & n779 ;
  assign n781 = ~n740 & ~n780 ;
  assign n782 = n454 & ~n723 ;
  assign n783 = ~n716 & ~n782 ;
  assign n784 = n707 & n783 ;
  assign n785 = n781 & n784 ;
  assign n786 = n732 & ~n785 ;
  assign n787 = n689 & ~n786 ;
  assign n788 = n674 & n787 ;
  assign n789 = n686 & ~n788 ;
  assign n790 = n592 & ~n789 ;
  assign n791 = ~n592 & n789 ;
  assign n792 = ~n790 & ~n791 ;
  assign n793 = n308 & ~n792 ;
  assign n794 = ~n358 & ~n793 ;
  assign n795 = ~n586 & ~n587 ;
  assign n319 = n312 & ~n318 ;
  assign n796 = ~n312 & n318 ;
  assign n797 = ~n319 & ~n796 ;
  assign n798 = n795 & n797 ;
  assign n799 = ~n794 & n798 ;
  assign n328 = ~n322 & n327 ;
  assign n329 = n319 & n328 ;
  assign n330 = ~n308 & ~n329 ;
  assign n331 = ~n322 & ~n327 ;
  assign n332 = n319 & ~n331 ;
  assign n333 = ~n330 & n332 ;
  assign n357 = n333 & n356 ;
  assign n909 = ~n331 & n796 ;
  assign n910 = n319 & n322 ;
  assign n911 = ~n308 & n910 ;
  assign n912 = ~n909 & ~n911 ;
  assign n913 = n233 & ~n912 ;
  assign n914 = ~n357 & ~n913 ;
  assign n915 = ~n799 & n914 ;
  assign n800 = n555 & n662 ;
  assign n801 = n537 & ~n671 ;
  assign n802 = ~n800 & ~n801 ;
  assign n803 = ~n546 & ~n646 ;
  assign n804 = n546 & n646 ;
  assign n805 = ~n526 & ~n654 ;
  assign n806 = ~n804 & n805 ;
  assign n807 = ~n803 & ~n806 ;
  assign n808 = n802 & ~n807 ;
  assign n809 = ~n555 & ~n662 ;
  assign n810 = ~n537 & n671 ;
  assign n811 = ~n809 & ~n810 ;
  assign n812 = ~n800 & ~n811 ;
  assign n813 = ~n808 & ~n812 ;
  assign n814 = n526 & n654 ;
  assign n815 = ~n804 & ~n814 ;
  assign n816 = n802 & n815 ;
  assign n817 = n504 & n602 ;
  assign n818 = n495 & n612 ;
  assign n819 = ~n817 & ~n818 ;
  assign n820 = n513 & n622 ;
  assign n821 = ~n513 & ~n622 ;
  assign n822 = ~n474 & ~n630 ;
  assign n823 = ~n821 & ~n822 ;
  assign n824 = ~n820 & ~n823 ;
  assign n825 = n819 & n824 ;
  assign n826 = ~n495 & ~n612 ;
  assign n827 = ~n504 & ~n602 ;
  assign n828 = ~n818 & n827 ;
  assign n829 = ~n826 & ~n828 ;
  assign n830 = ~n825 & n829 ;
  assign n831 = n816 & ~n830 ;
  assign n832 = n813 & ~n831 ;
  assign n833 = n474 & n630 ;
  assign n834 = ~n820 & ~n833 ;
  assign n835 = n819 & n834 ;
  assign n836 = n465 & n705 ;
  assign n837 = n483 & n698 ;
  assign n838 = ~n836 & ~n837 ;
  assign n839 = ~n445 & ~n715 ;
  assign n840 = n445 & n715 ;
  assign n841 = ~n454 & ~n723 ;
  assign n842 = ~n840 & n841 ;
  assign n843 = ~n839 & ~n842 ;
  assign n844 = n838 & ~n843 ;
  assign n845 = ~n465 & ~n705 ;
  assign n846 = ~n483 & ~n698 ;
  assign n847 = ~n845 & ~n846 ;
  assign n848 = ~n836 & ~n847 ;
  assign n849 = ~n844 & ~n848 ;
  assign n852 = ~n382 & ~n761 ;
  assign n853 = ~n389 & ~n747 ;
  assign n854 = n389 & n747 ;
  assign n855 = ~n396 & ~n751 ;
  assign n856 = ~n854 & n855 ;
  assign n857 = ~n853 & ~n856 ;
  assign n858 = ~n852 & n857 ;
  assign n859 = n425 & n772 ;
  assign n860 = n382 & n761 ;
  assign n861 = ~n859 & ~n860 ;
  assign n862 = n434 & n739 ;
  assign n863 = n861 & ~n862 ;
  assign n864 = ~n858 & n863 ;
  assign n865 = ~n434 & ~n739 ;
  assign n866 = ~n425 & ~n772 ;
  assign n867 = ~n865 & ~n866 ;
  assign n868 = ~n862 & ~n867 ;
  assign n869 = ~n864 & ~n868 ;
  assign n850 = n454 & n723 ;
  assign n851 = ~n840 & ~n850 ;
  assign n870 = n838 & n851 ;
  assign n871 = ~n869 & n870 ;
  assign n872 = n849 & ~n871 ;
  assign n873 = n835 & ~n872 ;
  assign n874 = n816 & n873 ;
  assign n875 = n832 & ~n874 ;
  assign n876 = n592 & ~n875 ;
  assign n877 = ~n592 & n875 ;
  assign n878 = ~n876 & ~n877 ;
  assign n879 = n308 & n878 ;
  assign n880 = ~n358 & ~n879 ;
  assign n881 = ~n795 & ~n796 ;
  assign n882 = ~n880 & n881 ;
  assign n883 = n747 & n751 ;
  assign n884 = n761 & n883 ;
  assign n885 = n772 & n884 ;
  assign n886 = n739 & n885 ;
  assign n887 = n723 & n886 ;
  assign n888 = n715 & n887 ;
  assign n889 = n698 & n888 ;
  assign n890 = n630 & n705 ;
  assign n891 = n889 & n890 ;
  assign n892 = n602 & n622 ;
  assign n893 = n612 & n654 ;
  assign n894 = n892 & n893 ;
  assign n895 = n891 & n894 ;
  assign n896 = n646 & n895 ;
  assign n897 = ~n671 & n896 ;
  assign n898 = n662 & n897 ;
  assign n899 = n356 & ~n898 ;
  assign n900 = ~n356 & n646 ;
  assign n901 = n662 & ~n671 ;
  assign n902 = n900 & n901 ;
  assign n903 = n895 & n902 ;
  assign n904 = ~n899 & ~n903 ;
  assign n905 = n308 & n904 ;
  assign n906 = ~n358 & ~n905 ;
  assign n907 = n319 & n331 ;
  assign n908 = ~n906 & n907 ;
  assign n916 = ~n882 & ~n908 ;
  assign n917 = n915 & n916 ;
  assign n918 = ~n589 & n917 ;
  assign n919 = n292 & ~n918 ;
  assign n920 = ~n291 & ~n919 ;
  assign n921 = \state_reg[0]/NET0131  & ~n920 ;
  assign n217 = \reg3_reg[17]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n260 = \state_reg[0]/NET0131  & n259 ;
  assign n261 = n233 & n260 ;
  assign n922 = ~n217 & ~n261 ;
  assign n923 = ~n921 & n922 ;
  assign n927 = n398 & n401 ;
  assign n928 = ~\reg3_reg[23]/NET0131  & ~n927 ;
  assign n929 = n398 & n402 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = n378 & n930 ;
  assign n926 = \reg2_reg[23]/NET0131  & n372 ;
  assign n924 = \reg0_reg[23]/NET0131  & n376 ;
  assign n925 = \reg1_reg[23]/NET0131  & n374 ;
  assign n932 = ~n924 & ~n925 ;
  assign n933 = ~n926 & n932 ;
  assign n934 = ~n931 & n933 ;
  assign n935 = \reg3_reg[25]/NET0131  & n404 ;
  assign n936 = \reg3_reg[26]/NET0131  & n935 ;
  assign n937 = \reg3_reg[27]/NET0131  & n936 ;
  assign n938 = ~\reg3_reg[28]/NET0131  & ~n937 ;
  assign n939 = \reg3_reg[28]/NET0131  & n937 ;
  assign n940 = ~n938 & ~n939 ;
  assign n941 = ~n308 & n940 ;
  assign n942 = \datai[27]_pad  & ~n348 ;
  assign n946 = ~\reg3_reg[27]/NET0131  & ~n936 ;
  assign n947 = ~n937 & ~n946 ;
  assign n948 = n378 & n947 ;
  assign n945 = \reg2_reg[27]/NET0131  & n372 ;
  assign n943 = \reg1_reg[27]/NET0131  & n374 ;
  assign n944 = \reg0_reg[27]/NET0131  & n376 ;
  assign n949 = ~n943 & ~n944 ;
  assign n950 = ~n945 & n949 ;
  assign n951 = ~n948 & n950 ;
  assign n952 = n942 & n951 ;
  assign n953 = \datai[26]_pad  & ~n348 ;
  assign n957 = ~\reg3_reg[26]/NET0131  & ~n935 ;
  assign n958 = ~n936 & ~n957 ;
  assign n959 = n378 & n958 ;
  assign n956 = \reg0_reg[26]/NET0131  & n376 ;
  assign n954 = \reg2_reg[26]/NET0131  & n372 ;
  assign n955 = \reg1_reg[26]/NET0131  & n374 ;
  assign n960 = ~n954 & ~n955 ;
  assign n961 = ~n956 & n960 ;
  assign n962 = ~n959 & n961 ;
  assign n963 = n953 & n962 ;
  assign n964 = ~n952 & ~n963 ;
  assign n965 = \datai[25]_pad  & ~n348 ;
  assign n969 = ~\reg3_reg[25]/NET0131  & ~n404 ;
  assign n970 = ~n935 & ~n969 ;
  assign n971 = n378 & n970 ;
  assign n968 = \reg2_reg[25]/NET0131  & n372 ;
  assign n966 = \reg0_reg[25]/NET0131  & n376 ;
  assign n967 = \reg1_reg[25]/NET0131  & n374 ;
  assign n972 = ~n966 & ~n967 ;
  assign n973 = ~n968 & n972 ;
  assign n974 = ~n971 & n973 ;
  assign n975 = n965 & n974 ;
  assign n976 = \datai[24]_pad  & ~n348 ;
  assign n980 = ~\reg3_reg[24]/NET0131  & ~n929 ;
  assign n981 = ~n404 & ~n980 ;
  assign n982 = n378 & n981 ;
  assign n979 = \reg2_reg[24]/NET0131  & n372 ;
  assign n977 = \reg1_reg[24]/NET0131  & n374 ;
  assign n978 = \reg0_reg[24]/NET0131  & n376 ;
  assign n983 = ~n977 & ~n978 ;
  assign n984 = ~n979 & n983 ;
  assign n985 = ~n982 & n984 ;
  assign n986 = n976 & n985 ;
  assign n987 = ~n975 & ~n986 ;
  assign n988 = n964 & n987 ;
  assign n989 = \datai[23]_pad  & ~n348 ;
  assign n990 = n934 & n989 ;
  assign n991 = \datai[22]_pad  & ~n348 ;
  assign n995 = n398 & n400 ;
  assign n996 = ~\reg3_reg[22]/NET0131  & ~n995 ;
  assign n997 = ~n927 & ~n996 ;
  assign n998 = n378 & n997 ;
  assign n994 = \reg1_reg[22]/NET0131  & n374 ;
  assign n992 = \reg0_reg[22]/NET0131  & n376 ;
  assign n993 = \reg2_reg[22]/NET0131  & n372 ;
  assign n999 = ~n992 & ~n993 ;
  assign n1000 = ~n994 & n999 ;
  assign n1001 = ~n998 & n1000 ;
  assign n1002 = n991 & n1001 ;
  assign n1003 = ~n990 & ~n1002 ;
  assign n1004 = \datai[21]_pad  & ~n348 ;
  assign n1008 = n398 & n399 ;
  assign n1009 = ~\reg3_reg[21]/NET0131  & ~n1008 ;
  assign n1010 = ~n995 & ~n1009 ;
  assign n1011 = n378 & n1010 ;
  assign n1007 = \reg2_reg[21]/NET0131  & n372 ;
  assign n1005 = \reg1_reg[21]/NET0131  & n374 ;
  assign n1006 = \reg0_reg[21]/NET0131  & n376 ;
  assign n1012 = ~n1005 & ~n1006 ;
  assign n1013 = ~n1007 & n1012 ;
  assign n1014 = ~n1011 & n1013 ;
  assign n1015 = n1004 & n1014 ;
  assign n1016 = \datai[20]_pad  & ~n348 ;
  assign n1020 = \reg3_reg[19]/NET0131  & n398 ;
  assign n1021 = ~\reg3_reg[20]/NET0131  & ~n1020 ;
  assign n1022 = ~n1008 & ~n1021 ;
  assign n1023 = n378 & n1022 ;
  assign n1019 = \reg1_reg[20]/NET0131  & n374 ;
  assign n1017 = \reg0_reg[20]/NET0131  & n376 ;
  assign n1018 = \reg2_reg[20]/NET0131  & n372 ;
  assign n1024 = ~n1017 & ~n1018 ;
  assign n1025 = ~n1019 & n1024 ;
  assign n1026 = ~n1023 & n1025 ;
  assign n1027 = n1016 & n1026 ;
  assign n1028 = ~n1015 & ~n1027 ;
  assign n1029 = n1003 & n1028 ;
  assign n1030 = n988 & n1029 ;
  assign n1031 = \IR_reg[31]/NET0131  & ~n250 ;
  assign n1032 = ~n282 & ~n1031 ;
  assign n1033 = \IR_reg[18]/NET0131  & ~n1032 ;
  assign n1034 = ~\IR_reg[18]/NET0131  & n1032 ;
  assign n1035 = ~n1033 & ~n1034 ;
  assign n1036 = n348 & ~n1035 ;
  assign n1037 = ~\datai[18]_pad  & ~n348 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = n576 & n1038 ;
  assign n1043 = ~\reg3_reg[19]/NET0131  & ~n398 ;
  assign n1044 = ~n1020 & ~n1043 ;
  assign n1045 = n378 & n1044 ;
  assign n1042 = \reg0_reg[19]/NET0131  & n376 ;
  assign n1040 = \reg1_reg[19]/NET0131  & n374 ;
  assign n1041 = \reg2_reg[19]/NET0131  & n372 ;
  assign n1046 = ~n1040 & ~n1041 ;
  assign n1047 = ~n1042 & n1046 ;
  assign n1048 = ~n1045 & n1047 ;
  assign n1049 = n327 & n348 ;
  assign n1050 = \datai[19]_pad  & ~n348 ;
  assign n1051 = ~n1049 & ~n1050 ;
  assign n1052 = n1048 & ~n1051 ;
  assign n1053 = ~n1039 & ~n1052 ;
  assign n1054 = n356 & n566 ;
  assign n1055 = ~n663 & ~n1054 ;
  assign n1056 = n1053 & n1055 ;
  assign n1074 = ~n603 & ~n623 ;
  assign n1075 = ~n631 & ~n728 ;
  assign n1076 = ~n687 & ~n1075 ;
  assign n1077 = n1074 & n1076 ;
  assign n1078 = ~n603 & n624 ;
  assign n1079 = ~n636 & ~n1078 ;
  assign n1080 = ~n1077 & n1079 ;
  assign n1081 = ~n699 & ~n716 ;
  assign n1082 = ~n753 & ~n754 ;
  assign n1083 = n775 & ~n1082 ;
  assign n1084 = ~n762 & ~n777 ;
  assign n1085 = ~n773 & ~n1084 ;
  assign n1086 = ~n1083 & ~n1085 ;
  assign n1087 = ~n740 & ~n782 ;
  assign n1088 = ~n1086 & n1087 ;
  assign n1089 = n1081 & n1088 ;
  assign n1090 = ~n724 & ~n778 ;
  assign n1091 = ~n782 & ~n1090 ;
  assign n1092 = n1081 & n1091 ;
  assign n1093 = ~n699 & n717 ;
  assign n1094 = ~n729 & ~n1093 ;
  assign n1095 = ~n1092 & n1094 ;
  assign n1096 = ~n1089 & n1095 ;
  assign n1097 = ~n687 & ~n706 ;
  assign n1098 = n1074 & n1097 ;
  assign n1099 = ~n1096 & n1098 ;
  assign n1100 = n1080 & ~n1099 ;
  assign n1057 = ~n647 & ~n672 ;
  assign n1101 = ~n613 & ~n655 ;
  assign n1102 = n1057 & n1101 ;
  assign n1103 = ~n1100 & n1102 ;
  assign n1104 = n1056 & n1103 ;
  assign n1058 = n635 & ~n655 ;
  assign n1059 = ~n677 & ~n1058 ;
  assign n1060 = n1057 & ~n1059 ;
  assign n1061 = ~n676 & ~n682 ;
  assign n1062 = ~n672 & ~n1061 ;
  assign n1063 = ~n1060 & ~n1062 ;
  assign n1064 = n1056 & ~n1063 ;
  assign n1065 = ~n356 & ~n566 ;
  assign n1066 = ~n681 & ~n1065 ;
  assign n1067 = ~n1054 & ~n1066 ;
  assign n1068 = n1053 & n1067 ;
  assign n1069 = ~n1048 & n1051 ;
  assign n1070 = ~n576 & ~n1038 ;
  assign n1071 = ~n1069 & ~n1070 ;
  assign n1072 = ~n1052 & ~n1071 ;
  assign n1073 = ~n1068 & ~n1072 ;
  assign n1105 = ~n1064 & n1073 ;
  assign n1106 = ~n1104 & n1105 ;
  assign n1107 = n1030 & ~n1106 ;
  assign n1108 = ~n1004 & ~n1014 ;
  assign n1109 = ~n1016 & ~n1026 ;
  assign n1110 = ~n1108 & ~n1109 ;
  assign n1111 = ~n1015 & ~n1110 ;
  assign n1112 = n1003 & n1111 ;
  assign n1113 = ~n934 & ~n989 ;
  assign n1114 = ~n991 & ~n1001 ;
  assign n1115 = ~n990 & n1114 ;
  assign n1116 = ~n1113 & ~n1115 ;
  assign n1117 = ~n1112 & n1116 ;
  assign n1118 = n988 & ~n1117 ;
  assign n1119 = ~n953 & ~n962 ;
  assign n1120 = ~n942 & ~n951 ;
  assign n1121 = ~n1119 & ~n1120 ;
  assign n1122 = ~n965 & ~n974 ;
  assign n1123 = ~n976 & ~n985 ;
  assign n1124 = ~n1122 & ~n1123 ;
  assign n1125 = ~n975 & ~n1124 ;
  assign n1126 = ~n963 & n1125 ;
  assign n1127 = n1121 & ~n1126 ;
  assign n1128 = ~n952 & ~n1127 ;
  assign n1129 = ~n1118 & ~n1128 ;
  assign n1130 = ~n1107 & n1129 ;
  assign n1131 = \datai[28]_pad  & ~n348 ;
  assign n1135 = n378 & n940 ;
  assign n1134 = \reg2_reg[28]/NET0131  & n372 ;
  assign n1132 = \reg1_reg[28]/NET0131  & n374 ;
  assign n1133 = \reg0_reg[28]/NET0131  & n376 ;
  assign n1136 = ~n1132 & ~n1133 ;
  assign n1137 = ~n1134 & n1136 ;
  assign n1138 = ~n1135 & n1137 ;
  assign n1139 = ~n1131 & n1138 ;
  assign n1140 = n1131 & ~n1138 ;
  assign n1141 = ~n1139 & ~n1140 ;
  assign n1142 = ~n1130 & n1141 ;
  assign n1143 = n1130 & ~n1141 ;
  assign n1144 = ~n1142 & ~n1143 ;
  assign n1145 = n308 & ~n1144 ;
  assign n1146 = ~n941 & ~n1145 ;
  assign n1147 = n798 & ~n1146 ;
  assign n1148 = ~n814 & ~n818 ;
  assign n1149 = ~n801 & ~n804 ;
  assign n1150 = n1148 & n1149 ;
  assign n1151 = ~n590 & ~n800 ;
  assign n1152 = n1048 & n1051 ;
  assign n1153 = n576 & ~n1038 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = n1151 & n1154 ;
  assign n1156 = n1150 & n1155 ;
  assign n1157 = ~n817 & ~n820 ;
  assign n1158 = ~n822 & ~n845 ;
  assign n1159 = ~n833 & ~n1158 ;
  assign n1160 = n1157 & n1159 ;
  assign n1161 = ~n817 & n821 ;
  assign n1162 = ~n827 & ~n1161 ;
  assign n1163 = ~n1160 & n1162 ;
  assign n1164 = ~n837 & ~n840 ;
  assign n1165 = ~n857 & n861 ;
  assign n1166 = ~n852 & ~n866 ;
  assign n1167 = ~n859 & ~n1166 ;
  assign n1168 = ~n1165 & ~n1167 ;
  assign n1169 = ~n850 & ~n862 ;
  assign n1170 = ~n1168 & n1169 ;
  assign n1171 = n1164 & n1170 ;
  assign n1172 = ~n850 & n865 ;
  assign n1173 = ~n841 & ~n1172 ;
  assign n1174 = n1164 & ~n1173 ;
  assign n1175 = ~n837 & n839 ;
  assign n1176 = ~n846 & ~n1175 ;
  assign n1177 = ~n1174 & n1176 ;
  assign n1178 = ~n1171 & n1177 ;
  assign n1179 = ~n833 & ~n836 ;
  assign n1180 = n1157 & n1179 ;
  assign n1181 = ~n1178 & n1180 ;
  assign n1182 = n1163 & ~n1181 ;
  assign n1183 = n1156 & ~n1182 ;
  assign n1184 = ~n814 & n826 ;
  assign n1185 = ~n805 & ~n1184 ;
  assign n1186 = n1149 & ~n1185 ;
  assign n1187 = ~n801 & n803 ;
  assign n1188 = ~n810 & ~n1187 ;
  assign n1189 = ~n1186 & n1188 ;
  assign n1190 = n1155 & ~n1189 ;
  assign n1191 = ~n590 & n809 ;
  assign n1192 = ~n591 & ~n1191 ;
  assign n1193 = n1154 & ~n1192 ;
  assign n1194 = ~n1048 & ~n1051 ;
  assign n1195 = ~n576 & n1038 ;
  assign n1196 = ~n1152 & n1195 ;
  assign n1197 = ~n1194 & ~n1196 ;
  assign n1198 = ~n1193 & n1197 ;
  assign n1199 = ~n1190 & n1198 ;
  assign n1200 = ~n1183 & n1199 ;
  assign n1201 = ~n1004 & n1014 ;
  assign n1202 = ~n1016 & n1026 ;
  assign n1203 = ~n1201 & ~n1202 ;
  assign n1204 = n934 & ~n989 ;
  assign n1205 = ~n991 & n1001 ;
  assign n1206 = ~n1204 & ~n1205 ;
  assign n1207 = n1203 & n1206 ;
  assign n1208 = ~n942 & n951 ;
  assign n1209 = ~n953 & n962 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1211 = ~n976 & n985 ;
  assign n1212 = ~n965 & n974 ;
  assign n1213 = ~n1211 & ~n1212 ;
  assign n1214 = n1210 & n1213 ;
  assign n1215 = n1207 & n1214 ;
  assign n1216 = ~n1200 & n1215 ;
  assign n1217 = n1004 & ~n1014 ;
  assign n1218 = n1016 & ~n1026 ;
  assign n1219 = ~n1201 & n1218 ;
  assign n1220 = ~n1217 & ~n1219 ;
  assign n1221 = n1206 & ~n1220 ;
  assign n1222 = ~n934 & n989 ;
  assign n1223 = n991 & ~n1001 ;
  assign n1224 = ~n1204 & n1223 ;
  assign n1225 = ~n1222 & ~n1224 ;
  assign n1226 = ~n1221 & n1225 ;
  assign n1227 = n1214 & ~n1226 ;
  assign n1228 = n942 & ~n951 ;
  assign n1229 = n953 & ~n962 ;
  assign n1230 = n965 & ~n974 ;
  assign n1231 = n976 & ~n985 ;
  assign n1232 = ~n1212 & n1231 ;
  assign n1233 = ~n1230 & ~n1232 ;
  assign n1234 = ~n1229 & n1233 ;
  assign n1235 = n1210 & ~n1234 ;
  assign n1236 = ~n1228 & ~n1235 ;
  assign n1237 = ~n1227 & n1236 ;
  assign n1238 = ~n1216 & n1237 ;
  assign n1239 = n1141 & n1238 ;
  assign n1240 = ~n1141 & ~n1238 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = n308 & ~n1241 ;
  assign n1243 = ~n941 & ~n1242 ;
  assign n1244 = n881 & ~n1243 ;
  assign n1245 = ~n953 & ~n965 ;
  assign n1246 = ~n1038 & n1051 ;
  assign n1247 = n903 & n1246 ;
  assign n1248 = ~n991 & ~n1004 ;
  assign n1249 = ~n1016 & n1248 ;
  assign n1250 = ~n989 & n1249 ;
  assign n1251 = ~n976 & n1250 ;
  assign n1252 = n1247 & n1251 ;
  assign n1253 = n1245 & n1252 ;
  assign n1254 = ~n942 & n1253 ;
  assign n1255 = n1131 & ~n1254 ;
  assign n1256 = ~n942 & ~n1131 ;
  assign n1257 = n1245 & n1256 ;
  assign n1258 = n1252 & n1257 ;
  assign n1259 = ~n1255 & ~n1258 ;
  assign n1260 = n308 & n1259 ;
  assign n1261 = ~n941 & ~n1260 ;
  assign n1262 = n907 & ~n1261 ;
  assign n1263 = ~n1001 & ~n1014 ;
  assign n1264 = ~n934 & ~n1026 ;
  assign n1265 = n1263 & n1264 ;
  assign n1266 = ~n985 & ~n1048 ;
  assign n1267 = n1265 & n1266 ;
  assign n1268 = ~n974 & n1267 ;
  assign n1269 = ~n951 & ~n962 ;
  assign n1270 = n578 & ~n1138 ;
  assign n1271 = n1269 & n1270 ;
  assign n1272 = n1268 & n1271 ;
  assign n1273 = n559 & n1272 ;
  assign n1276 = \reg1_reg[29]/NET0131  & n374 ;
  assign n1274 = \reg0_reg[29]/NET0131  & n376 ;
  assign n1275 = \reg2_reg[29]/NET0131  & n372 ;
  assign n1277 = ~n1274 & ~n1275 ;
  assign n1278 = ~n1276 & n1277 ;
  assign n1279 = ~n409 & n1278 ;
  assign n1280 = ~n1273 & ~n1279 ;
  assign n1281 = n1273 & n1279 ;
  assign n1282 = ~n1280 & ~n1281 ;
  assign n1283 = ~n341 & ~n1282 ;
  assign n1284 = n341 & ~n951 ;
  assign n1285 = ~n1283 & ~n1284 ;
  assign n1286 = n308 & ~n1285 ;
  assign n1287 = ~n941 & ~n1286 ;
  assign n1288 = n588 & ~n1287 ;
  assign n1289 = ~n912 & n940 ;
  assign n1290 = n333 & n1131 ;
  assign n1291 = ~n1289 & ~n1290 ;
  assign n1292 = ~n1288 & n1291 ;
  assign n1293 = ~n1262 & n1292 ;
  assign n1294 = ~n1244 & n1293 ;
  assign n1295 = ~n1147 & n1294 ;
  assign n1296 = n292 & ~n1295 ;
  assign n1297 = n290 & n940 ;
  assign n1298 = ~n1296 & ~n1297 ;
  assign n1299 = \state_reg[0]/NET0131  & ~n1298 ;
  assign n1300 = \reg3_reg[28]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1301 = n260 & n940 ;
  assign n1302 = ~n1300 & ~n1301 ;
  assign n1303 = ~n1299 & n1302 ;
  assign n1304 = ~n308 & n947 ;
  assign n1305 = ~n590 & ~n1153 ;
  assign n1306 = n802 & n1305 ;
  assign n1307 = n851 & ~n869 ;
  assign n1308 = n843 & ~n1307 ;
  assign n1309 = n834 & n838 ;
  assign n1310 = ~n1308 & n1309 ;
  assign n1311 = n834 & n848 ;
  assign n1312 = ~n824 & ~n1311 ;
  assign n1313 = ~n1310 & n1312 ;
  assign n1314 = n815 & n819 ;
  assign n1315 = ~n1313 & n1314 ;
  assign n1316 = n1306 & n1315 ;
  assign n1317 = n815 & ~n829 ;
  assign n1318 = n807 & ~n1317 ;
  assign n1319 = n1306 & ~n1318 ;
  assign n1320 = n812 & n1305 ;
  assign n1321 = n591 & ~n1153 ;
  assign n1322 = ~n1195 & ~n1321 ;
  assign n1323 = ~n1320 & n1322 ;
  assign n1324 = ~n1319 & n1323 ;
  assign n1325 = ~n1316 & n1324 ;
  assign n1326 = ~n1201 & ~n1205 ;
  assign n1327 = ~n1152 & ~n1202 ;
  assign n1328 = n1326 & n1327 ;
  assign n1329 = ~n1204 & ~n1211 ;
  assign n1330 = ~n1209 & ~n1212 ;
  assign n1331 = n1329 & n1330 ;
  assign n1332 = n1328 & n1331 ;
  assign n1333 = ~n1325 & n1332 ;
  assign n1334 = n1194 & ~n1202 ;
  assign n1335 = ~n1218 & ~n1334 ;
  assign n1336 = n1326 & ~n1335 ;
  assign n1337 = ~n1205 & n1217 ;
  assign n1338 = ~n1223 & ~n1337 ;
  assign n1339 = ~n1336 & n1338 ;
  assign n1340 = n1331 & ~n1339 ;
  assign n1341 = ~n1229 & ~n1230 ;
  assign n1342 = ~n1211 & n1222 ;
  assign n1343 = ~n1231 & ~n1342 ;
  assign n1344 = ~n1212 & ~n1343 ;
  assign n1345 = n1341 & ~n1344 ;
  assign n1346 = ~n1209 & ~n1345 ;
  assign n1347 = ~n1340 & ~n1346 ;
  assign n1348 = ~n1333 & n1347 ;
  assign n1349 = ~n1208 & ~n1228 ;
  assign n1350 = n1348 & n1349 ;
  assign n1351 = ~n1348 & ~n1349 ;
  assign n1352 = ~n1350 & ~n1351 ;
  assign n1353 = n308 & ~n1352 ;
  assign n1354 = ~n1304 & ~n1353 ;
  assign n1355 = n881 & ~n1354 ;
  assign n1356 = n781 & n783 ;
  assign n1357 = ~n726 & ~n1356 ;
  assign n1358 = n688 & n707 ;
  assign n1359 = ~n1357 & n1358 ;
  assign n1360 = n688 & n731 ;
  assign n1361 = ~n633 & ~n1360 ;
  assign n1362 = ~n1359 & n1361 ;
  assign n1363 = ~n1039 & ~n1054 ;
  assign n1364 = n673 & n1363 ;
  assign n1365 = n614 & n656 ;
  assign n1366 = n1364 & n1365 ;
  assign n1367 = ~n1362 & n1366 ;
  assign n1368 = n638 & n656 ;
  assign n1369 = ~n679 & ~n1368 ;
  assign n1370 = n1364 & ~n1369 ;
  assign n1371 = n684 & n1363 ;
  assign n1372 = ~n1065 & ~n1070 ;
  assign n1373 = ~n1039 & ~n1372 ;
  assign n1374 = ~n1371 & ~n1373 ;
  assign n1375 = ~n1370 & n1374 ;
  assign n1376 = ~n1367 & n1375 ;
  assign n1377 = ~n1027 & ~n1052 ;
  assign n1378 = ~n1002 & ~n1015 ;
  assign n1379 = n1377 & n1378 ;
  assign n1380 = ~n986 & ~n990 ;
  assign n1381 = ~n963 & ~n975 ;
  assign n1382 = n1380 & n1381 ;
  assign n1383 = n1379 & n1382 ;
  assign n1384 = ~n1376 & n1383 ;
  assign n1387 = ~n1069 & ~n1109 ;
  assign n1388 = ~n1027 & ~n1387 ;
  assign n1389 = n1378 & n1388 ;
  assign n1390 = ~n1108 & ~n1114 ;
  assign n1391 = ~n1002 & ~n1390 ;
  assign n1392 = ~n1389 & ~n1391 ;
  assign n1393 = n1382 & ~n1392 ;
  assign n1385 = ~n1119 & ~n1122 ;
  assign n1386 = ~n963 & ~n1385 ;
  assign n1394 = ~n986 & n1113 ;
  assign n1395 = ~n1123 & ~n1394 ;
  assign n1396 = n1381 & ~n1395 ;
  assign n1397 = ~n1386 & ~n1396 ;
  assign n1398 = ~n1393 & n1397 ;
  assign n1399 = ~n1384 & n1398 ;
  assign n1400 = n1349 & ~n1399 ;
  assign n1401 = ~n1349 & n1399 ;
  assign n1402 = ~n1400 & ~n1401 ;
  assign n1403 = n308 & ~n1402 ;
  assign n1404 = ~n1304 & ~n1403 ;
  assign n1405 = n798 & ~n1404 ;
  assign n1406 = n578 & ~n1048 ;
  assign n1407 = n558 & n1406 ;
  assign n1408 = n516 & n1407 ;
  assign n1409 = n1265 & n1408 ;
  assign n1410 = ~n974 & ~n985 ;
  assign n1411 = n1269 & n1410 ;
  assign n1412 = n1409 & n1411 ;
  assign n1413 = n1138 & ~n1412 ;
  assign n1414 = ~n1138 & n1412 ;
  assign n1415 = ~n1413 & ~n1414 ;
  assign n1416 = ~n341 & ~n1415 ;
  assign n1417 = n341 & n962 ;
  assign n1418 = ~n1416 & ~n1417 ;
  assign n1419 = n308 & n1418 ;
  assign n1420 = ~n1304 & ~n1419 ;
  assign n1421 = n588 & ~n1420 ;
  assign n1426 = n942 & ~n1253 ;
  assign n1427 = ~n1254 & ~n1426 ;
  assign n1428 = n907 & n1427 ;
  assign n1429 = n308 & n1428 ;
  assign n1422 = n319 & ~n328 ;
  assign n1423 = ~n308 & n1422 ;
  assign n1424 = ~n909 & ~n1423 ;
  assign n1425 = n947 & ~n1424 ;
  assign n1430 = n333 & n942 ;
  assign n1431 = ~n1425 & ~n1430 ;
  assign n1432 = ~n1429 & n1431 ;
  assign n1433 = ~n1421 & n1432 ;
  assign n1434 = ~n1405 & n1433 ;
  assign n1435 = ~n1355 & n1434 ;
  assign n1436 = n292 & ~n1435 ;
  assign n1437 = n290 & n947 ;
  assign n1438 = ~n1436 & ~n1437 ;
  assign n1439 = \state_reg[0]/NET0131  & ~n1438 ;
  assign n1440 = \reg3_reg[27]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1441 = n260 & n947 ;
  assign n1442 = ~n1440 & ~n1441 ;
  assign n1443 = ~n1439 & n1442 ;
  assign n1444 = n300 & ~n307 ;
  assign n1445 = \reg0_reg[27]/NET0131  & ~n1444 ;
  assign n1446 = ~n1352 & n1444 ;
  assign n1447 = ~n1445 & ~n1446 ;
  assign n1448 = n881 & ~n1447 ;
  assign n1449 = ~n1402 & n1444 ;
  assign n1450 = ~n1445 & ~n1449 ;
  assign n1451 = n798 & ~n1450 ;
  assign n1452 = n588 & n1418 ;
  assign n1453 = n910 & n942 ;
  assign n1454 = ~n1428 & ~n1453 ;
  assign n1455 = ~n1452 & n1454 ;
  assign n1456 = n1444 & ~n1455 ;
  assign n1457 = n910 & ~n1444 ;
  assign n1458 = ~n329 & ~n909 ;
  assign n1459 = ~n1457 & n1458 ;
  assign n1460 = n331 & ~n797 ;
  assign n1461 = ~n1444 & n1460 ;
  assign n1462 = n1459 & ~n1461 ;
  assign n1463 = \reg0_reg[27]/NET0131  & ~n1462 ;
  assign n1464 = ~n1456 & ~n1463 ;
  assign n1465 = ~n1451 & n1464 ;
  assign n1466 = ~n1448 & n1465 ;
  assign n1467 = n292 & ~n1466 ;
  assign n1468 = \reg0_reg[27]/NET0131  & n290 ;
  assign n1469 = ~n1467 & ~n1468 ;
  assign n1470 = \state_reg[0]/NET0131  & ~n1469 ;
  assign n1471 = \state_reg[0]/NET0131  & ~n259 ;
  assign n1472 = \reg0_reg[27]/NET0131  & ~n1471 ;
  assign n1473 = ~n1470 & ~n1472 ;
  assign n1474 = \reg0_reg[28]/NET0131  & ~n1444 ;
  assign n1475 = ~n1144 & n1444 ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1477 = n798 & ~n1476 ;
  assign n1478 = ~n1241 & n1444 ;
  assign n1479 = ~n1474 & ~n1478 ;
  assign n1480 = n881 & ~n1479 ;
  assign n1481 = n907 & n1259 ;
  assign n1482 = n910 & n1131 ;
  assign n1483 = n588 & ~n1285 ;
  assign n1484 = ~n1482 & ~n1483 ;
  assign n1485 = ~n1481 & n1484 ;
  assign n1486 = n1444 & ~n1485 ;
  assign n1487 = \reg0_reg[28]/NET0131  & ~n1462 ;
  assign n1488 = ~n1486 & ~n1487 ;
  assign n1489 = ~n1480 & n1488 ;
  assign n1490 = ~n1477 & n1489 ;
  assign n1491 = n292 & ~n1490 ;
  assign n1492 = \reg0_reg[28]/NET0131  & n290 ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1494 = \state_reg[0]/NET0131  & ~n1493 ;
  assign n1495 = \reg0_reg[28]/NET0131  & ~n1471 ;
  assign n1496 = ~n1494 & ~n1495 ;
  assign n1497 = ~n300 & ~n307 ;
  assign n1498 = \reg1_reg[27]/NET0131  & ~n1497 ;
  assign n1499 = ~n1352 & n1497 ;
  assign n1500 = ~n1498 & ~n1499 ;
  assign n1501 = n881 & ~n1500 ;
  assign n1502 = ~n1402 & n1497 ;
  assign n1503 = ~n1498 & ~n1502 ;
  assign n1504 = n798 & ~n1503 ;
  assign n1505 = ~n1455 & n1497 ;
  assign n1506 = n1422 & ~n1497 ;
  assign n1507 = n1458 & ~n1506 ;
  assign n1508 = n588 & ~n1497 ;
  assign n1509 = n1507 & ~n1508 ;
  assign n1510 = \reg1_reg[27]/NET0131  & ~n1509 ;
  assign n1511 = ~n1505 & ~n1510 ;
  assign n1512 = ~n1504 & n1511 ;
  assign n1513 = ~n1501 & n1512 ;
  assign n1514 = n292 & ~n1513 ;
  assign n1515 = \reg1_reg[27]/NET0131  & n290 ;
  assign n1516 = ~n1514 & ~n1515 ;
  assign n1517 = \state_reg[0]/NET0131  & ~n1516 ;
  assign n1518 = \reg1_reg[27]/NET0131  & ~n1471 ;
  assign n1519 = ~n1517 & ~n1518 ;
  assign n1520 = \reg1_reg[28]/NET0131  & ~n1497 ;
  assign n1521 = ~n1144 & n1497 ;
  assign n1522 = ~n1520 & ~n1521 ;
  assign n1523 = n798 & ~n1522 ;
  assign n1524 = ~n1241 & n1497 ;
  assign n1525 = ~n1520 & ~n1524 ;
  assign n1526 = n881 & ~n1525 ;
  assign n1527 = ~n1485 & n1497 ;
  assign n1528 = n910 & ~n1497 ;
  assign n1529 = n1458 & ~n1528 ;
  assign n1530 = n907 & ~n1497 ;
  assign n1531 = n1529 & ~n1530 ;
  assign n1532 = ~n1508 & n1531 ;
  assign n1533 = \reg1_reg[28]/NET0131  & ~n1532 ;
  assign n1534 = ~n1527 & ~n1533 ;
  assign n1535 = ~n1526 & n1534 ;
  assign n1536 = ~n1523 & n1535 ;
  assign n1537 = n292 & ~n1536 ;
  assign n1538 = \reg1_reg[28]/NET0131  & n290 ;
  assign n1539 = ~n1537 & ~n1538 ;
  assign n1540 = \state_reg[0]/NET0131  & ~n1539 ;
  assign n1541 = \reg1_reg[28]/NET0131  & ~n1471 ;
  assign n1542 = ~n1540 & ~n1541 ;
  assign n1543 = n300 & n307 ;
  assign n1544 = \reg2_reg[27]/NET0131  & ~n1543 ;
  assign n1545 = ~n1352 & n1543 ;
  assign n1546 = ~n1544 & ~n1545 ;
  assign n1547 = n881 & ~n1546 ;
  assign n1548 = ~n1402 & n1543 ;
  assign n1549 = ~n1544 & ~n1548 ;
  assign n1550 = n798 & ~n1549 ;
  assign n1551 = n1418 & n1543 ;
  assign n1552 = ~n1544 & ~n1551 ;
  assign n1553 = n588 & ~n1552 ;
  assign n1554 = n1427 & n1543 ;
  assign n1555 = ~n1544 & ~n1554 ;
  assign n1556 = n907 & ~n1555 ;
  assign n1559 = n910 & ~n1543 ;
  assign n1560 = ~n909 & ~n1559 ;
  assign n1561 = \reg2_reg[27]/NET0131  & ~n1560 ;
  assign n1557 = n329 & n947 ;
  assign n1558 = n1453 & n1543 ;
  assign n1562 = ~n1557 & ~n1558 ;
  assign n1563 = ~n1561 & n1562 ;
  assign n1564 = ~n1556 & n1563 ;
  assign n1565 = ~n1553 & n1564 ;
  assign n1566 = ~n1550 & n1565 ;
  assign n1567 = ~n1547 & n1566 ;
  assign n1568 = n292 & ~n1567 ;
  assign n1569 = \reg2_reg[27]/NET0131  & n290 ;
  assign n1570 = ~n1568 & ~n1569 ;
  assign n1571 = \state_reg[0]/NET0131  & ~n1570 ;
  assign n1572 = \reg2_reg[27]/NET0131  & ~n1471 ;
  assign n1573 = ~n1571 & ~n1572 ;
  assign n1574 = \reg2_reg[28]/NET0131  & ~n1543 ;
  assign n1575 = ~n1144 & n1543 ;
  assign n1576 = ~n1574 & ~n1575 ;
  assign n1577 = n798 & ~n1576 ;
  assign n1578 = ~n1241 & n1543 ;
  assign n1579 = ~n1574 & ~n1578 ;
  assign n1580 = n881 & ~n1579 ;
  assign n1581 = ~n1485 & n1543 ;
  assign n1582 = n329 & n940 ;
  assign n1583 = n588 & ~n1543 ;
  assign n1584 = n907 & ~n1543 ;
  assign n1585 = n1560 & ~n1584 ;
  assign n1586 = ~n1583 & n1585 ;
  assign n1587 = \reg2_reg[28]/NET0131  & ~n1586 ;
  assign n1588 = ~n1582 & ~n1587 ;
  assign n1589 = ~n1581 & n1588 ;
  assign n1590 = ~n1580 & n1589 ;
  assign n1591 = ~n1577 & n1590 ;
  assign n1592 = n292 & ~n1591 ;
  assign n1593 = \reg2_reg[28]/NET0131  & n290 ;
  assign n1594 = ~n1592 & ~n1593 ;
  assign n1595 = \state_reg[0]/NET0131  & ~n1594 ;
  assign n1596 = \reg2_reg[28]/NET0131  & ~n1471 ;
  assign n1597 = ~n1595 & ~n1596 ;
  assign n1600 = n290 & n533 ;
  assign n1602 = ~n308 & n533 ;
  assign n1619 = n516 & ~n526 ;
  assign n1620 = ~n546 & n1619 ;
  assign n1621 = ~n537 & n1620 ;
  assign n1622 = n555 & ~n1621 ;
  assign n1623 = ~n559 & ~n1622 ;
  assign n1624 = ~n341 & ~n1623 ;
  assign n1625 = n341 & n546 ;
  assign n1626 = ~n1624 & ~n1625 ;
  assign n1627 = n308 & n1626 ;
  assign n1628 = ~n1602 & ~n1627 ;
  assign n1629 = n588 & ~n1628 ;
  assign n1603 = ~n801 & ~n810 ;
  assign n1612 = ~n1315 & n1318 ;
  assign n1613 = n1603 & n1612 ;
  assign n1614 = ~n1603 & ~n1612 ;
  assign n1615 = ~n1613 & ~n1614 ;
  assign n1616 = n308 & ~n1615 ;
  assign n1617 = ~n1602 & ~n1616 ;
  assign n1618 = n881 & ~n1617 ;
  assign n1604 = ~n1362 & n1365 ;
  assign n1605 = n1369 & ~n1604 ;
  assign n1606 = n1603 & n1605 ;
  assign n1607 = ~n1603 & ~n1605 ;
  assign n1608 = ~n1606 & ~n1607 ;
  assign n1609 = n308 & n1608 ;
  assign n1610 = ~n1602 & ~n1609 ;
  assign n1611 = n798 & ~n1610 ;
  assign n1630 = n671 & ~n896 ;
  assign n1631 = ~n897 & ~n1630 ;
  assign n1632 = n308 & n1631 ;
  assign n1633 = ~n1602 & ~n1632 ;
  assign n1634 = n907 & ~n1633 ;
  assign n1601 = n333 & n671 ;
  assign n1635 = n533 & ~n912 ;
  assign n1636 = ~n1601 & ~n1635 ;
  assign n1637 = ~n1634 & n1636 ;
  assign n1638 = ~n1611 & n1637 ;
  assign n1639 = ~n1618 & n1638 ;
  assign n1640 = ~n1629 & n1639 ;
  assign n1641 = n292 & ~n1640 ;
  assign n1642 = ~n1600 & ~n1641 ;
  assign n1643 = \state_reg[0]/NET0131  & ~n1642 ;
  assign n1598 = n260 & n533 ;
  assign n1599 = \reg3_reg[15]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1644 = ~n1598 & ~n1599 ;
  assign n1645 = ~n1643 & n1644 ;
  assign n1648 = n290 & n500 ;
  assign n1650 = ~n308 & n500 ;
  assign n1651 = ~n817 & ~n827 ;
  assign n1652 = ~n1362 & n1651 ;
  assign n1653 = n1362 & ~n1651 ;
  assign n1654 = ~n1652 & ~n1653 ;
  assign n1655 = n308 & ~n1654 ;
  assign n1656 = ~n1650 & ~n1655 ;
  assign n1657 = n798 & ~n1656 ;
  assign n1673 = n622 & n891 ;
  assign n1674 = ~n602 & ~n1673 ;
  assign n1675 = n891 & n892 ;
  assign n1676 = ~n1674 & ~n1675 ;
  assign n1677 = n308 & n1676 ;
  assign n1678 = ~n1650 & ~n1677 ;
  assign n1679 = n907 & ~n1678 ;
  assign n1649 = n333 & ~n602 ;
  assign n1680 = n500 & ~n912 ;
  assign n1681 = ~n1649 & ~n1680 ;
  assign n1682 = ~n1679 & n1681 ;
  assign n1683 = ~n1657 & n1682 ;
  assign n1658 = n486 & n514 ;
  assign n1659 = n495 & ~n1658 ;
  assign n1660 = ~n516 & ~n1659 ;
  assign n1661 = ~n341 & ~n1660 ;
  assign n1662 = n341 & n513 ;
  assign n1663 = ~n1661 & ~n1662 ;
  assign n1664 = n308 & n1663 ;
  assign n1665 = ~n1650 & ~n1664 ;
  assign n1666 = n588 & ~n1665 ;
  assign n1667 = ~n1313 & n1651 ;
  assign n1668 = n1313 & ~n1651 ;
  assign n1669 = ~n1667 & ~n1668 ;
  assign n1670 = n308 & n1669 ;
  assign n1671 = ~n1650 & ~n1670 ;
  assign n1672 = n881 & ~n1671 ;
  assign n1684 = ~n1666 & ~n1672 ;
  assign n1685 = n1683 & n1684 ;
  assign n1686 = n292 & ~n1685 ;
  assign n1687 = ~n1648 & ~n1686 ;
  assign n1688 = \state_reg[0]/NET0131  & ~n1687 ;
  assign n1646 = \reg3_reg[11]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1647 = n260 & n500 ;
  assign n1689 = ~n1646 & ~n1647 ;
  assign n1690 = ~n1688 & n1689 ;
  assign n1693 = n290 & n488 ;
  assign n1696 = ~n308 & n488 ;
  assign n1697 = ~n818 & ~n826 ;
  assign n1698 = ~n1100 & n1697 ;
  assign n1699 = n1100 & ~n1697 ;
  assign n1700 = ~n1698 & ~n1699 ;
  assign n1701 = n308 & ~n1700 ;
  assign n1702 = ~n1696 & ~n1701 ;
  assign n1703 = n798 & ~n1702 ;
  assign n1718 = ~n612 & ~n1675 ;
  assign n1719 = n612 & n1675 ;
  assign n1720 = ~n1718 & ~n1719 ;
  assign n1721 = n308 & n1720 ;
  assign n1722 = ~n1696 & ~n1721 ;
  assign n1723 = n907 & ~n1722 ;
  assign n1694 = n333 & ~n612 ;
  assign n1695 = n488 & ~n912 ;
  assign n1724 = ~n1694 & ~n1695 ;
  assign n1725 = ~n1723 & n1724 ;
  assign n1726 = ~n1703 & n1725 ;
  assign n1704 = ~n1182 & n1697 ;
  assign n1705 = n1182 & ~n1697 ;
  assign n1706 = ~n1704 & ~n1705 ;
  assign n1707 = n308 & n1706 ;
  assign n1708 = ~n1696 & ~n1707 ;
  assign n1709 = n881 & ~n1708 ;
  assign n1710 = ~n516 & n526 ;
  assign n1711 = ~n1619 & ~n1710 ;
  assign n1712 = ~n341 & ~n1711 ;
  assign n1713 = n341 & n504 ;
  assign n1714 = ~n1712 & ~n1713 ;
  assign n1715 = n308 & n1714 ;
  assign n1716 = ~n1696 & ~n1715 ;
  assign n1717 = n588 & ~n1716 ;
  assign n1727 = ~n1709 & ~n1717 ;
  assign n1728 = n1726 & n1727 ;
  assign n1729 = n292 & ~n1728 ;
  assign n1730 = ~n1693 & ~n1729 ;
  assign n1731 = \state_reg[0]/NET0131  & ~n1730 ;
  assign n1691 = n260 & n488 ;
  assign n1692 = \reg3_reg[12]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1732 = ~n1691 & ~n1692 ;
  assign n1733 = ~n1731 & n1732 ;
  assign n1738 = ~n308 & n1044 ;
  assign n1739 = ~n1152 & ~n1194 ;
  assign n1740 = ~n1325 & n1739 ;
  assign n1741 = n1325 & ~n1739 ;
  assign n1742 = ~n1740 & ~n1741 ;
  assign n1743 = n308 & n1742 ;
  assign n1744 = ~n1738 & ~n1743 ;
  assign n1745 = n881 & ~n1744 ;
  assign n1746 = ~n1376 & n1739 ;
  assign n1747 = n1376 & ~n1739 ;
  assign n1748 = ~n1746 & ~n1747 ;
  assign n1749 = n308 & ~n1748 ;
  assign n1750 = ~n1738 & ~n1749 ;
  assign n1751 = n798 & ~n1750 ;
  assign n1752 = ~n1026 & n1408 ;
  assign n1753 = n1026 & ~n1408 ;
  assign n1754 = ~n1752 & ~n1753 ;
  assign n1755 = ~n341 & ~n1754 ;
  assign n1756 = n341 & n576 ;
  assign n1757 = n588 & ~n1756 ;
  assign n1758 = ~n1755 & n1757 ;
  assign n1759 = n903 & ~n1038 ;
  assign n1760 = ~n1051 & ~n1759 ;
  assign n1761 = n907 & ~n1247 ;
  assign n1762 = ~n1760 & n1761 ;
  assign n1763 = ~n1758 & ~n1762 ;
  assign n1764 = n308 & ~n1763 ;
  assign n1735 = ~n308 & n1460 ;
  assign n1736 = n912 & ~n1735 ;
  assign n1737 = n1044 & ~n1736 ;
  assign n1765 = n333 & ~n1051 ;
  assign n1766 = ~n1737 & ~n1765 ;
  assign n1767 = ~n1764 & n1766 ;
  assign n1768 = ~n1751 & n1767 ;
  assign n1769 = ~n1745 & n1768 ;
  assign n1770 = n292 & ~n1769 ;
  assign n1771 = n290 & n1044 ;
  assign n1772 = ~n1770 & ~n1771 ;
  assign n1773 = \state_reg[0]/NET0131  & ~n1772 ;
  assign n1734 = n260 & n1044 ;
  assign n1774 = \reg3_reg[19]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1775 = ~n1734 & ~n1774 ;
  assign n1776 = ~n1773 & n1775 ;
  assign n1779 = n290 & n981 ;
  assign n1780 = ~n308 & n981 ;
  assign n1781 = ~n1211 & ~n1231 ;
  assign n1782 = n1156 & n1181 ;
  assign n1783 = n1150 & ~n1163 ;
  assign n1784 = n1189 & ~n1783 ;
  assign n1785 = n1155 & ~n1784 ;
  assign n1786 = n1198 & ~n1785 ;
  assign n1787 = ~n1782 & n1786 ;
  assign n1788 = n1207 & ~n1787 ;
  assign n1789 = n1226 & ~n1788 ;
  assign n1790 = n1781 & n1789 ;
  assign n1791 = ~n1781 & ~n1789 ;
  assign n1792 = ~n1790 & ~n1791 ;
  assign n1793 = n308 & ~n1792 ;
  assign n1794 = ~n1780 & ~n1793 ;
  assign n1795 = n881 & ~n1794 ;
  assign n1819 = n1029 & n1102 ;
  assign n1820 = n1056 & n1819 ;
  assign n1821 = n1099 & n1820 ;
  assign n1814 = ~n1080 & n1102 ;
  assign n1815 = n1063 & ~n1814 ;
  assign n1816 = n1056 & ~n1815 ;
  assign n1817 = n1073 & ~n1816 ;
  assign n1818 = n1029 & ~n1817 ;
  assign n1822 = n1117 & ~n1818 ;
  assign n1823 = ~n1821 & n1822 ;
  assign n1824 = n1781 & ~n1823 ;
  assign n1825 = ~n1781 & n1823 ;
  assign n1826 = ~n1824 & ~n1825 ;
  assign n1827 = n308 & ~n1826 ;
  assign n1828 = ~n1780 & ~n1827 ;
  assign n1829 = n798 & ~n1828 ;
  assign n1804 = n341 & ~n934 ;
  assign n1806 = n579 & n1267 ;
  assign n1807 = n974 & ~n1806 ;
  assign n1805 = n579 & n1268 ;
  assign n1808 = ~n341 & ~n1805 ;
  assign n1809 = ~n1807 & n1808 ;
  assign n1810 = ~n1804 & ~n1809 ;
  assign n1811 = n308 & ~n1810 ;
  assign n1812 = ~n1780 & ~n1811 ;
  assign n1813 = n588 & ~n1812 ;
  assign n1796 = n1247 & n1250 ;
  assign n1797 = n976 & ~n1796 ;
  assign n1798 = ~n1252 & ~n1797 ;
  assign n1799 = n308 & n1798 ;
  assign n1800 = ~n1780 & ~n1799 ;
  assign n1801 = n907 & ~n1800 ;
  assign n1802 = n333 & n976 ;
  assign n1803 = ~n912 & n981 ;
  assign n1830 = ~n1802 & ~n1803 ;
  assign n1831 = ~n1801 & n1830 ;
  assign n1832 = ~n1813 & n1831 ;
  assign n1833 = ~n1829 & n1832 ;
  assign n1834 = ~n1795 & n1833 ;
  assign n1835 = n292 & ~n1834 ;
  assign n1836 = ~n1779 & ~n1835 ;
  assign n1837 = \state_reg[0]/NET0131  & ~n1836 ;
  assign n1777 = n260 & n981 ;
  assign n1778 = \reg3_reg[24]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1838 = ~n1777 & ~n1778 ;
  assign n1839 = ~n1837 & n1838 ;
  assign n1842 = n290 & n930 ;
  assign n1843 = ~n308 & n930 ;
  assign n1844 = ~n1204 & ~n1222 ;
  assign n1856 = n1306 & n1328 ;
  assign n1857 = ~n1612 & n1856 ;
  assign n1858 = ~n1323 & n1328 ;
  assign n1859 = n1339 & ~n1858 ;
  assign n1860 = ~n1857 & n1859 ;
  assign n1861 = n1844 & n1860 ;
  assign n1862 = ~n1844 & ~n1860 ;
  assign n1863 = ~n1861 & ~n1862 ;
  assign n1864 = n308 & ~n1863 ;
  assign n1865 = ~n1843 & ~n1864 ;
  assign n1866 = n881 & ~n1865 ;
  assign n1845 = n1364 & n1379 ;
  assign n1846 = ~n1605 & n1845 ;
  assign n1847 = ~n1374 & n1379 ;
  assign n1848 = n1392 & ~n1847 ;
  assign n1849 = ~n1846 & n1848 ;
  assign n1850 = n1844 & ~n1849 ;
  assign n1851 = ~n1844 & n1849 ;
  assign n1852 = ~n1850 & ~n1851 ;
  assign n1853 = n308 & ~n1852 ;
  assign n1854 = ~n1843 & ~n1853 ;
  assign n1855 = n798 & ~n1854 ;
  assign n1868 = ~n985 & n1409 ;
  assign n1869 = n985 & ~n1409 ;
  assign n1870 = ~n1868 & ~n1869 ;
  assign n1871 = ~n341 & ~n1870 ;
  assign n1872 = n341 & n1001 ;
  assign n1873 = ~n1871 & ~n1872 ;
  assign n1874 = n308 & n1873 ;
  assign n1875 = ~n1843 & ~n1874 ;
  assign n1876 = n588 & ~n1875 ;
  assign n1877 = n1247 & n1249 ;
  assign n1878 = n989 & ~n1877 ;
  assign n1879 = ~n1796 & ~n1878 ;
  assign n1880 = n308 & n1879 ;
  assign n1881 = ~n1843 & ~n1880 ;
  assign n1882 = n907 & ~n1881 ;
  assign n1867 = n333 & n989 ;
  assign n1883 = ~n912 & n930 ;
  assign n1884 = ~n1867 & ~n1883 ;
  assign n1885 = ~n1882 & n1884 ;
  assign n1886 = ~n1876 & n1885 ;
  assign n1887 = ~n1855 & n1886 ;
  assign n1888 = ~n1866 & n1887 ;
  assign n1889 = n292 & ~n1888 ;
  assign n1890 = ~n1842 & ~n1889 ;
  assign n1891 = \state_reg[0]/NET0131  & ~n1890 ;
  assign n1840 = \reg3_reg[23]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1841 = n260 & n930 ;
  assign n1892 = ~n1840 & ~n1841 ;
  assign n1893 = ~n1891 & n1892 ;
  assign n1894 = \reg0_reg[15]/NET0131  & ~n1471 ;
  assign n1895 = \reg0_reg[15]/NET0131  & n290 ;
  assign n1900 = \reg0_reg[15]/NET0131  & ~n1444 ;
  assign n1907 = n1444 & n1626 ;
  assign n1908 = ~n1900 & ~n1907 ;
  assign n1909 = n588 & ~n1908 ;
  assign n1904 = n1444 & ~n1615 ;
  assign n1905 = ~n1900 & ~n1904 ;
  assign n1906 = n881 & ~n1905 ;
  assign n1901 = n1444 & n1608 ;
  assign n1902 = ~n1900 & ~n1901 ;
  assign n1903 = n798 & ~n1902 ;
  assign n1896 = n671 & n910 ;
  assign n1897 = n907 & n1631 ;
  assign n1898 = ~n1896 & ~n1897 ;
  assign n1899 = n1444 & ~n1898 ;
  assign n1910 = n907 & ~n1444 ;
  assign n1911 = n1459 & ~n1910 ;
  assign n1912 = \reg0_reg[15]/NET0131  & ~n1911 ;
  assign n1913 = ~n1899 & ~n1912 ;
  assign n1914 = ~n1903 & n1913 ;
  assign n1915 = ~n1906 & n1914 ;
  assign n1916 = ~n1909 & n1915 ;
  assign n1917 = n292 & ~n1916 ;
  assign n1918 = ~n1895 & ~n1917 ;
  assign n1919 = \state_reg[0]/NET0131  & ~n1918 ;
  assign n1920 = ~n1894 & ~n1919 ;
  assign n1921 = \reg0_reg[23]/NET0131  & ~n1471 ;
  assign n1922 = \reg0_reg[23]/NET0131  & n290 ;
  assign n1923 = \reg0_reg[23]/NET0131  & ~n1444 ;
  assign n1927 = n1444 & ~n1863 ;
  assign n1928 = ~n1923 & ~n1927 ;
  assign n1929 = n881 & ~n1928 ;
  assign n1924 = n1444 & ~n1852 ;
  assign n1925 = ~n1923 & ~n1924 ;
  assign n1926 = n798 & ~n1925 ;
  assign n1934 = n1444 & n1873 ;
  assign n1935 = ~n1923 & ~n1934 ;
  assign n1936 = n588 & ~n1935 ;
  assign n1930 = n910 & n989 ;
  assign n1931 = n907 & n1879 ;
  assign n1932 = ~n1930 & ~n1931 ;
  assign n1933 = n1444 & ~n1932 ;
  assign n1937 = \reg0_reg[23]/NET0131  & ~n1911 ;
  assign n1938 = ~n1933 & ~n1937 ;
  assign n1939 = ~n1936 & n1938 ;
  assign n1940 = ~n1926 & n1939 ;
  assign n1941 = ~n1929 & n1940 ;
  assign n1942 = n292 & ~n1941 ;
  assign n1943 = ~n1922 & ~n1942 ;
  assign n1944 = \state_reg[0]/NET0131  & ~n1943 ;
  assign n1945 = ~n1921 & ~n1944 ;
  assign n1946 = \reg0_reg[24]/NET0131  & ~n1471 ;
  assign n1947 = \reg0_reg[24]/NET0131  & n290 ;
  assign n1951 = n798 & ~n1826 ;
  assign n1950 = n588 & ~n1810 ;
  assign n1948 = n907 & n1798 ;
  assign n1949 = n910 & n976 ;
  assign n1952 = ~n1948 & ~n1949 ;
  assign n1953 = ~n1950 & n1952 ;
  assign n1954 = ~n1951 & n1953 ;
  assign n1955 = n1444 & ~n1954 ;
  assign n1956 = ~n588 & ~n798 ;
  assign n1957 = ~n1444 & ~n1956 ;
  assign n1958 = n1911 & ~n1957 ;
  assign n1959 = \reg0_reg[24]/NET0131  & ~n1958 ;
  assign n1961 = n1444 & n1792 ;
  assign n1960 = ~\reg0_reg[24]/NET0131  & ~n1444 ;
  assign n1962 = n881 & ~n1960 ;
  assign n1963 = ~n1961 & n1962 ;
  assign n1964 = ~n1959 & ~n1963 ;
  assign n1965 = ~n1955 & n1964 ;
  assign n1966 = n292 & ~n1965 ;
  assign n1967 = ~n1947 & ~n1966 ;
  assign n1968 = \state_reg[0]/NET0131  & ~n1967 ;
  assign n1969 = ~n1946 & ~n1968 ;
  assign n1970 = \reg1_reg[15]/NET0131  & ~n1471 ;
  assign n1971 = \reg1_reg[15]/NET0131  & n290 ;
  assign n1973 = \reg1_reg[15]/NET0131  & ~n1497 ;
  assign n1980 = n1497 & n1626 ;
  assign n1981 = ~n1973 & ~n1980 ;
  assign n1982 = n588 & ~n1981 ;
  assign n1977 = n1497 & ~n1615 ;
  assign n1978 = ~n1973 & ~n1977 ;
  assign n1979 = n881 & ~n1978 ;
  assign n1974 = n1497 & n1608 ;
  assign n1975 = ~n1973 & ~n1974 ;
  assign n1976 = n798 & ~n1975 ;
  assign n1972 = n1497 & ~n1898 ;
  assign n1983 = \reg1_reg[15]/NET0131  & ~n1507 ;
  assign n1984 = ~n1972 & ~n1983 ;
  assign n1985 = ~n1976 & n1984 ;
  assign n1986 = ~n1979 & n1985 ;
  assign n1987 = ~n1982 & n1986 ;
  assign n1988 = n292 & ~n1987 ;
  assign n1989 = ~n1971 & ~n1988 ;
  assign n1990 = \state_reg[0]/NET0131  & ~n1989 ;
  assign n1991 = ~n1970 & ~n1990 ;
  assign n1992 = \reg1_reg[23]/NET0131  & ~n1471 ;
  assign n1993 = \reg1_reg[23]/NET0131  & n290 ;
  assign n1994 = \reg1_reg[23]/NET0131  & ~n1497 ;
  assign n1998 = n1497 & ~n1863 ;
  assign n1999 = ~n1994 & ~n1998 ;
  assign n2000 = n881 & ~n1999 ;
  assign n1995 = n1497 & ~n1852 ;
  assign n1996 = ~n1994 & ~n1995 ;
  assign n1997 = n798 & ~n1996 ;
  assign n2002 = n1497 & n1873 ;
  assign n2003 = ~n1994 & ~n2002 ;
  assign n2004 = n588 & ~n2003 ;
  assign n2001 = n1497 & ~n1932 ;
  assign n2005 = \reg1_reg[23]/NET0131  & ~n1507 ;
  assign n2006 = ~n2001 & ~n2005 ;
  assign n2007 = ~n2004 & n2006 ;
  assign n2008 = ~n1997 & n2007 ;
  assign n2009 = ~n2000 & n2008 ;
  assign n2010 = n292 & ~n2009 ;
  assign n2011 = ~n1993 & ~n2010 ;
  assign n2012 = \state_reg[0]/NET0131  & ~n2011 ;
  assign n2013 = ~n1992 & ~n2012 ;
  assign n2014 = \reg1_reg[24]/NET0131  & ~n1471 ;
  assign n2015 = \reg1_reg[24]/NET0131  & n290 ;
  assign n2016 = n1497 & ~n1954 ;
  assign n2017 = n798 & ~n1497 ;
  assign n2018 = n1507 & ~n2017 ;
  assign n2019 = ~n1508 & n2018 ;
  assign n2020 = \reg1_reg[24]/NET0131  & ~n2019 ;
  assign n2022 = n1497 & n1792 ;
  assign n2021 = ~\reg1_reg[24]/NET0131  & ~n1497 ;
  assign n2023 = n881 & ~n2021 ;
  assign n2024 = ~n2022 & n2023 ;
  assign n2025 = ~n2020 & ~n2024 ;
  assign n2026 = ~n2016 & n2025 ;
  assign n2027 = n292 & ~n2026 ;
  assign n2028 = ~n2015 & ~n2027 ;
  assign n2029 = \state_reg[0]/NET0131  & ~n2028 ;
  assign n2030 = ~n2014 & ~n2029 ;
  assign n2031 = \reg2_reg[15]/NET0131  & ~n1471 ;
  assign n2032 = \reg2_reg[15]/NET0131  & n290 ;
  assign n2034 = \reg2_reg[15]/NET0131  & ~n1543 ;
  assign n2035 = n1543 & n1626 ;
  assign n2036 = ~n2034 & ~n2035 ;
  assign n2037 = n588 & ~n2036 ;
  assign n2041 = n1543 & ~n1615 ;
  assign n2042 = ~n2034 & ~n2041 ;
  assign n2043 = n881 & ~n2042 ;
  assign n2038 = n1543 & n1608 ;
  assign n2039 = ~n2034 & ~n2038 ;
  assign n2040 = n798 & ~n2039 ;
  assign n2033 = n1543 & ~n1898 ;
  assign n2044 = n329 & n533 ;
  assign n2045 = n1422 & ~n1543 ;
  assign n2046 = ~n909 & ~n2045 ;
  assign n2047 = \reg2_reg[15]/NET0131  & ~n2046 ;
  assign n2048 = ~n2044 & ~n2047 ;
  assign n2049 = ~n2033 & n2048 ;
  assign n2050 = ~n2040 & n2049 ;
  assign n2051 = ~n2043 & n2050 ;
  assign n2052 = ~n2037 & n2051 ;
  assign n2053 = n292 & ~n2052 ;
  assign n2054 = ~n2032 & ~n2053 ;
  assign n2055 = \state_reg[0]/NET0131  & ~n2054 ;
  assign n2056 = ~n2031 & ~n2055 ;
  assign n2057 = \reg2_reg[23]/NET0131  & ~n1471 ;
  assign n2058 = \reg2_reg[23]/NET0131  & n290 ;
  assign n2059 = \reg2_reg[23]/NET0131  & ~n1543 ;
  assign n2063 = n1543 & ~n1863 ;
  assign n2064 = ~n2059 & ~n2063 ;
  assign n2065 = n881 & ~n2064 ;
  assign n2060 = n1543 & ~n1852 ;
  assign n2061 = ~n2059 & ~n2060 ;
  assign n2062 = n798 & ~n2061 ;
  assign n2067 = n1543 & n1873 ;
  assign n2068 = ~n2059 & ~n2067 ;
  assign n2069 = n588 & ~n2068 ;
  assign n2070 = n1543 & ~n1932 ;
  assign n2066 = n329 & n930 ;
  assign n2071 = \reg2_reg[23]/NET0131  & ~n2046 ;
  assign n2072 = ~n2066 & ~n2071 ;
  assign n2073 = ~n2070 & n2072 ;
  assign n2074 = ~n2069 & n2073 ;
  assign n2075 = ~n2062 & n2074 ;
  assign n2076 = ~n2065 & n2075 ;
  assign n2077 = n292 & ~n2076 ;
  assign n2078 = ~n2058 & ~n2077 ;
  assign n2079 = \state_reg[0]/NET0131  & ~n2078 ;
  assign n2080 = ~n2057 & ~n2079 ;
  assign n2081 = \reg2_reg[29]/NET0131  & n290 ;
  assign n2082 = \reg2_reg[29]/NET0131  & ~n1543 ;
  assign n2083 = n341 & ~n1138 ;
  assign n2086 = ~n1279 & n1414 ;
  assign n2089 = \reg0_reg[30]/NET0131  & n376 ;
  assign n2087 = \reg1_reg[30]/NET0131  & n374 ;
  assign n2088 = \reg2_reg[30]/NET0131  & n372 ;
  assign n2090 = ~n2087 & ~n2088 ;
  assign n2091 = ~n2089 & n2090 ;
  assign n2092 = ~n409 & n2091 ;
  assign n2094 = n2086 & ~n2092 ;
  assign n2084 = ~\B_reg/NET0131  & ~n341 ;
  assign n2085 = ~n348 & ~n2084 ;
  assign n2093 = ~n2086 & n2092 ;
  assign n2095 = ~n2085 & ~n2093 ;
  assign n2096 = ~n2094 & n2095 ;
  assign n2097 = ~n2083 & ~n2096 ;
  assign n2098 = n1543 & ~n2097 ;
  assign n2099 = ~n2082 & ~n2098 ;
  assign n2100 = n588 & ~n2099 ;
  assign n2101 = \datai[29]_pad  & ~n348 ;
  assign n2102 = n1279 & n2101 ;
  assign n2103 = ~n1279 & ~n2101 ;
  assign n2104 = ~n2102 & ~n2103 ;
  assign n2137 = n689 & n785 ;
  assign n2138 = n689 & ~n732 ;
  assign n2139 = n639 & ~n2138 ;
  assign n2140 = ~n2137 & n2139 ;
  assign n2141 = n1363 & n1377 ;
  assign n2142 = n674 & n2141 ;
  assign n2143 = ~n2140 & n2142 ;
  assign n2144 = ~n685 & n2141 ;
  assign n2145 = n1373 & n1377 ;
  assign n2146 = ~n1388 & ~n2145 ;
  assign n2147 = ~n2144 & n2146 ;
  assign n2148 = ~n2143 & n2147 ;
  assign n2149 = n1378 & n1380 ;
  assign n2150 = n1131 & n1138 ;
  assign n2151 = ~n952 & ~n2150 ;
  assign n2152 = n1381 & n2151 ;
  assign n2153 = n2149 & n2152 ;
  assign n2154 = ~n2148 & n2153 ;
  assign n2156 = n1380 & n1391 ;
  assign n2157 = n1395 & ~n2156 ;
  assign n2158 = n2152 & ~n2157 ;
  assign n2160 = n1386 & n2151 ;
  assign n2155 = n1120 & ~n2150 ;
  assign n2159 = ~n1131 & ~n1138 ;
  assign n2161 = ~n2155 & ~n2159 ;
  assign n2162 = ~n2160 & n2161 ;
  assign n2163 = ~n2158 & n2162 ;
  assign n2164 = ~n2154 & n2163 ;
  assign n2165 = ~n2104 & n2164 ;
  assign n2166 = n2104 & ~n2164 ;
  assign n2167 = ~n2165 & ~n2166 ;
  assign n2168 = n1543 & n2167 ;
  assign n2169 = ~n2082 & ~n2168 ;
  assign n2170 = n798 & ~n2169 ;
  assign n2105 = n835 & n871 ;
  assign n2106 = n835 & ~n849 ;
  assign n2107 = n830 & ~n2106 ;
  assign n2108 = ~n2105 & n2107 ;
  assign n2109 = n1305 & n1327 ;
  assign n2110 = n816 & n2109 ;
  assign n2111 = ~n2108 & n2110 ;
  assign n2112 = ~n813 & n2109 ;
  assign n2113 = ~n1322 & n1327 ;
  assign n2114 = n1335 & ~n2113 ;
  assign n2115 = ~n2112 & n2114 ;
  assign n2116 = ~n2111 & n2115 ;
  assign n2117 = n1326 & n1329 ;
  assign n2118 = ~n1139 & ~n1212 ;
  assign n2119 = n1210 & n2118 ;
  assign n2120 = n2117 & n2119 ;
  assign n2121 = ~n2116 & n2120 ;
  assign n2125 = n1210 & ~n1341 ;
  assign n2126 = ~n1228 & ~n2125 ;
  assign n2127 = ~n1139 & ~n2126 ;
  assign n2122 = n1329 & ~n1338 ;
  assign n2123 = n1343 & ~n2122 ;
  assign n2124 = n2119 & ~n2123 ;
  assign n2128 = ~n1140 & ~n2124 ;
  assign n2129 = ~n2127 & n2128 ;
  assign n2130 = ~n2121 & n2129 ;
  assign n2131 = ~n2104 & n2130 ;
  assign n2132 = n2104 & ~n2130 ;
  assign n2133 = ~n2131 & ~n2132 ;
  assign n2134 = n1543 & ~n2133 ;
  assign n2135 = ~n2082 & ~n2134 ;
  assign n2136 = n881 & ~n2135 ;
  assign n2171 = n1258 & ~n2101 ;
  assign n2172 = ~n1258 & n2101 ;
  assign n2173 = ~n2171 & ~n2172 ;
  assign n2174 = n1543 & n2173 ;
  assign n2175 = ~n2082 & ~n2174 ;
  assign n2176 = n907 & ~n2175 ;
  assign n2180 = \reg2_reg[29]/NET0131  & ~n1560 ;
  assign n2177 = n329 & n408 ;
  assign n2178 = n910 & n2101 ;
  assign n2179 = n1543 & n2178 ;
  assign n2181 = ~n2177 & ~n2179 ;
  assign n2182 = ~n2180 & n2181 ;
  assign n2183 = ~n2176 & n2182 ;
  assign n2184 = ~n2136 & n2183 ;
  assign n2185 = ~n2170 & n2184 ;
  assign n2186 = ~n2100 & n2185 ;
  assign n2187 = n292 & ~n2186 ;
  assign n2188 = ~n2081 & ~n2187 ;
  assign n2189 = \state_reg[0]/NET0131  & ~n2188 ;
  assign n2190 = \reg2_reg[29]/NET0131  & ~n1471 ;
  assign n2191 = ~n2189 & ~n2190 ;
  assign n2194 = n290 & n542 ;
  assign n2196 = ~n308 & n542 ;
  assign n2197 = n537 & ~n1620 ;
  assign n2198 = ~n1621 & ~n2197 ;
  assign n2199 = ~n341 & ~n2198 ;
  assign n2200 = n341 & n526 ;
  assign n2201 = ~n2199 & ~n2200 ;
  assign n2202 = n308 & n2201 ;
  assign n2203 = ~n2196 & ~n2202 ;
  assign n2204 = n588 & ~n2203 ;
  assign n2216 = ~n647 & ~n676 ;
  assign n2223 = ~n1170 & n1173 ;
  assign n2224 = n1164 & n1179 ;
  assign n2225 = ~n2223 & n2224 ;
  assign n2226 = ~n1176 & n1179 ;
  assign n2227 = ~n1159 & ~n2226 ;
  assign n2228 = ~n2225 & n2227 ;
  assign n2229 = n1148 & n1157 ;
  assign n2230 = ~n2228 & n2229 ;
  assign n2231 = n1148 & ~n1162 ;
  assign n2232 = n1185 & ~n2231 ;
  assign n2233 = ~n2230 & n2232 ;
  assign n2234 = n2216 & n2233 ;
  assign n2235 = ~n2216 & ~n2233 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = n308 & n2236 ;
  assign n2238 = ~n2196 & ~n2237 ;
  assign n2239 = n881 & ~n2238 ;
  assign n2205 = ~n1079 & n1101 ;
  assign n2206 = n1059 & ~n2205 ;
  assign n2207 = n1074 & n1101 ;
  assign n2208 = ~n1094 & n1097 ;
  assign n2209 = ~n1076 & ~n2208 ;
  assign n2210 = n1081 & n1097 ;
  assign n2211 = ~n1088 & ~n1091 ;
  assign n2212 = n2210 & ~n2211 ;
  assign n2213 = n2209 & ~n2212 ;
  assign n2214 = n2207 & ~n2213 ;
  assign n2215 = n2206 & ~n2214 ;
  assign n2217 = n2215 & n2216 ;
  assign n2218 = ~n2215 & ~n2216 ;
  assign n2219 = ~n2217 & ~n2218 ;
  assign n2220 = n308 & ~n2219 ;
  assign n2221 = ~n2196 & ~n2220 ;
  assign n2222 = n798 & ~n2221 ;
  assign n2240 = ~n646 & ~n895 ;
  assign n2241 = ~n896 & ~n2240 ;
  assign n2242 = n308 & n2241 ;
  assign n2243 = ~n2196 & ~n2242 ;
  assign n2244 = n907 & ~n2243 ;
  assign n2195 = n333 & ~n646 ;
  assign n2245 = n542 & ~n912 ;
  assign n2246 = ~n2195 & ~n2245 ;
  assign n2247 = ~n2244 & n2246 ;
  assign n2248 = ~n2222 & n2247 ;
  assign n2249 = ~n2239 & n2248 ;
  assign n2250 = ~n2204 & n2249 ;
  assign n2251 = n292 & ~n2250 ;
  assign n2252 = ~n2194 & ~n2251 ;
  assign n2253 = \state_reg[0]/NET0131  & ~n2252 ;
  assign n2192 = \reg3_reg[14]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2193 = n260 & n542 ;
  assign n2254 = ~n2192 & ~n2193 ;
  assign n2255 = ~n2253 & n2254 ;
  assign n2258 = n290 & n551 ;
  assign n2260 = ~n308 & n551 ;
  assign n2261 = ~n663 & ~n681 ;
  assign n2269 = n1150 & ~n1182 ;
  assign n2270 = n1189 & ~n2269 ;
  assign n2271 = n2261 & n2270 ;
  assign n2272 = ~n2261 & ~n2270 ;
  assign n2273 = ~n2271 & ~n2272 ;
  assign n2274 = n308 & n2273 ;
  assign n2275 = ~n2260 & ~n2274 ;
  assign n2276 = n881 & ~n2275 ;
  assign n2262 = n1063 & ~n1103 ;
  assign n2263 = n2261 & n2262 ;
  assign n2264 = ~n2261 & ~n2262 ;
  assign n2265 = ~n2263 & ~n2264 ;
  assign n2266 = n308 & ~n2265 ;
  assign n2267 = ~n2260 & ~n2266 ;
  assign n2268 = n798 & ~n2267 ;
  assign n2277 = ~n559 & n566 ;
  assign n2278 = ~n567 & ~n2277 ;
  assign n2279 = ~n341 & ~n2278 ;
  assign n2280 = n341 & n537 ;
  assign n2281 = ~n2279 & ~n2280 ;
  assign n2282 = n308 & n2281 ;
  assign n2283 = ~n2260 & ~n2282 ;
  assign n2284 = n588 & ~n2283 ;
  assign n2285 = ~n662 & ~n897 ;
  assign n2286 = ~n898 & ~n2285 ;
  assign n2287 = n308 & n2286 ;
  assign n2288 = ~n2260 & ~n2287 ;
  assign n2289 = n907 & ~n2288 ;
  assign n2259 = n333 & ~n662 ;
  assign n2290 = n551 & ~n912 ;
  assign n2291 = ~n2259 & ~n2290 ;
  assign n2292 = ~n2289 & n2291 ;
  assign n2293 = ~n2284 & n2292 ;
  assign n2294 = ~n2268 & n2293 ;
  assign n2295 = ~n2276 & n2294 ;
  assign n2296 = n292 & ~n2295 ;
  assign n2297 = ~n2258 & ~n2296 ;
  assign n2298 = \state_reg[0]/NET0131  & ~n2297 ;
  assign n2256 = \reg3_reg[16]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2257 = n260 & n551 ;
  assign n2299 = ~n2256 & ~n2257 ;
  assign n2300 = ~n2298 & n2299 ;
  assign n2303 = n290 & n479 ;
  assign n2308 = ~n308 & n479 ;
  assign n2309 = n456 & ~n483 ;
  assign n2310 = n465 & ~n2309 ;
  assign n2311 = ~n465 & n2309 ;
  assign n2312 = ~n2310 & ~n2311 ;
  assign n2313 = ~n341 & ~n2312 ;
  assign n2314 = n341 & n445 ;
  assign n2315 = ~n2313 & ~n2314 ;
  assign n2316 = n308 & n2315 ;
  assign n2317 = ~n2308 & ~n2316 ;
  assign n2318 = n588 & ~n2317 ;
  assign n2319 = ~n837 & ~n846 ;
  assign n2326 = ~n1357 & n2319 ;
  assign n2327 = n1357 & ~n2319 ;
  assign n2328 = ~n2326 & ~n2327 ;
  assign n2329 = n308 & ~n2328 ;
  assign n2330 = ~n2308 & ~n2329 ;
  assign n2331 = n798 & ~n2330 ;
  assign n2320 = ~n1308 & n2319 ;
  assign n2321 = n1308 & ~n2319 ;
  assign n2322 = ~n2320 & ~n2321 ;
  assign n2323 = n308 & n2322 ;
  assign n2324 = ~n2308 & ~n2323 ;
  assign n2325 = n881 & ~n2324 ;
  assign n2304 = ~n698 & ~n888 ;
  assign n2305 = ~n889 & n907 ;
  assign n2306 = ~n2304 & n2305 ;
  assign n2307 = n308 & n2306 ;
  assign n2332 = n479 & ~n1424 ;
  assign n2333 = n333 & ~n698 ;
  assign n2334 = ~n2332 & ~n2333 ;
  assign n2335 = ~n2307 & n2334 ;
  assign n2336 = ~n2325 & n2335 ;
  assign n2337 = ~n2331 & n2336 ;
  assign n2338 = ~n2318 & n2337 ;
  assign n2339 = n292 & ~n2338 ;
  assign n2340 = ~n2303 & ~n2339 ;
  assign n2341 = \state_reg[0]/NET0131  & ~n2340 ;
  assign n2301 = \reg3_reg[7]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2302 = n260 & n479 ;
  assign n2342 = ~n2301 & ~n2302 ;
  assign n2343 = ~n2341 & n2342 ;
  assign n2346 = n290 & n1022 ;
  assign n2348 = ~n308 & n1022 ;
  assign n2349 = ~n1202 & ~n1218 ;
  assign n2350 = ~n1106 & n2349 ;
  assign n2351 = n1106 & ~n2349 ;
  assign n2352 = ~n2350 & ~n2351 ;
  assign n2353 = n308 & ~n2352 ;
  assign n2354 = ~n2348 & ~n2353 ;
  assign n2355 = n798 & ~n2354 ;
  assign n2362 = ~n1014 & n1752 ;
  assign n2363 = n1014 & ~n1752 ;
  assign n2364 = ~n2362 & ~n2363 ;
  assign n2365 = ~n341 & ~n2364 ;
  assign n2366 = n341 & n1048 ;
  assign n2367 = ~n2365 & ~n2366 ;
  assign n2368 = n308 & n2367 ;
  assign n2369 = ~n2348 & ~n2368 ;
  assign n2370 = n588 & ~n2369 ;
  assign n2356 = n1200 & n2349 ;
  assign n2357 = ~n1200 & ~n2349 ;
  assign n2358 = ~n2356 & ~n2357 ;
  assign n2359 = n308 & ~n2358 ;
  assign n2360 = ~n2348 & ~n2359 ;
  assign n2361 = n881 & ~n2360 ;
  assign n2371 = ~n1016 & n1247 ;
  assign n2372 = n1016 & ~n1247 ;
  assign n2373 = ~n2371 & ~n2372 ;
  assign n2374 = n308 & n2373 ;
  assign n2375 = ~n2348 & ~n2374 ;
  assign n2376 = n907 & ~n2375 ;
  assign n2347 = n333 & n1016 ;
  assign n2377 = ~n912 & n1022 ;
  assign n2378 = ~n2347 & ~n2377 ;
  assign n2379 = ~n2376 & n2378 ;
  assign n2380 = ~n2361 & n2379 ;
  assign n2381 = ~n2370 & n2380 ;
  assign n2382 = ~n2355 & n2381 ;
  assign n2383 = n292 & ~n2382 ;
  assign n2384 = ~n2346 & ~n2383 ;
  assign n2385 = \state_reg[0]/NET0131  & ~n2384 ;
  assign n2344 = n260 & n1022 ;
  assign n2345 = \reg3_reg[20]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2386 = ~n2344 & ~n2345 ;
  assign n2387 = ~n2385 & n2386 ;
  assign n2388 = ~n329 & ~n1543 ;
  assign n2389 = \state_reg[0]/NET0131  & n292 ;
  assign n2390 = ~n909 & n2389 ;
  assign n2391 = ~n2388 & n2390 ;
  assign n2392 = \reg2_reg[31]/NET0131  & ~n2391 ;
  assign n2393 = \datai[31]_pad  & ~n348 ;
  assign n2403 = \datai[30]_pad  & ~n348 ;
  assign n2404 = n2171 & ~n2403 ;
  assign n2406 = ~n2393 & n2404 ;
  assign n2405 = n2393 & ~n2404 ;
  assign n2407 = n907 & ~n2405 ;
  assign n2408 = ~n2406 & n2407 ;
  assign n2394 = n910 & n2393 ;
  assign n2395 = ~n962 & n1805 ;
  assign n2396 = ~n951 & n2395 ;
  assign n2397 = ~n1279 & ~n2092 ;
  assign n2398 = ~n1138 & n2397 ;
  assign n2399 = n2396 & n2398 ;
  assign n2400 = n588 & ~n2085 ;
  assign n2401 = ~n415 & n2400 ;
  assign n2402 = ~n2399 & n2401 ;
  assign n2409 = ~n2394 & ~n2402 ;
  assign n2410 = ~n2408 & n2409 ;
  assign n2411 = n1543 & ~n2410 ;
  assign n2412 = ~n2177 & ~n2411 ;
  assign n2413 = n2389 & ~n2412 ;
  assign n2414 = ~n2392 & ~n2413 ;
  assign n2415 = ~n308 & n958 ;
  assign n2416 = ~n1209 & ~n1229 ;
  assign n2417 = n1151 & ~n1188 ;
  assign n2418 = n1192 & ~n2417 ;
  assign n2419 = n1149 & n1151 ;
  assign n2420 = ~n2233 & n2419 ;
  assign n2421 = n2418 & ~n2420 ;
  assign n2422 = n1206 & n1213 ;
  assign n2423 = n1154 & n1203 ;
  assign n2424 = n2422 & n2423 ;
  assign n2425 = ~n2421 & n2424 ;
  assign n2427 = ~n1197 & n1203 ;
  assign n2428 = n1220 & ~n2427 ;
  assign n2429 = n2422 & ~n2428 ;
  assign n2426 = n1213 & ~n1225 ;
  assign n2430 = n1233 & ~n2426 ;
  assign n2431 = ~n2429 & n2430 ;
  assign n2432 = ~n2425 & n2431 ;
  assign n2433 = n2416 & n2432 ;
  assign n2434 = ~n2416 & ~n2432 ;
  assign n2435 = ~n2433 & ~n2434 ;
  assign n2436 = n308 & ~n2435 ;
  assign n2437 = ~n2415 & ~n2436 ;
  assign n2438 = n881 & ~n2437 ;
  assign n2439 = n951 & ~n2395 ;
  assign n2440 = ~n2396 & ~n2439 ;
  assign n2441 = ~n341 & ~n2440 ;
  assign n2442 = n341 & n974 ;
  assign n2443 = ~n2441 & ~n2442 ;
  assign n2444 = n308 & n2443 ;
  assign n2445 = ~n2415 & ~n2444 ;
  assign n2446 = n588 & ~n2445 ;
  assign n2450 = ~n965 & n1252 ;
  assign n2451 = n953 & ~n2450 ;
  assign n2452 = ~n1253 & ~n2451 ;
  assign n2453 = n308 & n2452 ;
  assign n2454 = ~n2415 & ~n2453 ;
  assign n2455 = n907 & ~n2454 ;
  assign n2462 = n1085 & n1087 ;
  assign n2463 = ~n1091 & ~n2462 ;
  assign n2464 = n2210 & ~n2463 ;
  assign n2465 = n1087 & n2210 ;
  assign n2466 = n1083 & n2465 ;
  assign n2467 = n2209 & ~n2466 ;
  assign n2468 = ~n2464 & n2467 ;
  assign n2458 = n1055 & n1057 ;
  assign n2469 = n2207 & n2458 ;
  assign n2470 = ~n2468 & n2469 ;
  assign n2459 = ~n2206 & n2458 ;
  assign n2460 = n1055 & n1062 ;
  assign n2461 = ~n1067 & ~n2460 ;
  assign n2471 = ~n2459 & n2461 ;
  assign n2472 = ~n2470 & n2471 ;
  assign n2456 = n987 & n1003 ;
  assign n2457 = n1028 & n1053 ;
  assign n2473 = n2456 & n2457 ;
  assign n2474 = ~n2472 & n2473 ;
  assign n2476 = n1028 & n1072 ;
  assign n2477 = ~n1111 & ~n2476 ;
  assign n2478 = n2456 & ~n2477 ;
  assign n2475 = n987 & ~n1116 ;
  assign n2479 = ~n1125 & ~n2475 ;
  assign n2480 = ~n2478 & n2479 ;
  assign n2481 = ~n2474 & n2480 ;
  assign n2482 = n2416 & ~n2481 ;
  assign n2483 = ~n2416 & n2481 ;
  assign n2484 = ~n2482 & ~n2483 ;
  assign n2485 = n798 & ~n2484 ;
  assign n2486 = n308 & n2485 ;
  assign n2447 = ~n308 & n798 ;
  assign n2448 = n912 & ~n2447 ;
  assign n2449 = n958 & ~n2448 ;
  assign n2487 = n333 & n953 ;
  assign n2488 = ~n2449 & ~n2487 ;
  assign n2489 = ~n2486 & n2488 ;
  assign n2490 = ~n2455 & n2489 ;
  assign n2491 = ~n2446 & n2490 ;
  assign n2492 = ~n2438 & n2491 ;
  assign n2493 = n292 & ~n2492 ;
  assign n2494 = n290 & n958 ;
  assign n2495 = ~n2493 & ~n2494 ;
  assign n2496 = \state_reg[0]/NET0131  & ~n2495 ;
  assign n2497 = \reg3_reg[26]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2498 = n260 & n958 ;
  assign n2499 = ~n2497 & ~n2498 ;
  assign n2500 = ~n2496 & n2499 ;
  assign n2501 = \reg0_reg[19]/NET0131  & ~n1471 ;
  assign n2502 = \reg0_reg[19]/NET0131  & n290 ;
  assign n2506 = \reg0_reg[19]/NET0131  & ~n1444 ;
  assign n2507 = n1444 & n1742 ;
  assign n2508 = ~n2506 & ~n2507 ;
  assign n2509 = n881 & ~n2508 ;
  assign n2510 = n1444 & ~n1748 ;
  assign n2511 = ~n2506 & ~n2510 ;
  assign n2512 = n798 & ~n2511 ;
  assign n2503 = n910 & ~n1051 ;
  assign n2504 = n1763 & ~n2503 ;
  assign n2505 = n1444 & ~n2504 ;
  assign n2513 = \reg0_reg[19]/NET0131  & ~n1462 ;
  assign n2514 = ~n2505 & ~n2513 ;
  assign n2515 = ~n2512 & n2514 ;
  assign n2516 = ~n2509 & n2515 ;
  assign n2517 = n292 & ~n2516 ;
  assign n2518 = ~n2502 & ~n2517 ;
  assign n2519 = \state_reg[0]/NET0131  & ~n2518 ;
  assign n2520 = ~n2501 & ~n2519 ;
  assign n2521 = \reg0_reg[20]/NET0131  & ~n1471 ;
  assign n2522 = \reg0_reg[20]/NET0131  & n290 ;
  assign n2527 = \reg0_reg[20]/NET0131  & ~n1444 ;
  assign n2528 = n1444 & ~n2352 ;
  assign n2529 = ~n2527 & ~n2528 ;
  assign n2530 = n798 & ~n2529 ;
  assign n2534 = n1444 & n2367 ;
  assign n2535 = ~n2527 & ~n2534 ;
  assign n2536 = n588 & ~n2535 ;
  assign n2531 = n1444 & ~n2358 ;
  assign n2532 = ~n2527 & ~n2531 ;
  assign n2533 = n881 & ~n2532 ;
  assign n2523 = n910 & n1016 ;
  assign n2524 = n907 & n2373 ;
  assign n2525 = ~n2523 & ~n2524 ;
  assign n2526 = n1444 & ~n2525 ;
  assign n2537 = \reg0_reg[20]/NET0131  & ~n1911 ;
  assign n2538 = ~n2526 & ~n2537 ;
  assign n2539 = ~n2533 & n2538 ;
  assign n2540 = ~n2536 & n2539 ;
  assign n2541 = ~n2530 & n2540 ;
  assign n2542 = n292 & ~n2541 ;
  assign n2543 = ~n2522 & ~n2542 ;
  assign n2544 = \state_reg[0]/NET0131  & ~n2543 ;
  assign n2545 = ~n2521 & ~n2544 ;
  assign n2546 = \reg0_reg[29]/NET0131  & ~n1444 ;
  assign n2547 = n1444 & ~n2097 ;
  assign n2548 = ~n2546 & ~n2547 ;
  assign n2549 = n588 & ~n2548 ;
  assign n2553 = n1444 & ~n2133 ;
  assign n2554 = ~n2546 & ~n2553 ;
  assign n2555 = n881 & ~n2554 ;
  assign n2550 = n1444 & n2167 ;
  assign n2551 = ~n2546 & ~n2550 ;
  assign n2552 = n798 & ~n2551 ;
  assign n2556 = n1444 & n2173 ;
  assign n2557 = ~n2546 & ~n2556 ;
  assign n2558 = n907 & ~n2557 ;
  assign n2559 = \reg0_reg[29]/NET0131  & ~n1459 ;
  assign n2560 = n1444 & n2178 ;
  assign n2561 = ~n2559 & ~n2560 ;
  assign n2562 = ~n2558 & n2561 ;
  assign n2563 = ~n2552 & n2562 ;
  assign n2564 = ~n2555 & n2563 ;
  assign n2565 = ~n2549 & n2564 ;
  assign n2566 = n292 & ~n2565 ;
  assign n2567 = \reg0_reg[29]/NET0131  & n290 ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = \state_reg[0]/NET0131  & ~n2568 ;
  assign n2570 = \reg0_reg[29]/NET0131  & ~n1471 ;
  assign n2571 = ~n2569 & ~n2570 ;
  assign n2572 = \reg1_reg[12]/NET0131  & ~n1471 ;
  assign n2573 = \reg1_reg[12]/NET0131  & n290 ;
  assign n2577 = \reg1_reg[12]/NET0131  & ~n1497 ;
  assign n2578 = n1497 & ~n1700 ;
  assign n2579 = ~n2577 & ~n2578 ;
  assign n2580 = n798 & ~n2579 ;
  assign n2587 = n1497 & n1720 ;
  assign n2588 = ~n2577 & ~n2587 ;
  assign n2589 = n907 & ~n2588 ;
  assign n2574 = \reg1_reg[12]/NET0131  & ~n1529 ;
  assign n2575 = ~n612 & n910 ;
  assign n2576 = n1497 & n2575 ;
  assign n2590 = ~n2574 & ~n2576 ;
  assign n2591 = ~n2589 & n2590 ;
  assign n2592 = ~n2580 & n2591 ;
  assign n2581 = n1497 & n1706 ;
  assign n2582 = ~n2577 & ~n2581 ;
  assign n2583 = n881 & ~n2582 ;
  assign n2584 = n1497 & n1714 ;
  assign n2585 = ~n2577 & ~n2584 ;
  assign n2586 = n588 & ~n2585 ;
  assign n2593 = ~n2583 & ~n2586 ;
  assign n2594 = n2592 & n2593 ;
  assign n2595 = n292 & ~n2594 ;
  assign n2596 = ~n2573 & ~n2595 ;
  assign n2597 = \state_reg[0]/NET0131  & ~n2596 ;
  assign n2598 = ~n2572 & ~n2597 ;
  assign n2599 = \reg1_reg[19]/NET0131  & ~n1471 ;
  assign n2600 = \reg1_reg[19]/NET0131  & n290 ;
  assign n2602 = \reg1_reg[19]/NET0131  & ~n1497 ;
  assign n2603 = n1497 & n1742 ;
  assign n2604 = ~n2602 & ~n2603 ;
  assign n2605 = n881 & ~n2604 ;
  assign n2606 = n1497 & ~n1748 ;
  assign n2607 = ~n2602 & ~n2606 ;
  assign n2608 = n798 & ~n2607 ;
  assign n2601 = n1497 & ~n2504 ;
  assign n2609 = \reg1_reg[19]/NET0131  & ~n1509 ;
  assign n2610 = ~n2601 & ~n2609 ;
  assign n2611 = ~n2608 & n2610 ;
  assign n2612 = ~n2605 & n2611 ;
  assign n2613 = n292 & ~n2612 ;
  assign n2614 = ~n2600 & ~n2613 ;
  assign n2615 = \state_reg[0]/NET0131  & ~n2614 ;
  assign n2616 = ~n2599 & ~n2615 ;
  assign n2617 = \reg1_reg[20]/NET0131  & ~n1471 ;
  assign n2618 = \reg1_reg[20]/NET0131  & n290 ;
  assign n2620 = \reg1_reg[20]/NET0131  & ~n1497 ;
  assign n2621 = n1497 & ~n2352 ;
  assign n2622 = ~n2620 & ~n2621 ;
  assign n2623 = n798 & ~n2622 ;
  assign n2627 = n1497 & n2367 ;
  assign n2628 = ~n2620 & ~n2627 ;
  assign n2629 = n588 & ~n2628 ;
  assign n2624 = n1497 & ~n2358 ;
  assign n2625 = ~n2620 & ~n2624 ;
  assign n2626 = n881 & ~n2625 ;
  assign n2619 = n1497 & ~n2525 ;
  assign n2630 = \reg1_reg[20]/NET0131  & ~n1507 ;
  assign n2631 = ~n2619 & ~n2630 ;
  assign n2632 = ~n2626 & n2631 ;
  assign n2633 = ~n2629 & n2632 ;
  assign n2634 = ~n2623 & n2633 ;
  assign n2635 = n292 & ~n2634 ;
  assign n2636 = ~n2618 & ~n2635 ;
  assign n2637 = \state_reg[0]/NET0131  & ~n2636 ;
  assign n2638 = ~n2617 & ~n2637 ;
  assign n2639 = \reg1_reg[26]/NET0131  & ~n1497 ;
  assign n2640 = n1497 & ~n2435 ;
  assign n2641 = ~n2639 & ~n2640 ;
  assign n2642 = n881 & ~n2641 ;
  assign n2643 = n1497 & n2443 ;
  assign n2644 = ~n2639 & ~n2643 ;
  assign n2645 = n588 & ~n2644 ;
  assign n2647 = n907 & n2452 ;
  assign n2646 = n910 & n953 ;
  assign n2648 = ~n2485 & ~n2646 ;
  assign n2649 = ~n2647 & n2648 ;
  assign n2650 = n1497 & ~n2649 ;
  assign n2651 = n1531 & ~n2017 ;
  assign n2652 = \reg1_reg[26]/NET0131  & ~n2651 ;
  assign n2653 = ~n2650 & ~n2652 ;
  assign n2654 = ~n2645 & n2653 ;
  assign n2655 = ~n2642 & n2654 ;
  assign n2656 = n292 & ~n2655 ;
  assign n2657 = \reg1_reg[26]/NET0131  & n290 ;
  assign n2658 = ~n2656 & ~n2657 ;
  assign n2659 = \state_reg[0]/NET0131  & ~n2658 ;
  assign n2660 = \reg1_reg[26]/NET0131  & ~n1471 ;
  assign n2661 = ~n2659 & ~n2660 ;
  assign n2662 = \reg1_reg[29]/NET0131  & ~n1497 ;
  assign n2663 = n1497 & ~n2097 ;
  assign n2664 = ~n2662 & ~n2663 ;
  assign n2665 = n588 & ~n2664 ;
  assign n2669 = n1497 & ~n2133 ;
  assign n2670 = ~n2662 & ~n2669 ;
  assign n2671 = n881 & ~n2670 ;
  assign n2666 = n1497 & n2167 ;
  assign n2667 = ~n2662 & ~n2666 ;
  assign n2668 = n798 & ~n2667 ;
  assign n2672 = n1497 & n2173 ;
  assign n2673 = ~n2662 & ~n2672 ;
  assign n2674 = n907 & ~n2673 ;
  assign n2675 = \reg1_reg[29]/NET0131  & ~n1529 ;
  assign n2676 = n1497 & n2178 ;
  assign n2677 = ~n2675 & ~n2676 ;
  assign n2678 = ~n2674 & n2677 ;
  assign n2679 = ~n2668 & n2678 ;
  assign n2680 = ~n2671 & n2679 ;
  assign n2681 = ~n2665 & n2680 ;
  assign n2682 = n292 & ~n2681 ;
  assign n2683 = \reg1_reg[29]/NET0131  & n290 ;
  assign n2684 = ~n2682 & ~n2683 ;
  assign n2685 = \state_reg[0]/NET0131  & ~n2684 ;
  assign n2686 = \reg1_reg[29]/NET0131  & ~n1471 ;
  assign n2687 = ~n2685 & ~n2686 ;
  assign n2688 = \reg2_reg[12]/NET0131  & ~n1471 ;
  assign n2689 = \reg2_reg[12]/NET0131  & n290 ;
  assign n2691 = \reg2_reg[12]/NET0131  & ~n1543 ;
  assign n2692 = n1543 & ~n1700 ;
  assign n2693 = ~n2691 & ~n2692 ;
  assign n2694 = n798 & ~n2693 ;
  assign n2701 = n1543 & n1720 ;
  assign n2702 = ~n2691 & ~n2701 ;
  assign n2703 = n907 & ~n2702 ;
  assign n2690 = \reg2_reg[12]/NET0131  & ~n1560 ;
  assign n2704 = n329 & n488 ;
  assign n2705 = n1543 & n2575 ;
  assign n2706 = ~n2704 & ~n2705 ;
  assign n2707 = ~n2690 & n2706 ;
  assign n2708 = ~n2703 & n2707 ;
  assign n2709 = ~n2694 & n2708 ;
  assign n2695 = n1543 & n1706 ;
  assign n2696 = ~n2691 & ~n2695 ;
  assign n2697 = n881 & ~n2696 ;
  assign n2698 = n1543 & n1714 ;
  assign n2699 = ~n2691 & ~n2698 ;
  assign n2700 = n588 & ~n2699 ;
  assign n2710 = ~n2697 & ~n2700 ;
  assign n2711 = n2709 & n2710 ;
  assign n2712 = n292 & ~n2711 ;
  assign n2713 = ~n2689 & ~n2712 ;
  assign n2714 = \state_reg[0]/NET0131  & ~n2713 ;
  assign n2715 = ~n2688 & ~n2714 ;
  assign n2716 = \reg2_reg[19]/NET0131  & ~n1471 ;
  assign n2717 = \reg2_reg[19]/NET0131  & n290 ;
  assign n2724 = n881 & n1742 ;
  assign n2723 = n798 & ~n1748 ;
  assign n2725 = n2504 & ~n2723 ;
  assign n2726 = ~n2724 & n2725 ;
  assign n2727 = n1543 & ~n2726 ;
  assign n2718 = n329 & n1044 ;
  assign n2719 = ~n588 & ~n797 ;
  assign n2720 = ~n1543 & ~n2719 ;
  assign n2721 = n2046 & ~n2720 ;
  assign n2722 = \reg2_reg[19]/NET0131  & ~n2721 ;
  assign n2728 = ~n2718 & ~n2722 ;
  assign n2729 = ~n2727 & n2728 ;
  assign n2730 = n292 & ~n2729 ;
  assign n2731 = ~n2717 & ~n2730 ;
  assign n2732 = \state_reg[0]/NET0131  & ~n2731 ;
  assign n2733 = ~n2716 & ~n2732 ;
  assign n2734 = \reg2_reg[20]/NET0131  & ~n1471 ;
  assign n2735 = \reg2_reg[20]/NET0131  & n290 ;
  assign n2737 = \reg2_reg[20]/NET0131  & ~n1543 ;
  assign n2738 = n1543 & ~n2352 ;
  assign n2739 = ~n2737 & ~n2738 ;
  assign n2740 = n798 & ~n2739 ;
  assign n2744 = n1543 & n2367 ;
  assign n2745 = ~n2737 & ~n2744 ;
  assign n2746 = n588 & ~n2745 ;
  assign n2741 = n1543 & ~n2358 ;
  assign n2742 = ~n2737 & ~n2741 ;
  assign n2743 = n881 & ~n2742 ;
  assign n2748 = n1543 & ~n2525 ;
  assign n2736 = \reg2_reg[20]/NET0131  & ~n2046 ;
  assign n2747 = n329 & n1022 ;
  assign n2749 = ~n2736 & ~n2747 ;
  assign n2750 = ~n2748 & n2749 ;
  assign n2751 = ~n2743 & n2750 ;
  assign n2752 = ~n2746 & n2751 ;
  assign n2753 = ~n2740 & n2752 ;
  assign n2754 = n292 & ~n2753 ;
  assign n2755 = ~n2735 & ~n2754 ;
  assign n2756 = \state_reg[0]/NET0131  & ~n2755 ;
  assign n2757 = ~n2734 & ~n2756 ;
  assign n2758 = \reg0_reg[12]/NET0131  & ~n1471 ;
  assign n2759 = \reg0_reg[12]/NET0131  & n290 ;
  assign n2762 = \reg0_reg[12]/NET0131  & ~n1444 ;
  assign n2763 = n1444 & n1706 ;
  assign n2764 = ~n2762 & ~n2763 ;
  assign n2765 = n881 & ~n2764 ;
  assign n2772 = n1444 & n1720 ;
  assign n2773 = ~n2762 & ~n2772 ;
  assign n2774 = n907 & ~n2773 ;
  assign n2760 = \reg0_reg[12]/NET0131  & ~n1459 ;
  assign n2761 = n1444 & n2575 ;
  assign n2775 = ~n2760 & ~n2761 ;
  assign n2776 = ~n2774 & n2775 ;
  assign n2777 = ~n2765 & n2776 ;
  assign n2766 = n1444 & ~n1700 ;
  assign n2767 = ~n2762 & ~n2766 ;
  assign n2768 = n798 & ~n2767 ;
  assign n2769 = n1444 & n1714 ;
  assign n2770 = ~n2762 & ~n2769 ;
  assign n2771 = n588 & ~n2770 ;
  assign n2778 = ~n2768 & ~n2771 ;
  assign n2779 = n2777 & n2778 ;
  assign n2780 = n292 & ~n2779 ;
  assign n2781 = ~n2759 & ~n2780 ;
  assign n2782 = \state_reg[0]/NET0131  & ~n2781 ;
  assign n2783 = ~n2758 & ~n2782 ;
  assign n2786 = ~n308 & n572 ;
  assign n2787 = ~n1153 & ~n1195 ;
  assign n2788 = n2421 & n2787 ;
  assign n2789 = ~n2421 & ~n2787 ;
  assign n2790 = ~n2788 & ~n2789 ;
  assign n2791 = n308 & ~n2790 ;
  assign n2792 = ~n2786 & ~n2791 ;
  assign n2793 = n881 & ~n2792 ;
  assign n2794 = ~n579 & n1048 ;
  assign n2795 = ~n1408 & ~n2794 ;
  assign n2796 = ~n341 & ~n2795 ;
  assign n2797 = n341 & n566 ;
  assign n2798 = ~n2796 & ~n2797 ;
  assign n2799 = n308 & n2798 ;
  assign n2800 = ~n2786 & ~n2799 ;
  assign n2801 = n588 & ~n2800 ;
  assign n2802 = ~n903 & n1038 ;
  assign n2803 = n907 & ~n1759 ;
  assign n2804 = ~n2802 & n2803 ;
  assign n2806 = ~n2472 & ~n2787 ;
  assign n2805 = n2472 & n2787 ;
  assign n2807 = n798 & ~n2805 ;
  assign n2808 = ~n2806 & n2807 ;
  assign n2809 = ~n2804 & ~n2808 ;
  assign n2810 = n308 & ~n2809 ;
  assign n2785 = n333 & n1038 ;
  assign n2811 = ~n798 & ~n907 ;
  assign n2812 = ~n308 & ~n2811 ;
  assign n2813 = n912 & ~n2812 ;
  assign n2814 = n572 & ~n2813 ;
  assign n2815 = ~n2785 & ~n2814 ;
  assign n2816 = ~n2810 & n2815 ;
  assign n2817 = ~n2801 & n2816 ;
  assign n2818 = ~n2793 & n2817 ;
  assign n2819 = n292 & ~n2818 ;
  assign n2820 = n290 & n572 ;
  assign n2821 = ~n2819 & ~n2820 ;
  assign n2822 = \state_reg[0]/NET0131  & ~n2821 ;
  assign n2784 = n260 & n572 ;
  assign n2823 = \reg3_reg[18]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2824 = ~n2784 & ~n2823 ;
  assign n2825 = ~n2822 & n2824 ;
  assign n2826 = \reg2_reg[25]/NET0131  & ~n1471 ;
  assign n2827 = \reg2_reg[25]/NET0131  & n290 ;
  assign n2828 = \reg2_reg[25]/NET0131  & ~n1543 ;
  assign n2851 = ~n974 & n1868 ;
  assign n2852 = ~n962 & ~n2851 ;
  assign n2853 = n962 & n2851 ;
  assign n2854 = ~n2852 & ~n2853 ;
  assign n2855 = ~n341 & ~n2854 ;
  assign n2856 = n341 & ~n985 ;
  assign n2857 = ~n2855 & ~n2856 ;
  assign n2858 = n1543 & ~n2857 ;
  assign n2859 = ~n2828 & ~n2858 ;
  assign n2860 = n588 & ~n2859 ;
  assign n2829 = ~n1212 & ~n1230 ;
  assign n2862 = n787 & n2142 ;
  assign n2861 = ~n686 & n2141 ;
  assign n2863 = n2146 & ~n2861 ;
  assign n2864 = ~n2862 & n2863 ;
  assign n2865 = n2149 & ~n2864 ;
  assign n2866 = n2157 & ~n2865 ;
  assign n2867 = n2829 & ~n2866 ;
  assign n2868 = ~n2829 & n2866 ;
  assign n2869 = ~n2867 & ~n2868 ;
  assign n2870 = n1543 & ~n2869 ;
  assign n2871 = ~n2828 & ~n2870 ;
  assign n2872 = n798 & ~n2871 ;
  assign n2831 = n873 & n2110 ;
  assign n2830 = ~n832 & n2109 ;
  assign n2832 = n2114 & ~n2830 ;
  assign n2833 = ~n2831 & n2832 ;
  assign n2834 = n2117 & ~n2833 ;
  assign n2835 = n2123 & ~n2834 ;
  assign n2836 = n2829 & n2835 ;
  assign n2837 = ~n2829 & ~n2835 ;
  assign n2838 = ~n2836 & ~n2837 ;
  assign n2839 = n1543 & ~n2838 ;
  assign n2840 = ~n2828 & ~n2839 ;
  assign n2841 = n881 & ~n2840 ;
  assign n2843 = n965 & ~n1252 ;
  assign n2844 = ~n2450 & ~n2843 ;
  assign n2845 = n1543 & n2844 ;
  assign n2846 = ~n2828 & ~n2845 ;
  assign n2847 = n907 & ~n2846 ;
  assign n2842 = \reg2_reg[25]/NET0131  & ~n1560 ;
  assign n2848 = n329 & n970 ;
  assign n2849 = n910 & n965 ;
  assign n2850 = n1543 & n2849 ;
  assign n2873 = ~n2848 & ~n2850 ;
  assign n2874 = ~n2842 & n2873 ;
  assign n2875 = ~n2847 & n2874 ;
  assign n2876 = ~n2841 & n2875 ;
  assign n2877 = ~n2872 & n2876 ;
  assign n2878 = ~n2860 & n2877 ;
  assign n2879 = n292 & ~n2878 ;
  assign n2880 = ~n2827 & ~n2879 ;
  assign n2881 = \state_reg[0]/NET0131  & ~n2880 ;
  assign n2882 = ~n2826 & ~n2881 ;
  assign n2883 = ~n308 & n997 ;
  assign n2884 = ~n1205 & ~n1223 ;
  assign n2885 = ~n2215 & n2458 ;
  assign n2886 = n2461 & ~n2885 ;
  assign n2887 = n2457 & ~n2886 ;
  assign n2888 = n2477 & ~n2887 ;
  assign n2889 = n2884 & n2888 ;
  assign n2890 = ~n2884 & ~n2888 ;
  assign n2891 = ~n2889 & ~n2890 ;
  assign n2892 = n308 & n2891 ;
  assign n2893 = ~n2883 & ~n2892 ;
  assign n2894 = n798 & ~n2893 ;
  assign n2895 = n2420 & n2423 ;
  assign n2896 = ~n2418 & n2423 ;
  assign n2897 = n2428 & ~n2896 ;
  assign n2898 = ~n2895 & n2897 ;
  assign n2899 = n2884 & n2898 ;
  assign n2900 = ~n2884 & ~n2898 ;
  assign n2901 = ~n2899 & ~n2900 ;
  assign n2902 = n308 & ~n2901 ;
  assign n2903 = ~n2883 & ~n2902 ;
  assign n2904 = n881 & ~n2903 ;
  assign n2906 = n341 & ~n1014 ;
  assign n2907 = n1263 & n1752 ;
  assign n2908 = n934 & ~n2907 ;
  assign n2909 = ~n341 & ~n1409 ;
  assign n2910 = ~n2908 & n2909 ;
  assign n2911 = ~n2906 & ~n2910 ;
  assign n2912 = n588 & ~n2911 ;
  assign n2913 = ~n1004 & n2371 ;
  assign n2914 = n991 & ~n2913 ;
  assign n2915 = n907 & ~n1877 ;
  assign n2916 = ~n2914 & n2915 ;
  assign n2917 = ~n2912 & ~n2916 ;
  assign n2918 = n308 & ~n2917 ;
  assign n2905 = n997 & ~n1736 ;
  assign n2919 = n333 & n991 ;
  assign n2920 = ~n2905 & ~n2919 ;
  assign n2921 = ~n2918 & n2920 ;
  assign n2922 = ~n2904 & n2921 ;
  assign n2923 = ~n2894 & n2922 ;
  assign n2924 = n292 & ~n2923 ;
  assign n2925 = n290 & n997 ;
  assign n2926 = ~n2924 & ~n2925 ;
  assign n2927 = \state_reg[0]/NET0131  & ~n2926 ;
  assign n2928 = \reg3_reg[22]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2929 = n260 & n997 ;
  assign n2930 = ~n2928 & ~n2929 ;
  assign n2931 = ~n2927 & n2930 ;
  assign n2932 = \reg2_reg[30]/NET0131  & ~n1471 ;
  assign n2933 = \reg2_reg[30]/NET0131  & n290 ;
  assign n2941 = ~n2171 & n2403 ;
  assign n2942 = ~n2404 & ~n2941 ;
  assign n2943 = n1543 & ~n2942 ;
  assign n2944 = ~\reg2_reg[30]/NET0131  & ~n1543 ;
  assign n2945 = n907 & ~n2944 ;
  assign n2946 = ~n2943 & n2945 ;
  assign n2938 = n910 & n2403 ;
  assign n2939 = ~n2402 & ~n2938 ;
  assign n2940 = n1543 & ~n2939 ;
  assign n2934 = n319 & ~n322 ;
  assign n2935 = ~n1543 & ~n2934 ;
  assign n2936 = ~n909 & ~n2935 ;
  assign n2937 = \reg2_reg[30]/NET0131  & ~n2936 ;
  assign n2947 = ~n2177 & ~n2937 ;
  assign n2948 = ~n2940 & n2947 ;
  assign n2949 = ~n2946 & n2948 ;
  assign n2950 = n292 & ~n2949 ;
  assign n2951 = ~n2933 & ~n2950 ;
  assign n2952 = \state_reg[0]/NET0131  & ~n2951 ;
  assign n2953 = ~n2932 & ~n2952 ;
  assign n2954 = \reg0_reg[16]/NET0131  & ~n1471 ;
  assign n2955 = \reg0_reg[16]/NET0131  & n290 ;
  assign n2960 = \reg0_reg[16]/NET0131  & ~n1444 ;
  assign n2964 = n1444 & n2273 ;
  assign n2965 = ~n2960 & ~n2964 ;
  assign n2966 = n881 & ~n2965 ;
  assign n2961 = n1444 & ~n2265 ;
  assign n2962 = ~n2960 & ~n2961 ;
  assign n2963 = n798 & ~n2962 ;
  assign n2967 = n1444 & n2281 ;
  assign n2968 = ~n2960 & ~n2967 ;
  assign n2969 = n588 & ~n2968 ;
  assign n2956 = ~n662 & n910 ;
  assign n2957 = n907 & n2286 ;
  assign n2958 = ~n2956 & ~n2957 ;
  assign n2959 = n1444 & ~n2958 ;
  assign n2970 = \reg0_reg[16]/NET0131  & ~n1911 ;
  assign n2971 = ~n2959 & ~n2970 ;
  assign n2972 = ~n2969 & n2971 ;
  assign n2973 = ~n2963 & n2972 ;
  assign n2974 = ~n2966 & n2973 ;
  assign n2975 = n292 & ~n2974 ;
  assign n2976 = ~n2955 & ~n2975 ;
  assign n2977 = \state_reg[0]/NET0131  & ~n2976 ;
  assign n2978 = ~n2954 & ~n2977 ;
  assign n2979 = \reg2_reg[7]/NET0131  & ~n1471 ;
  assign n2980 = \reg2_reg[7]/NET0131  & n290 ;
  assign n2982 = \reg2_reg[7]/NET0131  & ~n1543 ;
  assign n2983 = n1543 & n2315 ;
  assign n2984 = ~n2982 & ~n2983 ;
  assign n2985 = n588 & ~n2984 ;
  assign n2989 = n1543 & ~n2328 ;
  assign n2990 = ~n2982 & ~n2989 ;
  assign n2991 = n798 & ~n2990 ;
  assign n2986 = n1543 & n2322 ;
  assign n2987 = ~n2982 & ~n2986 ;
  assign n2988 = n881 & ~n2987 ;
  assign n2993 = ~n698 & n910 ;
  assign n2994 = ~n2306 & ~n2993 ;
  assign n2995 = n1543 & ~n2994 ;
  assign n2981 = \reg2_reg[7]/NET0131  & ~n1585 ;
  assign n2992 = n329 & n479 ;
  assign n2996 = ~n2981 & ~n2992 ;
  assign n2997 = ~n2995 & n2996 ;
  assign n2998 = ~n2988 & n2997 ;
  assign n2999 = ~n2991 & n2998 ;
  assign n3000 = ~n2985 & n2999 ;
  assign n3001 = n292 & ~n3000 ;
  assign n3002 = ~n2980 & ~n3001 ;
  assign n3003 = \state_reg[0]/NET0131  & ~n3002 ;
  assign n3004 = ~n2979 & ~n3003 ;
  assign n3005 = \reg0_reg[22]/NET0131  & ~n1444 ;
  assign n3006 = n1444 & n2891 ;
  assign n3007 = ~n3005 & ~n3006 ;
  assign n3008 = n798 & ~n3007 ;
  assign n3009 = n1444 & ~n2901 ;
  assign n3010 = ~n3005 & ~n3009 ;
  assign n3011 = n881 & ~n3010 ;
  assign n3012 = n910 & n991 ;
  assign n3013 = n2917 & ~n3012 ;
  assign n3014 = n1444 & ~n3013 ;
  assign n3015 = \reg0_reg[22]/NET0131  & ~n1462 ;
  assign n3016 = ~n3014 & ~n3015 ;
  assign n3017 = ~n3011 & n3016 ;
  assign n3018 = ~n3008 & n3017 ;
  assign n3019 = n292 & ~n3018 ;
  assign n3020 = \reg0_reg[22]/NET0131  & n290 ;
  assign n3021 = ~n3019 & ~n3020 ;
  assign n3022 = \state_reg[0]/NET0131  & ~n3021 ;
  assign n3023 = \reg0_reg[22]/NET0131  & ~n1471 ;
  assign n3024 = ~n3022 & ~n3023 ;
  assign n3025 = \reg0_reg[26]/NET0131  & ~n1444 ;
  assign n3026 = n1444 & ~n2435 ;
  assign n3027 = ~n3025 & ~n3026 ;
  assign n3028 = n881 & ~n3027 ;
  assign n3029 = n1444 & n2443 ;
  assign n3030 = ~n3025 & ~n3029 ;
  assign n3031 = n588 & ~n3030 ;
  assign n3032 = n1444 & ~n2649 ;
  assign n3033 = ~n798 & ~n1422 ;
  assign n3034 = ~n1444 & ~n3033 ;
  assign n3035 = n1458 & ~n3034 ;
  assign n3036 = \reg0_reg[26]/NET0131  & ~n3035 ;
  assign n3037 = ~n3032 & ~n3036 ;
  assign n3038 = ~n3031 & n3037 ;
  assign n3039 = ~n3028 & n3038 ;
  assign n3040 = n292 & ~n3039 ;
  assign n3041 = \reg0_reg[26]/NET0131  & n290 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3043 = \state_reg[0]/NET0131  & ~n3042 ;
  assign n3044 = \reg0_reg[26]/NET0131  & ~n1471 ;
  assign n3045 = ~n3043 & ~n3044 ;
  assign n3046 = n907 & n2942 ;
  assign n3047 = n2939 & ~n3046 ;
  assign n3048 = n1444 & n2389 ;
  assign n3049 = ~n3047 & n3048 ;
  assign n3050 = n1458 & n3048 ;
  assign n3051 = \reg0_reg[30]/NET0131  & ~n3050 ;
  assign n3052 = ~n3049 & ~n3051 ;
  assign n3053 = ~n2410 & n3048 ;
  assign n3054 = \reg0_reg[31]/NET0131  & ~n3050 ;
  assign n3055 = ~n3053 & ~n3054 ;
  assign n3056 = \reg0_reg[7]/NET0131  & ~n1471 ;
  assign n3057 = \reg0_reg[7]/NET0131  & n290 ;
  assign n3059 = \reg0_reg[7]/NET0131  & ~n1444 ;
  assign n3060 = n1444 & n2315 ;
  assign n3061 = ~n3059 & ~n3060 ;
  assign n3062 = n588 & ~n3061 ;
  assign n3066 = n1444 & ~n2328 ;
  assign n3067 = ~n3059 & ~n3066 ;
  assign n3068 = n798 & ~n3067 ;
  assign n3063 = n1444 & n2322 ;
  assign n3064 = ~n3059 & ~n3063 ;
  assign n3065 = n881 & ~n3064 ;
  assign n3058 = \reg0_reg[7]/NET0131  & ~n1911 ;
  assign n3069 = n1444 & ~n2994 ;
  assign n3070 = ~n3058 & ~n3069 ;
  assign n3071 = ~n3065 & n3070 ;
  assign n3072 = ~n3068 & n3071 ;
  assign n3073 = ~n3062 & n3072 ;
  assign n3074 = n292 & ~n3073 ;
  assign n3075 = ~n3057 & ~n3074 ;
  assign n3076 = \state_reg[0]/NET0131  & ~n3075 ;
  assign n3077 = ~n3056 & ~n3076 ;
  assign n3078 = \reg0_reg[8]/NET0131  & ~n1471 ;
  assign n3079 = \reg0_reg[8]/NET0131  & n290 ;
  assign n3081 = \reg0_reg[8]/NET0131  & ~n1444 ;
  assign n3095 = n341 & ~n483 ;
  assign n3096 = n474 & ~n2311 ;
  assign n3097 = ~n341 & ~n486 ;
  assign n3098 = ~n3096 & n3097 ;
  assign n3099 = ~n3095 & ~n3098 ;
  assign n3100 = n1444 & ~n3099 ;
  assign n3101 = ~n3081 & ~n3100 ;
  assign n3102 = n588 & ~n3101 ;
  assign n3082 = ~n706 & ~n728 ;
  assign n3089 = n1178 & n3082 ;
  assign n3090 = ~n1178 & ~n3082 ;
  assign n3091 = ~n3089 & ~n3090 ;
  assign n3092 = n1444 & n3091 ;
  assign n3093 = ~n3081 & ~n3092 ;
  assign n3094 = n881 & ~n3093 ;
  assign n3083 = n1096 & n3082 ;
  assign n3084 = ~n1096 & ~n3082 ;
  assign n3085 = ~n3083 & ~n3084 ;
  assign n3086 = n1444 & ~n3085 ;
  assign n3087 = ~n3081 & ~n3086 ;
  assign n3088 = n798 & ~n3087 ;
  assign n3103 = ~n705 & ~n889 ;
  assign n3104 = n705 & n889 ;
  assign n3105 = ~n3103 & ~n3104 ;
  assign n3106 = n1444 & n3105 ;
  assign n3107 = ~n3081 & ~n3106 ;
  assign n3108 = n907 & ~n3107 ;
  assign n3080 = \reg0_reg[8]/NET0131  & ~n1459 ;
  assign n3109 = ~n705 & n910 ;
  assign n3110 = n1444 & n3109 ;
  assign n3111 = ~n3080 & ~n3110 ;
  assign n3112 = ~n3108 & n3111 ;
  assign n3113 = ~n3088 & n3112 ;
  assign n3114 = ~n3094 & n3113 ;
  assign n3115 = ~n3102 & n3114 ;
  assign n3116 = n292 & ~n3115 ;
  assign n3117 = ~n3079 & ~n3116 ;
  assign n3118 = \state_reg[0]/NET0131  & ~n3117 ;
  assign n3119 = ~n3078 & ~n3118 ;
  assign n3120 = \reg1_reg[11]/NET0131  & ~n1471 ;
  assign n3121 = \reg1_reg[11]/NET0131  & n290 ;
  assign n3123 = \reg1_reg[11]/NET0131  & ~n1497 ;
  assign n3124 = n1497 & ~n1654 ;
  assign n3125 = ~n3123 & ~n3124 ;
  assign n3126 = n798 & ~n3125 ;
  assign n3133 = n1497 & n1676 ;
  assign n3134 = ~n3123 & ~n3133 ;
  assign n3135 = n907 & ~n3134 ;
  assign n3122 = \reg1_reg[11]/NET0131  & ~n1529 ;
  assign n3136 = ~n602 & n910 ;
  assign n3137 = n1497 & n3136 ;
  assign n3138 = ~n3122 & ~n3137 ;
  assign n3139 = ~n3135 & n3138 ;
  assign n3140 = ~n3126 & n3139 ;
  assign n3127 = n1497 & n1663 ;
  assign n3128 = ~n3123 & ~n3127 ;
  assign n3129 = n588 & ~n3128 ;
  assign n3130 = n1497 & n1669 ;
  assign n3131 = ~n3123 & ~n3130 ;
  assign n3132 = n881 & ~n3131 ;
  assign n3141 = ~n3129 & ~n3132 ;
  assign n3142 = n3140 & n3141 ;
  assign n3143 = n292 & ~n3142 ;
  assign n3144 = ~n3121 & ~n3143 ;
  assign n3145 = \state_reg[0]/NET0131  & ~n3144 ;
  assign n3146 = ~n3120 & ~n3145 ;
  assign n3147 = \reg1_reg[14]/NET0131  & ~n1471 ;
  assign n3148 = \reg1_reg[14]/NET0131  & n290 ;
  assign n3150 = \reg1_reg[14]/NET0131  & ~n1497 ;
  assign n3151 = n1497 & n2201 ;
  assign n3152 = ~n3150 & ~n3151 ;
  assign n3153 = n588 & ~n3152 ;
  assign n3157 = n1497 & n2236 ;
  assign n3158 = ~n3150 & ~n3157 ;
  assign n3159 = n881 & ~n3158 ;
  assign n3154 = n1497 & ~n2219 ;
  assign n3155 = ~n3150 & ~n3154 ;
  assign n3156 = n798 & ~n3155 ;
  assign n3149 = \reg1_reg[14]/NET0131  & ~n1507 ;
  assign n3160 = ~n646 & n910 ;
  assign n3161 = n907 & n2241 ;
  assign n3162 = ~n3160 & ~n3161 ;
  assign n3163 = n1497 & ~n3162 ;
  assign n3164 = ~n3149 & ~n3163 ;
  assign n3165 = ~n3156 & n3164 ;
  assign n3166 = ~n3159 & n3165 ;
  assign n3167 = ~n3153 & n3166 ;
  assign n3168 = n292 & ~n3167 ;
  assign n3169 = ~n3148 & ~n3168 ;
  assign n3170 = \state_reg[0]/NET0131  & ~n3169 ;
  assign n3171 = ~n3147 & ~n3170 ;
  assign n3172 = \reg1_reg[16]/NET0131  & ~n1471 ;
  assign n3173 = \reg1_reg[16]/NET0131  & n290 ;
  assign n3175 = \reg1_reg[16]/NET0131  & ~n1497 ;
  assign n3179 = n1497 & n2273 ;
  assign n3180 = ~n3175 & ~n3179 ;
  assign n3181 = n881 & ~n3180 ;
  assign n3176 = n1497 & ~n2265 ;
  assign n3177 = ~n3175 & ~n3176 ;
  assign n3178 = n798 & ~n3177 ;
  assign n3182 = n1497 & n2281 ;
  assign n3183 = ~n3175 & ~n3182 ;
  assign n3184 = n588 & ~n3183 ;
  assign n3174 = n1497 & ~n2958 ;
  assign n3185 = \reg1_reg[16]/NET0131  & ~n1507 ;
  assign n3186 = ~n3174 & ~n3185 ;
  assign n3187 = ~n3184 & n3186 ;
  assign n3188 = ~n3178 & n3187 ;
  assign n3189 = ~n3181 & n3188 ;
  assign n3190 = n292 & ~n3189 ;
  assign n3191 = ~n3173 & ~n3190 ;
  assign n3192 = \state_reg[0]/NET0131  & ~n3191 ;
  assign n3193 = ~n3172 & ~n3192 ;
  assign n3194 = \reg1_reg[22]/NET0131  & ~n1497 ;
  assign n3195 = n1497 & n2891 ;
  assign n3196 = ~n3194 & ~n3195 ;
  assign n3197 = n798 & ~n3196 ;
  assign n3198 = n1497 & ~n2901 ;
  assign n3199 = ~n3194 & ~n3198 ;
  assign n3200 = n881 & ~n3199 ;
  assign n3201 = n1497 & ~n3013 ;
  assign n3202 = \reg1_reg[22]/NET0131  & ~n1509 ;
  assign n3203 = ~n3201 & ~n3202 ;
  assign n3204 = ~n3200 & n3203 ;
  assign n3205 = ~n3197 & n3204 ;
  assign n3206 = n292 & ~n3205 ;
  assign n3207 = \reg1_reg[22]/NET0131  & n290 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = \state_reg[0]/NET0131  & ~n3208 ;
  assign n3210 = \reg1_reg[22]/NET0131  & ~n1471 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3212 = n1497 & n2389 ;
  assign n3213 = ~n2410 & n3212 ;
  assign n3214 = n1458 & n3212 ;
  assign n3215 = \reg1_reg[31]/NET0131  & ~n3214 ;
  assign n3216 = ~n3213 & ~n3215 ;
  assign n3217 = \reg1_reg[30]/NET0131  & ~n1471 ;
  assign n3218 = n1497 & ~n3047 ;
  assign n3219 = n1458 & n1497 ;
  assign n3220 = \reg1_reg[30]/NET0131  & ~n3219 ;
  assign n3221 = ~n3218 & ~n3220 ;
  assign n3222 = n292 & ~n3221 ;
  assign n3223 = \reg1_reg[30]/NET0131  & n290 ;
  assign n3224 = ~n3222 & ~n3223 ;
  assign n3225 = \state_reg[0]/NET0131  & ~n3224 ;
  assign n3226 = ~n3217 & ~n3225 ;
  assign n3227 = \reg1_reg[7]/NET0131  & ~n1471 ;
  assign n3228 = \reg1_reg[7]/NET0131  & n290 ;
  assign n3230 = \reg1_reg[7]/NET0131  & ~n1497 ;
  assign n3231 = n1497 & n2315 ;
  assign n3232 = ~n3230 & ~n3231 ;
  assign n3233 = n588 & ~n3232 ;
  assign n3237 = n1497 & n2322 ;
  assign n3238 = ~n3230 & ~n3237 ;
  assign n3239 = n881 & ~n3238 ;
  assign n3234 = n1497 & ~n2328 ;
  assign n3235 = ~n3230 & ~n3234 ;
  assign n3236 = n798 & ~n3235 ;
  assign n3229 = \reg1_reg[7]/NET0131  & ~n1531 ;
  assign n3240 = n1497 & ~n2994 ;
  assign n3241 = ~n3229 & ~n3240 ;
  assign n3242 = ~n3236 & n3241 ;
  assign n3243 = ~n3239 & n3242 ;
  assign n3244 = ~n3233 & n3243 ;
  assign n3245 = n292 & ~n3244 ;
  assign n3246 = ~n3228 & ~n3245 ;
  assign n3247 = \state_reg[0]/NET0131  & ~n3246 ;
  assign n3248 = ~n3227 & ~n3247 ;
  assign n3249 = \reg0_reg[11]/NET0131  & ~n1471 ;
  assign n3250 = \reg0_reg[11]/NET0131  & n290 ;
  assign n3252 = \reg0_reg[11]/NET0131  & ~n1444 ;
  assign n3253 = n1444 & ~n1654 ;
  assign n3254 = ~n3252 & ~n3253 ;
  assign n3255 = n798 & ~n3254 ;
  assign n3262 = n1444 & n1676 ;
  assign n3263 = ~n3252 & ~n3262 ;
  assign n3264 = n907 & ~n3263 ;
  assign n3251 = \reg0_reg[11]/NET0131  & ~n1459 ;
  assign n3265 = n1444 & n3136 ;
  assign n3266 = ~n3251 & ~n3265 ;
  assign n3267 = ~n3264 & n3266 ;
  assign n3268 = ~n3255 & n3267 ;
  assign n3256 = n1444 & n1663 ;
  assign n3257 = ~n3252 & ~n3256 ;
  assign n3258 = n588 & ~n3257 ;
  assign n3259 = n1444 & n1669 ;
  assign n3260 = ~n3252 & ~n3259 ;
  assign n3261 = n881 & ~n3260 ;
  assign n3269 = ~n3258 & ~n3261 ;
  assign n3270 = n3268 & n3269 ;
  assign n3271 = n292 & ~n3270 ;
  assign n3272 = ~n3250 & ~n3271 ;
  assign n3273 = \state_reg[0]/NET0131  & ~n3272 ;
  assign n3274 = ~n3249 & ~n3273 ;
  assign n3275 = \reg2_reg[14]/NET0131  & ~n1471 ;
  assign n3276 = \reg2_reg[14]/NET0131  & n290 ;
  assign n3278 = \reg2_reg[14]/NET0131  & ~n1543 ;
  assign n3279 = n1543 & n2201 ;
  assign n3280 = ~n3278 & ~n3279 ;
  assign n3281 = n588 & ~n3280 ;
  assign n3285 = n1543 & n2236 ;
  assign n3286 = ~n3278 & ~n3285 ;
  assign n3287 = n881 & ~n3286 ;
  assign n3282 = n1543 & ~n2219 ;
  assign n3283 = ~n3278 & ~n3282 ;
  assign n3284 = n798 & ~n3283 ;
  assign n3289 = n1543 & ~n3162 ;
  assign n3277 = \reg2_reg[14]/NET0131  & ~n2046 ;
  assign n3288 = n329 & n542 ;
  assign n3290 = ~n3277 & ~n3288 ;
  assign n3291 = ~n3289 & n3290 ;
  assign n3292 = ~n3284 & n3291 ;
  assign n3293 = ~n3287 & n3292 ;
  assign n3294 = ~n3281 & n3293 ;
  assign n3295 = n292 & ~n3294 ;
  assign n3296 = ~n3276 & ~n3295 ;
  assign n3297 = \state_reg[0]/NET0131  & ~n3296 ;
  assign n3298 = ~n3275 & ~n3297 ;
  assign n3299 = \reg2_reg[16]/NET0131  & ~n1471 ;
  assign n3300 = \reg2_reg[16]/NET0131  & n290 ;
  assign n3302 = \reg2_reg[16]/NET0131  & ~n1543 ;
  assign n3306 = n1543 & n2273 ;
  assign n3307 = ~n3302 & ~n3306 ;
  assign n3308 = n881 & ~n3307 ;
  assign n3303 = n1543 & ~n2265 ;
  assign n3304 = ~n3302 & ~n3303 ;
  assign n3305 = n798 & ~n3304 ;
  assign n3309 = n1543 & n2281 ;
  assign n3310 = ~n3302 & ~n3309 ;
  assign n3311 = n588 & ~n3310 ;
  assign n3301 = n1543 & ~n2958 ;
  assign n3312 = n329 & n551 ;
  assign n3313 = \reg2_reg[16]/NET0131  & ~n2046 ;
  assign n3314 = ~n3312 & ~n3313 ;
  assign n3315 = ~n3301 & n3314 ;
  assign n3316 = ~n3311 & n3315 ;
  assign n3317 = ~n3305 & n3316 ;
  assign n3318 = ~n3308 & n3317 ;
  assign n3319 = n292 & ~n3318 ;
  assign n3320 = ~n3300 & ~n3319 ;
  assign n3321 = \state_reg[0]/NET0131  & ~n3320 ;
  assign n3322 = ~n3299 & ~n3321 ;
  assign n3323 = \reg2_reg[22]/NET0131  & ~n1543 ;
  assign n3324 = n1543 & n2891 ;
  assign n3325 = ~n3323 & ~n3324 ;
  assign n3326 = n798 & ~n3325 ;
  assign n3327 = n1543 & ~n2901 ;
  assign n3328 = ~n3323 & ~n3327 ;
  assign n3329 = n881 & ~n3328 ;
  assign n3330 = n1543 & ~n3013 ;
  assign n3331 = n329 & n997 ;
  assign n3332 = ~n1583 & n2046 ;
  assign n3333 = \reg2_reg[22]/NET0131  & ~n3332 ;
  assign n3334 = ~n3331 & ~n3333 ;
  assign n3335 = ~n3330 & n3334 ;
  assign n3336 = ~n3329 & n3335 ;
  assign n3337 = ~n3326 & n3336 ;
  assign n3338 = n292 & ~n3337 ;
  assign n3339 = \reg2_reg[22]/NET0131  & n290 ;
  assign n3340 = ~n3338 & ~n3339 ;
  assign n3341 = \state_reg[0]/NET0131  & ~n3340 ;
  assign n3342 = \reg2_reg[22]/NET0131  & ~n1471 ;
  assign n3343 = ~n3341 & ~n3342 ;
  assign n3344 = \reg0_reg[14]/NET0131  & ~n1471 ;
  assign n3345 = \reg0_reg[14]/NET0131  & n290 ;
  assign n3347 = \reg0_reg[14]/NET0131  & ~n1444 ;
  assign n3348 = n1444 & n2201 ;
  assign n3349 = ~n3347 & ~n3348 ;
  assign n3350 = n588 & ~n3349 ;
  assign n3354 = n1444 & n2236 ;
  assign n3355 = ~n3347 & ~n3354 ;
  assign n3356 = n881 & ~n3355 ;
  assign n3351 = n1444 & ~n2219 ;
  assign n3352 = ~n3347 & ~n3351 ;
  assign n3353 = n798 & ~n3352 ;
  assign n3346 = \reg0_reg[14]/NET0131  & ~n1911 ;
  assign n3357 = n1444 & ~n3162 ;
  assign n3358 = ~n3346 & ~n3357 ;
  assign n3359 = ~n3353 & n3358 ;
  assign n3360 = ~n3356 & n3359 ;
  assign n3361 = ~n3350 & n3360 ;
  assign n3362 = n292 & ~n3361 ;
  assign n3363 = ~n3345 & ~n3362 ;
  assign n3364 = \state_reg[0]/NET0131  & ~n3363 ;
  assign n3365 = ~n3344 & ~n3364 ;
  assign n3366 = \reg3_reg[1]/NET0131  & ~n1471 ;
  assign n3367 = \reg3_reg[1]/NET0131  & n290 ;
  assign n3372 = ~n747 & ~n751 ;
  assign n3373 = ~n883 & ~n3372 ;
  assign n3374 = n907 & n3373 ;
  assign n3375 = n382 & ~n417 ;
  assign n3376 = ~n418 & ~n3375 ;
  assign n3377 = ~n341 & ~n3376 ;
  assign n3378 = n341 & n396 ;
  assign n3379 = n588 & ~n3378 ;
  assign n3380 = ~n3377 & n3379 ;
  assign n3381 = ~n748 & ~n754 ;
  assign n3383 = ~n752 & n3381 ;
  assign n3382 = n752 & ~n3381 ;
  assign n3384 = n798 & ~n3382 ;
  assign n3385 = ~n3383 & n3384 ;
  assign n3387 = n855 & ~n3381 ;
  assign n3386 = ~n855 & n3381 ;
  assign n3388 = n881 & ~n3386 ;
  assign n3389 = ~n3387 & n3388 ;
  assign n3390 = ~n3385 & ~n3389 ;
  assign n3391 = ~n3380 & n3390 ;
  assign n3392 = ~n3374 & n3391 ;
  assign n3393 = n308 & ~n3392 ;
  assign n3368 = ~n308 & ~n332 ;
  assign n3369 = n912 & ~n3368 ;
  assign n3370 = \reg3_reg[1]/NET0131  & ~n3369 ;
  assign n3371 = n333 & ~n747 ;
  assign n3394 = ~n3370 & ~n3371 ;
  assign n3395 = ~n3393 & n3394 ;
  assign n3396 = n292 & ~n3395 ;
  assign n3397 = ~n3367 & ~n3396 ;
  assign n3398 = \state_reg[0]/NET0131  & ~n3397 ;
  assign n3399 = ~n3366 & ~n3398 ;
  assign n3400 = \reg3_reg[2]/NET0131  & ~n1471 ;
  assign n3401 = \reg3_reg[2]/NET0131  & n290 ;
  assign n3423 = \reg3_reg[2]/NET0131  & ~n308 ;
  assign n3424 = n418 & ~n425 ;
  assign n3425 = ~n418 & n425 ;
  assign n3426 = ~n3424 & ~n3425 ;
  assign n3427 = ~n341 & ~n3426 ;
  assign n3428 = n341 & n389 ;
  assign n3429 = ~n3427 & ~n3428 ;
  assign n3430 = n308 & n3429 ;
  assign n3431 = ~n3423 & ~n3430 ;
  assign n3432 = n588 & ~n3431 ;
  assign n3411 = ~n762 & ~n774 ;
  assign n3417 = ~n1082 & n3411 ;
  assign n3416 = n1082 & ~n3411 ;
  assign n3418 = n798 & ~n3416 ;
  assign n3419 = ~n3417 & n3418 ;
  assign n3408 = ~n761 & ~n883 ;
  assign n3409 = ~n884 & n907 ;
  assign n3410 = ~n3408 & n3409 ;
  assign n3413 = ~n857 & ~n3411 ;
  assign n3412 = n857 & n3411 ;
  assign n3414 = n881 & ~n3412 ;
  assign n3415 = ~n3413 & n3414 ;
  assign n3420 = ~n3410 & ~n3415 ;
  assign n3421 = ~n3419 & n3420 ;
  assign n3422 = n308 & ~n3421 ;
  assign n3433 = n308 & ~n761 ;
  assign n3434 = ~n3423 & ~n3433 ;
  assign n3435 = n910 & ~n3434 ;
  assign n3402 = n329 & ~n761 ;
  assign n3403 = ~n318 & n331 ;
  assign n3404 = ~n797 & ~n3403 ;
  assign n3405 = ~n308 & ~n3404 ;
  assign n3406 = ~n909 & ~n3405 ;
  assign n3407 = \reg3_reg[2]/NET0131  & ~n3406 ;
  assign n3436 = ~n3402 & ~n3407 ;
  assign n3437 = ~n3435 & n3436 ;
  assign n3438 = ~n3422 & n3437 ;
  assign n3439 = ~n3432 & n3438 ;
  assign n3440 = n292 & ~n3439 ;
  assign n3441 = ~n3401 & ~n3440 ;
  assign n3442 = \state_reg[0]/NET0131  & ~n3441 ;
  assign n3443 = ~n3400 & ~n3442 ;
  assign n3446 = n290 & n441 ;
  assign n3448 = ~n308 & n441 ;
  assign n3449 = ~n456 & n483 ;
  assign n3450 = ~n2309 & ~n3449 ;
  assign n3451 = ~n341 & ~n3450 ;
  assign n3452 = n341 & n454 ;
  assign n3453 = ~n3451 & ~n3452 ;
  assign n3454 = n308 & n3453 ;
  assign n3455 = ~n3448 & ~n3454 ;
  assign n3456 = n588 & ~n3455 ;
  assign n3457 = ~n839 & ~n840 ;
  assign n3464 = ~n2223 & n3457 ;
  assign n3465 = n2223 & ~n3457 ;
  assign n3466 = ~n3464 & ~n3465 ;
  assign n3467 = n308 & n3466 ;
  assign n3468 = ~n3448 & ~n3467 ;
  assign n3469 = n881 & ~n3468 ;
  assign n3458 = ~n2211 & n3457 ;
  assign n3459 = n2211 & ~n3457 ;
  assign n3460 = ~n3458 & ~n3459 ;
  assign n3461 = n308 & ~n3460 ;
  assign n3462 = ~n3448 & ~n3461 ;
  assign n3463 = n798 & ~n3462 ;
  assign n3470 = ~n715 & ~n887 ;
  assign n3471 = ~n888 & n907 ;
  assign n3472 = ~n3470 & n3471 ;
  assign n3473 = n308 & n3472 ;
  assign n3447 = n441 & ~n1424 ;
  assign n3474 = n333 & ~n715 ;
  assign n3475 = ~n3447 & ~n3474 ;
  assign n3476 = ~n3473 & n3475 ;
  assign n3477 = ~n3463 & n3476 ;
  assign n3478 = ~n3469 & n3477 ;
  assign n3479 = ~n3456 & n3478 ;
  assign n3480 = n292 & ~n3479 ;
  assign n3481 = ~n3446 & ~n3480 ;
  assign n3482 = \state_reg[0]/NET0131  & ~n3481 ;
  assign n3444 = \reg3_reg[6]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3445 = n260 & n441 ;
  assign n3483 = ~n3444 & ~n3445 ;
  assign n3484 = ~n3482 & n3483 ;
  assign n3487 = n290 & n460 ;
  assign n3489 = ~n308 & n460 ;
  assign n3496 = n308 & ~n3099 ;
  assign n3497 = ~n3489 & ~n3496 ;
  assign n3498 = n588 & ~n3497 ;
  assign n3493 = n308 & n3091 ;
  assign n3494 = ~n3489 & ~n3493 ;
  assign n3495 = n881 & ~n3494 ;
  assign n3490 = n308 & ~n3085 ;
  assign n3491 = ~n3489 & ~n3490 ;
  assign n3492 = n798 & ~n3491 ;
  assign n3499 = n308 & n3105 ;
  assign n3500 = ~n3489 & ~n3499 ;
  assign n3501 = n907 & ~n3500 ;
  assign n3488 = n333 & ~n705 ;
  assign n3502 = n460 & ~n912 ;
  assign n3503 = ~n3488 & ~n3502 ;
  assign n3504 = ~n3501 & n3503 ;
  assign n3505 = ~n3492 & n3504 ;
  assign n3506 = ~n3495 & n3505 ;
  assign n3507 = ~n3498 & n3506 ;
  assign n3508 = n292 & ~n3507 ;
  assign n3509 = ~n3487 & ~n3508 ;
  assign n3510 = \state_reg[0]/NET0131  & ~n3509 ;
  assign n3485 = \reg3_reg[8]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3486 = n260 & n460 ;
  assign n3511 = ~n3485 & ~n3486 ;
  assign n3512 = ~n3510 & n3511 ;
  assign n3515 = n290 & n469 ;
  assign n3517 = ~n308 & n469 ;
  assign n3518 = n486 & ~n513 ;
  assign n3519 = ~n486 & n513 ;
  assign n3520 = ~n3518 & ~n3519 ;
  assign n3521 = ~n341 & ~n3520 ;
  assign n3522 = n341 & n465 ;
  assign n3523 = ~n3521 & ~n3522 ;
  assign n3524 = n308 & n3523 ;
  assign n3525 = ~n3517 & ~n3524 ;
  assign n3526 = n588 & ~n3525 ;
  assign n3527 = ~n631 & ~n687 ;
  assign n3534 = n786 & n3527 ;
  assign n3535 = ~n786 & ~n3527 ;
  assign n3536 = ~n3534 & ~n3535 ;
  assign n3537 = n308 & ~n3536 ;
  assign n3538 = ~n3517 & ~n3537 ;
  assign n3539 = n798 & ~n3538 ;
  assign n3528 = n872 & n3527 ;
  assign n3529 = ~n872 & ~n3527 ;
  assign n3530 = ~n3528 & ~n3529 ;
  assign n3531 = n308 & n3530 ;
  assign n3532 = ~n3517 & ~n3531 ;
  assign n3533 = n881 & ~n3532 ;
  assign n3540 = ~n630 & ~n3104 ;
  assign n3541 = ~n891 & ~n3540 ;
  assign n3542 = n308 & n3541 ;
  assign n3543 = ~n3517 & ~n3542 ;
  assign n3544 = n907 & ~n3543 ;
  assign n3516 = n333 & ~n630 ;
  assign n3545 = n469 & ~n912 ;
  assign n3546 = ~n3516 & ~n3545 ;
  assign n3547 = ~n3544 & n3546 ;
  assign n3548 = ~n3533 & n3547 ;
  assign n3549 = ~n3539 & n3548 ;
  assign n3550 = ~n3526 & n3549 ;
  assign n3551 = n292 & ~n3550 ;
  assign n3552 = ~n3515 & ~n3551 ;
  assign n3553 = \state_reg[0]/NET0131  & ~n3552 ;
  assign n3513 = \reg3_reg[9]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3514 = n260 & n469 ;
  assign n3554 = ~n3513 & ~n3514 ;
  assign n3555 = ~n3553 & n3554 ;
  assign n3558 = n290 & n970 ;
  assign n3559 = ~n308 & n970 ;
  assign n3568 = n308 & ~n2857 ;
  assign n3569 = ~n3559 & ~n3568 ;
  assign n3570 = n588 & ~n3569 ;
  assign n3571 = n308 & ~n2838 ;
  assign n3572 = ~n3559 & ~n3571 ;
  assign n3573 = n881 & ~n3572 ;
  assign n3560 = n308 & ~n2869 ;
  assign n3561 = ~n3559 & ~n3560 ;
  assign n3562 = n798 & ~n3561 ;
  assign n3564 = n308 & n2844 ;
  assign n3565 = ~n3559 & ~n3564 ;
  assign n3566 = n907 & ~n3565 ;
  assign n3563 = n333 & n965 ;
  assign n3567 = ~n912 & n970 ;
  assign n3574 = ~n3563 & ~n3567 ;
  assign n3575 = ~n3566 & n3574 ;
  assign n3576 = ~n3562 & n3575 ;
  assign n3577 = ~n3573 & n3576 ;
  assign n3578 = ~n3570 & n3577 ;
  assign n3579 = n292 & ~n3578 ;
  assign n3580 = ~n3558 & ~n3579 ;
  assign n3581 = \state_reg[0]/NET0131  & ~n3580 ;
  assign n3556 = \reg3_reg[25]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3557 = n260 & n970 ;
  assign n3582 = ~n3556 & ~n3557 ;
  assign n3583 = ~n3581 & n3582 ;
  assign n3590 = \reg2_reg[3]/NET0131  & ~n1543 ;
  assign n3591 = n341 & ~n382 ;
  assign n3592 = n434 & ~n3424 ;
  assign n3593 = ~n341 & ~n436 ;
  assign n3594 = ~n3592 & n3593 ;
  assign n3595 = ~n3591 & ~n3594 ;
  assign n3596 = n1543 & ~n3595 ;
  assign n3597 = ~n3590 & ~n3596 ;
  assign n3598 = n588 & ~n3597 ;
  assign n3599 = ~n858 & ~n860 ;
  assign n3600 = ~n859 & ~n866 ;
  assign n3601 = n3599 & ~n3600 ;
  assign n3602 = ~n3599 & n3600 ;
  assign n3603 = ~n3601 & ~n3602 ;
  assign n3604 = n1543 & ~n3603 ;
  assign n3605 = ~n3590 & ~n3604 ;
  assign n3606 = n881 & ~n3605 ;
  assign n3607 = ~n764 & ~n774 ;
  assign n3608 = ~n3600 & n3607 ;
  assign n3609 = n3600 & ~n3607 ;
  assign n3610 = ~n3608 & ~n3609 ;
  assign n3611 = n1543 & n3610 ;
  assign n3612 = ~n3590 & ~n3611 ;
  assign n3613 = n798 & ~n3612 ;
  assign n3584 = ~n772 & n910 ;
  assign n3585 = ~n772 & ~n884 ;
  assign n3586 = ~n885 & n907 ;
  assign n3587 = ~n3585 & n3586 ;
  assign n3588 = ~n3584 & ~n3587 ;
  assign n3589 = n1543 & ~n3588 ;
  assign n3614 = ~\reg3_reg[3]/NET0131  & n329 ;
  assign n3615 = \reg2_reg[3]/NET0131  & ~n2046 ;
  assign n3616 = ~n3614 & ~n3615 ;
  assign n3617 = ~n3589 & n3616 ;
  assign n3618 = ~n3613 & n3617 ;
  assign n3619 = ~n3606 & n3618 ;
  assign n3620 = ~n3598 & n3619 ;
  assign n3621 = n292 & ~n3620 ;
  assign n3622 = \reg2_reg[3]/NET0131  & n290 ;
  assign n3623 = ~n3621 & ~n3622 ;
  assign n3624 = \state_reg[0]/NET0131  & ~n3623 ;
  assign n3625 = \reg2_reg[3]/NET0131  & ~n1471 ;
  assign n3626 = ~n3624 & ~n3625 ;
  assign n3630 = \reg0_reg[18]/NET0131  & ~n1444 ;
  assign n3631 = n1444 & ~n2790 ;
  assign n3632 = ~n3630 & ~n3631 ;
  assign n3633 = n881 & ~n3632 ;
  assign n3634 = n1444 & n2798 ;
  assign n3635 = ~n3630 & ~n3634 ;
  assign n3636 = n588 & ~n3635 ;
  assign n3627 = n910 & n1038 ;
  assign n3628 = n2809 & ~n3627 ;
  assign n3629 = n1444 & ~n3628 ;
  assign n3637 = \reg0_reg[18]/NET0131  & ~n3035 ;
  assign n3638 = ~n3629 & ~n3637 ;
  assign n3639 = ~n3636 & n3638 ;
  assign n3640 = ~n3633 & n3639 ;
  assign n3641 = n292 & ~n3640 ;
  assign n3642 = \reg0_reg[18]/NET0131  & n290 ;
  assign n3643 = ~n3641 & ~n3642 ;
  assign n3644 = \state_reg[0]/NET0131  & ~n3643 ;
  assign n3645 = \reg0_reg[18]/NET0131  & ~n1471 ;
  assign n3646 = ~n3644 & ~n3645 ;
  assign n3647 = \reg0_reg[25]/NET0131  & ~n1471 ;
  assign n3648 = \reg0_reg[25]/NET0131  & n290 ;
  assign n3649 = \reg0_reg[25]/NET0131  & ~n1444 ;
  assign n3658 = n1444 & ~n2857 ;
  assign n3659 = ~n3649 & ~n3658 ;
  assign n3660 = n588 & ~n3659 ;
  assign n3661 = n1444 & ~n2838 ;
  assign n3662 = ~n3649 & ~n3661 ;
  assign n3663 = n881 & ~n3662 ;
  assign n3650 = n1444 & ~n2869 ;
  assign n3651 = ~n3649 & ~n3650 ;
  assign n3652 = n798 & ~n3651 ;
  assign n3654 = n1444 & n2844 ;
  assign n3655 = ~n3649 & ~n3654 ;
  assign n3656 = n907 & ~n3655 ;
  assign n3653 = \reg0_reg[25]/NET0131  & ~n1459 ;
  assign n3657 = n1444 & n2849 ;
  assign n3664 = ~n3653 & ~n3657 ;
  assign n3665 = ~n3656 & n3664 ;
  assign n3666 = ~n3652 & n3665 ;
  assign n3667 = ~n3663 & n3666 ;
  assign n3668 = ~n3660 & n3667 ;
  assign n3669 = n292 & ~n3668 ;
  assign n3670 = ~n3648 & ~n3669 ;
  assign n3671 = \state_reg[0]/NET0131  & ~n3670 ;
  assign n3672 = ~n3647 & ~n3671 ;
  assign n3676 = \reg0_reg[3]/NET0131  & ~n1444 ;
  assign n3677 = n1444 & ~n3595 ;
  assign n3678 = ~n3676 & ~n3677 ;
  assign n3679 = n588 & ~n3678 ;
  assign n3680 = n1444 & ~n3603 ;
  assign n3681 = ~n3676 & ~n3680 ;
  assign n3682 = n881 & ~n3681 ;
  assign n3673 = n798 & n3610 ;
  assign n3674 = n3588 & ~n3673 ;
  assign n3675 = n1444 & ~n3674 ;
  assign n3683 = \reg0_reg[3]/NET0131  & ~n3035 ;
  assign n3684 = ~n3675 & ~n3683 ;
  assign n3685 = ~n3682 & n3684 ;
  assign n3686 = ~n3679 & n3685 ;
  assign n3687 = n292 & ~n3686 ;
  assign n3688 = \reg0_reg[3]/NET0131  & n290 ;
  assign n3689 = ~n3687 & ~n3688 ;
  assign n3690 = \state_reg[0]/NET0131  & ~n3689 ;
  assign n3691 = \reg0_reg[3]/NET0131  & ~n1471 ;
  assign n3692 = ~n3690 & ~n3691 ;
  assign n3705 = \reg1_reg[10]/NET0131  & ~n1497 ;
  assign n3706 = n504 & ~n3518 ;
  assign n3707 = ~n1658 & ~n3706 ;
  assign n3708 = ~n341 & ~n3707 ;
  assign n3709 = n341 & n474 ;
  assign n3710 = ~n3708 & ~n3709 ;
  assign n3711 = n1497 & n3710 ;
  assign n3712 = ~n3705 & ~n3711 ;
  assign n3713 = n588 & ~n3712 ;
  assign n3697 = ~n820 & ~n821 ;
  assign n3714 = ~n2228 & n3697 ;
  assign n3715 = n2228 & ~n3697 ;
  assign n3716 = ~n3714 & ~n3715 ;
  assign n3717 = n1497 & n3716 ;
  assign n3718 = ~n3705 & ~n3717 ;
  assign n3719 = n881 & ~n3718 ;
  assign n3699 = n2468 & n3697 ;
  assign n3698 = ~n2468 & ~n3697 ;
  assign n3700 = n798 & ~n3698 ;
  assign n3701 = ~n3699 & n3700 ;
  assign n3693 = ~n622 & ~n891 ;
  assign n3694 = ~n1673 & ~n3693 ;
  assign n3695 = n907 & n3694 ;
  assign n3696 = ~n622 & n910 ;
  assign n3702 = ~n3695 & ~n3696 ;
  assign n3703 = ~n3701 & n3702 ;
  assign n3704 = n1497 & ~n3703 ;
  assign n3720 = \reg1_reg[10]/NET0131  & ~n2018 ;
  assign n3721 = ~n3704 & ~n3720 ;
  assign n3722 = ~n3719 & n3721 ;
  assign n3723 = ~n3713 & n3722 ;
  assign n3724 = n292 & ~n3723 ;
  assign n3725 = \reg1_reg[10]/NET0131  & n290 ;
  assign n3726 = ~n3724 & ~n3725 ;
  assign n3727 = \state_reg[0]/NET0131  & ~n3726 ;
  assign n3728 = \reg1_reg[10]/NET0131  & ~n1471 ;
  assign n3729 = ~n3727 & ~n3728 ;
  assign n3730 = \reg1_reg[25]/NET0131  & ~n1471 ;
  assign n3731 = \reg1_reg[25]/NET0131  & n290 ;
  assign n3732 = \reg1_reg[25]/NET0131  & ~n1497 ;
  assign n3741 = n1497 & ~n2857 ;
  assign n3742 = ~n3732 & ~n3741 ;
  assign n3743 = n588 & ~n3742 ;
  assign n3744 = n1497 & ~n2838 ;
  assign n3745 = ~n3732 & ~n3744 ;
  assign n3746 = n881 & ~n3745 ;
  assign n3733 = n1497 & ~n2869 ;
  assign n3734 = ~n3732 & ~n3733 ;
  assign n3735 = n798 & ~n3734 ;
  assign n3737 = n1497 & n2844 ;
  assign n3738 = ~n3732 & ~n3737 ;
  assign n3739 = n907 & ~n3738 ;
  assign n3736 = \reg1_reg[25]/NET0131  & ~n1529 ;
  assign n3740 = n1497 & n2849 ;
  assign n3747 = ~n3736 & ~n3740 ;
  assign n3748 = ~n3739 & n3747 ;
  assign n3749 = ~n3735 & n3748 ;
  assign n3750 = ~n3746 & n3749 ;
  assign n3751 = ~n3743 & n3750 ;
  assign n3752 = n292 & ~n3751 ;
  assign n3753 = ~n3731 & ~n3752 ;
  assign n3754 = \state_reg[0]/NET0131  & ~n3753 ;
  assign n3755 = ~n3730 & ~n3754 ;
  assign n3757 = \reg1_reg[3]/NET0131  & ~n1497 ;
  assign n3758 = n1497 & ~n3595 ;
  assign n3759 = ~n3757 & ~n3758 ;
  assign n3760 = n588 & ~n3759 ;
  assign n3761 = n1497 & ~n3603 ;
  assign n3762 = ~n3757 & ~n3761 ;
  assign n3763 = n881 & ~n3762 ;
  assign n3756 = n1497 & ~n3674 ;
  assign n3764 = \reg1_reg[3]/NET0131  & ~n2018 ;
  assign n3765 = ~n3756 & ~n3764 ;
  assign n3766 = ~n3763 & n3765 ;
  assign n3767 = ~n3760 & n3766 ;
  assign n3768 = n292 & ~n3767 ;
  assign n3769 = \reg1_reg[3]/NET0131  & n290 ;
  assign n3770 = ~n3768 & ~n3769 ;
  assign n3771 = \state_reg[0]/NET0131  & ~n3770 ;
  assign n3772 = \reg1_reg[3]/NET0131  & ~n1471 ;
  assign n3773 = ~n3771 & ~n3772 ;
  assign n3774 = \reg2_reg[10]/NET0131  & ~n1471 ;
  assign n3775 = \reg2_reg[10]/NET0131  & n290 ;
  assign n3777 = \reg2_reg[10]/NET0131  & ~n1543 ;
  assign n3778 = n1543 & n3710 ;
  assign n3779 = ~n3777 & ~n3778 ;
  assign n3780 = n588 & ~n3779 ;
  assign n3782 = n1543 & n3716 ;
  assign n3783 = ~n3777 & ~n3782 ;
  assign n3784 = n881 & ~n3783 ;
  assign n3776 = n1543 & ~n3703 ;
  assign n3781 = n329 & n508 ;
  assign n3785 = ~n1543 & ~n2811 ;
  assign n3786 = n1560 & ~n3785 ;
  assign n3787 = \reg2_reg[10]/NET0131  & ~n3786 ;
  assign n3788 = ~n3781 & ~n3787 ;
  assign n3789 = ~n3776 & n3788 ;
  assign n3790 = ~n3784 & n3789 ;
  assign n3791 = ~n3780 & n3790 ;
  assign n3792 = n292 & ~n3791 ;
  assign n3793 = ~n3775 & ~n3792 ;
  assign n3794 = \state_reg[0]/NET0131  & ~n3793 ;
  assign n3795 = ~n3774 & ~n3794 ;
  assign n3797 = \reg0_reg[10]/NET0131  & ~n1444 ;
  assign n3798 = n1444 & n3710 ;
  assign n3799 = ~n3797 & ~n3798 ;
  assign n3800 = n588 & ~n3799 ;
  assign n3801 = n1444 & n3716 ;
  assign n3802 = ~n3797 & ~n3801 ;
  assign n3803 = n881 & ~n3802 ;
  assign n3796 = \reg0_reg[10]/NET0131  & ~n3035 ;
  assign n3804 = n1444 & ~n3703 ;
  assign n3805 = ~n3796 & ~n3804 ;
  assign n3806 = ~n3803 & n3805 ;
  assign n3807 = ~n3800 & n3806 ;
  assign n3808 = n292 & ~n3807 ;
  assign n3809 = \reg0_reg[10]/NET0131  & n290 ;
  assign n3810 = ~n3808 & ~n3809 ;
  assign n3811 = \state_reg[0]/NET0131  & ~n3810 ;
  assign n3812 = \reg0_reg[10]/NET0131  & ~n1471 ;
  assign n3813 = ~n3811 & ~n3812 ;
  assign n3814 = \reg2_reg[18]/NET0131  & ~n1471 ;
  assign n3815 = \reg2_reg[18]/NET0131  & n290 ;
  assign n3817 = \reg2_reg[18]/NET0131  & ~n1543 ;
  assign n3818 = n1543 & ~n2790 ;
  assign n3819 = ~n3817 & ~n3818 ;
  assign n3820 = n881 & ~n3819 ;
  assign n3822 = n1543 & n2798 ;
  assign n3823 = ~n3817 & ~n3822 ;
  assign n3824 = n588 & ~n3823 ;
  assign n3816 = n1543 & ~n3628 ;
  assign n3821 = n329 & n572 ;
  assign n3825 = \reg2_reg[18]/NET0131  & ~n3786 ;
  assign n3826 = ~n3821 & ~n3825 ;
  assign n3827 = ~n3816 & n3826 ;
  assign n3828 = ~n3824 & n3827 ;
  assign n3829 = ~n3820 & n3828 ;
  assign n3830 = n292 & ~n3829 ;
  assign n3831 = ~n3815 & ~n3830 ;
  assign n3832 = \state_reg[0]/NET0131  & ~n3831 ;
  assign n3833 = ~n3814 & ~n3832 ;
  assign n3834 = n290 & n427 ;
  assign n3849 = ~n740 & ~n778 ;
  assign n3855 = n1086 & ~n3849 ;
  assign n3854 = ~n1086 & n3849 ;
  assign n3856 = n798 & ~n3854 ;
  assign n3857 = ~n3855 & n3856 ;
  assign n3846 = ~n739 & ~n885 ;
  assign n3847 = ~n886 & n907 ;
  assign n3848 = ~n3846 & n3847 ;
  assign n3851 = ~n1168 & ~n3849 ;
  assign n3850 = n1168 & n3849 ;
  assign n3852 = n881 & ~n3850 ;
  assign n3853 = ~n3851 & n3852 ;
  assign n3858 = ~n3848 & ~n3853 ;
  assign n3859 = ~n3857 & n3858 ;
  assign n3860 = n308 & ~n3859 ;
  assign n3836 = ~n436 & n454 ;
  assign n3837 = n436 & ~n454 ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = ~n341 & ~n3838 ;
  assign n3840 = n341 & n425 ;
  assign n3841 = ~n3839 & ~n3840 ;
  assign n3842 = n308 & ~n3841 ;
  assign n3843 = ~n308 & ~n427 ;
  assign n3844 = n588 & ~n3843 ;
  assign n3845 = ~n3842 & n3844 ;
  assign n3835 = n333 & ~n739 ;
  assign n3861 = ~n308 & n797 ;
  assign n3862 = n1424 & ~n3861 ;
  assign n3863 = n427 & ~n3862 ;
  assign n3864 = ~n3835 & ~n3863 ;
  assign n3865 = ~n3845 & n3864 ;
  assign n3866 = ~n3860 & n3865 ;
  assign n3867 = n292 & ~n3866 ;
  assign n3868 = ~n3834 & ~n3867 ;
  assign n3869 = \state_reg[0]/NET0131  & ~n3868 ;
  assign n3870 = \state_reg[0]/NET0131  & ~n427 ;
  assign n3871 = ~\reg3_reg[4]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3872 = ~n3870 & ~n3871 ;
  assign n3873 = ~n1471 & n3872 ;
  assign n3874 = ~n3869 & ~n3873 ;
  assign n3875 = \reg2_reg[6]/NET0131  & ~n1471 ;
  assign n3876 = \reg2_reg[6]/NET0131  & n290 ;
  assign n3878 = \reg2_reg[6]/NET0131  & ~n1543 ;
  assign n3879 = n1543 & n3453 ;
  assign n3880 = ~n3878 & ~n3879 ;
  assign n3881 = n588 & ~n3880 ;
  assign n3885 = n1543 & n3466 ;
  assign n3886 = ~n3878 & ~n3885 ;
  assign n3887 = n881 & ~n3886 ;
  assign n3882 = n1543 & ~n3460 ;
  assign n3883 = ~n3878 & ~n3882 ;
  assign n3884 = n798 & ~n3883 ;
  assign n3889 = ~n715 & n910 ;
  assign n3890 = ~n3472 & ~n3889 ;
  assign n3891 = n1543 & ~n3890 ;
  assign n3877 = \reg2_reg[6]/NET0131  & ~n1585 ;
  assign n3888 = n329 & n441 ;
  assign n3892 = ~n3877 & ~n3888 ;
  assign n3893 = ~n3891 & n3892 ;
  assign n3894 = ~n3884 & n3893 ;
  assign n3895 = ~n3887 & n3894 ;
  assign n3896 = ~n3881 & n3895 ;
  assign n3897 = n292 & ~n3896 ;
  assign n3898 = ~n3876 & ~n3897 ;
  assign n3899 = \state_reg[0]/NET0131  & ~n3898 ;
  assign n3900 = ~n3875 & ~n3899 ;
  assign n3901 = \reg2_reg[8]/NET0131  & ~n1471 ;
  assign n3902 = \reg2_reg[8]/NET0131  & n290 ;
  assign n3904 = \reg2_reg[8]/NET0131  & ~n1543 ;
  assign n3911 = n1543 & ~n3099 ;
  assign n3912 = ~n3904 & ~n3911 ;
  assign n3913 = n588 & ~n3912 ;
  assign n3908 = n1543 & n3091 ;
  assign n3909 = ~n3904 & ~n3908 ;
  assign n3910 = n881 & ~n3909 ;
  assign n3905 = n1543 & ~n3085 ;
  assign n3906 = ~n3904 & ~n3905 ;
  assign n3907 = n798 & ~n3906 ;
  assign n3914 = n1543 & n3105 ;
  assign n3915 = ~n3904 & ~n3914 ;
  assign n3916 = n907 & ~n3915 ;
  assign n3918 = \reg2_reg[8]/NET0131  & ~n1560 ;
  assign n3903 = n1543 & n3109 ;
  assign n3917 = n329 & n460 ;
  assign n3919 = ~n3903 & ~n3917 ;
  assign n3920 = ~n3918 & n3919 ;
  assign n3921 = ~n3916 & n3920 ;
  assign n3922 = ~n3907 & n3921 ;
  assign n3923 = ~n3910 & n3922 ;
  assign n3924 = ~n3913 & n3923 ;
  assign n3925 = n292 & ~n3924 ;
  assign n3926 = ~n3902 & ~n3925 ;
  assign n3927 = \state_reg[0]/NET0131  & ~n3926 ;
  assign n3928 = ~n3901 & ~n3927 ;
  assign n3929 = \reg0_reg[17]/NET0131  & ~n1471 ;
  assign n3930 = \reg0_reg[17]/NET0131  & n290 ;
  assign n3933 = \reg0_reg[17]/NET0131  & ~n1444 ;
  assign n3934 = n583 & n1444 ;
  assign n3935 = ~n3933 & ~n3934 ;
  assign n3936 = n588 & ~n3935 ;
  assign n3937 = ~n792 & n1444 ;
  assign n3938 = ~n3933 & ~n3937 ;
  assign n3939 = n798 & ~n3938 ;
  assign n3931 = n356 & n910 ;
  assign n3932 = n1444 & n3931 ;
  assign n3946 = \reg0_reg[17]/NET0131  & ~n1459 ;
  assign n3947 = ~n3932 & ~n3946 ;
  assign n3948 = ~n3939 & n3947 ;
  assign n3940 = n878 & n1444 ;
  assign n3941 = ~n3933 & ~n3940 ;
  assign n3942 = n881 & ~n3941 ;
  assign n3943 = n904 & n1444 ;
  assign n3944 = ~n3933 & ~n3943 ;
  assign n3945 = n907 & ~n3944 ;
  assign n3949 = ~n3942 & ~n3945 ;
  assign n3950 = n3948 & n3949 ;
  assign n3951 = ~n3936 & n3950 ;
  assign n3952 = n292 & ~n3951 ;
  assign n3953 = ~n3930 & ~n3952 ;
  assign n3954 = \state_reg[0]/NET0131  & ~n3953 ;
  assign n3955 = ~n3929 & ~n3954 ;
  assign n3956 = ~n747 & n910 ;
  assign n3957 = n3392 & ~n3956 ;
  assign n3958 = n3048 & ~n3957 ;
  assign n3959 = ~n588 & ~n881 ;
  assign n3960 = ~n797 & n3959 ;
  assign n3961 = ~n1444 & ~n3960 ;
  assign n3962 = n2389 & ~n3961 ;
  assign n3963 = n1911 & n3962 ;
  assign n3964 = \reg0_reg[1]/NET0131  & ~n3963 ;
  assign n3965 = ~n3958 & ~n3964 ;
  assign n3966 = \reg0_reg[21]/NET0131  & ~n1471 ;
  assign n3967 = \reg0_reg[21]/NET0131  & n290 ;
  assign n3968 = ~n332 & ~n909 ;
  assign n3969 = ~n1444 & n3968 ;
  assign n3970 = n1459 & ~n3969 ;
  assign n3971 = \reg0_reg[21]/NET0131  & ~n3970 ;
  assign n3972 = n910 & n1004 ;
  assign n3982 = n1004 & ~n2371 ;
  assign n3983 = n907 & ~n2913 ;
  assign n3984 = ~n3982 & n3983 ;
  assign n3973 = ~n1201 & ~n1217 ;
  assign n3975 = ~n2116 & n3973 ;
  assign n3974 = n2116 & ~n3973 ;
  assign n3976 = n881 & ~n3974 ;
  assign n3977 = ~n3975 & n3976 ;
  assign n3979 = ~n2148 & ~n3973 ;
  assign n3978 = n2148 & n3973 ;
  assign n3980 = n798 & ~n3978 ;
  assign n3981 = ~n3979 & n3980 ;
  assign n3985 = ~n3977 & ~n3981 ;
  assign n3986 = ~n3984 & n3985 ;
  assign n3987 = ~n3972 & n3986 ;
  assign n3988 = n1001 & ~n2362 ;
  assign n3989 = ~n2907 & ~n3988 ;
  assign n3990 = ~n341 & ~n3989 ;
  assign n3991 = n341 & n1026 ;
  assign n3992 = ~n3990 & ~n3991 ;
  assign n3993 = n588 & n3992 ;
  assign n3994 = n3987 & ~n3993 ;
  assign n3995 = n1444 & ~n3994 ;
  assign n3996 = ~n3971 & ~n3995 ;
  assign n3997 = n292 & ~n3996 ;
  assign n3998 = ~n3967 & ~n3997 ;
  assign n3999 = \state_reg[0]/NET0131  & ~n3998 ;
  assign n4000 = ~n3966 & ~n3999 ;
  assign n4001 = n2389 & n3970 ;
  assign n4002 = \reg0_reg[2]/NET0131  & ~n4001 ;
  assign n4003 = ~n761 & n910 ;
  assign n4004 = n3421 & ~n4003 ;
  assign n4005 = n588 & n3429 ;
  assign n4006 = n4004 & ~n4005 ;
  assign n4007 = n2389 & ~n4006 ;
  assign n4008 = n1444 & n4007 ;
  assign n4009 = ~n4002 & ~n4008 ;
  assign n4010 = \reg0_reg[4]/NET0131  & ~n4001 ;
  assign n4012 = n588 & n3841 ;
  assign n4011 = ~n739 & n910 ;
  assign n4013 = n3859 & ~n4011 ;
  assign n4014 = ~n4012 & n4013 ;
  assign n4015 = n2389 & ~n4014 ;
  assign n4016 = n1444 & n4015 ;
  assign n4017 = ~n4010 & ~n4016 ;
  assign n4018 = \reg0_reg[5]/NET0131  & ~n1471 ;
  assign n4019 = \reg0_reg[5]/NET0131  & n290 ;
  assign n4021 = \reg0_reg[5]/NET0131  & ~n1444 ;
  assign n4022 = n341 & ~n434 ;
  assign n4023 = n445 & ~n3837 ;
  assign n4024 = ~n341 & ~n456 ;
  assign n4025 = ~n4023 & n4024 ;
  assign n4026 = ~n4022 & ~n4025 ;
  assign n4027 = n1444 & ~n4026 ;
  assign n4028 = ~n4021 & ~n4027 ;
  assign n4029 = n588 & ~n4028 ;
  assign n4030 = ~n724 & ~n782 ;
  assign n4037 = n781 & n4030 ;
  assign n4038 = ~n781 & ~n4030 ;
  assign n4039 = ~n4037 & ~n4038 ;
  assign n4040 = n1444 & n4039 ;
  assign n4041 = ~n4021 & ~n4040 ;
  assign n4042 = n798 & ~n4041 ;
  assign n4031 = n869 & n4030 ;
  assign n4032 = ~n869 & ~n4030 ;
  assign n4033 = ~n4031 & ~n4032 ;
  assign n4034 = n1444 & n4033 ;
  assign n4035 = ~n4021 & ~n4034 ;
  assign n4036 = n881 & ~n4035 ;
  assign n4020 = \reg0_reg[5]/NET0131  & ~n1911 ;
  assign n4043 = ~n723 & n910 ;
  assign n4044 = ~n723 & ~n886 ;
  assign n4045 = ~n887 & n907 ;
  assign n4046 = ~n4044 & n4045 ;
  assign n4047 = ~n4043 & ~n4046 ;
  assign n4048 = n1444 & ~n4047 ;
  assign n4049 = ~n4020 & ~n4048 ;
  assign n4050 = ~n4036 & n4049 ;
  assign n4051 = ~n4042 & n4050 ;
  assign n4052 = ~n4029 & n4051 ;
  assign n4053 = n292 & ~n4052 ;
  assign n4054 = ~n4019 & ~n4053 ;
  assign n4055 = \state_reg[0]/NET0131  & ~n4054 ;
  assign n4056 = ~n4018 & ~n4055 ;
  assign n4057 = \reg0_reg[6]/NET0131  & ~n1471 ;
  assign n4058 = \reg0_reg[6]/NET0131  & n290 ;
  assign n4060 = \reg0_reg[6]/NET0131  & ~n1444 ;
  assign n4061 = n1444 & n3453 ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = n588 & ~n4062 ;
  assign n4067 = n1444 & n3466 ;
  assign n4068 = ~n4060 & ~n4067 ;
  assign n4069 = n881 & ~n4068 ;
  assign n4064 = n1444 & ~n3460 ;
  assign n4065 = ~n4060 & ~n4064 ;
  assign n4066 = n798 & ~n4065 ;
  assign n4059 = \reg0_reg[6]/NET0131  & ~n1911 ;
  assign n4070 = n1444 & ~n3890 ;
  assign n4071 = ~n4059 & ~n4070 ;
  assign n4072 = ~n4066 & n4071 ;
  assign n4073 = ~n4069 & n4072 ;
  assign n4074 = ~n4063 & n4073 ;
  assign n4075 = n292 & ~n4074 ;
  assign n4076 = ~n4058 & ~n4075 ;
  assign n4077 = \state_reg[0]/NET0131  & ~n4076 ;
  assign n4078 = ~n4057 & ~n4077 ;
  assign n4079 = \reg0_reg[9]/NET0131  & ~n1471 ;
  assign n4080 = \reg0_reg[9]/NET0131  & n290 ;
  assign n4083 = \reg0_reg[9]/NET0131  & ~n1444 ;
  assign n4084 = n1444 & n3523 ;
  assign n4085 = ~n4083 & ~n4084 ;
  assign n4086 = n588 & ~n4085 ;
  assign n4090 = n1444 & ~n3536 ;
  assign n4091 = ~n4083 & ~n4090 ;
  assign n4092 = n798 & ~n4091 ;
  assign n4087 = n1444 & n3530 ;
  assign n4088 = ~n4083 & ~n4087 ;
  assign n4089 = n881 & ~n4088 ;
  assign n4093 = n1444 & n3541 ;
  assign n4094 = ~n4083 & ~n4093 ;
  assign n4095 = n907 & ~n4094 ;
  assign n4081 = ~n630 & n910 ;
  assign n4082 = n1444 & n4081 ;
  assign n4096 = \reg0_reg[9]/NET0131  & ~n1459 ;
  assign n4097 = ~n4082 & ~n4096 ;
  assign n4098 = ~n4095 & n4097 ;
  assign n4099 = ~n4089 & n4098 ;
  assign n4100 = ~n4092 & n4099 ;
  assign n4101 = ~n4086 & n4100 ;
  assign n4102 = n292 & ~n4101 ;
  assign n4103 = ~n4080 & ~n4102 ;
  assign n4104 = \state_reg[0]/NET0131  & ~n4103 ;
  assign n4105 = ~n4079 & ~n4104 ;
  assign n4106 = \reg1_reg[17]/NET0131  & ~n1471 ;
  assign n4107 = \reg1_reg[17]/NET0131  & n290 ;
  assign n4109 = \reg1_reg[17]/NET0131  & ~n1497 ;
  assign n4110 = n583 & n1497 ;
  assign n4111 = ~n4109 & ~n4110 ;
  assign n4112 = n588 & ~n4111 ;
  assign n4113 = ~n792 & n1497 ;
  assign n4114 = ~n4109 & ~n4113 ;
  assign n4115 = n798 & ~n4114 ;
  assign n4108 = n1497 & n3931 ;
  assign n4122 = \reg1_reg[17]/NET0131  & ~n1529 ;
  assign n4123 = ~n4108 & ~n4122 ;
  assign n4124 = ~n4115 & n4123 ;
  assign n4116 = n878 & n1497 ;
  assign n4117 = ~n4109 & ~n4116 ;
  assign n4118 = n881 & ~n4117 ;
  assign n4119 = n904 & n1497 ;
  assign n4120 = ~n4109 & ~n4119 ;
  assign n4121 = n907 & ~n4120 ;
  assign n4125 = ~n4118 & ~n4121 ;
  assign n4126 = n4124 & n4125 ;
  assign n4127 = ~n4112 & n4126 ;
  assign n4128 = n292 & ~n4127 ;
  assign n4129 = ~n4107 & ~n4128 ;
  assign n4130 = \state_reg[0]/NET0131  & ~n4129 ;
  assign n4131 = ~n4106 & ~n4130 ;
  assign n4132 = n3212 & ~n3957 ;
  assign n4133 = ~n1497 & ~n3960 ;
  assign n4134 = n1507 & n2389 ;
  assign n4135 = ~n4133 & n4134 ;
  assign n4136 = \reg1_reg[1]/NET0131  & ~n4135 ;
  assign n4137 = ~n4132 & ~n4136 ;
  assign n4138 = ~n1497 & n3968 ;
  assign n4139 = n1529 & ~n4138 ;
  assign n4140 = n2389 & n4139 ;
  assign n4141 = \reg1_reg[2]/NET0131  & ~n4140 ;
  assign n4142 = n1497 & n4007 ;
  assign n4143 = ~n4141 & ~n4142 ;
  assign n4144 = ~n1497 & ~n2719 ;
  assign n4145 = n2389 & ~n4144 ;
  assign n4146 = n1531 & n4145 ;
  assign n4147 = \reg1_reg[4]/NET0131  & ~n4146 ;
  assign n4148 = n1497 & n4015 ;
  assign n4149 = ~n4147 & ~n4148 ;
  assign n4150 = \reg1_reg[5]/NET0131  & ~n1471 ;
  assign n4151 = \reg1_reg[5]/NET0131  & n290 ;
  assign n4153 = \reg1_reg[5]/NET0131  & ~n1497 ;
  assign n4154 = n1497 & ~n4026 ;
  assign n4155 = ~n4153 & ~n4154 ;
  assign n4156 = n588 & ~n4155 ;
  assign n4160 = n1497 & n4039 ;
  assign n4161 = ~n4153 & ~n4160 ;
  assign n4162 = n798 & ~n4161 ;
  assign n4157 = n1497 & n4033 ;
  assign n4158 = ~n4153 & ~n4157 ;
  assign n4159 = n881 & ~n4158 ;
  assign n4152 = \reg1_reg[5]/NET0131  & ~n1531 ;
  assign n4163 = n1497 & ~n4047 ;
  assign n4164 = ~n4152 & ~n4163 ;
  assign n4165 = ~n4159 & n4164 ;
  assign n4166 = ~n4162 & n4165 ;
  assign n4167 = ~n4156 & n4166 ;
  assign n4168 = n292 & ~n4167 ;
  assign n4169 = ~n4151 & ~n4168 ;
  assign n4170 = \state_reg[0]/NET0131  & ~n4169 ;
  assign n4171 = ~n4150 & ~n4170 ;
  assign n4172 = \reg1_reg[6]/NET0131  & ~n1471 ;
  assign n4173 = \reg1_reg[6]/NET0131  & n290 ;
  assign n4175 = \reg1_reg[6]/NET0131  & ~n1497 ;
  assign n4176 = n1497 & n3453 ;
  assign n4177 = ~n4175 & ~n4176 ;
  assign n4178 = n588 & ~n4177 ;
  assign n4182 = n1497 & n3466 ;
  assign n4183 = ~n4175 & ~n4182 ;
  assign n4184 = n881 & ~n4183 ;
  assign n4179 = n1497 & ~n3460 ;
  assign n4180 = ~n4175 & ~n4179 ;
  assign n4181 = n798 & ~n4180 ;
  assign n4174 = \reg1_reg[6]/NET0131  & ~n1531 ;
  assign n4185 = n1497 & ~n3890 ;
  assign n4186 = ~n4174 & ~n4185 ;
  assign n4187 = ~n4181 & n4186 ;
  assign n4188 = ~n4184 & n4187 ;
  assign n4189 = ~n4178 & n4188 ;
  assign n4190 = n292 & ~n4189 ;
  assign n4191 = ~n4173 & ~n4190 ;
  assign n4192 = \state_reg[0]/NET0131  & ~n4191 ;
  assign n4193 = ~n4172 & ~n4192 ;
  assign n4194 = \reg1_reg[8]/NET0131  & ~n1471 ;
  assign n4195 = \reg1_reg[8]/NET0131  & n290 ;
  assign n4197 = \reg1_reg[8]/NET0131  & ~n1497 ;
  assign n4204 = n1497 & ~n3099 ;
  assign n4205 = ~n4197 & ~n4204 ;
  assign n4206 = n588 & ~n4205 ;
  assign n4201 = n1497 & n3091 ;
  assign n4202 = ~n4197 & ~n4201 ;
  assign n4203 = n881 & ~n4202 ;
  assign n4198 = n1497 & ~n3085 ;
  assign n4199 = ~n4197 & ~n4198 ;
  assign n4200 = n798 & ~n4199 ;
  assign n4207 = n1497 & n3105 ;
  assign n4208 = ~n4197 & ~n4207 ;
  assign n4209 = n907 & ~n4208 ;
  assign n4196 = n1497 & n3109 ;
  assign n4210 = \reg1_reg[8]/NET0131  & ~n1529 ;
  assign n4211 = ~n4196 & ~n4210 ;
  assign n4212 = ~n4209 & n4211 ;
  assign n4213 = ~n4200 & n4212 ;
  assign n4214 = ~n4203 & n4213 ;
  assign n4215 = ~n4206 & n4214 ;
  assign n4216 = n292 & ~n4215 ;
  assign n4217 = ~n4195 & ~n4216 ;
  assign n4218 = \state_reg[0]/NET0131  & ~n4217 ;
  assign n4219 = ~n4194 & ~n4218 ;
  assign n4220 = \reg1_reg[9]/NET0131  & ~n1471 ;
  assign n4221 = \reg1_reg[9]/NET0131  & n290 ;
  assign n4223 = \reg1_reg[9]/NET0131  & ~n1497 ;
  assign n4224 = n1497 & n3523 ;
  assign n4225 = ~n4223 & ~n4224 ;
  assign n4226 = n588 & ~n4225 ;
  assign n4230 = n1497 & ~n3536 ;
  assign n4231 = ~n4223 & ~n4230 ;
  assign n4232 = n798 & ~n4231 ;
  assign n4227 = n1497 & n3530 ;
  assign n4228 = ~n4223 & ~n4227 ;
  assign n4229 = n881 & ~n4228 ;
  assign n4233 = n1497 & n3541 ;
  assign n4234 = ~n4223 & ~n4233 ;
  assign n4235 = n907 & ~n4234 ;
  assign n4222 = n1497 & n4081 ;
  assign n4236 = \reg1_reg[9]/NET0131  & ~n1529 ;
  assign n4237 = ~n4222 & ~n4236 ;
  assign n4238 = ~n4235 & n4237 ;
  assign n4239 = ~n4229 & n4238 ;
  assign n4240 = ~n4232 & n4239 ;
  assign n4241 = ~n4226 & n4240 ;
  assign n4242 = n292 & ~n4241 ;
  assign n4243 = ~n4221 & ~n4242 ;
  assign n4244 = \state_reg[0]/NET0131  & ~n4243 ;
  assign n4245 = ~n4220 & ~n4244 ;
  assign n4246 = \reg3_reg[0]/NET0131  & ~n1471 ;
  assign n4247 = \reg3_reg[0]/NET0131  & n290 ;
  assign n4248 = ~n751 & n1422 ;
  assign n4249 = n389 & ~n416 ;
  assign n4250 = ~n341 & ~n417 ;
  assign n4251 = ~n4249 & n4250 ;
  assign n4252 = n588 & n4251 ;
  assign n4253 = ~n4248 & ~n4252 ;
  assign n4254 = ~n396 & n751 ;
  assign n4255 = ~n752 & ~n4254 ;
  assign n4256 = n797 & ~n4255 ;
  assign n4257 = n4253 & ~n4256 ;
  assign n4258 = n308 & ~n4257 ;
  assign n4259 = n329 & ~n751 ;
  assign n4260 = ~n330 & ~n909 ;
  assign n4261 = \reg3_reg[0]/NET0131  & ~n4260 ;
  assign n4262 = ~n4259 & ~n4261 ;
  assign n4263 = ~n4258 & n4262 ;
  assign n4264 = n292 & ~n4263 ;
  assign n4265 = ~n4247 & ~n4264 ;
  assign n4266 = \state_reg[0]/NET0131  & ~n4265 ;
  assign n4267 = ~n4246 & ~n4266 ;
  assign n4269 = n290 & n1010 ;
  assign n4275 = n308 & ~n3992 ;
  assign n4274 = ~n308 & ~n1010 ;
  assign n4276 = n588 & ~n4274 ;
  assign n4277 = ~n4275 & n4276 ;
  assign n4271 = n308 & ~n3986 ;
  assign n4270 = n333 & n1004 ;
  assign n4272 = n912 & ~n3405 ;
  assign n4273 = n1010 & ~n4272 ;
  assign n4278 = ~n4270 & ~n4273 ;
  assign n4279 = ~n4271 & n4278 ;
  assign n4280 = ~n4277 & n4279 ;
  assign n4281 = n292 & ~n4280 ;
  assign n4282 = ~n4269 & ~n4281 ;
  assign n4283 = \state_reg[0]/NET0131  & ~n4282 ;
  assign n4268 = \reg3_reg[21]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n4284 = n260 & n1010 ;
  assign n4285 = ~n4268 & ~n4284 ;
  assign n4286 = ~n4283 & n4285 ;
  assign n4287 = \reg2_reg[4]/NET0131  & ~n1471 ;
  assign n4288 = \reg2_reg[4]/NET0131  & n290 ;
  assign n4290 = n1543 & ~n4014 ;
  assign n4289 = n329 & n427 ;
  assign n4291 = ~n1543 & ~n3959 ;
  assign n4292 = n3786 & ~n4291 ;
  assign n4293 = \reg2_reg[4]/NET0131  & ~n4292 ;
  assign n4294 = ~n4289 & ~n4293 ;
  assign n4295 = ~n4290 & n4294 ;
  assign n4296 = n292 & ~n4295 ;
  assign n4297 = ~n4288 & ~n4296 ;
  assign n4298 = \state_reg[0]/NET0131  & ~n4297 ;
  assign n4299 = ~n4287 & ~n4298 ;
  assign n4300 = \reg2_reg[5]/NET0131  & ~n1471 ;
  assign n4301 = \reg2_reg[5]/NET0131  & n290 ;
  assign n4303 = \reg2_reg[5]/NET0131  & ~n1543 ;
  assign n4304 = n1543 & ~n4026 ;
  assign n4305 = ~n4303 & ~n4304 ;
  assign n4306 = n588 & ~n4305 ;
  assign n4310 = n1543 & n4039 ;
  assign n4311 = ~n4303 & ~n4310 ;
  assign n4312 = n798 & ~n4311 ;
  assign n4307 = n1543 & n4033 ;
  assign n4308 = ~n4303 & ~n4307 ;
  assign n4309 = n881 & ~n4308 ;
  assign n4314 = n1543 & ~n4047 ;
  assign n4302 = \reg2_reg[5]/NET0131  & ~n1585 ;
  assign n4313 = n329 & n447 ;
  assign n4315 = ~n4302 & ~n4313 ;
  assign n4316 = ~n4314 & n4315 ;
  assign n4317 = ~n4309 & n4316 ;
  assign n4318 = ~n4312 & n4317 ;
  assign n4319 = ~n4306 & n4318 ;
  assign n4320 = n292 & ~n4319 ;
  assign n4321 = ~n4301 & ~n4320 ;
  assign n4322 = \state_reg[0]/NET0131  & ~n4321 ;
  assign n4323 = ~n4300 & ~n4322 ;
  assign n4324 = \reg2_reg[9]/NET0131  & ~n1471 ;
  assign n4325 = \reg2_reg[9]/NET0131  & n290 ;
  assign n4327 = \reg2_reg[9]/NET0131  & ~n1543 ;
  assign n4328 = n1543 & n3523 ;
  assign n4329 = ~n4327 & ~n4328 ;
  assign n4330 = n588 & ~n4329 ;
  assign n4334 = n1543 & n3530 ;
  assign n4335 = ~n4327 & ~n4334 ;
  assign n4336 = n881 & ~n4335 ;
  assign n4331 = n1543 & ~n3536 ;
  assign n4332 = ~n4327 & ~n4331 ;
  assign n4333 = n798 & ~n4332 ;
  assign n4337 = n1543 & n3541 ;
  assign n4338 = ~n4327 & ~n4337 ;
  assign n4339 = n907 & ~n4338 ;
  assign n4341 = \reg2_reg[9]/NET0131  & ~n1560 ;
  assign n4326 = n1543 & n4081 ;
  assign n4340 = n329 & n469 ;
  assign n4342 = ~n4326 & ~n4340 ;
  assign n4343 = ~n4341 & n4342 ;
  assign n4344 = ~n4339 & n4343 ;
  assign n4345 = ~n4333 & n4344 ;
  assign n4346 = ~n4336 & n4345 ;
  assign n4347 = ~n4330 & n4346 ;
  assign n4348 = n292 & ~n4347 ;
  assign n4349 = ~n4325 & ~n4348 ;
  assign n4350 = \state_reg[0]/NET0131  & ~n4349 ;
  assign n4351 = ~n4324 & ~n4350 ;
  assign n4352 = \reg1_reg[21]/NET0131  & ~n1471 ;
  assign n4353 = \reg1_reg[21]/NET0131  & n290 ;
  assign n4354 = \reg1_reg[21]/NET0131  & ~n4139 ;
  assign n4355 = n1497 & ~n3994 ;
  assign n4356 = ~n4354 & ~n4355 ;
  assign n4357 = n292 & ~n4356 ;
  assign n4358 = ~n4353 & ~n4357 ;
  assign n4359 = \state_reg[0]/NET0131  & ~n4358 ;
  assign n4360 = ~n4352 & ~n4359 ;
  assign n4361 = \reg2_reg[1]/NET0131  & ~n1471 ;
  assign n4362 = \reg2_reg[1]/NET0131  & n290 ;
  assign n4366 = n3391 & ~n3956 ;
  assign n4367 = n1543 & ~n4366 ;
  assign n4364 = n1560 & ~n2720 ;
  assign n4365 = \reg2_reg[1]/NET0131  & ~n4364 ;
  assign n4363 = \reg3_reg[1]/NET0131  & n329 ;
  assign n4369 = n1543 & ~n3373 ;
  assign n4368 = ~\reg2_reg[1]/NET0131  & ~n1543 ;
  assign n4370 = n907 & ~n4368 ;
  assign n4371 = ~n4369 & n4370 ;
  assign n4372 = ~n4363 & ~n4371 ;
  assign n4373 = ~n4365 & n4372 ;
  assign n4374 = ~n4367 & n4373 ;
  assign n4375 = n292 & ~n4374 ;
  assign n4376 = ~n4362 & ~n4375 ;
  assign n4377 = \state_reg[0]/NET0131  & ~n4376 ;
  assign n4378 = ~n4361 & ~n4377 ;
  assign n4379 = n3212 & ~n4257 ;
  assign n4380 = n1507 & n4145 ;
  assign n4381 = \reg1_reg[0]/NET0131  & ~n4380 ;
  assign n4382 = ~n4379 & ~n4381 ;
  assign n4383 = \reg1_reg[13]/NET0131  & ~n1471 ;
  assign n4384 = \reg1_reg[13]/NET0131  & n290 ;
  assign n4394 = ~n654 & n910 ;
  assign n4395 = ~n805 & ~n814 ;
  assign n4401 = n2108 & ~n4395 ;
  assign n4400 = ~n2108 & n4395 ;
  assign n4402 = n881 & ~n4400 ;
  assign n4403 = ~n4401 & n4402 ;
  assign n4397 = n2140 & n4395 ;
  assign n4396 = ~n2140 & ~n4395 ;
  assign n4398 = n798 & ~n4396 ;
  assign n4399 = ~n4397 & n4398 ;
  assign n4404 = ~n654 & ~n1719 ;
  assign n4405 = ~n895 & n907 ;
  assign n4406 = ~n4404 & n4405 ;
  assign n4407 = ~n4399 & ~n4406 ;
  assign n4408 = ~n4403 & n4407 ;
  assign n4409 = ~n4394 & n4408 ;
  assign n4410 = n1497 & ~n4409 ;
  assign n4385 = n546 & ~n1619 ;
  assign n4386 = ~n1620 & ~n4385 ;
  assign n4387 = ~n341 & ~n4386 ;
  assign n4388 = n341 & n495 ;
  assign n4389 = ~n4387 & ~n4388 ;
  assign n4390 = n1497 & ~n4389 ;
  assign n4391 = ~\reg1_reg[13]/NET0131  & ~n1497 ;
  assign n4392 = n588 & ~n4391 ;
  assign n4393 = ~n4390 & n4392 ;
  assign n4411 = ~n910 & n3404 ;
  assign n4412 = ~n1497 & ~n4411 ;
  assign n4413 = n1458 & ~n4412 ;
  assign n4414 = \reg1_reg[13]/NET0131  & ~n4413 ;
  assign n4415 = ~n4393 & ~n4414 ;
  assign n4416 = ~n4410 & n4415 ;
  assign n4417 = n292 & ~n4416 ;
  assign n4418 = ~n4384 & ~n4417 ;
  assign n4419 = \state_reg[0]/NET0131  & ~n4418 ;
  assign n4420 = ~n4383 & ~n4419 ;
  assign n4421 = n1444 & ~n4251 ;
  assign n4422 = n588 & ~n4421 ;
  assign n4424 = ~n319 & ~n4255 ;
  assign n4425 = n1444 & ~n4424 ;
  assign n4426 = ~n329 & ~n796 ;
  assign n4427 = ~n4425 & n4426 ;
  assign n4423 = \reg0_reg[0]/NET0131  & ~n1458 ;
  assign n4428 = n2389 & ~n4248 ;
  assign n4429 = ~n4423 & n4428 ;
  assign n4430 = ~n4427 & n4429 ;
  assign n4431 = ~n4422 & n4430 ;
  assign n4432 = ~\reg0_reg[0]/NET0131  & ~n3048 ;
  assign n4433 = ~n4431 & ~n4432 ;
  assign n4434 = n2389 & n3332 ;
  assign n4435 = \reg2_reg[0]/NET0131  & ~n4434 ;
  assign n4436 = n1543 & ~n4253 ;
  assign n4437 = \reg3_reg[0]/NET0131  & n329 ;
  assign n4439 = n1543 & n4255 ;
  assign n4438 = ~\reg2_reg[0]/NET0131  & ~n1543 ;
  assign n4440 = n797 & ~n4438 ;
  assign n4441 = ~n4439 & n4440 ;
  assign n4442 = ~n4437 & ~n4441 ;
  assign n4443 = ~n4436 & n4442 ;
  assign n4444 = n2389 & ~n4443 ;
  assign n4445 = ~n4435 & ~n4444 ;
  assign n4446 = \reg2_reg[13]/NET0131  & ~n1471 ;
  assign n4447 = \reg2_reg[13]/NET0131  & n290 ;
  assign n4449 = n588 & n4389 ;
  assign n4450 = n4408 & ~n4449 ;
  assign n4451 = ~n4394 & n4450 ;
  assign n4452 = n1543 & ~n4451 ;
  assign n4448 = n329 & n519 ;
  assign n4453 = n1585 & ~n2720 ;
  assign n4454 = \reg2_reg[13]/NET0131  & ~n4453 ;
  assign n4455 = ~n4448 & ~n4454 ;
  assign n4456 = ~n4452 & n4455 ;
  assign n4457 = n292 & ~n4456 ;
  assign n4458 = ~n4447 & ~n4457 ;
  assign n4459 = \state_reg[0]/NET0131  & ~n4458 ;
  assign n4460 = ~n4446 & ~n4459 ;
  assign n4461 = n3048 & ~n4451 ;
  assign n4462 = \reg0_reg[13]/NET0131  & ~n4001 ;
  assign n4463 = ~n4461 & ~n4462 ;
  assign n4464 = ~\reg3_reg[2]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n4467 = n341 & ~n347 ;
  assign n4466 = ~\IR_reg[0]/NET0131  & ~\reg1_reg[0]/NET0131  ;
  assign n4468 = \IR_reg[0]/NET0131  & \reg1_reg[0]/NET0131  ;
  assign n4469 = ~n4466 & ~n4468 ;
  assign n4470 = n4467 & n4469 ;
  assign n4471 = n341 & n347 ;
  assign n4472 = ~\IR_reg[0]/NET0131  & ~\reg2_reg[0]/NET0131  ;
  assign n4473 = \IR_reg[0]/NET0131  & \reg2_reg[0]/NET0131  ;
  assign n4474 = ~n4472 & ~n4473 ;
  assign n4475 = n4471 & n4474 ;
  assign n4476 = ~n4470 & ~n4475 ;
  assign n4465 = \IR_reg[0]/NET0131  & ~n341 ;
  assign n4477 = n289 & ~n4465 ;
  assign n4478 = n4476 & n4477 ;
  assign n4479 = ~\addr[2]_pad  & ~n289 ;
  assign n4480 = n796 & n4479 ;
  assign n4481 = ~n4478 & ~n4480 ;
  assign n4482 = ~n259 & ~n4481 ;
  assign n4508 = ~n259 & n796 ;
  assign n4509 = ~n290 & ~n4508 ;
  assign n4483 = ~n341 & n347 ;
  assign n4484 = ~n759 & n4483 ;
  assign n4485 = \reg2_reg[2]/NET0131  & ~n759 ;
  assign n4486 = ~\reg2_reg[2]/NET0131  & n759 ;
  assign n4487 = ~n4485 & ~n4486 ;
  assign n4488 = ~\reg2_reg[1]/NET0131  & ~n744 ;
  assign n4489 = \reg2_reg[1]/NET0131  & n744 ;
  assign n4490 = ~n4473 & ~n4489 ;
  assign n4491 = ~n4488 & ~n4490 ;
  assign n4492 = ~n4487 & ~n4491 ;
  assign n4493 = n4487 & n4491 ;
  assign n4494 = ~n4492 & ~n4493 ;
  assign n4495 = n4471 & n4494 ;
  assign n4510 = ~n4484 & ~n4495 ;
  assign n4496 = \reg1_reg[2]/NET0131  & ~n759 ;
  assign n4497 = ~\reg1_reg[2]/NET0131  & n759 ;
  assign n4498 = ~n4496 & ~n4497 ;
  assign n4499 = ~\reg1_reg[1]/NET0131  & ~n744 ;
  assign n4500 = \reg1_reg[1]/NET0131  & n744 ;
  assign n4501 = ~n4468 & ~n4500 ;
  assign n4502 = ~n4499 & ~n4501 ;
  assign n4503 = ~n4498 & ~n4502 ;
  assign n4504 = n4498 & n4502 ;
  assign n4505 = ~n4503 & ~n4504 ;
  assign n4506 = n4467 & n4505 ;
  assign n4507 = \addr[2]_pad  & n348 ;
  assign n4511 = ~n4506 & ~n4507 ;
  assign n4512 = n4510 & n4511 ;
  assign n4513 = n4509 & n4512 ;
  assign n4514 = ~n4482 & ~n4513 ;
  assign n4515 = \state_reg[0]/NET0131  & ~n4514 ;
  assign n4516 = ~n4464 & ~n4515 ;
  assign n4517 = ~\addr[4]_pad  & ~n289 ;
  assign n4518 = n796 & n4517 ;
  assign n4519 = ~n4478 & ~n4518 ;
  assign n4520 = ~n259 & ~n4519 ;
  assign n4536 = \reg2_reg[4]/NET0131  & ~n736 ;
  assign n4537 = ~\reg2_reg[4]/NET0131  & n736 ;
  assign n4538 = ~n4536 & ~n4537 ;
  assign n4539 = ~\reg2_reg[3]/NET0131  & ~n769 ;
  assign n4540 = \reg2_reg[3]/NET0131  & n769 ;
  assign n4541 = ~n4485 & ~n4491 ;
  assign n4542 = ~n4486 & ~n4541 ;
  assign n4543 = ~n4540 & ~n4542 ;
  assign n4544 = ~n4539 & ~n4543 ;
  assign n4546 = n4538 & n4544 ;
  assign n4545 = ~n4538 & ~n4544 ;
  assign n4547 = n4471 & ~n4545 ;
  assign n4548 = ~n4546 & n4547 ;
  assign n4521 = \reg1_reg[4]/NET0131  & ~n736 ;
  assign n4522 = ~\reg1_reg[4]/NET0131  & n736 ;
  assign n4523 = ~n4521 & ~n4522 ;
  assign n4524 = ~\reg1_reg[3]/NET0131  & ~n769 ;
  assign n4525 = \reg1_reg[3]/NET0131  & n769 ;
  assign n4526 = ~n4496 & ~n4502 ;
  assign n4527 = ~n4497 & ~n4526 ;
  assign n4528 = ~n4525 & ~n4527 ;
  assign n4529 = ~n4524 & ~n4528 ;
  assign n4531 = n4523 & n4529 ;
  assign n4530 = ~n4523 & ~n4529 ;
  assign n4532 = n4467 & ~n4530 ;
  assign n4533 = ~n4531 & n4532 ;
  assign n4534 = ~n736 & n4483 ;
  assign n4535 = \addr[4]_pad  & n348 ;
  assign n4549 = ~n4534 & ~n4535 ;
  assign n4550 = ~n4533 & n4549 ;
  assign n4551 = ~n4548 & n4550 ;
  assign n4552 = n4509 & n4551 ;
  assign n4553 = ~n4520 & ~n4552 ;
  assign n4554 = \state_reg[0]/NET0131  & ~n4553 ;
  assign n4555 = ~n3871 & ~n4554 ;
  assign n4556 = ~\addr[12]_pad  & n796 ;
  assign n4557 = n2389 & ~n4556 ;
  assign n4558 = ~n260 & ~n4557 ;
  assign n4601 = \reg1_reg[12]/NET0131  & n609 ;
  assign n4602 = ~\reg1_reg[12]/NET0131  & ~n609 ;
  assign n4603 = ~n4601 & ~n4602 ;
  assign n4604 = ~\reg1_reg[11]/NET0131  & ~n599 ;
  assign n4605 = \reg1_reg[11]/NET0131  & n599 ;
  assign n4606 = ~\reg1_reg[10]/NET0131  & ~n619 ;
  assign n4607 = ~\reg1_reg[9]/NET0131  & n627 ;
  assign n4608 = \reg1_reg[7]/NET0131  & n695 ;
  assign n4609 = ~\reg1_reg[6]/NET0131  & ~n712 ;
  assign n4610 = \reg1_reg[6]/NET0131  & n712 ;
  assign n4611 = ~\reg1_reg[5]/NET0131  & ~n721 ;
  assign n4612 = \reg1_reg[5]/NET0131  & n721 ;
  assign n4613 = ~n4521 & ~n4529 ;
  assign n4614 = ~n4522 & ~n4613 ;
  assign n4615 = ~n4612 & ~n4614 ;
  assign n4616 = ~n4611 & ~n4615 ;
  assign n4617 = ~n4610 & ~n4616 ;
  assign n4618 = ~n4609 & ~n4617 ;
  assign n4619 = ~n4608 & ~n4618 ;
  assign n4620 = ~\reg1_reg[8]/NET0131  & ~n702 ;
  assign n4621 = ~\reg1_reg[7]/NET0131  & ~n695 ;
  assign n4622 = ~n4620 & ~n4621 ;
  assign n4623 = ~n4619 & n4622 ;
  assign n4624 = \reg1_reg[9]/NET0131  & ~n627 ;
  assign n4625 = \reg1_reg[8]/NET0131  & n702 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = ~n4623 & n4626 ;
  assign n4628 = ~n4607 & ~n4627 ;
  assign n4629 = \reg1_reg[10]/NET0131  & n619 ;
  assign n4630 = ~n4628 & ~n4629 ;
  assign n4631 = ~n4606 & ~n4630 ;
  assign n4632 = ~n4605 & ~n4631 ;
  assign n4633 = ~n4604 & ~n4632 ;
  assign n4635 = ~n4603 & ~n4633 ;
  assign n4634 = n4603 & n4633 ;
  assign n4636 = n4467 & ~n4634 ;
  assign n4637 = ~n4635 & n4636 ;
  assign n4563 = \reg2_reg[12]/NET0131  & n609 ;
  assign n4564 = ~\reg2_reg[12]/NET0131  & ~n609 ;
  assign n4565 = ~n4563 & ~n4564 ;
  assign n4566 = ~\reg2_reg[11]/NET0131  & ~n599 ;
  assign n4567 = \reg2_reg[10]/NET0131  & n619 ;
  assign n4568 = \reg2_reg[11]/NET0131  & n599 ;
  assign n4569 = ~n4567 & ~n4568 ;
  assign n4570 = ~n4566 & ~n4569 ;
  assign n4571 = ~\reg2_reg[10]/NET0131  & ~n619 ;
  assign n4572 = ~n4566 & ~n4571 ;
  assign n4573 = ~\reg2_reg[9]/NET0131  & n627 ;
  assign n4576 = ~\reg2_reg[8]/NET0131  & ~n702 ;
  assign n4577 = ~\reg2_reg[7]/NET0131  & ~n695 ;
  assign n4578 = \reg2_reg[7]/NET0131  & n695 ;
  assign n4579 = ~\reg2_reg[6]/NET0131  & ~n712 ;
  assign n4580 = \reg2_reg[6]/NET0131  & n712 ;
  assign n4581 = ~\reg2_reg[5]/NET0131  & ~n721 ;
  assign n4582 = \reg2_reg[5]/NET0131  & n721 ;
  assign n4583 = ~n4536 & ~n4544 ;
  assign n4584 = ~n4537 & ~n4583 ;
  assign n4585 = ~n4582 & ~n4584 ;
  assign n4586 = ~n4581 & ~n4585 ;
  assign n4587 = ~n4580 & ~n4586 ;
  assign n4588 = ~n4579 & ~n4587 ;
  assign n4589 = ~n4578 & ~n4588 ;
  assign n4590 = ~n4577 & ~n4589 ;
  assign n4591 = ~n4576 & n4590 ;
  assign n4574 = \reg2_reg[8]/NET0131  & n702 ;
  assign n4575 = \reg2_reg[9]/NET0131  & ~n627 ;
  assign n4592 = ~n4574 & ~n4575 ;
  assign n4593 = ~n4591 & n4592 ;
  assign n4594 = ~n4573 & ~n4593 ;
  assign n4595 = n4572 & n4594 ;
  assign n4596 = ~n4570 & ~n4595 ;
  assign n4598 = ~n4565 & n4596 ;
  assign n4597 = n4565 & ~n4596 ;
  assign n4599 = n4471 & ~n4597 ;
  assign n4600 = ~n4598 & n4599 ;
  assign n4559 = n609 & n4483 ;
  assign n4560 = n796 & n2389 ;
  assign n4561 = ~n348 & ~n4560 ;
  assign n4562 = \addr[12]_pad  & ~n4561 ;
  assign n4638 = ~n4559 & ~n4562 ;
  assign n4639 = ~n4600 & n4638 ;
  assign n4640 = ~n4637 & n4639 ;
  assign n4641 = ~n4558 & ~n4640 ;
  assign n4642 = ~n1692 & ~n4641 ;
  assign n4643 = ~\addr[13]_pad  & n796 ;
  assign n4644 = n2389 & ~n4643 ;
  assign n4646 = ~n260 & ~n4644 ;
  assign n4653 = \reg1_reg[13]/NET0131  & n651 ;
  assign n4648 = ~n4604 & ~n4606 ;
  assign n4649 = ~n4630 & n4648 ;
  assign n4650 = ~n4601 & ~n4605 ;
  assign n4651 = ~n4649 & n4650 ;
  assign n4652 = ~n4602 & ~n4651 ;
  assign n4654 = ~\reg1_reg[13]/NET0131  & ~n651 ;
  assign n4657 = n4652 & ~n4654 ;
  assign n4658 = ~n4653 & n4657 ;
  assign n4655 = ~n4653 & ~n4654 ;
  assign n4656 = ~n4652 & ~n4655 ;
  assign n4659 = n4467 & ~n4656 ;
  assign n4660 = ~n4658 & n4659 ;
  assign n4662 = \reg2_reg[13]/NET0131  & n651 ;
  assign n4663 = ~\reg2_reg[13]/NET0131  & ~n651 ;
  assign n4664 = ~n4662 & ~n4663 ;
  assign n4665 = ~n4576 & ~n4577 ;
  assign n4666 = n4588 & n4665 ;
  assign n4667 = ~n4576 & n4578 ;
  assign n4668 = ~n4574 & ~n4667 ;
  assign n4669 = ~n4666 & n4668 ;
  assign n4670 = ~n4573 & ~n4669 ;
  assign n4671 = ~n4567 & ~n4575 ;
  assign n4672 = ~n4670 & n4671 ;
  assign n4673 = n4572 & ~n4672 ;
  assign n4674 = ~n4563 & ~n4568 ;
  assign n4675 = ~n4673 & n4674 ;
  assign n4676 = ~n4564 & ~n4675 ;
  assign n4678 = ~n4664 & ~n4676 ;
  assign n4677 = n4664 & n4676 ;
  assign n4679 = n4471 & ~n4677 ;
  assign n4680 = ~n4678 & n4679 ;
  assign n4647 = n651 & n4483 ;
  assign n4661 = \addr[13]_pad  & n348 ;
  assign n4681 = ~n4647 & ~n4661 ;
  assign n4682 = ~n4680 & n4681 ;
  assign n4683 = ~n4660 & n4682 ;
  assign n4684 = ~n4646 & ~n4683 ;
  assign n4645 = n796 & n4644 ;
  assign n4685 = \reg3_reg[13]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n4686 = ~n4645 & ~n4685 ;
  assign n4687 = ~n4684 & n4686 ;
  assign n4688 = ~\addr[14]_pad  & n796 ;
  assign n4689 = n2389 & ~n4688 ;
  assign n4690 = ~n260 & ~n4689 ;
  assign n4705 = \reg1_reg[14]/NET0131  & ~n643 ;
  assign n4706 = ~\reg1_reg[14]/NET0131  & n643 ;
  assign n4707 = ~n4705 & ~n4706 ;
  assign n4708 = ~n4602 & n4633 ;
  assign n4709 = ~n4601 & ~n4653 ;
  assign n4710 = ~n4708 & n4709 ;
  assign n4711 = ~n4654 & ~n4710 ;
  assign n4713 = ~n4707 & ~n4711 ;
  assign n4712 = n4707 & n4711 ;
  assign n4714 = n4467 & ~n4712 ;
  assign n4715 = ~n4713 & n4714 ;
  assign n4693 = \reg2_reg[14]/NET0131  & ~n643 ;
  assign n4694 = ~\reg2_reg[14]/NET0131  & n643 ;
  assign n4695 = ~n4693 & ~n4694 ;
  assign n4696 = ~n4564 & ~n4663 ;
  assign n4697 = ~n4596 & n4696 ;
  assign n4698 = n4563 & ~n4663 ;
  assign n4699 = ~n4662 & ~n4698 ;
  assign n4700 = ~n4697 & n4699 ;
  assign n4702 = ~n4695 & n4700 ;
  assign n4701 = n4695 & ~n4700 ;
  assign n4703 = n4471 & ~n4701 ;
  assign n4704 = ~n4702 & n4703 ;
  assign n4691 = \addr[14]_pad  & ~n4561 ;
  assign n4692 = ~n643 & n4483 ;
  assign n4716 = ~n4691 & ~n4692 ;
  assign n4717 = ~n4704 & n4716 ;
  assign n4718 = ~n4715 & n4717 ;
  assign n4719 = ~n4690 & ~n4718 ;
  assign n4720 = ~n2192 & ~n4719 ;
  assign n4721 = ~\addr[15]_pad  & n796 ;
  assign n4722 = n2389 & ~n4721 ;
  assign n4723 = ~n260 & ~n4722 ;
  assign n4738 = \reg1_reg[15]/NET0131  & n668 ;
  assign n4739 = ~\reg1_reg[15]/NET0131  & ~n668 ;
  assign n4740 = ~n4738 & ~n4739 ;
  assign n4741 = ~n4653 & ~n4705 ;
  assign n4742 = ~n4657 & n4741 ;
  assign n4743 = ~n4706 & ~n4742 ;
  assign n4745 = ~n4740 & ~n4743 ;
  assign n4744 = n4740 & n4743 ;
  assign n4746 = n4467 & ~n4744 ;
  assign n4747 = ~n4745 & n4746 ;
  assign n4726 = \reg2_reg[15]/NET0131  & n668 ;
  assign n4727 = ~\reg2_reg[15]/NET0131  & ~n668 ;
  assign n4728 = ~n4726 & ~n4727 ;
  assign n4729 = ~n4694 & n4696 ;
  assign n4730 = ~n4675 & n4729 ;
  assign n4731 = n4662 & ~n4694 ;
  assign n4732 = ~n4693 & ~n4731 ;
  assign n4733 = ~n4730 & n4732 ;
  assign n4735 = ~n4728 & n4733 ;
  assign n4734 = n4728 & ~n4733 ;
  assign n4736 = n4471 & ~n4734 ;
  assign n4737 = ~n4735 & n4736 ;
  assign n4724 = \addr[15]_pad  & ~n4561 ;
  assign n4725 = n668 & n4483 ;
  assign n4748 = ~n4724 & ~n4725 ;
  assign n4749 = ~n4737 & n4748 ;
  assign n4750 = ~n4747 & n4749 ;
  assign n4751 = ~n4723 & ~n4750 ;
  assign n4752 = ~n1599 & ~n4751 ;
  assign n4753 = ~\addr[17]_pad  & n796 ;
  assign n4754 = n2389 & ~n4753 ;
  assign n4756 = ~n260 & ~n4754 ;
  assign n4757 = \reg1_reg[17]/NET0131  & n353 ;
  assign n4758 = ~\reg1_reg[17]/NET0131  & ~n353 ;
  assign n4759 = ~n4757 & ~n4758 ;
  assign n4760 = ~\reg1_reg[16]/NET0131  & ~n660 ;
  assign n4761 = ~n4739 & n4743 ;
  assign n4762 = \reg1_reg[16]/NET0131  & n660 ;
  assign n4763 = ~n4738 & ~n4762 ;
  assign n4764 = ~n4761 & n4763 ;
  assign n4765 = ~n4760 & ~n4764 ;
  assign n4767 = n4759 & n4765 ;
  assign n4766 = ~n4759 & ~n4765 ;
  assign n4768 = n4467 & ~n4766 ;
  assign n4769 = ~n4767 & n4768 ;
  assign n4772 = \reg2_reg[17]/NET0131  & n353 ;
  assign n4773 = ~\reg2_reg[17]/NET0131  & ~n353 ;
  assign n4774 = ~n4772 & ~n4773 ;
  assign n4775 = ~\reg2_reg[16]/NET0131  & ~n660 ;
  assign n4776 = ~n4727 & ~n4733 ;
  assign n4777 = \reg2_reg[16]/NET0131  & n660 ;
  assign n4778 = ~n4726 & ~n4777 ;
  assign n4779 = ~n4776 & n4778 ;
  assign n4780 = ~n4775 & ~n4779 ;
  assign n4782 = ~n4774 & ~n4780 ;
  assign n4781 = n4774 & n4780 ;
  assign n4783 = n4471 & ~n4781 ;
  assign n4784 = ~n4782 & n4783 ;
  assign n4770 = n353 & n4483 ;
  assign n4771 = \addr[17]_pad  & n348 ;
  assign n4785 = ~n4770 & ~n4771 ;
  assign n4786 = ~n4784 & n4785 ;
  assign n4787 = ~n4769 & n4786 ;
  assign n4788 = ~n4756 & ~n4787 ;
  assign n4755 = n796 & n4754 ;
  assign n4789 = ~n217 & ~n4755 ;
  assign n4790 = ~n4788 & n4789 ;
  assign n4791 = ~\addr[18]_pad  & n796 ;
  assign n4792 = n2389 & ~n4791 ;
  assign n4793 = ~n260 & ~n4792 ;
  assign n4811 = \reg1_reg[18]/NET0131  & n1035 ;
  assign n4812 = ~\reg1_reg[18]/NET0131  & ~n1035 ;
  assign n4813 = ~n4811 & ~n4812 ;
  assign n4814 = ~n4706 & n4711 ;
  assign n4815 = ~n4705 & ~n4738 ;
  assign n4816 = ~n4814 & n4815 ;
  assign n4817 = ~n4739 & ~n4816 ;
  assign n4818 = ~n4760 & n4817 ;
  assign n4819 = ~n4757 & ~n4762 ;
  assign n4820 = ~n4818 & n4819 ;
  assign n4821 = ~n4758 & ~n4820 ;
  assign n4823 = n4813 & n4821 ;
  assign n4822 = ~n4813 & ~n4821 ;
  assign n4824 = n4467 & ~n4822 ;
  assign n4825 = ~n4823 & n4824 ;
  assign n4796 = \reg2_reg[18]/NET0131  & n1035 ;
  assign n4797 = ~\reg2_reg[18]/NET0131  & ~n1035 ;
  assign n4798 = ~n4796 & ~n4797 ;
  assign n4799 = ~n4694 & ~n4700 ;
  assign n4800 = ~n4693 & ~n4726 ;
  assign n4801 = ~n4799 & n4800 ;
  assign n4802 = ~n4727 & ~n4801 ;
  assign n4803 = ~n4775 & n4802 ;
  assign n4804 = ~n4772 & ~n4777 ;
  assign n4805 = ~n4803 & n4804 ;
  assign n4806 = ~n4773 & ~n4805 ;
  assign n4808 = ~n4798 & ~n4806 ;
  assign n4807 = n4798 & n4806 ;
  assign n4809 = n4471 & ~n4807 ;
  assign n4810 = ~n4808 & n4809 ;
  assign n4794 = n1035 & n4483 ;
  assign n4795 = \addr[18]_pad  & n348 ;
  assign n4826 = ~n4794 & ~n4795 ;
  assign n4827 = ~n4810 & n4826 ;
  assign n4828 = ~n4825 & n4827 ;
  assign n4829 = ~n4793 & ~n4828 ;
  assign n4830 = n796 & n4792 ;
  assign n4831 = ~n2823 & ~n4830 ;
  assign n4832 = ~n4829 & n4831 ;
  assign n4833 = ~\addr[19]_pad  & n796 ;
  assign n4834 = n2389 & ~n4833 ;
  assign n4835 = ~n260 & ~n4834 ;
  assign n4849 = ~n4757 & ~n4765 ;
  assign n4850 = ~n4758 & ~n4812 ;
  assign n4851 = ~n4849 & n4850 ;
  assign n4852 = ~n4811 & ~n4851 ;
  assign n4853 = \reg1_reg[19]/NET0131  & n327 ;
  assign n4854 = ~\reg1_reg[19]/NET0131  & ~n327 ;
  assign n4855 = ~n4853 & ~n4854 ;
  assign n4857 = ~n4852 & n4855 ;
  assign n4856 = n4852 & ~n4855 ;
  assign n4858 = n4467 & ~n4856 ;
  assign n4859 = ~n4857 & n4858 ;
  assign n4838 = ~n4773 & n4780 ;
  assign n4839 = ~n4772 & ~n4796 ;
  assign n4840 = ~n4838 & n4839 ;
  assign n4841 = ~n4797 & ~n4840 ;
  assign n4842 = \reg2_reg[19]/NET0131  & ~n4841 ;
  assign n4843 = ~\reg2_reg[19]/NET0131  & n4841 ;
  assign n4844 = ~n4842 & ~n4843 ;
  assign n4846 = ~n327 & n4844 ;
  assign n4845 = n327 & ~n4844 ;
  assign n4847 = n4471 & ~n4845 ;
  assign n4848 = ~n4846 & n4847 ;
  assign n4836 = \addr[19]_pad  & n348 ;
  assign n4837 = n327 & n4483 ;
  assign n4860 = ~n4836 & ~n4837 ;
  assign n4861 = ~n4848 & n4860 ;
  assign n4862 = ~n4859 & n4861 ;
  assign n4863 = ~n4835 & ~n4862 ;
  assign n4864 = n796 & n4834 ;
  assign n4865 = ~n1774 & ~n4864 ;
  assign n4866 = ~n4863 & n4865 ;
  assign n4867 = \reg3_reg[1]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n4868 = ~\addr[1]_pad  & n796 ;
  assign n4869 = n2389 & ~n4868 ;
  assign n4870 = ~n260 & ~n4869 ;
  assign n4871 = \addr[1]_pad  & ~n4561 ;
  assign n4878 = ~n4488 & ~n4489 ;
  assign n4879 = ~n4473 & ~n4878 ;
  assign n4880 = n4473 & n4878 ;
  assign n4881 = ~n4879 & ~n4880 ;
  assign n4882 = n4471 & n4881 ;
  assign n4872 = ~n4499 & ~n4500 ;
  assign n4873 = ~n4468 & ~n4872 ;
  assign n4874 = n4468 & n4872 ;
  assign n4875 = ~n4873 & ~n4874 ;
  assign n4876 = n4467 & n4875 ;
  assign n4877 = n744 & n4483 ;
  assign n4883 = ~n4876 & ~n4877 ;
  assign n4884 = ~n4882 & n4883 ;
  assign n4885 = ~n4871 & n4884 ;
  assign n4886 = ~n4870 & ~n4885 ;
  assign n4887 = ~n4867 & ~n4886 ;
  assign n4888 = \reg3_reg[3]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n4889 = ~\addr[3]_pad  & n796 ;
  assign n4890 = n2389 & ~n4889 ;
  assign n4891 = ~n260 & ~n4890 ;
  assign n4892 = \addr[3]_pad  & ~n4561 ;
  assign n4899 = ~n4524 & ~n4525 ;
  assign n4900 = ~n4527 & ~n4899 ;
  assign n4901 = n4527 & n4899 ;
  assign n4902 = ~n4900 & ~n4901 ;
  assign n4903 = n4467 & n4902 ;
  assign n4893 = ~n4539 & ~n4540 ;
  assign n4894 = ~n4542 & ~n4893 ;
  assign n4895 = n4542 & n4893 ;
  assign n4896 = ~n4894 & ~n4895 ;
  assign n4897 = n4471 & n4896 ;
  assign n4898 = n769 & n4483 ;
  assign n4904 = ~n4897 & ~n4898 ;
  assign n4905 = ~n4903 & n4904 ;
  assign n4906 = ~n4892 & n4905 ;
  assign n4907 = ~n4891 & ~n4906 ;
  assign n4908 = ~n4888 & ~n4907 ;
  assign n4918 = ~n4581 & ~n4582 ;
  assign n4920 = n4584 & n4918 ;
  assign n4919 = ~n4584 & ~n4918 ;
  assign n4921 = n4471 & ~n4919 ;
  assign n4922 = ~n4920 & n4921 ;
  assign n4912 = ~n4611 & ~n4612 ;
  assign n4914 = n4614 & n4912 ;
  assign n4913 = ~n4614 & ~n4912 ;
  assign n4915 = n4467 & ~n4913 ;
  assign n4916 = ~n4914 & n4915 ;
  assign n4911 = n721 & n4483 ;
  assign n4917 = \addr[5]_pad  & n348 ;
  assign n4923 = ~n4911 & ~n4917 ;
  assign n4924 = ~n4916 & n4923 ;
  assign n4925 = ~n4922 & n4924 ;
  assign n4926 = \state_reg[0]/NET0131  & n4509 ;
  assign n4927 = ~n4925 & n4926 ;
  assign n4909 = \addr[5]_pad  & n4560 ;
  assign n4910 = \reg3_reg[5]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n4928 = ~n4909 & ~n4910 ;
  assign n4929 = ~n4927 & n4928 ;
  assign n4930 = ~\addr[6]_pad  & n796 ;
  assign n4931 = n2389 & ~n4930 ;
  assign n4932 = ~n260 & ~n4931 ;
  assign n4933 = \addr[6]_pad  & ~n4561 ;
  assign n4944 = n712 & n4483 ;
  assign n4945 = ~n4933 & ~n4944 ;
  assign n4934 = ~n4609 & ~n4610 ;
  assign n4936 = n4616 & n4934 ;
  assign n4935 = ~n4616 & ~n4934 ;
  assign n4937 = n4467 & ~n4935 ;
  assign n4938 = ~n4936 & n4937 ;
  assign n4939 = ~n4579 & ~n4580 ;
  assign n4941 = n4586 & n4939 ;
  assign n4940 = ~n4586 & ~n4939 ;
  assign n4942 = n4471 & ~n4940 ;
  assign n4943 = ~n4941 & n4942 ;
  assign n4946 = ~n4938 & ~n4943 ;
  assign n4947 = n4945 & n4946 ;
  assign n4948 = ~n4932 & ~n4947 ;
  assign n4949 = ~n3444 & ~n4948 ;
  assign n4950 = ~\addr[7]_pad  & n796 ;
  assign n4951 = n2389 & ~n4950 ;
  assign n4953 = ~n260 & ~n4951 ;
  assign n4961 = ~n4608 & ~n4621 ;
  assign n4963 = n4618 & n4961 ;
  assign n4962 = ~n4618 & ~n4961 ;
  assign n4964 = n4467 & ~n4962 ;
  assign n4965 = ~n4963 & n4964 ;
  assign n4956 = ~n4577 & ~n4578 ;
  assign n4958 = n4588 & n4956 ;
  assign n4957 = ~n4588 & ~n4956 ;
  assign n4959 = n4471 & ~n4957 ;
  assign n4960 = ~n4958 & n4959 ;
  assign n4954 = n695 & n4483 ;
  assign n4955 = \addr[7]_pad  & n348 ;
  assign n4966 = ~n4954 & ~n4955 ;
  assign n4967 = ~n4960 & n4966 ;
  assign n4968 = ~n4965 & n4967 ;
  assign n4969 = ~n4953 & ~n4968 ;
  assign n4952 = n796 & n4951 ;
  assign n4970 = ~n2301 & ~n4952 ;
  assign n4971 = ~n4969 & n4970 ;
  assign n4972 = ~\addr[8]_pad  & n796 ;
  assign n4973 = n2389 & ~n4972 ;
  assign n4974 = ~n260 & ~n4973 ;
  assign n4982 = ~n4619 & ~n4621 ;
  assign n4983 = ~n4620 & ~n4625 ;
  assign n4985 = n4982 & n4983 ;
  assign n4984 = ~n4982 & ~n4983 ;
  assign n4986 = n4467 & ~n4984 ;
  assign n4987 = ~n4985 & n4986 ;
  assign n4977 = ~n4574 & ~n4576 ;
  assign n4979 = n4590 & n4977 ;
  assign n4978 = ~n4590 & ~n4977 ;
  assign n4980 = n4471 & ~n4978 ;
  assign n4981 = ~n4979 & n4980 ;
  assign n4975 = n702 & n4483 ;
  assign n4976 = \addr[8]_pad  & ~n4561 ;
  assign n4988 = ~n4975 & ~n4976 ;
  assign n4989 = ~n4981 & n4988 ;
  assign n4990 = ~n4987 & n4989 ;
  assign n4991 = ~n4974 & ~n4990 ;
  assign n4992 = ~n3485 & ~n4991 ;
  assign n4993 = ~\addr[9]_pad  & n796 ;
  assign n4994 = n2389 & ~n4993 ;
  assign n4995 = ~n260 & ~n4994 ;
  assign n4996 = ~n4623 & ~n4625 ;
  assign n4997 = ~n4607 & ~n4624 ;
  assign n4999 = n4996 & ~n4997 ;
  assign n4998 = ~n4996 & n4997 ;
  assign n5000 = n4467 & ~n4998 ;
  assign n5001 = ~n4999 & n5000 ;
  assign n5004 = ~n4573 & ~n4575 ;
  assign n5006 = ~n4669 & n5004 ;
  assign n5005 = n4669 & ~n5004 ;
  assign n5007 = n4471 & ~n5005 ;
  assign n5008 = ~n5006 & n5007 ;
  assign n5002 = ~n627 & n4483 ;
  assign n5003 = \addr[9]_pad  & ~n4561 ;
  assign n5009 = ~n5002 & ~n5003 ;
  assign n5010 = ~n5008 & n5009 ;
  assign n5011 = ~n5001 & n5010 ;
  assign n5012 = ~n4995 & ~n5011 ;
  assign n5013 = ~n3513 & ~n5012 ;
  assign n5014 = ~\addr[11]_pad  & n796 ;
  assign n5015 = n2389 & ~n5014 ;
  assign n5017 = ~n260 & ~n5015 ;
  assign n5021 = ~n4605 & n4649 ;
  assign n5019 = ~n4604 & ~n4605 ;
  assign n5020 = ~n4631 & ~n5019 ;
  assign n5022 = n4467 & ~n5020 ;
  assign n5023 = ~n5021 & n5022 ;
  assign n5028 = ~n4568 & n4673 ;
  assign n5025 = ~n4566 & ~n4568 ;
  assign n5026 = ~n4571 & ~n4672 ;
  assign n5027 = ~n5025 & ~n5026 ;
  assign n5029 = n4471 & ~n5027 ;
  assign n5030 = ~n5028 & n5029 ;
  assign n5018 = n599 & n4483 ;
  assign n5024 = \addr[11]_pad  & n348 ;
  assign n5031 = ~n5018 & ~n5024 ;
  assign n5032 = ~n5030 & n5031 ;
  assign n5033 = ~n5023 & n5032 ;
  assign n5034 = ~n5017 & ~n5033 ;
  assign n5016 = n796 & n5015 ;
  assign n5035 = ~n1646 & ~n5016 ;
  assign n5036 = ~n5034 & n5035 ;
  assign n5037 = ~n348 & n4509 ;
  assign n5038 = \state_reg[0]/NET0131  & ~n5037 ;
  assign n5039 = \reg3_reg[0]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n5040 = ~\addr[0]_pad  & n796 ;
  assign n5041 = n2389 & ~n5040 ;
  assign n5042 = ~n260 & ~n5041 ;
  assign n5044 = \addr[0]_pad  & ~n4561 ;
  assign n5043 = n347 & n4465 ;
  assign n5045 = n4476 & ~n5043 ;
  assign n5046 = ~n5044 & n5045 ;
  assign n5047 = ~n5042 & ~n5046 ;
  assign n5048 = ~n5039 & ~n5047 ;
  assign n5049 = \reg3_reg[10]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n5050 = ~\addr[10]_pad  & n796 ;
  assign n5051 = n2389 & ~n5050 ;
  assign n5052 = ~n260 & ~n5051 ;
  assign n5060 = ~n4567 & ~n4571 ;
  assign n5062 = ~n4594 & ~n5060 ;
  assign n5061 = n4594 & n5060 ;
  assign n5063 = n4471 & ~n5061 ;
  assign n5064 = ~n5062 & n5063 ;
  assign n5055 = ~n4606 & ~n4629 ;
  assign n5057 = ~n4628 & ~n5055 ;
  assign n5056 = n4628 & n5055 ;
  assign n5058 = n4467 & ~n5056 ;
  assign n5059 = ~n5057 & n5058 ;
  assign n5053 = \addr[10]_pad  & ~n4561 ;
  assign n5054 = n619 & n4483 ;
  assign n5065 = ~n5053 & ~n5054 ;
  assign n5066 = ~n5059 & n5065 ;
  assign n5067 = ~n5064 & n5066 ;
  assign n5068 = ~n5052 & ~n5067 ;
  assign n5069 = ~n5049 & ~n5068 ;
  assign n5070 = ~\addr[16]_pad  & n796 ;
  assign n5071 = n2389 & ~n5070 ;
  assign n5073 = ~n260 & ~n5071 ;
  assign n5075 = ~n4760 & ~n4762 ;
  assign n5077 = n4817 & n5075 ;
  assign n5076 = ~n4817 & ~n5075 ;
  assign n5078 = n4467 & ~n5076 ;
  assign n5079 = ~n5077 & n5078 ;
  assign n5081 = ~n4775 & ~n4777 ;
  assign n5083 = n4802 & n5081 ;
  assign n5082 = ~n4802 & ~n5081 ;
  assign n5084 = n4471 & ~n5082 ;
  assign n5085 = ~n5083 & n5084 ;
  assign n5074 = \addr[16]_pad  & n348 ;
  assign n5080 = n660 & n4483 ;
  assign n5086 = ~n5074 & ~n5080 ;
  assign n5087 = ~n5085 & n5086 ;
  assign n5088 = ~n5079 & n5087 ;
  assign n5089 = ~n5073 & ~n5088 ;
  assign n5072 = n796 & n5071 ;
  assign n5090 = ~n2256 & ~n5072 ;
  assign n5091 = ~n5089 & n5090 ;
  assign n5092 = \state_reg[0]/NET0131  & n290 ;
  assign n5093 = \datao[15]_pad  & ~n289 ;
  assign n5094 = n289 & ~n537 ;
  assign n5095 = ~n5093 & ~n5094 ;
  assign n5096 = \datao[28]_pad  & ~n289 ;
  assign n5097 = n289 & ~n1138 ;
  assign n5098 = ~n5096 & ~n5097 ;
  assign n5099 = \datao[8]_pad  & ~n289 ;
  assign n5100 = n289 & ~n465 ;
  assign n5101 = ~n5099 & ~n5100 ;
  assign n5102 = \state_reg[0]/NET0131  & n347 ;
  assign n5103 = \datai[27]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5104 = ~n5102 & ~n5103 ;
  assign n5105 = \state_reg[0]/NET0131  & n371 ;
  assign n5106 = \datai[30]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5107 = ~n5105 & ~n5106 ;
  assign n5108 = \state_reg[0]/NET0131  & n341 ;
  assign n5109 = \datai[28]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5110 = ~n5108 & ~n5109 ;
  assign n5111 = \state_reg[0]/NET0131  & n365 ;
  assign n5112 = \datai[29]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5113 = ~n5111 & ~n5112 ;
  assign n5114 = ~\datai[31]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5115 = ~\IR_reg[29]/NET0131  & ~\IR_reg[30]/NET0131  ;
  assign n5116 = \IR_reg[31]/NET0131  & n5115 ;
  assign n5117 = n361 & n5116 ;
  assign n5118 = \state_reg[0]/NET0131  & ~n5117 ;
  assign n5119 = ~n5114 & ~n5118 ;
  assign n5120 = \state_reg[0]/NET0131  & ~n668 ;
  assign n5121 = ~\datai[15]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5122 = ~n5120 & ~n5121 ;
  assign n5123 = \datai[23]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5124 = ~n260 & ~n5123 ;
  assign n5125 = \state_reg[0]/NET0131  & n287 ;
  assign n5126 = \datai[24]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5127 = ~n5125 & ~n5126 ;
  assign n5128 = \state_reg[0]/NET0131  & ~n353 ;
  assign n5129 = ~\datai[17]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5130 = ~n5128 & ~n5129 ;
  assign n5131 = \state_reg[0]/NET0131  & ~n312 ;
  assign n5132 = \datai[22]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5133 = ~n5131 & ~n5132 ;
  assign n5134 = \state_reg[0]/NET0131  & n327 ;
  assign n5135 = \datai[19]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5136 = ~n5134 & ~n5135 ;
  assign n5137 = ~\datai[16]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5138 = \state_reg[0]/NET0131  & ~n660 ;
  assign n5139 = ~n5137 & ~n5138 ;
  assign n5140 = \state_reg[0]/NET0131  & n318 ;
  assign n5141 = \datai[21]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5142 = ~n5140 & ~n5141 ;
  assign n5143 = ~\datai[20]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5144 = \state_reg[0]/NET0131  & ~n322 ;
  assign n5145 = ~n5143 & ~n5144 ;
  assign n5146 = \datai[26]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5147 = \state_reg[0]/NET0131  & ~n272 ;
  assign n5148 = ~n5146 & ~n5147 ;
  assign n5149 = \datai[25]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5150 = \state_reg[0]/NET0131  & ~n281 ;
  assign n5151 = ~n5149 & ~n5150 ;
  assign n5152 = \state_reg[0]/NET0131  & n599 ;
  assign n5153 = \datai[11]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5154 = ~n5152 & ~n5153 ;
  assign n5155 = \state_reg[0]/NET0131  & n651 ;
  assign n5156 = \datai[13]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5157 = ~n5155 & ~n5156 ;
  assign n5158 = \datai[14]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5159 = \state_reg[0]/NET0131  & ~n643 ;
  assign n5160 = ~n5158 & ~n5159 ;
  assign n5161 = \state_reg[0]/NET0131  & n609 ;
  assign n5162 = \datai[12]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5163 = ~n5161 & ~n5162 ;
  assign n5164 = \state_reg[0]/NET0131  & ~n1035 ;
  assign n5165 = ~\datai[18]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5166 = ~n5164 & ~n5165 ;
  assign n5167 = \state_reg[0]/NET0131  & ~n627 ;
  assign n5168 = \datai[9]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5169 = ~n5167 & ~n5168 ;
  assign n5170 = \state_reg[0]/NET0131  & n695 ;
  assign n5171 = \datai[7]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5172 = ~n5170 & ~n5171 ;
  assign n5173 = \state_reg[0]/NET0131  & n619 ;
  assign n5174 = \datai[10]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5175 = ~n5173 & ~n5174 ;
  assign n5176 = \state_reg[0]/NET0131  & n702 ;
  assign n5177 = \datai[8]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5178 = ~n5176 & ~n5177 ;
  assign n5179 = \state_reg[0]/NET0131  & n712 ;
  assign n5180 = \datai[6]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5181 = ~n5179 & ~n5180 ;
  assign n5182 = \state_reg[0]/NET0131  & ~n736 ;
  assign n5183 = \datai[4]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5184 = ~n5182 & ~n5183 ;
  assign n5185 = ~\datai[5]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5186 = \state_reg[0]/NET0131  & ~n721 ;
  assign n5187 = ~n5185 & ~n5186 ;
  assign n5188 = \state_reg[0]/NET0131  & n769 ;
  assign n5189 = \datai[3]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5190 = ~n5188 & ~n5189 ;
  assign n5191 = \datai[2]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5192 = \state_reg[0]/NET0131  & ~n759 ;
  assign n5193 = ~n5191 & ~n5192 ;
  assign n5194 = \state_reg[0]/NET0131  & n744 ;
  assign n5195 = \datai[1]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5196 = ~n5194 & ~n5195 ;
  assign n5197 = \reg2_reg[24]/NET0131  & ~n2390 ;
  assign n5199 = \reg2_reg[24]/NET0131  & ~n1543 ;
  assign n5203 = n1543 & ~n1792 ;
  assign n5204 = ~n5199 & ~n5203 ;
  assign n5205 = n881 & ~n5204 ;
  assign n5209 = n1543 & ~n1826 ;
  assign n5210 = ~n5199 & ~n5209 ;
  assign n5211 = n798 & ~n5210 ;
  assign n5200 = n1543 & ~n1810 ;
  assign n5201 = ~n5199 & ~n5200 ;
  assign n5202 = n588 & ~n5201 ;
  assign n5206 = n1543 & n1798 ;
  assign n5207 = ~n5199 & ~n5206 ;
  assign n5208 = n907 & ~n5207 ;
  assign n5198 = n329 & n981 ;
  assign n5212 = n976 & n1543 ;
  assign n5213 = ~n5199 & ~n5212 ;
  assign n5214 = n910 & ~n5213 ;
  assign n5215 = ~n5198 & ~n5214 ;
  assign n5216 = ~n5208 & n5215 ;
  assign n5217 = ~n5202 & n5216 ;
  assign n5218 = ~n5211 & n5217 ;
  assign n5219 = ~n5205 & n5218 ;
  assign n5220 = n2389 & ~n5219 ;
  assign n5221 = ~n5197 & ~n5220 ;
  assign n5224 = ~\reg3_reg[3]/NET0131  & ~n308 ;
  assign n5225 = n308 & ~n3595 ;
  assign n5226 = ~n5224 & ~n5225 ;
  assign n5227 = n588 & ~n5226 ;
  assign n5228 = n308 & ~n3603 ;
  assign n5229 = ~n5224 & ~n5228 ;
  assign n5230 = n881 & ~n5229 ;
  assign n5231 = n308 & n3610 ;
  assign n5232 = ~n5224 & ~n5231 ;
  assign n5233 = n798 & ~n5232 ;
  assign n5223 = n308 & ~n3588 ;
  assign n5234 = n329 & ~n772 ;
  assign n5235 = ~\reg3_reg[3]/NET0131  & ~n1424 ;
  assign n5236 = ~n5234 & ~n5235 ;
  assign n5237 = ~n5223 & n5236 ;
  assign n5238 = ~n5233 & n5237 ;
  assign n5239 = ~n5230 & n5238 ;
  assign n5240 = ~n5227 & n5239 ;
  assign n5241 = n292 & ~n5240 ;
  assign n5242 = ~\reg3_reg[3]/NET0131  & n290 ;
  assign n5243 = ~n5241 & ~n5242 ;
  assign n5244 = \state_reg[0]/NET0131  & ~n5243 ;
  assign n5222 = ~\reg3_reg[3]/NET0131  & n260 ;
  assign n5245 = ~n4888 & ~n5222 ;
  assign n5246 = ~n5244 & n5245 ;
  assign n5247 = \reg2_reg[11]/NET0131  & ~n2390 ;
  assign n5249 = \reg2_reg[11]/NET0131  & ~n1543 ;
  assign n5250 = n1543 & n1663 ;
  assign n5251 = ~n5249 & ~n5250 ;
  assign n5252 = n588 & ~n5251 ;
  assign n5259 = n1543 & n1676 ;
  assign n5260 = ~n5249 & ~n5259 ;
  assign n5261 = n907 & ~n5260 ;
  assign n5248 = n329 & n500 ;
  assign n5262 = ~n602 & n1543 ;
  assign n5263 = ~n5249 & ~n5262 ;
  assign n5264 = n910 & ~n5263 ;
  assign n5265 = ~n5248 & ~n5264 ;
  assign n5266 = ~n5261 & n5265 ;
  assign n5267 = ~n5252 & n5266 ;
  assign n5253 = n1543 & ~n1654 ;
  assign n5254 = ~n5249 & ~n5253 ;
  assign n5255 = n798 & ~n5254 ;
  assign n5256 = n1543 & n1669 ;
  assign n5257 = ~n5249 & ~n5256 ;
  assign n5258 = n881 & ~n5257 ;
  assign n5268 = ~n5255 & ~n5258 ;
  assign n5269 = n5267 & n5268 ;
  assign n5270 = n2389 & ~n5269 ;
  assign n5271 = ~n5247 & ~n5270 ;
  assign n5273 = n290 & n519 ;
  assign n5275 = n308 & ~n4450 ;
  assign n5274 = n333 & ~n654 ;
  assign n5276 = n519 & ~n3369 ;
  assign n5277 = ~n5274 & ~n5276 ;
  assign n5278 = ~n5275 & n5277 ;
  assign n5279 = n292 & ~n5278 ;
  assign n5280 = ~n5273 & ~n5279 ;
  assign n5281 = \state_reg[0]/NET0131  & ~n5280 ;
  assign n5272 = n260 & n519 ;
  assign n5282 = ~n4685 & ~n5272 ;
  assign n5283 = ~n5281 & n5282 ;
  assign n5285 = n290 & n508 ;
  assign n5287 = ~n308 & n508 ;
  assign n5288 = n308 & n3710 ;
  assign n5289 = ~n5287 & ~n5288 ;
  assign n5290 = n588 & ~n5289 ;
  assign n5291 = n308 & n3716 ;
  assign n5292 = ~n5287 & ~n5291 ;
  assign n5293 = n881 & ~n5292 ;
  assign n5294 = n308 & n3694 ;
  assign n5295 = ~n5287 & ~n5294 ;
  assign n5296 = n907 & ~n5295 ;
  assign n5297 = n308 & n3701 ;
  assign n5286 = n333 & ~n622 ;
  assign n5298 = n508 & ~n2448 ;
  assign n5299 = ~n5286 & ~n5298 ;
  assign n5300 = ~n5297 & n5299 ;
  assign n5301 = ~n5296 & n5300 ;
  assign n5302 = ~n5293 & n5301 ;
  assign n5303 = ~n5290 & n5302 ;
  assign n5304 = n292 & ~n5303 ;
  assign n5305 = ~n5285 & ~n5304 ;
  assign n5306 = \state_reg[0]/NET0131  & ~n5305 ;
  assign n5284 = n260 & n508 ;
  assign n5307 = ~n5049 & ~n5284 ;
  assign n5308 = ~n5306 & n5307 ;
  assign n5310 = n290 & n447 ;
  assign n5312 = ~n308 & n447 ;
  assign n5313 = n308 & ~n4026 ;
  assign n5314 = ~n5312 & ~n5313 ;
  assign n5315 = n588 & ~n5314 ;
  assign n5319 = n308 & n4033 ;
  assign n5320 = ~n5312 & ~n5319 ;
  assign n5321 = n881 & ~n5320 ;
  assign n5316 = n308 & n4039 ;
  assign n5317 = ~n5312 & ~n5316 ;
  assign n5318 = n798 & ~n5317 ;
  assign n5322 = n308 & n4046 ;
  assign n5311 = n447 & ~n1424 ;
  assign n5323 = n333 & ~n723 ;
  assign n5324 = ~n5311 & ~n5323 ;
  assign n5325 = ~n5322 & n5324 ;
  assign n5326 = ~n5318 & n5325 ;
  assign n5327 = ~n5321 & n5326 ;
  assign n5328 = ~n5315 & n5327 ;
  assign n5329 = n292 & ~n5328 ;
  assign n5330 = ~n5310 & ~n5329 ;
  assign n5331 = \state_reg[0]/NET0131  & ~n5330 ;
  assign n5309 = n260 & n447 ;
  assign n5332 = ~n4910 & ~n5309 ;
  assign n5333 = ~n5331 & n5332 ;
  assign n5334 = \reg2_reg[17]/NET0131  & ~n2390 ;
  assign n5336 = \reg2_reg[17]/NET0131  & ~n1543 ;
  assign n5337 = n583 & n1543 ;
  assign n5338 = ~n5336 & ~n5337 ;
  assign n5339 = n588 & ~n5338 ;
  assign n5340 = ~n792 & n1543 ;
  assign n5341 = ~n5336 & ~n5340 ;
  assign n5342 = n798 & ~n5341 ;
  assign n5335 = n233 & n329 ;
  assign n5349 = n356 & n1543 ;
  assign n5350 = ~n5336 & ~n5349 ;
  assign n5351 = n910 & ~n5350 ;
  assign n5352 = ~n5335 & ~n5351 ;
  assign n5353 = ~n5342 & n5352 ;
  assign n5343 = n878 & n1543 ;
  assign n5344 = ~n5336 & ~n5343 ;
  assign n5345 = n881 & ~n5344 ;
  assign n5346 = n904 & n1543 ;
  assign n5347 = ~n5336 & ~n5346 ;
  assign n5348 = n907 & ~n5347 ;
  assign n5354 = ~n5345 & ~n5348 ;
  assign n5355 = n5353 & n5354 ;
  assign n5356 = ~n5339 & n5355 ;
  assign n5357 = n2389 & ~n5356 ;
  assign n5358 = ~n5334 & ~n5357 ;
  assign n5359 = \reg2_reg[2]/NET0131  & ~n2390 ;
  assign n5361 = \reg2_reg[2]/NET0131  & ~n1543 ;
  assign n5362 = n1543 & n3429 ;
  assign n5363 = ~n5361 & ~n5362 ;
  assign n5364 = n588 & ~n5363 ;
  assign n5365 = n1543 & ~n4004 ;
  assign n5360 = \reg3_reg[2]/NET0131  & n329 ;
  assign n5366 = ~n881 & n3033 ;
  assign n5367 = n5361 & ~n5366 ;
  assign n5368 = ~n5360 & ~n5367 ;
  assign n5369 = ~n5365 & n5368 ;
  assign n5370 = ~n5364 & n5369 ;
  assign n5371 = n2389 & ~n5370 ;
  assign n5372 = ~n5359 & ~n5371 ;
  assign n5373 = \reg2_reg[21]/NET0131  & ~n2390 ;
  assign n5376 = \reg2_reg[21]/NET0131  & ~n1543 ;
  assign n5377 = n1543 & n3992 ;
  assign n5378 = ~n5376 & ~n5377 ;
  assign n5379 = n588 & ~n5378 ;
  assign n5375 = n1543 & ~n3987 ;
  assign n5374 = n329 & n1010 ;
  assign n5380 = ~n4411 & n5376 ;
  assign n5381 = ~n5374 & ~n5380 ;
  assign n5382 = ~n5375 & n5381 ;
  assign n5383 = ~n5379 & n5382 ;
  assign n5384 = n2389 & ~n5383 ;
  assign n5385 = ~n5373 & ~n5384 ;
  assign n5386 = \reg2_reg[26]/NET0131  & ~n2390 ;
  assign n5388 = \reg2_reg[26]/NET0131  & ~n1543 ;
  assign n5389 = n1543 & ~n2435 ;
  assign n5390 = ~n5388 & ~n5389 ;
  assign n5391 = n881 & ~n5390 ;
  assign n5392 = n1543 & n2443 ;
  assign n5393 = ~n5388 & ~n5392 ;
  assign n5394 = n588 & ~n5393 ;
  assign n5395 = n1543 & n2452 ;
  assign n5396 = ~n5388 & ~n5395 ;
  assign n5397 = n907 & ~n5396 ;
  assign n5398 = n1543 & ~n2484 ;
  assign n5399 = ~n5388 & ~n5398 ;
  assign n5400 = n798 & ~n5399 ;
  assign n5387 = n329 & n958 ;
  assign n5401 = n953 & n1543 ;
  assign n5402 = ~n5388 & ~n5401 ;
  assign n5403 = n910 & ~n5402 ;
  assign n5404 = ~n5387 & ~n5403 ;
  assign n5405 = ~n5400 & n5404 ;
  assign n5406 = ~n5397 & n5405 ;
  assign n5407 = ~n5394 & n5406 ;
  assign n5408 = ~n5391 & n5407 ;
  assign n5409 = n2389 & ~n5408 ;
  assign n5410 = ~n5386 & ~n5409 ;
  assign n5411 = \reg1_reg[18]/NET0131  & ~n1497 ;
  assign n5412 = ~n2790 & n3212 ;
  assign n5413 = ~n5411 & ~n5412 ;
  assign n5414 = n881 & ~n5413 ;
  assign n5415 = n588 & n2798 ;
  assign n5416 = n3628 & ~n5415 ;
  assign n5417 = n3212 & ~n5416 ;
  assign n5418 = n2019 & n2389 ;
  assign n5419 = \reg1_reg[18]/NET0131  & ~n5418 ;
  assign n5420 = ~n5417 & ~n5419 ;
  assign n5421 = ~n5414 & n5420 ;
  assign n5422 = ~n289 & n4471 ;
  assign n5423 = n588 & n5422 ;
  assign n5424 = ~n259 & ~n5423 ;
  assign n5425 = \state_reg[0]/NET0131  & ~n5424 ;
  assign n5426 = \B_reg/NET0131  & ~n5425 ;
  assign n5521 = ~n987 & n1385 ;
  assign n5522 = n964 & ~n5521 ;
  assign n5523 = ~n1120 & ~n5522 ;
  assign n5448 = ~n1028 & n1390 ;
  assign n5449 = n1003 & ~n5448 ;
  assign n5450 = ~n1113 & ~n5449 ;
  assign n5434 = n632 & ~n1097 ;
  assign n5435 = n1074 & ~n5434 ;
  assign n5436 = ~n636 & ~n5435 ;
  assign n5437 = n678 & ~n1101 ;
  assign n5438 = n1057 & ~n5437 ;
  assign n5439 = ~n682 & ~n5438 ;
  assign n5440 = ~n5436 & ~n5439 ;
  assign n5525 = n1063 & ~n5440 ;
  assign n5526 = ~n748 & n4254 ;
  assign n5527 = n763 & ~n5526 ;
  assign n5528 = n775 & ~n5527 ;
  assign n5529 = n779 & ~n5528 ;
  assign n5530 = n1087 & ~n5529 ;
  assign n5531 = n725 & ~n5530 ;
  assign n5532 = n1081 & ~n5531 ;
  assign n5533 = n632 & n637 ;
  assign n5534 = ~n682 & n730 ;
  assign n5535 = n5533 & n5534 ;
  assign n5536 = n678 & n5535 ;
  assign n5537 = ~n5532 & n5536 ;
  assign n5538 = ~n5525 & ~n5537 ;
  assign n5539 = n1066 & ~n1070 ;
  assign n5540 = ~n5538 & n5539 ;
  assign n5524 = ~n1055 & n1372 ;
  assign n5541 = n1053 & ~n5524 ;
  assign n5542 = ~n5540 & n5541 ;
  assign n5543 = ~n1113 & n1387 ;
  assign n5544 = n1390 & n5543 ;
  assign n5545 = ~n5542 & n5544 ;
  assign n5546 = ~n5450 & ~n5545 ;
  assign n5547 = n1121 & n1124 ;
  assign n5548 = ~n5546 & n5547 ;
  assign n5549 = ~n5523 & ~n5548 ;
  assign n5430 = ~n2103 & ~n2159 ;
  assign n5427 = ~n2092 & ~n2403 ;
  assign n5469 = n415 & n2393 ;
  assign n5470 = ~n5427 & ~n5469 ;
  assign n5550 = n5430 & n5470 ;
  assign n5551 = ~n5549 & n5550 ;
  assign n5458 = ~n415 & ~n2393 ;
  assign n5471 = n2092 & n2403 ;
  assign n5475 = ~n5458 & ~n5471 ;
  assign n5432 = ~n2102 & ~n2150 ;
  assign n5552 = ~n2103 & ~n5427 ;
  assign n5553 = ~n5432 & n5552 ;
  assign n5554 = n5475 & ~n5553 ;
  assign n5555 = ~n5469 & ~n5554 ;
  assign n5556 = ~n5551 & ~n5555 ;
  assign n5558 = n327 & ~n5556 ;
  assign n5557 = ~n327 & n5556 ;
  assign n5559 = n586 & ~n5557 ;
  assign n5560 = ~n5558 & n5559 ;
  assign n5428 = ~n415 & ~n5427 ;
  assign n5429 = n2393 & ~n5428 ;
  assign n5431 = ~n2102 & ~n5430 ;
  assign n5433 = n1030 & n1056 ;
  assign n5441 = ~n717 & n2211 ;
  assign n5442 = n1081 & ~n5441 ;
  assign n5443 = ~n729 & ~n1814 ;
  assign n5444 = ~n5442 & n5443 ;
  assign n5445 = n5440 & ~n5444 ;
  assign n5446 = n1063 & ~n5445 ;
  assign n5447 = n5433 & ~n5446 ;
  assign n5451 = n1073 & n1117 ;
  assign n5452 = n988 & ~n5450 ;
  assign n5453 = ~n5451 & n5452 ;
  assign n5454 = ~n1128 & ~n5453 ;
  assign n5455 = ~n5447 & n5454 ;
  assign n5456 = n5432 & ~n5455 ;
  assign n5457 = ~n5431 & ~n5456 ;
  assign n5459 = ~n415 & ~n2092 ;
  assign n5460 = n2403 & ~n5459 ;
  assign n5461 = ~n5458 & ~n5460 ;
  assign n5462 = ~n5457 & n5461 ;
  assign n5463 = ~n5429 & ~n5462 ;
  assign n5465 = n327 & n5463 ;
  assign n5464 = ~n327 & ~n5463 ;
  assign n5466 = n318 & n322 ;
  assign n5467 = ~n5464 & n5466 ;
  assign n5468 = ~n5465 & n5467 ;
  assign n5472 = n5431 & ~n5471 ;
  assign n5473 = n5470 & ~n5472 ;
  assign n5474 = ~n5458 & ~n5473 ;
  assign n5476 = ~n2262 & n5433 ;
  assign n5477 = n5454 & ~n5476 ;
  assign n5478 = n5432 & n5475 ;
  assign n5479 = ~n5477 & n5478 ;
  assign n5480 = ~n5474 & ~n5479 ;
  assign n5483 = n3403 & n5480 ;
  assign n5481 = ~n318 & n328 ;
  assign n5482 = ~n5480 & n5481 ;
  assign n5484 = \B_reg/NET0131  & ~n312 ;
  assign n5503 = ~n1781 & ~n1844 ;
  assign n5504 = n2261 & ~n2349 ;
  assign n5507 = n5503 & n5504 ;
  assign n5486 = ~n2319 & n3082 ;
  assign n5487 = n3381 & n3411 ;
  assign n5494 = n5486 & n5487 ;
  assign n5485 = ~n1651 & ~n1697 ;
  assign n5495 = ~n592 & n5485 ;
  assign n5501 = n5494 & n5495 ;
  assign n5490 = n3849 & n4030 ;
  assign n5491 = n4255 & ~n4395 ;
  assign n5492 = n5490 & n5491 ;
  assign n5488 = ~n3457 & n3527 ;
  assign n5489 = ~n3600 & ~n3697 ;
  assign n5493 = n5488 & n5489 ;
  assign n5502 = n5492 & n5493 ;
  assign n5508 = n5501 & n5502 ;
  assign n5511 = n5507 & n5508 ;
  assign n5505 = ~n2829 & ~n2884 ;
  assign n5506 = ~n3973 & n5505 ;
  assign n5512 = ~n1349 & n5506 ;
  assign n5513 = n5511 & n5512 ;
  assign n5498 = ~n2787 & n5470 ;
  assign n5499 = n5475 & n5498 ;
  assign n5496 = ~n1603 & ~n1739 ;
  assign n5497 = n2104 & n2216 ;
  assign n5500 = n5496 & n5497 ;
  assign n5509 = n5499 & n5500 ;
  assign n5510 = ~n2416 & n5509 ;
  assign n5514 = ~n1141 & n5510 ;
  assign n5515 = n5513 & n5514 ;
  assign n5517 = ~n327 & ~n5515 ;
  assign n5516 = n327 & n5515 ;
  assign n5518 = ~n318 & n322 ;
  assign n5519 = ~n5516 & n5518 ;
  assign n5520 = ~n5517 & n5519 ;
  assign n5561 = ~n5484 & ~n5520 ;
  assign n5562 = ~n5482 & n5561 ;
  assign n5563 = ~n5483 & n5562 ;
  assign n5564 = ~n5468 & n5563 ;
  assign n5565 = ~n5560 & n5564 ;
  assign n5566 = n260 & ~n5565 ;
  assign n5567 = ~n5426 & ~n5566 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g22/_0_  = ~n923 ;
  assign \g32_dup/_0_  = ~n934 ;
  assign \g35904/_0_  = ~n1303 ;
  assign \g35905/_0_  = ~n1443 ;
  assign \g35906/_0_  = ~n1473 ;
  assign \g35907/_0_  = ~n1496 ;
  assign \g35908/_0_  = ~n1519 ;
  assign \g35909/_0_  = ~n1542 ;
  assign \g35910/_0_  = ~n1573 ;
  assign \g35911/_0_  = ~n1597 ;
  assign \g35932/_0_  = ~n1645 ;
  assign \g35955/_0_  = ~n1690 ;
  assign \g35956/_0_  = ~n1733 ;
  assign \g35957/_0_  = ~n1776 ;
  assign \g35962/_0_  = ~n1839 ;
  assign \g35967/_0_  = ~n1893 ;
  assign \g35968/_0_  = ~n1920 ;
  assign \g35971/_0_  = ~n1945 ;
  assign \g35972/_0_  = ~n1969 ;
  assign \g35973/_0_  = ~n1991 ;
  assign \g35974/_0_  = ~n2013 ;
  assign \g35975/_0_  = ~n2030 ;
  assign \g35976/_0_  = ~n2056 ;
  assign \g35977/_0_  = ~n2080 ;
  assign \g35978/_0_  = ~n2191 ;
  assign \g36015/_0_  = ~n2255 ;
  assign \g36016/_0_  = ~n2300 ;
  assign \g36018/_0_  = ~n2343 ;
  assign \g36022/_0_  = ~n2387 ;
  assign \g36023/_0_  = ~n2414 ;
  assign \g36025/_0_  = ~n2500 ;
  assign \g36029/_0_  = ~n2520 ;
  assign \g36030/_0_  = ~n2545 ;
  assign \g36031/_0_  = ~n2571 ;
  assign \g36032/_0_  = ~n2598 ;
  assign \g36033/_0_  = ~n2616 ;
  assign \g36034/_0_  = ~n2638 ;
  assign \g36035/_0_  = ~n2661 ;
  assign \g36036/_0_  = ~n2687 ;
  assign \g36038/_0_  = ~n2715 ;
  assign \g36039/_0_  = ~n2733 ;
  assign \g36040/_0_  = ~n2757 ;
  assign \g36041/_0_  = ~n2783 ;
  assign \g36073/_0_  = ~n2825 ;
  assign \g36087/_0_  = ~n2882 ;
  assign \g36091/_0_  = ~n2931 ;
  assign \g36092/_0_  = ~n2953 ;
  assign \g36093/_0_  = ~n2978 ;
  assign \g36094/_0_  = ~n3004 ;
  assign \g36096/_0_  = ~n3024 ;
  assign \g36097/_0_  = ~n3045 ;
  assign \g36098/_0_  = ~n3052 ;
  assign \g36099/_0_  = ~n3055 ;
  assign \g36100/_0_  = ~n3077 ;
  assign \g36101/_0_  = ~n3119 ;
  assign \g36102/_0_  = ~n3146 ;
  assign \g36103/_0_  = ~n3171 ;
  assign \g36104/_0_  = ~n3193 ;
  assign \g36105/_0_  = ~n3211 ;
  assign \g36106/_0_  = ~n3216 ;
  assign \g36107/_0_  = ~n3226 ;
  assign \g36108/_0_  = ~n3248 ;
  assign \g36109/_0_  = ~n3274 ;
  assign \g36110/_0_  = ~n3298 ;
  assign \g36111/_0_  = ~n3322 ;
  assign \g36112/_0_  = ~n3343 ;
  assign \g36113/_0_  = ~n3365 ;
  assign \g36165/_0_  = ~n3399 ;
  assign \g36169/_0_  = ~n3443 ;
  assign \g36170/_0_  = ~n3484 ;
  assign \g36171/_0_  = ~n3512 ;
  assign \g36172/_0_  = ~n3555 ;
  assign \g36198/_0_  = ~n3583 ;
  assign \g36199/_0_  = ~n3626 ;
  assign \g36200/_0_  = ~n3646 ;
  assign \g36201/_0_  = ~n3672 ;
  assign \g36202/_0_  = ~n3692 ;
  assign \g36203/_0_  = ~n3729 ;
  assign \g36205/_0_  = ~n3755 ;
  assign \g36206/_0_  = ~n3773 ;
  assign \g36207/_0_  = ~n3795 ;
  assign \g36208/_0_  = ~n3813 ;
  assign \g36209/_0_  = ~n3833 ;
  assign \g36240/_0_  = ~n3874 ;
  assign \g36281/_0_  = ~n3900 ;
  assign \g36282/_0_  = ~n3928 ;
  assign \g36283/_0_  = ~n3955 ;
  assign \g36284/_0_  = ~n3965 ;
  assign \g36285/_0_  = ~n4000 ;
  assign \g36286/_0_  = ~n4009 ;
  assign \g36287/_0_  = ~n4017 ;
  assign \g36288/_0_  = ~n4056 ;
  assign \g36289/_0_  = ~n4078 ;
  assign \g36290/_0_  = ~n4105 ;
  assign \g36291/_0_  = ~n4131 ;
  assign \g36292/_0_  = ~n4137 ;
  assign \g36293/_0_  = ~n4143 ;
  assign \g36294/_0_  = ~n4149 ;
  assign \g36295/_0_  = ~n4171 ;
  assign \g36296/_0_  = ~n4193 ;
  assign \g36297/_0_  = ~n4219 ;
  assign \g36298/_0_  = ~n4245 ;
  assign \g36330/_0_  = ~n4267 ;
  assign \g36385/_0_  = ~n4286 ;
  assign \g36390/_0_  = ~n4299 ;
  assign \g36391/_0_  = ~n4323 ;
  assign \g36392/_0_  = ~n4351 ;
  assign \g36393/_0_  = ~n4360 ;
  assign \g36394/_0_  = ~n4378 ;
  assign \g36470/_0_  = ~n4382 ;
  assign \g36471/_0_  = ~n4420 ;
  assign \g36472/_0_  = n4433 ;
  assign \g36473/_0_  = ~n4445 ;
  assign \g36474/_0_  = ~n4460 ;
  assign \g36475/_0_  = ~n4463 ;
  assign \g38/_0_  = ~n546 ;
  assign \g38399/_0_  = n4516 ;
  assign \g38400/_0_  = n4555 ;
  assign \g39639/_0_  = ~n4642 ;
  assign \g39641/_0_  = ~n4687 ;
  assign \g39644/_0_  = ~n4720 ;
  assign \g39647/_0_  = ~n4752 ;
  assign \g39648/_0_  = ~n4790 ;
  assign \g39650/_0_  = ~n4832 ;
  assign \g39654/_0_  = ~n4866 ;
  assign \g39658/_0_  = ~n4887 ;
  assign \g39660/_0_  = ~n4908 ;
  assign \g39662/_0_  = ~n4929 ;
  assign \g39663/_0_  = ~n4949 ;
  assign \g39665/_0_  = ~n4971 ;
  assign \g39666/_0_  = ~n4992 ;
  assign \g39667/_0_  = ~n5013 ;
  assign \g39730/_0_  = ~n5036 ;
  assign \g39796/_0_  = ~n5038 ;
  assign \g39930/_0_  = ~n5048 ;
  assign \g39931/_0_  = ~n5069 ;
  assign \g39932/_0_  = ~n5091 ;
  assign \g40045/_0_  = ~n300 ;
  assign \g40150/u3_syn_4  = n2389 ;
  assign \g40608/_0_  = n307 ;
  assign \g41017/u3_syn_4  = n5092 ;
  assign \g42159/_0_  = ~n5095 ;
  assign \g42169/_0_  = ~n5098 ;
  assign \g42174/_0_  = ~n5101 ;
  assign \g42483/_0_  = ~n1279 ;
  assign \g42736/_0_  = ~n434 ;
  assign \g42746/_0_  = ~n526 ;
  assign \g42755/_0_  = ~n425 ;
  assign \g42767/_0_  = ~n389 ;
  assign \g42776/_0_  = ~n483 ;
  assign \g42871_dup/_1_  = ~n1014 ;
  assign \g42908/_0_  = ~n985 ;
  assign \g42938/_0_  = ~n513 ;
  assign \g42969/_0_  = ~n495 ;
  assign \g43022/_0_  = ~n1026 ;
  assign \g44035/_1__syn_2  = n1471 ;
  assign \g44227/_3_  = ~n5104 ;
  assign \g44260/_3_  = ~n5107 ;
  assign \g44261/_3_  = ~n5110 ;
  assign \g44262/_3_  = ~n5113 ;
  assign \g44311/_3_  = n5119 ;
  assign \g44378/_3_  = n5122 ;
  assign \g44379/_3_  = ~n5124 ;
  assign \g44383/_3_  = ~n5127 ;
  assign \g44384/_3_  = n5130 ;
  assign \g44385/_3_  = ~n5133 ;
  assign \g44386/_3_  = ~n5136 ;
  assign \g44390/_3_  = n5139 ;
  assign \g44391/_3_  = ~n5142 ;
  assign \g44492/_3_  = n5145 ;
  assign \g44493/_3_  = ~n5148 ;
  assign \g44494/_3_  = ~n5151 ;
  assign \g44495/_3_  = ~n5154 ;
  assign \g44496/_3_  = ~n5157 ;
  assign \g44497/_3_  = ~n5160 ;
  assign \g44498/_3_  = ~n5163 ;
  assign \g44499/_3_  = n5166 ;
  assign \g44575/_3_  = ~n5169 ;
  assign \g44589/_3_  = ~n5172 ;
  assign \g44596/_3_  = ~n5175 ;
  assign \g44615/_3_  = ~n5178 ;
  assign \g44795/_3_  = ~n5181 ;
  assign \g44803/_3_  = ~n5184 ;
  assign \g44804/_3_  = n5187 ;
  assign \g44888/_3_  = ~n5190 ;
  assign \g44889/_3_  = ~n5193 ;
  assign \g45004/_3_  = ~n5196 ;
  assign \g46129/_0_  = ~n396 ;
  assign \g46133/_0_  = ~n415 ;
  assign \g46265/_2_  = ~n454 ;
  assign \g46313/_0_  = ~n5221 ;
  assign \g46372/_0_  = ~n5246 ;
  assign \g46377/_0_  = ~n5271 ;
  assign \g46399/_0_  = ~n5283 ;
  assign \g46405/_0_  = ~n5308 ;
  assign \g46427/_0_  = ~n5333 ;
  assign \g46461/_0_  = ~n5358 ;
  assign \g46526/_0_  = ~n5372 ;
  assign \g46576/_0_  = ~n555 ;
  assign \g46608/_0_  = ~n382 ;
  assign \g46697/_0_  = ~n1001 ;
  assign \g46778/_0_  = ~n445 ;
  assign \g47007/_0_  = ~n474 ;
  assign \g47023/_0_  = ~n5385 ;
  assign \g47077/_1_  = ~n576 ;
  assign \g47097/_0_  = ~n1048 ;
  assign \g47109/_1_  = ~n962 ;
  assign \g47142_dup/_1_  = ~n504 ;
  assign \g47256/_0_  = ~n951 ;
  assign \g47328/_0_  = ~n5410 ;
  assign \g47373/_0_  = ~n5421 ;
  assign \g47465/_0_  = ~n2092 ;
  assign \g47518/_0_  = ~n5567 ;
  assign \g47556/_1_  = ~n974 ;
  assign \g56/_0_  = ~n566 ;
  assign \state_reg[0]/NET0131_syn_2  = ~\state_reg[0]/NET0131  ;
endmodule
