module top (\C_0_pad , \C_10_pad , \C_11_pad , \C_12_pad , \C_13_pad , \C_14_pad , \C_15_pad , \C_16_pad , \C_17_pad , \C_18_pad , \C_19_pad , \C_1_pad , \C_20_pad , \C_21_pad , \C_22_pad , \C_23_pad , \C_24_pad , \C_25_pad , \C_26_pad , \C_27_pad , \C_28_pad , \C_29_pad , \C_2_pad , \C_30_pad , \C_31_pad , \C_32_pad , \C_3_pad , \C_4_pad , \C_5_pad , \C_6_pad , \C_7_pad , \C_8_pad , \C_9_pad , \P_0_pad , \X_10_reg/NET0131 , \X_11_reg/NET0131 , \X_12_reg/NET0131 , \X_13_reg/NET0131 , \X_14_reg/NET0131 , \X_15_reg/NET0131 , \X_16_reg/NET0131 , \X_17_reg/NET0131 , \X_18_reg/NET0131 , \X_19_reg/NET0131 , \X_1_reg/NET0131 , \X_20_reg/NET0131 , \X_21_reg/NET0131 , \X_22_reg/NET0131 , \X_23_reg/NET0131 , \X_24_reg/NET0131 , \X_25_reg/NET0131 , \X_26_reg/NET0131 , \X_27_reg/NET0131 , \X_28_reg/NET0131 , \X_29_reg/NET0131 , \X_2_reg/NET0131 , \X_30_reg/P0002 , \X_31_reg/P0002 , \X_32_reg/P0002 , \X_3_reg/NET0131 , \X_4_reg/NET0131 , \X_5_reg/NET0131 , \X_6_reg/NET0131 , \X_7_reg/NET0131 , \X_8_reg/NET0131 , \X_9_reg/NET0131 , \X_30_reg/P0000 , \X_31_reg/P0000 , \X_32_reg/P0000 , Z_pad, \_al_n0 , \_al_n1 , \g1375/_1_ , \g1387/_0_ , \g1398/_0_ , \g1400/_0_ , \g1419/_0_ , \g1433/_0_ , \g1443/_0_ , \g1457/_0_ , \g1458/_0_ , \g1468/_0_ , \g1483/_0_ , \g1486/_0_ , \g1493/_0_ , \g1504/_0_ , \g1505/_0_ , \g1512/_0_ , \g1525/_0_ , \g1535/_0_ , \g1544/_0_ , \g1565/_0_ , \g1871/_0_ , \g1900/_0_ , \g1955/_0_ , \g1961/_0_ , \g1991/_0_ , \g2026/_0_ , \g2040/_0_ , \g2046/_0_ , \g2051/_1_ , \g2098/_0_ , \g21/_0_ , \g2101/_0_ );
	input \C_0_pad  ;
	input \C_10_pad  ;
	input \C_11_pad  ;
	input \C_12_pad  ;
	input \C_13_pad  ;
	input \C_14_pad  ;
	input \C_15_pad  ;
	input \C_16_pad  ;
	input \C_17_pad  ;
	input \C_18_pad  ;
	input \C_19_pad  ;
	input \C_1_pad  ;
	input \C_20_pad  ;
	input \C_21_pad  ;
	input \C_22_pad  ;
	input \C_23_pad  ;
	input \C_24_pad  ;
	input \C_25_pad  ;
	input \C_26_pad  ;
	input \C_27_pad  ;
	input \C_28_pad  ;
	input \C_29_pad  ;
	input \C_2_pad  ;
	input \C_30_pad  ;
	input \C_31_pad  ;
	input \C_32_pad  ;
	input \C_3_pad  ;
	input \C_4_pad  ;
	input \C_5_pad  ;
	input \C_6_pad  ;
	input \C_7_pad  ;
	input \C_8_pad  ;
	input \C_9_pad  ;
	input \P_0_pad  ;
	input \X_10_reg/NET0131  ;
	input \X_11_reg/NET0131  ;
	input \X_12_reg/NET0131  ;
	input \X_13_reg/NET0131  ;
	input \X_14_reg/NET0131  ;
	input \X_15_reg/NET0131  ;
	input \X_16_reg/NET0131  ;
	input \X_17_reg/NET0131  ;
	input \X_18_reg/NET0131  ;
	input \X_19_reg/NET0131  ;
	input \X_1_reg/NET0131  ;
	input \X_20_reg/NET0131  ;
	input \X_21_reg/NET0131  ;
	input \X_22_reg/NET0131  ;
	input \X_23_reg/NET0131  ;
	input \X_24_reg/NET0131  ;
	input \X_25_reg/NET0131  ;
	input \X_26_reg/NET0131  ;
	input \X_27_reg/NET0131  ;
	input \X_28_reg/NET0131  ;
	input \X_29_reg/NET0131  ;
	input \X_2_reg/NET0131  ;
	input \X_30_reg/P0002  ;
	input \X_31_reg/P0002  ;
	input \X_32_reg/P0002  ;
	input \X_3_reg/NET0131  ;
	input \X_4_reg/NET0131  ;
	input \X_5_reg/NET0131  ;
	input \X_6_reg/NET0131  ;
	input \X_7_reg/NET0131  ;
	input \X_8_reg/NET0131  ;
	input \X_9_reg/NET0131  ;
	output \X_30_reg/P0000  ;
	output \X_31_reg/P0000  ;
	output \X_32_reg/P0000  ;
	output Z_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1375/_1_  ;
	output \g1387/_0_  ;
	output \g1398/_0_  ;
	output \g1400/_0_  ;
	output \g1419/_0_  ;
	output \g1433/_0_  ;
	output \g1443/_0_  ;
	output \g1457/_0_  ;
	output \g1458/_0_  ;
	output \g1468/_0_  ;
	output \g1483/_0_  ;
	output \g1486/_0_  ;
	output \g1493/_0_  ;
	output \g1504/_0_  ;
	output \g1505/_0_  ;
	output \g1512/_0_  ;
	output \g1525/_0_  ;
	output \g1535/_0_  ;
	output \g1544/_0_  ;
	output \g1565/_0_  ;
	output \g1871/_0_  ;
	output \g1900/_0_  ;
	output \g1955/_0_  ;
	output \g1961/_0_  ;
	output \g1991/_0_  ;
	output \g2026/_0_  ;
	output \g2040/_0_  ;
	output \g2046/_0_  ;
	output \g2051/_1_  ;
	output \g2098/_0_  ;
	output \g21/_0_  ;
	output \g2101/_0_  ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w121_ ;
	wire _w119_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w75_ ;
	wire _w73_ ;
	wire _w71_ ;
	wire _w76_ ;
	wire _w122_ ;
	wire _w63_ ;
	wire _w190_ ;
	wire _w92_ ;
	wire _w74_ ;
	wire _w120_ ;
	wire _w61_ ;
	wire _w188_ ;
	wire _w90_ ;
	wire _w72_ ;
	wire _w118_ ;
	wire _w59_ ;
	wire _w186_ ;
	wire _w88_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w89_ ;
	wire _w91_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w187_ ;
	wire _w189_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\X_30_reg/P0002 ,
		_w59_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\X_31_reg/P0002 ,
		_w61_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\X_32_reg/P0002 ,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w71_
	);
	LUT3 #(
		.INIT('h01)
	) name4 (
		\X_4_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		\X_20_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		_w75_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		\X_19_reg/NET0131 ,
		\X_1_reg/NET0131 ,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w77_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\X_10_reg/NET0131 ,
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('h0001)
	) name11 (
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		\X_15_reg/NET0131 ,
		\X_16_reg/NET0131 ,
		_w79_
	);
	LUT4 #(
		.INIT('h8000)
	) name12 (
		_w78_,
		_w79_,
		_w74_,
		_w76_,
		_w80_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\C_21_pad ,
		\X_21_reg/NET0131 ,
		_w81_
	);
	LUT3 #(
		.INIT('h20)
	) name14 (
		\C_23_pad ,
		\X_22_reg/NET0131 ,
		\X_23_reg/NET0131 ,
		_w82_
	);
	LUT3 #(
		.INIT('h13)
	) name15 (
		\C_22_pad ,
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		_w83_
	);
	LUT3 #(
		.INIT('h45)
	) name16 (
		_w81_,
		_w82_,
		_w83_,
		_w84_
	);
	LUT3 #(
		.INIT('h80)
	) name17 (
		_w73_,
		_w80_,
		_w84_,
		_w85_
	);
	LUT3 #(
		.INIT('h01)
	) name18 (
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w86_
	);
	LUT3 #(
		.INIT('h80)
	) name19 (
		_w86_,
		_w71_,
		_w72_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\C_14_pad ,
		\X_14_reg/NET0131 ,
		_w88_
	);
	LUT4 #(
		.INIT('h0200)
	) name21 (
		\C_16_pad ,
		\X_14_reg/NET0131 ,
		\X_15_reg/NET0131 ,
		\X_16_reg/NET0131 ,
		_w89_
	);
	LUT4 #(
		.INIT('h4440)
	) name22 (
		\X_13_reg/NET0131 ,
		_w78_,
		_w88_,
		_w89_,
		_w90_
	);
	LUT4 #(
		.INIT('h0001)
	) name23 (
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\C_5_pad ,
		\X_5_reg/NET0131 ,
		_w92_
	);
	LUT3 #(
		.INIT('h15)
	) name25 (
		\C_0_pad ,
		_w91_,
		_w92_,
		_w93_
	);
	LUT3 #(
		.INIT('h70)
	) name26 (
		_w87_,
		_w90_,
		_w93_,
		_w94_
	);
	LUT3 #(
		.INIT('h8a)
	) name27 (
		\P_0_pad ,
		_w85_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		_w96_
	);
	LUT4 #(
		.INIT('h0800)
	) name29 (
		\C_24_pad ,
		\P_0_pad ,
		\X_23_reg/NET0131 ,
		\X_24_reg/NET0131 ,
		_w97_
	);
	LUT4 #(
		.INIT('h8000)
	) name30 (
		_w73_,
		_w80_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h8000)
	) name31 (
		\P_0_pad ,
		_w86_,
		_w71_,
		_w72_,
		_w99_
	);
	LUT4 #(
		.INIT('h535f)
	) name32 (
		\C_11_pad ,
		\C_12_pad ,
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		_w100_
	);
	LUT4 #(
		.INIT('h335f)
	) name33 (
		\C_10_pad ,
		\C_9_pad ,
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w101_
	);
	LUT3 #(
		.INIT('hd0)
	) name34 (
		_w77_,
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w99_,
		_w102_,
		_w103_
	);
	LUT3 #(
		.INIT('h20)
	) name36 (
		\C_8_pad ,
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w104_
	);
	LUT3 #(
		.INIT('h13)
	) name37 (
		\C_7_pad ,
		\X_6_reg/NET0131 ,
		\X_7_reg/NET0131 ,
		_w105_
	);
	LUT4 #(
		.INIT('h080c)
	) name38 (
		\C_6_pad ,
		\P_0_pad ,
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w106_
	);
	LUT4 #(
		.INIT('h8a00)
	) name39 (
		_w91_,
		_w104_,
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\C_2_pad ,
		\X_2_reg/NET0131 ,
		_w109_
	);
	LUT4 #(
		.INIT('h0200)
	) name42 (
		\C_4_pad ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w110_
	);
	LUT3 #(
		.INIT('ha8)
	) name43 (
		_w108_,
		_w109_,
		_w110_,
		_w111_
	);
	LUT3 #(
		.INIT('h80)
	) name44 (
		\C_1_pad ,
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w112_
	);
	LUT3 #(
		.INIT('h20)
	) name45 (
		\C_3_pad ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w113_
	);
	LUT3 #(
		.INIT('h13)
	) name46 (
		_w108_,
		_w112_,
		_w113_,
		_w114_
	);
	LUT3 #(
		.INIT('h10)
	) name47 (
		_w111_,
		_w107_,
		_w114_,
		_w115_
	);
	LUT3 #(
		.INIT('h10)
	) name48 (
		_w103_,
		_w98_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\C_17_pad ,
		\X_17_reg/NET0131 ,
		_w117_
	);
	LUT4 #(
		.INIT('h535f)
	) name50 (
		\C_19_pad ,
		\C_20_pad ,
		\X_19_reg/NET0131 ,
		\X_20_reg/NET0131 ,
		_w118_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name51 (
		_w79_,
		_w75_,
		_w117_,
		_w118_,
		_w119_
	);
	LUT3 #(
		.INIT('h20)
	) name52 (
		\C_18_pad ,
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\C_13_pad ,
		\X_13_reg/NET0131 ,
		_w121_
	);
	LUT4 #(
		.INIT('h0200)
	) name54 (
		\C_15_pad ,
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		\X_15_reg/NET0131 ,
		_w122_
	);
	LUT4 #(
		.INIT('h0103)
	) name55 (
		_w79_,
		_w121_,
		_w122_,
		_w120_,
		_w123_
	);
	LUT4 #(
		.INIT('h8a00)
	) name56 (
		_w78_,
		_w119_,
		_w123_,
		_w99_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\C_25_pad ,
		\X_25_reg/NET0131 ,
		_w125_
	);
	LUT3 #(
		.INIT('h20)
	) name58 (
		\C_28_pad ,
		\X_27_reg/NET0131 ,
		\X_28_reg/NET0131 ,
		_w126_
	);
	LUT3 #(
		.INIT('h13)
	) name59 (
		\C_27_pad ,
		\X_26_reg/NET0131 ,
		\X_27_reg/NET0131 ,
		_w127_
	);
	LUT3 #(
		.INIT('h23)
	) name60 (
		\C_26_pad ,
		\X_25_reg/NET0131 ,
		\X_26_reg/NET0131 ,
		_w128_
	);
	LUT4 #(
		.INIT('h1055)
	) name61 (
		_w125_,
		_w126_,
		_w127_,
		_w128_,
		_w129_
	);
	LUT4 #(
		.INIT('h535f)
	) name62 (
		\C_31_pad ,
		\C_32_pad ,
		\X_31_reg/P0002 ,
		\X_32_reg/P0002 ,
		_w130_
	);
	LUT3 #(
		.INIT('h13)
	) name63 (
		\C_30_pad ,
		\X_29_reg/NET0131 ,
		\X_30_reg/P0002 ,
		_w131_
	);
	LUT3 #(
		.INIT('he0)
	) name64 (
		\X_30_reg/P0002 ,
		_w130_,
		_w131_,
		_w132_
	);
	LUT3 #(
		.INIT('h01)
	) name65 (
		\X_26_reg/NET0131 ,
		\X_27_reg/NET0131 ,
		\X_28_reg/NET0131 ,
		_w133_
	);
	LUT4 #(
		.INIT('h080c)
	) name66 (
		\C_29_pad ,
		\P_0_pad ,
		\X_25_reg/NET0131 ,
		\X_29_reg/NET0131 ,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name68 (
		\P_0_pad ,
		_w129_,
		_w132_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\X_23_reg/NET0131 ,
		\X_24_reg/NET0131 ,
		_w137_
	);
	LUT4 #(
		.INIT('h8000)
	) name70 (
		_w73_,
		_w80_,
		_w96_,
		_w137_,
		_w138_
	);
	LUT3 #(
		.INIT('h45)
	) name71 (
		_w124_,
		_w136_,
		_w138_,
		_w139_
	);
	LUT3 #(
		.INIT('hbf)
	) name72 (
		_w95_,
		_w116_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w141_
	);
	LUT4 #(
		.INIT('h8000)
	) name74 (
		\X_10_reg/NET0131 ,
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w142_
	);
	LUT4 #(
		.INIT('h8000)
	) name75 (
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT3 #(
		.INIT('h80)
	) name77 (
		\X_14_reg/NET0131 ,
		\X_15_reg/NET0131 ,
		\X_16_reg/NET0131 ,
		_w145_
	);
	LUT3 #(
		.INIT('h80)
	) name78 (
		\X_20_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		_w147_
	);
	LUT4 #(
		.INIT('h8000)
	) name80 (
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		\X_19_reg/NET0131 ,
		\X_1_reg/NET0131 ,
		_w148_
	);
	LUT3 #(
		.INIT('h80)
	) name81 (
		_w145_,
		_w146_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		_w150_
	);
	LUT3 #(
		.INIT('h80)
	) name83 (
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		\X_23_reg/NET0131 ,
		_w151_
	);
	LUT4 #(
		.INIT('h8000)
	) name84 (
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		\X_23_reg/NET0131 ,
		\X_24_reg/NET0131 ,
		_w152_
	);
	LUT3 #(
		.INIT('h80)
	) name85 (
		\P_0_pad ,
		\X_13_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w153_
	);
	LUT4 #(
		.INIT('h8000)
	) name86 (
		\P_0_pad ,
		\X_13_reg/NET0131 ,
		\X_25_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w152_,
		_w154_,
		_w155_
	);
	LUT3 #(
		.INIT('h80)
	) name88 (
		_w144_,
		_w149_,
		_w155_,
		_w156_
	);
	LUT4 #(
		.INIT('h8000)
	) name89 (
		\X_26_reg/NET0131 ,
		_w144_,
		_w149_,
		_w155_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\X_27_reg/NET0131 ,
		\X_28_reg/NET0131 ,
		_w158_
	);
	LUT3 #(
		.INIT('h80)
	) name91 (
		\X_29_reg/NET0131 ,
		_w157_,
		_w158_,
		_w159_
	);
	LUT4 #(
		.INIT('h8000)
	) name92 (
		\X_29_reg/NET0131 ,
		\X_30_reg/P0002 ,
		_w157_,
		_w158_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\X_31_reg/P0002 ,
		_w160_,
		_w161_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name94 (
		\X_26_reg/NET0131 ,
		_w144_,
		_w149_,
		_w155_,
		_w162_
	);
	LUT3 #(
		.INIT('h80)
	) name95 (
		_w144_,
		_w149_,
		_w153_,
		_w163_
	);
	LUT3 #(
		.INIT('h6c)
	) name96 (
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h6)
	) name97 (
		\X_27_reg/NET0131 ,
		_w157_,
		_w165_
	);
	LUT3 #(
		.INIT('h6a)
	) name98 (
		\X_23_reg/NET0131 ,
		_w150_,
		_w163_,
		_w166_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name99 (
		\X_21_reg/NET0131 ,
		_w144_,
		_w149_,
		_w153_,
		_w167_
	);
	LUT4 #(
		.INIT('h8000)
	) name100 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w168_
	);
	LUT4 #(
		.INIT('h8000)
	) name101 (
		\X_4_reg/NET0131 ,
		_w142_,
		_w143_,
		_w168_,
		_w169_
	);
	LUT3 #(
		.INIT('h80)
	) name102 (
		\X_13_reg/NET0131 ,
		_w145_,
		_w169_,
		_w170_
	);
	LUT4 #(
		.INIT('h8000)
	) name103 (
		\X_13_reg/NET0131 ,
		_w145_,
		_w147_,
		_w169_,
		_w171_
	);
	LUT2 #(
		.INIT('h6)
	) name104 (
		\X_19_reg/NET0131 ,
		_w171_,
		_w172_
	);
	LUT4 #(
		.INIT('h8000)
	) name105 (
		\X_4_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w168_,
		_w173_
	);
	LUT4 #(
		.INIT('h1333)
	) name106 (
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		_w142_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w169_,
		_w174_,
		_w175_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name108 (
		\X_13_reg/NET0131 ,
		\X_17_reg/NET0131 ,
		_w145_,
		_w169_,
		_w176_
	);
	LUT4 #(
		.INIT('h8000)
	) name109 (
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		\X_15_reg/NET0131 ,
		_w169_,
		_w177_
	);
	LUT4 #(
		.INIT('h78f0)
	) name110 (
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		\X_15_reg/NET0131 ,
		_w169_,
		_w178_
	);
	LUT2 #(
		.INIT('h6)
	) name111 (
		\X_13_reg/NET0131 ,
		_w169_,
		_w179_
	);
	LUT4 #(
		.INIT('h78f0)
	) name112 (
		\X_4_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w168_,
		_w180_
	);
	LUT3 #(
		.INIT('h6a)
	) name113 (
		\X_11_reg/NET0131 ,
		_w142_,
		_w173_,
		_w181_
	);
	LUT2 #(
		.INIT('h6)
	) name114 (
		\X_4_reg/NET0131 ,
		_w168_,
		_w182_
	);
	LUT3 #(
		.INIT('h6a)
	) name115 (
		\X_9_reg/NET0131 ,
		_w141_,
		_w173_,
		_w183_
	);
	LUT2 #(
		.INIT('h6)
	) name116 (
		\X_7_reg/NET0131 ,
		_w173_,
		_w184_
	);
	LUT3 #(
		.INIT('h6c)
	) name117 (
		\X_4_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		_w168_,
		_w185_
	);
	LUT4 #(
		.INIT('h7f80)
	) name118 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w186_
	);
	LUT3 #(
		.INIT('h78)
	) name119 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w187_
	);
	LUT2 #(
		.INIT('h6)
	) name120 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w188_
	);
	LUT3 #(
		.INIT('h6c)
	) name121 (
		\X_19_reg/NET0131 ,
		\X_20_reg/NET0131 ,
		_w171_,
		_w189_
	);
	LUT3 #(
		.INIT('h6c)
	) name122 (
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		_w169_,
		_w190_
	);
	LUT3 #(
		.INIT('h6c)
	) name123 (
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		_w170_,
		_w191_
	);
	LUT4 #(
		.INIT('h8000)
	) name124 (
		_w144_,
		_w149_,
		_w153_,
		_w152_,
		_w192_
	);
	LUT3 #(
		.INIT('h6a)
	) name125 (
		\X_24_reg/NET0131 ,
		_w151_,
		_w163_,
		_w193_
	);
	LUT3 #(
		.INIT('h32)
	) name126 (
		\X_25_reg/NET0131 ,
		_w156_,
		_w192_,
		_w194_
	);
	LUT3 #(
		.INIT('h6a)
	) name127 (
		\X_29_reg/NET0131 ,
		_w157_,
		_w158_,
		_w195_
	);
	LUT3 #(
		.INIT('h6c)
	) name128 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w173_,
		_w196_
	);
	LUT3 #(
		.INIT('h6c)
	) name129 (
		\X_27_reg/NET0131 ,
		\X_28_reg/NET0131 ,
		_w157_,
		_w197_
	);
	LUT3 #(
		.INIT('h32)
	) name130 (
		\X_16_reg/NET0131 ,
		_w170_,
		_w177_,
		_w198_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name131 (
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w141_,
		_w173_,
		_w199_
	);
	assign \X_30_reg/P0000  = _w59_ ;
	assign \X_31_reg/P0000  = _w61_ ;
	assign \X_32_reg/P0000  = _w63_ ;
	assign Z_pad = _w140_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1375/_1_  = _w161_ ;
	assign \g1387/_0_  = _w162_ ;
	assign \g1398/_0_  = _w164_ ;
	assign \g1400/_0_  = _w165_ ;
	assign \g1419/_0_  = _w166_ ;
	assign \g1433/_0_  = _w167_ ;
	assign \g1443/_0_  = _w172_ ;
	assign \g1457/_0_  = _w175_ ;
	assign \g1458/_0_  = _w176_ ;
	assign \g1468/_0_  = _w178_ ;
	assign \g1483/_0_  = _w179_ ;
	assign \g1486/_0_  = _w180_ ;
	assign \g1493/_0_  = _w181_ ;
	assign \g1504/_0_  = _w182_ ;
	assign \g1505/_0_  = _w183_ ;
	assign \g1512/_0_  = _w184_ ;
	assign \g1525/_0_  = _w185_ ;
	assign \g1535/_0_  = _w186_ ;
	assign \g1544/_0_  = _w187_ ;
	assign \g1565/_0_  = _w188_ ;
	assign \g1871/_0_  = _w189_ ;
	assign \g1900/_0_  = _w190_ ;
	assign \g1955/_0_  = _w191_ ;
	assign \g1961/_0_  = _w193_ ;
	assign \g1991/_0_  = _w194_ ;
	assign \g2026/_0_  = _w195_ ;
	assign \g2040/_0_  = _w196_ ;
	assign \g2046/_0_  = _w160_ ;
	assign \g2051/_1_  = _w159_ ;
	assign \g2098/_0_  = _w197_ ;
	assign \g21/_0_  = _w198_ ;
	assign \g2101/_0_  = _w199_ ;
endmodule;