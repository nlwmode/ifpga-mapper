module top (a_pad, b_pad, d_pad, \e0_pad , f_pad, \g0_pad , g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, \a0_pad , \b0_pad , \c0_pad , \d0_pad , \f0_pad , \h0_pad , t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad);
	input a_pad ;
	input b_pad ;
	input d_pad ;
	input \e0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	output \a0_pad  ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \d0_pad  ;
	output \f0_pad  ;
	output \h0_pad  ;
	output t_pad ;
	output u_pad ;
	output v_pad ;
	output w_pad ;
	output x_pad ;
	output y_pad ;
	output z_pad ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	LUT3 #(
		.INIT('h80)
	) name0 (
		g_pad,
		h_pad,
		i_pad,
		_w21_
	);
	LUT4 #(
		.INIT('h0080)
	) name1 (
		g_pad,
		h_pad,
		i_pad,
		j_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		k_pad,
		l_pad,
		_w23_
	);
	LUT3 #(
		.INIT('hb0)
	) name3 (
		d_pad,
		\e0_pad ,
		q_pad,
		_w24_
	);
	LUT4 #(
		.INIT('h40f0)
	) name4 (
		d_pad,
		\e0_pad ,
		\g0_pad ,
		q_pad,
		_w25_
	);
	LUT4 #(
		.INIT('h9cff)
	) name5 (
		k_pad,
		l_pad,
		_w22_,
		_w25_,
		_w26_
	);
	LUT4 #(
		.INIT('h6aff)
	) name6 (
		m_pad,
		_w22_,
		_w23_,
		_w25_,
		_w27_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name7 (
		m_pad,
		n_pad,
		_w22_,
		_w23_,
		_w28_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		k_pad,
		l_pad,
		m_pad,
		n_pad,
		_w29_
	);
	LUT3 #(
		.INIT('h4c)
	) name9 (
		_w22_,
		_w25_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('hb)
	) name10 (
		_w28_,
		_w30_,
		_w31_
	);
	LUT4 #(
		.INIT('hb000)
	) name11 (
		d_pad,
		\e0_pad ,
		o_pad,
		q_pad,
		_w32_
	);
	LUT4 #(
		.INIT('h0c08)
	) name12 (
		a_pad,
		_w22_,
		_w24_,
		_w29_,
		_w33_
	);
	LUT3 #(
		.INIT('ha8)
	) name13 (
		\g0_pad ,
		_w32_,
		_w33_,
		_w34_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name14 (
		d_pad,
		\e0_pad ,
		\g0_pad ,
		q_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\g0_pad ,
		r_pad,
		_w36_
	);
	LUT3 #(
		.INIT('h27)
	) name16 (
		b_pad,
		\e0_pad ,
		o_pad,
		_w37_
	);
	LUT4 #(
		.INIT('h7277)
	) name17 (
		f_pad,
		\g0_pad ,
		p_pad,
		s_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		g_pad,
		_w25_,
		_w39_
	);
	LUT2 #(
		.INIT('h6)
	) name19 (
		g_pad,
		h_pad,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w25_,
		_w40_,
		_w41_
	);
	LUT3 #(
		.INIT('h78)
	) name21 (
		g_pad,
		h_pad,
		i_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w25_,
		_w42_,
		_w43_
	);
	LUT3 #(
		.INIT('h6f)
	) name23 (
		j_pad,
		_w21_,
		_w25_,
		_w44_
	);
	LUT3 #(
		.INIT('h6f)
	) name24 (
		k_pad,
		_w22_,
		_w25_,
		_w45_
	);
	assign \a0_pad  = _w26_ ;
	assign \b0_pad  = _w27_ ;
	assign \c0_pad  = _w31_ ;
	assign \d0_pad  = _w34_ ;
	assign \f0_pad  = _w35_ ;
	assign \h0_pad  = _w36_ ;
	assign t_pad = _w37_ ;
	assign u_pad = _w38_ ;
	assign v_pad = _w39_ ;
	assign w_pad = _w41_ ;
	assign x_pad = _w43_ ;
	assign y_pad = _w44_ ;
	assign z_pad = _w45_ ;
endmodule;