module top( \m0_addr_i[0]_pad  , \m0_addr_i[10]_pad  , \m0_addr_i[11]_pad  , \m0_addr_i[12]_pad  , \m0_addr_i[13]_pad  , \m0_addr_i[14]_pad  , \m0_addr_i[15]_pad  , \m0_addr_i[16]_pad  , \m0_addr_i[17]_pad  , \m0_addr_i[18]_pad  , \m0_addr_i[19]_pad  , \m0_addr_i[1]_pad  , \m0_addr_i[20]_pad  , \m0_addr_i[21]_pad  , \m0_addr_i[22]_pad  , \m0_addr_i[23]_pad  , \m0_addr_i[24]_pad  , \m0_addr_i[25]_pad  , \m0_addr_i[26]_pad  , \m0_addr_i[27]_pad  , \m0_addr_i[28]_pad  , \m0_addr_i[29]_pad  , \m0_addr_i[2]_pad  , \m0_addr_i[30]_pad  , \m0_addr_i[31]_pad  , \m0_addr_i[3]_pad  , \m0_addr_i[4]_pad  , \m0_addr_i[5]_pad  , \m0_addr_i[6]_pad  , \m0_addr_i[7]_pad  , \m0_addr_i[8]_pad  , \m0_addr_i[9]_pad  , \m0_cyc_i_pad  , \m0_data_i[0]_pad  , \m0_data_i[10]_pad  , \m0_data_i[11]_pad  , \m0_data_i[12]_pad  , \m0_data_i[13]_pad  , \m0_data_i[14]_pad  , \m0_data_i[15]_pad  , \m0_data_i[16]_pad  , \m0_data_i[17]_pad  , \m0_data_i[18]_pad  , \m0_data_i[19]_pad  , \m0_data_i[1]_pad  , \m0_data_i[20]_pad  , \m0_data_i[21]_pad  , \m0_data_i[22]_pad  , \m0_data_i[23]_pad  , \m0_data_i[24]_pad  , \m0_data_i[25]_pad  , \m0_data_i[26]_pad  , \m0_data_i[27]_pad  , \m0_data_i[28]_pad  , \m0_data_i[29]_pad  , \m0_data_i[2]_pad  , \m0_data_i[30]_pad  , \m0_data_i[31]_pad  , \m0_data_i[3]_pad  , \m0_data_i[4]_pad  , \m0_data_i[5]_pad  , \m0_data_i[6]_pad  , \m0_data_i[7]_pad  , \m0_data_i[8]_pad  , \m0_data_i[9]_pad  , \m0_s0_cyc_o_reg/NET0131  , \m0_s10_cyc_o_reg/NET0131  , \m0_s11_cyc_o_reg/NET0131  , \m0_s12_cyc_o_reg/NET0131  , \m0_s13_cyc_o_reg/NET0131  , \m0_s14_cyc_o_reg/NET0131  , \m0_s15_cyc_o_reg/NET0131  , \m0_s1_cyc_o_reg/NET0131  , \m0_s2_cyc_o_reg/NET0131  , \m0_s3_cyc_o_reg/NET0131  , \m0_s4_cyc_o_reg/NET0131  , \m0_s5_cyc_o_reg/NET0131  , \m0_s6_cyc_o_reg/NET0131  , \m0_s7_cyc_o_reg/NET0131  , \m0_s8_cyc_o_reg/NET0131  , \m0_s9_cyc_o_reg/NET0131  , \m0_sel_i[0]_pad  , \m0_sel_i[1]_pad  , \m0_sel_i[2]_pad  , \m0_sel_i[3]_pad  , \m0_stb_i_pad  , \m0_we_i_pad  , \m1_addr_i[0]_pad  , \m1_addr_i[10]_pad  , \m1_addr_i[11]_pad  , \m1_addr_i[12]_pad  , \m1_addr_i[13]_pad  , \m1_addr_i[14]_pad  , \m1_addr_i[15]_pad  , \m1_addr_i[16]_pad  , \m1_addr_i[17]_pad  , \m1_addr_i[18]_pad  , \m1_addr_i[19]_pad  , \m1_addr_i[1]_pad  , \m1_addr_i[20]_pad  , \m1_addr_i[21]_pad  , \m1_addr_i[22]_pad  , \m1_addr_i[23]_pad  , \m1_addr_i[24]_pad  , \m1_addr_i[25]_pad  , \m1_addr_i[26]_pad  , \m1_addr_i[27]_pad  , \m1_addr_i[28]_pad  , \m1_addr_i[29]_pad  , \m1_addr_i[2]_pad  , \m1_addr_i[30]_pad  , \m1_addr_i[31]_pad  , \m1_addr_i[3]_pad  , \m1_addr_i[4]_pad  , \m1_addr_i[5]_pad  , \m1_addr_i[6]_pad  , \m1_addr_i[7]_pad  , \m1_addr_i[8]_pad  , \m1_addr_i[9]_pad  , \m1_cyc_i_pad  , \m1_data_i[0]_pad  , \m1_data_i[10]_pad  , \m1_data_i[11]_pad  , \m1_data_i[12]_pad  , \m1_data_i[13]_pad  , \m1_data_i[14]_pad  , \m1_data_i[15]_pad  , \m1_data_i[16]_pad  , \m1_data_i[17]_pad  , \m1_data_i[18]_pad  , \m1_data_i[19]_pad  , \m1_data_i[1]_pad  , \m1_data_i[20]_pad  , \m1_data_i[21]_pad  , \m1_data_i[22]_pad  , \m1_data_i[23]_pad  , \m1_data_i[24]_pad  , \m1_data_i[25]_pad  , \m1_data_i[26]_pad  , \m1_data_i[27]_pad  , \m1_data_i[28]_pad  , \m1_data_i[29]_pad  , \m1_data_i[2]_pad  , \m1_data_i[30]_pad  , \m1_data_i[31]_pad  , \m1_data_i[3]_pad  , \m1_data_i[4]_pad  , \m1_data_i[5]_pad  , \m1_data_i[6]_pad  , \m1_data_i[7]_pad  , \m1_data_i[8]_pad  , \m1_data_i[9]_pad  , \m1_s0_cyc_o_reg/NET0131  , \m1_s10_cyc_o_reg/NET0131  , \m1_s11_cyc_o_reg/NET0131  , \m1_s12_cyc_o_reg/NET0131  , \m1_s13_cyc_o_reg/NET0131  , \m1_s14_cyc_o_reg/NET0131  , \m1_s15_cyc_o_reg/NET0131  , \m1_s1_cyc_o_reg/NET0131  , \m1_s2_cyc_o_reg/NET0131  , \m1_s3_cyc_o_reg/NET0131  , \m1_s4_cyc_o_reg/NET0131  , \m1_s5_cyc_o_reg/NET0131  , \m1_s6_cyc_o_reg/NET0131  , \m1_s7_cyc_o_reg/NET0131  , \m1_s8_cyc_o_reg/NET0131  , \m1_s9_cyc_o_reg/NET0131  , \m1_sel_i[0]_pad  , \m1_sel_i[1]_pad  , \m1_sel_i[2]_pad  , \m1_sel_i[3]_pad  , \m1_stb_i_pad  , \m1_we_i_pad  , \m2_addr_i[0]_pad  , \m2_addr_i[10]_pad  , \m2_addr_i[11]_pad  , \m2_addr_i[12]_pad  , \m2_addr_i[13]_pad  , \m2_addr_i[14]_pad  , \m2_addr_i[15]_pad  , \m2_addr_i[16]_pad  , \m2_addr_i[17]_pad  , \m2_addr_i[18]_pad  , \m2_addr_i[19]_pad  , \m2_addr_i[1]_pad  , \m2_addr_i[20]_pad  , \m2_addr_i[21]_pad  , \m2_addr_i[22]_pad  , \m2_addr_i[23]_pad  , \m2_addr_i[24]_pad  , \m2_addr_i[25]_pad  , \m2_addr_i[26]_pad  , \m2_addr_i[27]_pad  , \m2_addr_i[28]_pad  , \m2_addr_i[29]_pad  , \m2_addr_i[2]_pad  , \m2_addr_i[30]_pad  , \m2_addr_i[31]_pad  , \m2_addr_i[3]_pad  , \m2_addr_i[4]_pad  , \m2_addr_i[5]_pad  , \m2_addr_i[6]_pad  , \m2_addr_i[7]_pad  , \m2_addr_i[8]_pad  , \m2_addr_i[9]_pad  , \m2_cyc_i_pad  , \m2_data_i[0]_pad  , \m2_data_i[10]_pad  , \m2_data_i[11]_pad  , \m2_data_i[12]_pad  , \m2_data_i[13]_pad  , \m2_data_i[14]_pad  , \m2_data_i[15]_pad  , \m2_data_i[16]_pad  , \m2_data_i[17]_pad  , \m2_data_i[18]_pad  , \m2_data_i[19]_pad  , \m2_data_i[1]_pad  , \m2_data_i[20]_pad  , \m2_data_i[21]_pad  , \m2_data_i[22]_pad  , \m2_data_i[23]_pad  , \m2_data_i[24]_pad  , \m2_data_i[25]_pad  , \m2_data_i[26]_pad  , \m2_data_i[27]_pad  , \m2_data_i[28]_pad  , \m2_data_i[29]_pad  , \m2_data_i[2]_pad  , \m2_data_i[30]_pad  , \m2_data_i[31]_pad  , \m2_data_i[3]_pad  , \m2_data_i[4]_pad  , \m2_data_i[5]_pad  , \m2_data_i[6]_pad  , \m2_data_i[7]_pad  , \m2_data_i[8]_pad  , \m2_data_i[9]_pad  , \m2_s0_cyc_o_reg/NET0131  , \m2_s10_cyc_o_reg/NET0131  , \m2_s11_cyc_o_reg/NET0131  , \m2_s12_cyc_o_reg/NET0131  , \m2_s13_cyc_o_reg/NET0131  , \m2_s14_cyc_o_reg/NET0131  , \m2_s15_cyc_o_reg/NET0131  , \m2_s1_cyc_o_reg/NET0131  , \m2_s2_cyc_o_reg/NET0131  , \m2_s3_cyc_o_reg/NET0131  , \m2_s4_cyc_o_reg/NET0131  , \m2_s5_cyc_o_reg/NET0131  , \m2_s6_cyc_o_reg/NET0131  , \m2_s7_cyc_o_reg/NET0131  , \m2_s8_cyc_o_reg/NET0131  , \m2_s9_cyc_o_reg/NET0131  , \m2_sel_i[0]_pad  , \m2_sel_i[1]_pad  , \m2_sel_i[2]_pad  , \m2_sel_i[3]_pad  , \m2_stb_i_pad  , \m2_we_i_pad  , \m3_addr_i[0]_pad  , \m3_addr_i[10]_pad  , \m3_addr_i[11]_pad  , \m3_addr_i[12]_pad  , \m3_addr_i[13]_pad  , \m3_addr_i[14]_pad  , \m3_addr_i[15]_pad  , \m3_addr_i[16]_pad  , \m3_addr_i[17]_pad  , \m3_addr_i[18]_pad  , \m3_addr_i[19]_pad  , \m3_addr_i[1]_pad  , \m3_addr_i[20]_pad  , \m3_addr_i[21]_pad  , \m3_addr_i[22]_pad  , \m3_addr_i[23]_pad  , \m3_addr_i[24]_pad  , \m3_addr_i[25]_pad  , \m3_addr_i[26]_pad  , \m3_addr_i[27]_pad  , \m3_addr_i[28]_pad  , \m3_addr_i[29]_pad  , \m3_addr_i[2]_pad  , \m3_addr_i[30]_pad  , \m3_addr_i[31]_pad  , \m3_addr_i[3]_pad  , \m3_addr_i[4]_pad  , \m3_addr_i[5]_pad  , \m3_addr_i[6]_pad  , \m3_addr_i[7]_pad  , \m3_addr_i[8]_pad  , \m3_addr_i[9]_pad  , \m3_cyc_i_pad  , \m3_data_i[0]_pad  , \m3_data_i[10]_pad  , \m3_data_i[11]_pad  , \m3_data_i[12]_pad  , \m3_data_i[13]_pad  , \m3_data_i[14]_pad  , \m3_data_i[15]_pad  , \m3_data_i[16]_pad  , \m3_data_i[17]_pad  , \m3_data_i[18]_pad  , \m3_data_i[19]_pad  , \m3_data_i[1]_pad  , \m3_data_i[20]_pad  , \m3_data_i[21]_pad  , \m3_data_i[22]_pad  , \m3_data_i[23]_pad  , \m3_data_i[24]_pad  , \m3_data_i[25]_pad  , \m3_data_i[26]_pad  , \m3_data_i[27]_pad  , \m3_data_i[28]_pad  , \m3_data_i[29]_pad  , \m3_data_i[2]_pad  , \m3_data_i[30]_pad  , \m3_data_i[31]_pad  , \m3_data_i[3]_pad  , \m3_data_i[4]_pad  , \m3_data_i[5]_pad  , \m3_data_i[6]_pad  , \m3_data_i[7]_pad  , \m3_data_i[8]_pad  , \m3_data_i[9]_pad  , \m3_s0_cyc_o_reg/NET0131  , \m3_s10_cyc_o_reg/NET0131  , \m3_s11_cyc_o_reg/NET0131  , \m3_s12_cyc_o_reg/NET0131  , \m3_s13_cyc_o_reg/NET0131  , \m3_s14_cyc_o_reg/NET0131  , \m3_s15_cyc_o_reg/NET0131  , \m3_s1_cyc_o_reg/NET0131  , \m3_s2_cyc_o_reg/NET0131  , \m3_s3_cyc_o_reg/NET0131  , \m3_s4_cyc_o_reg/NET0131  , \m3_s5_cyc_o_reg/NET0131  , \m3_s6_cyc_o_reg/NET0131  , \m3_s7_cyc_o_reg/NET0131  , \m3_s8_cyc_o_reg/NET0131  , \m3_s9_cyc_o_reg/NET0131  , \m3_sel_i[0]_pad  , \m3_sel_i[1]_pad  , \m3_sel_i[2]_pad  , \m3_sel_i[3]_pad  , \m3_stb_i_pad  , \m3_we_i_pad  , \m4_addr_i[0]_pad  , \m4_addr_i[10]_pad  , \m4_addr_i[11]_pad  , \m4_addr_i[12]_pad  , \m4_addr_i[13]_pad  , \m4_addr_i[14]_pad  , \m4_addr_i[15]_pad  , \m4_addr_i[16]_pad  , \m4_addr_i[17]_pad  , \m4_addr_i[18]_pad  , \m4_addr_i[19]_pad  , \m4_addr_i[1]_pad  , \m4_addr_i[20]_pad  , \m4_addr_i[21]_pad  , \m4_addr_i[22]_pad  , \m4_addr_i[23]_pad  , \m4_addr_i[24]_pad  , \m4_addr_i[25]_pad  , \m4_addr_i[26]_pad  , \m4_addr_i[27]_pad  , \m4_addr_i[28]_pad  , \m4_addr_i[29]_pad  , \m4_addr_i[2]_pad  , \m4_addr_i[30]_pad  , \m4_addr_i[31]_pad  , \m4_addr_i[3]_pad  , \m4_addr_i[4]_pad  , \m4_addr_i[5]_pad  , \m4_addr_i[6]_pad  , \m4_addr_i[7]_pad  , \m4_addr_i[8]_pad  , \m4_addr_i[9]_pad  , \m4_cyc_i_pad  , \m4_data_i[0]_pad  , \m4_data_i[10]_pad  , \m4_data_i[11]_pad  , \m4_data_i[12]_pad  , \m4_data_i[13]_pad  , \m4_data_i[14]_pad  , \m4_data_i[15]_pad  , \m4_data_i[16]_pad  , \m4_data_i[17]_pad  , \m4_data_i[18]_pad  , \m4_data_i[19]_pad  , \m4_data_i[1]_pad  , \m4_data_i[20]_pad  , \m4_data_i[21]_pad  , \m4_data_i[22]_pad  , \m4_data_i[23]_pad  , \m4_data_i[24]_pad  , \m4_data_i[25]_pad  , \m4_data_i[26]_pad  , \m4_data_i[27]_pad  , \m4_data_i[28]_pad  , \m4_data_i[29]_pad  , \m4_data_i[2]_pad  , \m4_data_i[30]_pad  , \m4_data_i[31]_pad  , \m4_data_i[3]_pad  , \m4_data_i[4]_pad  , \m4_data_i[5]_pad  , \m4_data_i[6]_pad  , \m4_data_i[7]_pad  , \m4_data_i[8]_pad  , \m4_data_i[9]_pad  , \m4_s0_cyc_o_reg/NET0131  , \m4_s10_cyc_o_reg/NET0131  , \m4_s11_cyc_o_reg/NET0131  , \m4_s12_cyc_o_reg/NET0131  , \m4_s13_cyc_o_reg/NET0131  , \m4_s14_cyc_o_reg/NET0131  , \m4_s15_cyc_o_reg/NET0131  , \m4_s1_cyc_o_reg/NET0131  , \m4_s2_cyc_o_reg/NET0131  , \m4_s3_cyc_o_reg/NET0131  , \m4_s4_cyc_o_reg/NET0131  , \m4_s5_cyc_o_reg/NET0131  , \m4_s6_cyc_o_reg/NET0131  , \m4_s7_cyc_o_reg/NET0131  , \m4_s8_cyc_o_reg/NET0131  , \m4_s9_cyc_o_reg/NET0131  , \m4_sel_i[0]_pad  , \m4_sel_i[1]_pad  , \m4_sel_i[2]_pad  , \m4_sel_i[3]_pad  , \m4_stb_i_pad  , \m4_we_i_pad  , \m5_addr_i[0]_pad  , \m5_addr_i[10]_pad  , \m5_addr_i[11]_pad  , \m5_addr_i[12]_pad  , \m5_addr_i[13]_pad  , \m5_addr_i[14]_pad  , \m5_addr_i[15]_pad  , \m5_addr_i[16]_pad  , \m5_addr_i[17]_pad  , \m5_addr_i[18]_pad  , \m5_addr_i[19]_pad  , \m5_addr_i[1]_pad  , \m5_addr_i[20]_pad  , \m5_addr_i[21]_pad  , \m5_addr_i[22]_pad  , \m5_addr_i[23]_pad  , \m5_addr_i[24]_pad  , \m5_addr_i[25]_pad  , \m5_addr_i[26]_pad  , \m5_addr_i[27]_pad  , \m5_addr_i[28]_pad  , \m5_addr_i[29]_pad  , \m5_addr_i[2]_pad  , \m5_addr_i[30]_pad  , \m5_addr_i[31]_pad  , \m5_addr_i[3]_pad  , \m5_addr_i[4]_pad  , \m5_addr_i[5]_pad  , \m5_addr_i[6]_pad  , \m5_addr_i[7]_pad  , \m5_addr_i[8]_pad  , \m5_addr_i[9]_pad  , \m5_cyc_i_pad  , \m5_data_i[0]_pad  , \m5_data_i[10]_pad  , \m5_data_i[11]_pad  , \m5_data_i[12]_pad  , \m5_data_i[13]_pad  , \m5_data_i[14]_pad  , \m5_data_i[15]_pad  , \m5_data_i[16]_pad  , \m5_data_i[17]_pad  , \m5_data_i[18]_pad  , \m5_data_i[19]_pad  , \m5_data_i[1]_pad  , \m5_data_i[20]_pad  , \m5_data_i[21]_pad  , \m5_data_i[22]_pad  , \m5_data_i[23]_pad  , \m5_data_i[24]_pad  , \m5_data_i[25]_pad  , \m5_data_i[26]_pad  , \m5_data_i[27]_pad  , \m5_data_i[28]_pad  , \m5_data_i[29]_pad  , \m5_data_i[2]_pad  , \m5_data_i[30]_pad  , \m5_data_i[31]_pad  , \m5_data_i[3]_pad  , \m5_data_i[4]_pad  , \m5_data_i[5]_pad  , \m5_data_i[6]_pad  , \m5_data_i[7]_pad  , \m5_data_i[8]_pad  , \m5_data_i[9]_pad  , \m5_s0_cyc_o_reg/NET0131  , \m5_s10_cyc_o_reg/NET0131  , \m5_s11_cyc_o_reg/NET0131  , \m5_s12_cyc_o_reg/NET0131  , \m5_s13_cyc_o_reg/NET0131  , \m5_s14_cyc_o_reg/NET0131  , \m5_s15_cyc_o_reg/NET0131  , \m5_s1_cyc_o_reg/NET0131  , \m5_s2_cyc_o_reg/NET0131  , \m5_s3_cyc_o_reg/NET0131  , \m5_s4_cyc_o_reg/NET0131  , \m5_s5_cyc_o_reg/NET0131  , \m5_s6_cyc_o_reg/NET0131  , \m5_s7_cyc_o_reg/NET0131  , \m5_s8_cyc_o_reg/NET0131  , \m5_s9_cyc_o_reg/NET0131  , \m5_sel_i[0]_pad  , \m5_sel_i[1]_pad  , \m5_sel_i[2]_pad  , \m5_sel_i[3]_pad  , \m5_stb_i_pad  , \m5_we_i_pad  , \m6_addr_i[0]_pad  , \m6_addr_i[10]_pad  , \m6_addr_i[11]_pad  , \m6_addr_i[12]_pad  , \m6_addr_i[13]_pad  , \m6_addr_i[14]_pad  , \m6_addr_i[15]_pad  , \m6_addr_i[16]_pad  , \m6_addr_i[17]_pad  , \m6_addr_i[18]_pad  , \m6_addr_i[19]_pad  , \m6_addr_i[1]_pad  , \m6_addr_i[20]_pad  , \m6_addr_i[21]_pad  , \m6_addr_i[22]_pad  , \m6_addr_i[23]_pad  , \m6_addr_i[24]_pad  , \m6_addr_i[25]_pad  , \m6_addr_i[26]_pad  , \m6_addr_i[27]_pad  , \m6_addr_i[28]_pad  , \m6_addr_i[29]_pad  , \m6_addr_i[2]_pad  , \m6_addr_i[30]_pad  , \m6_addr_i[31]_pad  , \m6_addr_i[3]_pad  , \m6_addr_i[4]_pad  , \m6_addr_i[5]_pad  , \m6_addr_i[6]_pad  , \m6_addr_i[7]_pad  , \m6_addr_i[8]_pad  , \m6_addr_i[9]_pad  , \m6_cyc_i_pad  , \m6_data_i[0]_pad  , \m6_data_i[10]_pad  , \m6_data_i[11]_pad  , \m6_data_i[12]_pad  , \m6_data_i[13]_pad  , \m6_data_i[14]_pad  , \m6_data_i[15]_pad  , \m6_data_i[16]_pad  , \m6_data_i[17]_pad  , \m6_data_i[18]_pad  , \m6_data_i[19]_pad  , \m6_data_i[1]_pad  , \m6_data_i[20]_pad  , \m6_data_i[21]_pad  , \m6_data_i[22]_pad  , \m6_data_i[23]_pad  , \m6_data_i[24]_pad  , \m6_data_i[25]_pad  , \m6_data_i[26]_pad  , \m6_data_i[27]_pad  , \m6_data_i[28]_pad  , \m6_data_i[29]_pad  , \m6_data_i[2]_pad  , \m6_data_i[30]_pad  , \m6_data_i[31]_pad  , \m6_data_i[3]_pad  , \m6_data_i[4]_pad  , \m6_data_i[5]_pad  , \m6_data_i[6]_pad  , \m6_data_i[7]_pad  , \m6_data_i[8]_pad  , \m6_data_i[9]_pad  , \m6_s0_cyc_o_reg/NET0131  , \m6_s10_cyc_o_reg/NET0131  , \m6_s11_cyc_o_reg/NET0131  , \m6_s12_cyc_o_reg/NET0131  , \m6_s13_cyc_o_reg/NET0131  , \m6_s14_cyc_o_reg/NET0131  , \m6_s15_cyc_o_reg/NET0131  , \m6_s1_cyc_o_reg/NET0131  , \m6_s2_cyc_o_reg/NET0131  , \m6_s3_cyc_o_reg/NET0131  , \m6_s4_cyc_o_reg/NET0131  , \m6_s5_cyc_o_reg/NET0131  , \m6_s6_cyc_o_reg/NET0131  , \m6_s7_cyc_o_reg/NET0131  , \m6_s8_cyc_o_reg/NET0131  , \m6_s9_cyc_o_reg/NET0131  , \m6_sel_i[0]_pad  , \m6_sel_i[1]_pad  , \m6_sel_i[2]_pad  , \m6_sel_i[3]_pad  , \m6_stb_i_pad  , \m6_we_i_pad  , \m7_addr_i[0]_pad  , \m7_addr_i[10]_pad  , \m7_addr_i[11]_pad  , \m7_addr_i[12]_pad  , \m7_addr_i[13]_pad  , \m7_addr_i[14]_pad  , \m7_addr_i[15]_pad  , \m7_addr_i[16]_pad  , \m7_addr_i[17]_pad  , \m7_addr_i[18]_pad  , \m7_addr_i[19]_pad  , \m7_addr_i[1]_pad  , \m7_addr_i[20]_pad  , \m7_addr_i[21]_pad  , \m7_addr_i[22]_pad  , \m7_addr_i[23]_pad  , \m7_addr_i[24]_pad  , \m7_addr_i[25]_pad  , \m7_addr_i[26]_pad  , \m7_addr_i[27]_pad  , \m7_addr_i[28]_pad  , \m7_addr_i[29]_pad  , \m7_addr_i[2]_pad  , \m7_addr_i[30]_pad  , \m7_addr_i[31]_pad  , \m7_addr_i[3]_pad  , \m7_addr_i[4]_pad  , \m7_addr_i[5]_pad  , \m7_addr_i[6]_pad  , \m7_addr_i[7]_pad  , \m7_addr_i[8]_pad  , \m7_addr_i[9]_pad  , \m7_cyc_i_pad  , \m7_data_i[0]_pad  , \m7_data_i[10]_pad  , \m7_data_i[11]_pad  , \m7_data_i[12]_pad  , \m7_data_i[13]_pad  , \m7_data_i[14]_pad  , \m7_data_i[15]_pad  , \m7_data_i[16]_pad  , \m7_data_i[17]_pad  , \m7_data_i[18]_pad  , \m7_data_i[19]_pad  , \m7_data_i[1]_pad  , \m7_data_i[20]_pad  , \m7_data_i[21]_pad  , \m7_data_i[22]_pad  , \m7_data_i[23]_pad  , \m7_data_i[24]_pad  , \m7_data_i[25]_pad  , \m7_data_i[26]_pad  , \m7_data_i[27]_pad  , \m7_data_i[28]_pad  , \m7_data_i[29]_pad  , \m7_data_i[2]_pad  , \m7_data_i[30]_pad  , \m7_data_i[31]_pad  , \m7_data_i[3]_pad  , \m7_data_i[4]_pad  , \m7_data_i[5]_pad  , \m7_data_i[6]_pad  , \m7_data_i[7]_pad  , \m7_data_i[8]_pad  , \m7_data_i[9]_pad  , \m7_s0_cyc_o_reg/NET0131  , \m7_s10_cyc_o_reg/NET0131  , \m7_s11_cyc_o_reg/NET0131  , \m7_s12_cyc_o_reg/NET0131  , \m7_s13_cyc_o_reg/NET0131  , \m7_s14_cyc_o_reg/NET0131  , \m7_s15_cyc_o_reg/NET0131  , \m7_s1_cyc_o_reg/NET0131  , \m7_s2_cyc_o_reg/NET0131  , \m7_s3_cyc_o_reg/NET0131  , \m7_s4_cyc_o_reg/NET0131  , \m7_s5_cyc_o_reg/NET0131  , \m7_s6_cyc_o_reg/NET0131  , \m7_s7_cyc_o_reg/NET0131  , \m7_s8_cyc_o_reg/NET0131  , \m7_s9_cyc_o_reg/NET0131  , \m7_sel_i[0]_pad  , \m7_sel_i[1]_pad  , \m7_sel_i[2]_pad  , \m7_sel_i[3]_pad  , \m7_stb_i_pad  , \m7_we_i_pad  , \rf_conf0_reg[0]/NET0131  , \rf_conf0_reg[10]/NET0131  , \rf_conf0_reg[11]/NET0131  , \rf_conf0_reg[12]/NET0131  , \rf_conf0_reg[13]/NET0131  , \rf_conf0_reg[14]/NET0131  , \rf_conf0_reg[15]/NET0131  , \rf_conf0_reg[1]/NET0131  , \rf_conf0_reg[2]/NET0131  , \rf_conf0_reg[3]/NET0131  , \rf_conf0_reg[4]/NET0131  , \rf_conf0_reg[5]/NET0131  , \rf_conf0_reg[6]/NET0131  , \rf_conf0_reg[7]/NET0131  , \rf_conf0_reg[8]/NET0131  , \rf_conf0_reg[9]/NET0131  , \rf_conf10_reg[0]/NET0131  , \rf_conf10_reg[10]/NET0131  , \rf_conf10_reg[11]/NET0131  , \rf_conf10_reg[12]/NET0131  , \rf_conf10_reg[13]/NET0131  , \rf_conf10_reg[14]/NET0131  , \rf_conf10_reg[15]/NET0131  , \rf_conf10_reg[1]/NET0131  , \rf_conf10_reg[2]/NET0131  , \rf_conf10_reg[3]/NET0131  , \rf_conf10_reg[4]/NET0131  , \rf_conf10_reg[5]/NET0131  , \rf_conf10_reg[6]/NET0131  , \rf_conf10_reg[7]/NET0131  , \rf_conf10_reg[8]/NET0131  , \rf_conf10_reg[9]/NET0131  , \rf_conf11_reg[0]/NET0131  , \rf_conf11_reg[10]/NET0131  , \rf_conf11_reg[11]/NET0131  , \rf_conf11_reg[12]/NET0131  , \rf_conf11_reg[13]/NET0131  , \rf_conf11_reg[14]/NET0131  , \rf_conf11_reg[15]/NET0131  , \rf_conf11_reg[1]/NET0131  , \rf_conf11_reg[2]/NET0131  , \rf_conf11_reg[3]/NET0131  , \rf_conf11_reg[4]/NET0131  , \rf_conf11_reg[5]/NET0131  , \rf_conf11_reg[6]/NET0131  , \rf_conf11_reg[7]/NET0131  , \rf_conf11_reg[8]/NET0131  , \rf_conf11_reg[9]/NET0131  , \rf_conf12_reg[0]/NET0131  , \rf_conf12_reg[10]/NET0131  , \rf_conf12_reg[11]/NET0131  , \rf_conf12_reg[12]/NET0131  , \rf_conf12_reg[13]/NET0131  , \rf_conf12_reg[14]/NET0131  , \rf_conf12_reg[15]/NET0131  , \rf_conf12_reg[1]/NET0131  , \rf_conf12_reg[2]/NET0131  , \rf_conf12_reg[3]/NET0131  , \rf_conf12_reg[4]/NET0131  , \rf_conf12_reg[5]/NET0131  , \rf_conf12_reg[6]/NET0131  , \rf_conf12_reg[7]/NET0131  , \rf_conf12_reg[8]/NET0131  , \rf_conf12_reg[9]/NET0131  , \rf_conf13_reg[0]/NET0131  , \rf_conf13_reg[10]/NET0131  , \rf_conf13_reg[11]/NET0131  , \rf_conf13_reg[12]/NET0131  , \rf_conf13_reg[13]/NET0131  , \rf_conf13_reg[14]/NET0131  , \rf_conf13_reg[15]/NET0131  , \rf_conf13_reg[1]/NET0131  , \rf_conf13_reg[2]/NET0131  , \rf_conf13_reg[3]/NET0131  , \rf_conf13_reg[4]/NET0131  , \rf_conf13_reg[5]/NET0131  , \rf_conf13_reg[6]/NET0131  , \rf_conf13_reg[7]/NET0131  , \rf_conf13_reg[8]/NET0131  , \rf_conf13_reg[9]/NET0131  , \rf_conf14_reg[0]/NET0131  , \rf_conf14_reg[10]/NET0131  , \rf_conf14_reg[11]/NET0131  , \rf_conf14_reg[12]/NET0131  , \rf_conf14_reg[13]/NET0131  , \rf_conf14_reg[14]/NET0131  , \rf_conf14_reg[15]/NET0131  , \rf_conf14_reg[1]/NET0131  , \rf_conf14_reg[2]/NET0131  , \rf_conf14_reg[3]/NET0131  , \rf_conf14_reg[4]/NET0131  , \rf_conf14_reg[5]/NET0131  , \rf_conf14_reg[6]/NET0131  , \rf_conf14_reg[7]/NET0131  , \rf_conf14_reg[8]/NET0131  , \rf_conf14_reg[9]/NET0131  , \rf_conf15_reg[0]/NET0131  , \rf_conf15_reg[10]/NET0131  , \rf_conf15_reg[11]/NET0131  , \rf_conf15_reg[12]/NET0131  , \rf_conf15_reg[13]/NET0131  , \rf_conf15_reg[14]/NET0131  , \rf_conf15_reg[15]/NET0131  , \rf_conf15_reg[1]/NET0131  , \rf_conf15_reg[2]/NET0131  , \rf_conf15_reg[3]/NET0131  , \rf_conf15_reg[4]/NET0131  , \rf_conf15_reg[5]/NET0131  , \rf_conf15_reg[6]/NET0131  , \rf_conf15_reg[7]/NET0131  , \rf_conf15_reg[8]/NET0131  , \rf_conf15_reg[9]/NET0131  , \rf_conf1_reg[0]/NET0131  , \rf_conf1_reg[10]/NET0131  , \rf_conf1_reg[11]/NET0131  , \rf_conf1_reg[12]/NET0131  , \rf_conf1_reg[13]/NET0131  , \rf_conf1_reg[14]/NET0131  , \rf_conf1_reg[15]/NET0131  , \rf_conf1_reg[1]/NET0131  , \rf_conf1_reg[2]/NET0131  , \rf_conf1_reg[3]/NET0131  , \rf_conf1_reg[4]/NET0131  , \rf_conf1_reg[5]/NET0131  , \rf_conf1_reg[6]/NET0131  , \rf_conf1_reg[7]/NET0131  , \rf_conf1_reg[8]/NET0131  , \rf_conf1_reg[9]/NET0131  , \rf_conf2_reg[0]/NET0131  , \rf_conf2_reg[10]/NET0131  , \rf_conf2_reg[11]/NET0131  , \rf_conf2_reg[12]/NET0131  , \rf_conf2_reg[13]/NET0131  , \rf_conf2_reg[14]/NET0131  , \rf_conf2_reg[15]/NET0131  , \rf_conf2_reg[1]/NET0131  , \rf_conf2_reg[2]/NET0131  , \rf_conf2_reg[3]/NET0131  , \rf_conf2_reg[4]/NET0131  , \rf_conf2_reg[5]/NET0131  , \rf_conf2_reg[6]/NET0131  , \rf_conf2_reg[7]/NET0131  , \rf_conf2_reg[8]/NET0131  , \rf_conf2_reg[9]/NET0131  , \rf_conf3_reg[0]/NET0131  , \rf_conf3_reg[10]/NET0131  , \rf_conf3_reg[11]/NET0131  , \rf_conf3_reg[12]/NET0131  , \rf_conf3_reg[13]/NET0131  , \rf_conf3_reg[14]/NET0131  , \rf_conf3_reg[15]/NET0131  , \rf_conf3_reg[1]/NET0131  , \rf_conf3_reg[2]/NET0131  , \rf_conf3_reg[3]/NET0131  , \rf_conf3_reg[4]/NET0131  , \rf_conf3_reg[5]/NET0131  , \rf_conf3_reg[6]/NET0131  , \rf_conf3_reg[7]/NET0131  , \rf_conf3_reg[8]/NET0131  , \rf_conf3_reg[9]/NET0131  , \rf_conf4_reg[0]/NET0131  , \rf_conf4_reg[10]/NET0131  , \rf_conf4_reg[11]/NET0131  , \rf_conf4_reg[12]/NET0131  , \rf_conf4_reg[13]/NET0131  , \rf_conf4_reg[14]/NET0131  , \rf_conf4_reg[15]/NET0131  , \rf_conf4_reg[1]/NET0131  , \rf_conf4_reg[2]/NET0131  , \rf_conf4_reg[3]/NET0131  , \rf_conf4_reg[4]/NET0131  , \rf_conf4_reg[5]/NET0131  , \rf_conf4_reg[6]/NET0131  , \rf_conf4_reg[7]/NET0131  , \rf_conf4_reg[8]/NET0131  , \rf_conf4_reg[9]/NET0131  , \rf_conf5_reg[0]/NET0131  , \rf_conf5_reg[10]/NET0131  , \rf_conf5_reg[11]/NET0131  , \rf_conf5_reg[12]/NET0131  , \rf_conf5_reg[13]/NET0131  , \rf_conf5_reg[14]/NET0131  , \rf_conf5_reg[15]/NET0131  , \rf_conf5_reg[1]/NET0131  , \rf_conf5_reg[2]/NET0131  , \rf_conf5_reg[3]/NET0131  , \rf_conf5_reg[4]/NET0131  , \rf_conf5_reg[5]/NET0131  , \rf_conf5_reg[6]/NET0131  , \rf_conf5_reg[7]/NET0131  , \rf_conf5_reg[8]/NET0131  , \rf_conf5_reg[9]/NET0131  , \rf_conf6_reg[0]/NET0131  , \rf_conf6_reg[10]/NET0131  , \rf_conf6_reg[11]/NET0131  , \rf_conf6_reg[12]/NET0131  , \rf_conf6_reg[13]/NET0131  , \rf_conf6_reg[14]/NET0131  , \rf_conf6_reg[15]/NET0131  , \rf_conf6_reg[1]/NET0131  , \rf_conf6_reg[2]/NET0131  , \rf_conf6_reg[3]/NET0131  , \rf_conf6_reg[4]/NET0131  , \rf_conf6_reg[5]/NET0131  , \rf_conf6_reg[6]/NET0131  , \rf_conf6_reg[7]/NET0131  , \rf_conf6_reg[8]/NET0131  , \rf_conf6_reg[9]/NET0131  , \rf_conf7_reg[0]/NET0131  , \rf_conf7_reg[10]/NET0131  , \rf_conf7_reg[11]/NET0131  , \rf_conf7_reg[12]/NET0131  , \rf_conf7_reg[13]/NET0131  , \rf_conf7_reg[14]/NET0131  , \rf_conf7_reg[15]/NET0131  , \rf_conf7_reg[1]/NET0131  , \rf_conf7_reg[2]/NET0131  , \rf_conf7_reg[3]/NET0131  , \rf_conf7_reg[4]/NET0131  , \rf_conf7_reg[5]/NET0131  , \rf_conf7_reg[6]/NET0131  , \rf_conf7_reg[7]/NET0131  , \rf_conf7_reg[8]/NET0131  , \rf_conf7_reg[9]/NET0131  , \rf_conf8_reg[0]/NET0131  , \rf_conf8_reg[10]/NET0131  , \rf_conf8_reg[11]/NET0131  , \rf_conf8_reg[12]/NET0131  , \rf_conf8_reg[13]/NET0131  , \rf_conf8_reg[14]/NET0131  , \rf_conf8_reg[15]/NET0131  , \rf_conf8_reg[1]/NET0131  , \rf_conf8_reg[2]/NET0131  , \rf_conf8_reg[3]/NET0131  , \rf_conf8_reg[4]/NET0131  , \rf_conf8_reg[5]/NET0131  , \rf_conf8_reg[6]/NET0131  , \rf_conf8_reg[7]/NET0131  , \rf_conf8_reg[8]/NET0131  , \rf_conf8_reg[9]/NET0131  , \rf_conf9_reg[0]/NET0131  , \rf_conf9_reg[10]/NET0131  , \rf_conf9_reg[11]/NET0131  , \rf_conf9_reg[12]/NET0131  , \rf_conf9_reg[13]/NET0131  , \rf_conf9_reg[14]/NET0131  , \rf_conf9_reg[15]/NET0131  , \rf_conf9_reg[1]/NET0131  , \rf_conf9_reg[2]/NET0131  , \rf_conf9_reg[3]/NET0131  , \rf_conf9_reg[4]/NET0131  , \rf_conf9_reg[5]/NET0131  , \rf_conf9_reg[6]/NET0131  , \rf_conf9_reg[7]/NET0131  , \rf_conf9_reg[8]/NET0131  , \rf_conf9_reg[9]/NET0131  , \rf_rf_ack_reg/P0001  , \rf_rf_dout_reg[0]/P0001  , \rf_rf_dout_reg[10]/P0001  , \rf_rf_dout_reg[11]/P0001  , \rf_rf_dout_reg[12]/P0001  , \rf_rf_dout_reg[13]/P0001  , \rf_rf_dout_reg[14]/P0001  , \rf_rf_dout_reg[15]/P0001  , \rf_rf_dout_reg[1]/P0001  , \rf_rf_dout_reg[2]/P0001  , \rf_rf_dout_reg[3]/P0001  , \rf_rf_dout_reg[4]/P0001  , \rf_rf_dout_reg[5]/P0001  , \rf_rf_dout_reg[6]/P0001  , \rf_rf_dout_reg[7]/P0001  , \rf_rf_dout_reg[8]/P0001  , \rf_rf_dout_reg[9]/P0001  , \rf_rf_we_reg/P0001  , rst_i_pad , \s0_ack_i_pad  , \s0_data_i[0]_pad  , \s0_data_i[10]_pad  , \s0_data_i[11]_pad  , \s0_data_i[12]_pad  , \s0_data_i[13]_pad  , \s0_data_i[14]_pad  , \s0_data_i[15]_pad  , \s0_data_i[16]_pad  , \s0_data_i[17]_pad  , \s0_data_i[18]_pad  , \s0_data_i[19]_pad  , \s0_data_i[1]_pad  , \s0_data_i[20]_pad  , \s0_data_i[21]_pad  , \s0_data_i[22]_pad  , \s0_data_i[23]_pad  , \s0_data_i[24]_pad  , \s0_data_i[25]_pad  , \s0_data_i[26]_pad  , \s0_data_i[27]_pad  , \s0_data_i[28]_pad  , \s0_data_i[29]_pad  , \s0_data_i[2]_pad  , \s0_data_i[30]_pad  , \s0_data_i[31]_pad  , \s0_data_i[3]_pad  , \s0_data_i[4]_pad  , \s0_data_i[5]_pad  , \s0_data_i[6]_pad  , \s0_data_i[7]_pad  , \s0_data_i[8]_pad  , \s0_data_i[9]_pad  , \s0_err_i_pad  , \s0_m0_cyc_r_reg/P0001  , \s0_m1_cyc_r_reg/P0001  , \s0_m2_cyc_r_reg/P0001  , \s0_m3_cyc_r_reg/P0001  , \s0_m4_cyc_r_reg/P0001  , \s0_m5_cyc_r_reg/P0001  , \s0_m6_cyc_r_reg/P0001  , \s0_m7_cyc_r_reg/P0001  , \s0_msel_arb0_state_reg[0]/NET0131  , \s0_msel_arb0_state_reg[1]/NET0131  , \s0_msel_arb0_state_reg[2]/NET0131  , \s0_msel_arb1_state_reg[0]/NET0131  , \s0_msel_arb1_state_reg[1]/NET0131  , \s0_msel_arb1_state_reg[2]/NET0131  , \s0_msel_arb2_state_reg[0]/NET0131  , \s0_msel_arb2_state_reg[1]/NET0131  , \s0_msel_arb2_state_reg[2]/NET0131  , \s0_msel_arb3_state_reg[0]/NET0131  , \s0_msel_arb3_state_reg[1]/NET0131  , \s0_msel_arb3_state_reg[2]/NET0131  , \s0_msel_pri_out_reg[0]/NET0131  , \s0_msel_pri_out_reg[1]/NET0131  , \s0_next_reg/P0001  , \s0_rty_i_pad  , \s10_ack_i_pad  , \s10_data_i[0]_pad  , \s10_data_i[10]_pad  , \s10_data_i[11]_pad  , \s10_data_i[12]_pad  , \s10_data_i[13]_pad  , \s10_data_i[14]_pad  , \s10_data_i[15]_pad  , \s10_data_i[16]_pad  , \s10_data_i[17]_pad  , \s10_data_i[18]_pad  , \s10_data_i[19]_pad  , \s10_data_i[1]_pad  , \s10_data_i[20]_pad  , \s10_data_i[21]_pad  , \s10_data_i[22]_pad  , \s10_data_i[23]_pad  , \s10_data_i[24]_pad  , \s10_data_i[25]_pad  , \s10_data_i[26]_pad  , \s10_data_i[27]_pad  , \s10_data_i[28]_pad  , \s10_data_i[29]_pad  , \s10_data_i[2]_pad  , \s10_data_i[30]_pad  , \s10_data_i[31]_pad  , \s10_data_i[3]_pad  , \s10_data_i[4]_pad  , \s10_data_i[5]_pad  , \s10_data_i[6]_pad  , \s10_data_i[7]_pad  , \s10_data_i[8]_pad  , \s10_data_i[9]_pad  , \s10_err_i_pad  , \s10_m0_cyc_r_reg/P0001  , \s10_m1_cyc_r_reg/P0001  , \s10_m2_cyc_r_reg/P0001  , \s10_m3_cyc_r_reg/P0001  , \s10_m4_cyc_r_reg/P0001  , \s10_m5_cyc_r_reg/P0001  , \s10_m6_cyc_r_reg/P0001  , \s10_m7_cyc_r_reg/P0001  , \s10_msel_arb0_state_reg[0]/NET0131  , \s10_msel_arb0_state_reg[1]/NET0131  , \s10_msel_arb0_state_reg[2]/NET0131  , \s10_msel_arb1_state_reg[0]/NET0131  , \s10_msel_arb1_state_reg[1]/NET0131  , \s10_msel_arb1_state_reg[2]/NET0131  , \s10_msel_arb2_state_reg[0]/NET0131  , \s10_msel_arb2_state_reg[1]/NET0131  , \s10_msel_arb2_state_reg[2]/NET0131  , \s10_msel_arb3_state_reg[0]/NET0131  , \s10_msel_arb3_state_reg[1]/NET0131  , \s10_msel_arb3_state_reg[2]/NET0131  , \s10_msel_pri_out_reg[0]/NET0131  , \s10_msel_pri_out_reg[1]/NET0131  , \s10_next_reg/P0001  , \s10_rty_i_pad  , \s11_ack_i_pad  , \s11_data_i[0]_pad  , \s11_data_i[10]_pad  , \s11_data_i[11]_pad  , \s11_data_i[12]_pad  , \s11_data_i[13]_pad  , \s11_data_i[14]_pad  , \s11_data_i[15]_pad  , \s11_data_i[16]_pad  , \s11_data_i[17]_pad  , \s11_data_i[18]_pad  , \s11_data_i[19]_pad  , \s11_data_i[1]_pad  , \s11_data_i[20]_pad  , \s11_data_i[21]_pad  , \s11_data_i[22]_pad  , \s11_data_i[23]_pad  , \s11_data_i[24]_pad  , \s11_data_i[25]_pad  , \s11_data_i[26]_pad  , \s11_data_i[27]_pad  , \s11_data_i[28]_pad  , \s11_data_i[29]_pad  , \s11_data_i[2]_pad  , \s11_data_i[30]_pad  , \s11_data_i[31]_pad  , \s11_data_i[3]_pad  , \s11_data_i[4]_pad  , \s11_data_i[5]_pad  , \s11_data_i[6]_pad  , \s11_data_i[7]_pad  , \s11_data_i[8]_pad  , \s11_data_i[9]_pad  , \s11_err_i_pad  , \s11_m0_cyc_r_reg/P0001  , \s11_m1_cyc_r_reg/P0001  , \s11_m2_cyc_r_reg/P0001  , \s11_m3_cyc_r_reg/P0001  , \s11_m4_cyc_r_reg/P0001  , \s11_m5_cyc_r_reg/P0001  , \s11_m6_cyc_r_reg/P0001  , \s11_m7_cyc_r_reg/P0001  , \s11_msel_arb0_state_reg[0]/NET0131  , \s11_msel_arb0_state_reg[1]/NET0131  , \s11_msel_arb0_state_reg[2]/NET0131  , \s11_msel_arb1_state_reg[0]/NET0131  , \s11_msel_arb1_state_reg[1]/NET0131  , \s11_msel_arb1_state_reg[2]/NET0131  , \s11_msel_arb2_state_reg[0]/NET0131  , \s11_msel_arb2_state_reg[1]/NET0131  , \s11_msel_arb2_state_reg[2]/NET0131  , \s11_msel_arb3_state_reg[0]/NET0131  , \s11_msel_arb3_state_reg[1]/NET0131  , \s11_msel_arb3_state_reg[2]/NET0131  , \s11_msel_pri_out_reg[0]/NET0131  , \s11_msel_pri_out_reg[1]/NET0131  , \s11_next_reg/P0001  , \s11_rty_i_pad  , \s12_ack_i_pad  , \s12_data_i[0]_pad  , \s12_data_i[10]_pad  , \s12_data_i[11]_pad  , \s12_data_i[12]_pad  , \s12_data_i[13]_pad  , \s12_data_i[14]_pad  , \s12_data_i[15]_pad  , \s12_data_i[16]_pad  , \s12_data_i[17]_pad  , \s12_data_i[18]_pad  , \s12_data_i[19]_pad  , \s12_data_i[1]_pad  , \s12_data_i[20]_pad  , \s12_data_i[21]_pad  , \s12_data_i[22]_pad  , \s12_data_i[23]_pad  , \s12_data_i[24]_pad  , \s12_data_i[25]_pad  , \s12_data_i[26]_pad  , \s12_data_i[27]_pad  , \s12_data_i[28]_pad  , \s12_data_i[29]_pad  , \s12_data_i[2]_pad  , \s12_data_i[30]_pad  , \s12_data_i[31]_pad  , \s12_data_i[3]_pad  , \s12_data_i[4]_pad  , \s12_data_i[5]_pad  , \s12_data_i[6]_pad  , \s12_data_i[7]_pad  , \s12_data_i[8]_pad  , \s12_data_i[9]_pad  , \s12_err_i_pad  , \s12_m0_cyc_r_reg/P0001  , \s12_m1_cyc_r_reg/P0001  , \s12_m2_cyc_r_reg/P0001  , \s12_m3_cyc_r_reg/P0001  , \s12_m4_cyc_r_reg/P0001  , \s12_m5_cyc_r_reg/P0001  , \s12_m6_cyc_r_reg/P0001  , \s12_m7_cyc_r_reg/P0001  , \s12_msel_arb0_state_reg[0]/NET0131  , \s12_msel_arb0_state_reg[1]/NET0131  , \s12_msel_arb0_state_reg[2]/NET0131  , \s12_msel_arb1_state_reg[0]/NET0131  , \s12_msel_arb1_state_reg[1]/NET0131  , \s12_msel_arb1_state_reg[2]/NET0131  , \s12_msel_arb2_state_reg[0]/NET0131  , \s12_msel_arb2_state_reg[1]/NET0131  , \s12_msel_arb2_state_reg[2]/NET0131  , \s12_msel_arb3_state_reg[0]/NET0131  , \s12_msel_arb3_state_reg[1]/NET0131  , \s12_msel_arb3_state_reg[2]/NET0131  , \s12_msel_pri_out_reg[0]/NET0131  , \s12_msel_pri_out_reg[1]/NET0131  , \s12_next_reg/P0001  , \s12_rty_i_pad  , \s13_ack_i_pad  , \s13_data_i[0]_pad  , \s13_data_i[10]_pad  , \s13_data_i[11]_pad  , \s13_data_i[12]_pad  , \s13_data_i[13]_pad  , \s13_data_i[14]_pad  , \s13_data_i[15]_pad  , \s13_data_i[16]_pad  , \s13_data_i[17]_pad  , \s13_data_i[18]_pad  , \s13_data_i[19]_pad  , \s13_data_i[1]_pad  , \s13_data_i[20]_pad  , \s13_data_i[21]_pad  , \s13_data_i[22]_pad  , \s13_data_i[23]_pad  , \s13_data_i[24]_pad  , \s13_data_i[25]_pad  , \s13_data_i[26]_pad  , \s13_data_i[27]_pad  , \s13_data_i[28]_pad  , \s13_data_i[29]_pad  , \s13_data_i[2]_pad  , \s13_data_i[30]_pad  , \s13_data_i[31]_pad  , \s13_data_i[3]_pad  , \s13_data_i[4]_pad  , \s13_data_i[5]_pad  , \s13_data_i[6]_pad  , \s13_data_i[7]_pad  , \s13_data_i[8]_pad  , \s13_data_i[9]_pad  , \s13_err_i_pad  , \s13_m0_cyc_r_reg/P0001  , \s13_m1_cyc_r_reg/P0001  , \s13_m2_cyc_r_reg/P0001  , \s13_m3_cyc_r_reg/P0001  , \s13_m4_cyc_r_reg/P0001  , \s13_m5_cyc_r_reg/P0001  , \s13_m6_cyc_r_reg/P0001  , \s13_m7_cyc_r_reg/P0001  , \s13_msel_arb0_state_reg[0]/NET0131  , \s13_msel_arb0_state_reg[1]/NET0131  , \s13_msel_arb0_state_reg[2]/NET0131  , \s13_msel_arb1_state_reg[0]/NET0131  , \s13_msel_arb1_state_reg[1]/NET0131  , \s13_msel_arb1_state_reg[2]/NET0131  , \s13_msel_arb2_state_reg[0]/NET0131  , \s13_msel_arb2_state_reg[1]/NET0131  , \s13_msel_arb2_state_reg[2]/NET0131  , \s13_msel_arb3_state_reg[0]/NET0131  , \s13_msel_arb3_state_reg[1]/NET0131  , \s13_msel_arb3_state_reg[2]/NET0131  , \s13_msel_pri_out_reg[0]/NET0131  , \s13_msel_pri_out_reg[1]/NET0131  , \s13_next_reg/P0001  , \s13_rty_i_pad  , \s14_ack_i_pad  , \s14_data_i[0]_pad  , \s14_data_i[10]_pad  , \s14_data_i[11]_pad  , \s14_data_i[12]_pad  , \s14_data_i[13]_pad  , \s14_data_i[14]_pad  , \s14_data_i[15]_pad  , \s14_data_i[16]_pad  , \s14_data_i[17]_pad  , \s14_data_i[18]_pad  , \s14_data_i[19]_pad  , \s14_data_i[1]_pad  , \s14_data_i[20]_pad  , \s14_data_i[21]_pad  , \s14_data_i[22]_pad  , \s14_data_i[23]_pad  , \s14_data_i[24]_pad  , \s14_data_i[25]_pad  , \s14_data_i[26]_pad  , \s14_data_i[27]_pad  , \s14_data_i[28]_pad  , \s14_data_i[29]_pad  , \s14_data_i[2]_pad  , \s14_data_i[30]_pad  , \s14_data_i[31]_pad  , \s14_data_i[3]_pad  , \s14_data_i[4]_pad  , \s14_data_i[5]_pad  , \s14_data_i[6]_pad  , \s14_data_i[7]_pad  , \s14_data_i[8]_pad  , \s14_data_i[9]_pad  , \s14_err_i_pad  , \s14_m0_cyc_r_reg/P0001  , \s14_m1_cyc_r_reg/P0001  , \s14_m2_cyc_r_reg/P0001  , \s14_m3_cyc_r_reg/P0001  , \s14_m4_cyc_r_reg/P0001  , \s14_m5_cyc_r_reg/P0001  , \s14_m6_cyc_r_reg/P0001  , \s14_m7_cyc_r_reg/P0001  , \s14_msel_arb0_state_reg[0]/NET0131  , \s14_msel_arb0_state_reg[1]/NET0131  , \s14_msel_arb0_state_reg[2]/NET0131  , \s14_msel_arb1_state_reg[0]/NET0131  , \s14_msel_arb1_state_reg[1]/NET0131  , \s14_msel_arb1_state_reg[2]/NET0131  , \s14_msel_arb2_state_reg[0]/NET0131  , \s14_msel_arb2_state_reg[1]/NET0131  , \s14_msel_arb2_state_reg[2]/NET0131  , \s14_msel_arb3_state_reg[0]/NET0131  , \s14_msel_arb3_state_reg[1]/NET0131  , \s14_msel_arb3_state_reg[2]/NET0131  , \s14_msel_pri_out_reg[0]/NET0131  , \s14_msel_pri_out_reg[1]/NET0131  , \s14_next_reg/P0001  , \s14_rty_i_pad  , \s15_ack_i_pad  , \s15_data_i[0]_pad  , \s15_data_i[10]_pad  , \s15_data_i[11]_pad  , \s15_data_i[12]_pad  , \s15_data_i[13]_pad  , \s15_data_i[14]_pad  , \s15_data_i[15]_pad  , \s15_data_i[16]_pad  , \s15_data_i[17]_pad  , \s15_data_i[18]_pad  , \s15_data_i[19]_pad  , \s15_data_i[1]_pad  , \s15_data_i[20]_pad  , \s15_data_i[21]_pad  , \s15_data_i[22]_pad  , \s15_data_i[23]_pad  , \s15_data_i[24]_pad  , \s15_data_i[25]_pad  , \s15_data_i[26]_pad  , \s15_data_i[27]_pad  , \s15_data_i[28]_pad  , \s15_data_i[29]_pad  , \s15_data_i[2]_pad  , \s15_data_i[30]_pad  , \s15_data_i[31]_pad  , \s15_data_i[3]_pad  , \s15_data_i[4]_pad  , \s15_data_i[5]_pad  , \s15_data_i[6]_pad  , \s15_data_i[7]_pad  , \s15_data_i[8]_pad  , \s15_data_i[9]_pad  , \s15_err_i_pad  , \s15_m0_cyc_r_reg/P0001  , \s15_m1_cyc_r_reg/P0001  , \s15_m2_cyc_r_reg/P0001  , \s15_m3_cyc_r_reg/P0001  , \s15_m4_cyc_r_reg/P0001  , \s15_m5_cyc_r_reg/P0001  , \s15_m6_cyc_r_reg/P0001  , \s15_m7_cyc_r_reg/P0001  , \s15_msel_arb0_state_reg[0]/NET0131  , \s15_msel_arb0_state_reg[1]/NET0131  , \s15_msel_arb0_state_reg[2]/NET0131  , \s15_msel_arb1_state_reg[0]/NET0131  , \s15_msel_arb1_state_reg[1]/NET0131  , \s15_msel_arb1_state_reg[2]/NET0131  , \s15_msel_arb2_state_reg[0]/NET0131  , \s15_msel_arb2_state_reg[1]/NET0131  , \s15_msel_arb2_state_reg[2]/NET0131  , \s15_msel_arb3_state_reg[0]/NET0131  , \s15_msel_arb3_state_reg[1]/NET0131  , \s15_msel_arb3_state_reg[2]/NET0131  , \s15_msel_pri_out_reg[0]/NET0131  , \s15_msel_pri_out_reg[1]/NET0131  , \s15_next_reg/P0001  , \s15_rty_i_pad  , \s1_ack_i_pad  , \s1_data_i[0]_pad  , \s1_data_i[10]_pad  , \s1_data_i[11]_pad  , \s1_data_i[12]_pad  , \s1_data_i[13]_pad  , \s1_data_i[14]_pad  , \s1_data_i[15]_pad  , \s1_data_i[16]_pad  , \s1_data_i[17]_pad  , \s1_data_i[18]_pad  , \s1_data_i[19]_pad  , \s1_data_i[1]_pad  , \s1_data_i[20]_pad  , \s1_data_i[21]_pad  , \s1_data_i[22]_pad  , \s1_data_i[23]_pad  , \s1_data_i[24]_pad  , \s1_data_i[25]_pad  , \s1_data_i[26]_pad  , \s1_data_i[27]_pad  , \s1_data_i[28]_pad  , \s1_data_i[29]_pad  , \s1_data_i[2]_pad  , \s1_data_i[30]_pad  , \s1_data_i[31]_pad  , \s1_data_i[3]_pad  , \s1_data_i[4]_pad  , \s1_data_i[5]_pad  , \s1_data_i[6]_pad  , \s1_data_i[7]_pad  , \s1_data_i[8]_pad  , \s1_data_i[9]_pad  , \s1_err_i_pad  , \s1_m0_cyc_r_reg/P0001  , \s1_m1_cyc_r_reg/P0001  , \s1_m2_cyc_r_reg/P0001  , \s1_m3_cyc_r_reg/P0001  , \s1_m4_cyc_r_reg/P0001  , \s1_m5_cyc_r_reg/P0001  , \s1_m6_cyc_r_reg/P0001  , \s1_m7_cyc_r_reg/P0001  , \s1_msel_arb0_state_reg[0]/NET0131  , \s1_msel_arb0_state_reg[1]/NET0131  , \s1_msel_arb0_state_reg[2]/NET0131  , \s1_msel_arb1_state_reg[0]/NET0131  , \s1_msel_arb1_state_reg[1]/NET0131  , \s1_msel_arb1_state_reg[2]/NET0131  , \s1_msel_arb2_state_reg[0]/NET0131  , \s1_msel_arb2_state_reg[1]/NET0131  , \s1_msel_arb2_state_reg[2]/NET0131  , \s1_msel_arb3_state_reg[0]/NET0131  , \s1_msel_arb3_state_reg[1]/NET0131  , \s1_msel_arb3_state_reg[2]/NET0131  , \s1_msel_pri_out_reg[0]/NET0131  , \s1_msel_pri_out_reg[1]/NET0131  , \s1_next_reg/P0001  , \s1_rty_i_pad  , \s2_ack_i_pad  , \s2_data_i[0]_pad  , \s2_data_i[10]_pad  , \s2_data_i[11]_pad  , \s2_data_i[12]_pad  , \s2_data_i[13]_pad  , \s2_data_i[14]_pad  , \s2_data_i[15]_pad  , \s2_data_i[16]_pad  , \s2_data_i[17]_pad  , \s2_data_i[18]_pad  , \s2_data_i[19]_pad  , \s2_data_i[1]_pad  , \s2_data_i[20]_pad  , \s2_data_i[21]_pad  , \s2_data_i[22]_pad  , \s2_data_i[23]_pad  , \s2_data_i[24]_pad  , \s2_data_i[25]_pad  , \s2_data_i[26]_pad  , \s2_data_i[27]_pad  , \s2_data_i[28]_pad  , \s2_data_i[29]_pad  , \s2_data_i[2]_pad  , \s2_data_i[30]_pad  , \s2_data_i[31]_pad  , \s2_data_i[3]_pad  , \s2_data_i[4]_pad  , \s2_data_i[5]_pad  , \s2_data_i[6]_pad  , \s2_data_i[7]_pad  , \s2_data_i[8]_pad  , \s2_data_i[9]_pad  , \s2_err_i_pad  , \s2_m0_cyc_r_reg/P0001  , \s2_m1_cyc_r_reg/P0001  , \s2_m2_cyc_r_reg/P0001  , \s2_m3_cyc_r_reg/P0001  , \s2_m4_cyc_r_reg/P0001  , \s2_m5_cyc_r_reg/P0001  , \s2_m6_cyc_r_reg/P0001  , \s2_m7_cyc_r_reg/P0001  , \s2_msel_arb0_state_reg[0]/NET0131  , \s2_msel_arb0_state_reg[1]/NET0131  , \s2_msel_arb0_state_reg[2]/NET0131  , \s2_msel_arb1_state_reg[0]/NET0131  , \s2_msel_arb1_state_reg[1]/NET0131  , \s2_msel_arb1_state_reg[2]/NET0131  , \s2_msel_arb2_state_reg[0]/NET0131  , \s2_msel_arb2_state_reg[1]/NET0131  , \s2_msel_arb2_state_reg[2]/NET0131  , \s2_msel_arb3_state_reg[0]/NET0131  , \s2_msel_arb3_state_reg[1]/NET0131  , \s2_msel_arb3_state_reg[2]/NET0131  , \s2_msel_pri_out_reg[0]/NET0131  , \s2_msel_pri_out_reg[1]/NET0131  , \s2_next_reg/P0001  , \s2_rty_i_pad  , \s3_ack_i_pad  , \s3_data_i[0]_pad  , \s3_data_i[10]_pad  , \s3_data_i[11]_pad  , \s3_data_i[12]_pad  , \s3_data_i[13]_pad  , \s3_data_i[14]_pad  , \s3_data_i[15]_pad  , \s3_data_i[16]_pad  , \s3_data_i[17]_pad  , \s3_data_i[18]_pad  , \s3_data_i[19]_pad  , \s3_data_i[1]_pad  , \s3_data_i[20]_pad  , \s3_data_i[21]_pad  , \s3_data_i[22]_pad  , \s3_data_i[23]_pad  , \s3_data_i[24]_pad  , \s3_data_i[25]_pad  , \s3_data_i[26]_pad  , \s3_data_i[27]_pad  , \s3_data_i[28]_pad  , \s3_data_i[29]_pad  , \s3_data_i[2]_pad  , \s3_data_i[30]_pad  , \s3_data_i[31]_pad  , \s3_data_i[3]_pad  , \s3_data_i[4]_pad  , \s3_data_i[5]_pad  , \s3_data_i[6]_pad  , \s3_data_i[7]_pad  , \s3_data_i[8]_pad  , \s3_data_i[9]_pad  , \s3_err_i_pad  , \s3_m0_cyc_r_reg/P0001  , \s3_m1_cyc_r_reg/P0001  , \s3_m2_cyc_r_reg/P0001  , \s3_m3_cyc_r_reg/P0001  , \s3_m4_cyc_r_reg/P0001  , \s3_m5_cyc_r_reg/P0001  , \s3_m6_cyc_r_reg/P0001  , \s3_m7_cyc_r_reg/P0001  , \s3_msel_arb0_state_reg[0]/NET0131  , \s3_msel_arb0_state_reg[1]/NET0131  , \s3_msel_arb0_state_reg[2]/NET0131  , \s3_msel_arb1_state_reg[0]/NET0131  , \s3_msel_arb1_state_reg[1]/NET0131  , \s3_msel_arb1_state_reg[2]/NET0131  , \s3_msel_arb2_state_reg[0]/NET0131  , \s3_msel_arb2_state_reg[1]/NET0131  , \s3_msel_arb2_state_reg[2]/NET0131  , \s3_msel_arb3_state_reg[0]/NET0131  , \s3_msel_arb3_state_reg[1]/NET0131  , \s3_msel_arb3_state_reg[2]/NET0131  , \s3_msel_pri_out_reg[0]/NET0131  , \s3_msel_pri_out_reg[1]/NET0131  , \s3_next_reg/P0001  , \s3_rty_i_pad  , \s4_ack_i_pad  , \s4_data_i[0]_pad  , \s4_data_i[10]_pad  , \s4_data_i[11]_pad  , \s4_data_i[12]_pad  , \s4_data_i[13]_pad  , \s4_data_i[14]_pad  , \s4_data_i[15]_pad  , \s4_data_i[16]_pad  , \s4_data_i[17]_pad  , \s4_data_i[18]_pad  , \s4_data_i[19]_pad  , \s4_data_i[1]_pad  , \s4_data_i[20]_pad  , \s4_data_i[21]_pad  , \s4_data_i[22]_pad  , \s4_data_i[23]_pad  , \s4_data_i[24]_pad  , \s4_data_i[25]_pad  , \s4_data_i[26]_pad  , \s4_data_i[27]_pad  , \s4_data_i[28]_pad  , \s4_data_i[29]_pad  , \s4_data_i[2]_pad  , \s4_data_i[30]_pad  , \s4_data_i[31]_pad  , \s4_data_i[3]_pad  , \s4_data_i[4]_pad  , \s4_data_i[5]_pad  , \s4_data_i[6]_pad  , \s4_data_i[7]_pad  , \s4_data_i[8]_pad  , \s4_data_i[9]_pad  , \s4_err_i_pad  , \s4_m0_cyc_r_reg/P0001  , \s4_m1_cyc_r_reg/P0001  , \s4_m2_cyc_r_reg/P0001  , \s4_m3_cyc_r_reg/P0001  , \s4_m4_cyc_r_reg/P0001  , \s4_m5_cyc_r_reg/P0001  , \s4_m6_cyc_r_reg/P0001  , \s4_m7_cyc_r_reg/P0001  , \s4_msel_arb0_state_reg[0]/NET0131  , \s4_msel_arb0_state_reg[1]/NET0131  , \s4_msel_arb0_state_reg[2]/NET0131  , \s4_msel_arb1_state_reg[0]/NET0131  , \s4_msel_arb1_state_reg[1]/NET0131  , \s4_msel_arb1_state_reg[2]/NET0131  , \s4_msel_arb2_state_reg[0]/NET0131  , \s4_msel_arb2_state_reg[1]/NET0131  , \s4_msel_arb2_state_reg[2]/NET0131  , \s4_msel_arb3_state_reg[0]/NET0131  , \s4_msel_arb3_state_reg[1]/NET0131  , \s4_msel_arb3_state_reg[2]/NET0131  , \s4_msel_pri_out_reg[0]/NET0131  , \s4_msel_pri_out_reg[1]/NET0131  , \s4_next_reg/P0001  , \s4_rty_i_pad  , \s5_ack_i_pad  , \s5_data_i[0]_pad  , \s5_data_i[10]_pad  , \s5_data_i[11]_pad  , \s5_data_i[12]_pad  , \s5_data_i[13]_pad  , \s5_data_i[14]_pad  , \s5_data_i[15]_pad  , \s5_data_i[16]_pad  , \s5_data_i[17]_pad  , \s5_data_i[18]_pad  , \s5_data_i[19]_pad  , \s5_data_i[1]_pad  , \s5_data_i[20]_pad  , \s5_data_i[21]_pad  , \s5_data_i[22]_pad  , \s5_data_i[23]_pad  , \s5_data_i[24]_pad  , \s5_data_i[25]_pad  , \s5_data_i[26]_pad  , \s5_data_i[27]_pad  , \s5_data_i[28]_pad  , \s5_data_i[29]_pad  , \s5_data_i[2]_pad  , \s5_data_i[30]_pad  , \s5_data_i[31]_pad  , \s5_data_i[3]_pad  , \s5_data_i[4]_pad  , \s5_data_i[5]_pad  , \s5_data_i[6]_pad  , \s5_data_i[7]_pad  , \s5_data_i[8]_pad  , \s5_data_i[9]_pad  , \s5_err_i_pad  , \s5_m0_cyc_r_reg/P0001  , \s5_m1_cyc_r_reg/P0001  , \s5_m2_cyc_r_reg/P0001  , \s5_m3_cyc_r_reg/P0001  , \s5_m4_cyc_r_reg/P0001  , \s5_m5_cyc_r_reg/P0001  , \s5_m6_cyc_r_reg/P0001  , \s5_m7_cyc_r_reg/P0001  , \s5_msel_arb0_state_reg[0]/NET0131  , \s5_msel_arb0_state_reg[1]/NET0131  , \s5_msel_arb0_state_reg[2]/NET0131  , \s5_msel_arb1_state_reg[0]/NET0131  , \s5_msel_arb1_state_reg[1]/NET0131  , \s5_msel_arb1_state_reg[2]/NET0131  , \s5_msel_arb2_state_reg[0]/NET0131  , \s5_msel_arb2_state_reg[1]/NET0131  , \s5_msel_arb2_state_reg[2]/NET0131  , \s5_msel_arb3_state_reg[0]/NET0131  , \s5_msel_arb3_state_reg[1]/NET0131  , \s5_msel_arb3_state_reg[2]/NET0131  , \s5_msel_pri_out_reg[0]/NET0131  , \s5_msel_pri_out_reg[1]/NET0131  , \s5_next_reg/P0001  , \s5_rty_i_pad  , \s6_ack_i_pad  , \s6_data_i[0]_pad  , \s6_data_i[10]_pad  , \s6_data_i[11]_pad  , \s6_data_i[12]_pad  , \s6_data_i[13]_pad  , \s6_data_i[14]_pad  , \s6_data_i[15]_pad  , \s6_data_i[16]_pad  , \s6_data_i[17]_pad  , \s6_data_i[18]_pad  , \s6_data_i[19]_pad  , \s6_data_i[1]_pad  , \s6_data_i[20]_pad  , \s6_data_i[21]_pad  , \s6_data_i[22]_pad  , \s6_data_i[23]_pad  , \s6_data_i[24]_pad  , \s6_data_i[25]_pad  , \s6_data_i[26]_pad  , \s6_data_i[27]_pad  , \s6_data_i[28]_pad  , \s6_data_i[29]_pad  , \s6_data_i[2]_pad  , \s6_data_i[30]_pad  , \s6_data_i[31]_pad  , \s6_data_i[3]_pad  , \s6_data_i[4]_pad  , \s6_data_i[5]_pad  , \s6_data_i[6]_pad  , \s6_data_i[7]_pad  , \s6_data_i[8]_pad  , \s6_data_i[9]_pad  , \s6_err_i_pad  , \s6_m0_cyc_r_reg/P0001  , \s6_m1_cyc_r_reg/P0001  , \s6_m2_cyc_r_reg/P0001  , \s6_m3_cyc_r_reg/P0001  , \s6_m4_cyc_r_reg/P0001  , \s6_m5_cyc_r_reg/P0001  , \s6_m6_cyc_r_reg/P0001  , \s6_m7_cyc_r_reg/P0001  , \s6_msel_arb0_state_reg[0]/NET0131  , \s6_msel_arb0_state_reg[1]/NET0131  , \s6_msel_arb0_state_reg[2]/NET0131  , \s6_msel_arb1_state_reg[0]/NET0131  , \s6_msel_arb1_state_reg[1]/NET0131  , \s6_msel_arb1_state_reg[2]/NET0131  , \s6_msel_arb2_state_reg[0]/NET0131  , \s6_msel_arb2_state_reg[1]/NET0131  , \s6_msel_arb2_state_reg[2]/NET0131  , \s6_msel_arb3_state_reg[0]/NET0131  , \s6_msel_arb3_state_reg[1]/NET0131  , \s6_msel_arb3_state_reg[2]/NET0131  , \s6_msel_pri_out_reg[0]/NET0131  , \s6_msel_pri_out_reg[1]/NET0131  , \s6_next_reg/P0001  , \s6_rty_i_pad  , \s7_ack_i_pad  , \s7_data_i[0]_pad  , \s7_data_i[10]_pad  , \s7_data_i[11]_pad  , \s7_data_i[12]_pad  , \s7_data_i[13]_pad  , \s7_data_i[14]_pad  , \s7_data_i[15]_pad  , \s7_data_i[16]_pad  , \s7_data_i[17]_pad  , \s7_data_i[18]_pad  , \s7_data_i[19]_pad  , \s7_data_i[1]_pad  , \s7_data_i[20]_pad  , \s7_data_i[21]_pad  , \s7_data_i[22]_pad  , \s7_data_i[23]_pad  , \s7_data_i[24]_pad  , \s7_data_i[25]_pad  , \s7_data_i[26]_pad  , \s7_data_i[27]_pad  , \s7_data_i[28]_pad  , \s7_data_i[29]_pad  , \s7_data_i[2]_pad  , \s7_data_i[30]_pad  , \s7_data_i[31]_pad  , \s7_data_i[3]_pad  , \s7_data_i[4]_pad  , \s7_data_i[5]_pad  , \s7_data_i[6]_pad  , \s7_data_i[7]_pad  , \s7_data_i[8]_pad  , \s7_data_i[9]_pad  , \s7_err_i_pad  , \s7_m0_cyc_r_reg/P0001  , \s7_m1_cyc_r_reg/P0001  , \s7_m2_cyc_r_reg/P0001  , \s7_m3_cyc_r_reg/P0001  , \s7_m4_cyc_r_reg/P0001  , \s7_m5_cyc_r_reg/P0001  , \s7_m6_cyc_r_reg/P0001  , \s7_m7_cyc_r_reg/P0001  , \s7_msel_arb0_state_reg[0]/NET0131  , \s7_msel_arb0_state_reg[1]/NET0131  , \s7_msel_arb0_state_reg[2]/NET0131  , \s7_msel_arb1_state_reg[0]/NET0131  , \s7_msel_arb1_state_reg[1]/NET0131  , \s7_msel_arb1_state_reg[2]/NET0131  , \s7_msel_arb2_state_reg[0]/NET0131  , \s7_msel_arb2_state_reg[1]/NET0131  , \s7_msel_arb2_state_reg[2]/NET0131  , \s7_msel_arb3_state_reg[0]/NET0131  , \s7_msel_arb3_state_reg[1]/NET0131  , \s7_msel_arb3_state_reg[2]/NET0131  , \s7_msel_pri_out_reg[0]/NET0131  , \s7_msel_pri_out_reg[1]/NET0131  , \s7_next_reg/P0001  , \s7_rty_i_pad  , \s8_ack_i_pad  , \s8_data_i[0]_pad  , \s8_data_i[10]_pad  , \s8_data_i[11]_pad  , \s8_data_i[12]_pad  , \s8_data_i[13]_pad  , \s8_data_i[14]_pad  , \s8_data_i[15]_pad  , \s8_data_i[16]_pad  , \s8_data_i[17]_pad  , \s8_data_i[18]_pad  , \s8_data_i[19]_pad  , \s8_data_i[1]_pad  , \s8_data_i[20]_pad  , \s8_data_i[21]_pad  , \s8_data_i[22]_pad  , \s8_data_i[23]_pad  , \s8_data_i[24]_pad  , \s8_data_i[25]_pad  , \s8_data_i[26]_pad  , \s8_data_i[27]_pad  , \s8_data_i[28]_pad  , \s8_data_i[29]_pad  , \s8_data_i[2]_pad  , \s8_data_i[30]_pad  , \s8_data_i[31]_pad  , \s8_data_i[3]_pad  , \s8_data_i[4]_pad  , \s8_data_i[5]_pad  , \s8_data_i[6]_pad  , \s8_data_i[7]_pad  , \s8_data_i[8]_pad  , \s8_data_i[9]_pad  , \s8_err_i_pad  , \s8_m0_cyc_r_reg/P0001  , \s8_m1_cyc_r_reg/P0001  , \s8_m2_cyc_r_reg/P0001  , \s8_m3_cyc_r_reg/P0001  , \s8_m4_cyc_r_reg/P0001  , \s8_m5_cyc_r_reg/P0001  , \s8_m6_cyc_r_reg/P0001  , \s8_m7_cyc_r_reg/P0001  , \s8_msel_arb0_state_reg[0]/NET0131  , \s8_msel_arb0_state_reg[1]/NET0131  , \s8_msel_arb0_state_reg[2]/NET0131  , \s8_msel_arb1_state_reg[0]/NET0131  , \s8_msel_arb1_state_reg[1]/NET0131  , \s8_msel_arb1_state_reg[2]/NET0131  , \s8_msel_arb2_state_reg[0]/NET0131  , \s8_msel_arb2_state_reg[1]/NET0131  , \s8_msel_arb2_state_reg[2]/NET0131  , \s8_msel_arb3_state_reg[0]/NET0131  , \s8_msel_arb3_state_reg[1]/NET0131  , \s8_msel_arb3_state_reg[2]/NET0131  , \s8_msel_pri_out_reg[0]/NET0131  , \s8_msel_pri_out_reg[1]/NET0131  , \s8_next_reg/P0001  , \s8_rty_i_pad  , \s9_ack_i_pad  , \s9_data_i[0]_pad  , \s9_data_i[10]_pad  , \s9_data_i[11]_pad  , \s9_data_i[12]_pad  , \s9_data_i[13]_pad  , \s9_data_i[14]_pad  , \s9_data_i[15]_pad  , \s9_data_i[16]_pad  , \s9_data_i[17]_pad  , \s9_data_i[18]_pad  , \s9_data_i[19]_pad  , \s9_data_i[1]_pad  , \s9_data_i[20]_pad  , \s9_data_i[21]_pad  , \s9_data_i[22]_pad  , \s9_data_i[23]_pad  , \s9_data_i[24]_pad  , \s9_data_i[25]_pad  , \s9_data_i[26]_pad  , \s9_data_i[27]_pad  , \s9_data_i[28]_pad  , \s9_data_i[29]_pad  , \s9_data_i[2]_pad  , \s9_data_i[30]_pad  , \s9_data_i[31]_pad  , \s9_data_i[3]_pad  , \s9_data_i[4]_pad  , \s9_data_i[5]_pad  , \s9_data_i[6]_pad  , \s9_data_i[7]_pad  , \s9_data_i[8]_pad  , \s9_data_i[9]_pad  , \s9_err_i_pad  , \s9_m0_cyc_r_reg/P0001  , \s9_m1_cyc_r_reg/P0001  , \s9_m2_cyc_r_reg/P0001  , \s9_m3_cyc_r_reg/P0001  , \s9_m4_cyc_r_reg/P0001  , \s9_m5_cyc_r_reg/P0001  , \s9_m6_cyc_r_reg/P0001  , \s9_m7_cyc_r_reg/P0001  , \s9_msel_arb0_state_reg[0]/NET0131  , \s9_msel_arb0_state_reg[1]/NET0131  , \s9_msel_arb0_state_reg[2]/NET0131  , \s9_msel_arb1_state_reg[0]/NET0131  , \s9_msel_arb1_state_reg[1]/NET0131  , \s9_msel_arb1_state_reg[2]/NET0131  , \s9_msel_arb2_state_reg[0]/NET0131  , \s9_msel_arb2_state_reg[1]/NET0131  , \s9_msel_arb2_state_reg[2]/NET0131  , \s9_msel_arb3_state_reg[0]/NET0131  , \s9_msel_arb3_state_reg[1]/NET0131  , \s9_msel_arb3_state_reg[2]/NET0131  , \s9_msel_pri_out_reg[0]/NET0131  , \s9_msel_pri_out_reg[1]/NET0131  , \s9_next_reg/P0001  , \s9_rty_i_pad  , \_al_n0  , \_al_n1  , \g106655/_1_  , \g106703/_1_  , \g69412/_0_  , \g69413/_0_  , \g69417/_1_  , \g69418/_0_  , \g69420/_1_  , \g69421/_0_  , \g69423/_1_  , \g69424/_0_  , \g69426/_1_  , \g69428/_1_  , \g69430/_1_  , \g69432/_1_  , \g69434/_1_  , \g69436/_1_  , \g69438/_1_  , \g69757/_2_  , \g69758/_2_  , \g69759/_2_  , \g69760/_2_  , \g69761/_0_  , \g69762/_2_  , \g69763/_2_  , \g69764/_2_  , \g69765/_2_  , \g69766/_2_  , \g69767/_0_  , \g69768/_0_  , \g69769/_0_  , \g69770/_0_  , \g69771/_0_  , \g69772/_0_  , \g70206/_0_  , \g70392/_0_  , \g70393/_0_  , \g70394/_0_  , \g70395/_0_  , \g70396/_0_  , \g70397/_0_  , \g70398/_0_  , \g70399/_0_  , \g70400/_0_  , \g70401/_0_  , \g70402/_0_  , \g70403/_0_  , \g70404/_0_  , \g70405/_0_  , \g70406/_0_  , \g70407/_0_  , \g70408/_0_  , \g70409/_0_  , \g70410/_0_  , \g70411/_0_  , \g70412/_0_  , \g70413/_0_  , \g70414/_0_  , \g70415/_0_  , \g70416/_0_  , \g70417/_0_  , \g70418/_0_  , \g70419/_0_  , \g70420/_0_  , \g70421/_0_  , \g70422/_0_  , \g70423/_0_  , \g70424/_0_  , \g70425/_0_  , \g70426/_0_  , \g70427/_0_  , \g70428/_0_  , \g70429/_0_  , \g70430/_0_  , \g70431/_0_  , \g70432/_0_  , \g70433/_0_  , \g70434/_0_  , \g70435/_0_  , \g70436/_0_  , \g70437/_0_  , \g70438/_0_  , \g70439/_0_  , \g70440/_0_  , \g70441/_0_  , \g70442/_0_  , \g70443/_0_  , \g70444/_0_  , \g70445/_0_  , \g70446/_0_  , \g70447/_0_  , \g70448/_0_  , \g70449/_0_  , \g70450/_0_  , \g70451/_0_  , \g70452/_0_  , \g70453/_0_  , \g70454/_0_  , \g70455/_0_  , \g70456/_0_  , \g70457/_0_  , \g70458/_0_  , \g70459/_0_  , \g70460/_0_  , \g70461/_0_  , \g70462/_0_  , \g70463/_0_  , \g70464/_0_  , \g70465/_0_  , \g70466/_0_  , \g70467/_0_  , \g70468/_0_  , \g70469/_0_  , \g70470/_0_  , \g70471/_0_  , \g70472/_0_  , \g70473/_0_  , \g70474/_0_  , \g70475/_0_  , \g70476/_0_  , \g70477/_0_  , \g70478/_0_  , \g70479/_0_  , \g70480/_0_  , \g70481/_0_  , \g70482/_0_  , \g70483/_0_  , \g70484/_0_  , \g70485/_0_  , \g70486/_0_  , \g70487/_0_  , \g70488/_0_  , \g70489/_0_  , \g70490/_0_  , \g70491/_0_  , \g70492/_0_  , \g70493/_0_  , \g70494/_0_  , \g70495/_0_  , \g70496/_0_  , \g70497/_0_  , \g70498/_0_  , \g70499/_0_  , \g70500/_0_  , \g70501/_0_  , \g70502/_0_  , \g70503/_0_  , \g70504/_0_  , \g70505/_0_  , \g70506/_0_  , \g70507/_0_  , \g70508/_0_  , \g70509/_0_  , \g70510/_0_  , \g70511/_0_  , \g70513/_0_  , \g70515/_0_  , \g70516/_0_  , \g70517/_0_  , \g70518/_0_  , \g70519/_0_  , \g70521/_0_  , \g70522/_0_  , \g70524/_0_  , \g70557/_0_  , \g70559/_0_  , \g70560/_0_  , \g70561/_0_  , \g70562/_0_  , \g70563/_0_  , \g70564/_0_  , \g70565/_0_  , \g70566/_0_  , \g70567/_0_  , \g70568/_0_  , \g70569/_0_  , \g70570/_0_  , \g70571/_0_  , \g70572/_0_  , \g70573/_0_  , \g70574/_0_  , \g70575/_0_  , \g70576/_0_  , \g70577/_0_  , \g70578/_0_  , \g70579/_0_  , \g70580/_0_  , \g70581/_0_  , \g70582/_0_  , \g70583/_0_  , \g70584/_0_  , \g70585/_0_  , \g70586/_0_  , \g70587/_0_  , \g70588/_0_  , \g70589/_0_  , \g70590/_0_  , \g70591/_0_  , \g70592/_0_  , \g70593/_0_  , \g70594/_0_  , \g70595/_0_  , \g70596/_0_  , \g70597/_0_  , \g70598/_0_  , \g70599/_0_  , \g70600/_0_  , \g70601/_0_  , \g70602/_0_  , \g70603/_0_  , \g70604/_0_  , \g70605/_0_  , \g70606/_0_  , \g70607/_0_  , \g70608/_0_  , \g70609/_0_  , \g70610/_0_  , \g70611/_0_  , \g70612/_0_  , \g70613/_0_  , \g70614/_0_  , \g70615/_0_  , \g70616/_0_  , \g70617/_0_  , \g70618/_0_  , \g70619/_0_  , \g70620/_0_  , \g70621/_0_  , \g70622/_0_  , \g70623/_0_  , \g70624/_0_  , \g70625/_0_  , \g70626/_0_  , \g70627/_0_  , \g70628/_0_  , \g70629/_0_  , \g70630/_0_  , \g70631/_0_  , \g70632/_0_  , \g70633/_0_  , \g70634/_0_  , \g70635/_0_  , \g70636/_0_  , \g70637/_0_  , \g70638/_0_  , \g70639/_0_  , \g70640/_0_  , \g70641/_0_  , \g70642/_0_  , \g70643/_0_  , \g70644/_0_  , \g70645/_0_  , \g70646/_0_  , \g70647/_0_  , \g70648/_0_  , \g70649/_0_  , \g70650/_0_  , \g70651/_0_  , \g70652/_0_  , \g70653/_0_  , \g70654/_0_  , \g70655/_0_  , \g70656/_0_  , \g70657/_0_  , \g70658/_0_  , \g70659/_0_  , \g70660/_0_  , \g70661/_0_  , \g70662/_0_  , \g70663/_0_  , \g70664/_0_  , \g70665/_0_  , \g70666/_0_  , \g70667/_0_  , \g70668/_0_  , \g70669/_0_  , \g70670/_0_  , \g70671/_0_  , \g70672/_0_  , \g70673/_0_  , \g70674/_0_  , \g70675/_0_  , \g70676/_0_  , \g70677/_0_  , \g70678/_0_  , \g70679/_0_  , \g70680/_0_  , \g70681/_0_  , \g70682/_0_  , \g70683/_0_  , \g70684/_0_  , \g70685/_0_  , \g70686/_0_  , \g70687/_0_  , \g70688/_0_  , \g70689/_0_  , \g70690/_0_  , \g70691/_0_  , \g70692/_0_  , \g70693/_0_  , \g70694/_0_  , \g70695/_0_  , \g70696/_0_  , \g70697/_0_  , \g70698/_0_  , \g70699/_0_  , \g70700/_0_  , \g70701/_0_  , \g70702/_0_  , \g70703/_0_  , \g70704/_0_  , \g70705/_0_  , \g70706/_0_  , \g70707/_0_  , \g70708/_0_  , \g70709/_0_  , \g70710/_0_  , \g70711/_0_  , \g70712/_0_  , \g70713/_0_  , \g70714/_0_  , \g70715/_0_  , \g70716/_0_  , \g70717/_0_  , \g70718/_0_  , \g70719/_0_  , \g70720/_0_  , \g70721/_0_  , \g70722/_0_  , \g70723/_0_  , \g70724/_0_  , \g70725/_0_  , \g70726/_0_  , \g70727/_0_  , \g70728/_0_  , \g70729/_0_  , \g70730/_0_  , \g70731/_0_  , \g70732/_0_  , \g70733/_0_  , \g70734/_0_  , \g70735/_0_  , \g70736/_0_  , \g70737/_0_  , \g70738/_0_  , \g70739/_0_  , \g70740/_0_  , \g70741/_0_  , \g70742/_0_  , \g70743/_0_  , \g70744/_0_  , \g70745/_0_  , \g70746/_0_  , \g70747/_0_  , \g70748/_0_  , \g70749/_0_  , \g70750/_0_  , \g70751/_0_  , \g70752/_0_  , \g70753/_0_  , \g70754/_0_  , \g70755/_0_  , \g70756/_0_  , \g70757/_0_  , \g70758/_0_  , \g70759/_0_  , \g70760/_0_  , \g70761/_0_  , \g70762/_0_  , \g70763/_0_  , \g70764/_0_  , \g70765/_0_  , \g70766/_0_  , \g70767/_0_  , \g70768/_0_  , \g70769/_0_  , \g70770/_0_  , \g70771/_0_  , \g70772/_0_  , \g70773/_0_  , \g70774/_0_  , \g70775/_0_  , \g70776/_0_  , \g70777/_0_  , \g70778/_0_  , \g70779/_0_  , \g70780/_0_  , \g70781/_0_  , \g70782/_0_  , \g70783/_0_  , \g70784/_0_  , \g70785/_0_  , \g70786/_0_  , \g70787/_0_  , \g70788/_0_  , \g70789/_0_  , \g70790/_0_  , \g70791/_0_  , \g70792/_0_  , \g70793/_0_  , \g70794/_0_  , \g70795/_0_  , \g70796/_0_  , \g70797/_0_  , \g70798/_0_  , \g70799/_0_  , \g70800/_0_  , \g70801/_0_  , \g70802/_0_  , \g70803/_0_  , \g70804/_0_  , \g70805/_0_  , \g70806/_0_  , \g70807/_0_  , \g70808/_0_  , \g70809/_0_  , \g70810/_0_  , \g70811/_0_  , \g70812/_0_  , \g70813/_0_  , \g70814/_0_  , \g70815/_0_  , \g70816/_0_  , \g70817/_0_  , \g70818/_0_  , \g70819/_0_  , \g70820/_0_  , \g70821/_0_  , \g70822/_0_  , \g70823/_0_  , \g70824/_0_  , \g70825/_0_  , \g70826/_0_  , \g70827/_0_  , \g70828/_0_  , \g70829/_0_  , \g70830/_0_  , \g70831/_0_  , \g70832/_0_  , \g70833/_0_  , \g70834/_0_  , \g70835/_0_  , \g70836/_0_  , \g70837/_0_  , \g70838/_0_  , \g70839/_0_  , \g70840/_0_  , \g70841/_0_  , \g70842/_0_  , \g70843/_0_  , \g70844/_0_  , \g70845/_0_  , \g70846/_0_  , \g70847/_0_  , \g70848/_0_  , \g70849/_0_  , \g70850/_0_  , \g70851/_0_  , \g70852/_0_  , \g70853/_0_  , \g70854/_0_  , \g70855/_0_  , \g70856/_0_  , \g70857/_0_  , \g70858/_0_  , \g70859/_0_  , \g70860/_0_  , \g70861/_0_  , \g71404/_0_  , \g71407/_0_  , \g72631/_0_  , \g72631/_1_  , \g72633/_0_  , \g72642/_0_  , \g72649/_0_  , \g72649/_1_  , \g72652/_0_  , \g72660/_0_  , \g72666/_0_  , \g72666/_1_  , \g72671/_0_  , \g72681/_0_  , \g72681/_1_  , \g72689/_0_  , \g72696/_0_  , \g72696/_1_  , \g72698/_0_  , \g72707/_0_  , \g72715/_0_  , \g72715/_1_  , \g72718/_0_  , \g72726/_0_  , \g72732/_0_  , \g72732/_1_  , \g72736/_0_  , \g72743/_0_  , \g72745/_0_  , \g72745/_1_  , \g72752/_0_  , \g72752/_1_  , \g72756/_0_  , \g72763/_0_  , \g72763/_1_  , \g72765/_0_  , \g72767/_0_  , \g72767/_1_  , \g72769/_0_  , \g72769/_1_  , \g72772/_0_  , \g72772/_1_  , \g72774/_0_  , \g72774/_1_  , \g72790/_0_  , \g72790/_1_  , \g72797/_0_  , \g73807/_0_  , \g73820/_0_  , \g73832/_0_  , \g73844/_0_  , \g73856/_0_  , \g73871/_0_  , \g73883/_0_  , \g73895/_0_  , \g73905/_3_  , \g73910/_0_  , \g73922/_0_  , \g73934/_0_  , \g73946/_0_  , \g73958/_0_  , \g73970/_0_  , \g73982/_0_  , \g87036/_0_  , \g87042/_0_  , \g87043/_0_  , \g87044/_0_  , \g87045/_0_  , \g87046/_0_  , \g87047/_0_  , \g87048/_0_  , \g87049/_0_  , \g87050/_0_  , \g87051/_0_  , \g87052/_0_  , \g87053/_0_  , \g87054/_0_  , \g87055/_0_  , \g87062/_0_  , \g88572/_0_  , \g88681/_0_  , \g88682/_0_  , \g88683/_0_  , \g88684/_0_  , \g88685/_0_  , \g88686/_0_  , \g88687/_0_  , \g88688/_0_  , \g88689/_0_  , \g88690/_0_  , \g88691/_0_  , \g88692/_0_  , \g88693/_0_  , \g88695/_0_  , \g88697/_0_  , \g88698/_0_  , \g88700/_0_  , \g88701/_0_  , \g88703/_0_  , \g88704/_0_  , \g88705/_0_  , \g88706/_0_  , \g88707/_0_  , \g88709/_0_  , \g88710/_0_  , \g88711/_0_  , \g88712/_0_  , \g88713/_0_  , \g88714/_0_  , \g88716/_0_  , \g88717/_0_  , \g88718/_0_  , \g88719/_0_  , \g88720/_0_  , \g88722/_0_  , \g88723/_0_  , \g88724/_0_  , \g88725/_0_  , \g88726/_0_  , \g88727/_0_  , \g88728/_0_  , \g88729/_0_  , \g88731/_0_  , \g88732/_0_  , \g88733/_0_  , \g88734/_0_  , \g88736/_0_  , \g88737/_0_  , \g88738/_0_  , \g88739/_0_  , \g88740/_0_  , \g88741/_0_  , \g88742/_0_  , \g88743/_0_  , \g88744/_0_  , \g88745/_0_  , \g88746/_0_  , \g88748/_0_  , \g88749/_0_  , \g88750/_0_  , \g88752/_0_  , \g88753/_0_  , \g88754/_0_  , \g88755/_0_  , \g88756/_0_  , \g88757/_0_  , \g88759/_0_  , \g88760/_0_  , \g88761/_0_  , \g88762/_0_  , \g88764/_0_  , \g88765/_0_  , \g88766/_0_  , \g88768/_0_  , \g88769/_0_  , \g88770/_0_  , \g88771/_0_  , \g88772/_0_  , \g88773/_0_  , \g88775/_0_  , \g88776/_0_  , \g88777/_0_  , \g88778/_0_  , \g88779/_0_  , \g88780/_0_  , \g88782/_0_  , \g88783/_0_  , \g88784/_0_  , \g88785/_0_  , \g88786/_0_  , \g88787/_0_  , \g88789/_0_  , \g88790/_0_  , \g88791/_0_  , \g88792/_0_  , \g88793/_0_  , \g88795/_0_  , \g88796/_0_  , \g88797/_0_  , \g88799/_0_  , \g88800/_0_  , \g88801/_0_  , \g88802/_0_  , \g88806/_0_  , \g88807/_0_  , \g88808/_0_  , \g88809/_0_  , \g88810/_0_  , \g88813/_0_  , \g88814/_0_  , \g88815/_0_  , \m0_ack_o_pad  , \m0_data_o[0]_pad  , \m0_data_o[10]_pad  , \m0_data_o[11]_pad  , \m0_data_o[12]_pad  , \m0_data_o[13]_pad  , \m0_data_o[14]_pad  , \m0_data_o[15]_pad  , \m0_data_o[16]_pad  , \m0_data_o[17]_pad  , \m0_data_o[18]_pad  , \m0_data_o[19]_pad  , \m0_data_o[1]_pad  , \m0_data_o[20]_pad  , \m0_data_o[21]_pad  , \m0_data_o[22]_pad  , \m0_data_o[23]_pad  , \m0_data_o[24]_pad  , \m0_data_o[25]_pad  , \m0_data_o[26]_pad  , \m0_data_o[27]_pad  , \m0_data_o[28]_pad  , \m0_data_o[29]_pad  , \m0_data_o[2]_pad  , \m0_data_o[30]_pad  , \m0_data_o[31]_pad  , \m0_data_o[3]_pad  , \m0_data_o[4]_pad  , \m0_data_o[5]_pad  , \m0_data_o[6]_pad  , \m0_data_o[7]_pad  , \m0_data_o[8]_pad  , \m0_data_o[9]_pad  , \m0_err_o_pad  , \m0_rty_o_pad  , \m1_ack_o_pad  , \m1_data_o[0]_pad  , \m1_data_o[10]_pad  , \m1_data_o[11]_pad  , \m1_data_o[12]_pad  , \m1_data_o[13]_pad  , \m1_data_o[14]_pad  , \m1_data_o[15]_pad  , \m1_data_o[16]_pad  , \m1_data_o[17]_pad  , \m1_data_o[18]_pad  , \m1_data_o[19]_pad  , \m1_data_o[1]_pad  , \m1_data_o[20]_pad  , \m1_data_o[21]_pad  , \m1_data_o[22]_pad  , \m1_data_o[23]_pad  , \m1_data_o[24]_pad  , \m1_data_o[25]_pad  , \m1_data_o[26]_pad  , \m1_data_o[27]_pad  , \m1_data_o[28]_pad  , \m1_data_o[29]_pad  , \m1_data_o[2]_pad  , \m1_data_o[30]_pad  , \m1_data_o[31]_pad  , \m1_data_o[3]_pad  , \m1_data_o[4]_pad  , \m1_data_o[5]_pad  , \m1_data_o[6]_pad  , \m1_data_o[7]_pad  , \m1_data_o[8]_pad  , \m1_data_o[9]_pad  , \m1_err_o_pad  , \m1_rty_o_pad  , \m2_ack_o_pad  , \m2_data_o[0]_pad  , \m2_data_o[10]_pad  , \m2_data_o[11]_pad  , \m2_data_o[12]_pad  , \m2_data_o[13]_pad  , \m2_data_o[14]_pad  , \m2_data_o[15]_pad  , \m2_data_o[16]_pad  , \m2_data_o[17]_pad  , \m2_data_o[18]_pad  , \m2_data_o[19]_pad  , \m2_data_o[1]_pad  , \m2_data_o[20]_pad  , \m2_data_o[21]_pad  , \m2_data_o[22]_pad  , \m2_data_o[23]_pad  , \m2_data_o[24]_pad  , \m2_data_o[25]_pad  , \m2_data_o[26]_pad  , \m2_data_o[27]_pad  , \m2_data_o[28]_pad  , \m2_data_o[29]_pad  , \m2_data_o[2]_pad  , \m2_data_o[30]_pad  , \m2_data_o[31]_pad  , \m2_data_o[3]_pad  , \m2_data_o[4]_pad  , \m2_data_o[5]_pad  , \m2_data_o[6]_pad  , \m2_data_o[7]_pad  , \m2_data_o[8]_pad  , \m2_data_o[9]_pad  , \m2_err_o_pad  , \m2_rty_o_pad  , \m3_ack_o_pad  , \m3_data_o[0]_pad  , \m3_data_o[10]_pad  , \m3_data_o[11]_pad  , \m3_data_o[12]_pad  , \m3_data_o[13]_pad  , \m3_data_o[14]_pad  , \m3_data_o[15]_pad  , \m3_data_o[16]_pad  , \m3_data_o[17]_pad  , \m3_data_o[18]_pad  , \m3_data_o[19]_pad  , \m3_data_o[1]_pad  , \m3_data_o[20]_pad  , \m3_data_o[21]_pad  , \m3_data_o[22]_pad  , \m3_data_o[23]_pad  , \m3_data_o[24]_pad  , \m3_data_o[25]_pad  , \m3_data_o[26]_pad  , \m3_data_o[27]_pad  , \m3_data_o[28]_pad  , \m3_data_o[29]_pad  , \m3_data_o[2]_pad  , \m3_data_o[30]_pad  , \m3_data_o[31]_pad  , \m3_data_o[3]_pad  , \m3_data_o[4]_pad  , \m3_data_o[5]_pad  , \m3_data_o[6]_pad  , \m3_data_o[7]_pad  , \m3_data_o[8]_pad  , \m3_data_o[9]_pad  , \m3_err_o_pad  , \m3_rty_o_pad  , \m4_ack_o_pad  , \m4_data_o[0]_pad  , \m4_data_o[10]_pad  , \m4_data_o[11]_pad  , \m4_data_o[12]_pad  , \m4_data_o[13]_pad  , \m4_data_o[14]_pad  , \m4_data_o[15]_pad  , \m4_data_o[16]_pad  , \m4_data_o[17]_pad  , \m4_data_o[18]_pad  , \m4_data_o[19]_pad  , \m4_data_o[1]_pad  , \m4_data_o[20]_pad  , \m4_data_o[21]_pad  , \m4_data_o[22]_pad  , \m4_data_o[23]_pad  , \m4_data_o[24]_pad  , \m4_data_o[25]_pad  , \m4_data_o[26]_pad  , \m4_data_o[27]_pad  , \m4_data_o[28]_pad  , \m4_data_o[29]_pad  , \m4_data_o[2]_pad  , \m4_data_o[30]_pad  , \m4_data_o[31]_pad  , \m4_data_o[3]_pad  , \m4_data_o[4]_pad  , \m4_data_o[5]_pad  , \m4_data_o[6]_pad  , \m4_data_o[7]_pad  , \m4_data_o[8]_pad  , \m4_data_o[9]_pad  , \m4_err_o_pad  , \m4_rty_o_pad  , \m5_ack_o_pad  , \m5_data_o[0]_pad  , \m5_data_o[10]_pad  , \m5_data_o[11]_pad  , \m5_data_o[12]_pad  , \m5_data_o[13]_pad  , \m5_data_o[14]_pad  , \m5_data_o[15]_pad  , \m5_data_o[16]_pad  , \m5_data_o[17]_pad  , \m5_data_o[18]_pad  , \m5_data_o[19]_pad  , \m5_data_o[1]_pad  , \m5_data_o[20]_pad  , \m5_data_o[21]_pad  , \m5_data_o[22]_pad  , \m5_data_o[23]_pad  , \m5_data_o[24]_pad  , \m5_data_o[25]_pad  , \m5_data_o[26]_pad  , \m5_data_o[27]_pad  , \m5_data_o[28]_pad  , \m5_data_o[29]_pad  , \m5_data_o[2]_pad  , \m5_data_o[30]_pad  , \m5_data_o[31]_pad  , \m5_data_o[3]_pad  , \m5_data_o[4]_pad  , \m5_data_o[5]_pad  , \m5_data_o[6]_pad  , \m5_data_o[7]_pad  , \m5_data_o[8]_pad  , \m5_data_o[9]_pad  , \m5_err_o_pad  , \m5_rty_o_pad  , \m6_ack_o_pad  , \m6_data_o[0]_pad  , \m6_data_o[10]_pad  , \m6_data_o[11]_pad  , \m6_data_o[12]_pad  , \m6_data_o[13]_pad  , \m6_data_o[14]_pad  , \m6_data_o[15]_pad  , \m6_data_o[16]_pad  , \m6_data_o[17]_pad  , \m6_data_o[18]_pad  , \m6_data_o[19]_pad  , \m6_data_o[1]_pad  , \m6_data_o[20]_pad  , \m6_data_o[21]_pad  , \m6_data_o[22]_pad  , \m6_data_o[23]_pad  , \m6_data_o[24]_pad  , \m6_data_o[25]_pad  , \m6_data_o[26]_pad  , \m6_data_o[27]_pad  , \m6_data_o[28]_pad  , \m6_data_o[29]_pad  , \m6_data_o[2]_pad  , \m6_data_o[30]_pad  , \m6_data_o[31]_pad  , \m6_data_o[3]_pad  , \m6_data_o[4]_pad  , \m6_data_o[5]_pad  , \m6_data_o[6]_pad  , \m6_data_o[7]_pad  , \m6_data_o[8]_pad  , \m6_data_o[9]_pad  , \m6_err_o_pad  , \m6_rty_o_pad  , \m7_ack_o_pad  , \m7_data_o[0]_pad  , \m7_data_o[10]_pad  , \m7_data_o[11]_pad  , \m7_data_o[12]_pad  , \m7_data_o[13]_pad  , \m7_data_o[14]_pad  , \m7_data_o[15]_pad  , \m7_data_o[16]_pad  , \m7_data_o[17]_pad  , \m7_data_o[18]_pad  , \m7_data_o[19]_pad  , \m7_data_o[1]_pad  , \m7_data_o[20]_pad  , \m7_data_o[21]_pad  , \m7_data_o[22]_pad  , \m7_data_o[23]_pad  , \m7_data_o[24]_pad  , \m7_data_o[25]_pad  , \m7_data_o[26]_pad  , \m7_data_o[27]_pad  , \m7_data_o[28]_pad  , \m7_data_o[29]_pad  , \m7_data_o[2]_pad  , \m7_data_o[30]_pad  , \m7_data_o[31]_pad  , \m7_data_o[3]_pad  , \m7_data_o[4]_pad  , \m7_data_o[5]_pad  , \m7_data_o[6]_pad  , \m7_data_o[7]_pad  , \m7_data_o[8]_pad  , \m7_data_o[9]_pad  , \m7_err_o_pad  , \m7_rty_o_pad  , \s0_addr_o[0]_pad  , \s0_addr_o[10]_pad  , \s0_addr_o[11]_pad  , \s0_addr_o[12]_pad  , \s0_addr_o[13]_pad  , \s0_addr_o[14]_pad  , \s0_addr_o[15]_pad  , \s0_addr_o[16]_pad  , \s0_addr_o[17]_pad  , \s0_addr_o[18]_pad  , \s0_addr_o[19]_pad  , \s0_addr_o[1]_pad  , \s0_addr_o[20]_pad  , \s0_addr_o[21]_pad  , \s0_addr_o[22]_pad  , \s0_addr_o[23]_pad  , \s0_addr_o[24]_pad  , \s0_addr_o[25]_pad  , \s0_addr_o[26]_pad  , \s0_addr_o[27]_pad  , \s0_addr_o[28]_pad  , \s0_addr_o[29]_pad  , \s0_addr_o[2]_pad  , \s0_addr_o[30]_pad  , \s0_addr_o[31]_pad  , \s0_addr_o[3]_pad  , \s0_addr_o[4]_pad  , \s0_addr_o[5]_pad  , \s0_addr_o[6]_pad  , \s0_addr_o[7]_pad  , \s0_addr_o[8]_pad  , \s0_addr_o[9]_pad  , \s0_data_o[0]_pad  , \s0_data_o[10]_pad  , \s0_data_o[11]_pad  , \s0_data_o[12]_pad  , \s0_data_o[13]_pad  , \s0_data_o[14]_pad  , \s0_data_o[15]_pad  , \s0_data_o[16]_pad  , \s0_data_o[17]_pad  , \s0_data_o[18]_pad  , \s0_data_o[19]_pad  , \s0_data_o[1]_pad  , \s0_data_o[20]_pad  , \s0_data_o[21]_pad  , \s0_data_o[22]_pad  , \s0_data_o[23]_pad  , \s0_data_o[24]_pad  , \s0_data_o[25]_pad  , \s0_data_o[26]_pad  , \s0_data_o[27]_pad  , \s0_data_o[28]_pad  , \s0_data_o[29]_pad  , \s0_data_o[2]_pad  , \s0_data_o[30]_pad  , \s0_data_o[31]_pad  , \s0_data_o[3]_pad  , \s0_data_o[4]_pad  , \s0_data_o[5]_pad  , \s0_data_o[6]_pad  , \s0_data_o[7]_pad  , \s0_data_o[8]_pad  , \s0_data_o[9]_pad  , \s0_sel_o[0]_pad  , \s0_sel_o[1]_pad  , \s0_sel_o[2]_pad  , \s0_sel_o[3]_pad  , \s0_stb_o_pad  , \s0_we_o_pad  , \s10_addr_o[0]_pad  , \s10_addr_o[10]_pad  , \s10_addr_o[11]_pad  , \s10_addr_o[12]_pad  , \s10_addr_o[13]_pad  , \s10_addr_o[14]_pad  , \s10_addr_o[15]_pad  , \s10_addr_o[16]_pad  , \s10_addr_o[17]_pad  , \s10_addr_o[18]_pad  , \s10_addr_o[19]_pad  , \s10_addr_o[1]_pad  , \s10_addr_o[20]_pad  , \s10_addr_o[21]_pad  , \s10_addr_o[22]_pad  , \s10_addr_o[23]_pad  , \s10_addr_o[24]_pad  , \s10_addr_o[25]_pad  , \s10_addr_o[26]_pad  , \s10_addr_o[27]_pad  , \s10_addr_o[28]_pad  , \s10_addr_o[29]_pad  , \s10_addr_o[2]_pad  , \s10_addr_o[30]_pad  , \s10_addr_o[31]_pad  , \s10_addr_o[3]_pad  , \s10_addr_o[4]_pad  , \s10_addr_o[5]_pad  , \s10_addr_o[6]_pad  , \s10_addr_o[7]_pad  , \s10_addr_o[8]_pad  , \s10_addr_o[9]_pad  , \s10_data_o[0]_pad  , \s10_data_o[10]_pad  , \s10_data_o[11]_pad  , \s10_data_o[12]_pad  , \s10_data_o[13]_pad  , \s10_data_o[14]_pad  , \s10_data_o[15]_pad  , \s10_data_o[16]_pad  , \s10_data_o[17]_pad  , \s10_data_o[18]_pad  , \s10_data_o[19]_pad  , \s10_data_o[1]_pad  , \s10_data_o[20]_pad  , \s10_data_o[21]_pad  , \s10_data_o[22]_pad  , \s10_data_o[23]_pad  , \s10_data_o[24]_pad  , \s10_data_o[25]_pad  , \s10_data_o[26]_pad  , \s10_data_o[27]_pad  , \s10_data_o[28]_pad  , \s10_data_o[29]_pad  , \s10_data_o[2]_pad  , \s10_data_o[30]_pad  , \s10_data_o[31]_pad  , \s10_data_o[3]_pad  , \s10_data_o[4]_pad  , \s10_data_o[5]_pad  , \s10_data_o[6]_pad  , \s10_data_o[7]_pad  , \s10_data_o[8]_pad  , \s10_data_o[9]_pad  , \s10_sel_o[0]_pad  , \s10_sel_o[1]_pad  , \s10_sel_o[2]_pad  , \s10_sel_o[3]_pad  , \s10_stb_o_pad  , \s10_we_o_pad  , \s11_addr_o[0]_pad  , \s11_addr_o[10]_pad  , \s11_addr_o[11]_pad  , \s11_addr_o[12]_pad  , \s11_addr_o[13]_pad  , \s11_addr_o[14]_pad  , \s11_addr_o[15]_pad  , \s11_addr_o[16]_pad  , \s11_addr_o[17]_pad  , \s11_addr_o[18]_pad  , \s11_addr_o[19]_pad  , \s11_addr_o[1]_pad  , \s11_addr_o[20]_pad  , \s11_addr_o[21]_pad  , \s11_addr_o[22]_pad  , \s11_addr_o[23]_pad  , \s11_addr_o[24]_pad  , \s11_addr_o[25]_pad  , \s11_addr_o[26]_pad  , \s11_addr_o[27]_pad  , \s11_addr_o[28]_pad  , \s11_addr_o[29]_pad  , \s11_addr_o[2]_pad  , \s11_addr_o[30]_pad  , \s11_addr_o[31]_pad  , \s11_addr_o[3]_pad  , \s11_addr_o[4]_pad  , \s11_addr_o[5]_pad  , \s11_addr_o[6]_pad  , \s11_addr_o[7]_pad  , \s11_addr_o[8]_pad  , \s11_addr_o[9]_pad  , \s11_data_o[0]_pad  , \s11_data_o[10]_pad  , \s11_data_o[11]_pad  , \s11_data_o[12]_pad  , \s11_data_o[13]_pad  , \s11_data_o[14]_pad  , \s11_data_o[15]_pad  , \s11_data_o[16]_pad  , \s11_data_o[17]_pad  , \s11_data_o[18]_pad  , \s11_data_o[19]_pad  , \s11_data_o[1]_pad  , \s11_data_o[20]_pad  , \s11_data_o[21]_pad  , \s11_data_o[22]_pad  , \s11_data_o[23]_pad  , \s11_data_o[24]_pad  , \s11_data_o[25]_pad  , \s11_data_o[26]_pad  , \s11_data_o[27]_pad  , \s11_data_o[28]_pad  , \s11_data_o[29]_pad  , \s11_data_o[2]_pad  , \s11_data_o[30]_pad  , \s11_data_o[31]_pad  , \s11_data_o[3]_pad  , \s11_data_o[4]_pad  , \s11_data_o[5]_pad  , \s11_data_o[6]_pad  , \s11_data_o[7]_pad  , \s11_data_o[8]_pad  , \s11_data_o[9]_pad  , \s11_sel_o[0]_pad  , \s11_sel_o[1]_pad  , \s11_sel_o[2]_pad  , \s11_sel_o[3]_pad  , \s11_stb_o_pad  , \s11_we_o_pad  , \s12_addr_o[0]_pad  , \s12_addr_o[10]_pad  , \s12_addr_o[11]_pad  , \s12_addr_o[12]_pad  , \s12_addr_o[13]_pad  , \s12_addr_o[14]_pad  , \s12_addr_o[15]_pad  , \s12_addr_o[16]_pad  , \s12_addr_o[17]_pad  , \s12_addr_o[18]_pad  , \s12_addr_o[19]_pad  , \s12_addr_o[1]_pad  , \s12_addr_o[20]_pad  , \s12_addr_o[21]_pad  , \s12_addr_o[22]_pad  , \s12_addr_o[23]_pad  , \s12_addr_o[24]_pad  , \s12_addr_o[25]_pad  , \s12_addr_o[26]_pad  , \s12_addr_o[27]_pad  , \s12_addr_o[28]_pad  , \s12_addr_o[29]_pad  , \s12_addr_o[2]_pad  , \s12_addr_o[30]_pad  , \s12_addr_o[31]_pad  , \s12_addr_o[3]_pad  , \s12_addr_o[4]_pad  , \s12_addr_o[5]_pad  , \s12_addr_o[6]_pad  , \s12_addr_o[7]_pad  , \s12_addr_o[8]_pad  , \s12_addr_o[9]_pad  , \s12_data_o[0]_pad  , \s12_data_o[10]_pad  , \s12_data_o[11]_pad  , \s12_data_o[12]_pad  , \s12_data_o[13]_pad  , \s12_data_o[14]_pad  , \s12_data_o[15]_pad  , \s12_data_o[16]_pad  , \s12_data_o[17]_pad  , \s12_data_o[18]_pad  , \s12_data_o[19]_pad  , \s12_data_o[1]_pad  , \s12_data_o[20]_pad  , \s12_data_o[21]_pad  , \s12_data_o[22]_pad  , \s12_data_o[23]_pad  , \s12_data_o[24]_pad  , \s12_data_o[25]_pad  , \s12_data_o[26]_pad  , \s12_data_o[27]_pad  , \s12_data_o[28]_pad  , \s12_data_o[29]_pad  , \s12_data_o[2]_pad  , \s12_data_o[30]_pad  , \s12_data_o[31]_pad  , \s12_data_o[3]_pad  , \s12_data_o[4]_pad  , \s12_data_o[5]_pad  , \s12_data_o[6]_pad  , \s12_data_o[7]_pad  , \s12_data_o[8]_pad  , \s12_data_o[9]_pad  , \s12_sel_o[0]_pad  , \s12_sel_o[1]_pad  , \s12_sel_o[2]_pad  , \s12_sel_o[3]_pad  , \s12_stb_o_pad  , \s12_we_o_pad  , \s13_addr_o[0]_pad  , \s13_addr_o[10]_pad  , \s13_addr_o[11]_pad  , \s13_addr_o[12]_pad  , \s13_addr_o[13]_pad  , \s13_addr_o[14]_pad  , \s13_addr_o[15]_pad  , \s13_addr_o[16]_pad  , \s13_addr_o[17]_pad  , \s13_addr_o[18]_pad  , \s13_addr_o[19]_pad  , \s13_addr_o[1]_pad  , \s13_addr_o[20]_pad  , \s13_addr_o[21]_pad  , \s13_addr_o[22]_pad  , \s13_addr_o[23]_pad  , \s13_addr_o[24]_pad  , \s13_addr_o[25]_pad  , \s13_addr_o[26]_pad  , \s13_addr_o[27]_pad  , \s13_addr_o[28]_pad  , \s13_addr_o[29]_pad  , \s13_addr_o[2]_pad  , \s13_addr_o[30]_pad  , \s13_addr_o[31]_pad  , \s13_addr_o[3]_pad  , \s13_addr_o[4]_pad  , \s13_addr_o[5]_pad  , \s13_addr_o[6]_pad  , \s13_addr_o[7]_pad  , \s13_addr_o[8]_pad  , \s13_addr_o[9]_pad  , \s13_data_o[0]_pad  , \s13_data_o[10]_pad  , \s13_data_o[11]_pad  , \s13_data_o[12]_pad  , \s13_data_o[13]_pad  , \s13_data_o[14]_pad  , \s13_data_o[15]_pad  , \s13_data_o[16]_pad  , \s13_data_o[17]_pad  , \s13_data_o[18]_pad  , \s13_data_o[19]_pad  , \s13_data_o[1]_pad  , \s13_data_o[20]_pad  , \s13_data_o[21]_pad  , \s13_data_o[22]_pad  , \s13_data_o[23]_pad  , \s13_data_o[24]_pad  , \s13_data_o[25]_pad  , \s13_data_o[26]_pad  , \s13_data_o[27]_pad  , \s13_data_o[28]_pad  , \s13_data_o[29]_pad  , \s13_data_o[2]_pad  , \s13_data_o[30]_pad  , \s13_data_o[31]_pad  , \s13_data_o[3]_pad  , \s13_data_o[4]_pad  , \s13_data_o[5]_pad  , \s13_data_o[6]_pad  , \s13_data_o[7]_pad  , \s13_data_o[8]_pad  , \s13_data_o[9]_pad  , \s13_sel_o[0]_pad  , \s13_sel_o[1]_pad  , \s13_sel_o[2]_pad  , \s13_sel_o[3]_pad  , \s13_stb_o_pad  , \s13_we_o_pad  , \s14_addr_o[0]_pad  , \s14_addr_o[10]_pad  , \s14_addr_o[11]_pad  , \s14_addr_o[12]_pad  , \s14_addr_o[13]_pad  , \s14_addr_o[14]_pad  , \s14_addr_o[15]_pad  , \s14_addr_o[16]_pad  , \s14_addr_o[17]_pad  , \s14_addr_o[18]_pad  , \s14_addr_o[19]_pad  , \s14_addr_o[1]_pad  , \s14_addr_o[20]_pad  , \s14_addr_o[21]_pad  , \s14_addr_o[22]_pad  , \s14_addr_o[23]_pad  , \s14_addr_o[24]_pad  , \s14_addr_o[25]_pad  , \s14_addr_o[26]_pad  , \s14_addr_o[27]_pad  , \s14_addr_o[28]_pad  , \s14_addr_o[29]_pad  , \s14_addr_o[2]_pad  , \s14_addr_o[30]_pad  , \s14_addr_o[31]_pad  , \s14_addr_o[3]_pad  , \s14_addr_o[4]_pad  , \s14_addr_o[5]_pad  , \s14_addr_o[6]_pad  , \s14_addr_o[7]_pad  , \s14_addr_o[8]_pad  , \s14_addr_o[9]_pad  , \s14_data_o[0]_pad  , \s14_data_o[10]_pad  , \s14_data_o[11]_pad  , \s14_data_o[12]_pad  , \s14_data_o[13]_pad  , \s14_data_o[14]_pad  , \s14_data_o[15]_pad  , \s14_data_o[16]_pad  , \s14_data_o[17]_pad  , \s14_data_o[18]_pad  , \s14_data_o[19]_pad  , \s14_data_o[1]_pad  , \s14_data_o[20]_pad  , \s14_data_o[21]_pad  , \s14_data_o[22]_pad  , \s14_data_o[23]_pad  , \s14_data_o[24]_pad  , \s14_data_o[25]_pad  , \s14_data_o[26]_pad  , \s14_data_o[27]_pad  , \s14_data_o[28]_pad  , \s14_data_o[29]_pad  , \s14_data_o[2]_pad  , \s14_data_o[30]_pad  , \s14_data_o[31]_pad  , \s14_data_o[3]_pad  , \s14_data_o[4]_pad  , \s14_data_o[5]_pad  , \s14_data_o[6]_pad  , \s14_data_o[7]_pad  , \s14_data_o[8]_pad  , \s14_data_o[9]_pad  , \s14_sel_o[0]_pad  , \s14_sel_o[1]_pad  , \s14_sel_o[2]_pad  , \s14_sel_o[3]_pad  , \s14_stb_o_pad  , \s14_we_o_pad  , \s15_addr_o[0]_pad  , \s15_addr_o[10]_pad  , \s15_addr_o[11]_pad  , \s15_addr_o[12]_pad  , \s15_addr_o[13]_pad  , \s15_addr_o[14]_pad  , \s15_addr_o[15]_pad  , \s15_addr_o[16]_pad  , \s15_addr_o[17]_pad  , \s15_addr_o[18]_pad  , \s15_addr_o[19]_pad  , \s15_addr_o[1]_pad  , \s15_addr_o[20]_pad  , \s15_addr_o[21]_pad  , \s15_addr_o[22]_pad  , \s15_addr_o[23]_pad  , \s15_addr_o[24]_pad  , \s15_addr_o[25]_pad  , \s15_addr_o[26]_pad  , \s15_addr_o[27]_pad  , \s15_addr_o[28]_pad  , \s15_addr_o[29]_pad  , \s15_addr_o[2]_pad  , \s15_addr_o[30]_pad  , \s15_addr_o[31]_pad  , \s15_addr_o[3]_pad  , \s15_addr_o[4]_pad  , \s15_addr_o[6]_pad  , \s15_addr_o[7]_pad  , \s15_addr_o[8]_pad  , \s15_addr_o[9]_pad  , \s15_cyc_o_pad  , \s15_data_o[0]_pad  , \s15_data_o[10]_pad  , \s15_data_o[11]_pad  , \s15_data_o[12]_pad  , \s15_data_o[13]_pad  , \s15_data_o[14]_pad  , \s15_data_o[15]_pad  , \s15_data_o[16]_pad  , \s15_data_o[17]_pad  , \s15_data_o[18]_pad  , \s15_data_o[19]_pad  , \s15_data_o[1]_pad  , \s15_data_o[20]_pad  , \s15_data_o[21]_pad  , \s15_data_o[22]_pad  , \s15_data_o[23]_pad  , \s15_data_o[24]_pad  , \s15_data_o[25]_pad  , \s15_data_o[26]_pad  , \s15_data_o[27]_pad  , \s15_data_o[28]_pad  , \s15_data_o[29]_pad  , \s15_data_o[2]_pad  , \s15_data_o[30]_pad  , \s15_data_o[31]_pad  , \s15_data_o[3]_pad  , \s15_data_o[4]_pad  , \s15_data_o[5]_pad  , \s15_data_o[6]_pad  , \s15_data_o[7]_pad  , \s15_data_o[8]_pad  , \s15_data_o[9]_pad  , \s15_sel_o[0]_pad  , \s15_sel_o[1]_pad  , \s15_sel_o[2]_pad  , \s15_sel_o[3]_pad  , \s15_stb_o_pad  , \s15_we_o_pad  , \s1_addr_o[0]_pad  , \s1_addr_o[10]_pad  , \s1_addr_o[11]_pad  , \s1_addr_o[12]_pad  , \s1_addr_o[13]_pad  , \s1_addr_o[14]_pad  , \s1_addr_o[15]_pad  , \s1_addr_o[16]_pad  , \s1_addr_o[17]_pad  , \s1_addr_o[18]_pad  , \s1_addr_o[19]_pad  , \s1_addr_o[1]_pad  , \s1_addr_o[20]_pad  , \s1_addr_o[21]_pad  , \s1_addr_o[22]_pad  , \s1_addr_o[23]_pad  , \s1_addr_o[24]_pad  , \s1_addr_o[25]_pad  , \s1_addr_o[26]_pad  , \s1_addr_o[27]_pad  , \s1_addr_o[28]_pad  , \s1_addr_o[29]_pad  , \s1_addr_o[2]_pad  , \s1_addr_o[30]_pad  , \s1_addr_o[31]_pad  , \s1_addr_o[3]_pad  , \s1_addr_o[4]_pad  , \s1_addr_o[5]_pad  , \s1_addr_o[6]_pad  , \s1_addr_o[7]_pad  , \s1_addr_o[8]_pad  , \s1_addr_o[9]_pad  , \s1_data_o[0]_pad  , \s1_data_o[10]_pad  , \s1_data_o[11]_pad  , \s1_data_o[12]_pad  , \s1_data_o[13]_pad  , \s1_data_o[14]_pad  , \s1_data_o[15]_pad  , \s1_data_o[16]_pad  , \s1_data_o[17]_pad  , \s1_data_o[18]_pad  , \s1_data_o[19]_pad  , \s1_data_o[1]_pad  , \s1_data_o[20]_pad  , \s1_data_o[21]_pad  , \s1_data_o[22]_pad  , \s1_data_o[23]_pad  , \s1_data_o[24]_pad  , \s1_data_o[25]_pad  , \s1_data_o[26]_pad  , \s1_data_o[27]_pad  , \s1_data_o[28]_pad  , \s1_data_o[29]_pad  , \s1_data_o[2]_pad  , \s1_data_o[30]_pad  , \s1_data_o[31]_pad  , \s1_data_o[3]_pad  , \s1_data_o[4]_pad  , \s1_data_o[5]_pad  , \s1_data_o[6]_pad  , \s1_data_o[7]_pad  , \s1_data_o[8]_pad  , \s1_data_o[9]_pad  , \s1_sel_o[0]_pad  , \s1_sel_o[1]_pad  , \s1_sel_o[2]_pad  , \s1_sel_o[3]_pad  , \s1_stb_o_pad  , \s1_we_o_pad  , \s2_addr_o[0]_pad  , \s2_addr_o[10]_pad  , \s2_addr_o[11]_pad  , \s2_addr_o[12]_pad  , \s2_addr_o[13]_pad  , \s2_addr_o[14]_pad  , \s2_addr_o[15]_pad  , \s2_addr_o[16]_pad  , \s2_addr_o[17]_pad  , \s2_addr_o[18]_pad  , \s2_addr_o[19]_pad  , \s2_addr_o[1]_pad  , \s2_addr_o[20]_pad  , \s2_addr_o[21]_pad  , \s2_addr_o[22]_pad  , \s2_addr_o[23]_pad  , \s2_addr_o[24]_pad  , \s2_addr_o[25]_pad  , \s2_addr_o[26]_pad  , \s2_addr_o[27]_pad  , \s2_addr_o[28]_pad  , \s2_addr_o[29]_pad  , \s2_addr_o[2]_pad  , \s2_addr_o[30]_pad  , \s2_addr_o[31]_pad  , \s2_addr_o[3]_pad  , \s2_addr_o[4]_pad  , \s2_addr_o[5]_pad  , \s2_addr_o[6]_pad  , \s2_addr_o[7]_pad  , \s2_addr_o[8]_pad  , \s2_addr_o[9]_pad  , \s2_data_o[0]_pad  , \s2_data_o[10]_pad  , \s2_data_o[11]_pad  , \s2_data_o[12]_pad  , \s2_data_o[13]_pad  , \s2_data_o[14]_pad  , \s2_data_o[15]_pad  , \s2_data_o[16]_pad  , \s2_data_o[17]_pad  , \s2_data_o[18]_pad  , \s2_data_o[19]_pad  , \s2_data_o[1]_pad  , \s2_data_o[20]_pad  , \s2_data_o[21]_pad  , \s2_data_o[22]_pad  , \s2_data_o[23]_pad  , \s2_data_o[24]_pad  , \s2_data_o[25]_pad  , \s2_data_o[26]_pad  , \s2_data_o[27]_pad  , \s2_data_o[28]_pad  , \s2_data_o[29]_pad  , \s2_data_o[2]_pad  , \s2_data_o[30]_pad  , \s2_data_o[31]_pad  , \s2_data_o[3]_pad  , \s2_data_o[4]_pad  , \s2_data_o[5]_pad  , \s2_data_o[6]_pad  , \s2_data_o[7]_pad  , \s2_data_o[8]_pad  , \s2_data_o[9]_pad  , \s2_sel_o[0]_pad  , \s2_sel_o[1]_pad  , \s2_sel_o[2]_pad  , \s2_sel_o[3]_pad  , \s2_stb_o_pad  , \s2_we_o_pad  , \s3_addr_o[0]_pad  , \s3_addr_o[10]_pad  , \s3_addr_o[11]_pad  , \s3_addr_o[12]_pad  , \s3_addr_o[13]_pad  , \s3_addr_o[14]_pad  , \s3_addr_o[15]_pad  , \s3_addr_o[16]_pad  , \s3_addr_o[17]_pad  , \s3_addr_o[18]_pad  , \s3_addr_o[19]_pad  , \s3_addr_o[1]_pad  , \s3_addr_o[20]_pad  , \s3_addr_o[21]_pad  , \s3_addr_o[22]_pad  , \s3_addr_o[23]_pad  , \s3_addr_o[24]_pad  , \s3_addr_o[25]_pad  , \s3_addr_o[26]_pad  , \s3_addr_o[27]_pad  , \s3_addr_o[28]_pad  , \s3_addr_o[29]_pad  , \s3_addr_o[2]_pad  , \s3_addr_o[30]_pad  , \s3_addr_o[31]_pad  , \s3_addr_o[3]_pad  , \s3_addr_o[4]_pad  , \s3_addr_o[5]_pad  , \s3_addr_o[6]_pad  , \s3_addr_o[7]_pad  , \s3_addr_o[8]_pad  , \s3_addr_o[9]_pad  , \s3_data_o[0]_pad  , \s3_data_o[10]_pad  , \s3_data_o[11]_pad  , \s3_data_o[12]_pad  , \s3_data_o[13]_pad  , \s3_data_o[14]_pad  , \s3_data_o[15]_pad  , \s3_data_o[16]_pad  , \s3_data_o[17]_pad  , \s3_data_o[18]_pad  , \s3_data_o[19]_pad  , \s3_data_o[1]_pad  , \s3_data_o[20]_pad  , \s3_data_o[21]_pad  , \s3_data_o[22]_pad  , \s3_data_o[23]_pad  , \s3_data_o[24]_pad  , \s3_data_o[25]_pad  , \s3_data_o[26]_pad  , \s3_data_o[27]_pad  , \s3_data_o[28]_pad  , \s3_data_o[29]_pad  , \s3_data_o[2]_pad  , \s3_data_o[30]_pad  , \s3_data_o[31]_pad  , \s3_data_o[3]_pad  , \s3_data_o[4]_pad  , \s3_data_o[5]_pad  , \s3_data_o[6]_pad  , \s3_data_o[7]_pad  , \s3_data_o[8]_pad  , \s3_data_o[9]_pad  , \s3_sel_o[0]_pad  , \s3_sel_o[1]_pad  , \s3_sel_o[2]_pad  , \s3_sel_o[3]_pad  , \s3_stb_o_pad  , \s3_we_o_pad  , \s4_addr_o[0]_pad  , \s4_addr_o[10]_pad  , \s4_addr_o[11]_pad  , \s4_addr_o[12]_pad  , \s4_addr_o[13]_pad  , \s4_addr_o[14]_pad  , \s4_addr_o[15]_pad  , \s4_addr_o[16]_pad  , \s4_addr_o[17]_pad  , \s4_addr_o[18]_pad  , \s4_addr_o[19]_pad  , \s4_addr_o[1]_pad  , \s4_addr_o[20]_pad  , \s4_addr_o[21]_pad  , \s4_addr_o[22]_pad  , \s4_addr_o[23]_pad  , \s4_addr_o[24]_pad  , \s4_addr_o[25]_pad  , \s4_addr_o[26]_pad  , \s4_addr_o[27]_pad  , \s4_addr_o[28]_pad  , \s4_addr_o[29]_pad  , \s4_addr_o[2]_pad  , \s4_addr_o[30]_pad  , \s4_addr_o[31]_pad  , \s4_addr_o[3]_pad  , \s4_addr_o[4]_pad  , \s4_addr_o[5]_pad  , \s4_addr_o[6]_pad  , \s4_addr_o[7]_pad  , \s4_addr_o[8]_pad  , \s4_addr_o[9]_pad  , \s4_data_o[0]_pad  , \s4_data_o[10]_pad  , \s4_data_o[11]_pad  , \s4_data_o[12]_pad  , \s4_data_o[13]_pad  , \s4_data_o[14]_pad  , \s4_data_o[15]_pad  , \s4_data_o[16]_pad  , \s4_data_o[17]_pad  , \s4_data_o[18]_pad  , \s4_data_o[19]_pad  , \s4_data_o[1]_pad  , \s4_data_o[20]_pad  , \s4_data_o[21]_pad  , \s4_data_o[22]_pad  , \s4_data_o[23]_pad  , \s4_data_o[24]_pad  , \s4_data_o[25]_pad  , \s4_data_o[26]_pad  , \s4_data_o[27]_pad  , \s4_data_o[28]_pad  , \s4_data_o[29]_pad  , \s4_data_o[2]_pad  , \s4_data_o[30]_pad  , \s4_data_o[31]_pad  , \s4_data_o[3]_pad  , \s4_data_o[4]_pad  , \s4_data_o[5]_pad  , \s4_data_o[6]_pad  , \s4_data_o[7]_pad  , \s4_data_o[8]_pad  , \s4_data_o[9]_pad  , \s4_sel_o[0]_pad  , \s4_sel_o[1]_pad  , \s4_sel_o[2]_pad  , \s4_sel_o[3]_pad  , \s4_stb_o_pad  , \s4_we_o_pad  , \s5_addr_o[0]_pad  , \s5_addr_o[10]_pad  , \s5_addr_o[11]_pad  , \s5_addr_o[12]_pad  , \s5_addr_o[13]_pad  , \s5_addr_o[14]_pad  , \s5_addr_o[15]_pad  , \s5_addr_o[16]_pad  , \s5_addr_o[17]_pad  , \s5_addr_o[18]_pad  , \s5_addr_o[19]_pad  , \s5_addr_o[1]_pad  , \s5_addr_o[20]_pad  , \s5_addr_o[21]_pad  , \s5_addr_o[22]_pad  , \s5_addr_o[23]_pad  , \s5_addr_o[24]_pad  , \s5_addr_o[25]_pad  , \s5_addr_o[26]_pad  , \s5_addr_o[27]_pad  , \s5_addr_o[28]_pad  , \s5_addr_o[29]_pad  , \s5_addr_o[2]_pad  , \s5_addr_o[30]_pad  , \s5_addr_o[31]_pad  , \s5_addr_o[3]_pad  , \s5_addr_o[4]_pad  , \s5_addr_o[5]_pad  , \s5_addr_o[6]_pad  , \s5_addr_o[7]_pad  , \s5_addr_o[8]_pad  , \s5_addr_o[9]_pad  , \s5_data_o[0]_pad  , \s5_data_o[10]_pad  , \s5_data_o[11]_pad  , \s5_data_o[12]_pad  , \s5_data_o[13]_pad  , \s5_data_o[14]_pad  , \s5_data_o[15]_pad  , \s5_data_o[16]_pad  , \s5_data_o[17]_pad  , \s5_data_o[18]_pad  , \s5_data_o[19]_pad  , \s5_data_o[1]_pad  , \s5_data_o[20]_pad  , \s5_data_o[21]_pad  , \s5_data_o[22]_pad  , \s5_data_o[23]_pad  , \s5_data_o[24]_pad  , \s5_data_o[25]_pad  , \s5_data_o[26]_pad  , \s5_data_o[27]_pad  , \s5_data_o[28]_pad  , \s5_data_o[29]_pad  , \s5_data_o[2]_pad  , \s5_data_o[30]_pad  , \s5_data_o[31]_pad  , \s5_data_o[3]_pad  , \s5_data_o[4]_pad  , \s5_data_o[5]_pad  , \s5_data_o[6]_pad  , \s5_data_o[7]_pad  , \s5_data_o[8]_pad  , \s5_data_o[9]_pad  , \s5_sel_o[0]_pad  , \s5_sel_o[1]_pad  , \s5_sel_o[2]_pad  , \s5_sel_o[3]_pad  , \s5_stb_o_pad  , \s5_we_o_pad  , \s6_addr_o[0]_pad  , \s6_addr_o[10]_pad  , \s6_addr_o[11]_pad  , \s6_addr_o[12]_pad  , \s6_addr_o[13]_pad  , \s6_addr_o[14]_pad  , \s6_addr_o[15]_pad  , \s6_addr_o[16]_pad  , \s6_addr_o[17]_pad  , \s6_addr_o[18]_pad  , \s6_addr_o[19]_pad  , \s6_addr_o[1]_pad  , \s6_addr_o[20]_pad  , \s6_addr_o[21]_pad  , \s6_addr_o[22]_pad  , \s6_addr_o[23]_pad  , \s6_addr_o[24]_pad  , \s6_addr_o[25]_pad  , \s6_addr_o[26]_pad  , \s6_addr_o[27]_pad  , \s6_addr_o[28]_pad  , \s6_addr_o[29]_pad  , \s6_addr_o[2]_pad  , \s6_addr_o[30]_pad  , \s6_addr_o[31]_pad  , \s6_addr_o[3]_pad  , \s6_addr_o[4]_pad  , \s6_addr_o[5]_pad  , \s6_addr_o[6]_pad  , \s6_addr_o[7]_pad  , \s6_addr_o[8]_pad  , \s6_addr_o[9]_pad  , \s6_data_o[0]_pad  , \s6_data_o[10]_pad  , \s6_data_o[11]_pad  , \s6_data_o[12]_pad  , \s6_data_o[13]_pad  , \s6_data_o[14]_pad  , \s6_data_o[15]_pad  , \s6_data_o[16]_pad  , \s6_data_o[17]_pad  , \s6_data_o[18]_pad  , \s6_data_o[19]_pad  , \s6_data_o[1]_pad  , \s6_data_o[20]_pad  , \s6_data_o[21]_pad  , \s6_data_o[22]_pad  , \s6_data_o[23]_pad  , \s6_data_o[24]_pad  , \s6_data_o[25]_pad  , \s6_data_o[26]_pad  , \s6_data_o[27]_pad  , \s6_data_o[28]_pad  , \s6_data_o[29]_pad  , \s6_data_o[2]_pad  , \s6_data_o[30]_pad  , \s6_data_o[31]_pad  , \s6_data_o[3]_pad  , \s6_data_o[4]_pad  , \s6_data_o[5]_pad  , \s6_data_o[6]_pad  , \s6_data_o[7]_pad  , \s6_data_o[8]_pad  , \s6_data_o[9]_pad  , \s6_sel_o[0]_pad  , \s6_sel_o[1]_pad  , \s6_sel_o[2]_pad  , \s6_sel_o[3]_pad  , \s6_stb_o_pad  , \s6_we_o_pad  , \s7_addr_o[0]_pad  , \s7_addr_o[10]_pad  , \s7_addr_o[11]_pad  , \s7_addr_o[12]_pad  , \s7_addr_o[13]_pad  , \s7_addr_o[14]_pad  , \s7_addr_o[15]_pad  , \s7_addr_o[16]_pad  , \s7_addr_o[17]_pad  , \s7_addr_o[18]_pad  , \s7_addr_o[19]_pad  , \s7_addr_o[1]_pad  , \s7_addr_o[20]_pad  , \s7_addr_o[21]_pad  , \s7_addr_o[22]_pad  , \s7_addr_o[23]_pad  , \s7_addr_o[24]_pad  , \s7_addr_o[25]_pad  , \s7_addr_o[26]_pad  , \s7_addr_o[27]_pad  , \s7_addr_o[28]_pad  , \s7_addr_o[29]_pad  , \s7_addr_o[2]_pad  , \s7_addr_o[30]_pad  , \s7_addr_o[31]_pad  , \s7_addr_o[3]_pad  , \s7_addr_o[4]_pad  , \s7_addr_o[5]_pad  , \s7_addr_o[6]_pad  , \s7_addr_o[7]_pad  , \s7_addr_o[8]_pad  , \s7_addr_o[9]_pad  , \s7_data_o[0]_pad  , \s7_data_o[10]_pad  , \s7_data_o[11]_pad  , \s7_data_o[12]_pad  , \s7_data_o[13]_pad  , \s7_data_o[14]_pad  , \s7_data_o[15]_pad  , \s7_data_o[16]_pad  , \s7_data_o[17]_pad  , \s7_data_o[18]_pad  , \s7_data_o[19]_pad  , \s7_data_o[1]_pad  , \s7_data_o[20]_pad  , \s7_data_o[21]_pad  , \s7_data_o[22]_pad  , \s7_data_o[23]_pad  , \s7_data_o[24]_pad  , \s7_data_o[25]_pad  , \s7_data_o[26]_pad  , \s7_data_o[27]_pad  , \s7_data_o[28]_pad  , \s7_data_o[29]_pad  , \s7_data_o[2]_pad  , \s7_data_o[30]_pad  , \s7_data_o[31]_pad  , \s7_data_o[3]_pad  , \s7_data_o[4]_pad  , \s7_data_o[5]_pad  , \s7_data_o[6]_pad  , \s7_data_o[7]_pad  , \s7_data_o[8]_pad  , \s7_data_o[9]_pad  , \s7_sel_o[0]_pad  , \s7_sel_o[1]_pad  , \s7_sel_o[2]_pad  , \s7_sel_o[3]_pad  , \s7_stb_o_pad  , \s7_we_o_pad  , \s8_addr_o[0]_pad  , \s8_addr_o[10]_pad  , \s8_addr_o[11]_pad  , \s8_addr_o[12]_pad  , \s8_addr_o[13]_pad  , \s8_addr_o[14]_pad  , \s8_addr_o[15]_pad  , \s8_addr_o[16]_pad  , \s8_addr_o[17]_pad  , \s8_addr_o[18]_pad  , \s8_addr_o[19]_pad  , \s8_addr_o[1]_pad  , \s8_addr_o[20]_pad  , \s8_addr_o[21]_pad  , \s8_addr_o[22]_pad  , \s8_addr_o[23]_pad  , \s8_addr_o[24]_pad  , \s8_addr_o[25]_pad  , \s8_addr_o[26]_pad  , \s8_addr_o[27]_pad  , \s8_addr_o[28]_pad  , \s8_addr_o[29]_pad  , \s8_addr_o[2]_pad  , \s8_addr_o[30]_pad  , \s8_addr_o[31]_pad  , \s8_addr_o[3]_pad  , \s8_addr_o[4]_pad  , \s8_addr_o[5]_pad  , \s8_addr_o[6]_pad  , \s8_addr_o[7]_pad  , \s8_addr_o[8]_pad  , \s8_addr_o[9]_pad  , \s8_data_o[0]_pad  , \s8_data_o[10]_pad  , \s8_data_o[11]_pad  , \s8_data_o[12]_pad  , \s8_data_o[13]_pad  , \s8_data_o[14]_pad  , \s8_data_o[15]_pad  , \s8_data_o[16]_pad  , \s8_data_o[17]_pad  , \s8_data_o[18]_pad  , \s8_data_o[19]_pad  , \s8_data_o[1]_pad  , \s8_data_o[20]_pad  , \s8_data_o[21]_pad  , \s8_data_o[22]_pad  , \s8_data_o[23]_pad  , \s8_data_o[24]_pad  , \s8_data_o[25]_pad  , \s8_data_o[26]_pad  , \s8_data_o[27]_pad  , \s8_data_o[28]_pad  , \s8_data_o[29]_pad  , \s8_data_o[2]_pad  , \s8_data_o[30]_pad  , \s8_data_o[31]_pad  , \s8_data_o[3]_pad  , \s8_data_o[4]_pad  , \s8_data_o[5]_pad  , \s8_data_o[6]_pad  , \s8_data_o[7]_pad  , \s8_data_o[8]_pad  , \s8_data_o[9]_pad  , \s8_sel_o[0]_pad  , \s8_sel_o[1]_pad  , \s8_sel_o[2]_pad  , \s8_sel_o[3]_pad  , \s8_stb_o_pad  , \s8_we_o_pad  , \s9_addr_o[0]_pad  , \s9_addr_o[10]_pad  , \s9_addr_o[11]_pad  , \s9_addr_o[12]_pad  , \s9_addr_o[13]_pad  , \s9_addr_o[14]_pad  , \s9_addr_o[15]_pad  , \s9_addr_o[16]_pad  , \s9_addr_o[17]_pad  , \s9_addr_o[18]_pad  , \s9_addr_o[19]_pad  , \s9_addr_o[1]_pad  , \s9_addr_o[20]_pad  , \s9_addr_o[21]_pad  , \s9_addr_o[22]_pad  , \s9_addr_o[23]_pad  , \s9_addr_o[24]_pad  , \s9_addr_o[25]_pad  , \s9_addr_o[26]_pad  , \s9_addr_o[27]_pad  , \s9_addr_o[28]_pad  , \s9_addr_o[29]_pad  , \s9_addr_o[2]_pad  , \s9_addr_o[30]_pad  , \s9_addr_o[31]_pad  , \s9_addr_o[3]_pad  , \s9_addr_o[4]_pad  , \s9_addr_o[5]_pad  , \s9_addr_o[6]_pad  , \s9_addr_o[7]_pad  , \s9_addr_o[8]_pad  , \s9_addr_o[9]_pad  , \s9_data_o[0]_pad  , \s9_data_o[10]_pad  , \s9_data_o[11]_pad  , \s9_data_o[12]_pad  , \s9_data_o[13]_pad  , \s9_data_o[14]_pad  , \s9_data_o[15]_pad  , \s9_data_o[16]_pad  , \s9_data_o[17]_pad  , \s9_data_o[18]_pad  , \s9_data_o[19]_pad  , \s9_data_o[1]_pad  , \s9_data_o[20]_pad  , \s9_data_o[21]_pad  , \s9_data_o[22]_pad  , \s9_data_o[23]_pad  , \s9_data_o[24]_pad  , \s9_data_o[25]_pad  , \s9_data_o[26]_pad  , \s9_data_o[27]_pad  , \s9_data_o[28]_pad  , \s9_data_o[29]_pad  , \s9_data_o[2]_pad  , \s9_data_o[30]_pad  , \s9_data_o[31]_pad  , \s9_data_o[3]_pad  , \s9_data_o[4]_pad  , \s9_data_o[5]_pad  , \s9_data_o[6]_pad  , \s9_data_o[7]_pad  , \s9_data_o[8]_pad  , \s9_data_o[9]_pad  , \s9_sel_o[0]_pad  , \s9_sel_o[1]_pad  , \s9_sel_o[2]_pad  , \s9_sel_o[3]_pad  , \s9_stb_o_pad  , \s9_we_o_pad  );
  input \m0_addr_i[0]_pad  ;
  input \m0_addr_i[10]_pad  ;
  input \m0_addr_i[11]_pad  ;
  input \m0_addr_i[12]_pad  ;
  input \m0_addr_i[13]_pad  ;
  input \m0_addr_i[14]_pad  ;
  input \m0_addr_i[15]_pad  ;
  input \m0_addr_i[16]_pad  ;
  input \m0_addr_i[17]_pad  ;
  input \m0_addr_i[18]_pad  ;
  input \m0_addr_i[19]_pad  ;
  input \m0_addr_i[1]_pad  ;
  input \m0_addr_i[20]_pad  ;
  input \m0_addr_i[21]_pad  ;
  input \m0_addr_i[22]_pad  ;
  input \m0_addr_i[23]_pad  ;
  input \m0_addr_i[24]_pad  ;
  input \m0_addr_i[25]_pad  ;
  input \m0_addr_i[26]_pad  ;
  input \m0_addr_i[27]_pad  ;
  input \m0_addr_i[28]_pad  ;
  input \m0_addr_i[29]_pad  ;
  input \m0_addr_i[2]_pad  ;
  input \m0_addr_i[30]_pad  ;
  input \m0_addr_i[31]_pad  ;
  input \m0_addr_i[3]_pad  ;
  input \m0_addr_i[4]_pad  ;
  input \m0_addr_i[5]_pad  ;
  input \m0_addr_i[6]_pad  ;
  input \m0_addr_i[7]_pad  ;
  input \m0_addr_i[8]_pad  ;
  input \m0_addr_i[9]_pad  ;
  input \m0_cyc_i_pad  ;
  input \m0_data_i[0]_pad  ;
  input \m0_data_i[10]_pad  ;
  input \m0_data_i[11]_pad  ;
  input \m0_data_i[12]_pad  ;
  input \m0_data_i[13]_pad  ;
  input \m0_data_i[14]_pad  ;
  input \m0_data_i[15]_pad  ;
  input \m0_data_i[16]_pad  ;
  input \m0_data_i[17]_pad  ;
  input \m0_data_i[18]_pad  ;
  input \m0_data_i[19]_pad  ;
  input \m0_data_i[1]_pad  ;
  input \m0_data_i[20]_pad  ;
  input \m0_data_i[21]_pad  ;
  input \m0_data_i[22]_pad  ;
  input \m0_data_i[23]_pad  ;
  input \m0_data_i[24]_pad  ;
  input \m0_data_i[25]_pad  ;
  input \m0_data_i[26]_pad  ;
  input \m0_data_i[27]_pad  ;
  input \m0_data_i[28]_pad  ;
  input \m0_data_i[29]_pad  ;
  input \m0_data_i[2]_pad  ;
  input \m0_data_i[30]_pad  ;
  input \m0_data_i[31]_pad  ;
  input \m0_data_i[3]_pad  ;
  input \m0_data_i[4]_pad  ;
  input \m0_data_i[5]_pad  ;
  input \m0_data_i[6]_pad  ;
  input \m0_data_i[7]_pad  ;
  input \m0_data_i[8]_pad  ;
  input \m0_data_i[9]_pad  ;
  input \m0_s0_cyc_o_reg/NET0131  ;
  input \m0_s10_cyc_o_reg/NET0131  ;
  input \m0_s11_cyc_o_reg/NET0131  ;
  input \m0_s12_cyc_o_reg/NET0131  ;
  input \m0_s13_cyc_o_reg/NET0131  ;
  input \m0_s14_cyc_o_reg/NET0131  ;
  input \m0_s15_cyc_o_reg/NET0131  ;
  input \m0_s1_cyc_o_reg/NET0131  ;
  input \m0_s2_cyc_o_reg/NET0131  ;
  input \m0_s3_cyc_o_reg/NET0131  ;
  input \m0_s4_cyc_o_reg/NET0131  ;
  input \m0_s5_cyc_o_reg/NET0131  ;
  input \m0_s6_cyc_o_reg/NET0131  ;
  input \m0_s7_cyc_o_reg/NET0131  ;
  input \m0_s8_cyc_o_reg/NET0131  ;
  input \m0_s9_cyc_o_reg/NET0131  ;
  input \m0_sel_i[0]_pad  ;
  input \m0_sel_i[1]_pad  ;
  input \m0_sel_i[2]_pad  ;
  input \m0_sel_i[3]_pad  ;
  input \m0_stb_i_pad  ;
  input \m0_we_i_pad  ;
  input \m1_addr_i[0]_pad  ;
  input \m1_addr_i[10]_pad  ;
  input \m1_addr_i[11]_pad  ;
  input \m1_addr_i[12]_pad  ;
  input \m1_addr_i[13]_pad  ;
  input \m1_addr_i[14]_pad  ;
  input \m1_addr_i[15]_pad  ;
  input \m1_addr_i[16]_pad  ;
  input \m1_addr_i[17]_pad  ;
  input \m1_addr_i[18]_pad  ;
  input \m1_addr_i[19]_pad  ;
  input \m1_addr_i[1]_pad  ;
  input \m1_addr_i[20]_pad  ;
  input \m1_addr_i[21]_pad  ;
  input \m1_addr_i[22]_pad  ;
  input \m1_addr_i[23]_pad  ;
  input \m1_addr_i[24]_pad  ;
  input \m1_addr_i[25]_pad  ;
  input \m1_addr_i[26]_pad  ;
  input \m1_addr_i[27]_pad  ;
  input \m1_addr_i[28]_pad  ;
  input \m1_addr_i[29]_pad  ;
  input \m1_addr_i[2]_pad  ;
  input \m1_addr_i[30]_pad  ;
  input \m1_addr_i[31]_pad  ;
  input \m1_addr_i[3]_pad  ;
  input \m1_addr_i[4]_pad  ;
  input \m1_addr_i[5]_pad  ;
  input \m1_addr_i[6]_pad  ;
  input \m1_addr_i[7]_pad  ;
  input \m1_addr_i[8]_pad  ;
  input \m1_addr_i[9]_pad  ;
  input \m1_cyc_i_pad  ;
  input \m1_data_i[0]_pad  ;
  input \m1_data_i[10]_pad  ;
  input \m1_data_i[11]_pad  ;
  input \m1_data_i[12]_pad  ;
  input \m1_data_i[13]_pad  ;
  input \m1_data_i[14]_pad  ;
  input \m1_data_i[15]_pad  ;
  input \m1_data_i[16]_pad  ;
  input \m1_data_i[17]_pad  ;
  input \m1_data_i[18]_pad  ;
  input \m1_data_i[19]_pad  ;
  input \m1_data_i[1]_pad  ;
  input \m1_data_i[20]_pad  ;
  input \m1_data_i[21]_pad  ;
  input \m1_data_i[22]_pad  ;
  input \m1_data_i[23]_pad  ;
  input \m1_data_i[24]_pad  ;
  input \m1_data_i[25]_pad  ;
  input \m1_data_i[26]_pad  ;
  input \m1_data_i[27]_pad  ;
  input \m1_data_i[28]_pad  ;
  input \m1_data_i[29]_pad  ;
  input \m1_data_i[2]_pad  ;
  input \m1_data_i[30]_pad  ;
  input \m1_data_i[31]_pad  ;
  input \m1_data_i[3]_pad  ;
  input \m1_data_i[4]_pad  ;
  input \m1_data_i[5]_pad  ;
  input \m1_data_i[6]_pad  ;
  input \m1_data_i[7]_pad  ;
  input \m1_data_i[8]_pad  ;
  input \m1_data_i[9]_pad  ;
  input \m1_s0_cyc_o_reg/NET0131  ;
  input \m1_s10_cyc_o_reg/NET0131  ;
  input \m1_s11_cyc_o_reg/NET0131  ;
  input \m1_s12_cyc_o_reg/NET0131  ;
  input \m1_s13_cyc_o_reg/NET0131  ;
  input \m1_s14_cyc_o_reg/NET0131  ;
  input \m1_s15_cyc_o_reg/NET0131  ;
  input \m1_s1_cyc_o_reg/NET0131  ;
  input \m1_s2_cyc_o_reg/NET0131  ;
  input \m1_s3_cyc_o_reg/NET0131  ;
  input \m1_s4_cyc_o_reg/NET0131  ;
  input \m1_s5_cyc_o_reg/NET0131  ;
  input \m1_s6_cyc_o_reg/NET0131  ;
  input \m1_s7_cyc_o_reg/NET0131  ;
  input \m1_s8_cyc_o_reg/NET0131  ;
  input \m1_s9_cyc_o_reg/NET0131  ;
  input \m1_sel_i[0]_pad  ;
  input \m1_sel_i[1]_pad  ;
  input \m1_sel_i[2]_pad  ;
  input \m1_sel_i[3]_pad  ;
  input \m1_stb_i_pad  ;
  input \m1_we_i_pad  ;
  input \m2_addr_i[0]_pad  ;
  input \m2_addr_i[10]_pad  ;
  input \m2_addr_i[11]_pad  ;
  input \m2_addr_i[12]_pad  ;
  input \m2_addr_i[13]_pad  ;
  input \m2_addr_i[14]_pad  ;
  input \m2_addr_i[15]_pad  ;
  input \m2_addr_i[16]_pad  ;
  input \m2_addr_i[17]_pad  ;
  input \m2_addr_i[18]_pad  ;
  input \m2_addr_i[19]_pad  ;
  input \m2_addr_i[1]_pad  ;
  input \m2_addr_i[20]_pad  ;
  input \m2_addr_i[21]_pad  ;
  input \m2_addr_i[22]_pad  ;
  input \m2_addr_i[23]_pad  ;
  input \m2_addr_i[24]_pad  ;
  input \m2_addr_i[25]_pad  ;
  input \m2_addr_i[26]_pad  ;
  input \m2_addr_i[27]_pad  ;
  input \m2_addr_i[28]_pad  ;
  input \m2_addr_i[29]_pad  ;
  input \m2_addr_i[2]_pad  ;
  input \m2_addr_i[30]_pad  ;
  input \m2_addr_i[31]_pad  ;
  input \m2_addr_i[3]_pad  ;
  input \m2_addr_i[4]_pad  ;
  input \m2_addr_i[5]_pad  ;
  input \m2_addr_i[6]_pad  ;
  input \m2_addr_i[7]_pad  ;
  input \m2_addr_i[8]_pad  ;
  input \m2_addr_i[9]_pad  ;
  input \m2_cyc_i_pad  ;
  input \m2_data_i[0]_pad  ;
  input \m2_data_i[10]_pad  ;
  input \m2_data_i[11]_pad  ;
  input \m2_data_i[12]_pad  ;
  input \m2_data_i[13]_pad  ;
  input \m2_data_i[14]_pad  ;
  input \m2_data_i[15]_pad  ;
  input \m2_data_i[16]_pad  ;
  input \m2_data_i[17]_pad  ;
  input \m2_data_i[18]_pad  ;
  input \m2_data_i[19]_pad  ;
  input \m2_data_i[1]_pad  ;
  input \m2_data_i[20]_pad  ;
  input \m2_data_i[21]_pad  ;
  input \m2_data_i[22]_pad  ;
  input \m2_data_i[23]_pad  ;
  input \m2_data_i[24]_pad  ;
  input \m2_data_i[25]_pad  ;
  input \m2_data_i[26]_pad  ;
  input \m2_data_i[27]_pad  ;
  input \m2_data_i[28]_pad  ;
  input \m2_data_i[29]_pad  ;
  input \m2_data_i[2]_pad  ;
  input \m2_data_i[30]_pad  ;
  input \m2_data_i[31]_pad  ;
  input \m2_data_i[3]_pad  ;
  input \m2_data_i[4]_pad  ;
  input \m2_data_i[5]_pad  ;
  input \m2_data_i[6]_pad  ;
  input \m2_data_i[7]_pad  ;
  input \m2_data_i[8]_pad  ;
  input \m2_data_i[9]_pad  ;
  input \m2_s0_cyc_o_reg/NET0131  ;
  input \m2_s10_cyc_o_reg/NET0131  ;
  input \m2_s11_cyc_o_reg/NET0131  ;
  input \m2_s12_cyc_o_reg/NET0131  ;
  input \m2_s13_cyc_o_reg/NET0131  ;
  input \m2_s14_cyc_o_reg/NET0131  ;
  input \m2_s15_cyc_o_reg/NET0131  ;
  input \m2_s1_cyc_o_reg/NET0131  ;
  input \m2_s2_cyc_o_reg/NET0131  ;
  input \m2_s3_cyc_o_reg/NET0131  ;
  input \m2_s4_cyc_o_reg/NET0131  ;
  input \m2_s5_cyc_o_reg/NET0131  ;
  input \m2_s6_cyc_o_reg/NET0131  ;
  input \m2_s7_cyc_o_reg/NET0131  ;
  input \m2_s8_cyc_o_reg/NET0131  ;
  input \m2_s9_cyc_o_reg/NET0131  ;
  input \m2_sel_i[0]_pad  ;
  input \m2_sel_i[1]_pad  ;
  input \m2_sel_i[2]_pad  ;
  input \m2_sel_i[3]_pad  ;
  input \m2_stb_i_pad  ;
  input \m2_we_i_pad  ;
  input \m3_addr_i[0]_pad  ;
  input \m3_addr_i[10]_pad  ;
  input \m3_addr_i[11]_pad  ;
  input \m3_addr_i[12]_pad  ;
  input \m3_addr_i[13]_pad  ;
  input \m3_addr_i[14]_pad  ;
  input \m3_addr_i[15]_pad  ;
  input \m3_addr_i[16]_pad  ;
  input \m3_addr_i[17]_pad  ;
  input \m3_addr_i[18]_pad  ;
  input \m3_addr_i[19]_pad  ;
  input \m3_addr_i[1]_pad  ;
  input \m3_addr_i[20]_pad  ;
  input \m3_addr_i[21]_pad  ;
  input \m3_addr_i[22]_pad  ;
  input \m3_addr_i[23]_pad  ;
  input \m3_addr_i[24]_pad  ;
  input \m3_addr_i[25]_pad  ;
  input \m3_addr_i[26]_pad  ;
  input \m3_addr_i[27]_pad  ;
  input \m3_addr_i[28]_pad  ;
  input \m3_addr_i[29]_pad  ;
  input \m3_addr_i[2]_pad  ;
  input \m3_addr_i[30]_pad  ;
  input \m3_addr_i[31]_pad  ;
  input \m3_addr_i[3]_pad  ;
  input \m3_addr_i[4]_pad  ;
  input \m3_addr_i[5]_pad  ;
  input \m3_addr_i[6]_pad  ;
  input \m3_addr_i[7]_pad  ;
  input \m3_addr_i[8]_pad  ;
  input \m3_addr_i[9]_pad  ;
  input \m3_cyc_i_pad  ;
  input \m3_data_i[0]_pad  ;
  input \m3_data_i[10]_pad  ;
  input \m3_data_i[11]_pad  ;
  input \m3_data_i[12]_pad  ;
  input \m3_data_i[13]_pad  ;
  input \m3_data_i[14]_pad  ;
  input \m3_data_i[15]_pad  ;
  input \m3_data_i[16]_pad  ;
  input \m3_data_i[17]_pad  ;
  input \m3_data_i[18]_pad  ;
  input \m3_data_i[19]_pad  ;
  input \m3_data_i[1]_pad  ;
  input \m3_data_i[20]_pad  ;
  input \m3_data_i[21]_pad  ;
  input \m3_data_i[22]_pad  ;
  input \m3_data_i[23]_pad  ;
  input \m3_data_i[24]_pad  ;
  input \m3_data_i[25]_pad  ;
  input \m3_data_i[26]_pad  ;
  input \m3_data_i[27]_pad  ;
  input \m3_data_i[28]_pad  ;
  input \m3_data_i[29]_pad  ;
  input \m3_data_i[2]_pad  ;
  input \m3_data_i[30]_pad  ;
  input \m3_data_i[31]_pad  ;
  input \m3_data_i[3]_pad  ;
  input \m3_data_i[4]_pad  ;
  input \m3_data_i[5]_pad  ;
  input \m3_data_i[6]_pad  ;
  input \m3_data_i[7]_pad  ;
  input \m3_data_i[8]_pad  ;
  input \m3_data_i[9]_pad  ;
  input \m3_s0_cyc_o_reg/NET0131  ;
  input \m3_s10_cyc_o_reg/NET0131  ;
  input \m3_s11_cyc_o_reg/NET0131  ;
  input \m3_s12_cyc_o_reg/NET0131  ;
  input \m3_s13_cyc_o_reg/NET0131  ;
  input \m3_s14_cyc_o_reg/NET0131  ;
  input \m3_s15_cyc_o_reg/NET0131  ;
  input \m3_s1_cyc_o_reg/NET0131  ;
  input \m3_s2_cyc_o_reg/NET0131  ;
  input \m3_s3_cyc_o_reg/NET0131  ;
  input \m3_s4_cyc_o_reg/NET0131  ;
  input \m3_s5_cyc_o_reg/NET0131  ;
  input \m3_s6_cyc_o_reg/NET0131  ;
  input \m3_s7_cyc_o_reg/NET0131  ;
  input \m3_s8_cyc_o_reg/NET0131  ;
  input \m3_s9_cyc_o_reg/NET0131  ;
  input \m3_sel_i[0]_pad  ;
  input \m3_sel_i[1]_pad  ;
  input \m3_sel_i[2]_pad  ;
  input \m3_sel_i[3]_pad  ;
  input \m3_stb_i_pad  ;
  input \m3_we_i_pad  ;
  input \m4_addr_i[0]_pad  ;
  input \m4_addr_i[10]_pad  ;
  input \m4_addr_i[11]_pad  ;
  input \m4_addr_i[12]_pad  ;
  input \m4_addr_i[13]_pad  ;
  input \m4_addr_i[14]_pad  ;
  input \m4_addr_i[15]_pad  ;
  input \m4_addr_i[16]_pad  ;
  input \m4_addr_i[17]_pad  ;
  input \m4_addr_i[18]_pad  ;
  input \m4_addr_i[19]_pad  ;
  input \m4_addr_i[1]_pad  ;
  input \m4_addr_i[20]_pad  ;
  input \m4_addr_i[21]_pad  ;
  input \m4_addr_i[22]_pad  ;
  input \m4_addr_i[23]_pad  ;
  input \m4_addr_i[24]_pad  ;
  input \m4_addr_i[25]_pad  ;
  input \m4_addr_i[26]_pad  ;
  input \m4_addr_i[27]_pad  ;
  input \m4_addr_i[28]_pad  ;
  input \m4_addr_i[29]_pad  ;
  input \m4_addr_i[2]_pad  ;
  input \m4_addr_i[30]_pad  ;
  input \m4_addr_i[31]_pad  ;
  input \m4_addr_i[3]_pad  ;
  input \m4_addr_i[4]_pad  ;
  input \m4_addr_i[5]_pad  ;
  input \m4_addr_i[6]_pad  ;
  input \m4_addr_i[7]_pad  ;
  input \m4_addr_i[8]_pad  ;
  input \m4_addr_i[9]_pad  ;
  input \m4_cyc_i_pad  ;
  input \m4_data_i[0]_pad  ;
  input \m4_data_i[10]_pad  ;
  input \m4_data_i[11]_pad  ;
  input \m4_data_i[12]_pad  ;
  input \m4_data_i[13]_pad  ;
  input \m4_data_i[14]_pad  ;
  input \m4_data_i[15]_pad  ;
  input \m4_data_i[16]_pad  ;
  input \m4_data_i[17]_pad  ;
  input \m4_data_i[18]_pad  ;
  input \m4_data_i[19]_pad  ;
  input \m4_data_i[1]_pad  ;
  input \m4_data_i[20]_pad  ;
  input \m4_data_i[21]_pad  ;
  input \m4_data_i[22]_pad  ;
  input \m4_data_i[23]_pad  ;
  input \m4_data_i[24]_pad  ;
  input \m4_data_i[25]_pad  ;
  input \m4_data_i[26]_pad  ;
  input \m4_data_i[27]_pad  ;
  input \m4_data_i[28]_pad  ;
  input \m4_data_i[29]_pad  ;
  input \m4_data_i[2]_pad  ;
  input \m4_data_i[30]_pad  ;
  input \m4_data_i[31]_pad  ;
  input \m4_data_i[3]_pad  ;
  input \m4_data_i[4]_pad  ;
  input \m4_data_i[5]_pad  ;
  input \m4_data_i[6]_pad  ;
  input \m4_data_i[7]_pad  ;
  input \m4_data_i[8]_pad  ;
  input \m4_data_i[9]_pad  ;
  input \m4_s0_cyc_o_reg/NET0131  ;
  input \m4_s10_cyc_o_reg/NET0131  ;
  input \m4_s11_cyc_o_reg/NET0131  ;
  input \m4_s12_cyc_o_reg/NET0131  ;
  input \m4_s13_cyc_o_reg/NET0131  ;
  input \m4_s14_cyc_o_reg/NET0131  ;
  input \m4_s15_cyc_o_reg/NET0131  ;
  input \m4_s1_cyc_o_reg/NET0131  ;
  input \m4_s2_cyc_o_reg/NET0131  ;
  input \m4_s3_cyc_o_reg/NET0131  ;
  input \m4_s4_cyc_o_reg/NET0131  ;
  input \m4_s5_cyc_o_reg/NET0131  ;
  input \m4_s6_cyc_o_reg/NET0131  ;
  input \m4_s7_cyc_o_reg/NET0131  ;
  input \m4_s8_cyc_o_reg/NET0131  ;
  input \m4_s9_cyc_o_reg/NET0131  ;
  input \m4_sel_i[0]_pad  ;
  input \m4_sel_i[1]_pad  ;
  input \m4_sel_i[2]_pad  ;
  input \m4_sel_i[3]_pad  ;
  input \m4_stb_i_pad  ;
  input \m4_we_i_pad  ;
  input \m5_addr_i[0]_pad  ;
  input \m5_addr_i[10]_pad  ;
  input \m5_addr_i[11]_pad  ;
  input \m5_addr_i[12]_pad  ;
  input \m5_addr_i[13]_pad  ;
  input \m5_addr_i[14]_pad  ;
  input \m5_addr_i[15]_pad  ;
  input \m5_addr_i[16]_pad  ;
  input \m5_addr_i[17]_pad  ;
  input \m5_addr_i[18]_pad  ;
  input \m5_addr_i[19]_pad  ;
  input \m5_addr_i[1]_pad  ;
  input \m5_addr_i[20]_pad  ;
  input \m5_addr_i[21]_pad  ;
  input \m5_addr_i[22]_pad  ;
  input \m5_addr_i[23]_pad  ;
  input \m5_addr_i[24]_pad  ;
  input \m5_addr_i[25]_pad  ;
  input \m5_addr_i[26]_pad  ;
  input \m5_addr_i[27]_pad  ;
  input \m5_addr_i[28]_pad  ;
  input \m5_addr_i[29]_pad  ;
  input \m5_addr_i[2]_pad  ;
  input \m5_addr_i[30]_pad  ;
  input \m5_addr_i[31]_pad  ;
  input \m5_addr_i[3]_pad  ;
  input \m5_addr_i[4]_pad  ;
  input \m5_addr_i[5]_pad  ;
  input \m5_addr_i[6]_pad  ;
  input \m5_addr_i[7]_pad  ;
  input \m5_addr_i[8]_pad  ;
  input \m5_addr_i[9]_pad  ;
  input \m5_cyc_i_pad  ;
  input \m5_data_i[0]_pad  ;
  input \m5_data_i[10]_pad  ;
  input \m5_data_i[11]_pad  ;
  input \m5_data_i[12]_pad  ;
  input \m5_data_i[13]_pad  ;
  input \m5_data_i[14]_pad  ;
  input \m5_data_i[15]_pad  ;
  input \m5_data_i[16]_pad  ;
  input \m5_data_i[17]_pad  ;
  input \m5_data_i[18]_pad  ;
  input \m5_data_i[19]_pad  ;
  input \m5_data_i[1]_pad  ;
  input \m5_data_i[20]_pad  ;
  input \m5_data_i[21]_pad  ;
  input \m5_data_i[22]_pad  ;
  input \m5_data_i[23]_pad  ;
  input \m5_data_i[24]_pad  ;
  input \m5_data_i[25]_pad  ;
  input \m5_data_i[26]_pad  ;
  input \m5_data_i[27]_pad  ;
  input \m5_data_i[28]_pad  ;
  input \m5_data_i[29]_pad  ;
  input \m5_data_i[2]_pad  ;
  input \m5_data_i[30]_pad  ;
  input \m5_data_i[31]_pad  ;
  input \m5_data_i[3]_pad  ;
  input \m5_data_i[4]_pad  ;
  input \m5_data_i[5]_pad  ;
  input \m5_data_i[6]_pad  ;
  input \m5_data_i[7]_pad  ;
  input \m5_data_i[8]_pad  ;
  input \m5_data_i[9]_pad  ;
  input \m5_s0_cyc_o_reg/NET0131  ;
  input \m5_s10_cyc_o_reg/NET0131  ;
  input \m5_s11_cyc_o_reg/NET0131  ;
  input \m5_s12_cyc_o_reg/NET0131  ;
  input \m5_s13_cyc_o_reg/NET0131  ;
  input \m5_s14_cyc_o_reg/NET0131  ;
  input \m5_s15_cyc_o_reg/NET0131  ;
  input \m5_s1_cyc_o_reg/NET0131  ;
  input \m5_s2_cyc_o_reg/NET0131  ;
  input \m5_s3_cyc_o_reg/NET0131  ;
  input \m5_s4_cyc_o_reg/NET0131  ;
  input \m5_s5_cyc_o_reg/NET0131  ;
  input \m5_s6_cyc_o_reg/NET0131  ;
  input \m5_s7_cyc_o_reg/NET0131  ;
  input \m5_s8_cyc_o_reg/NET0131  ;
  input \m5_s9_cyc_o_reg/NET0131  ;
  input \m5_sel_i[0]_pad  ;
  input \m5_sel_i[1]_pad  ;
  input \m5_sel_i[2]_pad  ;
  input \m5_sel_i[3]_pad  ;
  input \m5_stb_i_pad  ;
  input \m5_we_i_pad  ;
  input \m6_addr_i[0]_pad  ;
  input \m6_addr_i[10]_pad  ;
  input \m6_addr_i[11]_pad  ;
  input \m6_addr_i[12]_pad  ;
  input \m6_addr_i[13]_pad  ;
  input \m6_addr_i[14]_pad  ;
  input \m6_addr_i[15]_pad  ;
  input \m6_addr_i[16]_pad  ;
  input \m6_addr_i[17]_pad  ;
  input \m6_addr_i[18]_pad  ;
  input \m6_addr_i[19]_pad  ;
  input \m6_addr_i[1]_pad  ;
  input \m6_addr_i[20]_pad  ;
  input \m6_addr_i[21]_pad  ;
  input \m6_addr_i[22]_pad  ;
  input \m6_addr_i[23]_pad  ;
  input \m6_addr_i[24]_pad  ;
  input \m6_addr_i[25]_pad  ;
  input \m6_addr_i[26]_pad  ;
  input \m6_addr_i[27]_pad  ;
  input \m6_addr_i[28]_pad  ;
  input \m6_addr_i[29]_pad  ;
  input \m6_addr_i[2]_pad  ;
  input \m6_addr_i[30]_pad  ;
  input \m6_addr_i[31]_pad  ;
  input \m6_addr_i[3]_pad  ;
  input \m6_addr_i[4]_pad  ;
  input \m6_addr_i[5]_pad  ;
  input \m6_addr_i[6]_pad  ;
  input \m6_addr_i[7]_pad  ;
  input \m6_addr_i[8]_pad  ;
  input \m6_addr_i[9]_pad  ;
  input \m6_cyc_i_pad  ;
  input \m6_data_i[0]_pad  ;
  input \m6_data_i[10]_pad  ;
  input \m6_data_i[11]_pad  ;
  input \m6_data_i[12]_pad  ;
  input \m6_data_i[13]_pad  ;
  input \m6_data_i[14]_pad  ;
  input \m6_data_i[15]_pad  ;
  input \m6_data_i[16]_pad  ;
  input \m6_data_i[17]_pad  ;
  input \m6_data_i[18]_pad  ;
  input \m6_data_i[19]_pad  ;
  input \m6_data_i[1]_pad  ;
  input \m6_data_i[20]_pad  ;
  input \m6_data_i[21]_pad  ;
  input \m6_data_i[22]_pad  ;
  input \m6_data_i[23]_pad  ;
  input \m6_data_i[24]_pad  ;
  input \m6_data_i[25]_pad  ;
  input \m6_data_i[26]_pad  ;
  input \m6_data_i[27]_pad  ;
  input \m6_data_i[28]_pad  ;
  input \m6_data_i[29]_pad  ;
  input \m6_data_i[2]_pad  ;
  input \m6_data_i[30]_pad  ;
  input \m6_data_i[31]_pad  ;
  input \m6_data_i[3]_pad  ;
  input \m6_data_i[4]_pad  ;
  input \m6_data_i[5]_pad  ;
  input \m6_data_i[6]_pad  ;
  input \m6_data_i[7]_pad  ;
  input \m6_data_i[8]_pad  ;
  input \m6_data_i[9]_pad  ;
  input \m6_s0_cyc_o_reg/NET0131  ;
  input \m6_s10_cyc_o_reg/NET0131  ;
  input \m6_s11_cyc_o_reg/NET0131  ;
  input \m6_s12_cyc_o_reg/NET0131  ;
  input \m6_s13_cyc_o_reg/NET0131  ;
  input \m6_s14_cyc_o_reg/NET0131  ;
  input \m6_s15_cyc_o_reg/NET0131  ;
  input \m6_s1_cyc_o_reg/NET0131  ;
  input \m6_s2_cyc_o_reg/NET0131  ;
  input \m6_s3_cyc_o_reg/NET0131  ;
  input \m6_s4_cyc_o_reg/NET0131  ;
  input \m6_s5_cyc_o_reg/NET0131  ;
  input \m6_s6_cyc_o_reg/NET0131  ;
  input \m6_s7_cyc_o_reg/NET0131  ;
  input \m6_s8_cyc_o_reg/NET0131  ;
  input \m6_s9_cyc_o_reg/NET0131  ;
  input \m6_sel_i[0]_pad  ;
  input \m6_sel_i[1]_pad  ;
  input \m6_sel_i[2]_pad  ;
  input \m6_sel_i[3]_pad  ;
  input \m6_stb_i_pad  ;
  input \m6_we_i_pad  ;
  input \m7_addr_i[0]_pad  ;
  input \m7_addr_i[10]_pad  ;
  input \m7_addr_i[11]_pad  ;
  input \m7_addr_i[12]_pad  ;
  input \m7_addr_i[13]_pad  ;
  input \m7_addr_i[14]_pad  ;
  input \m7_addr_i[15]_pad  ;
  input \m7_addr_i[16]_pad  ;
  input \m7_addr_i[17]_pad  ;
  input \m7_addr_i[18]_pad  ;
  input \m7_addr_i[19]_pad  ;
  input \m7_addr_i[1]_pad  ;
  input \m7_addr_i[20]_pad  ;
  input \m7_addr_i[21]_pad  ;
  input \m7_addr_i[22]_pad  ;
  input \m7_addr_i[23]_pad  ;
  input \m7_addr_i[24]_pad  ;
  input \m7_addr_i[25]_pad  ;
  input \m7_addr_i[26]_pad  ;
  input \m7_addr_i[27]_pad  ;
  input \m7_addr_i[28]_pad  ;
  input \m7_addr_i[29]_pad  ;
  input \m7_addr_i[2]_pad  ;
  input \m7_addr_i[30]_pad  ;
  input \m7_addr_i[31]_pad  ;
  input \m7_addr_i[3]_pad  ;
  input \m7_addr_i[4]_pad  ;
  input \m7_addr_i[5]_pad  ;
  input \m7_addr_i[6]_pad  ;
  input \m7_addr_i[7]_pad  ;
  input \m7_addr_i[8]_pad  ;
  input \m7_addr_i[9]_pad  ;
  input \m7_cyc_i_pad  ;
  input \m7_data_i[0]_pad  ;
  input \m7_data_i[10]_pad  ;
  input \m7_data_i[11]_pad  ;
  input \m7_data_i[12]_pad  ;
  input \m7_data_i[13]_pad  ;
  input \m7_data_i[14]_pad  ;
  input \m7_data_i[15]_pad  ;
  input \m7_data_i[16]_pad  ;
  input \m7_data_i[17]_pad  ;
  input \m7_data_i[18]_pad  ;
  input \m7_data_i[19]_pad  ;
  input \m7_data_i[1]_pad  ;
  input \m7_data_i[20]_pad  ;
  input \m7_data_i[21]_pad  ;
  input \m7_data_i[22]_pad  ;
  input \m7_data_i[23]_pad  ;
  input \m7_data_i[24]_pad  ;
  input \m7_data_i[25]_pad  ;
  input \m7_data_i[26]_pad  ;
  input \m7_data_i[27]_pad  ;
  input \m7_data_i[28]_pad  ;
  input \m7_data_i[29]_pad  ;
  input \m7_data_i[2]_pad  ;
  input \m7_data_i[30]_pad  ;
  input \m7_data_i[31]_pad  ;
  input \m7_data_i[3]_pad  ;
  input \m7_data_i[4]_pad  ;
  input \m7_data_i[5]_pad  ;
  input \m7_data_i[6]_pad  ;
  input \m7_data_i[7]_pad  ;
  input \m7_data_i[8]_pad  ;
  input \m7_data_i[9]_pad  ;
  input \m7_s0_cyc_o_reg/NET0131  ;
  input \m7_s10_cyc_o_reg/NET0131  ;
  input \m7_s11_cyc_o_reg/NET0131  ;
  input \m7_s12_cyc_o_reg/NET0131  ;
  input \m7_s13_cyc_o_reg/NET0131  ;
  input \m7_s14_cyc_o_reg/NET0131  ;
  input \m7_s15_cyc_o_reg/NET0131  ;
  input \m7_s1_cyc_o_reg/NET0131  ;
  input \m7_s2_cyc_o_reg/NET0131  ;
  input \m7_s3_cyc_o_reg/NET0131  ;
  input \m7_s4_cyc_o_reg/NET0131  ;
  input \m7_s5_cyc_o_reg/NET0131  ;
  input \m7_s6_cyc_o_reg/NET0131  ;
  input \m7_s7_cyc_o_reg/NET0131  ;
  input \m7_s8_cyc_o_reg/NET0131  ;
  input \m7_s9_cyc_o_reg/NET0131  ;
  input \m7_sel_i[0]_pad  ;
  input \m7_sel_i[1]_pad  ;
  input \m7_sel_i[2]_pad  ;
  input \m7_sel_i[3]_pad  ;
  input \m7_stb_i_pad  ;
  input \m7_we_i_pad  ;
  input \rf_conf0_reg[0]/NET0131  ;
  input \rf_conf0_reg[10]/NET0131  ;
  input \rf_conf0_reg[11]/NET0131  ;
  input \rf_conf0_reg[12]/NET0131  ;
  input \rf_conf0_reg[13]/NET0131  ;
  input \rf_conf0_reg[14]/NET0131  ;
  input \rf_conf0_reg[15]/NET0131  ;
  input \rf_conf0_reg[1]/NET0131  ;
  input \rf_conf0_reg[2]/NET0131  ;
  input \rf_conf0_reg[3]/NET0131  ;
  input \rf_conf0_reg[4]/NET0131  ;
  input \rf_conf0_reg[5]/NET0131  ;
  input \rf_conf0_reg[6]/NET0131  ;
  input \rf_conf0_reg[7]/NET0131  ;
  input \rf_conf0_reg[8]/NET0131  ;
  input \rf_conf0_reg[9]/NET0131  ;
  input \rf_conf10_reg[0]/NET0131  ;
  input \rf_conf10_reg[10]/NET0131  ;
  input \rf_conf10_reg[11]/NET0131  ;
  input \rf_conf10_reg[12]/NET0131  ;
  input \rf_conf10_reg[13]/NET0131  ;
  input \rf_conf10_reg[14]/NET0131  ;
  input \rf_conf10_reg[15]/NET0131  ;
  input \rf_conf10_reg[1]/NET0131  ;
  input \rf_conf10_reg[2]/NET0131  ;
  input \rf_conf10_reg[3]/NET0131  ;
  input \rf_conf10_reg[4]/NET0131  ;
  input \rf_conf10_reg[5]/NET0131  ;
  input \rf_conf10_reg[6]/NET0131  ;
  input \rf_conf10_reg[7]/NET0131  ;
  input \rf_conf10_reg[8]/NET0131  ;
  input \rf_conf10_reg[9]/NET0131  ;
  input \rf_conf11_reg[0]/NET0131  ;
  input \rf_conf11_reg[10]/NET0131  ;
  input \rf_conf11_reg[11]/NET0131  ;
  input \rf_conf11_reg[12]/NET0131  ;
  input \rf_conf11_reg[13]/NET0131  ;
  input \rf_conf11_reg[14]/NET0131  ;
  input \rf_conf11_reg[15]/NET0131  ;
  input \rf_conf11_reg[1]/NET0131  ;
  input \rf_conf11_reg[2]/NET0131  ;
  input \rf_conf11_reg[3]/NET0131  ;
  input \rf_conf11_reg[4]/NET0131  ;
  input \rf_conf11_reg[5]/NET0131  ;
  input \rf_conf11_reg[6]/NET0131  ;
  input \rf_conf11_reg[7]/NET0131  ;
  input \rf_conf11_reg[8]/NET0131  ;
  input \rf_conf11_reg[9]/NET0131  ;
  input \rf_conf12_reg[0]/NET0131  ;
  input \rf_conf12_reg[10]/NET0131  ;
  input \rf_conf12_reg[11]/NET0131  ;
  input \rf_conf12_reg[12]/NET0131  ;
  input \rf_conf12_reg[13]/NET0131  ;
  input \rf_conf12_reg[14]/NET0131  ;
  input \rf_conf12_reg[15]/NET0131  ;
  input \rf_conf12_reg[1]/NET0131  ;
  input \rf_conf12_reg[2]/NET0131  ;
  input \rf_conf12_reg[3]/NET0131  ;
  input \rf_conf12_reg[4]/NET0131  ;
  input \rf_conf12_reg[5]/NET0131  ;
  input \rf_conf12_reg[6]/NET0131  ;
  input \rf_conf12_reg[7]/NET0131  ;
  input \rf_conf12_reg[8]/NET0131  ;
  input \rf_conf12_reg[9]/NET0131  ;
  input \rf_conf13_reg[0]/NET0131  ;
  input \rf_conf13_reg[10]/NET0131  ;
  input \rf_conf13_reg[11]/NET0131  ;
  input \rf_conf13_reg[12]/NET0131  ;
  input \rf_conf13_reg[13]/NET0131  ;
  input \rf_conf13_reg[14]/NET0131  ;
  input \rf_conf13_reg[15]/NET0131  ;
  input \rf_conf13_reg[1]/NET0131  ;
  input \rf_conf13_reg[2]/NET0131  ;
  input \rf_conf13_reg[3]/NET0131  ;
  input \rf_conf13_reg[4]/NET0131  ;
  input \rf_conf13_reg[5]/NET0131  ;
  input \rf_conf13_reg[6]/NET0131  ;
  input \rf_conf13_reg[7]/NET0131  ;
  input \rf_conf13_reg[8]/NET0131  ;
  input \rf_conf13_reg[9]/NET0131  ;
  input \rf_conf14_reg[0]/NET0131  ;
  input \rf_conf14_reg[10]/NET0131  ;
  input \rf_conf14_reg[11]/NET0131  ;
  input \rf_conf14_reg[12]/NET0131  ;
  input \rf_conf14_reg[13]/NET0131  ;
  input \rf_conf14_reg[14]/NET0131  ;
  input \rf_conf14_reg[15]/NET0131  ;
  input \rf_conf14_reg[1]/NET0131  ;
  input \rf_conf14_reg[2]/NET0131  ;
  input \rf_conf14_reg[3]/NET0131  ;
  input \rf_conf14_reg[4]/NET0131  ;
  input \rf_conf14_reg[5]/NET0131  ;
  input \rf_conf14_reg[6]/NET0131  ;
  input \rf_conf14_reg[7]/NET0131  ;
  input \rf_conf14_reg[8]/NET0131  ;
  input \rf_conf14_reg[9]/NET0131  ;
  input \rf_conf15_reg[0]/NET0131  ;
  input \rf_conf15_reg[10]/NET0131  ;
  input \rf_conf15_reg[11]/NET0131  ;
  input \rf_conf15_reg[12]/NET0131  ;
  input \rf_conf15_reg[13]/NET0131  ;
  input \rf_conf15_reg[14]/NET0131  ;
  input \rf_conf15_reg[15]/NET0131  ;
  input \rf_conf15_reg[1]/NET0131  ;
  input \rf_conf15_reg[2]/NET0131  ;
  input \rf_conf15_reg[3]/NET0131  ;
  input \rf_conf15_reg[4]/NET0131  ;
  input \rf_conf15_reg[5]/NET0131  ;
  input \rf_conf15_reg[6]/NET0131  ;
  input \rf_conf15_reg[7]/NET0131  ;
  input \rf_conf15_reg[8]/NET0131  ;
  input \rf_conf15_reg[9]/NET0131  ;
  input \rf_conf1_reg[0]/NET0131  ;
  input \rf_conf1_reg[10]/NET0131  ;
  input \rf_conf1_reg[11]/NET0131  ;
  input \rf_conf1_reg[12]/NET0131  ;
  input \rf_conf1_reg[13]/NET0131  ;
  input \rf_conf1_reg[14]/NET0131  ;
  input \rf_conf1_reg[15]/NET0131  ;
  input \rf_conf1_reg[1]/NET0131  ;
  input \rf_conf1_reg[2]/NET0131  ;
  input \rf_conf1_reg[3]/NET0131  ;
  input \rf_conf1_reg[4]/NET0131  ;
  input \rf_conf1_reg[5]/NET0131  ;
  input \rf_conf1_reg[6]/NET0131  ;
  input \rf_conf1_reg[7]/NET0131  ;
  input \rf_conf1_reg[8]/NET0131  ;
  input \rf_conf1_reg[9]/NET0131  ;
  input \rf_conf2_reg[0]/NET0131  ;
  input \rf_conf2_reg[10]/NET0131  ;
  input \rf_conf2_reg[11]/NET0131  ;
  input \rf_conf2_reg[12]/NET0131  ;
  input \rf_conf2_reg[13]/NET0131  ;
  input \rf_conf2_reg[14]/NET0131  ;
  input \rf_conf2_reg[15]/NET0131  ;
  input \rf_conf2_reg[1]/NET0131  ;
  input \rf_conf2_reg[2]/NET0131  ;
  input \rf_conf2_reg[3]/NET0131  ;
  input \rf_conf2_reg[4]/NET0131  ;
  input \rf_conf2_reg[5]/NET0131  ;
  input \rf_conf2_reg[6]/NET0131  ;
  input \rf_conf2_reg[7]/NET0131  ;
  input \rf_conf2_reg[8]/NET0131  ;
  input \rf_conf2_reg[9]/NET0131  ;
  input \rf_conf3_reg[0]/NET0131  ;
  input \rf_conf3_reg[10]/NET0131  ;
  input \rf_conf3_reg[11]/NET0131  ;
  input \rf_conf3_reg[12]/NET0131  ;
  input \rf_conf3_reg[13]/NET0131  ;
  input \rf_conf3_reg[14]/NET0131  ;
  input \rf_conf3_reg[15]/NET0131  ;
  input \rf_conf3_reg[1]/NET0131  ;
  input \rf_conf3_reg[2]/NET0131  ;
  input \rf_conf3_reg[3]/NET0131  ;
  input \rf_conf3_reg[4]/NET0131  ;
  input \rf_conf3_reg[5]/NET0131  ;
  input \rf_conf3_reg[6]/NET0131  ;
  input \rf_conf3_reg[7]/NET0131  ;
  input \rf_conf3_reg[8]/NET0131  ;
  input \rf_conf3_reg[9]/NET0131  ;
  input \rf_conf4_reg[0]/NET0131  ;
  input \rf_conf4_reg[10]/NET0131  ;
  input \rf_conf4_reg[11]/NET0131  ;
  input \rf_conf4_reg[12]/NET0131  ;
  input \rf_conf4_reg[13]/NET0131  ;
  input \rf_conf4_reg[14]/NET0131  ;
  input \rf_conf4_reg[15]/NET0131  ;
  input \rf_conf4_reg[1]/NET0131  ;
  input \rf_conf4_reg[2]/NET0131  ;
  input \rf_conf4_reg[3]/NET0131  ;
  input \rf_conf4_reg[4]/NET0131  ;
  input \rf_conf4_reg[5]/NET0131  ;
  input \rf_conf4_reg[6]/NET0131  ;
  input \rf_conf4_reg[7]/NET0131  ;
  input \rf_conf4_reg[8]/NET0131  ;
  input \rf_conf4_reg[9]/NET0131  ;
  input \rf_conf5_reg[0]/NET0131  ;
  input \rf_conf5_reg[10]/NET0131  ;
  input \rf_conf5_reg[11]/NET0131  ;
  input \rf_conf5_reg[12]/NET0131  ;
  input \rf_conf5_reg[13]/NET0131  ;
  input \rf_conf5_reg[14]/NET0131  ;
  input \rf_conf5_reg[15]/NET0131  ;
  input \rf_conf5_reg[1]/NET0131  ;
  input \rf_conf5_reg[2]/NET0131  ;
  input \rf_conf5_reg[3]/NET0131  ;
  input \rf_conf5_reg[4]/NET0131  ;
  input \rf_conf5_reg[5]/NET0131  ;
  input \rf_conf5_reg[6]/NET0131  ;
  input \rf_conf5_reg[7]/NET0131  ;
  input \rf_conf5_reg[8]/NET0131  ;
  input \rf_conf5_reg[9]/NET0131  ;
  input \rf_conf6_reg[0]/NET0131  ;
  input \rf_conf6_reg[10]/NET0131  ;
  input \rf_conf6_reg[11]/NET0131  ;
  input \rf_conf6_reg[12]/NET0131  ;
  input \rf_conf6_reg[13]/NET0131  ;
  input \rf_conf6_reg[14]/NET0131  ;
  input \rf_conf6_reg[15]/NET0131  ;
  input \rf_conf6_reg[1]/NET0131  ;
  input \rf_conf6_reg[2]/NET0131  ;
  input \rf_conf6_reg[3]/NET0131  ;
  input \rf_conf6_reg[4]/NET0131  ;
  input \rf_conf6_reg[5]/NET0131  ;
  input \rf_conf6_reg[6]/NET0131  ;
  input \rf_conf6_reg[7]/NET0131  ;
  input \rf_conf6_reg[8]/NET0131  ;
  input \rf_conf6_reg[9]/NET0131  ;
  input \rf_conf7_reg[0]/NET0131  ;
  input \rf_conf7_reg[10]/NET0131  ;
  input \rf_conf7_reg[11]/NET0131  ;
  input \rf_conf7_reg[12]/NET0131  ;
  input \rf_conf7_reg[13]/NET0131  ;
  input \rf_conf7_reg[14]/NET0131  ;
  input \rf_conf7_reg[15]/NET0131  ;
  input \rf_conf7_reg[1]/NET0131  ;
  input \rf_conf7_reg[2]/NET0131  ;
  input \rf_conf7_reg[3]/NET0131  ;
  input \rf_conf7_reg[4]/NET0131  ;
  input \rf_conf7_reg[5]/NET0131  ;
  input \rf_conf7_reg[6]/NET0131  ;
  input \rf_conf7_reg[7]/NET0131  ;
  input \rf_conf7_reg[8]/NET0131  ;
  input \rf_conf7_reg[9]/NET0131  ;
  input \rf_conf8_reg[0]/NET0131  ;
  input \rf_conf8_reg[10]/NET0131  ;
  input \rf_conf8_reg[11]/NET0131  ;
  input \rf_conf8_reg[12]/NET0131  ;
  input \rf_conf8_reg[13]/NET0131  ;
  input \rf_conf8_reg[14]/NET0131  ;
  input \rf_conf8_reg[15]/NET0131  ;
  input \rf_conf8_reg[1]/NET0131  ;
  input \rf_conf8_reg[2]/NET0131  ;
  input \rf_conf8_reg[3]/NET0131  ;
  input \rf_conf8_reg[4]/NET0131  ;
  input \rf_conf8_reg[5]/NET0131  ;
  input \rf_conf8_reg[6]/NET0131  ;
  input \rf_conf8_reg[7]/NET0131  ;
  input \rf_conf8_reg[8]/NET0131  ;
  input \rf_conf8_reg[9]/NET0131  ;
  input \rf_conf9_reg[0]/NET0131  ;
  input \rf_conf9_reg[10]/NET0131  ;
  input \rf_conf9_reg[11]/NET0131  ;
  input \rf_conf9_reg[12]/NET0131  ;
  input \rf_conf9_reg[13]/NET0131  ;
  input \rf_conf9_reg[14]/NET0131  ;
  input \rf_conf9_reg[15]/NET0131  ;
  input \rf_conf9_reg[1]/NET0131  ;
  input \rf_conf9_reg[2]/NET0131  ;
  input \rf_conf9_reg[3]/NET0131  ;
  input \rf_conf9_reg[4]/NET0131  ;
  input \rf_conf9_reg[5]/NET0131  ;
  input \rf_conf9_reg[6]/NET0131  ;
  input \rf_conf9_reg[7]/NET0131  ;
  input \rf_conf9_reg[8]/NET0131  ;
  input \rf_conf9_reg[9]/NET0131  ;
  input \rf_rf_ack_reg/P0001  ;
  input \rf_rf_dout_reg[0]/P0001  ;
  input \rf_rf_dout_reg[10]/P0001  ;
  input \rf_rf_dout_reg[11]/P0001  ;
  input \rf_rf_dout_reg[12]/P0001  ;
  input \rf_rf_dout_reg[13]/P0001  ;
  input \rf_rf_dout_reg[14]/P0001  ;
  input \rf_rf_dout_reg[15]/P0001  ;
  input \rf_rf_dout_reg[1]/P0001  ;
  input \rf_rf_dout_reg[2]/P0001  ;
  input \rf_rf_dout_reg[3]/P0001  ;
  input \rf_rf_dout_reg[4]/P0001  ;
  input \rf_rf_dout_reg[5]/P0001  ;
  input \rf_rf_dout_reg[6]/P0001  ;
  input \rf_rf_dout_reg[7]/P0001  ;
  input \rf_rf_dout_reg[8]/P0001  ;
  input \rf_rf_dout_reg[9]/P0001  ;
  input \rf_rf_we_reg/P0001  ;
  input rst_i_pad ;
  input \s0_ack_i_pad  ;
  input \s0_data_i[0]_pad  ;
  input \s0_data_i[10]_pad  ;
  input \s0_data_i[11]_pad  ;
  input \s0_data_i[12]_pad  ;
  input \s0_data_i[13]_pad  ;
  input \s0_data_i[14]_pad  ;
  input \s0_data_i[15]_pad  ;
  input \s0_data_i[16]_pad  ;
  input \s0_data_i[17]_pad  ;
  input \s0_data_i[18]_pad  ;
  input \s0_data_i[19]_pad  ;
  input \s0_data_i[1]_pad  ;
  input \s0_data_i[20]_pad  ;
  input \s0_data_i[21]_pad  ;
  input \s0_data_i[22]_pad  ;
  input \s0_data_i[23]_pad  ;
  input \s0_data_i[24]_pad  ;
  input \s0_data_i[25]_pad  ;
  input \s0_data_i[26]_pad  ;
  input \s0_data_i[27]_pad  ;
  input \s0_data_i[28]_pad  ;
  input \s0_data_i[29]_pad  ;
  input \s0_data_i[2]_pad  ;
  input \s0_data_i[30]_pad  ;
  input \s0_data_i[31]_pad  ;
  input \s0_data_i[3]_pad  ;
  input \s0_data_i[4]_pad  ;
  input \s0_data_i[5]_pad  ;
  input \s0_data_i[6]_pad  ;
  input \s0_data_i[7]_pad  ;
  input \s0_data_i[8]_pad  ;
  input \s0_data_i[9]_pad  ;
  input \s0_err_i_pad  ;
  input \s0_m0_cyc_r_reg/P0001  ;
  input \s0_m1_cyc_r_reg/P0001  ;
  input \s0_m2_cyc_r_reg/P0001  ;
  input \s0_m3_cyc_r_reg/P0001  ;
  input \s0_m4_cyc_r_reg/P0001  ;
  input \s0_m5_cyc_r_reg/P0001  ;
  input \s0_m6_cyc_r_reg/P0001  ;
  input \s0_m7_cyc_r_reg/P0001  ;
  input \s0_msel_arb0_state_reg[0]/NET0131  ;
  input \s0_msel_arb0_state_reg[1]/NET0131  ;
  input \s0_msel_arb0_state_reg[2]/NET0131  ;
  input \s0_msel_arb1_state_reg[0]/NET0131  ;
  input \s0_msel_arb1_state_reg[1]/NET0131  ;
  input \s0_msel_arb1_state_reg[2]/NET0131  ;
  input \s0_msel_arb2_state_reg[0]/NET0131  ;
  input \s0_msel_arb2_state_reg[1]/NET0131  ;
  input \s0_msel_arb2_state_reg[2]/NET0131  ;
  input \s0_msel_arb3_state_reg[0]/NET0131  ;
  input \s0_msel_arb3_state_reg[1]/NET0131  ;
  input \s0_msel_arb3_state_reg[2]/NET0131  ;
  input \s0_msel_pri_out_reg[0]/NET0131  ;
  input \s0_msel_pri_out_reg[1]/NET0131  ;
  input \s0_next_reg/P0001  ;
  input \s0_rty_i_pad  ;
  input \s10_ack_i_pad  ;
  input \s10_data_i[0]_pad  ;
  input \s10_data_i[10]_pad  ;
  input \s10_data_i[11]_pad  ;
  input \s10_data_i[12]_pad  ;
  input \s10_data_i[13]_pad  ;
  input \s10_data_i[14]_pad  ;
  input \s10_data_i[15]_pad  ;
  input \s10_data_i[16]_pad  ;
  input \s10_data_i[17]_pad  ;
  input \s10_data_i[18]_pad  ;
  input \s10_data_i[19]_pad  ;
  input \s10_data_i[1]_pad  ;
  input \s10_data_i[20]_pad  ;
  input \s10_data_i[21]_pad  ;
  input \s10_data_i[22]_pad  ;
  input \s10_data_i[23]_pad  ;
  input \s10_data_i[24]_pad  ;
  input \s10_data_i[25]_pad  ;
  input \s10_data_i[26]_pad  ;
  input \s10_data_i[27]_pad  ;
  input \s10_data_i[28]_pad  ;
  input \s10_data_i[29]_pad  ;
  input \s10_data_i[2]_pad  ;
  input \s10_data_i[30]_pad  ;
  input \s10_data_i[31]_pad  ;
  input \s10_data_i[3]_pad  ;
  input \s10_data_i[4]_pad  ;
  input \s10_data_i[5]_pad  ;
  input \s10_data_i[6]_pad  ;
  input \s10_data_i[7]_pad  ;
  input \s10_data_i[8]_pad  ;
  input \s10_data_i[9]_pad  ;
  input \s10_err_i_pad  ;
  input \s10_m0_cyc_r_reg/P0001  ;
  input \s10_m1_cyc_r_reg/P0001  ;
  input \s10_m2_cyc_r_reg/P0001  ;
  input \s10_m3_cyc_r_reg/P0001  ;
  input \s10_m4_cyc_r_reg/P0001  ;
  input \s10_m5_cyc_r_reg/P0001  ;
  input \s10_m6_cyc_r_reg/P0001  ;
  input \s10_m7_cyc_r_reg/P0001  ;
  input \s10_msel_arb0_state_reg[0]/NET0131  ;
  input \s10_msel_arb0_state_reg[1]/NET0131  ;
  input \s10_msel_arb0_state_reg[2]/NET0131  ;
  input \s10_msel_arb1_state_reg[0]/NET0131  ;
  input \s10_msel_arb1_state_reg[1]/NET0131  ;
  input \s10_msel_arb1_state_reg[2]/NET0131  ;
  input \s10_msel_arb2_state_reg[0]/NET0131  ;
  input \s10_msel_arb2_state_reg[1]/NET0131  ;
  input \s10_msel_arb2_state_reg[2]/NET0131  ;
  input \s10_msel_arb3_state_reg[0]/NET0131  ;
  input \s10_msel_arb3_state_reg[1]/NET0131  ;
  input \s10_msel_arb3_state_reg[2]/NET0131  ;
  input \s10_msel_pri_out_reg[0]/NET0131  ;
  input \s10_msel_pri_out_reg[1]/NET0131  ;
  input \s10_next_reg/P0001  ;
  input \s10_rty_i_pad  ;
  input \s11_ack_i_pad  ;
  input \s11_data_i[0]_pad  ;
  input \s11_data_i[10]_pad  ;
  input \s11_data_i[11]_pad  ;
  input \s11_data_i[12]_pad  ;
  input \s11_data_i[13]_pad  ;
  input \s11_data_i[14]_pad  ;
  input \s11_data_i[15]_pad  ;
  input \s11_data_i[16]_pad  ;
  input \s11_data_i[17]_pad  ;
  input \s11_data_i[18]_pad  ;
  input \s11_data_i[19]_pad  ;
  input \s11_data_i[1]_pad  ;
  input \s11_data_i[20]_pad  ;
  input \s11_data_i[21]_pad  ;
  input \s11_data_i[22]_pad  ;
  input \s11_data_i[23]_pad  ;
  input \s11_data_i[24]_pad  ;
  input \s11_data_i[25]_pad  ;
  input \s11_data_i[26]_pad  ;
  input \s11_data_i[27]_pad  ;
  input \s11_data_i[28]_pad  ;
  input \s11_data_i[29]_pad  ;
  input \s11_data_i[2]_pad  ;
  input \s11_data_i[30]_pad  ;
  input \s11_data_i[31]_pad  ;
  input \s11_data_i[3]_pad  ;
  input \s11_data_i[4]_pad  ;
  input \s11_data_i[5]_pad  ;
  input \s11_data_i[6]_pad  ;
  input \s11_data_i[7]_pad  ;
  input \s11_data_i[8]_pad  ;
  input \s11_data_i[9]_pad  ;
  input \s11_err_i_pad  ;
  input \s11_m0_cyc_r_reg/P0001  ;
  input \s11_m1_cyc_r_reg/P0001  ;
  input \s11_m2_cyc_r_reg/P0001  ;
  input \s11_m3_cyc_r_reg/P0001  ;
  input \s11_m4_cyc_r_reg/P0001  ;
  input \s11_m5_cyc_r_reg/P0001  ;
  input \s11_m6_cyc_r_reg/P0001  ;
  input \s11_m7_cyc_r_reg/P0001  ;
  input \s11_msel_arb0_state_reg[0]/NET0131  ;
  input \s11_msel_arb0_state_reg[1]/NET0131  ;
  input \s11_msel_arb0_state_reg[2]/NET0131  ;
  input \s11_msel_arb1_state_reg[0]/NET0131  ;
  input \s11_msel_arb1_state_reg[1]/NET0131  ;
  input \s11_msel_arb1_state_reg[2]/NET0131  ;
  input \s11_msel_arb2_state_reg[0]/NET0131  ;
  input \s11_msel_arb2_state_reg[1]/NET0131  ;
  input \s11_msel_arb2_state_reg[2]/NET0131  ;
  input \s11_msel_arb3_state_reg[0]/NET0131  ;
  input \s11_msel_arb3_state_reg[1]/NET0131  ;
  input \s11_msel_arb3_state_reg[2]/NET0131  ;
  input \s11_msel_pri_out_reg[0]/NET0131  ;
  input \s11_msel_pri_out_reg[1]/NET0131  ;
  input \s11_next_reg/P0001  ;
  input \s11_rty_i_pad  ;
  input \s12_ack_i_pad  ;
  input \s12_data_i[0]_pad  ;
  input \s12_data_i[10]_pad  ;
  input \s12_data_i[11]_pad  ;
  input \s12_data_i[12]_pad  ;
  input \s12_data_i[13]_pad  ;
  input \s12_data_i[14]_pad  ;
  input \s12_data_i[15]_pad  ;
  input \s12_data_i[16]_pad  ;
  input \s12_data_i[17]_pad  ;
  input \s12_data_i[18]_pad  ;
  input \s12_data_i[19]_pad  ;
  input \s12_data_i[1]_pad  ;
  input \s12_data_i[20]_pad  ;
  input \s12_data_i[21]_pad  ;
  input \s12_data_i[22]_pad  ;
  input \s12_data_i[23]_pad  ;
  input \s12_data_i[24]_pad  ;
  input \s12_data_i[25]_pad  ;
  input \s12_data_i[26]_pad  ;
  input \s12_data_i[27]_pad  ;
  input \s12_data_i[28]_pad  ;
  input \s12_data_i[29]_pad  ;
  input \s12_data_i[2]_pad  ;
  input \s12_data_i[30]_pad  ;
  input \s12_data_i[31]_pad  ;
  input \s12_data_i[3]_pad  ;
  input \s12_data_i[4]_pad  ;
  input \s12_data_i[5]_pad  ;
  input \s12_data_i[6]_pad  ;
  input \s12_data_i[7]_pad  ;
  input \s12_data_i[8]_pad  ;
  input \s12_data_i[9]_pad  ;
  input \s12_err_i_pad  ;
  input \s12_m0_cyc_r_reg/P0001  ;
  input \s12_m1_cyc_r_reg/P0001  ;
  input \s12_m2_cyc_r_reg/P0001  ;
  input \s12_m3_cyc_r_reg/P0001  ;
  input \s12_m4_cyc_r_reg/P0001  ;
  input \s12_m5_cyc_r_reg/P0001  ;
  input \s12_m6_cyc_r_reg/P0001  ;
  input \s12_m7_cyc_r_reg/P0001  ;
  input \s12_msel_arb0_state_reg[0]/NET0131  ;
  input \s12_msel_arb0_state_reg[1]/NET0131  ;
  input \s12_msel_arb0_state_reg[2]/NET0131  ;
  input \s12_msel_arb1_state_reg[0]/NET0131  ;
  input \s12_msel_arb1_state_reg[1]/NET0131  ;
  input \s12_msel_arb1_state_reg[2]/NET0131  ;
  input \s12_msel_arb2_state_reg[0]/NET0131  ;
  input \s12_msel_arb2_state_reg[1]/NET0131  ;
  input \s12_msel_arb2_state_reg[2]/NET0131  ;
  input \s12_msel_arb3_state_reg[0]/NET0131  ;
  input \s12_msel_arb3_state_reg[1]/NET0131  ;
  input \s12_msel_arb3_state_reg[2]/NET0131  ;
  input \s12_msel_pri_out_reg[0]/NET0131  ;
  input \s12_msel_pri_out_reg[1]/NET0131  ;
  input \s12_next_reg/P0001  ;
  input \s12_rty_i_pad  ;
  input \s13_ack_i_pad  ;
  input \s13_data_i[0]_pad  ;
  input \s13_data_i[10]_pad  ;
  input \s13_data_i[11]_pad  ;
  input \s13_data_i[12]_pad  ;
  input \s13_data_i[13]_pad  ;
  input \s13_data_i[14]_pad  ;
  input \s13_data_i[15]_pad  ;
  input \s13_data_i[16]_pad  ;
  input \s13_data_i[17]_pad  ;
  input \s13_data_i[18]_pad  ;
  input \s13_data_i[19]_pad  ;
  input \s13_data_i[1]_pad  ;
  input \s13_data_i[20]_pad  ;
  input \s13_data_i[21]_pad  ;
  input \s13_data_i[22]_pad  ;
  input \s13_data_i[23]_pad  ;
  input \s13_data_i[24]_pad  ;
  input \s13_data_i[25]_pad  ;
  input \s13_data_i[26]_pad  ;
  input \s13_data_i[27]_pad  ;
  input \s13_data_i[28]_pad  ;
  input \s13_data_i[29]_pad  ;
  input \s13_data_i[2]_pad  ;
  input \s13_data_i[30]_pad  ;
  input \s13_data_i[31]_pad  ;
  input \s13_data_i[3]_pad  ;
  input \s13_data_i[4]_pad  ;
  input \s13_data_i[5]_pad  ;
  input \s13_data_i[6]_pad  ;
  input \s13_data_i[7]_pad  ;
  input \s13_data_i[8]_pad  ;
  input \s13_data_i[9]_pad  ;
  input \s13_err_i_pad  ;
  input \s13_m0_cyc_r_reg/P0001  ;
  input \s13_m1_cyc_r_reg/P0001  ;
  input \s13_m2_cyc_r_reg/P0001  ;
  input \s13_m3_cyc_r_reg/P0001  ;
  input \s13_m4_cyc_r_reg/P0001  ;
  input \s13_m5_cyc_r_reg/P0001  ;
  input \s13_m6_cyc_r_reg/P0001  ;
  input \s13_m7_cyc_r_reg/P0001  ;
  input \s13_msel_arb0_state_reg[0]/NET0131  ;
  input \s13_msel_arb0_state_reg[1]/NET0131  ;
  input \s13_msel_arb0_state_reg[2]/NET0131  ;
  input \s13_msel_arb1_state_reg[0]/NET0131  ;
  input \s13_msel_arb1_state_reg[1]/NET0131  ;
  input \s13_msel_arb1_state_reg[2]/NET0131  ;
  input \s13_msel_arb2_state_reg[0]/NET0131  ;
  input \s13_msel_arb2_state_reg[1]/NET0131  ;
  input \s13_msel_arb2_state_reg[2]/NET0131  ;
  input \s13_msel_arb3_state_reg[0]/NET0131  ;
  input \s13_msel_arb3_state_reg[1]/NET0131  ;
  input \s13_msel_arb3_state_reg[2]/NET0131  ;
  input \s13_msel_pri_out_reg[0]/NET0131  ;
  input \s13_msel_pri_out_reg[1]/NET0131  ;
  input \s13_next_reg/P0001  ;
  input \s13_rty_i_pad  ;
  input \s14_ack_i_pad  ;
  input \s14_data_i[0]_pad  ;
  input \s14_data_i[10]_pad  ;
  input \s14_data_i[11]_pad  ;
  input \s14_data_i[12]_pad  ;
  input \s14_data_i[13]_pad  ;
  input \s14_data_i[14]_pad  ;
  input \s14_data_i[15]_pad  ;
  input \s14_data_i[16]_pad  ;
  input \s14_data_i[17]_pad  ;
  input \s14_data_i[18]_pad  ;
  input \s14_data_i[19]_pad  ;
  input \s14_data_i[1]_pad  ;
  input \s14_data_i[20]_pad  ;
  input \s14_data_i[21]_pad  ;
  input \s14_data_i[22]_pad  ;
  input \s14_data_i[23]_pad  ;
  input \s14_data_i[24]_pad  ;
  input \s14_data_i[25]_pad  ;
  input \s14_data_i[26]_pad  ;
  input \s14_data_i[27]_pad  ;
  input \s14_data_i[28]_pad  ;
  input \s14_data_i[29]_pad  ;
  input \s14_data_i[2]_pad  ;
  input \s14_data_i[30]_pad  ;
  input \s14_data_i[31]_pad  ;
  input \s14_data_i[3]_pad  ;
  input \s14_data_i[4]_pad  ;
  input \s14_data_i[5]_pad  ;
  input \s14_data_i[6]_pad  ;
  input \s14_data_i[7]_pad  ;
  input \s14_data_i[8]_pad  ;
  input \s14_data_i[9]_pad  ;
  input \s14_err_i_pad  ;
  input \s14_m0_cyc_r_reg/P0001  ;
  input \s14_m1_cyc_r_reg/P0001  ;
  input \s14_m2_cyc_r_reg/P0001  ;
  input \s14_m3_cyc_r_reg/P0001  ;
  input \s14_m4_cyc_r_reg/P0001  ;
  input \s14_m5_cyc_r_reg/P0001  ;
  input \s14_m6_cyc_r_reg/P0001  ;
  input \s14_m7_cyc_r_reg/P0001  ;
  input \s14_msel_arb0_state_reg[0]/NET0131  ;
  input \s14_msel_arb0_state_reg[1]/NET0131  ;
  input \s14_msel_arb0_state_reg[2]/NET0131  ;
  input \s14_msel_arb1_state_reg[0]/NET0131  ;
  input \s14_msel_arb1_state_reg[1]/NET0131  ;
  input \s14_msel_arb1_state_reg[2]/NET0131  ;
  input \s14_msel_arb2_state_reg[0]/NET0131  ;
  input \s14_msel_arb2_state_reg[1]/NET0131  ;
  input \s14_msel_arb2_state_reg[2]/NET0131  ;
  input \s14_msel_arb3_state_reg[0]/NET0131  ;
  input \s14_msel_arb3_state_reg[1]/NET0131  ;
  input \s14_msel_arb3_state_reg[2]/NET0131  ;
  input \s14_msel_pri_out_reg[0]/NET0131  ;
  input \s14_msel_pri_out_reg[1]/NET0131  ;
  input \s14_next_reg/P0001  ;
  input \s14_rty_i_pad  ;
  input \s15_ack_i_pad  ;
  input \s15_data_i[0]_pad  ;
  input \s15_data_i[10]_pad  ;
  input \s15_data_i[11]_pad  ;
  input \s15_data_i[12]_pad  ;
  input \s15_data_i[13]_pad  ;
  input \s15_data_i[14]_pad  ;
  input \s15_data_i[15]_pad  ;
  input \s15_data_i[16]_pad  ;
  input \s15_data_i[17]_pad  ;
  input \s15_data_i[18]_pad  ;
  input \s15_data_i[19]_pad  ;
  input \s15_data_i[1]_pad  ;
  input \s15_data_i[20]_pad  ;
  input \s15_data_i[21]_pad  ;
  input \s15_data_i[22]_pad  ;
  input \s15_data_i[23]_pad  ;
  input \s15_data_i[24]_pad  ;
  input \s15_data_i[25]_pad  ;
  input \s15_data_i[26]_pad  ;
  input \s15_data_i[27]_pad  ;
  input \s15_data_i[28]_pad  ;
  input \s15_data_i[29]_pad  ;
  input \s15_data_i[2]_pad  ;
  input \s15_data_i[30]_pad  ;
  input \s15_data_i[31]_pad  ;
  input \s15_data_i[3]_pad  ;
  input \s15_data_i[4]_pad  ;
  input \s15_data_i[5]_pad  ;
  input \s15_data_i[6]_pad  ;
  input \s15_data_i[7]_pad  ;
  input \s15_data_i[8]_pad  ;
  input \s15_data_i[9]_pad  ;
  input \s15_err_i_pad  ;
  input \s15_m0_cyc_r_reg/P0001  ;
  input \s15_m1_cyc_r_reg/P0001  ;
  input \s15_m2_cyc_r_reg/P0001  ;
  input \s15_m3_cyc_r_reg/P0001  ;
  input \s15_m4_cyc_r_reg/P0001  ;
  input \s15_m5_cyc_r_reg/P0001  ;
  input \s15_m6_cyc_r_reg/P0001  ;
  input \s15_m7_cyc_r_reg/P0001  ;
  input \s15_msel_arb0_state_reg[0]/NET0131  ;
  input \s15_msel_arb0_state_reg[1]/NET0131  ;
  input \s15_msel_arb0_state_reg[2]/NET0131  ;
  input \s15_msel_arb1_state_reg[0]/NET0131  ;
  input \s15_msel_arb1_state_reg[1]/NET0131  ;
  input \s15_msel_arb1_state_reg[2]/NET0131  ;
  input \s15_msel_arb2_state_reg[0]/NET0131  ;
  input \s15_msel_arb2_state_reg[1]/NET0131  ;
  input \s15_msel_arb2_state_reg[2]/NET0131  ;
  input \s15_msel_arb3_state_reg[0]/NET0131  ;
  input \s15_msel_arb3_state_reg[1]/NET0131  ;
  input \s15_msel_arb3_state_reg[2]/NET0131  ;
  input \s15_msel_pri_out_reg[0]/NET0131  ;
  input \s15_msel_pri_out_reg[1]/NET0131  ;
  input \s15_next_reg/P0001  ;
  input \s15_rty_i_pad  ;
  input \s1_ack_i_pad  ;
  input \s1_data_i[0]_pad  ;
  input \s1_data_i[10]_pad  ;
  input \s1_data_i[11]_pad  ;
  input \s1_data_i[12]_pad  ;
  input \s1_data_i[13]_pad  ;
  input \s1_data_i[14]_pad  ;
  input \s1_data_i[15]_pad  ;
  input \s1_data_i[16]_pad  ;
  input \s1_data_i[17]_pad  ;
  input \s1_data_i[18]_pad  ;
  input \s1_data_i[19]_pad  ;
  input \s1_data_i[1]_pad  ;
  input \s1_data_i[20]_pad  ;
  input \s1_data_i[21]_pad  ;
  input \s1_data_i[22]_pad  ;
  input \s1_data_i[23]_pad  ;
  input \s1_data_i[24]_pad  ;
  input \s1_data_i[25]_pad  ;
  input \s1_data_i[26]_pad  ;
  input \s1_data_i[27]_pad  ;
  input \s1_data_i[28]_pad  ;
  input \s1_data_i[29]_pad  ;
  input \s1_data_i[2]_pad  ;
  input \s1_data_i[30]_pad  ;
  input \s1_data_i[31]_pad  ;
  input \s1_data_i[3]_pad  ;
  input \s1_data_i[4]_pad  ;
  input \s1_data_i[5]_pad  ;
  input \s1_data_i[6]_pad  ;
  input \s1_data_i[7]_pad  ;
  input \s1_data_i[8]_pad  ;
  input \s1_data_i[9]_pad  ;
  input \s1_err_i_pad  ;
  input \s1_m0_cyc_r_reg/P0001  ;
  input \s1_m1_cyc_r_reg/P0001  ;
  input \s1_m2_cyc_r_reg/P0001  ;
  input \s1_m3_cyc_r_reg/P0001  ;
  input \s1_m4_cyc_r_reg/P0001  ;
  input \s1_m5_cyc_r_reg/P0001  ;
  input \s1_m6_cyc_r_reg/P0001  ;
  input \s1_m7_cyc_r_reg/P0001  ;
  input \s1_msel_arb0_state_reg[0]/NET0131  ;
  input \s1_msel_arb0_state_reg[1]/NET0131  ;
  input \s1_msel_arb0_state_reg[2]/NET0131  ;
  input \s1_msel_arb1_state_reg[0]/NET0131  ;
  input \s1_msel_arb1_state_reg[1]/NET0131  ;
  input \s1_msel_arb1_state_reg[2]/NET0131  ;
  input \s1_msel_arb2_state_reg[0]/NET0131  ;
  input \s1_msel_arb2_state_reg[1]/NET0131  ;
  input \s1_msel_arb2_state_reg[2]/NET0131  ;
  input \s1_msel_arb3_state_reg[0]/NET0131  ;
  input \s1_msel_arb3_state_reg[1]/NET0131  ;
  input \s1_msel_arb3_state_reg[2]/NET0131  ;
  input \s1_msel_pri_out_reg[0]/NET0131  ;
  input \s1_msel_pri_out_reg[1]/NET0131  ;
  input \s1_next_reg/P0001  ;
  input \s1_rty_i_pad  ;
  input \s2_ack_i_pad  ;
  input \s2_data_i[0]_pad  ;
  input \s2_data_i[10]_pad  ;
  input \s2_data_i[11]_pad  ;
  input \s2_data_i[12]_pad  ;
  input \s2_data_i[13]_pad  ;
  input \s2_data_i[14]_pad  ;
  input \s2_data_i[15]_pad  ;
  input \s2_data_i[16]_pad  ;
  input \s2_data_i[17]_pad  ;
  input \s2_data_i[18]_pad  ;
  input \s2_data_i[19]_pad  ;
  input \s2_data_i[1]_pad  ;
  input \s2_data_i[20]_pad  ;
  input \s2_data_i[21]_pad  ;
  input \s2_data_i[22]_pad  ;
  input \s2_data_i[23]_pad  ;
  input \s2_data_i[24]_pad  ;
  input \s2_data_i[25]_pad  ;
  input \s2_data_i[26]_pad  ;
  input \s2_data_i[27]_pad  ;
  input \s2_data_i[28]_pad  ;
  input \s2_data_i[29]_pad  ;
  input \s2_data_i[2]_pad  ;
  input \s2_data_i[30]_pad  ;
  input \s2_data_i[31]_pad  ;
  input \s2_data_i[3]_pad  ;
  input \s2_data_i[4]_pad  ;
  input \s2_data_i[5]_pad  ;
  input \s2_data_i[6]_pad  ;
  input \s2_data_i[7]_pad  ;
  input \s2_data_i[8]_pad  ;
  input \s2_data_i[9]_pad  ;
  input \s2_err_i_pad  ;
  input \s2_m0_cyc_r_reg/P0001  ;
  input \s2_m1_cyc_r_reg/P0001  ;
  input \s2_m2_cyc_r_reg/P0001  ;
  input \s2_m3_cyc_r_reg/P0001  ;
  input \s2_m4_cyc_r_reg/P0001  ;
  input \s2_m5_cyc_r_reg/P0001  ;
  input \s2_m6_cyc_r_reg/P0001  ;
  input \s2_m7_cyc_r_reg/P0001  ;
  input \s2_msel_arb0_state_reg[0]/NET0131  ;
  input \s2_msel_arb0_state_reg[1]/NET0131  ;
  input \s2_msel_arb0_state_reg[2]/NET0131  ;
  input \s2_msel_arb1_state_reg[0]/NET0131  ;
  input \s2_msel_arb1_state_reg[1]/NET0131  ;
  input \s2_msel_arb1_state_reg[2]/NET0131  ;
  input \s2_msel_arb2_state_reg[0]/NET0131  ;
  input \s2_msel_arb2_state_reg[1]/NET0131  ;
  input \s2_msel_arb2_state_reg[2]/NET0131  ;
  input \s2_msel_arb3_state_reg[0]/NET0131  ;
  input \s2_msel_arb3_state_reg[1]/NET0131  ;
  input \s2_msel_arb3_state_reg[2]/NET0131  ;
  input \s2_msel_pri_out_reg[0]/NET0131  ;
  input \s2_msel_pri_out_reg[1]/NET0131  ;
  input \s2_next_reg/P0001  ;
  input \s2_rty_i_pad  ;
  input \s3_ack_i_pad  ;
  input \s3_data_i[0]_pad  ;
  input \s3_data_i[10]_pad  ;
  input \s3_data_i[11]_pad  ;
  input \s3_data_i[12]_pad  ;
  input \s3_data_i[13]_pad  ;
  input \s3_data_i[14]_pad  ;
  input \s3_data_i[15]_pad  ;
  input \s3_data_i[16]_pad  ;
  input \s3_data_i[17]_pad  ;
  input \s3_data_i[18]_pad  ;
  input \s3_data_i[19]_pad  ;
  input \s3_data_i[1]_pad  ;
  input \s3_data_i[20]_pad  ;
  input \s3_data_i[21]_pad  ;
  input \s3_data_i[22]_pad  ;
  input \s3_data_i[23]_pad  ;
  input \s3_data_i[24]_pad  ;
  input \s3_data_i[25]_pad  ;
  input \s3_data_i[26]_pad  ;
  input \s3_data_i[27]_pad  ;
  input \s3_data_i[28]_pad  ;
  input \s3_data_i[29]_pad  ;
  input \s3_data_i[2]_pad  ;
  input \s3_data_i[30]_pad  ;
  input \s3_data_i[31]_pad  ;
  input \s3_data_i[3]_pad  ;
  input \s3_data_i[4]_pad  ;
  input \s3_data_i[5]_pad  ;
  input \s3_data_i[6]_pad  ;
  input \s3_data_i[7]_pad  ;
  input \s3_data_i[8]_pad  ;
  input \s3_data_i[9]_pad  ;
  input \s3_err_i_pad  ;
  input \s3_m0_cyc_r_reg/P0001  ;
  input \s3_m1_cyc_r_reg/P0001  ;
  input \s3_m2_cyc_r_reg/P0001  ;
  input \s3_m3_cyc_r_reg/P0001  ;
  input \s3_m4_cyc_r_reg/P0001  ;
  input \s3_m5_cyc_r_reg/P0001  ;
  input \s3_m6_cyc_r_reg/P0001  ;
  input \s3_m7_cyc_r_reg/P0001  ;
  input \s3_msel_arb0_state_reg[0]/NET0131  ;
  input \s3_msel_arb0_state_reg[1]/NET0131  ;
  input \s3_msel_arb0_state_reg[2]/NET0131  ;
  input \s3_msel_arb1_state_reg[0]/NET0131  ;
  input \s3_msel_arb1_state_reg[1]/NET0131  ;
  input \s3_msel_arb1_state_reg[2]/NET0131  ;
  input \s3_msel_arb2_state_reg[0]/NET0131  ;
  input \s3_msel_arb2_state_reg[1]/NET0131  ;
  input \s3_msel_arb2_state_reg[2]/NET0131  ;
  input \s3_msel_arb3_state_reg[0]/NET0131  ;
  input \s3_msel_arb3_state_reg[1]/NET0131  ;
  input \s3_msel_arb3_state_reg[2]/NET0131  ;
  input \s3_msel_pri_out_reg[0]/NET0131  ;
  input \s3_msel_pri_out_reg[1]/NET0131  ;
  input \s3_next_reg/P0001  ;
  input \s3_rty_i_pad  ;
  input \s4_ack_i_pad  ;
  input \s4_data_i[0]_pad  ;
  input \s4_data_i[10]_pad  ;
  input \s4_data_i[11]_pad  ;
  input \s4_data_i[12]_pad  ;
  input \s4_data_i[13]_pad  ;
  input \s4_data_i[14]_pad  ;
  input \s4_data_i[15]_pad  ;
  input \s4_data_i[16]_pad  ;
  input \s4_data_i[17]_pad  ;
  input \s4_data_i[18]_pad  ;
  input \s4_data_i[19]_pad  ;
  input \s4_data_i[1]_pad  ;
  input \s4_data_i[20]_pad  ;
  input \s4_data_i[21]_pad  ;
  input \s4_data_i[22]_pad  ;
  input \s4_data_i[23]_pad  ;
  input \s4_data_i[24]_pad  ;
  input \s4_data_i[25]_pad  ;
  input \s4_data_i[26]_pad  ;
  input \s4_data_i[27]_pad  ;
  input \s4_data_i[28]_pad  ;
  input \s4_data_i[29]_pad  ;
  input \s4_data_i[2]_pad  ;
  input \s4_data_i[30]_pad  ;
  input \s4_data_i[31]_pad  ;
  input \s4_data_i[3]_pad  ;
  input \s4_data_i[4]_pad  ;
  input \s4_data_i[5]_pad  ;
  input \s4_data_i[6]_pad  ;
  input \s4_data_i[7]_pad  ;
  input \s4_data_i[8]_pad  ;
  input \s4_data_i[9]_pad  ;
  input \s4_err_i_pad  ;
  input \s4_m0_cyc_r_reg/P0001  ;
  input \s4_m1_cyc_r_reg/P0001  ;
  input \s4_m2_cyc_r_reg/P0001  ;
  input \s4_m3_cyc_r_reg/P0001  ;
  input \s4_m4_cyc_r_reg/P0001  ;
  input \s4_m5_cyc_r_reg/P0001  ;
  input \s4_m6_cyc_r_reg/P0001  ;
  input \s4_m7_cyc_r_reg/P0001  ;
  input \s4_msel_arb0_state_reg[0]/NET0131  ;
  input \s4_msel_arb0_state_reg[1]/NET0131  ;
  input \s4_msel_arb0_state_reg[2]/NET0131  ;
  input \s4_msel_arb1_state_reg[0]/NET0131  ;
  input \s4_msel_arb1_state_reg[1]/NET0131  ;
  input \s4_msel_arb1_state_reg[2]/NET0131  ;
  input \s4_msel_arb2_state_reg[0]/NET0131  ;
  input \s4_msel_arb2_state_reg[1]/NET0131  ;
  input \s4_msel_arb2_state_reg[2]/NET0131  ;
  input \s4_msel_arb3_state_reg[0]/NET0131  ;
  input \s4_msel_arb3_state_reg[1]/NET0131  ;
  input \s4_msel_arb3_state_reg[2]/NET0131  ;
  input \s4_msel_pri_out_reg[0]/NET0131  ;
  input \s4_msel_pri_out_reg[1]/NET0131  ;
  input \s4_next_reg/P0001  ;
  input \s4_rty_i_pad  ;
  input \s5_ack_i_pad  ;
  input \s5_data_i[0]_pad  ;
  input \s5_data_i[10]_pad  ;
  input \s5_data_i[11]_pad  ;
  input \s5_data_i[12]_pad  ;
  input \s5_data_i[13]_pad  ;
  input \s5_data_i[14]_pad  ;
  input \s5_data_i[15]_pad  ;
  input \s5_data_i[16]_pad  ;
  input \s5_data_i[17]_pad  ;
  input \s5_data_i[18]_pad  ;
  input \s5_data_i[19]_pad  ;
  input \s5_data_i[1]_pad  ;
  input \s5_data_i[20]_pad  ;
  input \s5_data_i[21]_pad  ;
  input \s5_data_i[22]_pad  ;
  input \s5_data_i[23]_pad  ;
  input \s5_data_i[24]_pad  ;
  input \s5_data_i[25]_pad  ;
  input \s5_data_i[26]_pad  ;
  input \s5_data_i[27]_pad  ;
  input \s5_data_i[28]_pad  ;
  input \s5_data_i[29]_pad  ;
  input \s5_data_i[2]_pad  ;
  input \s5_data_i[30]_pad  ;
  input \s5_data_i[31]_pad  ;
  input \s5_data_i[3]_pad  ;
  input \s5_data_i[4]_pad  ;
  input \s5_data_i[5]_pad  ;
  input \s5_data_i[6]_pad  ;
  input \s5_data_i[7]_pad  ;
  input \s5_data_i[8]_pad  ;
  input \s5_data_i[9]_pad  ;
  input \s5_err_i_pad  ;
  input \s5_m0_cyc_r_reg/P0001  ;
  input \s5_m1_cyc_r_reg/P0001  ;
  input \s5_m2_cyc_r_reg/P0001  ;
  input \s5_m3_cyc_r_reg/P0001  ;
  input \s5_m4_cyc_r_reg/P0001  ;
  input \s5_m5_cyc_r_reg/P0001  ;
  input \s5_m6_cyc_r_reg/P0001  ;
  input \s5_m7_cyc_r_reg/P0001  ;
  input \s5_msel_arb0_state_reg[0]/NET0131  ;
  input \s5_msel_arb0_state_reg[1]/NET0131  ;
  input \s5_msel_arb0_state_reg[2]/NET0131  ;
  input \s5_msel_arb1_state_reg[0]/NET0131  ;
  input \s5_msel_arb1_state_reg[1]/NET0131  ;
  input \s5_msel_arb1_state_reg[2]/NET0131  ;
  input \s5_msel_arb2_state_reg[0]/NET0131  ;
  input \s5_msel_arb2_state_reg[1]/NET0131  ;
  input \s5_msel_arb2_state_reg[2]/NET0131  ;
  input \s5_msel_arb3_state_reg[0]/NET0131  ;
  input \s5_msel_arb3_state_reg[1]/NET0131  ;
  input \s5_msel_arb3_state_reg[2]/NET0131  ;
  input \s5_msel_pri_out_reg[0]/NET0131  ;
  input \s5_msel_pri_out_reg[1]/NET0131  ;
  input \s5_next_reg/P0001  ;
  input \s5_rty_i_pad  ;
  input \s6_ack_i_pad  ;
  input \s6_data_i[0]_pad  ;
  input \s6_data_i[10]_pad  ;
  input \s6_data_i[11]_pad  ;
  input \s6_data_i[12]_pad  ;
  input \s6_data_i[13]_pad  ;
  input \s6_data_i[14]_pad  ;
  input \s6_data_i[15]_pad  ;
  input \s6_data_i[16]_pad  ;
  input \s6_data_i[17]_pad  ;
  input \s6_data_i[18]_pad  ;
  input \s6_data_i[19]_pad  ;
  input \s6_data_i[1]_pad  ;
  input \s6_data_i[20]_pad  ;
  input \s6_data_i[21]_pad  ;
  input \s6_data_i[22]_pad  ;
  input \s6_data_i[23]_pad  ;
  input \s6_data_i[24]_pad  ;
  input \s6_data_i[25]_pad  ;
  input \s6_data_i[26]_pad  ;
  input \s6_data_i[27]_pad  ;
  input \s6_data_i[28]_pad  ;
  input \s6_data_i[29]_pad  ;
  input \s6_data_i[2]_pad  ;
  input \s6_data_i[30]_pad  ;
  input \s6_data_i[31]_pad  ;
  input \s6_data_i[3]_pad  ;
  input \s6_data_i[4]_pad  ;
  input \s6_data_i[5]_pad  ;
  input \s6_data_i[6]_pad  ;
  input \s6_data_i[7]_pad  ;
  input \s6_data_i[8]_pad  ;
  input \s6_data_i[9]_pad  ;
  input \s6_err_i_pad  ;
  input \s6_m0_cyc_r_reg/P0001  ;
  input \s6_m1_cyc_r_reg/P0001  ;
  input \s6_m2_cyc_r_reg/P0001  ;
  input \s6_m3_cyc_r_reg/P0001  ;
  input \s6_m4_cyc_r_reg/P0001  ;
  input \s6_m5_cyc_r_reg/P0001  ;
  input \s6_m6_cyc_r_reg/P0001  ;
  input \s6_m7_cyc_r_reg/P0001  ;
  input \s6_msel_arb0_state_reg[0]/NET0131  ;
  input \s6_msel_arb0_state_reg[1]/NET0131  ;
  input \s6_msel_arb0_state_reg[2]/NET0131  ;
  input \s6_msel_arb1_state_reg[0]/NET0131  ;
  input \s6_msel_arb1_state_reg[1]/NET0131  ;
  input \s6_msel_arb1_state_reg[2]/NET0131  ;
  input \s6_msel_arb2_state_reg[0]/NET0131  ;
  input \s6_msel_arb2_state_reg[1]/NET0131  ;
  input \s6_msel_arb2_state_reg[2]/NET0131  ;
  input \s6_msel_arb3_state_reg[0]/NET0131  ;
  input \s6_msel_arb3_state_reg[1]/NET0131  ;
  input \s6_msel_arb3_state_reg[2]/NET0131  ;
  input \s6_msel_pri_out_reg[0]/NET0131  ;
  input \s6_msel_pri_out_reg[1]/NET0131  ;
  input \s6_next_reg/P0001  ;
  input \s6_rty_i_pad  ;
  input \s7_ack_i_pad  ;
  input \s7_data_i[0]_pad  ;
  input \s7_data_i[10]_pad  ;
  input \s7_data_i[11]_pad  ;
  input \s7_data_i[12]_pad  ;
  input \s7_data_i[13]_pad  ;
  input \s7_data_i[14]_pad  ;
  input \s7_data_i[15]_pad  ;
  input \s7_data_i[16]_pad  ;
  input \s7_data_i[17]_pad  ;
  input \s7_data_i[18]_pad  ;
  input \s7_data_i[19]_pad  ;
  input \s7_data_i[1]_pad  ;
  input \s7_data_i[20]_pad  ;
  input \s7_data_i[21]_pad  ;
  input \s7_data_i[22]_pad  ;
  input \s7_data_i[23]_pad  ;
  input \s7_data_i[24]_pad  ;
  input \s7_data_i[25]_pad  ;
  input \s7_data_i[26]_pad  ;
  input \s7_data_i[27]_pad  ;
  input \s7_data_i[28]_pad  ;
  input \s7_data_i[29]_pad  ;
  input \s7_data_i[2]_pad  ;
  input \s7_data_i[30]_pad  ;
  input \s7_data_i[31]_pad  ;
  input \s7_data_i[3]_pad  ;
  input \s7_data_i[4]_pad  ;
  input \s7_data_i[5]_pad  ;
  input \s7_data_i[6]_pad  ;
  input \s7_data_i[7]_pad  ;
  input \s7_data_i[8]_pad  ;
  input \s7_data_i[9]_pad  ;
  input \s7_err_i_pad  ;
  input \s7_m0_cyc_r_reg/P0001  ;
  input \s7_m1_cyc_r_reg/P0001  ;
  input \s7_m2_cyc_r_reg/P0001  ;
  input \s7_m3_cyc_r_reg/P0001  ;
  input \s7_m4_cyc_r_reg/P0001  ;
  input \s7_m5_cyc_r_reg/P0001  ;
  input \s7_m6_cyc_r_reg/P0001  ;
  input \s7_m7_cyc_r_reg/P0001  ;
  input \s7_msel_arb0_state_reg[0]/NET0131  ;
  input \s7_msel_arb0_state_reg[1]/NET0131  ;
  input \s7_msel_arb0_state_reg[2]/NET0131  ;
  input \s7_msel_arb1_state_reg[0]/NET0131  ;
  input \s7_msel_arb1_state_reg[1]/NET0131  ;
  input \s7_msel_arb1_state_reg[2]/NET0131  ;
  input \s7_msel_arb2_state_reg[0]/NET0131  ;
  input \s7_msel_arb2_state_reg[1]/NET0131  ;
  input \s7_msel_arb2_state_reg[2]/NET0131  ;
  input \s7_msel_arb3_state_reg[0]/NET0131  ;
  input \s7_msel_arb3_state_reg[1]/NET0131  ;
  input \s7_msel_arb3_state_reg[2]/NET0131  ;
  input \s7_msel_pri_out_reg[0]/NET0131  ;
  input \s7_msel_pri_out_reg[1]/NET0131  ;
  input \s7_next_reg/P0001  ;
  input \s7_rty_i_pad  ;
  input \s8_ack_i_pad  ;
  input \s8_data_i[0]_pad  ;
  input \s8_data_i[10]_pad  ;
  input \s8_data_i[11]_pad  ;
  input \s8_data_i[12]_pad  ;
  input \s8_data_i[13]_pad  ;
  input \s8_data_i[14]_pad  ;
  input \s8_data_i[15]_pad  ;
  input \s8_data_i[16]_pad  ;
  input \s8_data_i[17]_pad  ;
  input \s8_data_i[18]_pad  ;
  input \s8_data_i[19]_pad  ;
  input \s8_data_i[1]_pad  ;
  input \s8_data_i[20]_pad  ;
  input \s8_data_i[21]_pad  ;
  input \s8_data_i[22]_pad  ;
  input \s8_data_i[23]_pad  ;
  input \s8_data_i[24]_pad  ;
  input \s8_data_i[25]_pad  ;
  input \s8_data_i[26]_pad  ;
  input \s8_data_i[27]_pad  ;
  input \s8_data_i[28]_pad  ;
  input \s8_data_i[29]_pad  ;
  input \s8_data_i[2]_pad  ;
  input \s8_data_i[30]_pad  ;
  input \s8_data_i[31]_pad  ;
  input \s8_data_i[3]_pad  ;
  input \s8_data_i[4]_pad  ;
  input \s8_data_i[5]_pad  ;
  input \s8_data_i[6]_pad  ;
  input \s8_data_i[7]_pad  ;
  input \s8_data_i[8]_pad  ;
  input \s8_data_i[9]_pad  ;
  input \s8_err_i_pad  ;
  input \s8_m0_cyc_r_reg/P0001  ;
  input \s8_m1_cyc_r_reg/P0001  ;
  input \s8_m2_cyc_r_reg/P0001  ;
  input \s8_m3_cyc_r_reg/P0001  ;
  input \s8_m4_cyc_r_reg/P0001  ;
  input \s8_m5_cyc_r_reg/P0001  ;
  input \s8_m6_cyc_r_reg/P0001  ;
  input \s8_m7_cyc_r_reg/P0001  ;
  input \s8_msel_arb0_state_reg[0]/NET0131  ;
  input \s8_msel_arb0_state_reg[1]/NET0131  ;
  input \s8_msel_arb0_state_reg[2]/NET0131  ;
  input \s8_msel_arb1_state_reg[0]/NET0131  ;
  input \s8_msel_arb1_state_reg[1]/NET0131  ;
  input \s8_msel_arb1_state_reg[2]/NET0131  ;
  input \s8_msel_arb2_state_reg[0]/NET0131  ;
  input \s8_msel_arb2_state_reg[1]/NET0131  ;
  input \s8_msel_arb2_state_reg[2]/NET0131  ;
  input \s8_msel_arb3_state_reg[0]/NET0131  ;
  input \s8_msel_arb3_state_reg[1]/NET0131  ;
  input \s8_msel_arb3_state_reg[2]/NET0131  ;
  input \s8_msel_pri_out_reg[0]/NET0131  ;
  input \s8_msel_pri_out_reg[1]/NET0131  ;
  input \s8_next_reg/P0001  ;
  input \s8_rty_i_pad  ;
  input \s9_ack_i_pad  ;
  input \s9_data_i[0]_pad  ;
  input \s9_data_i[10]_pad  ;
  input \s9_data_i[11]_pad  ;
  input \s9_data_i[12]_pad  ;
  input \s9_data_i[13]_pad  ;
  input \s9_data_i[14]_pad  ;
  input \s9_data_i[15]_pad  ;
  input \s9_data_i[16]_pad  ;
  input \s9_data_i[17]_pad  ;
  input \s9_data_i[18]_pad  ;
  input \s9_data_i[19]_pad  ;
  input \s9_data_i[1]_pad  ;
  input \s9_data_i[20]_pad  ;
  input \s9_data_i[21]_pad  ;
  input \s9_data_i[22]_pad  ;
  input \s9_data_i[23]_pad  ;
  input \s9_data_i[24]_pad  ;
  input \s9_data_i[25]_pad  ;
  input \s9_data_i[26]_pad  ;
  input \s9_data_i[27]_pad  ;
  input \s9_data_i[28]_pad  ;
  input \s9_data_i[29]_pad  ;
  input \s9_data_i[2]_pad  ;
  input \s9_data_i[30]_pad  ;
  input \s9_data_i[31]_pad  ;
  input \s9_data_i[3]_pad  ;
  input \s9_data_i[4]_pad  ;
  input \s9_data_i[5]_pad  ;
  input \s9_data_i[6]_pad  ;
  input \s9_data_i[7]_pad  ;
  input \s9_data_i[8]_pad  ;
  input \s9_data_i[9]_pad  ;
  input \s9_err_i_pad  ;
  input \s9_m0_cyc_r_reg/P0001  ;
  input \s9_m1_cyc_r_reg/P0001  ;
  input \s9_m2_cyc_r_reg/P0001  ;
  input \s9_m3_cyc_r_reg/P0001  ;
  input \s9_m4_cyc_r_reg/P0001  ;
  input \s9_m5_cyc_r_reg/P0001  ;
  input \s9_m6_cyc_r_reg/P0001  ;
  input \s9_m7_cyc_r_reg/P0001  ;
  input \s9_msel_arb0_state_reg[0]/NET0131  ;
  input \s9_msel_arb0_state_reg[1]/NET0131  ;
  input \s9_msel_arb0_state_reg[2]/NET0131  ;
  input \s9_msel_arb1_state_reg[0]/NET0131  ;
  input \s9_msel_arb1_state_reg[1]/NET0131  ;
  input \s9_msel_arb1_state_reg[2]/NET0131  ;
  input \s9_msel_arb2_state_reg[0]/NET0131  ;
  input \s9_msel_arb2_state_reg[1]/NET0131  ;
  input \s9_msel_arb2_state_reg[2]/NET0131  ;
  input \s9_msel_arb3_state_reg[0]/NET0131  ;
  input \s9_msel_arb3_state_reg[1]/NET0131  ;
  input \s9_msel_arb3_state_reg[2]/NET0131  ;
  input \s9_msel_pri_out_reg[0]/NET0131  ;
  input \s9_msel_pri_out_reg[1]/NET0131  ;
  input \s9_next_reg/P0001  ;
  input \s9_rty_i_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g106655/_1_  ;
  output \g106703/_1_  ;
  output \g69412/_0_  ;
  output \g69413/_0_  ;
  output \g69417/_1_  ;
  output \g69418/_0_  ;
  output \g69420/_1_  ;
  output \g69421/_0_  ;
  output \g69423/_1_  ;
  output \g69424/_0_  ;
  output \g69426/_1_  ;
  output \g69428/_1_  ;
  output \g69430/_1_  ;
  output \g69432/_1_  ;
  output \g69434/_1_  ;
  output \g69436/_1_  ;
  output \g69438/_1_  ;
  output \g69757/_2_  ;
  output \g69758/_2_  ;
  output \g69759/_2_  ;
  output \g69760/_2_  ;
  output \g69761/_0_  ;
  output \g69762/_2_  ;
  output \g69763/_2_  ;
  output \g69764/_2_  ;
  output \g69765/_2_  ;
  output \g69766/_2_  ;
  output \g69767/_0_  ;
  output \g69768/_0_  ;
  output \g69769/_0_  ;
  output \g69770/_0_  ;
  output \g69771/_0_  ;
  output \g69772/_0_  ;
  output \g70206/_0_  ;
  output \g70392/_0_  ;
  output \g70393/_0_  ;
  output \g70394/_0_  ;
  output \g70395/_0_  ;
  output \g70396/_0_  ;
  output \g70397/_0_  ;
  output \g70398/_0_  ;
  output \g70399/_0_  ;
  output \g70400/_0_  ;
  output \g70401/_0_  ;
  output \g70402/_0_  ;
  output \g70403/_0_  ;
  output \g70404/_0_  ;
  output \g70405/_0_  ;
  output \g70406/_0_  ;
  output \g70407/_0_  ;
  output \g70408/_0_  ;
  output \g70409/_0_  ;
  output \g70410/_0_  ;
  output \g70411/_0_  ;
  output \g70412/_0_  ;
  output \g70413/_0_  ;
  output \g70414/_0_  ;
  output \g70415/_0_  ;
  output \g70416/_0_  ;
  output \g70417/_0_  ;
  output \g70418/_0_  ;
  output \g70419/_0_  ;
  output \g70420/_0_  ;
  output \g70421/_0_  ;
  output \g70422/_0_  ;
  output \g70423/_0_  ;
  output \g70424/_0_  ;
  output \g70425/_0_  ;
  output \g70426/_0_  ;
  output \g70427/_0_  ;
  output \g70428/_0_  ;
  output \g70429/_0_  ;
  output \g70430/_0_  ;
  output \g70431/_0_  ;
  output \g70432/_0_  ;
  output \g70433/_0_  ;
  output \g70434/_0_  ;
  output \g70435/_0_  ;
  output \g70436/_0_  ;
  output \g70437/_0_  ;
  output \g70438/_0_  ;
  output \g70439/_0_  ;
  output \g70440/_0_  ;
  output \g70441/_0_  ;
  output \g70442/_0_  ;
  output \g70443/_0_  ;
  output \g70444/_0_  ;
  output \g70445/_0_  ;
  output \g70446/_0_  ;
  output \g70447/_0_  ;
  output \g70448/_0_  ;
  output \g70449/_0_  ;
  output \g70450/_0_  ;
  output \g70451/_0_  ;
  output \g70452/_0_  ;
  output \g70453/_0_  ;
  output \g70454/_0_  ;
  output \g70455/_0_  ;
  output \g70456/_0_  ;
  output \g70457/_0_  ;
  output \g70458/_0_  ;
  output \g70459/_0_  ;
  output \g70460/_0_  ;
  output \g70461/_0_  ;
  output \g70462/_0_  ;
  output \g70463/_0_  ;
  output \g70464/_0_  ;
  output \g70465/_0_  ;
  output \g70466/_0_  ;
  output \g70467/_0_  ;
  output \g70468/_0_  ;
  output \g70469/_0_  ;
  output \g70470/_0_  ;
  output \g70471/_0_  ;
  output \g70472/_0_  ;
  output \g70473/_0_  ;
  output \g70474/_0_  ;
  output \g70475/_0_  ;
  output \g70476/_0_  ;
  output \g70477/_0_  ;
  output \g70478/_0_  ;
  output \g70479/_0_  ;
  output \g70480/_0_  ;
  output \g70481/_0_  ;
  output \g70482/_0_  ;
  output \g70483/_0_  ;
  output \g70484/_0_  ;
  output \g70485/_0_  ;
  output \g70486/_0_  ;
  output \g70487/_0_  ;
  output \g70488/_0_  ;
  output \g70489/_0_  ;
  output \g70490/_0_  ;
  output \g70491/_0_  ;
  output \g70492/_0_  ;
  output \g70493/_0_  ;
  output \g70494/_0_  ;
  output \g70495/_0_  ;
  output \g70496/_0_  ;
  output \g70497/_0_  ;
  output \g70498/_0_  ;
  output \g70499/_0_  ;
  output \g70500/_0_  ;
  output \g70501/_0_  ;
  output \g70502/_0_  ;
  output \g70503/_0_  ;
  output \g70504/_0_  ;
  output \g70505/_0_  ;
  output \g70506/_0_  ;
  output \g70507/_0_  ;
  output \g70508/_0_  ;
  output \g70509/_0_  ;
  output \g70510/_0_  ;
  output \g70511/_0_  ;
  output \g70513/_0_  ;
  output \g70515/_0_  ;
  output \g70516/_0_  ;
  output \g70517/_0_  ;
  output \g70518/_0_  ;
  output \g70519/_0_  ;
  output \g70521/_0_  ;
  output \g70522/_0_  ;
  output \g70524/_0_  ;
  output \g70557/_0_  ;
  output \g70559/_0_  ;
  output \g70560/_0_  ;
  output \g70561/_0_  ;
  output \g70562/_0_  ;
  output \g70563/_0_  ;
  output \g70564/_0_  ;
  output \g70565/_0_  ;
  output \g70566/_0_  ;
  output \g70567/_0_  ;
  output \g70568/_0_  ;
  output \g70569/_0_  ;
  output \g70570/_0_  ;
  output \g70571/_0_  ;
  output \g70572/_0_  ;
  output \g70573/_0_  ;
  output \g70574/_0_  ;
  output \g70575/_0_  ;
  output \g70576/_0_  ;
  output \g70577/_0_  ;
  output \g70578/_0_  ;
  output \g70579/_0_  ;
  output \g70580/_0_  ;
  output \g70581/_0_  ;
  output \g70582/_0_  ;
  output \g70583/_0_  ;
  output \g70584/_0_  ;
  output \g70585/_0_  ;
  output \g70586/_0_  ;
  output \g70587/_0_  ;
  output \g70588/_0_  ;
  output \g70589/_0_  ;
  output \g70590/_0_  ;
  output \g70591/_0_  ;
  output \g70592/_0_  ;
  output \g70593/_0_  ;
  output \g70594/_0_  ;
  output \g70595/_0_  ;
  output \g70596/_0_  ;
  output \g70597/_0_  ;
  output \g70598/_0_  ;
  output \g70599/_0_  ;
  output \g70600/_0_  ;
  output \g70601/_0_  ;
  output \g70602/_0_  ;
  output \g70603/_0_  ;
  output \g70604/_0_  ;
  output \g70605/_0_  ;
  output \g70606/_0_  ;
  output \g70607/_0_  ;
  output \g70608/_0_  ;
  output \g70609/_0_  ;
  output \g70610/_0_  ;
  output \g70611/_0_  ;
  output \g70612/_0_  ;
  output \g70613/_0_  ;
  output \g70614/_0_  ;
  output \g70615/_0_  ;
  output \g70616/_0_  ;
  output \g70617/_0_  ;
  output \g70618/_0_  ;
  output \g70619/_0_  ;
  output \g70620/_0_  ;
  output \g70621/_0_  ;
  output \g70622/_0_  ;
  output \g70623/_0_  ;
  output \g70624/_0_  ;
  output \g70625/_0_  ;
  output \g70626/_0_  ;
  output \g70627/_0_  ;
  output \g70628/_0_  ;
  output \g70629/_0_  ;
  output \g70630/_0_  ;
  output \g70631/_0_  ;
  output \g70632/_0_  ;
  output \g70633/_0_  ;
  output \g70634/_0_  ;
  output \g70635/_0_  ;
  output \g70636/_0_  ;
  output \g70637/_0_  ;
  output \g70638/_0_  ;
  output \g70639/_0_  ;
  output \g70640/_0_  ;
  output \g70641/_0_  ;
  output \g70642/_0_  ;
  output \g70643/_0_  ;
  output \g70644/_0_  ;
  output \g70645/_0_  ;
  output \g70646/_0_  ;
  output \g70647/_0_  ;
  output \g70648/_0_  ;
  output \g70649/_0_  ;
  output \g70650/_0_  ;
  output \g70651/_0_  ;
  output \g70652/_0_  ;
  output \g70653/_0_  ;
  output \g70654/_0_  ;
  output \g70655/_0_  ;
  output \g70656/_0_  ;
  output \g70657/_0_  ;
  output \g70658/_0_  ;
  output \g70659/_0_  ;
  output \g70660/_0_  ;
  output \g70661/_0_  ;
  output \g70662/_0_  ;
  output \g70663/_0_  ;
  output \g70664/_0_  ;
  output \g70665/_0_  ;
  output \g70666/_0_  ;
  output \g70667/_0_  ;
  output \g70668/_0_  ;
  output \g70669/_0_  ;
  output \g70670/_0_  ;
  output \g70671/_0_  ;
  output \g70672/_0_  ;
  output \g70673/_0_  ;
  output \g70674/_0_  ;
  output \g70675/_0_  ;
  output \g70676/_0_  ;
  output \g70677/_0_  ;
  output \g70678/_0_  ;
  output \g70679/_0_  ;
  output \g70680/_0_  ;
  output \g70681/_0_  ;
  output \g70682/_0_  ;
  output \g70683/_0_  ;
  output \g70684/_0_  ;
  output \g70685/_0_  ;
  output \g70686/_0_  ;
  output \g70687/_0_  ;
  output \g70688/_0_  ;
  output \g70689/_0_  ;
  output \g70690/_0_  ;
  output \g70691/_0_  ;
  output \g70692/_0_  ;
  output \g70693/_0_  ;
  output \g70694/_0_  ;
  output \g70695/_0_  ;
  output \g70696/_0_  ;
  output \g70697/_0_  ;
  output \g70698/_0_  ;
  output \g70699/_0_  ;
  output \g70700/_0_  ;
  output \g70701/_0_  ;
  output \g70702/_0_  ;
  output \g70703/_0_  ;
  output \g70704/_0_  ;
  output \g70705/_0_  ;
  output \g70706/_0_  ;
  output \g70707/_0_  ;
  output \g70708/_0_  ;
  output \g70709/_0_  ;
  output \g70710/_0_  ;
  output \g70711/_0_  ;
  output \g70712/_0_  ;
  output \g70713/_0_  ;
  output \g70714/_0_  ;
  output \g70715/_0_  ;
  output \g70716/_0_  ;
  output \g70717/_0_  ;
  output \g70718/_0_  ;
  output \g70719/_0_  ;
  output \g70720/_0_  ;
  output \g70721/_0_  ;
  output \g70722/_0_  ;
  output \g70723/_0_  ;
  output \g70724/_0_  ;
  output \g70725/_0_  ;
  output \g70726/_0_  ;
  output \g70727/_0_  ;
  output \g70728/_0_  ;
  output \g70729/_0_  ;
  output \g70730/_0_  ;
  output \g70731/_0_  ;
  output \g70732/_0_  ;
  output \g70733/_0_  ;
  output \g70734/_0_  ;
  output \g70735/_0_  ;
  output \g70736/_0_  ;
  output \g70737/_0_  ;
  output \g70738/_0_  ;
  output \g70739/_0_  ;
  output \g70740/_0_  ;
  output \g70741/_0_  ;
  output \g70742/_0_  ;
  output \g70743/_0_  ;
  output \g70744/_0_  ;
  output \g70745/_0_  ;
  output \g70746/_0_  ;
  output \g70747/_0_  ;
  output \g70748/_0_  ;
  output \g70749/_0_  ;
  output \g70750/_0_  ;
  output \g70751/_0_  ;
  output \g70752/_0_  ;
  output \g70753/_0_  ;
  output \g70754/_0_  ;
  output \g70755/_0_  ;
  output \g70756/_0_  ;
  output \g70757/_0_  ;
  output \g70758/_0_  ;
  output \g70759/_0_  ;
  output \g70760/_0_  ;
  output \g70761/_0_  ;
  output \g70762/_0_  ;
  output \g70763/_0_  ;
  output \g70764/_0_  ;
  output \g70765/_0_  ;
  output \g70766/_0_  ;
  output \g70767/_0_  ;
  output \g70768/_0_  ;
  output \g70769/_0_  ;
  output \g70770/_0_  ;
  output \g70771/_0_  ;
  output \g70772/_0_  ;
  output \g70773/_0_  ;
  output \g70774/_0_  ;
  output \g70775/_0_  ;
  output \g70776/_0_  ;
  output \g70777/_0_  ;
  output \g70778/_0_  ;
  output \g70779/_0_  ;
  output \g70780/_0_  ;
  output \g70781/_0_  ;
  output \g70782/_0_  ;
  output \g70783/_0_  ;
  output \g70784/_0_  ;
  output \g70785/_0_  ;
  output \g70786/_0_  ;
  output \g70787/_0_  ;
  output \g70788/_0_  ;
  output \g70789/_0_  ;
  output \g70790/_0_  ;
  output \g70791/_0_  ;
  output \g70792/_0_  ;
  output \g70793/_0_  ;
  output \g70794/_0_  ;
  output \g70795/_0_  ;
  output \g70796/_0_  ;
  output \g70797/_0_  ;
  output \g70798/_0_  ;
  output \g70799/_0_  ;
  output \g70800/_0_  ;
  output \g70801/_0_  ;
  output \g70802/_0_  ;
  output \g70803/_0_  ;
  output \g70804/_0_  ;
  output \g70805/_0_  ;
  output \g70806/_0_  ;
  output \g70807/_0_  ;
  output \g70808/_0_  ;
  output \g70809/_0_  ;
  output \g70810/_0_  ;
  output \g70811/_0_  ;
  output \g70812/_0_  ;
  output \g70813/_0_  ;
  output \g70814/_0_  ;
  output \g70815/_0_  ;
  output \g70816/_0_  ;
  output \g70817/_0_  ;
  output \g70818/_0_  ;
  output \g70819/_0_  ;
  output \g70820/_0_  ;
  output \g70821/_0_  ;
  output \g70822/_0_  ;
  output \g70823/_0_  ;
  output \g70824/_0_  ;
  output \g70825/_0_  ;
  output \g70826/_0_  ;
  output \g70827/_0_  ;
  output \g70828/_0_  ;
  output \g70829/_0_  ;
  output \g70830/_0_  ;
  output \g70831/_0_  ;
  output \g70832/_0_  ;
  output \g70833/_0_  ;
  output \g70834/_0_  ;
  output \g70835/_0_  ;
  output \g70836/_0_  ;
  output \g70837/_0_  ;
  output \g70838/_0_  ;
  output \g70839/_0_  ;
  output \g70840/_0_  ;
  output \g70841/_0_  ;
  output \g70842/_0_  ;
  output \g70843/_0_  ;
  output \g70844/_0_  ;
  output \g70845/_0_  ;
  output \g70846/_0_  ;
  output \g70847/_0_  ;
  output \g70848/_0_  ;
  output \g70849/_0_  ;
  output \g70850/_0_  ;
  output \g70851/_0_  ;
  output \g70852/_0_  ;
  output \g70853/_0_  ;
  output \g70854/_0_  ;
  output \g70855/_0_  ;
  output \g70856/_0_  ;
  output \g70857/_0_  ;
  output \g70858/_0_  ;
  output \g70859/_0_  ;
  output \g70860/_0_  ;
  output \g70861/_0_  ;
  output \g71404/_0_  ;
  output \g71407/_0_  ;
  output \g72631/_0_  ;
  output \g72631/_1_  ;
  output \g72633/_0_  ;
  output \g72642/_0_  ;
  output \g72649/_0_  ;
  output \g72649/_1_  ;
  output \g72652/_0_  ;
  output \g72660/_0_  ;
  output \g72666/_0_  ;
  output \g72666/_1_  ;
  output \g72671/_0_  ;
  output \g72681/_0_  ;
  output \g72681/_1_  ;
  output \g72689/_0_  ;
  output \g72696/_0_  ;
  output \g72696/_1_  ;
  output \g72698/_0_  ;
  output \g72707/_0_  ;
  output \g72715/_0_  ;
  output \g72715/_1_  ;
  output \g72718/_0_  ;
  output \g72726/_0_  ;
  output \g72732/_0_  ;
  output \g72732/_1_  ;
  output \g72736/_0_  ;
  output \g72743/_0_  ;
  output \g72745/_0_  ;
  output \g72745/_1_  ;
  output \g72752/_0_  ;
  output \g72752/_1_  ;
  output \g72756/_0_  ;
  output \g72763/_0_  ;
  output \g72763/_1_  ;
  output \g72765/_0_  ;
  output \g72767/_0_  ;
  output \g72767/_1_  ;
  output \g72769/_0_  ;
  output \g72769/_1_  ;
  output \g72772/_0_  ;
  output \g72772/_1_  ;
  output \g72774/_0_  ;
  output \g72774/_1_  ;
  output \g72790/_0_  ;
  output \g72790/_1_  ;
  output \g72797/_0_  ;
  output \g73807/_0_  ;
  output \g73820/_0_  ;
  output \g73832/_0_  ;
  output \g73844/_0_  ;
  output \g73856/_0_  ;
  output \g73871/_0_  ;
  output \g73883/_0_  ;
  output \g73895/_0_  ;
  output \g73905/_3_  ;
  output \g73910/_0_  ;
  output \g73922/_0_  ;
  output \g73934/_0_  ;
  output \g73946/_0_  ;
  output \g73958/_0_  ;
  output \g73970/_0_  ;
  output \g73982/_0_  ;
  output \g87036/_0_  ;
  output \g87042/_0_  ;
  output \g87043/_0_  ;
  output \g87044/_0_  ;
  output \g87045/_0_  ;
  output \g87046/_0_  ;
  output \g87047/_0_  ;
  output \g87048/_0_  ;
  output \g87049/_0_  ;
  output \g87050/_0_  ;
  output \g87051/_0_  ;
  output \g87052/_0_  ;
  output \g87053/_0_  ;
  output \g87054/_0_  ;
  output \g87055/_0_  ;
  output \g87062/_0_  ;
  output \g88572/_0_  ;
  output \g88681/_0_  ;
  output \g88682/_0_  ;
  output \g88683/_0_  ;
  output \g88684/_0_  ;
  output \g88685/_0_  ;
  output \g88686/_0_  ;
  output \g88687/_0_  ;
  output \g88688/_0_  ;
  output \g88689/_0_  ;
  output \g88690/_0_  ;
  output \g88691/_0_  ;
  output \g88692/_0_  ;
  output \g88693/_0_  ;
  output \g88695/_0_  ;
  output \g88697/_0_  ;
  output \g88698/_0_  ;
  output \g88700/_0_  ;
  output \g88701/_0_  ;
  output \g88703/_0_  ;
  output \g88704/_0_  ;
  output \g88705/_0_  ;
  output \g88706/_0_  ;
  output \g88707/_0_  ;
  output \g88709/_0_  ;
  output \g88710/_0_  ;
  output \g88711/_0_  ;
  output \g88712/_0_  ;
  output \g88713/_0_  ;
  output \g88714/_0_  ;
  output \g88716/_0_  ;
  output \g88717/_0_  ;
  output \g88718/_0_  ;
  output \g88719/_0_  ;
  output \g88720/_0_  ;
  output \g88722/_0_  ;
  output \g88723/_0_  ;
  output \g88724/_0_  ;
  output \g88725/_0_  ;
  output \g88726/_0_  ;
  output \g88727/_0_  ;
  output \g88728/_0_  ;
  output \g88729/_0_  ;
  output \g88731/_0_  ;
  output \g88732/_0_  ;
  output \g88733/_0_  ;
  output \g88734/_0_  ;
  output \g88736/_0_  ;
  output \g88737/_0_  ;
  output \g88738/_0_  ;
  output \g88739/_0_  ;
  output \g88740/_0_  ;
  output \g88741/_0_  ;
  output \g88742/_0_  ;
  output \g88743/_0_  ;
  output \g88744/_0_  ;
  output \g88745/_0_  ;
  output \g88746/_0_  ;
  output \g88748/_0_  ;
  output \g88749/_0_  ;
  output \g88750/_0_  ;
  output \g88752/_0_  ;
  output \g88753/_0_  ;
  output \g88754/_0_  ;
  output \g88755/_0_  ;
  output \g88756/_0_  ;
  output \g88757/_0_  ;
  output \g88759/_0_  ;
  output \g88760/_0_  ;
  output \g88761/_0_  ;
  output \g88762/_0_  ;
  output \g88764/_0_  ;
  output \g88765/_0_  ;
  output \g88766/_0_  ;
  output \g88768/_0_  ;
  output \g88769/_0_  ;
  output \g88770/_0_  ;
  output \g88771/_0_  ;
  output \g88772/_0_  ;
  output \g88773/_0_  ;
  output \g88775/_0_  ;
  output \g88776/_0_  ;
  output \g88777/_0_  ;
  output \g88778/_0_  ;
  output \g88779/_0_  ;
  output \g88780/_0_  ;
  output \g88782/_0_  ;
  output \g88783/_0_  ;
  output \g88784/_0_  ;
  output \g88785/_0_  ;
  output \g88786/_0_  ;
  output \g88787/_0_  ;
  output \g88789/_0_  ;
  output \g88790/_0_  ;
  output \g88791/_0_  ;
  output \g88792/_0_  ;
  output \g88793/_0_  ;
  output \g88795/_0_  ;
  output \g88796/_0_  ;
  output \g88797/_0_  ;
  output \g88799/_0_  ;
  output \g88800/_0_  ;
  output \g88801/_0_  ;
  output \g88802/_0_  ;
  output \g88806/_0_  ;
  output \g88807/_0_  ;
  output \g88808/_0_  ;
  output \g88809/_0_  ;
  output \g88810/_0_  ;
  output \g88813/_0_  ;
  output \g88814/_0_  ;
  output \g88815/_0_  ;
  output \m0_ack_o_pad  ;
  output \m0_data_o[0]_pad  ;
  output \m0_data_o[10]_pad  ;
  output \m0_data_o[11]_pad  ;
  output \m0_data_o[12]_pad  ;
  output \m0_data_o[13]_pad  ;
  output \m0_data_o[14]_pad  ;
  output \m0_data_o[15]_pad  ;
  output \m0_data_o[16]_pad  ;
  output \m0_data_o[17]_pad  ;
  output \m0_data_o[18]_pad  ;
  output \m0_data_o[19]_pad  ;
  output \m0_data_o[1]_pad  ;
  output \m0_data_o[20]_pad  ;
  output \m0_data_o[21]_pad  ;
  output \m0_data_o[22]_pad  ;
  output \m0_data_o[23]_pad  ;
  output \m0_data_o[24]_pad  ;
  output \m0_data_o[25]_pad  ;
  output \m0_data_o[26]_pad  ;
  output \m0_data_o[27]_pad  ;
  output \m0_data_o[28]_pad  ;
  output \m0_data_o[29]_pad  ;
  output \m0_data_o[2]_pad  ;
  output \m0_data_o[30]_pad  ;
  output \m0_data_o[31]_pad  ;
  output \m0_data_o[3]_pad  ;
  output \m0_data_o[4]_pad  ;
  output \m0_data_o[5]_pad  ;
  output \m0_data_o[6]_pad  ;
  output \m0_data_o[7]_pad  ;
  output \m0_data_o[8]_pad  ;
  output \m0_data_o[9]_pad  ;
  output \m0_err_o_pad  ;
  output \m0_rty_o_pad  ;
  output \m1_ack_o_pad  ;
  output \m1_data_o[0]_pad  ;
  output \m1_data_o[10]_pad  ;
  output \m1_data_o[11]_pad  ;
  output \m1_data_o[12]_pad  ;
  output \m1_data_o[13]_pad  ;
  output \m1_data_o[14]_pad  ;
  output \m1_data_o[15]_pad  ;
  output \m1_data_o[16]_pad  ;
  output \m1_data_o[17]_pad  ;
  output \m1_data_o[18]_pad  ;
  output \m1_data_o[19]_pad  ;
  output \m1_data_o[1]_pad  ;
  output \m1_data_o[20]_pad  ;
  output \m1_data_o[21]_pad  ;
  output \m1_data_o[22]_pad  ;
  output \m1_data_o[23]_pad  ;
  output \m1_data_o[24]_pad  ;
  output \m1_data_o[25]_pad  ;
  output \m1_data_o[26]_pad  ;
  output \m1_data_o[27]_pad  ;
  output \m1_data_o[28]_pad  ;
  output \m1_data_o[29]_pad  ;
  output \m1_data_o[2]_pad  ;
  output \m1_data_o[30]_pad  ;
  output \m1_data_o[31]_pad  ;
  output \m1_data_o[3]_pad  ;
  output \m1_data_o[4]_pad  ;
  output \m1_data_o[5]_pad  ;
  output \m1_data_o[6]_pad  ;
  output \m1_data_o[7]_pad  ;
  output \m1_data_o[8]_pad  ;
  output \m1_data_o[9]_pad  ;
  output \m1_err_o_pad  ;
  output \m1_rty_o_pad  ;
  output \m2_ack_o_pad  ;
  output \m2_data_o[0]_pad  ;
  output \m2_data_o[10]_pad  ;
  output \m2_data_o[11]_pad  ;
  output \m2_data_o[12]_pad  ;
  output \m2_data_o[13]_pad  ;
  output \m2_data_o[14]_pad  ;
  output \m2_data_o[15]_pad  ;
  output \m2_data_o[16]_pad  ;
  output \m2_data_o[17]_pad  ;
  output \m2_data_o[18]_pad  ;
  output \m2_data_o[19]_pad  ;
  output \m2_data_o[1]_pad  ;
  output \m2_data_o[20]_pad  ;
  output \m2_data_o[21]_pad  ;
  output \m2_data_o[22]_pad  ;
  output \m2_data_o[23]_pad  ;
  output \m2_data_o[24]_pad  ;
  output \m2_data_o[25]_pad  ;
  output \m2_data_o[26]_pad  ;
  output \m2_data_o[27]_pad  ;
  output \m2_data_o[28]_pad  ;
  output \m2_data_o[29]_pad  ;
  output \m2_data_o[2]_pad  ;
  output \m2_data_o[30]_pad  ;
  output \m2_data_o[31]_pad  ;
  output \m2_data_o[3]_pad  ;
  output \m2_data_o[4]_pad  ;
  output \m2_data_o[5]_pad  ;
  output \m2_data_o[6]_pad  ;
  output \m2_data_o[7]_pad  ;
  output \m2_data_o[8]_pad  ;
  output \m2_data_o[9]_pad  ;
  output \m2_err_o_pad  ;
  output \m2_rty_o_pad  ;
  output \m3_ack_o_pad  ;
  output \m3_data_o[0]_pad  ;
  output \m3_data_o[10]_pad  ;
  output \m3_data_o[11]_pad  ;
  output \m3_data_o[12]_pad  ;
  output \m3_data_o[13]_pad  ;
  output \m3_data_o[14]_pad  ;
  output \m3_data_o[15]_pad  ;
  output \m3_data_o[16]_pad  ;
  output \m3_data_o[17]_pad  ;
  output \m3_data_o[18]_pad  ;
  output \m3_data_o[19]_pad  ;
  output \m3_data_o[1]_pad  ;
  output \m3_data_o[20]_pad  ;
  output \m3_data_o[21]_pad  ;
  output \m3_data_o[22]_pad  ;
  output \m3_data_o[23]_pad  ;
  output \m3_data_o[24]_pad  ;
  output \m3_data_o[25]_pad  ;
  output \m3_data_o[26]_pad  ;
  output \m3_data_o[27]_pad  ;
  output \m3_data_o[28]_pad  ;
  output \m3_data_o[29]_pad  ;
  output \m3_data_o[2]_pad  ;
  output \m3_data_o[30]_pad  ;
  output \m3_data_o[31]_pad  ;
  output \m3_data_o[3]_pad  ;
  output \m3_data_o[4]_pad  ;
  output \m3_data_o[5]_pad  ;
  output \m3_data_o[6]_pad  ;
  output \m3_data_o[7]_pad  ;
  output \m3_data_o[8]_pad  ;
  output \m3_data_o[9]_pad  ;
  output \m3_err_o_pad  ;
  output \m3_rty_o_pad  ;
  output \m4_ack_o_pad  ;
  output \m4_data_o[0]_pad  ;
  output \m4_data_o[10]_pad  ;
  output \m4_data_o[11]_pad  ;
  output \m4_data_o[12]_pad  ;
  output \m4_data_o[13]_pad  ;
  output \m4_data_o[14]_pad  ;
  output \m4_data_o[15]_pad  ;
  output \m4_data_o[16]_pad  ;
  output \m4_data_o[17]_pad  ;
  output \m4_data_o[18]_pad  ;
  output \m4_data_o[19]_pad  ;
  output \m4_data_o[1]_pad  ;
  output \m4_data_o[20]_pad  ;
  output \m4_data_o[21]_pad  ;
  output \m4_data_o[22]_pad  ;
  output \m4_data_o[23]_pad  ;
  output \m4_data_o[24]_pad  ;
  output \m4_data_o[25]_pad  ;
  output \m4_data_o[26]_pad  ;
  output \m4_data_o[27]_pad  ;
  output \m4_data_o[28]_pad  ;
  output \m4_data_o[29]_pad  ;
  output \m4_data_o[2]_pad  ;
  output \m4_data_o[30]_pad  ;
  output \m4_data_o[31]_pad  ;
  output \m4_data_o[3]_pad  ;
  output \m4_data_o[4]_pad  ;
  output \m4_data_o[5]_pad  ;
  output \m4_data_o[6]_pad  ;
  output \m4_data_o[7]_pad  ;
  output \m4_data_o[8]_pad  ;
  output \m4_data_o[9]_pad  ;
  output \m4_err_o_pad  ;
  output \m4_rty_o_pad  ;
  output \m5_ack_o_pad  ;
  output \m5_data_o[0]_pad  ;
  output \m5_data_o[10]_pad  ;
  output \m5_data_o[11]_pad  ;
  output \m5_data_o[12]_pad  ;
  output \m5_data_o[13]_pad  ;
  output \m5_data_o[14]_pad  ;
  output \m5_data_o[15]_pad  ;
  output \m5_data_o[16]_pad  ;
  output \m5_data_o[17]_pad  ;
  output \m5_data_o[18]_pad  ;
  output \m5_data_o[19]_pad  ;
  output \m5_data_o[1]_pad  ;
  output \m5_data_o[20]_pad  ;
  output \m5_data_o[21]_pad  ;
  output \m5_data_o[22]_pad  ;
  output \m5_data_o[23]_pad  ;
  output \m5_data_o[24]_pad  ;
  output \m5_data_o[25]_pad  ;
  output \m5_data_o[26]_pad  ;
  output \m5_data_o[27]_pad  ;
  output \m5_data_o[28]_pad  ;
  output \m5_data_o[29]_pad  ;
  output \m5_data_o[2]_pad  ;
  output \m5_data_o[30]_pad  ;
  output \m5_data_o[31]_pad  ;
  output \m5_data_o[3]_pad  ;
  output \m5_data_o[4]_pad  ;
  output \m5_data_o[5]_pad  ;
  output \m5_data_o[6]_pad  ;
  output \m5_data_o[7]_pad  ;
  output \m5_data_o[8]_pad  ;
  output \m5_data_o[9]_pad  ;
  output \m5_err_o_pad  ;
  output \m5_rty_o_pad  ;
  output \m6_ack_o_pad  ;
  output \m6_data_o[0]_pad  ;
  output \m6_data_o[10]_pad  ;
  output \m6_data_o[11]_pad  ;
  output \m6_data_o[12]_pad  ;
  output \m6_data_o[13]_pad  ;
  output \m6_data_o[14]_pad  ;
  output \m6_data_o[15]_pad  ;
  output \m6_data_o[16]_pad  ;
  output \m6_data_o[17]_pad  ;
  output \m6_data_o[18]_pad  ;
  output \m6_data_o[19]_pad  ;
  output \m6_data_o[1]_pad  ;
  output \m6_data_o[20]_pad  ;
  output \m6_data_o[21]_pad  ;
  output \m6_data_o[22]_pad  ;
  output \m6_data_o[23]_pad  ;
  output \m6_data_o[24]_pad  ;
  output \m6_data_o[25]_pad  ;
  output \m6_data_o[26]_pad  ;
  output \m6_data_o[27]_pad  ;
  output \m6_data_o[28]_pad  ;
  output \m6_data_o[29]_pad  ;
  output \m6_data_o[2]_pad  ;
  output \m6_data_o[30]_pad  ;
  output \m6_data_o[31]_pad  ;
  output \m6_data_o[3]_pad  ;
  output \m6_data_o[4]_pad  ;
  output \m6_data_o[5]_pad  ;
  output \m6_data_o[6]_pad  ;
  output \m6_data_o[7]_pad  ;
  output \m6_data_o[8]_pad  ;
  output \m6_data_o[9]_pad  ;
  output \m6_err_o_pad  ;
  output \m6_rty_o_pad  ;
  output \m7_ack_o_pad  ;
  output \m7_data_o[0]_pad  ;
  output \m7_data_o[10]_pad  ;
  output \m7_data_o[11]_pad  ;
  output \m7_data_o[12]_pad  ;
  output \m7_data_o[13]_pad  ;
  output \m7_data_o[14]_pad  ;
  output \m7_data_o[15]_pad  ;
  output \m7_data_o[16]_pad  ;
  output \m7_data_o[17]_pad  ;
  output \m7_data_o[18]_pad  ;
  output \m7_data_o[19]_pad  ;
  output \m7_data_o[1]_pad  ;
  output \m7_data_o[20]_pad  ;
  output \m7_data_o[21]_pad  ;
  output \m7_data_o[22]_pad  ;
  output \m7_data_o[23]_pad  ;
  output \m7_data_o[24]_pad  ;
  output \m7_data_o[25]_pad  ;
  output \m7_data_o[26]_pad  ;
  output \m7_data_o[27]_pad  ;
  output \m7_data_o[28]_pad  ;
  output \m7_data_o[29]_pad  ;
  output \m7_data_o[2]_pad  ;
  output \m7_data_o[30]_pad  ;
  output \m7_data_o[31]_pad  ;
  output \m7_data_o[3]_pad  ;
  output \m7_data_o[4]_pad  ;
  output \m7_data_o[5]_pad  ;
  output \m7_data_o[6]_pad  ;
  output \m7_data_o[7]_pad  ;
  output \m7_data_o[8]_pad  ;
  output \m7_data_o[9]_pad  ;
  output \m7_err_o_pad  ;
  output \m7_rty_o_pad  ;
  output \s0_addr_o[0]_pad  ;
  output \s0_addr_o[10]_pad  ;
  output \s0_addr_o[11]_pad  ;
  output \s0_addr_o[12]_pad  ;
  output \s0_addr_o[13]_pad  ;
  output \s0_addr_o[14]_pad  ;
  output \s0_addr_o[15]_pad  ;
  output \s0_addr_o[16]_pad  ;
  output \s0_addr_o[17]_pad  ;
  output \s0_addr_o[18]_pad  ;
  output \s0_addr_o[19]_pad  ;
  output \s0_addr_o[1]_pad  ;
  output \s0_addr_o[20]_pad  ;
  output \s0_addr_o[21]_pad  ;
  output \s0_addr_o[22]_pad  ;
  output \s0_addr_o[23]_pad  ;
  output \s0_addr_o[24]_pad  ;
  output \s0_addr_o[25]_pad  ;
  output \s0_addr_o[26]_pad  ;
  output \s0_addr_o[27]_pad  ;
  output \s0_addr_o[28]_pad  ;
  output \s0_addr_o[29]_pad  ;
  output \s0_addr_o[2]_pad  ;
  output \s0_addr_o[30]_pad  ;
  output \s0_addr_o[31]_pad  ;
  output \s0_addr_o[3]_pad  ;
  output \s0_addr_o[4]_pad  ;
  output \s0_addr_o[5]_pad  ;
  output \s0_addr_o[6]_pad  ;
  output \s0_addr_o[7]_pad  ;
  output \s0_addr_o[8]_pad  ;
  output \s0_addr_o[9]_pad  ;
  output \s0_data_o[0]_pad  ;
  output \s0_data_o[10]_pad  ;
  output \s0_data_o[11]_pad  ;
  output \s0_data_o[12]_pad  ;
  output \s0_data_o[13]_pad  ;
  output \s0_data_o[14]_pad  ;
  output \s0_data_o[15]_pad  ;
  output \s0_data_o[16]_pad  ;
  output \s0_data_o[17]_pad  ;
  output \s0_data_o[18]_pad  ;
  output \s0_data_o[19]_pad  ;
  output \s0_data_o[1]_pad  ;
  output \s0_data_o[20]_pad  ;
  output \s0_data_o[21]_pad  ;
  output \s0_data_o[22]_pad  ;
  output \s0_data_o[23]_pad  ;
  output \s0_data_o[24]_pad  ;
  output \s0_data_o[25]_pad  ;
  output \s0_data_o[26]_pad  ;
  output \s0_data_o[27]_pad  ;
  output \s0_data_o[28]_pad  ;
  output \s0_data_o[29]_pad  ;
  output \s0_data_o[2]_pad  ;
  output \s0_data_o[30]_pad  ;
  output \s0_data_o[31]_pad  ;
  output \s0_data_o[3]_pad  ;
  output \s0_data_o[4]_pad  ;
  output \s0_data_o[5]_pad  ;
  output \s0_data_o[6]_pad  ;
  output \s0_data_o[7]_pad  ;
  output \s0_data_o[8]_pad  ;
  output \s0_data_o[9]_pad  ;
  output \s0_sel_o[0]_pad  ;
  output \s0_sel_o[1]_pad  ;
  output \s0_sel_o[2]_pad  ;
  output \s0_sel_o[3]_pad  ;
  output \s0_stb_o_pad  ;
  output \s0_we_o_pad  ;
  output \s10_addr_o[0]_pad  ;
  output \s10_addr_o[10]_pad  ;
  output \s10_addr_o[11]_pad  ;
  output \s10_addr_o[12]_pad  ;
  output \s10_addr_o[13]_pad  ;
  output \s10_addr_o[14]_pad  ;
  output \s10_addr_o[15]_pad  ;
  output \s10_addr_o[16]_pad  ;
  output \s10_addr_o[17]_pad  ;
  output \s10_addr_o[18]_pad  ;
  output \s10_addr_o[19]_pad  ;
  output \s10_addr_o[1]_pad  ;
  output \s10_addr_o[20]_pad  ;
  output \s10_addr_o[21]_pad  ;
  output \s10_addr_o[22]_pad  ;
  output \s10_addr_o[23]_pad  ;
  output \s10_addr_o[24]_pad  ;
  output \s10_addr_o[25]_pad  ;
  output \s10_addr_o[26]_pad  ;
  output \s10_addr_o[27]_pad  ;
  output \s10_addr_o[28]_pad  ;
  output \s10_addr_o[29]_pad  ;
  output \s10_addr_o[2]_pad  ;
  output \s10_addr_o[30]_pad  ;
  output \s10_addr_o[31]_pad  ;
  output \s10_addr_o[3]_pad  ;
  output \s10_addr_o[4]_pad  ;
  output \s10_addr_o[5]_pad  ;
  output \s10_addr_o[6]_pad  ;
  output \s10_addr_o[7]_pad  ;
  output \s10_addr_o[8]_pad  ;
  output \s10_addr_o[9]_pad  ;
  output \s10_data_o[0]_pad  ;
  output \s10_data_o[10]_pad  ;
  output \s10_data_o[11]_pad  ;
  output \s10_data_o[12]_pad  ;
  output \s10_data_o[13]_pad  ;
  output \s10_data_o[14]_pad  ;
  output \s10_data_o[15]_pad  ;
  output \s10_data_o[16]_pad  ;
  output \s10_data_o[17]_pad  ;
  output \s10_data_o[18]_pad  ;
  output \s10_data_o[19]_pad  ;
  output \s10_data_o[1]_pad  ;
  output \s10_data_o[20]_pad  ;
  output \s10_data_o[21]_pad  ;
  output \s10_data_o[22]_pad  ;
  output \s10_data_o[23]_pad  ;
  output \s10_data_o[24]_pad  ;
  output \s10_data_o[25]_pad  ;
  output \s10_data_o[26]_pad  ;
  output \s10_data_o[27]_pad  ;
  output \s10_data_o[28]_pad  ;
  output \s10_data_o[29]_pad  ;
  output \s10_data_o[2]_pad  ;
  output \s10_data_o[30]_pad  ;
  output \s10_data_o[31]_pad  ;
  output \s10_data_o[3]_pad  ;
  output \s10_data_o[4]_pad  ;
  output \s10_data_o[5]_pad  ;
  output \s10_data_o[6]_pad  ;
  output \s10_data_o[7]_pad  ;
  output \s10_data_o[8]_pad  ;
  output \s10_data_o[9]_pad  ;
  output \s10_sel_o[0]_pad  ;
  output \s10_sel_o[1]_pad  ;
  output \s10_sel_o[2]_pad  ;
  output \s10_sel_o[3]_pad  ;
  output \s10_stb_o_pad  ;
  output \s10_we_o_pad  ;
  output \s11_addr_o[0]_pad  ;
  output \s11_addr_o[10]_pad  ;
  output \s11_addr_o[11]_pad  ;
  output \s11_addr_o[12]_pad  ;
  output \s11_addr_o[13]_pad  ;
  output \s11_addr_o[14]_pad  ;
  output \s11_addr_o[15]_pad  ;
  output \s11_addr_o[16]_pad  ;
  output \s11_addr_o[17]_pad  ;
  output \s11_addr_o[18]_pad  ;
  output \s11_addr_o[19]_pad  ;
  output \s11_addr_o[1]_pad  ;
  output \s11_addr_o[20]_pad  ;
  output \s11_addr_o[21]_pad  ;
  output \s11_addr_o[22]_pad  ;
  output \s11_addr_o[23]_pad  ;
  output \s11_addr_o[24]_pad  ;
  output \s11_addr_o[25]_pad  ;
  output \s11_addr_o[26]_pad  ;
  output \s11_addr_o[27]_pad  ;
  output \s11_addr_o[28]_pad  ;
  output \s11_addr_o[29]_pad  ;
  output \s11_addr_o[2]_pad  ;
  output \s11_addr_o[30]_pad  ;
  output \s11_addr_o[31]_pad  ;
  output \s11_addr_o[3]_pad  ;
  output \s11_addr_o[4]_pad  ;
  output \s11_addr_o[5]_pad  ;
  output \s11_addr_o[6]_pad  ;
  output \s11_addr_o[7]_pad  ;
  output \s11_addr_o[8]_pad  ;
  output \s11_addr_o[9]_pad  ;
  output \s11_data_o[0]_pad  ;
  output \s11_data_o[10]_pad  ;
  output \s11_data_o[11]_pad  ;
  output \s11_data_o[12]_pad  ;
  output \s11_data_o[13]_pad  ;
  output \s11_data_o[14]_pad  ;
  output \s11_data_o[15]_pad  ;
  output \s11_data_o[16]_pad  ;
  output \s11_data_o[17]_pad  ;
  output \s11_data_o[18]_pad  ;
  output \s11_data_o[19]_pad  ;
  output \s11_data_o[1]_pad  ;
  output \s11_data_o[20]_pad  ;
  output \s11_data_o[21]_pad  ;
  output \s11_data_o[22]_pad  ;
  output \s11_data_o[23]_pad  ;
  output \s11_data_o[24]_pad  ;
  output \s11_data_o[25]_pad  ;
  output \s11_data_o[26]_pad  ;
  output \s11_data_o[27]_pad  ;
  output \s11_data_o[28]_pad  ;
  output \s11_data_o[29]_pad  ;
  output \s11_data_o[2]_pad  ;
  output \s11_data_o[30]_pad  ;
  output \s11_data_o[31]_pad  ;
  output \s11_data_o[3]_pad  ;
  output \s11_data_o[4]_pad  ;
  output \s11_data_o[5]_pad  ;
  output \s11_data_o[6]_pad  ;
  output \s11_data_o[7]_pad  ;
  output \s11_data_o[8]_pad  ;
  output \s11_data_o[9]_pad  ;
  output \s11_sel_o[0]_pad  ;
  output \s11_sel_o[1]_pad  ;
  output \s11_sel_o[2]_pad  ;
  output \s11_sel_o[3]_pad  ;
  output \s11_stb_o_pad  ;
  output \s11_we_o_pad  ;
  output \s12_addr_o[0]_pad  ;
  output \s12_addr_o[10]_pad  ;
  output \s12_addr_o[11]_pad  ;
  output \s12_addr_o[12]_pad  ;
  output \s12_addr_o[13]_pad  ;
  output \s12_addr_o[14]_pad  ;
  output \s12_addr_o[15]_pad  ;
  output \s12_addr_o[16]_pad  ;
  output \s12_addr_o[17]_pad  ;
  output \s12_addr_o[18]_pad  ;
  output \s12_addr_o[19]_pad  ;
  output \s12_addr_o[1]_pad  ;
  output \s12_addr_o[20]_pad  ;
  output \s12_addr_o[21]_pad  ;
  output \s12_addr_o[22]_pad  ;
  output \s12_addr_o[23]_pad  ;
  output \s12_addr_o[24]_pad  ;
  output \s12_addr_o[25]_pad  ;
  output \s12_addr_o[26]_pad  ;
  output \s12_addr_o[27]_pad  ;
  output \s12_addr_o[28]_pad  ;
  output \s12_addr_o[29]_pad  ;
  output \s12_addr_o[2]_pad  ;
  output \s12_addr_o[30]_pad  ;
  output \s12_addr_o[31]_pad  ;
  output \s12_addr_o[3]_pad  ;
  output \s12_addr_o[4]_pad  ;
  output \s12_addr_o[5]_pad  ;
  output \s12_addr_o[6]_pad  ;
  output \s12_addr_o[7]_pad  ;
  output \s12_addr_o[8]_pad  ;
  output \s12_addr_o[9]_pad  ;
  output \s12_data_o[0]_pad  ;
  output \s12_data_o[10]_pad  ;
  output \s12_data_o[11]_pad  ;
  output \s12_data_o[12]_pad  ;
  output \s12_data_o[13]_pad  ;
  output \s12_data_o[14]_pad  ;
  output \s12_data_o[15]_pad  ;
  output \s12_data_o[16]_pad  ;
  output \s12_data_o[17]_pad  ;
  output \s12_data_o[18]_pad  ;
  output \s12_data_o[19]_pad  ;
  output \s12_data_o[1]_pad  ;
  output \s12_data_o[20]_pad  ;
  output \s12_data_o[21]_pad  ;
  output \s12_data_o[22]_pad  ;
  output \s12_data_o[23]_pad  ;
  output \s12_data_o[24]_pad  ;
  output \s12_data_o[25]_pad  ;
  output \s12_data_o[26]_pad  ;
  output \s12_data_o[27]_pad  ;
  output \s12_data_o[28]_pad  ;
  output \s12_data_o[29]_pad  ;
  output \s12_data_o[2]_pad  ;
  output \s12_data_o[30]_pad  ;
  output \s12_data_o[31]_pad  ;
  output \s12_data_o[3]_pad  ;
  output \s12_data_o[4]_pad  ;
  output \s12_data_o[5]_pad  ;
  output \s12_data_o[6]_pad  ;
  output \s12_data_o[7]_pad  ;
  output \s12_data_o[8]_pad  ;
  output \s12_data_o[9]_pad  ;
  output \s12_sel_o[0]_pad  ;
  output \s12_sel_o[1]_pad  ;
  output \s12_sel_o[2]_pad  ;
  output \s12_sel_o[3]_pad  ;
  output \s12_stb_o_pad  ;
  output \s12_we_o_pad  ;
  output \s13_addr_o[0]_pad  ;
  output \s13_addr_o[10]_pad  ;
  output \s13_addr_o[11]_pad  ;
  output \s13_addr_o[12]_pad  ;
  output \s13_addr_o[13]_pad  ;
  output \s13_addr_o[14]_pad  ;
  output \s13_addr_o[15]_pad  ;
  output \s13_addr_o[16]_pad  ;
  output \s13_addr_o[17]_pad  ;
  output \s13_addr_o[18]_pad  ;
  output \s13_addr_o[19]_pad  ;
  output \s13_addr_o[1]_pad  ;
  output \s13_addr_o[20]_pad  ;
  output \s13_addr_o[21]_pad  ;
  output \s13_addr_o[22]_pad  ;
  output \s13_addr_o[23]_pad  ;
  output \s13_addr_o[24]_pad  ;
  output \s13_addr_o[25]_pad  ;
  output \s13_addr_o[26]_pad  ;
  output \s13_addr_o[27]_pad  ;
  output \s13_addr_o[28]_pad  ;
  output \s13_addr_o[29]_pad  ;
  output \s13_addr_o[2]_pad  ;
  output \s13_addr_o[30]_pad  ;
  output \s13_addr_o[31]_pad  ;
  output \s13_addr_o[3]_pad  ;
  output \s13_addr_o[4]_pad  ;
  output \s13_addr_o[5]_pad  ;
  output \s13_addr_o[6]_pad  ;
  output \s13_addr_o[7]_pad  ;
  output \s13_addr_o[8]_pad  ;
  output \s13_addr_o[9]_pad  ;
  output \s13_data_o[0]_pad  ;
  output \s13_data_o[10]_pad  ;
  output \s13_data_o[11]_pad  ;
  output \s13_data_o[12]_pad  ;
  output \s13_data_o[13]_pad  ;
  output \s13_data_o[14]_pad  ;
  output \s13_data_o[15]_pad  ;
  output \s13_data_o[16]_pad  ;
  output \s13_data_o[17]_pad  ;
  output \s13_data_o[18]_pad  ;
  output \s13_data_o[19]_pad  ;
  output \s13_data_o[1]_pad  ;
  output \s13_data_o[20]_pad  ;
  output \s13_data_o[21]_pad  ;
  output \s13_data_o[22]_pad  ;
  output \s13_data_o[23]_pad  ;
  output \s13_data_o[24]_pad  ;
  output \s13_data_o[25]_pad  ;
  output \s13_data_o[26]_pad  ;
  output \s13_data_o[27]_pad  ;
  output \s13_data_o[28]_pad  ;
  output \s13_data_o[29]_pad  ;
  output \s13_data_o[2]_pad  ;
  output \s13_data_o[30]_pad  ;
  output \s13_data_o[31]_pad  ;
  output \s13_data_o[3]_pad  ;
  output \s13_data_o[4]_pad  ;
  output \s13_data_o[5]_pad  ;
  output \s13_data_o[6]_pad  ;
  output \s13_data_o[7]_pad  ;
  output \s13_data_o[8]_pad  ;
  output \s13_data_o[9]_pad  ;
  output \s13_sel_o[0]_pad  ;
  output \s13_sel_o[1]_pad  ;
  output \s13_sel_o[2]_pad  ;
  output \s13_sel_o[3]_pad  ;
  output \s13_stb_o_pad  ;
  output \s13_we_o_pad  ;
  output \s14_addr_o[0]_pad  ;
  output \s14_addr_o[10]_pad  ;
  output \s14_addr_o[11]_pad  ;
  output \s14_addr_o[12]_pad  ;
  output \s14_addr_o[13]_pad  ;
  output \s14_addr_o[14]_pad  ;
  output \s14_addr_o[15]_pad  ;
  output \s14_addr_o[16]_pad  ;
  output \s14_addr_o[17]_pad  ;
  output \s14_addr_o[18]_pad  ;
  output \s14_addr_o[19]_pad  ;
  output \s14_addr_o[1]_pad  ;
  output \s14_addr_o[20]_pad  ;
  output \s14_addr_o[21]_pad  ;
  output \s14_addr_o[22]_pad  ;
  output \s14_addr_o[23]_pad  ;
  output \s14_addr_o[24]_pad  ;
  output \s14_addr_o[25]_pad  ;
  output \s14_addr_o[26]_pad  ;
  output \s14_addr_o[27]_pad  ;
  output \s14_addr_o[28]_pad  ;
  output \s14_addr_o[29]_pad  ;
  output \s14_addr_o[2]_pad  ;
  output \s14_addr_o[30]_pad  ;
  output \s14_addr_o[31]_pad  ;
  output \s14_addr_o[3]_pad  ;
  output \s14_addr_o[4]_pad  ;
  output \s14_addr_o[5]_pad  ;
  output \s14_addr_o[6]_pad  ;
  output \s14_addr_o[7]_pad  ;
  output \s14_addr_o[8]_pad  ;
  output \s14_addr_o[9]_pad  ;
  output \s14_data_o[0]_pad  ;
  output \s14_data_o[10]_pad  ;
  output \s14_data_o[11]_pad  ;
  output \s14_data_o[12]_pad  ;
  output \s14_data_o[13]_pad  ;
  output \s14_data_o[14]_pad  ;
  output \s14_data_o[15]_pad  ;
  output \s14_data_o[16]_pad  ;
  output \s14_data_o[17]_pad  ;
  output \s14_data_o[18]_pad  ;
  output \s14_data_o[19]_pad  ;
  output \s14_data_o[1]_pad  ;
  output \s14_data_o[20]_pad  ;
  output \s14_data_o[21]_pad  ;
  output \s14_data_o[22]_pad  ;
  output \s14_data_o[23]_pad  ;
  output \s14_data_o[24]_pad  ;
  output \s14_data_o[25]_pad  ;
  output \s14_data_o[26]_pad  ;
  output \s14_data_o[27]_pad  ;
  output \s14_data_o[28]_pad  ;
  output \s14_data_o[29]_pad  ;
  output \s14_data_o[2]_pad  ;
  output \s14_data_o[30]_pad  ;
  output \s14_data_o[31]_pad  ;
  output \s14_data_o[3]_pad  ;
  output \s14_data_o[4]_pad  ;
  output \s14_data_o[5]_pad  ;
  output \s14_data_o[6]_pad  ;
  output \s14_data_o[7]_pad  ;
  output \s14_data_o[8]_pad  ;
  output \s14_data_o[9]_pad  ;
  output \s14_sel_o[0]_pad  ;
  output \s14_sel_o[1]_pad  ;
  output \s14_sel_o[2]_pad  ;
  output \s14_sel_o[3]_pad  ;
  output \s14_stb_o_pad  ;
  output \s14_we_o_pad  ;
  output \s15_addr_o[0]_pad  ;
  output \s15_addr_o[10]_pad  ;
  output \s15_addr_o[11]_pad  ;
  output \s15_addr_o[12]_pad  ;
  output \s15_addr_o[13]_pad  ;
  output \s15_addr_o[14]_pad  ;
  output \s15_addr_o[15]_pad  ;
  output \s15_addr_o[16]_pad  ;
  output \s15_addr_o[17]_pad  ;
  output \s15_addr_o[18]_pad  ;
  output \s15_addr_o[19]_pad  ;
  output \s15_addr_o[1]_pad  ;
  output \s15_addr_o[20]_pad  ;
  output \s15_addr_o[21]_pad  ;
  output \s15_addr_o[22]_pad  ;
  output \s15_addr_o[23]_pad  ;
  output \s15_addr_o[24]_pad  ;
  output \s15_addr_o[25]_pad  ;
  output \s15_addr_o[26]_pad  ;
  output \s15_addr_o[27]_pad  ;
  output \s15_addr_o[28]_pad  ;
  output \s15_addr_o[29]_pad  ;
  output \s15_addr_o[2]_pad  ;
  output \s15_addr_o[30]_pad  ;
  output \s15_addr_o[31]_pad  ;
  output \s15_addr_o[3]_pad  ;
  output \s15_addr_o[4]_pad  ;
  output \s15_addr_o[6]_pad  ;
  output \s15_addr_o[7]_pad  ;
  output \s15_addr_o[8]_pad  ;
  output \s15_addr_o[9]_pad  ;
  output \s15_cyc_o_pad  ;
  output \s15_data_o[0]_pad  ;
  output \s15_data_o[10]_pad  ;
  output \s15_data_o[11]_pad  ;
  output \s15_data_o[12]_pad  ;
  output \s15_data_o[13]_pad  ;
  output \s15_data_o[14]_pad  ;
  output \s15_data_o[15]_pad  ;
  output \s15_data_o[16]_pad  ;
  output \s15_data_o[17]_pad  ;
  output \s15_data_o[18]_pad  ;
  output \s15_data_o[19]_pad  ;
  output \s15_data_o[1]_pad  ;
  output \s15_data_o[20]_pad  ;
  output \s15_data_o[21]_pad  ;
  output \s15_data_o[22]_pad  ;
  output \s15_data_o[23]_pad  ;
  output \s15_data_o[24]_pad  ;
  output \s15_data_o[25]_pad  ;
  output \s15_data_o[26]_pad  ;
  output \s15_data_o[27]_pad  ;
  output \s15_data_o[28]_pad  ;
  output \s15_data_o[29]_pad  ;
  output \s15_data_o[2]_pad  ;
  output \s15_data_o[30]_pad  ;
  output \s15_data_o[31]_pad  ;
  output \s15_data_o[3]_pad  ;
  output \s15_data_o[4]_pad  ;
  output \s15_data_o[5]_pad  ;
  output \s15_data_o[6]_pad  ;
  output \s15_data_o[7]_pad  ;
  output \s15_data_o[8]_pad  ;
  output \s15_data_o[9]_pad  ;
  output \s15_sel_o[0]_pad  ;
  output \s15_sel_o[1]_pad  ;
  output \s15_sel_o[2]_pad  ;
  output \s15_sel_o[3]_pad  ;
  output \s15_stb_o_pad  ;
  output \s15_we_o_pad  ;
  output \s1_addr_o[0]_pad  ;
  output \s1_addr_o[10]_pad  ;
  output \s1_addr_o[11]_pad  ;
  output \s1_addr_o[12]_pad  ;
  output \s1_addr_o[13]_pad  ;
  output \s1_addr_o[14]_pad  ;
  output \s1_addr_o[15]_pad  ;
  output \s1_addr_o[16]_pad  ;
  output \s1_addr_o[17]_pad  ;
  output \s1_addr_o[18]_pad  ;
  output \s1_addr_o[19]_pad  ;
  output \s1_addr_o[1]_pad  ;
  output \s1_addr_o[20]_pad  ;
  output \s1_addr_o[21]_pad  ;
  output \s1_addr_o[22]_pad  ;
  output \s1_addr_o[23]_pad  ;
  output \s1_addr_o[24]_pad  ;
  output \s1_addr_o[25]_pad  ;
  output \s1_addr_o[26]_pad  ;
  output \s1_addr_o[27]_pad  ;
  output \s1_addr_o[28]_pad  ;
  output \s1_addr_o[29]_pad  ;
  output \s1_addr_o[2]_pad  ;
  output \s1_addr_o[30]_pad  ;
  output \s1_addr_o[31]_pad  ;
  output \s1_addr_o[3]_pad  ;
  output \s1_addr_o[4]_pad  ;
  output \s1_addr_o[5]_pad  ;
  output \s1_addr_o[6]_pad  ;
  output \s1_addr_o[7]_pad  ;
  output \s1_addr_o[8]_pad  ;
  output \s1_addr_o[9]_pad  ;
  output \s1_data_o[0]_pad  ;
  output \s1_data_o[10]_pad  ;
  output \s1_data_o[11]_pad  ;
  output \s1_data_o[12]_pad  ;
  output \s1_data_o[13]_pad  ;
  output \s1_data_o[14]_pad  ;
  output \s1_data_o[15]_pad  ;
  output \s1_data_o[16]_pad  ;
  output \s1_data_o[17]_pad  ;
  output \s1_data_o[18]_pad  ;
  output \s1_data_o[19]_pad  ;
  output \s1_data_o[1]_pad  ;
  output \s1_data_o[20]_pad  ;
  output \s1_data_o[21]_pad  ;
  output \s1_data_o[22]_pad  ;
  output \s1_data_o[23]_pad  ;
  output \s1_data_o[24]_pad  ;
  output \s1_data_o[25]_pad  ;
  output \s1_data_o[26]_pad  ;
  output \s1_data_o[27]_pad  ;
  output \s1_data_o[28]_pad  ;
  output \s1_data_o[29]_pad  ;
  output \s1_data_o[2]_pad  ;
  output \s1_data_o[30]_pad  ;
  output \s1_data_o[31]_pad  ;
  output \s1_data_o[3]_pad  ;
  output \s1_data_o[4]_pad  ;
  output \s1_data_o[5]_pad  ;
  output \s1_data_o[6]_pad  ;
  output \s1_data_o[7]_pad  ;
  output \s1_data_o[8]_pad  ;
  output \s1_data_o[9]_pad  ;
  output \s1_sel_o[0]_pad  ;
  output \s1_sel_o[1]_pad  ;
  output \s1_sel_o[2]_pad  ;
  output \s1_sel_o[3]_pad  ;
  output \s1_stb_o_pad  ;
  output \s1_we_o_pad  ;
  output \s2_addr_o[0]_pad  ;
  output \s2_addr_o[10]_pad  ;
  output \s2_addr_o[11]_pad  ;
  output \s2_addr_o[12]_pad  ;
  output \s2_addr_o[13]_pad  ;
  output \s2_addr_o[14]_pad  ;
  output \s2_addr_o[15]_pad  ;
  output \s2_addr_o[16]_pad  ;
  output \s2_addr_o[17]_pad  ;
  output \s2_addr_o[18]_pad  ;
  output \s2_addr_o[19]_pad  ;
  output \s2_addr_o[1]_pad  ;
  output \s2_addr_o[20]_pad  ;
  output \s2_addr_o[21]_pad  ;
  output \s2_addr_o[22]_pad  ;
  output \s2_addr_o[23]_pad  ;
  output \s2_addr_o[24]_pad  ;
  output \s2_addr_o[25]_pad  ;
  output \s2_addr_o[26]_pad  ;
  output \s2_addr_o[27]_pad  ;
  output \s2_addr_o[28]_pad  ;
  output \s2_addr_o[29]_pad  ;
  output \s2_addr_o[2]_pad  ;
  output \s2_addr_o[30]_pad  ;
  output \s2_addr_o[31]_pad  ;
  output \s2_addr_o[3]_pad  ;
  output \s2_addr_o[4]_pad  ;
  output \s2_addr_o[5]_pad  ;
  output \s2_addr_o[6]_pad  ;
  output \s2_addr_o[7]_pad  ;
  output \s2_addr_o[8]_pad  ;
  output \s2_addr_o[9]_pad  ;
  output \s2_data_o[0]_pad  ;
  output \s2_data_o[10]_pad  ;
  output \s2_data_o[11]_pad  ;
  output \s2_data_o[12]_pad  ;
  output \s2_data_o[13]_pad  ;
  output \s2_data_o[14]_pad  ;
  output \s2_data_o[15]_pad  ;
  output \s2_data_o[16]_pad  ;
  output \s2_data_o[17]_pad  ;
  output \s2_data_o[18]_pad  ;
  output \s2_data_o[19]_pad  ;
  output \s2_data_o[1]_pad  ;
  output \s2_data_o[20]_pad  ;
  output \s2_data_o[21]_pad  ;
  output \s2_data_o[22]_pad  ;
  output \s2_data_o[23]_pad  ;
  output \s2_data_o[24]_pad  ;
  output \s2_data_o[25]_pad  ;
  output \s2_data_o[26]_pad  ;
  output \s2_data_o[27]_pad  ;
  output \s2_data_o[28]_pad  ;
  output \s2_data_o[29]_pad  ;
  output \s2_data_o[2]_pad  ;
  output \s2_data_o[30]_pad  ;
  output \s2_data_o[31]_pad  ;
  output \s2_data_o[3]_pad  ;
  output \s2_data_o[4]_pad  ;
  output \s2_data_o[5]_pad  ;
  output \s2_data_o[6]_pad  ;
  output \s2_data_o[7]_pad  ;
  output \s2_data_o[8]_pad  ;
  output \s2_data_o[9]_pad  ;
  output \s2_sel_o[0]_pad  ;
  output \s2_sel_o[1]_pad  ;
  output \s2_sel_o[2]_pad  ;
  output \s2_sel_o[3]_pad  ;
  output \s2_stb_o_pad  ;
  output \s2_we_o_pad  ;
  output \s3_addr_o[0]_pad  ;
  output \s3_addr_o[10]_pad  ;
  output \s3_addr_o[11]_pad  ;
  output \s3_addr_o[12]_pad  ;
  output \s3_addr_o[13]_pad  ;
  output \s3_addr_o[14]_pad  ;
  output \s3_addr_o[15]_pad  ;
  output \s3_addr_o[16]_pad  ;
  output \s3_addr_o[17]_pad  ;
  output \s3_addr_o[18]_pad  ;
  output \s3_addr_o[19]_pad  ;
  output \s3_addr_o[1]_pad  ;
  output \s3_addr_o[20]_pad  ;
  output \s3_addr_o[21]_pad  ;
  output \s3_addr_o[22]_pad  ;
  output \s3_addr_o[23]_pad  ;
  output \s3_addr_o[24]_pad  ;
  output \s3_addr_o[25]_pad  ;
  output \s3_addr_o[26]_pad  ;
  output \s3_addr_o[27]_pad  ;
  output \s3_addr_o[28]_pad  ;
  output \s3_addr_o[29]_pad  ;
  output \s3_addr_o[2]_pad  ;
  output \s3_addr_o[30]_pad  ;
  output \s3_addr_o[31]_pad  ;
  output \s3_addr_o[3]_pad  ;
  output \s3_addr_o[4]_pad  ;
  output \s3_addr_o[5]_pad  ;
  output \s3_addr_o[6]_pad  ;
  output \s3_addr_o[7]_pad  ;
  output \s3_addr_o[8]_pad  ;
  output \s3_addr_o[9]_pad  ;
  output \s3_data_o[0]_pad  ;
  output \s3_data_o[10]_pad  ;
  output \s3_data_o[11]_pad  ;
  output \s3_data_o[12]_pad  ;
  output \s3_data_o[13]_pad  ;
  output \s3_data_o[14]_pad  ;
  output \s3_data_o[15]_pad  ;
  output \s3_data_o[16]_pad  ;
  output \s3_data_o[17]_pad  ;
  output \s3_data_o[18]_pad  ;
  output \s3_data_o[19]_pad  ;
  output \s3_data_o[1]_pad  ;
  output \s3_data_o[20]_pad  ;
  output \s3_data_o[21]_pad  ;
  output \s3_data_o[22]_pad  ;
  output \s3_data_o[23]_pad  ;
  output \s3_data_o[24]_pad  ;
  output \s3_data_o[25]_pad  ;
  output \s3_data_o[26]_pad  ;
  output \s3_data_o[27]_pad  ;
  output \s3_data_o[28]_pad  ;
  output \s3_data_o[29]_pad  ;
  output \s3_data_o[2]_pad  ;
  output \s3_data_o[30]_pad  ;
  output \s3_data_o[31]_pad  ;
  output \s3_data_o[3]_pad  ;
  output \s3_data_o[4]_pad  ;
  output \s3_data_o[5]_pad  ;
  output \s3_data_o[6]_pad  ;
  output \s3_data_o[7]_pad  ;
  output \s3_data_o[8]_pad  ;
  output \s3_data_o[9]_pad  ;
  output \s3_sel_o[0]_pad  ;
  output \s3_sel_o[1]_pad  ;
  output \s3_sel_o[2]_pad  ;
  output \s3_sel_o[3]_pad  ;
  output \s3_stb_o_pad  ;
  output \s3_we_o_pad  ;
  output \s4_addr_o[0]_pad  ;
  output \s4_addr_o[10]_pad  ;
  output \s4_addr_o[11]_pad  ;
  output \s4_addr_o[12]_pad  ;
  output \s4_addr_o[13]_pad  ;
  output \s4_addr_o[14]_pad  ;
  output \s4_addr_o[15]_pad  ;
  output \s4_addr_o[16]_pad  ;
  output \s4_addr_o[17]_pad  ;
  output \s4_addr_o[18]_pad  ;
  output \s4_addr_o[19]_pad  ;
  output \s4_addr_o[1]_pad  ;
  output \s4_addr_o[20]_pad  ;
  output \s4_addr_o[21]_pad  ;
  output \s4_addr_o[22]_pad  ;
  output \s4_addr_o[23]_pad  ;
  output \s4_addr_o[24]_pad  ;
  output \s4_addr_o[25]_pad  ;
  output \s4_addr_o[26]_pad  ;
  output \s4_addr_o[27]_pad  ;
  output \s4_addr_o[28]_pad  ;
  output \s4_addr_o[29]_pad  ;
  output \s4_addr_o[2]_pad  ;
  output \s4_addr_o[30]_pad  ;
  output \s4_addr_o[31]_pad  ;
  output \s4_addr_o[3]_pad  ;
  output \s4_addr_o[4]_pad  ;
  output \s4_addr_o[5]_pad  ;
  output \s4_addr_o[6]_pad  ;
  output \s4_addr_o[7]_pad  ;
  output \s4_addr_o[8]_pad  ;
  output \s4_addr_o[9]_pad  ;
  output \s4_data_o[0]_pad  ;
  output \s4_data_o[10]_pad  ;
  output \s4_data_o[11]_pad  ;
  output \s4_data_o[12]_pad  ;
  output \s4_data_o[13]_pad  ;
  output \s4_data_o[14]_pad  ;
  output \s4_data_o[15]_pad  ;
  output \s4_data_o[16]_pad  ;
  output \s4_data_o[17]_pad  ;
  output \s4_data_o[18]_pad  ;
  output \s4_data_o[19]_pad  ;
  output \s4_data_o[1]_pad  ;
  output \s4_data_o[20]_pad  ;
  output \s4_data_o[21]_pad  ;
  output \s4_data_o[22]_pad  ;
  output \s4_data_o[23]_pad  ;
  output \s4_data_o[24]_pad  ;
  output \s4_data_o[25]_pad  ;
  output \s4_data_o[26]_pad  ;
  output \s4_data_o[27]_pad  ;
  output \s4_data_o[28]_pad  ;
  output \s4_data_o[29]_pad  ;
  output \s4_data_o[2]_pad  ;
  output \s4_data_o[30]_pad  ;
  output \s4_data_o[31]_pad  ;
  output \s4_data_o[3]_pad  ;
  output \s4_data_o[4]_pad  ;
  output \s4_data_o[5]_pad  ;
  output \s4_data_o[6]_pad  ;
  output \s4_data_o[7]_pad  ;
  output \s4_data_o[8]_pad  ;
  output \s4_data_o[9]_pad  ;
  output \s4_sel_o[0]_pad  ;
  output \s4_sel_o[1]_pad  ;
  output \s4_sel_o[2]_pad  ;
  output \s4_sel_o[3]_pad  ;
  output \s4_stb_o_pad  ;
  output \s4_we_o_pad  ;
  output \s5_addr_o[0]_pad  ;
  output \s5_addr_o[10]_pad  ;
  output \s5_addr_o[11]_pad  ;
  output \s5_addr_o[12]_pad  ;
  output \s5_addr_o[13]_pad  ;
  output \s5_addr_o[14]_pad  ;
  output \s5_addr_o[15]_pad  ;
  output \s5_addr_o[16]_pad  ;
  output \s5_addr_o[17]_pad  ;
  output \s5_addr_o[18]_pad  ;
  output \s5_addr_o[19]_pad  ;
  output \s5_addr_o[1]_pad  ;
  output \s5_addr_o[20]_pad  ;
  output \s5_addr_o[21]_pad  ;
  output \s5_addr_o[22]_pad  ;
  output \s5_addr_o[23]_pad  ;
  output \s5_addr_o[24]_pad  ;
  output \s5_addr_o[25]_pad  ;
  output \s5_addr_o[26]_pad  ;
  output \s5_addr_o[27]_pad  ;
  output \s5_addr_o[28]_pad  ;
  output \s5_addr_o[29]_pad  ;
  output \s5_addr_o[2]_pad  ;
  output \s5_addr_o[30]_pad  ;
  output \s5_addr_o[31]_pad  ;
  output \s5_addr_o[3]_pad  ;
  output \s5_addr_o[4]_pad  ;
  output \s5_addr_o[5]_pad  ;
  output \s5_addr_o[6]_pad  ;
  output \s5_addr_o[7]_pad  ;
  output \s5_addr_o[8]_pad  ;
  output \s5_addr_o[9]_pad  ;
  output \s5_data_o[0]_pad  ;
  output \s5_data_o[10]_pad  ;
  output \s5_data_o[11]_pad  ;
  output \s5_data_o[12]_pad  ;
  output \s5_data_o[13]_pad  ;
  output \s5_data_o[14]_pad  ;
  output \s5_data_o[15]_pad  ;
  output \s5_data_o[16]_pad  ;
  output \s5_data_o[17]_pad  ;
  output \s5_data_o[18]_pad  ;
  output \s5_data_o[19]_pad  ;
  output \s5_data_o[1]_pad  ;
  output \s5_data_o[20]_pad  ;
  output \s5_data_o[21]_pad  ;
  output \s5_data_o[22]_pad  ;
  output \s5_data_o[23]_pad  ;
  output \s5_data_o[24]_pad  ;
  output \s5_data_o[25]_pad  ;
  output \s5_data_o[26]_pad  ;
  output \s5_data_o[27]_pad  ;
  output \s5_data_o[28]_pad  ;
  output \s5_data_o[29]_pad  ;
  output \s5_data_o[2]_pad  ;
  output \s5_data_o[30]_pad  ;
  output \s5_data_o[31]_pad  ;
  output \s5_data_o[3]_pad  ;
  output \s5_data_o[4]_pad  ;
  output \s5_data_o[5]_pad  ;
  output \s5_data_o[6]_pad  ;
  output \s5_data_o[7]_pad  ;
  output \s5_data_o[8]_pad  ;
  output \s5_data_o[9]_pad  ;
  output \s5_sel_o[0]_pad  ;
  output \s5_sel_o[1]_pad  ;
  output \s5_sel_o[2]_pad  ;
  output \s5_sel_o[3]_pad  ;
  output \s5_stb_o_pad  ;
  output \s5_we_o_pad  ;
  output \s6_addr_o[0]_pad  ;
  output \s6_addr_o[10]_pad  ;
  output \s6_addr_o[11]_pad  ;
  output \s6_addr_o[12]_pad  ;
  output \s6_addr_o[13]_pad  ;
  output \s6_addr_o[14]_pad  ;
  output \s6_addr_o[15]_pad  ;
  output \s6_addr_o[16]_pad  ;
  output \s6_addr_o[17]_pad  ;
  output \s6_addr_o[18]_pad  ;
  output \s6_addr_o[19]_pad  ;
  output \s6_addr_o[1]_pad  ;
  output \s6_addr_o[20]_pad  ;
  output \s6_addr_o[21]_pad  ;
  output \s6_addr_o[22]_pad  ;
  output \s6_addr_o[23]_pad  ;
  output \s6_addr_o[24]_pad  ;
  output \s6_addr_o[25]_pad  ;
  output \s6_addr_o[26]_pad  ;
  output \s6_addr_o[27]_pad  ;
  output \s6_addr_o[28]_pad  ;
  output \s6_addr_o[29]_pad  ;
  output \s6_addr_o[2]_pad  ;
  output \s6_addr_o[30]_pad  ;
  output \s6_addr_o[31]_pad  ;
  output \s6_addr_o[3]_pad  ;
  output \s6_addr_o[4]_pad  ;
  output \s6_addr_o[5]_pad  ;
  output \s6_addr_o[6]_pad  ;
  output \s6_addr_o[7]_pad  ;
  output \s6_addr_o[8]_pad  ;
  output \s6_addr_o[9]_pad  ;
  output \s6_data_o[0]_pad  ;
  output \s6_data_o[10]_pad  ;
  output \s6_data_o[11]_pad  ;
  output \s6_data_o[12]_pad  ;
  output \s6_data_o[13]_pad  ;
  output \s6_data_o[14]_pad  ;
  output \s6_data_o[15]_pad  ;
  output \s6_data_o[16]_pad  ;
  output \s6_data_o[17]_pad  ;
  output \s6_data_o[18]_pad  ;
  output \s6_data_o[19]_pad  ;
  output \s6_data_o[1]_pad  ;
  output \s6_data_o[20]_pad  ;
  output \s6_data_o[21]_pad  ;
  output \s6_data_o[22]_pad  ;
  output \s6_data_o[23]_pad  ;
  output \s6_data_o[24]_pad  ;
  output \s6_data_o[25]_pad  ;
  output \s6_data_o[26]_pad  ;
  output \s6_data_o[27]_pad  ;
  output \s6_data_o[28]_pad  ;
  output \s6_data_o[29]_pad  ;
  output \s6_data_o[2]_pad  ;
  output \s6_data_o[30]_pad  ;
  output \s6_data_o[31]_pad  ;
  output \s6_data_o[3]_pad  ;
  output \s6_data_o[4]_pad  ;
  output \s6_data_o[5]_pad  ;
  output \s6_data_o[6]_pad  ;
  output \s6_data_o[7]_pad  ;
  output \s6_data_o[8]_pad  ;
  output \s6_data_o[9]_pad  ;
  output \s6_sel_o[0]_pad  ;
  output \s6_sel_o[1]_pad  ;
  output \s6_sel_o[2]_pad  ;
  output \s6_sel_o[3]_pad  ;
  output \s6_stb_o_pad  ;
  output \s6_we_o_pad  ;
  output \s7_addr_o[0]_pad  ;
  output \s7_addr_o[10]_pad  ;
  output \s7_addr_o[11]_pad  ;
  output \s7_addr_o[12]_pad  ;
  output \s7_addr_o[13]_pad  ;
  output \s7_addr_o[14]_pad  ;
  output \s7_addr_o[15]_pad  ;
  output \s7_addr_o[16]_pad  ;
  output \s7_addr_o[17]_pad  ;
  output \s7_addr_o[18]_pad  ;
  output \s7_addr_o[19]_pad  ;
  output \s7_addr_o[1]_pad  ;
  output \s7_addr_o[20]_pad  ;
  output \s7_addr_o[21]_pad  ;
  output \s7_addr_o[22]_pad  ;
  output \s7_addr_o[23]_pad  ;
  output \s7_addr_o[24]_pad  ;
  output \s7_addr_o[25]_pad  ;
  output \s7_addr_o[26]_pad  ;
  output \s7_addr_o[27]_pad  ;
  output \s7_addr_o[28]_pad  ;
  output \s7_addr_o[29]_pad  ;
  output \s7_addr_o[2]_pad  ;
  output \s7_addr_o[30]_pad  ;
  output \s7_addr_o[31]_pad  ;
  output \s7_addr_o[3]_pad  ;
  output \s7_addr_o[4]_pad  ;
  output \s7_addr_o[5]_pad  ;
  output \s7_addr_o[6]_pad  ;
  output \s7_addr_o[7]_pad  ;
  output \s7_addr_o[8]_pad  ;
  output \s7_addr_o[9]_pad  ;
  output \s7_data_o[0]_pad  ;
  output \s7_data_o[10]_pad  ;
  output \s7_data_o[11]_pad  ;
  output \s7_data_o[12]_pad  ;
  output \s7_data_o[13]_pad  ;
  output \s7_data_o[14]_pad  ;
  output \s7_data_o[15]_pad  ;
  output \s7_data_o[16]_pad  ;
  output \s7_data_o[17]_pad  ;
  output \s7_data_o[18]_pad  ;
  output \s7_data_o[19]_pad  ;
  output \s7_data_o[1]_pad  ;
  output \s7_data_o[20]_pad  ;
  output \s7_data_o[21]_pad  ;
  output \s7_data_o[22]_pad  ;
  output \s7_data_o[23]_pad  ;
  output \s7_data_o[24]_pad  ;
  output \s7_data_o[25]_pad  ;
  output \s7_data_o[26]_pad  ;
  output \s7_data_o[27]_pad  ;
  output \s7_data_o[28]_pad  ;
  output \s7_data_o[29]_pad  ;
  output \s7_data_o[2]_pad  ;
  output \s7_data_o[30]_pad  ;
  output \s7_data_o[31]_pad  ;
  output \s7_data_o[3]_pad  ;
  output \s7_data_o[4]_pad  ;
  output \s7_data_o[5]_pad  ;
  output \s7_data_o[6]_pad  ;
  output \s7_data_o[7]_pad  ;
  output \s7_data_o[8]_pad  ;
  output \s7_data_o[9]_pad  ;
  output \s7_sel_o[0]_pad  ;
  output \s7_sel_o[1]_pad  ;
  output \s7_sel_o[2]_pad  ;
  output \s7_sel_o[3]_pad  ;
  output \s7_stb_o_pad  ;
  output \s7_we_o_pad  ;
  output \s8_addr_o[0]_pad  ;
  output \s8_addr_o[10]_pad  ;
  output \s8_addr_o[11]_pad  ;
  output \s8_addr_o[12]_pad  ;
  output \s8_addr_o[13]_pad  ;
  output \s8_addr_o[14]_pad  ;
  output \s8_addr_o[15]_pad  ;
  output \s8_addr_o[16]_pad  ;
  output \s8_addr_o[17]_pad  ;
  output \s8_addr_o[18]_pad  ;
  output \s8_addr_o[19]_pad  ;
  output \s8_addr_o[1]_pad  ;
  output \s8_addr_o[20]_pad  ;
  output \s8_addr_o[21]_pad  ;
  output \s8_addr_o[22]_pad  ;
  output \s8_addr_o[23]_pad  ;
  output \s8_addr_o[24]_pad  ;
  output \s8_addr_o[25]_pad  ;
  output \s8_addr_o[26]_pad  ;
  output \s8_addr_o[27]_pad  ;
  output \s8_addr_o[28]_pad  ;
  output \s8_addr_o[29]_pad  ;
  output \s8_addr_o[2]_pad  ;
  output \s8_addr_o[30]_pad  ;
  output \s8_addr_o[31]_pad  ;
  output \s8_addr_o[3]_pad  ;
  output \s8_addr_o[4]_pad  ;
  output \s8_addr_o[5]_pad  ;
  output \s8_addr_o[6]_pad  ;
  output \s8_addr_o[7]_pad  ;
  output \s8_addr_o[8]_pad  ;
  output \s8_addr_o[9]_pad  ;
  output \s8_data_o[0]_pad  ;
  output \s8_data_o[10]_pad  ;
  output \s8_data_o[11]_pad  ;
  output \s8_data_o[12]_pad  ;
  output \s8_data_o[13]_pad  ;
  output \s8_data_o[14]_pad  ;
  output \s8_data_o[15]_pad  ;
  output \s8_data_o[16]_pad  ;
  output \s8_data_o[17]_pad  ;
  output \s8_data_o[18]_pad  ;
  output \s8_data_o[19]_pad  ;
  output \s8_data_o[1]_pad  ;
  output \s8_data_o[20]_pad  ;
  output \s8_data_o[21]_pad  ;
  output \s8_data_o[22]_pad  ;
  output \s8_data_o[23]_pad  ;
  output \s8_data_o[24]_pad  ;
  output \s8_data_o[25]_pad  ;
  output \s8_data_o[26]_pad  ;
  output \s8_data_o[27]_pad  ;
  output \s8_data_o[28]_pad  ;
  output \s8_data_o[29]_pad  ;
  output \s8_data_o[2]_pad  ;
  output \s8_data_o[30]_pad  ;
  output \s8_data_o[31]_pad  ;
  output \s8_data_o[3]_pad  ;
  output \s8_data_o[4]_pad  ;
  output \s8_data_o[5]_pad  ;
  output \s8_data_o[6]_pad  ;
  output \s8_data_o[7]_pad  ;
  output \s8_data_o[8]_pad  ;
  output \s8_data_o[9]_pad  ;
  output \s8_sel_o[0]_pad  ;
  output \s8_sel_o[1]_pad  ;
  output \s8_sel_o[2]_pad  ;
  output \s8_sel_o[3]_pad  ;
  output \s8_stb_o_pad  ;
  output \s8_we_o_pad  ;
  output \s9_addr_o[0]_pad  ;
  output \s9_addr_o[10]_pad  ;
  output \s9_addr_o[11]_pad  ;
  output \s9_addr_o[12]_pad  ;
  output \s9_addr_o[13]_pad  ;
  output \s9_addr_o[14]_pad  ;
  output \s9_addr_o[15]_pad  ;
  output \s9_addr_o[16]_pad  ;
  output \s9_addr_o[17]_pad  ;
  output \s9_addr_o[18]_pad  ;
  output \s9_addr_o[19]_pad  ;
  output \s9_addr_o[1]_pad  ;
  output \s9_addr_o[20]_pad  ;
  output \s9_addr_o[21]_pad  ;
  output \s9_addr_o[22]_pad  ;
  output \s9_addr_o[23]_pad  ;
  output \s9_addr_o[24]_pad  ;
  output \s9_addr_o[25]_pad  ;
  output \s9_addr_o[26]_pad  ;
  output \s9_addr_o[27]_pad  ;
  output \s9_addr_o[28]_pad  ;
  output \s9_addr_o[29]_pad  ;
  output \s9_addr_o[2]_pad  ;
  output \s9_addr_o[30]_pad  ;
  output \s9_addr_o[31]_pad  ;
  output \s9_addr_o[3]_pad  ;
  output \s9_addr_o[4]_pad  ;
  output \s9_addr_o[5]_pad  ;
  output \s9_addr_o[6]_pad  ;
  output \s9_addr_o[7]_pad  ;
  output \s9_addr_o[8]_pad  ;
  output \s9_addr_o[9]_pad  ;
  output \s9_data_o[0]_pad  ;
  output \s9_data_o[10]_pad  ;
  output \s9_data_o[11]_pad  ;
  output \s9_data_o[12]_pad  ;
  output \s9_data_o[13]_pad  ;
  output \s9_data_o[14]_pad  ;
  output \s9_data_o[15]_pad  ;
  output \s9_data_o[16]_pad  ;
  output \s9_data_o[17]_pad  ;
  output \s9_data_o[18]_pad  ;
  output \s9_data_o[19]_pad  ;
  output \s9_data_o[1]_pad  ;
  output \s9_data_o[20]_pad  ;
  output \s9_data_o[21]_pad  ;
  output \s9_data_o[22]_pad  ;
  output \s9_data_o[23]_pad  ;
  output \s9_data_o[24]_pad  ;
  output \s9_data_o[25]_pad  ;
  output \s9_data_o[26]_pad  ;
  output \s9_data_o[27]_pad  ;
  output \s9_data_o[28]_pad  ;
  output \s9_data_o[29]_pad  ;
  output \s9_data_o[2]_pad  ;
  output \s9_data_o[30]_pad  ;
  output \s9_data_o[31]_pad  ;
  output \s9_data_o[3]_pad  ;
  output \s9_data_o[4]_pad  ;
  output \s9_data_o[5]_pad  ;
  output \s9_data_o[6]_pad  ;
  output \s9_data_o[7]_pad  ;
  output \s9_data_o[8]_pad  ;
  output \s9_data_o[9]_pad  ;
  output \s9_sel_o[0]_pad  ;
  output \s9_sel_o[1]_pad  ;
  output \s9_sel_o[2]_pad  ;
  output \s9_sel_o[3]_pad  ;
  output \s9_stb_o_pad  ;
  output \s9_we_o_pad  ;
  wire n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 ;
  assign n1900 = \s15_msel_pri_out_reg[0]/NET0131  & ~\s15_msel_pri_out_reg[1]/NET0131  ;
  assign n1901 = \s15_msel_arb1_state_reg[2]/NET0131  & n1900 ;
  assign n1902 = ~\s15_msel_pri_out_reg[0]/NET0131  & \s15_msel_pri_out_reg[1]/NET0131  ;
  assign n1903 = \s15_msel_arb2_state_reg[2]/NET0131  & n1902 ;
  assign n1904 = ~n1901 & ~n1903 ;
  assign n1905 = ~\s15_msel_pri_out_reg[0]/NET0131  & ~\s15_msel_pri_out_reg[1]/NET0131  ;
  assign n1906 = \s15_msel_arb0_state_reg[2]/NET0131  & n1905 ;
  assign n1907 = \s15_msel_pri_out_reg[0]/NET0131  & \s15_msel_pri_out_reg[1]/NET0131  ;
  assign n1908 = \s15_msel_arb3_state_reg[2]/NET0131  & n1907 ;
  assign n1909 = ~n1906 & ~n1908 ;
  assign n1910 = n1904 & n1909 ;
  assign n1911 = \s15_msel_arb1_state_reg[0]/NET0131  & n1900 ;
  assign n1912 = \s15_msel_arb0_state_reg[0]/NET0131  & n1905 ;
  assign n1913 = ~n1911 & ~n1912 ;
  assign n1914 = \s15_msel_arb3_state_reg[0]/NET0131  & n1907 ;
  assign n1915 = \s15_msel_arb2_state_reg[0]/NET0131  & n1902 ;
  assign n1916 = ~n1914 & ~n1915 ;
  assign n1917 = n1913 & n1916 ;
  assign n1918 = ~n1910 & n1917 ;
  assign n1919 = \s15_msel_arb1_state_reg[1]/NET0131  & n1900 ;
  assign n1920 = \s15_msel_arb0_state_reg[1]/NET0131  & n1905 ;
  assign n1921 = ~n1919 & ~n1920 ;
  assign n1922 = \s15_msel_arb2_state_reg[1]/NET0131  & n1902 ;
  assign n1923 = \s15_msel_arb3_state_reg[1]/NET0131  & n1907 ;
  assign n1924 = ~n1922 & ~n1923 ;
  assign n1925 = n1921 & n1924 ;
  assign n1926 = \m4_addr_i[2]_pad  & n1925 ;
  assign n1927 = n1918 & n1926 ;
  assign n1928 = \m6_addr_i[2]_pad  & ~n1925 ;
  assign n1929 = n1918 & n1928 ;
  assign n1930 = ~n1927 & ~n1929 ;
  assign n1931 = n1910 & n1917 ;
  assign n1932 = \m2_addr_i[2]_pad  & ~n1925 ;
  assign n1933 = n1931 & n1932 ;
  assign n1934 = \m0_addr_i[2]_pad  & n1925 ;
  assign n1935 = n1931 & n1934 ;
  assign n1936 = ~n1933 & ~n1935 ;
  assign n1937 = n1930 & n1936 ;
  assign n1938 = ~n1917 & ~n1925 ;
  assign n1939 = \m7_addr_i[2]_pad  & ~n1910 ;
  assign n1940 = n1938 & n1939 ;
  assign n1941 = ~n1917 & n1925 ;
  assign n1942 = \m5_addr_i[2]_pad  & ~n1910 ;
  assign n1943 = n1941 & n1942 ;
  assign n1944 = ~n1940 & ~n1943 ;
  assign n1945 = \m1_addr_i[2]_pad  & n1910 ;
  assign n1946 = n1941 & n1945 ;
  assign n1947 = \m3_addr_i[2]_pad  & n1910 ;
  assign n1948 = n1938 & n1947 ;
  assign n1949 = ~n1946 & ~n1948 ;
  assign n1950 = n1944 & n1949 ;
  assign n1951 = n1937 & n1950 ;
  assign n1952 = \m7_addr_i[3]_pad  & ~n1910 ;
  assign n1953 = n1938 & n1952 ;
  assign n1954 = \m3_addr_i[3]_pad  & n1910 ;
  assign n1955 = n1938 & n1954 ;
  assign n1956 = ~n1953 & ~n1955 ;
  assign n1957 = \m6_addr_i[3]_pad  & ~n1925 ;
  assign n1958 = n1918 & n1957 ;
  assign n1959 = \m5_addr_i[3]_pad  & ~n1910 ;
  assign n1960 = n1941 & n1959 ;
  assign n1961 = ~n1958 & ~n1960 ;
  assign n1962 = n1956 & n1961 ;
  assign n1963 = \m4_addr_i[3]_pad  & n1925 ;
  assign n1964 = n1918 & n1963 ;
  assign n1965 = \m0_addr_i[3]_pad  & n1925 ;
  assign n1966 = n1931 & n1965 ;
  assign n1967 = ~n1964 & ~n1966 ;
  assign n1968 = \m1_addr_i[3]_pad  & n1910 ;
  assign n1969 = n1941 & n1968 ;
  assign n1970 = \m2_addr_i[3]_pad  & ~n1925 ;
  assign n1971 = n1931 & n1970 ;
  assign n1972 = ~n1969 & ~n1971 ;
  assign n1973 = n1967 & n1972 ;
  assign n1974 = n1962 & n1973 ;
  assign n1975 = ~n1951 & n1974 ;
  assign n1976 = \m6_addr_i[5]_pad  & ~n1925 ;
  assign n1977 = n1918 & n1976 ;
  assign n1978 = \m7_addr_i[5]_pad  & ~n1910 ;
  assign n1979 = n1938 & n1978 ;
  assign n1980 = ~n1977 & ~n1979 ;
  assign n1981 = \m4_addr_i[5]_pad  & n1925 ;
  assign n1982 = n1918 & n1981 ;
  assign n1983 = \m5_addr_i[5]_pad  & ~n1910 ;
  assign n1984 = n1941 & n1983 ;
  assign n1985 = ~n1982 & ~n1984 ;
  assign n1986 = n1980 & n1985 ;
  assign n1987 = \m0_addr_i[5]_pad  & n1925 ;
  assign n1988 = n1931 & n1987 ;
  assign n1989 = \m1_addr_i[5]_pad  & n1910 ;
  assign n1990 = n1941 & n1989 ;
  assign n1991 = ~n1988 & ~n1990 ;
  assign n1992 = \m2_addr_i[5]_pad  & ~n1925 ;
  assign n1993 = n1931 & n1992 ;
  assign n1994 = \m3_addr_i[5]_pad  & n1910 ;
  assign n1995 = n1938 & n1994 ;
  assign n1996 = ~n1993 & ~n1995 ;
  assign n1997 = n1991 & n1996 ;
  assign n1998 = n1986 & n1997 ;
  assign n1999 = \m1_addr_i[4]_pad  & n1910 ;
  assign n2000 = n1941 & n1999 ;
  assign n2001 = \m0_addr_i[4]_pad  & n1925 ;
  assign n2002 = n1931 & n2001 ;
  assign n2003 = ~n2000 & ~n2002 ;
  assign n2004 = \m4_addr_i[4]_pad  & n1925 ;
  assign n2005 = n1918 & n2004 ;
  assign n2006 = \m5_addr_i[4]_pad  & ~n1910 ;
  assign n2007 = n1941 & n2006 ;
  assign n2008 = ~n2005 & ~n2007 ;
  assign n2009 = n2003 & n2008 ;
  assign n2010 = \m6_addr_i[4]_pad  & ~n1925 ;
  assign n2011 = n1918 & n2010 ;
  assign n2012 = \m7_addr_i[4]_pad  & ~n1910 ;
  assign n2013 = n1938 & n2012 ;
  assign n2014 = ~n2011 & ~n2013 ;
  assign n2015 = \m3_addr_i[4]_pad  & n1910 ;
  assign n2016 = n1938 & n2015 ;
  assign n2017 = \m2_addr_i[4]_pad  & ~n1925 ;
  assign n2018 = n1931 & n2017 ;
  assign n2019 = ~n2016 & ~n2018 ;
  assign n2020 = n2014 & n2019 ;
  assign n2021 = n2009 & n2020 ;
  assign n2022 = n1998 & ~n2021 ;
  assign n2023 = n1975 & n2022 ;
  assign n2024 = \rf_conf5_reg[11]/NET0131  & n2023 ;
  assign n2025 = n1998 & n2021 ;
  assign n2026 = ~n1951 & ~n1974 ;
  assign n2027 = n2025 & n2026 ;
  assign n2028 = \rf_conf3_reg[11]/NET0131  & n2027 ;
  assign n2029 = ~n2024 & ~n2028 ;
  assign n2030 = n1951 & n1974 ;
  assign n2031 = ~n1998 & ~n2021 ;
  assign n2032 = n2030 & n2031 ;
  assign n2033 = \rf_conf12_reg[11]/NET0131  & n2032 ;
  assign n2034 = n1951 & ~n1974 ;
  assign n2035 = n2031 & n2034 ;
  assign n2036 = \rf_conf14_reg[11]/NET0131  & n2035 ;
  assign n2037 = ~n2033 & ~n2036 ;
  assign n2038 = n2029 & n2037 ;
  assign n2039 = n2025 & n2034 ;
  assign n2040 = \rf_conf2_reg[11]/NET0131  & n2039 ;
  assign n2041 = n1975 & n2025 ;
  assign n2042 = \rf_conf1_reg[11]/NET0131  & n2041 ;
  assign n2043 = ~n2040 & ~n2042 ;
  assign n2044 = n2025 & n2030 ;
  assign n2045 = \rf_conf0_reg[11]/NET0131  & n2044 ;
  assign n2046 = n2022 & n2030 ;
  assign n2047 = \rf_conf4_reg[11]/NET0131  & n2046 ;
  assign n2048 = ~n2045 & ~n2047 ;
  assign n2049 = n2043 & n2048 ;
  assign n2050 = n2038 & n2049 ;
  assign n2051 = n2022 & n2034 ;
  assign n2052 = \rf_conf6_reg[11]/NET0131  & n2051 ;
  assign n2053 = n2022 & n2026 ;
  assign n2054 = \rf_conf7_reg[11]/NET0131  & n2053 ;
  assign n2055 = ~n2052 & ~n2054 ;
  assign n2056 = ~n1998 & n2021 ;
  assign n2057 = n2030 & n2056 ;
  assign n2058 = \rf_conf8_reg[11]/NET0131  & n2057 ;
  assign n2059 = n2026 & n2056 ;
  assign n2060 = \rf_conf11_reg[11]/NET0131  & n2059 ;
  assign n2061 = ~n2058 & ~n2060 ;
  assign n2062 = n2055 & n2061 ;
  assign n2063 = n1975 & n2056 ;
  assign n2064 = \rf_conf9_reg[11]/NET0131  & n2063 ;
  assign n2065 = n2034 & n2056 ;
  assign n2066 = \rf_conf10_reg[11]/NET0131  & n2065 ;
  assign n2067 = ~n2064 & ~n2066 ;
  assign n2068 = n1975 & n2031 ;
  assign n2069 = \rf_conf13_reg[11]/NET0131  & n2068 ;
  assign n2070 = n2026 & n2031 ;
  assign n2071 = \rf_conf15_reg[11]/NET0131  & n2070 ;
  assign n2072 = ~n2069 & ~n2071 ;
  assign n2073 = n2067 & n2072 ;
  assign n2074 = n2062 & n2073 ;
  assign n2075 = n2050 & n2074 ;
  assign n2076 = \m5_s15_cyc_o_reg/NET0131  & \s15_m5_cyc_r_reg/P0001  ;
  assign n2077 = ~n1910 & n2076 ;
  assign n2078 = n1941 & n2077 ;
  assign n2079 = \m4_s15_cyc_o_reg/NET0131  & \s15_m4_cyc_r_reg/P0001  ;
  assign n2080 = n1925 & n2079 ;
  assign n2081 = n1918 & n2080 ;
  assign n2082 = ~n2078 & ~n2081 ;
  assign n2083 = \m2_s15_cyc_o_reg/NET0131  & \s15_m2_cyc_r_reg/P0001  ;
  assign n2084 = ~n1925 & n2083 ;
  assign n2085 = n1931 & n2084 ;
  assign n2086 = \m3_s15_cyc_o_reg/NET0131  & \s15_m3_cyc_r_reg/P0001  ;
  assign n2087 = n1910 & n2086 ;
  assign n2088 = n1938 & n2087 ;
  assign n2089 = ~n2085 & ~n2088 ;
  assign n2090 = n2082 & n2089 ;
  assign n2091 = \m0_s15_cyc_o_reg/NET0131  & \s15_m0_cyc_r_reg/P0001  ;
  assign n2092 = n1925 & n2091 ;
  assign n2093 = n1931 & n2092 ;
  assign n2094 = \m1_s15_cyc_o_reg/NET0131  & \s15_m1_cyc_r_reg/P0001  ;
  assign n2095 = n1910 & n2094 ;
  assign n2096 = n1941 & n2095 ;
  assign n2097 = ~n2093 & ~n2096 ;
  assign n2098 = \m6_s15_cyc_o_reg/NET0131  & \s15_m6_cyc_r_reg/P0001  ;
  assign n2099 = ~n1925 & n2098 ;
  assign n2100 = n1918 & n2099 ;
  assign n2101 = \m7_s15_cyc_o_reg/NET0131  & \s15_m7_cyc_r_reg/P0001  ;
  assign n2102 = ~n1910 & n2101 ;
  assign n2103 = n1938 & n2102 ;
  assign n2104 = ~n2100 & ~n2103 ;
  assign n2105 = n2097 & n2104 ;
  assign n2106 = n2090 & n2105 ;
  assign n2107 = \m3_addr_i[27]_pad  & n1910 ;
  assign n2108 = n1938 & n2107 ;
  assign n2109 = \m7_addr_i[27]_pad  & ~n1910 ;
  assign n2110 = n1938 & n2109 ;
  assign n2111 = ~n2108 & ~n2110 ;
  assign n2112 = \m4_addr_i[27]_pad  & n1925 ;
  assign n2113 = n1918 & n2112 ;
  assign n2114 = \m1_addr_i[27]_pad  & n1910 ;
  assign n2115 = n1941 & n2114 ;
  assign n2116 = ~n2113 & ~n2115 ;
  assign n2117 = n2111 & n2116 ;
  assign n2118 = \m0_addr_i[27]_pad  & n1925 ;
  assign n2119 = n1931 & n2118 ;
  assign n2120 = \m5_addr_i[27]_pad  & ~n1910 ;
  assign n2121 = n1941 & n2120 ;
  assign n2122 = ~n2119 & ~n2121 ;
  assign n2123 = \m2_addr_i[27]_pad  & ~n1925 ;
  assign n2124 = n1931 & n2123 ;
  assign n2125 = \m6_addr_i[27]_pad  & ~n1925 ;
  assign n2126 = n1918 & n2125 ;
  assign n2127 = ~n2124 & ~n2126 ;
  assign n2128 = n2122 & n2127 ;
  assign n2129 = n2117 & n2128 ;
  assign n2130 = \m2_addr_i[24]_pad  & ~n1925 ;
  assign n2131 = n1931 & n2130 ;
  assign n2132 = \m7_addr_i[24]_pad  & ~n1910 ;
  assign n2133 = n1938 & n2132 ;
  assign n2134 = ~n2131 & ~n2133 ;
  assign n2135 = \m0_addr_i[24]_pad  & n1925 ;
  assign n2136 = n1931 & n2135 ;
  assign n2137 = \m6_addr_i[24]_pad  & ~n1925 ;
  assign n2138 = n1918 & n2137 ;
  assign n2139 = ~n2136 & ~n2138 ;
  assign n2140 = n2134 & n2139 ;
  assign n2141 = \m1_addr_i[24]_pad  & n1910 ;
  assign n2142 = n1941 & n2141 ;
  assign n2143 = \m4_addr_i[24]_pad  & n1925 ;
  assign n2144 = n1918 & n2143 ;
  assign n2145 = ~n2142 & ~n2144 ;
  assign n2146 = \m5_addr_i[24]_pad  & ~n1910 ;
  assign n2147 = n1941 & n2146 ;
  assign n2148 = \m3_addr_i[24]_pad  & n1910 ;
  assign n2149 = n1938 & n2148 ;
  assign n2150 = ~n2147 & ~n2149 ;
  assign n2151 = n2145 & n2150 ;
  assign n2152 = n2140 & n2151 ;
  assign n2153 = ~n2129 & ~n2152 ;
  assign n2154 = ~n2106 & n2153 ;
  assign n2155 = \m1_addr_i[28]_pad  & \m1_addr_i[29]_pad  ;
  assign n2156 = \m1_addr_i[30]_pad  & \m1_addr_i[31]_pad  ;
  assign n2157 = n2155 & n2156 ;
  assign n2158 = \m1_stb_i_pad  & n2157 ;
  assign n2159 = n1910 & n2158 ;
  assign n2160 = n1941 & n2159 ;
  assign n2161 = \m0_addr_i[29]_pad  & \m0_addr_i[31]_pad  ;
  assign n2162 = \m0_addr_i[28]_pad  & \m0_addr_i[30]_pad  ;
  assign n2163 = n2161 & n2162 ;
  assign n2164 = \m0_stb_i_pad  & n2163 ;
  assign n2165 = n1925 & n2164 ;
  assign n2166 = n1931 & n2165 ;
  assign n2167 = ~n2160 & ~n2166 ;
  assign n2168 = \m7_addr_i[30]_pad  & \m7_addr_i[31]_pad  ;
  assign n2169 = \m7_addr_i[28]_pad  & \m7_addr_i[29]_pad  ;
  assign n2170 = n2168 & n2169 ;
  assign n2171 = \m7_stb_i_pad  & n2170 ;
  assign n2172 = ~n1910 & n2171 ;
  assign n2173 = n1938 & n2172 ;
  assign n2174 = \m6_addr_i[28]_pad  & \m6_addr_i[29]_pad  ;
  assign n2175 = \m6_addr_i[30]_pad  & \m6_addr_i[31]_pad  ;
  assign n2176 = n2174 & n2175 ;
  assign n2177 = \m6_stb_i_pad  & n2176 ;
  assign n2178 = ~n1925 & n2177 ;
  assign n2179 = n1918 & n2178 ;
  assign n2180 = ~n2173 & ~n2179 ;
  assign n2181 = n2167 & n2180 ;
  assign n2182 = \m2_addr_i[28]_pad  & \m2_addr_i[29]_pad  ;
  assign n2183 = \m2_addr_i[30]_pad  & \m2_addr_i[31]_pad  ;
  assign n2184 = n2182 & n2183 ;
  assign n2185 = \m2_stb_i_pad  & n2184 ;
  assign n2186 = ~n1925 & n2185 ;
  assign n2187 = n1931 & n2186 ;
  assign n2188 = \m3_addr_i[28]_pad  & \m3_addr_i[29]_pad  ;
  assign n2189 = \m3_addr_i[30]_pad  & \m3_addr_i[31]_pad  ;
  assign n2190 = n2188 & n2189 ;
  assign n2191 = \m3_stb_i_pad  & n2190 ;
  assign n2192 = n1910 & n2191 ;
  assign n2193 = n1938 & n2192 ;
  assign n2194 = ~n2187 & ~n2193 ;
  assign n2195 = \m4_addr_i[28]_pad  & \m4_addr_i[29]_pad  ;
  assign n2196 = \m4_addr_i[30]_pad  & \m4_addr_i[31]_pad  ;
  assign n2197 = n2195 & n2196 ;
  assign n2198 = \m4_stb_i_pad  & n2197 ;
  assign n2199 = n1925 & n2198 ;
  assign n2200 = n1918 & n2199 ;
  assign n2201 = \m5_addr_i[28]_pad  & \m5_addr_i[29]_pad  ;
  assign n2202 = \m5_addr_i[30]_pad  & \m5_addr_i[31]_pad  ;
  assign n2203 = n2201 & n2202 ;
  assign n2204 = \m5_stb_i_pad  & n2203 ;
  assign n2205 = ~n1910 & n2204 ;
  assign n2206 = n1941 & n2205 ;
  assign n2207 = ~n2200 & ~n2206 ;
  assign n2208 = n2194 & n2207 ;
  assign n2209 = n2181 & n2208 ;
  assign n2210 = \m7_addr_i[25]_pad  & ~n1910 ;
  assign n2211 = n1938 & n2210 ;
  assign n2212 = \m5_addr_i[25]_pad  & ~n1910 ;
  assign n2213 = n1941 & n2212 ;
  assign n2214 = ~n2211 & ~n2213 ;
  assign n2215 = \m6_addr_i[25]_pad  & ~n1925 ;
  assign n2216 = n1918 & n2215 ;
  assign n2217 = \m1_addr_i[25]_pad  & n1910 ;
  assign n2218 = n1941 & n2217 ;
  assign n2219 = ~n2216 & ~n2218 ;
  assign n2220 = n2214 & n2219 ;
  assign n2221 = \m3_addr_i[25]_pad  & n1910 ;
  assign n2222 = n1938 & n2221 ;
  assign n2223 = \m4_addr_i[25]_pad  & n1925 ;
  assign n2224 = n1918 & n2223 ;
  assign n2225 = ~n2222 & ~n2224 ;
  assign n2226 = \m0_addr_i[25]_pad  & n1925 ;
  assign n2227 = n1931 & n2226 ;
  assign n2228 = \m2_addr_i[25]_pad  & ~n1925 ;
  assign n2229 = n1931 & n2228 ;
  assign n2230 = ~n2227 & ~n2229 ;
  assign n2231 = n2225 & n2230 ;
  assign n2232 = n2220 & n2231 ;
  assign n2233 = \m1_addr_i[26]_pad  & n1910 ;
  assign n2234 = n1941 & n2233 ;
  assign n2235 = \m2_addr_i[26]_pad  & ~n1925 ;
  assign n2236 = n1931 & n2235 ;
  assign n2237 = ~n2234 & ~n2236 ;
  assign n2238 = \m7_addr_i[26]_pad  & ~n1910 ;
  assign n2239 = n1938 & n2238 ;
  assign n2240 = \m3_addr_i[26]_pad  & n1910 ;
  assign n2241 = n1938 & n2240 ;
  assign n2242 = ~n2239 & ~n2241 ;
  assign n2243 = n2237 & n2242 ;
  assign n2244 = \m6_addr_i[26]_pad  & ~n1925 ;
  assign n2245 = n1918 & n2244 ;
  assign n2246 = \m5_addr_i[26]_pad  & ~n1910 ;
  assign n2247 = n1941 & n2246 ;
  assign n2248 = ~n2245 & ~n2247 ;
  assign n2249 = \m4_addr_i[26]_pad  & n1925 ;
  assign n2250 = n1918 & n2249 ;
  assign n2251 = \m0_addr_i[26]_pad  & n1925 ;
  assign n2252 = n1931 & n2251 ;
  assign n2253 = ~n2250 & ~n2252 ;
  assign n2254 = n2248 & n2253 ;
  assign n2255 = n2243 & n2254 ;
  assign n2256 = ~n2232 & ~n2255 ;
  assign n2257 = ~n2209 & n2256 ;
  assign n2258 = n2154 & n2257 ;
  assign n2259 = ~n2075 & n2258 ;
  assign n2260 = \rf_conf8_reg[0]/NET0131  & n2057 ;
  assign n2261 = \rf_conf11_reg[0]/NET0131  & n2059 ;
  assign n2262 = ~n2260 & ~n2261 ;
  assign n2263 = \rf_conf6_reg[0]/NET0131  & n2051 ;
  assign n2264 = \rf_conf7_reg[0]/NET0131  & n2053 ;
  assign n2265 = ~n2263 & ~n2264 ;
  assign n2266 = n2262 & n2265 ;
  assign n2267 = \rf_conf12_reg[0]/NET0131  & n2032 ;
  assign n2268 = \rf_conf14_reg[0]/NET0131  & n2035 ;
  assign n2269 = ~n2267 & ~n2268 ;
  assign n2270 = \rf_conf5_reg[0]/NET0131  & n2023 ;
  assign n2271 = \rf_conf3_reg[0]/NET0131  & n2027 ;
  assign n2272 = ~n2270 & ~n2271 ;
  assign n2273 = n2269 & n2272 ;
  assign n2274 = n2266 & n2273 ;
  assign n2275 = \rf_conf2_reg[0]/NET0131  & n2039 ;
  assign n2276 = \rf_conf1_reg[0]/NET0131  & n2041 ;
  assign n2277 = ~n2275 & ~n2276 ;
  assign n2278 = \rf_conf15_reg[0]/NET0131  & n2070 ;
  assign n2279 = \rf_conf13_reg[0]/NET0131  & n2068 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = n2277 & n2280 ;
  assign n2282 = \rf_conf10_reg[0]/NET0131  & n2065 ;
  assign n2283 = \rf_conf9_reg[0]/NET0131  & n2063 ;
  assign n2284 = ~n2282 & ~n2283 ;
  assign n2285 = \rf_conf0_reg[0]/NET0131  & n2044 ;
  assign n2286 = \rf_conf4_reg[0]/NET0131  & n2046 ;
  assign n2287 = ~n2285 & ~n2286 ;
  assign n2288 = n2284 & n2287 ;
  assign n2289 = n2281 & n2288 ;
  assign n2290 = n2274 & n2289 ;
  assign n2291 = n2258 & ~n2290 ;
  assign n2292 = \rf_conf12_reg[10]/NET0131  & n2032 ;
  assign n2293 = \rf_conf14_reg[10]/NET0131  & n2035 ;
  assign n2294 = ~n2292 & ~n2293 ;
  assign n2295 = \rf_conf6_reg[10]/NET0131  & n2051 ;
  assign n2296 = \rf_conf7_reg[10]/NET0131  & n2053 ;
  assign n2297 = ~n2295 & ~n2296 ;
  assign n2298 = n2294 & n2297 ;
  assign n2299 = \rf_conf8_reg[10]/NET0131  & n2057 ;
  assign n2300 = \rf_conf11_reg[10]/NET0131  & n2059 ;
  assign n2301 = ~n2299 & ~n2300 ;
  assign n2302 = \rf_conf1_reg[10]/NET0131  & n2041 ;
  assign n2303 = \rf_conf2_reg[10]/NET0131  & n2039 ;
  assign n2304 = ~n2302 & ~n2303 ;
  assign n2305 = n2301 & n2304 ;
  assign n2306 = n2298 & n2305 ;
  assign n2307 = \rf_conf3_reg[10]/NET0131  & n2027 ;
  assign n2308 = \rf_conf5_reg[10]/NET0131  & n2023 ;
  assign n2309 = ~n2307 & ~n2308 ;
  assign n2310 = \rf_conf15_reg[10]/NET0131  & n2070 ;
  assign n2311 = \rf_conf13_reg[10]/NET0131  & n2068 ;
  assign n2312 = ~n2310 & ~n2311 ;
  assign n2313 = n2309 & n2312 ;
  assign n2314 = \rf_conf4_reg[10]/NET0131  & n2046 ;
  assign n2315 = \rf_conf0_reg[10]/NET0131  & n2044 ;
  assign n2316 = ~n2314 & ~n2315 ;
  assign n2317 = \rf_conf9_reg[10]/NET0131  & n2063 ;
  assign n2318 = \rf_conf10_reg[10]/NET0131  & n2065 ;
  assign n2319 = ~n2317 & ~n2318 ;
  assign n2320 = n2316 & n2319 ;
  assign n2321 = n2313 & n2320 ;
  assign n2322 = n2306 & n2321 ;
  assign n2323 = n2258 & ~n2322 ;
  assign n2324 = \rf_conf9_reg[12]/NET0131  & n2063 ;
  assign n2325 = \rf_conf10_reg[12]/NET0131  & n2065 ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2327 = \rf_conf14_reg[12]/NET0131  & n2035 ;
  assign n2328 = \rf_conf12_reg[12]/NET0131  & n2032 ;
  assign n2329 = ~n2327 & ~n2328 ;
  assign n2330 = n2326 & n2329 ;
  assign n2331 = \rf_conf0_reg[12]/NET0131  & n2044 ;
  assign n2332 = \rf_conf4_reg[12]/NET0131  & n2046 ;
  assign n2333 = ~n2331 & ~n2332 ;
  assign n2334 = \rf_conf13_reg[12]/NET0131  & n2068 ;
  assign n2335 = \rf_conf15_reg[12]/NET0131  & n2070 ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = n2333 & n2336 ;
  assign n2338 = n2330 & n2337 ;
  assign n2339 = \rf_conf6_reg[12]/NET0131  & n2051 ;
  assign n2340 = \rf_conf7_reg[12]/NET0131  & n2053 ;
  assign n2341 = ~n2339 & ~n2340 ;
  assign n2342 = \rf_conf8_reg[12]/NET0131  & n2057 ;
  assign n2343 = \rf_conf11_reg[12]/NET0131  & n2059 ;
  assign n2344 = ~n2342 & ~n2343 ;
  assign n2345 = n2341 & n2344 ;
  assign n2346 = \rf_conf5_reg[12]/NET0131  & n2023 ;
  assign n2347 = \rf_conf3_reg[12]/NET0131  & n2027 ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2349 = \rf_conf1_reg[12]/NET0131  & n2041 ;
  assign n2350 = \rf_conf2_reg[12]/NET0131  & n2039 ;
  assign n2351 = ~n2349 & ~n2350 ;
  assign n2352 = n2348 & n2351 ;
  assign n2353 = n2345 & n2352 ;
  assign n2354 = n2338 & n2353 ;
  assign n2355 = n2258 & ~n2354 ;
  assign n2356 = \rf_conf12_reg[13]/NET0131  & n2032 ;
  assign n2357 = \rf_conf14_reg[13]/NET0131  & n2035 ;
  assign n2358 = ~n2356 & ~n2357 ;
  assign n2359 = \rf_conf10_reg[13]/NET0131  & n2065 ;
  assign n2360 = \rf_conf9_reg[13]/NET0131  & n2063 ;
  assign n2361 = ~n2359 & ~n2360 ;
  assign n2362 = n2358 & n2361 ;
  assign n2363 = \rf_conf8_reg[13]/NET0131  & n2057 ;
  assign n2364 = \rf_conf11_reg[13]/NET0131  & n2059 ;
  assign n2365 = ~n2363 & ~n2364 ;
  assign n2366 = \rf_conf1_reg[13]/NET0131  & n2041 ;
  assign n2367 = \rf_conf2_reg[13]/NET0131  & n2039 ;
  assign n2368 = ~n2366 & ~n2367 ;
  assign n2369 = n2365 & n2368 ;
  assign n2370 = n2362 & n2369 ;
  assign n2371 = \rf_conf3_reg[13]/NET0131  & n2027 ;
  assign n2372 = \rf_conf5_reg[13]/NET0131  & n2023 ;
  assign n2373 = ~n2371 & ~n2372 ;
  assign n2374 = \rf_conf6_reg[13]/NET0131  & n2051 ;
  assign n2375 = \rf_conf7_reg[13]/NET0131  & n2053 ;
  assign n2376 = ~n2374 & ~n2375 ;
  assign n2377 = n2373 & n2376 ;
  assign n2378 = \rf_conf13_reg[13]/NET0131  & n2068 ;
  assign n2379 = \rf_conf15_reg[13]/NET0131  & n2070 ;
  assign n2380 = ~n2378 & ~n2379 ;
  assign n2381 = \rf_conf0_reg[13]/NET0131  & n2044 ;
  assign n2382 = \rf_conf4_reg[13]/NET0131  & n2046 ;
  assign n2383 = ~n2381 & ~n2382 ;
  assign n2384 = n2380 & n2383 ;
  assign n2385 = n2377 & n2384 ;
  assign n2386 = n2370 & n2385 ;
  assign n2387 = n2258 & ~n2386 ;
  assign n2388 = \rf_conf6_reg[14]/NET0131  & n2051 ;
  assign n2389 = \rf_conf7_reg[14]/NET0131  & n2053 ;
  assign n2390 = ~n2388 & ~n2389 ;
  assign n2391 = \rf_conf8_reg[14]/NET0131  & n2057 ;
  assign n2392 = \rf_conf11_reg[14]/NET0131  & n2059 ;
  assign n2393 = ~n2391 & ~n2392 ;
  assign n2394 = n2390 & n2393 ;
  assign n2395 = \rf_conf13_reg[14]/NET0131  & n2068 ;
  assign n2396 = \rf_conf15_reg[14]/NET0131  & n2070 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = \rf_conf4_reg[14]/NET0131  & n2046 ;
  assign n2399 = \rf_conf0_reg[14]/NET0131  & n2044 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = n2397 & n2400 ;
  assign n2402 = n2394 & n2401 ;
  assign n2403 = \rf_conf10_reg[14]/NET0131  & n2065 ;
  assign n2404 = \rf_conf9_reg[14]/NET0131  & n2063 ;
  assign n2405 = ~n2403 & ~n2404 ;
  assign n2406 = \rf_conf3_reg[14]/NET0131  & n2027 ;
  assign n2407 = \rf_conf2_reg[14]/NET0131  & n2039 ;
  assign n2408 = ~n2406 & ~n2407 ;
  assign n2409 = n2405 & n2408 ;
  assign n2410 = \rf_conf1_reg[14]/NET0131  & n2041 ;
  assign n2411 = \rf_conf14_reg[14]/NET0131  & n2035 ;
  assign n2412 = ~n2410 & ~n2411 ;
  assign n2413 = \rf_conf12_reg[14]/NET0131  & n2032 ;
  assign n2414 = \rf_conf5_reg[14]/NET0131  & n2023 ;
  assign n2415 = ~n2413 & ~n2414 ;
  assign n2416 = n2412 & n2415 ;
  assign n2417 = n2409 & n2416 ;
  assign n2418 = n2402 & n2417 ;
  assign n2419 = n2258 & ~n2418 ;
  assign n2420 = \rf_conf12_reg[15]/NET0131  & n2032 ;
  assign n2421 = \rf_conf14_reg[15]/NET0131  & n2035 ;
  assign n2422 = ~n2420 & ~n2421 ;
  assign n2423 = \rf_conf6_reg[15]/NET0131  & n2051 ;
  assign n2424 = \rf_conf7_reg[15]/NET0131  & n2053 ;
  assign n2425 = ~n2423 & ~n2424 ;
  assign n2426 = n2422 & n2425 ;
  assign n2427 = \rf_conf8_reg[15]/NET0131  & n2057 ;
  assign n2428 = \rf_conf11_reg[15]/NET0131  & n2059 ;
  assign n2429 = ~n2427 & ~n2428 ;
  assign n2430 = \rf_conf1_reg[15]/NET0131  & n2041 ;
  assign n2431 = \rf_conf2_reg[15]/NET0131  & n2039 ;
  assign n2432 = ~n2430 & ~n2431 ;
  assign n2433 = n2429 & n2432 ;
  assign n2434 = n2426 & n2433 ;
  assign n2435 = \rf_conf3_reg[15]/NET0131  & n2027 ;
  assign n2436 = \rf_conf5_reg[15]/NET0131  & n2023 ;
  assign n2437 = ~n2435 & ~n2436 ;
  assign n2438 = \rf_conf9_reg[15]/NET0131  & n2063 ;
  assign n2439 = \rf_conf10_reg[15]/NET0131  & n2065 ;
  assign n2440 = ~n2438 & ~n2439 ;
  assign n2441 = n2437 & n2440 ;
  assign n2442 = \rf_conf4_reg[15]/NET0131  & n2046 ;
  assign n2443 = \rf_conf0_reg[15]/NET0131  & n2044 ;
  assign n2444 = ~n2442 & ~n2443 ;
  assign n2445 = \rf_conf15_reg[15]/NET0131  & n2070 ;
  assign n2446 = \rf_conf13_reg[15]/NET0131  & n2068 ;
  assign n2447 = ~n2445 & ~n2446 ;
  assign n2448 = n2444 & n2447 ;
  assign n2449 = n2441 & n2448 ;
  assign n2450 = n2434 & n2449 ;
  assign n2451 = n2258 & ~n2450 ;
  assign n2452 = \rf_conf4_reg[1]/NET0131  & n2046 ;
  assign n2453 = \rf_conf0_reg[1]/NET0131  & n2044 ;
  assign n2454 = ~n2452 & ~n2453 ;
  assign n2455 = \rf_conf8_reg[1]/NET0131  & n2057 ;
  assign n2456 = \rf_conf11_reg[1]/NET0131  & n2059 ;
  assign n2457 = ~n2455 & ~n2456 ;
  assign n2458 = n2454 & n2457 ;
  assign n2459 = \rf_conf6_reg[1]/NET0131  & n2051 ;
  assign n2460 = \rf_conf7_reg[1]/NET0131  & n2053 ;
  assign n2461 = ~n2459 & ~n2460 ;
  assign n2462 = \rf_conf13_reg[1]/NET0131  & n2068 ;
  assign n2463 = \rf_conf15_reg[1]/NET0131  & n2070 ;
  assign n2464 = ~n2462 & ~n2463 ;
  assign n2465 = n2461 & n2464 ;
  assign n2466 = n2458 & n2465 ;
  assign n2467 = \rf_conf9_reg[1]/NET0131  & n2063 ;
  assign n2468 = \rf_conf10_reg[1]/NET0131  & n2065 ;
  assign n2469 = ~n2467 & ~n2468 ;
  assign n2470 = \rf_conf14_reg[1]/NET0131  & n2035 ;
  assign n2471 = \rf_conf12_reg[1]/NET0131  & n2032 ;
  assign n2472 = ~n2470 & ~n2471 ;
  assign n2473 = n2469 & n2472 ;
  assign n2474 = \rf_conf5_reg[1]/NET0131  & n2023 ;
  assign n2475 = \rf_conf3_reg[1]/NET0131  & n2027 ;
  assign n2476 = ~n2474 & ~n2475 ;
  assign n2477 = \rf_conf1_reg[1]/NET0131  & n2041 ;
  assign n2478 = \rf_conf2_reg[1]/NET0131  & n2039 ;
  assign n2479 = ~n2477 & ~n2478 ;
  assign n2480 = n2476 & n2479 ;
  assign n2481 = n2473 & n2480 ;
  assign n2482 = n2466 & n2481 ;
  assign n2483 = n2258 & ~n2482 ;
  assign n2484 = \rf_conf0_reg[2]/NET0131  & n2044 ;
  assign n2485 = \rf_conf4_reg[2]/NET0131  & n2046 ;
  assign n2486 = ~n2484 & ~n2485 ;
  assign n2487 = \rf_conf5_reg[2]/NET0131  & n2023 ;
  assign n2488 = \rf_conf3_reg[2]/NET0131  & n2027 ;
  assign n2489 = ~n2487 & ~n2488 ;
  assign n2490 = n2486 & n2489 ;
  assign n2491 = \rf_conf15_reg[2]/NET0131  & n2070 ;
  assign n2492 = \rf_conf13_reg[2]/NET0131  & n2068 ;
  assign n2493 = ~n2491 & ~n2492 ;
  assign n2494 = \rf_conf9_reg[2]/NET0131  & n2063 ;
  assign n2495 = \rf_conf10_reg[2]/NET0131  & n2065 ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = n2493 & n2496 ;
  assign n2498 = n2490 & n2497 ;
  assign n2499 = \rf_conf6_reg[2]/NET0131  & n2051 ;
  assign n2500 = \rf_conf7_reg[2]/NET0131  & n2053 ;
  assign n2501 = ~n2499 & ~n2500 ;
  assign n2502 = \rf_conf8_reg[2]/NET0131  & n2057 ;
  assign n2503 = \rf_conf11_reg[2]/NET0131  & n2059 ;
  assign n2504 = ~n2502 & ~n2503 ;
  assign n2505 = n2501 & n2504 ;
  assign n2506 = \rf_conf2_reg[2]/NET0131  & n2039 ;
  assign n2507 = \rf_conf1_reg[2]/NET0131  & n2041 ;
  assign n2508 = ~n2506 & ~n2507 ;
  assign n2509 = \rf_conf12_reg[2]/NET0131  & n2032 ;
  assign n2510 = \rf_conf14_reg[2]/NET0131  & n2035 ;
  assign n2511 = ~n2509 & ~n2510 ;
  assign n2512 = n2508 & n2511 ;
  assign n2513 = n2505 & n2512 ;
  assign n2514 = n2498 & n2513 ;
  assign n2515 = n2258 & ~n2514 ;
  assign n2516 = \rf_conf5_reg[3]/NET0131  & n2023 ;
  assign n2517 = \rf_conf3_reg[3]/NET0131  & n2027 ;
  assign n2518 = ~n2516 & ~n2517 ;
  assign n2519 = \rf_conf13_reg[3]/NET0131  & n2068 ;
  assign n2520 = \rf_conf15_reg[3]/NET0131  & n2070 ;
  assign n2521 = ~n2519 & ~n2520 ;
  assign n2522 = n2518 & n2521 ;
  assign n2523 = \rf_conf8_reg[3]/NET0131  & n2057 ;
  assign n2524 = \rf_conf11_reg[3]/NET0131  & n2059 ;
  assign n2525 = ~n2523 & ~n2524 ;
  assign n2526 = \rf_conf1_reg[3]/NET0131  & n2041 ;
  assign n2527 = \rf_conf2_reg[3]/NET0131  & n2039 ;
  assign n2528 = ~n2526 & ~n2527 ;
  assign n2529 = n2525 & n2528 ;
  assign n2530 = n2522 & n2529 ;
  assign n2531 = \rf_conf14_reg[3]/NET0131  & n2035 ;
  assign n2532 = \rf_conf12_reg[3]/NET0131  & n2032 ;
  assign n2533 = ~n2531 & ~n2532 ;
  assign n2534 = \rf_conf10_reg[3]/NET0131  & n2065 ;
  assign n2535 = \rf_conf9_reg[3]/NET0131  & n2063 ;
  assign n2536 = ~n2534 & ~n2535 ;
  assign n2537 = n2533 & n2536 ;
  assign n2538 = \rf_conf6_reg[3]/NET0131  & n2051 ;
  assign n2539 = \rf_conf7_reg[3]/NET0131  & n2053 ;
  assign n2540 = ~n2538 & ~n2539 ;
  assign n2541 = \rf_conf4_reg[3]/NET0131  & n2046 ;
  assign n2542 = \rf_conf0_reg[3]/NET0131  & n2044 ;
  assign n2543 = ~n2541 & ~n2542 ;
  assign n2544 = n2540 & n2543 ;
  assign n2545 = n2537 & n2544 ;
  assign n2546 = n2530 & n2545 ;
  assign n2547 = n2258 & ~n2546 ;
  assign n2548 = \rf_conf6_reg[4]/NET0131  & n2051 ;
  assign n2549 = \rf_conf7_reg[4]/NET0131  & n2053 ;
  assign n2550 = ~n2548 & ~n2549 ;
  assign n2551 = \rf_conf8_reg[4]/NET0131  & n2057 ;
  assign n2552 = \rf_conf11_reg[4]/NET0131  & n2059 ;
  assign n2553 = ~n2551 & ~n2552 ;
  assign n2554 = n2550 & n2553 ;
  assign n2555 = \rf_conf13_reg[4]/NET0131  & n2068 ;
  assign n2556 = \rf_conf15_reg[4]/NET0131  & n2070 ;
  assign n2557 = ~n2555 & ~n2556 ;
  assign n2558 = \rf_conf10_reg[4]/NET0131  & n2065 ;
  assign n2559 = \rf_conf9_reg[4]/NET0131  & n2063 ;
  assign n2560 = ~n2558 & ~n2559 ;
  assign n2561 = n2557 & n2560 ;
  assign n2562 = n2554 & n2561 ;
  assign n2563 = \rf_conf4_reg[4]/NET0131  & n2046 ;
  assign n2564 = \rf_conf0_reg[4]/NET0131  & n2044 ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = \rf_conf14_reg[4]/NET0131  & n2035 ;
  assign n2567 = \rf_conf12_reg[4]/NET0131  & n2032 ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = n2565 & n2568 ;
  assign n2570 = \rf_conf3_reg[4]/NET0131  & n2027 ;
  assign n2571 = \rf_conf5_reg[4]/NET0131  & n2023 ;
  assign n2572 = ~n2570 & ~n2571 ;
  assign n2573 = \rf_conf1_reg[4]/NET0131  & n2041 ;
  assign n2574 = \rf_conf2_reg[4]/NET0131  & n2039 ;
  assign n2575 = ~n2573 & ~n2574 ;
  assign n2576 = n2572 & n2575 ;
  assign n2577 = n2569 & n2576 ;
  assign n2578 = n2562 & n2577 ;
  assign n2579 = n2258 & ~n2578 ;
  assign n2580 = \rf_conf6_reg[5]/NET0131  & n2051 ;
  assign n2581 = \rf_conf7_reg[5]/NET0131  & n2053 ;
  assign n2582 = ~n2580 & ~n2581 ;
  assign n2583 = \rf_conf8_reg[5]/NET0131  & n2057 ;
  assign n2584 = \rf_conf11_reg[5]/NET0131  & n2059 ;
  assign n2585 = ~n2583 & ~n2584 ;
  assign n2586 = n2582 & n2585 ;
  assign n2587 = \rf_conf13_reg[5]/NET0131  & n2068 ;
  assign n2588 = \rf_conf15_reg[5]/NET0131  & n2070 ;
  assign n2589 = ~n2587 & ~n2588 ;
  assign n2590 = \rf_conf10_reg[5]/NET0131  & n2065 ;
  assign n2591 = \rf_conf9_reg[5]/NET0131  & n2063 ;
  assign n2592 = ~n2590 & ~n2591 ;
  assign n2593 = n2589 & n2592 ;
  assign n2594 = n2586 & n2593 ;
  assign n2595 = \rf_conf4_reg[5]/NET0131  & n2046 ;
  assign n2596 = \rf_conf0_reg[5]/NET0131  & n2044 ;
  assign n2597 = ~n2595 & ~n2596 ;
  assign n2598 = \rf_conf14_reg[5]/NET0131  & n2035 ;
  assign n2599 = \rf_conf12_reg[5]/NET0131  & n2032 ;
  assign n2600 = ~n2598 & ~n2599 ;
  assign n2601 = n2597 & n2600 ;
  assign n2602 = \rf_conf5_reg[5]/NET0131  & n2023 ;
  assign n2603 = \rf_conf3_reg[5]/NET0131  & n2027 ;
  assign n2604 = ~n2602 & ~n2603 ;
  assign n2605 = \rf_conf1_reg[5]/NET0131  & n2041 ;
  assign n2606 = \rf_conf2_reg[5]/NET0131  & n2039 ;
  assign n2607 = ~n2605 & ~n2606 ;
  assign n2608 = n2604 & n2607 ;
  assign n2609 = n2601 & n2608 ;
  assign n2610 = n2594 & n2609 ;
  assign n2611 = n2258 & ~n2610 ;
  assign n2612 = \rf_conf11_reg[6]/NET0131  & n2059 ;
  assign n2613 = \rf_conf15_reg[6]/NET0131  & n2070 ;
  assign n2614 = ~n2612 & ~n2613 ;
  assign n2615 = \rf_conf0_reg[6]/NET0131  & n2044 ;
  assign n2616 = \rf_conf4_reg[6]/NET0131  & n2046 ;
  assign n2617 = ~n2615 & ~n2616 ;
  assign n2618 = n2614 & n2617 ;
  assign n2619 = \rf_conf9_reg[6]/NET0131  & n2063 ;
  assign n2620 = \rf_conf6_reg[6]/NET0131  & n2051 ;
  assign n2621 = ~n2619 & ~n2620 ;
  assign n2622 = \rf_conf13_reg[6]/NET0131  & n2068 ;
  assign n2623 = \rf_conf8_reg[6]/NET0131  & n2057 ;
  assign n2624 = ~n2622 & ~n2623 ;
  assign n2625 = n2621 & n2624 ;
  assign n2626 = n2618 & n2625 ;
  assign n2627 = \rf_conf7_reg[6]/NET0131  & n2053 ;
  assign n2628 = \rf_conf10_reg[6]/NET0131  & n2065 ;
  assign n2629 = ~n2627 & ~n2628 ;
  assign n2630 = \rf_conf2_reg[6]/NET0131  & n2039 ;
  assign n2631 = \rf_conf1_reg[6]/NET0131  & n2041 ;
  assign n2632 = ~n2630 & ~n2631 ;
  assign n2633 = n2629 & n2632 ;
  assign n2634 = \rf_conf12_reg[6]/NET0131  & n2032 ;
  assign n2635 = \rf_conf14_reg[6]/NET0131  & n2035 ;
  assign n2636 = ~n2634 & ~n2635 ;
  assign n2637 = \rf_conf3_reg[6]/NET0131  & n2027 ;
  assign n2638 = \rf_conf5_reg[6]/NET0131  & n2023 ;
  assign n2639 = ~n2637 & ~n2638 ;
  assign n2640 = n2636 & n2639 ;
  assign n2641 = n2633 & n2640 ;
  assign n2642 = n2626 & n2641 ;
  assign n2643 = n2258 & ~n2642 ;
  assign n2644 = \rf_conf8_reg[7]/NET0131  & n2057 ;
  assign n2645 = \rf_conf11_reg[7]/NET0131  & n2059 ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = \rf_conf13_reg[7]/NET0131  & n2068 ;
  assign n2648 = \rf_conf15_reg[7]/NET0131  & n2070 ;
  assign n2649 = ~n2647 & ~n2648 ;
  assign n2650 = n2646 & n2649 ;
  assign n2651 = \rf_conf14_reg[7]/NET0131  & n2035 ;
  assign n2652 = \rf_conf12_reg[7]/NET0131  & n2032 ;
  assign n2653 = ~n2651 & ~n2652 ;
  assign n2654 = \rf_conf5_reg[7]/NET0131  & n2023 ;
  assign n2655 = \rf_conf3_reg[7]/NET0131  & n2027 ;
  assign n2656 = ~n2654 & ~n2655 ;
  assign n2657 = n2653 & n2656 ;
  assign n2658 = n2650 & n2657 ;
  assign n2659 = \rf_conf1_reg[7]/NET0131  & n2041 ;
  assign n2660 = \rf_conf2_reg[7]/NET0131  & n2039 ;
  assign n2661 = ~n2659 & ~n2660 ;
  assign n2662 = \rf_conf6_reg[7]/NET0131  & n2051 ;
  assign n2663 = \rf_conf7_reg[7]/NET0131  & n2053 ;
  assign n2664 = ~n2662 & ~n2663 ;
  assign n2665 = n2661 & n2664 ;
  assign n2666 = \rf_conf10_reg[7]/NET0131  & n2065 ;
  assign n2667 = \rf_conf9_reg[7]/NET0131  & n2063 ;
  assign n2668 = ~n2666 & ~n2667 ;
  assign n2669 = \rf_conf4_reg[7]/NET0131  & n2046 ;
  assign n2670 = \rf_conf0_reg[7]/NET0131  & n2044 ;
  assign n2671 = ~n2669 & ~n2670 ;
  assign n2672 = n2668 & n2671 ;
  assign n2673 = n2665 & n2672 ;
  assign n2674 = n2658 & n2673 ;
  assign n2675 = n2258 & ~n2674 ;
  assign n2676 = \rf_conf14_reg[8]/NET0131  & n2035 ;
  assign n2677 = \rf_conf12_reg[8]/NET0131  & n2032 ;
  assign n2678 = ~n2676 & ~n2677 ;
  assign n2679 = \rf_conf13_reg[8]/NET0131  & n2068 ;
  assign n2680 = \rf_conf15_reg[8]/NET0131  & n2070 ;
  assign n2681 = ~n2679 & ~n2680 ;
  assign n2682 = n2678 & n2681 ;
  assign n2683 = \rf_conf8_reg[8]/NET0131  & n2057 ;
  assign n2684 = \rf_conf11_reg[8]/NET0131  & n2059 ;
  assign n2685 = ~n2683 & ~n2684 ;
  assign n2686 = \rf_conf1_reg[8]/NET0131  & n2041 ;
  assign n2687 = \rf_conf2_reg[8]/NET0131  & n2039 ;
  assign n2688 = ~n2686 & ~n2687 ;
  assign n2689 = n2685 & n2688 ;
  assign n2690 = n2682 & n2689 ;
  assign n2691 = \rf_conf5_reg[8]/NET0131  & n2023 ;
  assign n2692 = \rf_conf3_reg[8]/NET0131  & n2027 ;
  assign n2693 = ~n2691 & ~n2692 ;
  assign n2694 = \rf_conf10_reg[8]/NET0131  & n2065 ;
  assign n2695 = \rf_conf9_reg[8]/NET0131  & n2063 ;
  assign n2696 = ~n2694 & ~n2695 ;
  assign n2697 = n2693 & n2696 ;
  assign n2698 = \rf_conf6_reg[8]/NET0131  & n2051 ;
  assign n2699 = \rf_conf7_reg[8]/NET0131  & n2053 ;
  assign n2700 = ~n2698 & ~n2699 ;
  assign n2701 = \rf_conf4_reg[8]/NET0131  & n2046 ;
  assign n2702 = \rf_conf0_reg[8]/NET0131  & n2044 ;
  assign n2703 = ~n2701 & ~n2702 ;
  assign n2704 = n2700 & n2703 ;
  assign n2705 = n2697 & n2704 ;
  assign n2706 = n2690 & n2705 ;
  assign n2707 = n2258 & ~n2706 ;
  assign n2708 = \rf_conf6_reg[9]/NET0131  & n2051 ;
  assign n2709 = \rf_conf7_reg[9]/NET0131  & n2053 ;
  assign n2710 = ~n2708 & ~n2709 ;
  assign n2711 = \rf_conf14_reg[9]/NET0131  & n2035 ;
  assign n2712 = \rf_conf12_reg[9]/NET0131  & n2032 ;
  assign n2713 = ~n2711 & ~n2712 ;
  assign n2714 = n2710 & n2713 ;
  assign n2715 = \rf_conf13_reg[9]/NET0131  & n2068 ;
  assign n2716 = \rf_conf15_reg[9]/NET0131  & n2070 ;
  assign n2717 = ~n2715 & ~n2716 ;
  assign n2718 = \rf_conf10_reg[9]/NET0131  & n2065 ;
  assign n2719 = \rf_conf9_reg[9]/NET0131  & n2063 ;
  assign n2720 = ~n2718 & ~n2719 ;
  assign n2721 = n2717 & n2720 ;
  assign n2722 = n2714 & n2721 ;
  assign n2723 = \rf_conf4_reg[9]/NET0131  & n2046 ;
  assign n2724 = \rf_conf0_reg[9]/NET0131  & n2044 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = \rf_conf8_reg[9]/NET0131  & n2057 ;
  assign n2727 = \rf_conf11_reg[9]/NET0131  & n2059 ;
  assign n2728 = ~n2726 & ~n2727 ;
  assign n2729 = n2725 & n2728 ;
  assign n2730 = \rf_conf5_reg[9]/NET0131  & n2023 ;
  assign n2731 = \rf_conf3_reg[9]/NET0131  & n2027 ;
  assign n2732 = ~n2730 & ~n2731 ;
  assign n2733 = \rf_conf1_reg[9]/NET0131  & n2041 ;
  assign n2734 = \rf_conf2_reg[9]/NET0131  & n2039 ;
  assign n2735 = ~n2733 & ~n2734 ;
  assign n2736 = n2732 & n2735 ;
  assign n2737 = n2729 & n2736 ;
  assign n2738 = n2722 & n2737 ;
  assign n2739 = n2258 & ~n2738 ;
  assign n2740 = \m5_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[10]/NET0131  ;
  assign n2741 = ~\rf_conf11_reg[11]/NET0131  & n2740 ;
  assign n2742 = \m4_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[8]/NET0131  ;
  assign n2743 = ~\rf_conf11_reg[9]/NET0131  & n2742 ;
  assign n2744 = ~n2741 & ~n2743 ;
  assign n2745 = \m7_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[14]/NET0131  ;
  assign n2746 = ~\rf_conf11_reg[15]/NET0131  & n2745 ;
  assign n2747 = \m6_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[12]/NET0131  ;
  assign n2748 = ~\rf_conf11_reg[13]/NET0131  & n2747 ;
  assign n2749 = ~n2746 & ~n2748 ;
  assign n2750 = \m1_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[2]/NET0131  ;
  assign n2751 = ~\rf_conf11_reg[3]/NET0131  & n2750 ;
  assign n2752 = \m0_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[0]/NET0131  ;
  assign n2753 = ~\rf_conf11_reg[1]/NET0131  & n2752 ;
  assign n2754 = ~n2751 & ~n2753 ;
  assign n2755 = n2749 & ~n2754 ;
  assign n2756 = n2744 & ~n2755 ;
  assign n2757 = \m3_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[6]/NET0131  ;
  assign n2758 = ~\rf_conf11_reg[7]/NET0131  & n2757 ;
  assign n2759 = ~\s11_msel_arb0_state_reg[2]/NET0131  & ~n2758 ;
  assign n2760 = ~n2756 & n2759 ;
  assign n2761 = \s11_msel_arb0_state_reg[2]/NET0131  & ~n2746 ;
  assign n2762 = \s11_msel_arb0_state_reg[1]/NET0131  & ~n2761 ;
  assign n2763 = \m2_s11_cyc_o_reg/NET0131  & ~\rf_conf11_reg[4]/NET0131  ;
  assign n2764 = ~\rf_conf11_reg[5]/NET0131  & n2763 ;
  assign n2765 = ~n2758 & ~n2764 ;
  assign n2766 = ~n2744 & n2765 ;
  assign n2767 = \s11_msel_arb0_state_reg[1]/NET0131  & n2754 ;
  assign n2768 = ~n2766 & n2767 ;
  assign n2769 = ~n2762 & ~n2768 ;
  assign n2770 = ~n2760 & ~n2769 ;
  assign n2771 = \s11_msel_arb0_state_reg[0]/NET0131  & n2770 ;
  assign n2772 = \s11_msel_arb0_state_reg[2]/NET0131  & ~n2749 ;
  assign n2773 = ~n2741 & n2772 ;
  assign n2774 = ~n2743 & ~n2749 ;
  assign n2775 = ~n2753 & ~n2765 ;
  assign n2776 = ~n2774 & ~n2775 ;
  assign n2777 = ~n2741 & ~n2751 ;
  assign n2778 = ~n2776 & n2777 ;
  assign n2779 = ~n2773 & ~n2778 ;
  assign n2780 = ~\s11_msel_arb0_state_reg[2]/NET0131  & ~n2751 ;
  assign n2781 = ~n2765 & n2780 ;
  assign n2782 = n2779 & ~n2781 ;
  assign n2783 = \s11_msel_arb0_state_reg[0]/NET0131  & ~\s11_msel_arb0_state_reg[1]/NET0131  ;
  assign n2784 = ~n2782 & n2783 ;
  assign n2785 = ~n2771 & ~n2784 ;
  assign n2786 = ~\s11_msel_arb0_state_reg[2]/NET0131  & n2766 ;
  assign n2787 = ~\s11_msel_arb0_state_reg[1]/NET0131  & ~\s11_msel_arb0_state_reg[2]/NET0131  ;
  assign n2788 = ~n2754 & n2787 ;
  assign n2789 = ~n2786 & ~n2788 ;
  assign n2790 = \s11_msel_arb0_state_reg[2]/NET0131  & n2755 ;
  assign n2791 = ~\s11_msel_arb0_state_reg[1]/NET0131  & \s11_msel_arb0_state_reg[2]/NET0131  ;
  assign n2792 = ~n2744 & n2791 ;
  assign n2793 = ~n2790 & ~n2792 ;
  assign n2794 = n2749 & n2765 ;
  assign n2795 = ~\s11_msel_arb0_state_reg[0]/NET0131  & ~n2794 ;
  assign n2796 = ~\s11_msel_arb0_state_reg[0]/NET0131  & n2744 ;
  assign n2797 = n2767 & n2796 ;
  assign n2798 = ~n2795 & ~n2797 ;
  assign n2799 = n2793 & ~n2798 ;
  assign n2800 = n2789 & n2799 ;
  assign n2801 = n2785 & ~n2800 ;
  assign n2802 = \m5_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[10]/NET0131  ;
  assign n2803 = ~\rf_conf12_reg[11]/NET0131  & n2802 ;
  assign n2804 = \m4_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[8]/NET0131  ;
  assign n2805 = ~\rf_conf12_reg[9]/NET0131  & n2804 ;
  assign n2806 = ~n2803 & ~n2805 ;
  assign n2807 = \m7_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[14]/NET0131  ;
  assign n2808 = ~\rf_conf12_reg[15]/NET0131  & n2807 ;
  assign n2809 = \m6_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[12]/NET0131  ;
  assign n2810 = ~\rf_conf12_reg[13]/NET0131  & n2809 ;
  assign n2811 = ~n2808 & ~n2810 ;
  assign n2812 = \m1_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[2]/NET0131  ;
  assign n2813 = ~\rf_conf12_reg[3]/NET0131  & n2812 ;
  assign n2814 = \m0_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[0]/NET0131  ;
  assign n2815 = ~\rf_conf12_reg[1]/NET0131  & n2814 ;
  assign n2816 = ~n2813 & ~n2815 ;
  assign n2817 = n2811 & ~n2816 ;
  assign n2818 = n2806 & ~n2817 ;
  assign n2819 = \m3_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[6]/NET0131  ;
  assign n2820 = ~\rf_conf12_reg[7]/NET0131  & n2819 ;
  assign n2821 = ~\s12_msel_arb0_state_reg[2]/NET0131  & ~n2820 ;
  assign n2822 = ~n2818 & n2821 ;
  assign n2823 = \s12_msel_arb0_state_reg[2]/NET0131  & ~n2808 ;
  assign n2824 = \s12_msel_arb0_state_reg[1]/NET0131  & ~n2823 ;
  assign n2825 = \m2_s12_cyc_o_reg/NET0131  & ~\rf_conf12_reg[4]/NET0131  ;
  assign n2826 = ~\rf_conf12_reg[5]/NET0131  & n2825 ;
  assign n2827 = ~n2820 & ~n2826 ;
  assign n2828 = ~n2806 & n2827 ;
  assign n2829 = \s12_msel_arb0_state_reg[1]/NET0131  & n2816 ;
  assign n2830 = ~n2828 & n2829 ;
  assign n2831 = ~n2824 & ~n2830 ;
  assign n2832 = ~n2822 & ~n2831 ;
  assign n2833 = \s12_msel_arb0_state_reg[0]/NET0131  & n2832 ;
  assign n2834 = \s12_msel_arb0_state_reg[2]/NET0131  & ~n2811 ;
  assign n2835 = ~n2803 & n2834 ;
  assign n2836 = ~n2805 & ~n2811 ;
  assign n2837 = ~n2815 & ~n2827 ;
  assign n2838 = ~n2836 & ~n2837 ;
  assign n2839 = ~n2803 & ~n2813 ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2841 = ~n2835 & ~n2840 ;
  assign n2842 = ~\s12_msel_arb0_state_reg[2]/NET0131  & ~n2813 ;
  assign n2843 = ~n2827 & n2842 ;
  assign n2844 = n2841 & ~n2843 ;
  assign n2845 = \s12_msel_arb0_state_reg[0]/NET0131  & ~\s12_msel_arb0_state_reg[1]/NET0131  ;
  assign n2846 = ~n2844 & n2845 ;
  assign n2847 = ~n2833 & ~n2846 ;
  assign n2848 = ~\s12_msel_arb0_state_reg[2]/NET0131  & n2828 ;
  assign n2849 = ~\s12_msel_arb0_state_reg[1]/NET0131  & ~\s12_msel_arb0_state_reg[2]/NET0131  ;
  assign n2850 = ~n2816 & n2849 ;
  assign n2851 = ~n2848 & ~n2850 ;
  assign n2852 = \s12_msel_arb0_state_reg[2]/NET0131  & n2817 ;
  assign n2853 = ~\s12_msel_arb0_state_reg[1]/NET0131  & \s12_msel_arb0_state_reg[2]/NET0131  ;
  assign n2854 = ~n2806 & n2853 ;
  assign n2855 = ~n2852 & ~n2854 ;
  assign n2856 = n2811 & n2827 ;
  assign n2857 = ~\s12_msel_arb0_state_reg[0]/NET0131  & ~n2856 ;
  assign n2858 = ~\s12_msel_arb0_state_reg[0]/NET0131  & n2806 ;
  assign n2859 = n2829 & n2858 ;
  assign n2860 = ~n2857 & ~n2859 ;
  assign n2861 = n2855 & ~n2860 ;
  assign n2862 = n2851 & n2861 ;
  assign n2863 = n2847 & ~n2862 ;
  assign n2864 = \m5_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[10]/NET0131  ;
  assign n2865 = ~\rf_conf13_reg[11]/NET0131  & n2864 ;
  assign n2866 = \m4_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[8]/NET0131  ;
  assign n2867 = ~\rf_conf13_reg[9]/NET0131  & n2866 ;
  assign n2868 = ~n2865 & ~n2867 ;
  assign n2869 = \m7_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[14]/NET0131  ;
  assign n2870 = ~\rf_conf13_reg[15]/NET0131  & n2869 ;
  assign n2871 = \m6_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[12]/NET0131  ;
  assign n2872 = ~\rf_conf13_reg[13]/NET0131  & n2871 ;
  assign n2873 = ~n2870 & ~n2872 ;
  assign n2874 = \m1_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[2]/NET0131  ;
  assign n2875 = ~\rf_conf13_reg[3]/NET0131  & n2874 ;
  assign n2876 = \m0_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[0]/NET0131  ;
  assign n2877 = ~\rf_conf13_reg[1]/NET0131  & n2876 ;
  assign n2878 = ~n2875 & ~n2877 ;
  assign n2879 = n2873 & ~n2878 ;
  assign n2880 = n2868 & ~n2879 ;
  assign n2881 = \m3_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[6]/NET0131  ;
  assign n2882 = ~\rf_conf13_reg[7]/NET0131  & n2881 ;
  assign n2883 = ~\s13_msel_arb0_state_reg[2]/NET0131  & ~n2882 ;
  assign n2884 = ~n2880 & n2883 ;
  assign n2885 = \s13_msel_arb0_state_reg[2]/NET0131  & ~n2870 ;
  assign n2886 = \s13_msel_arb0_state_reg[1]/NET0131  & ~n2885 ;
  assign n2887 = \m2_s13_cyc_o_reg/NET0131  & ~\rf_conf13_reg[4]/NET0131  ;
  assign n2888 = ~\rf_conf13_reg[5]/NET0131  & n2887 ;
  assign n2889 = ~n2882 & ~n2888 ;
  assign n2890 = ~n2868 & n2889 ;
  assign n2891 = \s13_msel_arb0_state_reg[1]/NET0131  & n2878 ;
  assign n2892 = ~n2890 & n2891 ;
  assign n2893 = ~n2886 & ~n2892 ;
  assign n2894 = ~n2884 & ~n2893 ;
  assign n2895 = \s13_msel_arb0_state_reg[0]/NET0131  & n2894 ;
  assign n2896 = \s13_msel_arb0_state_reg[2]/NET0131  & ~n2873 ;
  assign n2897 = ~n2865 & n2896 ;
  assign n2898 = ~n2867 & ~n2873 ;
  assign n2899 = ~n2877 & ~n2889 ;
  assign n2900 = ~n2898 & ~n2899 ;
  assign n2901 = ~n2865 & ~n2875 ;
  assign n2902 = ~n2900 & n2901 ;
  assign n2903 = ~n2897 & ~n2902 ;
  assign n2904 = ~\s13_msel_arb0_state_reg[2]/NET0131  & ~n2875 ;
  assign n2905 = ~n2889 & n2904 ;
  assign n2906 = n2903 & ~n2905 ;
  assign n2907 = \s13_msel_arb0_state_reg[0]/NET0131  & ~\s13_msel_arb0_state_reg[1]/NET0131  ;
  assign n2908 = ~n2906 & n2907 ;
  assign n2909 = ~n2895 & ~n2908 ;
  assign n2910 = ~\s13_msel_arb0_state_reg[2]/NET0131  & n2890 ;
  assign n2911 = ~\s13_msel_arb0_state_reg[1]/NET0131  & ~\s13_msel_arb0_state_reg[2]/NET0131  ;
  assign n2912 = ~n2878 & n2911 ;
  assign n2913 = ~n2910 & ~n2912 ;
  assign n2914 = \s13_msel_arb0_state_reg[2]/NET0131  & n2879 ;
  assign n2915 = ~\s13_msel_arb0_state_reg[1]/NET0131  & \s13_msel_arb0_state_reg[2]/NET0131  ;
  assign n2916 = ~n2868 & n2915 ;
  assign n2917 = ~n2914 & ~n2916 ;
  assign n2918 = n2873 & n2889 ;
  assign n2919 = ~\s13_msel_arb0_state_reg[0]/NET0131  & ~n2918 ;
  assign n2920 = ~\s13_msel_arb0_state_reg[0]/NET0131  & n2868 ;
  assign n2921 = n2891 & n2920 ;
  assign n2922 = ~n2919 & ~n2921 ;
  assign n2923 = n2917 & ~n2922 ;
  assign n2924 = n2913 & n2923 ;
  assign n2925 = n2909 & ~n2924 ;
  assign n2926 = \m5_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[10]/NET0131  ;
  assign n2927 = ~\rf_conf14_reg[11]/NET0131  & n2926 ;
  assign n2928 = \m4_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[8]/NET0131  ;
  assign n2929 = ~\rf_conf14_reg[9]/NET0131  & n2928 ;
  assign n2930 = ~n2927 & ~n2929 ;
  assign n2931 = \m7_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[14]/NET0131  ;
  assign n2932 = ~\rf_conf14_reg[15]/NET0131  & n2931 ;
  assign n2933 = \m6_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[12]/NET0131  ;
  assign n2934 = ~\rf_conf14_reg[13]/NET0131  & n2933 ;
  assign n2935 = ~n2932 & ~n2934 ;
  assign n2936 = \m1_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[2]/NET0131  ;
  assign n2937 = ~\rf_conf14_reg[3]/NET0131  & n2936 ;
  assign n2938 = \m0_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[0]/NET0131  ;
  assign n2939 = ~\rf_conf14_reg[1]/NET0131  & n2938 ;
  assign n2940 = ~n2937 & ~n2939 ;
  assign n2941 = n2935 & ~n2940 ;
  assign n2942 = n2930 & ~n2941 ;
  assign n2943 = \m3_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[6]/NET0131  ;
  assign n2944 = ~\rf_conf14_reg[7]/NET0131  & n2943 ;
  assign n2945 = ~\s14_msel_arb0_state_reg[2]/NET0131  & ~n2944 ;
  assign n2946 = ~n2942 & n2945 ;
  assign n2947 = \s14_msel_arb0_state_reg[2]/NET0131  & ~n2932 ;
  assign n2948 = \s14_msel_arb0_state_reg[1]/NET0131  & ~n2947 ;
  assign n2949 = \m2_s14_cyc_o_reg/NET0131  & ~\rf_conf14_reg[4]/NET0131  ;
  assign n2950 = ~\rf_conf14_reg[5]/NET0131  & n2949 ;
  assign n2951 = ~n2944 & ~n2950 ;
  assign n2952 = ~n2930 & n2951 ;
  assign n2953 = \s14_msel_arb0_state_reg[1]/NET0131  & n2940 ;
  assign n2954 = ~n2952 & n2953 ;
  assign n2955 = ~n2948 & ~n2954 ;
  assign n2956 = ~n2946 & ~n2955 ;
  assign n2957 = \s14_msel_arb0_state_reg[0]/NET0131  & n2956 ;
  assign n2958 = \s14_msel_arb0_state_reg[2]/NET0131  & ~n2935 ;
  assign n2959 = ~n2927 & n2958 ;
  assign n2960 = ~n2929 & ~n2935 ;
  assign n2961 = ~n2939 & ~n2951 ;
  assign n2962 = ~n2960 & ~n2961 ;
  assign n2963 = ~n2927 & ~n2937 ;
  assign n2964 = ~n2962 & n2963 ;
  assign n2965 = ~n2959 & ~n2964 ;
  assign n2966 = ~\s14_msel_arb0_state_reg[2]/NET0131  & ~n2937 ;
  assign n2967 = ~n2951 & n2966 ;
  assign n2968 = n2965 & ~n2967 ;
  assign n2969 = \s14_msel_arb0_state_reg[0]/NET0131  & ~\s14_msel_arb0_state_reg[1]/NET0131  ;
  assign n2970 = ~n2968 & n2969 ;
  assign n2971 = ~n2957 & ~n2970 ;
  assign n2972 = ~\s14_msel_arb0_state_reg[2]/NET0131  & n2952 ;
  assign n2973 = ~\s14_msel_arb0_state_reg[1]/NET0131  & ~\s14_msel_arb0_state_reg[2]/NET0131  ;
  assign n2974 = ~n2940 & n2973 ;
  assign n2975 = ~n2972 & ~n2974 ;
  assign n2976 = \s14_msel_arb0_state_reg[2]/NET0131  & n2941 ;
  assign n2977 = ~\s14_msel_arb0_state_reg[1]/NET0131  & \s14_msel_arb0_state_reg[2]/NET0131  ;
  assign n2978 = ~n2930 & n2977 ;
  assign n2979 = ~n2976 & ~n2978 ;
  assign n2980 = n2935 & n2951 ;
  assign n2981 = ~\s14_msel_arb0_state_reg[0]/NET0131  & ~n2980 ;
  assign n2982 = ~\s14_msel_arb0_state_reg[0]/NET0131  & n2930 ;
  assign n2983 = n2953 & n2982 ;
  assign n2984 = ~n2981 & ~n2983 ;
  assign n2985 = n2979 & ~n2984 ;
  assign n2986 = n2975 & n2985 ;
  assign n2987 = n2971 & ~n2986 ;
  assign n2988 = \m5_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[10]/NET0131  ;
  assign n2989 = ~\rf_conf15_reg[11]/NET0131  & n2988 ;
  assign n2990 = \m4_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[8]/NET0131  ;
  assign n2991 = ~\rf_conf15_reg[9]/NET0131  & n2990 ;
  assign n2992 = ~n2989 & ~n2991 ;
  assign n2993 = \m6_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[12]/NET0131  ;
  assign n2994 = ~\rf_conf15_reg[13]/NET0131  & n2993 ;
  assign n2995 = \m7_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[14]/NET0131  ;
  assign n2996 = ~\rf_conf15_reg[15]/NET0131  & n2995 ;
  assign n2997 = ~n2994 & ~n2996 ;
  assign n2998 = ~\s15_msel_arb0_state_reg[0]/NET0131  & ~\s15_msel_arb0_state_reg[1]/NET0131  ;
  assign n2999 = \s15_msel_arb0_state_reg[2]/NET0131  & n2998 ;
  assign n3000 = ~n2997 & n2999 ;
  assign n3001 = \m3_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[6]/NET0131  ;
  assign n3002 = ~\rf_conf15_reg[7]/NET0131  & n3001 ;
  assign n3003 = \m2_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[4]/NET0131  ;
  assign n3004 = ~\rf_conf15_reg[5]/NET0131  & n3003 ;
  assign n3005 = ~n3002 & ~n3004 ;
  assign n3006 = ~\s15_msel_arb0_state_reg[1]/NET0131  & n3005 ;
  assign n3007 = \m1_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[2]/NET0131  ;
  assign n3008 = ~\rf_conf15_reg[3]/NET0131  & n3007 ;
  assign n3009 = \m0_s15_cyc_o_reg/NET0131  & ~\rf_conf15_reg[0]/NET0131  ;
  assign n3010 = ~\rf_conf15_reg[1]/NET0131  & n3009 ;
  assign n3011 = ~n3008 & ~n3010 ;
  assign n3012 = n2999 & n3011 ;
  assign n3013 = ~n3006 & n3012 ;
  assign n3014 = ~n3000 & ~n3013 ;
  assign n3015 = n2997 & ~n3011 ;
  assign n3016 = \s15_msel_arb0_state_reg[0]/NET0131  & \s15_msel_arb0_state_reg[1]/NET0131  ;
  assign n3017 = ~\s15_msel_arb0_state_reg[2]/NET0131  & n3016 ;
  assign n3018 = ~n3002 & n3017 ;
  assign n3019 = ~n3015 & n3018 ;
  assign n3020 = n3014 & ~n3019 ;
  assign n3021 = n2992 & ~n3020 ;
  assign n3022 = ~n2992 & n3005 ;
  assign n3023 = \s15_msel_arb0_state_reg[1]/NET0131  & ~n2996 ;
  assign n3024 = ~n3022 & n3023 ;
  assign n3025 = ~\s15_msel_arb0_state_reg[1]/NET0131  & ~n2989 ;
  assign n3026 = ~n3005 & n3025 ;
  assign n3027 = ~n3024 & ~n3026 ;
  assign n3028 = \s15_msel_arb0_state_reg[0]/NET0131  & \s15_msel_arb0_state_reg[2]/NET0131  ;
  assign n3029 = n3011 & n3028 ;
  assign n3030 = ~n3027 & n3029 ;
  assign n3031 = ~\s15_msel_arb0_state_reg[2]/NET0131  & ~n3005 ;
  assign n3032 = n3015 & ~n3031 ;
  assign n3033 = \s15_msel_arb0_state_reg[2]/NET0131  & ~n2997 ;
  assign n3034 = n3022 & ~n3033 ;
  assign n3035 = ~\s15_msel_arb0_state_reg[0]/NET0131  & \s15_msel_arb0_state_reg[1]/NET0131  ;
  assign n3036 = ~n3034 & n3035 ;
  assign n3037 = ~n3032 & n3036 ;
  assign n3038 = n2992 & ~n2997 ;
  assign n3039 = n3005 & ~n3038 ;
  assign n3040 = \s15_msel_arb0_state_reg[0]/NET0131  & ~\s15_msel_arb0_state_reg[1]/NET0131  ;
  assign n3041 = ~\s15_msel_arb0_state_reg[2]/NET0131  & n3040 ;
  assign n3042 = ~n3008 & n3041 ;
  assign n3043 = ~\s15_msel_arb0_state_reg[2]/NET0131  & n2998 ;
  assign n3044 = n3011 & n3043 ;
  assign n3045 = ~n3042 & ~n3044 ;
  assign n3046 = ~n3039 & ~n3045 ;
  assign n3047 = \s15_msel_arb0_state_reg[2]/NET0131  & n3040 ;
  assign n3048 = ~n2989 & n3047 ;
  assign n3049 = ~n2997 & n3048 ;
  assign n3050 = n3002 & n3017 ;
  assign n3051 = \s15_msel_arb0_state_reg[2]/NET0131  & n3016 ;
  assign n3052 = n2996 & n3051 ;
  assign n3053 = ~n3050 & ~n3052 ;
  assign n3054 = ~n3049 & n3053 ;
  assign n3055 = ~n3046 & n3054 ;
  assign n3056 = ~n3037 & n3055 ;
  assign n3057 = ~n3030 & n3056 ;
  assign n3058 = ~n3021 & n3057 ;
  assign n3059 = \m5_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[10]/NET0131  ;
  assign n3060 = ~\rf_conf3_reg[11]/NET0131  & n3059 ;
  assign n3061 = \m4_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[8]/NET0131  ;
  assign n3062 = ~\rf_conf3_reg[9]/NET0131  & n3061 ;
  assign n3063 = ~n3060 & ~n3062 ;
  assign n3064 = \m7_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[14]/NET0131  ;
  assign n3065 = ~\rf_conf3_reg[15]/NET0131  & n3064 ;
  assign n3066 = \m6_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[12]/NET0131  ;
  assign n3067 = ~\rf_conf3_reg[13]/NET0131  & n3066 ;
  assign n3068 = ~n3065 & ~n3067 ;
  assign n3069 = \m1_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[2]/NET0131  ;
  assign n3070 = ~\rf_conf3_reg[3]/NET0131  & n3069 ;
  assign n3071 = \m0_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[0]/NET0131  ;
  assign n3072 = ~\rf_conf3_reg[1]/NET0131  & n3071 ;
  assign n3073 = ~n3070 & ~n3072 ;
  assign n3074 = n3068 & ~n3073 ;
  assign n3075 = n3063 & ~n3074 ;
  assign n3076 = \m3_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[6]/NET0131  ;
  assign n3077 = ~\rf_conf3_reg[7]/NET0131  & n3076 ;
  assign n3078 = ~\s3_msel_arb0_state_reg[2]/NET0131  & ~n3077 ;
  assign n3079 = ~n3075 & n3078 ;
  assign n3080 = \s3_msel_arb0_state_reg[2]/NET0131  & ~n3065 ;
  assign n3081 = \s3_msel_arb0_state_reg[1]/NET0131  & ~n3080 ;
  assign n3082 = \m2_s3_cyc_o_reg/NET0131  & ~\rf_conf3_reg[4]/NET0131  ;
  assign n3083 = ~\rf_conf3_reg[5]/NET0131  & n3082 ;
  assign n3084 = ~n3077 & ~n3083 ;
  assign n3085 = ~n3063 & n3084 ;
  assign n3086 = \s3_msel_arb0_state_reg[1]/NET0131  & n3073 ;
  assign n3087 = ~n3085 & n3086 ;
  assign n3088 = ~n3081 & ~n3087 ;
  assign n3089 = ~n3079 & ~n3088 ;
  assign n3090 = \s3_msel_arb0_state_reg[0]/NET0131  & n3089 ;
  assign n3091 = \s3_msel_arb0_state_reg[2]/NET0131  & ~n3068 ;
  assign n3092 = ~n3060 & n3091 ;
  assign n3093 = ~n3062 & ~n3068 ;
  assign n3094 = ~n3072 & ~n3084 ;
  assign n3095 = ~n3093 & ~n3094 ;
  assign n3096 = ~n3060 & ~n3070 ;
  assign n3097 = ~n3095 & n3096 ;
  assign n3098 = ~n3092 & ~n3097 ;
  assign n3099 = ~\s3_msel_arb0_state_reg[2]/NET0131  & ~n3070 ;
  assign n3100 = ~n3084 & n3099 ;
  assign n3101 = n3098 & ~n3100 ;
  assign n3102 = \s3_msel_arb0_state_reg[0]/NET0131  & ~\s3_msel_arb0_state_reg[1]/NET0131  ;
  assign n3103 = ~n3101 & n3102 ;
  assign n3104 = ~n3090 & ~n3103 ;
  assign n3105 = ~\s3_msel_arb0_state_reg[2]/NET0131  & n3085 ;
  assign n3106 = ~\s3_msel_arb0_state_reg[1]/NET0131  & ~\s3_msel_arb0_state_reg[2]/NET0131  ;
  assign n3107 = ~n3073 & n3106 ;
  assign n3108 = ~n3105 & ~n3107 ;
  assign n3109 = \s3_msel_arb0_state_reg[2]/NET0131  & n3074 ;
  assign n3110 = ~\s3_msel_arb0_state_reg[1]/NET0131  & \s3_msel_arb0_state_reg[2]/NET0131  ;
  assign n3111 = ~n3063 & n3110 ;
  assign n3112 = ~n3109 & ~n3111 ;
  assign n3113 = n3068 & n3084 ;
  assign n3114 = ~\s3_msel_arb0_state_reg[0]/NET0131  & ~n3113 ;
  assign n3115 = ~\s3_msel_arb0_state_reg[0]/NET0131  & n3063 ;
  assign n3116 = n3086 & n3115 ;
  assign n3117 = ~n3114 & ~n3116 ;
  assign n3118 = n3112 & ~n3117 ;
  assign n3119 = n3108 & n3118 ;
  assign n3120 = n3104 & ~n3119 ;
  assign n3121 = \m5_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[10]/NET0131  ;
  assign n3122 = ~\rf_conf4_reg[11]/NET0131  & n3121 ;
  assign n3123 = \m4_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[8]/NET0131  ;
  assign n3124 = ~\rf_conf4_reg[9]/NET0131  & n3123 ;
  assign n3125 = ~n3122 & ~n3124 ;
  assign n3126 = \m7_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[14]/NET0131  ;
  assign n3127 = ~\rf_conf4_reg[15]/NET0131  & n3126 ;
  assign n3128 = \m6_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[12]/NET0131  ;
  assign n3129 = ~\rf_conf4_reg[13]/NET0131  & n3128 ;
  assign n3130 = ~n3127 & ~n3129 ;
  assign n3131 = \m1_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[2]/NET0131  ;
  assign n3132 = ~\rf_conf4_reg[3]/NET0131  & n3131 ;
  assign n3133 = \m0_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[0]/NET0131  ;
  assign n3134 = ~\rf_conf4_reg[1]/NET0131  & n3133 ;
  assign n3135 = ~n3132 & ~n3134 ;
  assign n3136 = n3130 & ~n3135 ;
  assign n3137 = n3125 & ~n3136 ;
  assign n3138 = \m3_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[6]/NET0131  ;
  assign n3139 = ~\rf_conf4_reg[7]/NET0131  & n3138 ;
  assign n3140 = ~\s4_msel_arb0_state_reg[2]/NET0131  & ~n3139 ;
  assign n3141 = ~n3137 & n3140 ;
  assign n3142 = \s4_msel_arb0_state_reg[2]/NET0131  & ~n3127 ;
  assign n3143 = \s4_msel_arb0_state_reg[1]/NET0131  & ~n3142 ;
  assign n3144 = \m2_s4_cyc_o_reg/NET0131  & ~\rf_conf4_reg[4]/NET0131  ;
  assign n3145 = ~\rf_conf4_reg[5]/NET0131  & n3144 ;
  assign n3146 = ~n3139 & ~n3145 ;
  assign n3147 = ~n3125 & n3146 ;
  assign n3148 = \s4_msel_arb0_state_reg[1]/NET0131  & n3135 ;
  assign n3149 = ~n3147 & n3148 ;
  assign n3150 = ~n3143 & ~n3149 ;
  assign n3151 = ~n3141 & ~n3150 ;
  assign n3152 = \s4_msel_arb0_state_reg[0]/NET0131  & n3151 ;
  assign n3153 = \s4_msel_arb0_state_reg[2]/NET0131  & ~n3130 ;
  assign n3154 = ~n3122 & n3153 ;
  assign n3155 = ~n3124 & ~n3130 ;
  assign n3156 = ~n3134 & ~n3146 ;
  assign n3157 = ~n3155 & ~n3156 ;
  assign n3158 = ~n3122 & ~n3132 ;
  assign n3159 = ~n3157 & n3158 ;
  assign n3160 = ~n3154 & ~n3159 ;
  assign n3161 = ~\s4_msel_arb0_state_reg[2]/NET0131  & ~n3132 ;
  assign n3162 = ~n3146 & n3161 ;
  assign n3163 = n3160 & ~n3162 ;
  assign n3164 = \s4_msel_arb0_state_reg[0]/NET0131  & ~\s4_msel_arb0_state_reg[1]/NET0131  ;
  assign n3165 = ~n3163 & n3164 ;
  assign n3166 = ~n3152 & ~n3165 ;
  assign n3167 = ~\s4_msel_arb0_state_reg[2]/NET0131  & n3147 ;
  assign n3168 = ~\s4_msel_arb0_state_reg[1]/NET0131  & ~\s4_msel_arb0_state_reg[2]/NET0131  ;
  assign n3169 = ~n3135 & n3168 ;
  assign n3170 = ~n3167 & ~n3169 ;
  assign n3171 = \s4_msel_arb0_state_reg[2]/NET0131  & n3136 ;
  assign n3172 = ~\s4_msel_arb0_state_reg[1]/NET0131  & \s4_msel_arb0_state_reg[2]/NET0131  ;
  assign n3173 = ~n3125 & n3172 ;
  assign n3174 = ~n3171 & ~n3173 ;
  assign n3175 = n3130 & n3146 ;
  assign n3176 = ~\s4_msel_arb0_state_reg[0]/NET0131  & ~n3175 ;
  assign n3177 = ~\s4_msel_arb0_state_reg[0]/NET0131  & n3125 ;
  assign n3178 = n3148 & n3177 ;
  assign n3179 = ~n3176 & ~n3178 ;
  assign n3180 = n3174 & ~n3179 ;
  assign n3181 = n3170 & n3180 ;
  assign n3182 = n3166 & ~n3181 ;
  assign n3183 = \m5_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[10]/NET0131  ;
  assign n3184 = ~\rf_conf5_reg[11]/NET0131  & n3183 ;
  assign n3185 = \m4_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[8]/NET0131  ;
  assign n3186 = ~\rf_conf5_reg[9]/NET0131  & n3185 ;
  assign n3187 = ~n3184 & ~n3186 ;
  assign n3188 = \m7_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[14]/NET0131  ;
  assign n3189 = ~\rf_conf5_reg[15]/NET0131  & n3188 ;
  assign n3190 = \m6_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[12]/NET0131  ;
  assign n3191 = ~\rf_conf5_reg[13]/NET0131  & n3190 ;
  assign n3192 = ~n3189 & ~n3191 ;
  assign n3193 = \m1_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[2]/NET0131  ;
  assign n3194 = ~\rf_conf5_reg[3]/NET0131  & n3193 ;
  assign n3195 = \m0_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[0]/NET0131  ;
  assign n3196 = ~\rf_conf5_reg[1]/NET0131  & n3195 ;
  assign n3197 = ~n3194 & ~n3196 ;
  assign n3198 = n3192 & ~n3197 ;
  assign n3199 = n3187 & ~n3198 ;
  assign n3200 = \m3_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[6]/NET0131  ;
  assign n3201 = ~\rf_conf5_reg[7]/NET0131  & n3200 ;
  assign n3202 = ~\s5_msel_arb0_state_reg[2]/NET0131  & ~n3201 ;
  assign n3203 = ~n3199 & n3202 ;
  assign n3204 = \s5_msel_arb0_state_reg[2]/NET0131  & ~n3189 ;
  assign n3205 = \s5_msel_arb0_state_reg[1]/NET0131  & ~n3204 ;
  assign n3206 = \m2_s5_cyc_o_reg/NET0131  & ~\rf_conf5_reg[4]/NET0131  ;
  assign n3207 = ~\rf_conf5_reg[5]/NET0131  & n3206 ;
  assign n3208 = ~n3201 & ~n3207 ;
  assign n3209 = ~n3187 & n3208 ;
  assign n3210 = \s5_msel_arb0_state_reg[1]/NET0131  & n3197 ;
  assign n3211 = ~n3209 & n3210 ;
  assign n3212 = ~n3205 & ~n3211 ;
  assign n3213 = ~n3203 & ~n3212 ;
  assign n3214 = \s5_msel_arb0_state_reg[0]/NET0131  & n3213 ;
  assign n3215 = \s5_msel_arb0_state_reg[2]/NET0131  & ~n3192 ;
  assign n3216 = ~n3184 & n3215 ;
  assign n3217 = ~n3186 & ~n3192 ;
  assign n3218 = ~n3196 & ~n3208 ;
  assign n3219 = ~n3217 & ~n3218 ;
  assign n3220 = ~n3184 & ~n3194 ;
  assign n3221 = ~n3219 & n3220 ;
  assign n3222 = ~n3216 & ~n3221 ;
  assign n3223 = ~\s5_msel_arb0_state_reg[2]/NET0131  & ~n3194 ;
  assign n3224 = ~n3208 & n3223 ;
  assign n3225 = n3222 & ~n3224 ;
  assign n3226 = \s5_msel_arb0_state_reg[0]/NET0131  & ~\s5_msel_arb0_state_reg[1]/NET0131  ;
  assign n3227 = ~n3225 & n3226 ;
  assign n3228 = ~n3214 & ~n3227 ;
  assign n3229 = ~\s5_msel_arb0_state_reg[2]/NET0131  & n3209 ;
  assign n3230 = ~\s5_msel_arb0_state_reg[1]/NET0131  & ~\s5_msel_arb0_state_reg[2]/NET0131  ;
  assign n3231 = ~n3197 & n3230 ;
  assign n3232 = ~n3229 & ~n3231 ;
  assign n3233 = \s5_msel_arb0_state_reg[2]/NET0131  & n3198 ;
  assign n3234 = ~\s5_msel_arb0_state_reg[1]/NET0131  & \s5_msel_arb0_state_reg[2]/NET0131  ;
  assign n3235 = ~n3187 & n3234 ;
  assign n3236 = ~n3233 & ~n3235 ;
  assign n3237 = n3192 & n3208 ;
  assign n3238 = ~\s5_msel_arb0_state_reg[0]/NET0131  & ~n3237 ;
  assign n3239 = ~\s5_msel_arb0_state_reg[0]/NET0131  & n3187 ;
  assign n3240 = n3210 & n3239 ;
  assign n3241 = ~n3238 & ~n3240 ;
  assign n3242 = n3236 & ~n3241 ;
  assign n3243 = n3232 & n3242 ;
  assign n3244 = n3228 & ~n3243 ;
  assign n3245 = \m5_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[10]/NET0131  ;
  assign n3246 = ~\rf_conf6_reg[11]/NET0131  & n3245 ;
  assign n3247 = \m4_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[8]/NET0131  ;
  assign n3248 = ~\rf_conf6_reg[9]/NET0131  & n3247 ;
  assign n3249 = ~n3246 & ~n3248 ;
  assign n3250 = \m7_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[14]/NET0131  ;
  assign n3251 = ~\rf_conf6_reg[15]/NET0131  & n3250 ;
  assign n3252 = \m6_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[12]/NET0131  ;
  assign n3253 = ~\rf_conf6_reg[13]/NET0131  & n3252 ;
  assign n3254 = ~n3251 & ~n3253 ;
  assign n3255 = \m1_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[2]/NET0131  ;
  assign n3256 = ~\rf_conf6_reg[3]/NET0131  & n3255 ;
  assign n3257 = \m0_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[0]/NET0131  ;
  assign n3258 = ~\rf_conf6_reg[1]/NET0131  & n3257 ;
  assign n3259 = ~n3256 & ~n3258 ;
  assign n3260 = n3254 & ~n3259 ;
  assign n3261 = n3249 & ~n3260 ;
  assign n3262 = \m3_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[6]/NET0131  ;
  assign n3263 = ~\rf_conf6_reg[7]/NET0131  & n3262 ;
  assign n3264 = ~\s6_msel_arb0_state_reg[2]/NET0131  & ~n3263 ;
  assign n3265 = ~n3261 & n3264 ;
  assign n3266 = \s6_msel_arb0_state_reg[2]/NET0131  & ~n3251 ;
  assign n3267 = \s6_msel_arb0_state_reg[1]/NET0131  & ~n3266 ;
  assign n3268 = \m2_s6_cyc_o_reg/NET0131  & ~\rf_conf6_reg[4]/NET0131  ;
  assign n3269 = ~\rf_conf6_reg[5]/NET0131  & n3268 ;
  assign n3270 = ~n3263 & ~n3269 ;
  assign n3271 = ~n3249 & n3270 ;
  assign n3272 = \s6_msel_arb0_state_reg[1]/NET0131  & n3259 ;
  assign n3273 = ~n3271 & n3272 ;
  assign n3274 = ~n3267 & ~n3273 ;
  assign n3275 = ~n3265 & ~n3274 ;
  assign n3276 = \s6_msel_arb0_state_reg[0]/NET0131  & n3275 ;
  assign n3277 = \s6_msel_arb0_state_reg[2]/NET0131  & ~n3254 ;
  assign n3278 = ~n3246 & n3277 ;
  assign n3279 = ~n3248 & ~n3254 ;
  assign n3280 = ~n3258 & ~n3270 ;
  assign n3281 = ~n3279 & ~n3280 ;
  assign n3282 = ~n3246 & ~n3256 ;
  assign n3283 = ~n3281 & n3282 ;
  assign n3284 = ~n3278 & ~n3283 ;
  assign n3285 = ~\s6_msel_arb0_state_reg[2]/NET0131  & ~n3256 ;
  assign n3286 = ~n3270 & n3285 ;
  assign n3287 = n3284 & ~n3286 ;
  assign n3288 = \s6_msel_arb0_state_reg[0]/NET0131  & ~\s6_msel_arb0_state_reg[1]/NET0131  ;
  assign n3289 = ~n3287 & n3288 ;
  assign n3290 = ~n3276 & ~n3289 ;
  assign n3291 = ~\s6_msel_arb0_state_reg[2]/NET0131  & n3271 ;
  assign n3292 = ~\s6_msel_arb0_state_reg[1]/NET0131  & ~\s6_msel_arb0_state_reg[2]/NET0131  ;
  assign n3293 = ~n3259 & n3292 ;
  assign n3294 = ~n3291 & ~n3293 ;
  assign n3295 = \s6_msel_arb0_state_reg[2]/NET0131  & n3260 ;
  assign n3296 = ~\s6_msel_arb0_state_reg[1]/NET0131  & \s6_msel_arb0_state_reg[2]/NET0131  ;
  assign n3297 = ~n3249 & n3296 ;
  assign n3298 = ~n3295 & ~n3297 ;
  assign n3299 = n3254 & n3270 ;
  assign n3300 = ~\s6_msel_arb0_state_reg[0]/NET0131  & ~n3299 ;
  assign n3301 = ~\s6_msel_arb0_state_reg[0]/NET0131  & n3249 ;
  assign n3302 = n3272 & n3301 ;
  assign n3303 = ~n3300 & ~n3302 ;
  assign n3304 = n3298 & ~n3303 ;
  assign n3305 = n3294 & n3304 ;
  assign n3306 = n3290 & ~n3305 ;
  assign n3307 = \m5_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[10]/NET0131  ;
  assign n3308 = ~\rf_conf8_reg[11]/NET0131  & n3307 ;
  assign n3309 = \m4_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[8]/NET0131  ;
  assign n3310 = ~\rf_conf8_reg[9]/NET0131  & n3309 ;
  assign n3311 = ~n3308 & ~n3310 ;
  assign n3312 = \m7_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[14]/NET0131  ;
  assign n3313 = ~\rf_conf8_reg[15]/NET0131  & n3312 ;
  assign n3314 = \m6_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[12]/NET0131  ;
  assign n3315 = ~\rf_conf8_reg[13]/NET0131  & n3314 ;
  assign n3316 = ~n3313 & ~n3315 ;
  assign n3317 = \m1_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[2]/NET0131  ;
  assign n3318 = ~\rf_conf8_reg[3]/NET0131  & n3317 ;
  assign n3319 = \m0_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[0]/NET0131  ;
  assign n3320 = ~\rf_conf8_reg[1]/NET0131  & n3319 ;
  assign n3321 = ~n3318 & ~n3320 ;
  assign n3322 = n3316 & ~n3321 ;
  assign n3323 = n3311 & ~n3322 ;
  assign n3324 = \m3_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[6]/NET0131  ;
  assign n3325 = ~\rf_conf8_reg[7]/NET0131  & n3324 ;
  assign n3326 = ~\s8_msel_arb0_state_reg[2]/NET0131  & ~n3325 ;
  assign n3327 = ~n3323 & n3326 ;
  assign n3328 = \s8_msel_arb0_state_reg[2]/NET0131  & ~n3313 ;
  assign n3329 = \s8_msel_arb0_state_reg[1]/NET0131  & ~n3328 ;
  assign n3330 = \m2_s8_cyc_o_reg/NET0131  & ~\rf_conf8_reg[4]/NET0131  ;
  assign n3331 = ~\rf_conf8_reg[5]/NET0131  & n3330 ;
  assign n3332 = ~n3325 & ~n3331 ;
  assign n3333 = ~n3311 & n3332 ;
  assign n3334 = \s8_msel_arb0_state_reg[1]/NET0131  & n3321 ;
  assign n3335 = ~n3333 & n3334 ;
  assign n3336 = ~n3329 & ~n3335 ;
  assign n3337 = ~n3327 & ~n3336 ;
  assign n3338 = \s8_msel_arb0_state_reg[0]/NET0131  & n3337 ;
  assign n3339 = \s8_msel_arb0_state_reg[2]/NET0131  & ~n3316 ;
  assign n3340 = ~n3308 & n3339 ;
  assign n3341 = ~n3310 & ~n3316 ;
  assign n3342 = ~n3320 & ~n3332 ;
  assign n3343 = ~n3341 & ~n3342 ;
  assign n3344 = ~n3308 & ~n3318 ;
  assign n3345 = ~n3343 & n3344 ;
  assign n3346 = ~n3340 & ~n3345 ;
  assign n3347 = ~\s8_msel_arb0_state_reg[2]/NET0131  & ~n3318 ;
  assign n3348 = ~n3332 & n3347 ;
  assign n3349 = n3346 & ~n3348 ;
  assign n3350 = \s8_msel_arb0_state_reg[0]/NET0131  & ~\s8_msel_arb0_state_reg[1]/NET0131  ;
  assign n3351 = ~n3349 & n3350 ;
  assign n3352 = ~n3338 & ~n3351 ;
  assign n3353 = ~\s8_msel_arb0_state_reg[2]/NET0131  & n3333 ;
  assign n3354 = ~\s8_msel_arb0_state_reg[1]/NET0131  & ~\s8_msel_arb0_state_reg[2]/NET0131  ;
  assign n3355 = ~n3321 & n3354 ;
  assign n3356 = ~n3353 & ~n3355 ;
  assign n3357 = \s8_msel_arb0_state_reg[2]/NET0131  & n3322 ;
  assign n3358 = ~\s8_msel_arb0_state_reg[1]/NET0131  & \s8_msel_arb0_state_reg[2]/NET0131  ;
  assign n3359 = ~n3311 & n3358 ;
  assign n3360 = ~n3357 & ~n3359 ;
  assign n3361 = n3316 & n3332 ;
  assign n3362 = ~\s8_msel_arb0_state_reg[0]/NET0131  & ~n3361 ;
  assign n3363 = ~\s8_msel_arb0_state_reg[0]/NET0131  & n3311 ;
  assign n3364 = n3334 & n3363 ;
  assign n3365 = ~n3362 & ~n3364 ;
  assign n3366 = n3360 & ~n3365 ;
  assign n3367 = n3356 & n3366 ;
  assign n3368 = n3352 & ~n3367 ;
  assign n3369 = \m3_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[6]/NET0131  ;
  assign n3370 = ~\rf_conf1_reg[7]/NET0131  & n3369 ;
  assign n3371 = \m2_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[4]/NET0131  ;
  assign n3372 = ~\rf_conf1_reg[5]/NET0131  & n3371 ;
  assign n3373 = ~n3370 & ~n3372 ;
  assign n3374 = \m4_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[8]/NET0131  ;
  assign n3375 = ~\rf_conf1_reg[9]/NET0131  & n3374 ;
  assign n3376 = \m5_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[10]/NET0131  ;
  assign n3377 = ~\rf_conf1_reg[11]/NET0131  & n3376 ;
  assign n3378 = ~n3375 & ~n3377 ;
  assign n3379 = \m7_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[14]/NET0131  ;
  assign n3380 = ~\rf_conf1_reg[15]/NET0131  & n3379 ;
  assign n3381 = \m6_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[12]/NET0131  ;
  assign n3382 = ~\rf_conf1_reg[13]/NET0131  & n3381 ;
  assign n3383 = ~n3380 & ~n3382 ;
  assign n3384 = n3378 & ~n3383 ;
  assign n3385 = n3373 & ~n3384 ;
  assign n3386 = \m1_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[2]/NET0131  ;
  assign n3387 = ~\rf_conf1_reg[3]/NET0131  & n3386 ;
  assign n3388 = \m0_s1_cyc_o_reg/NET0131  & ~\rf_conf1_reg[0]/NET0131  ;
  assign n3389 = ~\rf_conf1_reg[1]/NET0131  & n3388 ;
  assign n3390 = ~n3387 & ~n3389 ;
  assign n3391 = ~\s1_msel_arb0_state_reg[1]/NET0131  & ~n3390 ;
  assign n3392 = ~\s1_msel_arb0_state_reg[2]/NET0131  & ~n3391 ;
  assign n3393 = ~n3385 & n3392 ;
  assign n3394 = \s1_msel_arb0_state_reg[2]/NET0131  & ~n3383 ;
  assign n3395 = \s1_msel_arb0_state_reg[1]/NET0131  & n3394 ;
  assign n3396 = n3373 & ~n3378 ;
  assign n3397 = \s1_msel_arb0_state_reg[1]/NET0131  & n3390 ;
  assign n3398 = ~n3396 & n3397 ;
  assign n3399 = ~n3395 & ~n3398 ;
  assign n3400 = ~n3393 & n3399 ;
  assign n3401 = ~\s1_msel_arb0_state_reg[0]/NET0131  & ~n3400 ;
  assign n3402 = \s1_msel_arb0_state_reg[0]/NET0131  & ~n3387 ;
  assign n3403 = ~\s1_msel_arb0_state_reg[2]/NET0131  & n3402 ;
  assign n3404 = ~n3385 & n3403 ;
  assign n3405 = ~\s1_msel_arb0_state_reg[1]/NET0131  & n3404 ;
  assign n3406 = ~\s1_msel_arb0_state_reg[0]/NET0131  & \s1_msel_arb0_state_reg[1]/NET0131  ;
  assign n3407 = n3373 & ~n3406 ;
  assign n3408 = n3390 & ~n3407 ;
  assign n3409 = n3383 & ~n3408 ;
  assign n3410 = ~\rf_conf1_reg[9]/NET0131  & ~\s1_msel_arb0_state_reg[0]/NET0131  ;
  assign n3411 = n3374 & n3410 ;
  assign n3412 = ~n3377 & ~n3411 ;
  assign n3413 = \s1_msel_arb0_state_reg[2]/NET0131  & n3412 ;
  assign n3414 = ~\s1_msel_arb0_state_reg[1]/NET0131  & n3413 ;
  assign n3415 = ~n3409 & n3414 ;
  assign n3416 = ~n3405 & ~n3415 ;
  assign n3417 = \s1_msel_arb0_state_reg[1]/NET0131  & ~\s1_msel_arb0_state_reg[2]/NET0131  ;
  assign n3418 = n3370 & n3417 ;
  assign n3419 = n3383 & ~n3390 ;
  assign n3420 = n3378 & n3417 ;
  assign n3421 = ~n3419 & n3420 ;
  assign n3422 = ~n3418 & ~n3421 ;
  assign n3423 = \s1_msel_arb0_state_reg[1]/NET0131  & \s1_msel_arb0_state_reg[2]/NET0131  ;
  assign n3424 = n3380 & n3423 ;
  assign n3425 = n3390 & n3423 ;
  assign n3426 = ~n3396 & n3425 ;
  assign n3427 = ~n3424 & ~n3426 ;
  assign n3428 = n3422 & n3427 ;
  assign n3429 = \s1_msel_arb0_state_reg[0]/NET0131  & ~n3428 ;
  assign n3430 = n3416 & ~n3429 ;
  assign n3431 = ~n3401 & n3430 ;
  assign n3432 = \m3_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[6]/NET0131  ;
  assign n3433 = ~\rf_conf2_reg[7]/NET0131  & n3432 ;
  assign n3434 = \m2_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[4]/NET0131  ;
  assign n3435 = ~\rf_conf2_reg[5]/NET0131  & n3434 ;
  assign n3436 = ~n3433 & ~n3435 ;
  assign n3437 = \m4_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[8]/NET0131  ;
  assign n3438 = ~\rf_conf2_reg[9]/NET0131  & n3437 ;
  assign n3439 = \m5_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[10]/NET0131  ;
  assign n3440 = ~\rf_conf2_reg[11]/NET0131  & n3439 ;
  assign n3441 = ~n3438 & ~n3440 ;
  assign n3442 = \m7_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[14]/NET0131  ;
  assign n3443 = ~\rf_conf2_reg[15]/NET0131  & n3442 ;
  assign n3444 = \m6_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[12]/NET0131  ;
  assign n3445 = ~\rf_conf2_reg[13]/NET0131  & n3444 ;
  assign n3446 = ~n3443 & ~n3445 ;
  assign n3447 = n3441 & ~n3446 ;
  assign n3448 = n3436 & ~n3447 ;
  assign n3449 = \m1_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[2]/NET0131  ;
  assign n3450 = ~\rf_conf2_reg[3]/NET0131  & n3449 ;
  assign n3451 = \m0_s2_cyc_o_reg/NET0131  & ~\rf_conf2_reg[0]/NET0131  ;
  assign n3452 = ~\rf_conf2_reg[1]/NET0131  & n3451 ;
  assign n3453 = ~n3450 & ~n3452 ;
  assign n3454 = ~\s2_msel_arb0_state_reg[1]/NET0131  & ~n3453 ;
  assign n3455 = ~\s2_msel_arb0_state_reg[2]/NET0131  & ~n3454 ;
  assign n3456 = ~n3448 & n3455 ;
  assign n3457 = \s2_msel_arb0_state_reg[2]/NET0131  & ~n3446 ;
  assign n3458 = \s2_msel_arb0_state_reg[1]/NET0131  & n3457 ;
  assign n3459 = n3436 & ~n3441 ;
  assign n3460 = \s2_msel_arb0_state_reg[1]/NET0131  & n3453 ;
  assign n3461 = ~n3459 & n3460 ;
  assign n3462 = ~n3458 & ~n3461 ;
  assign n3463 = ~n3456 & n3462 ;
  assign n3464 = ~\s2_msel_arb0_state_reg[0]/NET0131  & ~n3463 ;
  assign n3465 = \s2_msel_arb0_state_reg[0]/NET0131  & ~n3450 ;
  assign n3466 = ~\s2_msel_arb0_state_reg[2]/NET0131  & n3465 ;
  assign n3467 = ~n3448 & n3466 ;
  assign n3468 = ~\s2_msel_arb0_state_reg[1]/NET0131  & n3467 ;
  assign n3469 = ~\s2_msel_arb0_state_reg[0]/NET0131  & \s2_msel_arb0_state_reg[1]/NET0131  ;
  assign n3470 = n3436 & ~n3469 ;
  assign n3471 = n3453 & ~n3470 ;
  assign n3472 = n3446 & ~n3471 ;
  assign n3473 = ~\rf_conf2_reg[9]/NET0131  & ~\s2_msel_arb0_state_reg[0]/NET0131  ;
  assign n3474 = n3437 & n3473 ;
  assign n3475 = ~n3440 & ~n3474 ;
  assign n3476 = \s2_msel_arb0_state_reg[2]/NET0131  & n3475 ;
  assign n3477 = ~\s2_msel_arb0_state_reg[1]/NET0131  & n3476 ;
  assign n3478 = ~n3472 & n3477 ;
  assign n3479 = ~n3468 & ~n3478 ;
  assign n3480 = \s2_msel_arb0_state_reg[1]/NET0131  & ~\s2_msel_arb0_state_reg[2]/NET0131  ;
  assign n3481 = n3433 & n3480 ;
  assign n3482 = n3446 & ~n3453 ;
  assign n3483 = n3441 & n3480 ;
  assign n3484 = ~n3482 & n3483 ;
  assign n3485 = ~n3481 & ~n3484 ;
  assign n3486 = \s2_msel_arb0_state_reg[1]/NET0131  & \s2_msel_arb0_state_reg[2]/NET0131  ;
  assign n3487 = n3443 & n3486 ;
  assign n3488 = n3453 & n3486 ;
  assign n3489 = ~n3459 & n3488 ;
  assign n3490 = ~n3487 & ~n3489 ;
  assign n3491 = n3485 & n3490 ;
  assign n3492 = \s2_msel_arb0_state_reg[0]/NET0131  & ~n3491 ;
  assign n3493 = n3479 & ~n3492 ;
  assign n3494 = ~n3464 & n3493 ;
  assign n3495 = \m3_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[6]/NET0131  ;
  assign n3496 = ~\rf_conf7_reg[7]/NET0131  & n3495 ;
  assign n3497 = \m2_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[4]/NET0131  ;
  assign n3498 = ~\rf_conf7_reg[5]/NET0131  & n3497 ;
  assign n3499 = ~n3496 & ~n3498 ;
  assign n3500 = \m4_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[8]/NET0131  ;
  assign n3501 = ~\rf_conf7_reg[9]/NET0131  & n3500 ;
  assign n3502 = \m5_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[10]/NET0131  ;
  assign n3503 = ~\rf_conf7_reg[11]/NET0131  & n3502 ;
  assign n3504 = ~n3501 & ~n3503 ;
  assign n3505 = \m7_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[14]/NET0131  ;
  assign n3506 = ~\rf_conf7_reg[15]/NET0131  & n3505 ;
  assign n3507 = \m6_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[12]/NET0131  ;
  assign n3508 = ~\rf_conf7_reg[13]/NET0131  & n3507 ;
  assign n3509 = ~n3506 & ~n3508 ;
  assign n3510 = n3504 & ~n3509 ;
  assign n3511 = n3499 & ~n3510 ;
  assign n3512 = \m1_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[2]/NET0131  ;
  assign n3513 = ~\rf_conf7_reg[3]/NET0131  & n3512 ;
  assign n3514 = \m0_s7_cyc_o_reg/NET0131  & ~\rf_conf7_reg[0]/NET0131  ;
  assign n3515 = ~\rf_conf7_reg[1]/NET0131  & n3514 ;
  assign n3516 = ~n3513 & ~n3515 ;
  assign n3517 = ~\s7_msel_arb0_state_reg[1]/NET0131  & ~n3516 ;
  assign n3518 = ~\s7_msel_arb0_state_reg[2]/NET0131  & ~n3517 ;
  assign n3519 = ~n3511 & n3518 ;
  assign n3520 = \s7_msel_arb0_state_reg[2]/NET0131  & ~n3509 ;
  assign n3521 = \s7_msel_arb0_state_reg[1]/NET0131  & n3520 ;
  assign n3522 = n3499 & ~n3504 ;
  assign n3523 = \s7_msel_arb0_state_reg[1]/NET0131  & n3516 ;
  assign n3524 = ~n3522 & n3523 ;
  assign n3525 = ~n3521 & ~n3524 ;
  assign n3526 = ~n3519 & n3525 ;
  assign n3527 = ~\s7_msel_arb0_state_reg[0]/NET0131  & ~n3526 ;
  assign n3528 = \s7_msel_arb0_state_reg[0]/NET0131  & ~n3513 ;
  assign n3529 = ~\s7_msel_arb0_state_reg[2]/NET0131  & n3528 ;
  assign n3530 = ~n3511 & n3529 ;
  assign n3531 = ~\s7_msel_arb0_state_reg[1]/NET0131  & n3530 ;
  assign n3532 = ~\s7_msel_arb0_state_reg[0]/NET0131  & \s7_msel_arb0_state_reg[1]/NET0131  ;
  assign n3533 = n3499 & ~n3532 ;
  assign n3534 = n3516 & ~n3533 ;
  assign n3535 = n3509 & ~n3534 ;
  assign n3536 = ~\rf_conf7_reg[9]/NET0131  & ~\s7_msel_arb0_state_reg[0]/NET0131  ;
  assign n3537 = n3500 & n3536 ;
  assign n3538 = ~n3503 & ~n3537 ;
  assign n3539 = \s7_msel_arb0_state_reg[2]/NET0131  & n3538 ;
  assign n3540 = ~\s7_msel_arb0_state_reg[1]/NET0131  & n3539 ;
  assign n3541 = ~n3535 & n3540 ;
  assign n3542 = ~n3531 & ~n3541 ;
  assign n3543 = \s7_msel_arb0_state_reg[1]/NET0131  & ~\s7_msel_arb0_state_reg[2]/NET0131  ;
  assign n3544 = n3496 & n3543 ;
  assign n3545 = n3509 & ~n3516 ;
  assign n3546 = n3504 & n3543 ;
  assign n3547 = ~n3545 & n3546 ;
  assign n3548 = ~n3544 & ~n3547 ;
  assign n3549 = \s7_msel_arb0_state_reg[1]/NET0131  & \s7_msel_arb0_state_reg[2]/NET0131  ;
  assign n3550 = n3506 & n3549 ;
  assign n3551 = n3516 & n3549 ;
  assign n3552 = ~n3522 & n3551 ;
  assign n3553 = ~n3550 & ~n3552 ;
  assign n3554 = n3548 & n3553 ;
  assign n3555 = \s7_msel_arb0_state_reg[0]/NET0131  & ~n3554 ;
  assign n3556 = n3542 & ~n3555 ;
  assign n3557 = ~n3527 & n3556 ;
  assign n3558 = \m3_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[6]/NET0131  ;
  assign n3559 = ~\rf_conf9_reg[7]/NET0131  & n3558 ;
  assign n3560 = \m2_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[4]/NET0131  ;
  assign n3561 = ~\rf_conf9_reg[5]/NET0131  & n3560 ;
  assign n3562 = ~n3559 & ~n3561 ;
  assign n3563 = \m4_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[8]/NET0131  ;
  assign n3564 = ~\rf_conf9_reg[9]/NET0131  & n3563 ;
  assign n3565 = \m5_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[10]/NET0131  ;
  assign n3566 = ~\rf_conf9_reg[11]/NET0131  & n3565 ;
  assign n3567 = ~n3564 & ~n3566 ;
  assign n3568 = \m7_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[14]/NET0131  ;
  assign n3569 = ~\rf_conf9_reg[15]/NET0131  & n3568 ;
  assign n3570 = \m6_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[12]/NET0131  ;
  assign n3571 = ~\rf_conf9_reg[13]/NET0131  & n3570 ;
  assign n3572 = ~n3569 & ~n3571 ;
  assign n3573 = n3567 & ~n3572 ;
  assign n3574 = n3562 & ~n3573 ;
  assign n3575 = \m1_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[2]/NET0131  ;
  assign n3576 = ~\rf_conf9_reg[3]/NET0131  & n3575 ;
  assign n3577 = \m0_s9_cyc_o_reg/NET0131  & ~\rf_conf9_reg[0]/NET0131  ;
  assign n3578 = ~\rf_conf9_reg[1]/NET0131  & n3577 ;
  assign n3579 = ~n3576 & ~n3578 ;
  assign n3580 = ~\s9_msel_arb0_state_reg[1]/NET0131  & ~n3579 ;
  assign n3581 = ~\s9_msel_arb0_state_reg[2]/NET0131  & ~n3580 ;
  assign n3582 = ~n3574 & n3581 ;
  assign n3583 = \s9_msel_arb0_state_reg[2]/NET0131  & ~n3572 ;
  assign n3584 = \s9_msel_arb0_state_reg[1]/NET0131  & n3583 ;
  assign n3585 = n3562 & ~n3567 ;
  assign n3586 = \s9_msel_arb0_state_reg[1]/NET0131  & n3579 ;
  assign n3587 = ~n3585 & n3586 ;
  assign n3588 = ~n3584 & ~n3587 ;
  assign n3589 = ~n3582 & n3588 ;
  assign n3590 = ~\s9_msel_arb0_state_reg[0]/NET0131  & ~n3589 ;
  assign n3591 = \s9_msel_arb0_state_reg[0]/NET0131  & ~n3576 ;
  assign n3592 = ~\s9_msel_arb0_state_reg[2]/NET0131  & n3591 ;
  assign n3593 = ~n3574 & n3592 ;
  assign n3594 = ~\s9_msel_arb0_state_reg[1]/NET0131  & n3593 ;
  assign n3595 = ~\s9_msel_arb0_state_reg[0]/NET0131  & \s9_msel_arb0_state_reg[1]/NET0131  ;
  assign n3596 = n3562 & ~n3595 ;
  assign n3597 = n3579 & ~n3596 ;
  assign n3598 = n3572 & ~n3597 ;
  assign n3599 = ~\rf_conf9_reg[9]/NET0131  & ~\s9_msel_arb0_state_reg[0]/NET0131  ;
  assign n3600 = n3563 & n3599 ;
  assign n3601 = ~n3566 & ~n3600 ;
  assign n3602 = \s9_msel_arb0_state_reg[2]/NET0131  & n3601 ;
  assign n3603 = ~\s9_msel_arb0_state_reg[1]/NET0131  & n3602 ;
  assign n3604 = ~n3598 & n3603 ;
  assign n3605 = ~n3594 & ~n3604 ;
  assign n3606 = \s9_msel_arb0_state_reg[1]/NET0131  & ~\s9_msel_arb0_state_reg[2]/NET0131  ;
  assign n3607 = n3559 & n3606 ;
  assign n3608 = n3572 & ~n3579 ;
  assign n3609 = n3567 & n3606 ;
  assign n3610 = ~n3608 & n3609 ;
  assign n3611 = ~n3607 & ~n3610 ;
  assign n3612 = \s9_msel_arb0_state_reg[1]/NET0131  & \s9_msel_arb0_state_reg[2]/NET0131  ;
  assign n3613 = n3569 & n3612 ;
  assign n3614 = n3579 & n3612 ;
  assign n3615 = ~n3585 & n3614 ;
  assign n3616 = ~n3613 & ~n3615 ;
  assign n3617 = n3611 & n3616 ;
  assign n3618 = \s9_msel_arb0_state_reg[0]/NET0131  & ~n3617 ;
  assign n3619 = n3605 & ~n3618 ;
  assign n3620 = ~n3590 & n3619 ;
  assign n3621 = \m3_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[6]/NET0131  ;
  assign n3622 = ~\rf_conf0_reg[7]/NET0131  & n3621 ;
  assign n3623 = \m2_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[4]/NET0131  ;
  assign n3624 = ~\rf_conf0_reg[5]/NET0131  & n3623 ;
  assign n3625 = ~n3622 & ~n3624 ;
  assign n3626 = \m4_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[8]/NET0131  ;
  assign n3627 = ~\rf_conf0_reg[9]/NET0131  & n3626 ;
  assign n3628 = \m5_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[10]/NET0131  ;
  assign n3629 = ~\rf_conf0_reg[11]/NET0131  & n3628 ;
  assign n3630 = ~n3627 & ~n3629 ;
  assign n3631 = \m7_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[14]/NET0131  ;
  assign n3632 = ~\rf_conf0_reg[15]/NET0131  & n3631 ;
  assign n3633 = \m6_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[12]/NET0131  ;
  assign n3634 = ~\rf_conf0_reg[13]/NET0131  & n3633 ;
  assign n3635 = ~n3632 & ~n3634 ;
  assign n3636 = n3630 & ~n3635 ;
  assign n3637 = n3625 & ~n3636 ;
  assign n3638 = \m1_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[2]/NET0131  ;
  assign n3639 = ~\rf_conf0_reg[3]/NET0131  & n3638 ;
  assign n3640 = \m0_s0_cyc_o_reg/NET0131  & ~\rf_conf0_reg[0]/NET0131  ;
  assign n3641 = ~\rf_conf0_reg[1]/NET0131  & n3640 ;
  assign n3642 = ~n3639 & ~n3641 ;
  assign n3643 = ~\s0_msel_arb0_state_reg[1]/NET0131  & ~n3642 ;
  assign n3644 = ~\s0_msel_arb0_state_reg[2]/NET0131  & ~n3643 ;
  assign n3645 = ~n3637 & n3644 ;
  assign n3646 = \s0_msel_arb0_state_reg[2]/NET0131  & ~n3635 ;
  assign n3647 = \s0_msel_arb0_state_reg[1]/NET0131  & n3646 ;
  assign n3648 = n3625 & ~n3630 ;
  assign n3649 = \s0_msel_arb0_state_reg[1]/NET0131  & n3642 ;
  assign n3650 = ~n3648 & n3649 ;
  assign n3651 = ~n3647 & ~n3650 ;
  assign n3652 = ~n3645 & n3651 ;
  assign n3653 = ~\s0_msel_arb0_state_reg[0]/NET0131  & ~n3652 ;
  assign n3654 = \s0_msel_arb0_state_reg[0]/NET0131  & ~n3639 ;
  assign n3655 = ~\s0_msel_arb0_state_reg[2]/NET0131  & n3654 ;
  assign n3656 = ~n3637 & n3655 ;
  assign n3657 = ~\s0_msel_arb0_state_reg[1]/NET0131  & n3656 ;
  assign n3658 = ~\s0_msel_arb0_state_reg[0]/NET0131  & \s0_msel_arb0_state_reg[1]/NET0131  ;
  assign n3659 = n3625 & ~n3658 ;
  assign n3660 = n3642 & ~n3659 ;
  assign n3661 = n3635 & ~n3660 ;
  assign n3662 = ~\rf_conf0_reg[9]/NET0131  & ~\s0_msel_arb0_state_reg[0]/NET0131  ;
  assign n3663 = n3626 & n3662 ;
  assign n3664 = ~n3629 & ~n3663 ;
  assign n3665 = \s0_msel_arb0_state_reg[2]/NET0131  & n3664 ;
  assign n3666 = ~\s0_msel_arb0_state_reg[1]/NET0131  & n3665 ;
  assign n3667 = ~n3661 & n3666 ;
  assign n3668 = ~n3657 & ~n3667 ;
  assign n3669 = \s0_msel_arb0_state_reg[1]/NET0131  & ~\s0_msel_arb0_state_reg[2]/NET0131  ;
  assign n3670 = n3622 & n3669 ;
  assign n3671 = n3635 & ~n3642 ;
  assign n3672 = n3630 & n3669 ;
  assign n3673 = ~n3671 & n3672 ;
  assign n3674 = ~n3670 & ~n3673 ;
  assign n3675 = \s0_msel_arb0_state_reg[1]/NET0131  & \s0_msel_arb0_state_reg[2]/NET0131  ;
  assign n3676 = n3632 & n3675 ;
  assign n3677 = n3642 & n3675 ;
  assign n3678 = ~n3648 & n3677 ;
  assign n3679 = ~n3676 & ~n3678 ;
  assign n3680 = n3674 & n3679 ;
  assign n3681 = \s0_msel_arb0_state_reg[0]/NET0131  & ~n3680 ;
  assign n3682 = n3668 & ~n3681 ;
  assign n3683 = ~n3653 & n3682 ;
  assign n3684 = \m3_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[6]/NET0131  ;
  assign n3685 = ~\rf_conf10_reg[7]/NET0131  & n3684 ;
  assign n3686 = \m2_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[4]/NET0131  ;
  assign n3687 = ~\rf_conf10_reg[5]/NET0131  & n3686 ;
  assign n3688 = ~n3685 & ~n3687 ;
  assign n3689 = \m4_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[8]/NET0131  ;
  assign n3690 = ~\rf_conf10_reg[9]/NET0131  & n3689 ;
  assign n3691 = \m5_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[10]/NET0131  ;
  assign n3692 = ~\rf_conf10_reg[11]/NET0131  & n3691 ;
  assign n3693 = ~n3690 & ~n3692 ;
  assign n3694 = \m7_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[14]/NET0131  ;
  assign n3695 = ~\rf_conf10_reg[15]/NET0131  & n3694 ;
  assign n3696 = \m6_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[12]/NET0131  ;
  assign n3697 = ~\rf_conf10_reg[13]/NET0131  & n3696 ;
  assign n3698 = ~n3695 & ~n3697 ;
  assign n3699 = n3693 & ~n3698 ;
  assign n3700 = n3688 & ~n3699 ;
  assign n3701 = \m1_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[2]/NET0131  ;
  assign n3702 = ~\rf_conf10_reg[3]/NET0131  & n3701 ;
  assign n3703 = \m0_s10_cyc_o_reg/NET0131  & ~\rf_conf10_reg[0]/NET0131  ;
  assign n3704 = ~\rf_conf10_reg[1]/NET0131  & n3703 ;
  assign n3705 = ~n3702 & ~n3704 ;
  assign n3706 = ~\s10_msel_arb0_state_reg[1]/NET0131  & ~n3705 ;
  assign n3707 = ~\s10_msel_arb0_state_reg[2]/NET0131  & ~n3706 ;
  assign n3708 = ~n3700 & n3707 ;
  assign n3709 = \s10_msel_arb0_state_reg[2]/NET0131  & ~n3698 ;
  assign n3710 = \s10_msel_arb0_state_reg[1]/NET0131  & n3709 ;
  assign n3711 = n3688 & ~n3693 ;
  assign n3712 = \s10_msel_arb0_state_reg[1]/NET0131  & n3705 ;
  assign n3713 = ~n3711 & n3712 ;
  assign n3714 = ~n3710 & ~n3713 ;
  assign n3715 = ~n3708 & n3714 ;
  assign n3716 = ~\s10_msel_arb0_state_reg[0]/NET0131  & ~n3715 ;
  assign n3717 = \s10_msel_arb0_state_reg[0]/NET0131  & ~n3702 ;
  assign n3718 = ~\s10_msel_arb0_state_reg[2]/NET0131  & n3717 ;
  assign n3719 = ~n3700 & n3718 ;
  assign n3720 = ~\s10_msel_arb0_state_reg[1]/NET0131  & n3719 ;
  assign n3721 = ~\s10_msel_arb0_state_reg[0]/NET0131  & \s10_msel_arb0_state_reg[1]/NET0131  ;
  assign n3722 = n3688 & ~n3721 ;
  assign n3723 = n3705 & ~n3722 ;
  assign n3724 = n3698 & ~n3723 ;
  assign n3725 = ~\rf_conf10_reg[9]/NET0131  & ~\s10_msel_arb0_state_reg[0]/NET0131  ;
  assign n3726 = n3689 & n3725 ;
  assign n3727 = ~n3692 & ~n3726 ;
  assign n3728 = \s10_msel_arb0_state_reg[2]/NET0131  & n3727 ;
  assign n3729 = ~\s10_msel_arb0_state_reg[1]/NET0131  & n3728 ;
  assign n3730 = ~n3724 & n3729 ;
  assign n3731 = ~n3720 & ~n3730 ;
  assign n3732 = \s10_msel_arb0_state_reg[1]/NET0131  & ~\s10_msel_arb0_state_reg[2]/NET0131  ;
  assign n3733 = n3685 & n3732 ;
  assign n3734 = n3698 & ~n3705 ;
  assign n3735 = n3693 & n3732 ;
  assign n3736 = ~n3734 & n3735 ;
  assign n3737 = ~n3733 & ~n3736 ;
  assign n3738 = \s10_msel_arb0_state_reg[1]/NET0131  & \s10_msel_arb0_state_reg[2]/NET0131  ;
  assign n3739 = n3695 & n3738 ;
  assign n3740 = n3705 & n3738 ;
  assign n3741 = ~n3711 & n3740 ;
  assign n3742 = ~n3739 & ~n3741 ;
  assign n3743 = n3737 & n3742 ;
  assign n3744 = \s10_msel_arb0_state_reg[0]/NET0131  & ~n3743 ;
  assign n3745 = n3731 & ~n3744 ;
  assign n3746 = ~n3716 & n3745 ;
  assign n3747 = \m3_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[6]/NET0131  ;
  assign n3748 = ~\rf_conf15_reg[7]/NET0131  & n3747 ;
  assign n3749 = \m2_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[4]/NET0131  ;
  assign n3750 = ~\rf_conf15_reg[5]/NET0131  & n3749 ;
  assign n3751 = ~n3748 & ~n3750 ;
  assign n3752 = \m0_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[0]/NET0131  ;
  assign n3753 = ~\rf_conf15_reg[1]/NET0131  & n3752 ;
  assign n3754 = \m1_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[2]/NET0131  ;
  assign n3755 = ~\rf_conf15_reg[3]/NET0131  & n3754 ;
  assign n3756 = ~n3753 & ~n3755 ;
  assign n3757 = n3751 & n3756 ;
  assign n3758 = \m6_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[12]/NET0131  ;
  assign n3759 = ~\rf_conf15_reg[13]/NET0131  & n3758 ;
  assign n3760 = \m7_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[14]/NET0131  ;
  assign n3761 = ~\rf_conf15_reg[15]/NET0131  & n3760 ;
  assign n3762 = ~n3759 & ~n3761 ;
  assign n3763 = \m5_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[10]/NET0131  ;
  assign n3764 = ~\rf_conf15_reg[11]/NET0131  & n3763 ;
  assign n3765 = \m4_s15_cyc_o_reg/NET0131  & \rf_conf15_reg[8]/NET0131  ;
  assign n3766 = ~\rf_conf15_reg[9]/NET0131  & n3765 ;
  assign n3767 = ~n3764 & ~n3766 ;
  assign n3768 = n3762 & n3767 ;
  assign n3769 = n3757 & n3768 ;
  assign n3770 = \rf_conf15_reg[7]/NET0131  & n3001 ;
  assign n3771 = \rf_conf15_reg[5]/NET0131  & n3003 ;
  assign n3772 = ~n3770 & ~n3771 ;
  assign n3773 = \rf_conf15_reg[1]/NET0131  & n3009 ;
  assign n3774 = \rf_conf15_reg[3]/NET0131  & n3007 ;
  assign n3775 = ~n3773 & ~n3774 ;
  assign n3776 = n3772 & n3775 ;
  assign n3777 = \rf_conf15_reg[9]/NET0131  & n2990 ;
  assign n3778 = \rf_conf15_reg[11]/NET0131  & n2988 ;
  assign n3779 = ~n3777 & ~n3778 ;
  assign n3780 = \rf_conf15_reg[15]/NET0131  & n2995 ;
  assign n3781 = \rf_conf15_reg[13]/NET0131  & n2993 ;
  assign n3782 = ~n3780 & ~n3781 ;
  assign n3783 = n3779 & n3782 ;
  assign n3784 = \s15_next_reg/P0001  & n3783 ;
  assign n3785 = n3776 & n3784 ;
  assign n3786 = ~n3769 & n3785 ;
  assign n3787 = \s15_msel_pri_out_reg[0]/NET0131  & ~\s15_next_reg/P0001  ;
  assign n3788 = \rf_conf15_reg[7]/NET0131  & n3747 ;
  assign n3789 = \rf_conf15_reg[5]/NET0131  & n3749 ;
  assign n3790 = ~n3788 & ~n3789 ;
  assign n3791 = \rf_conf15_reg[1]/NET0131  & n3752 ;
  assign n3792 = \rf_conf15_reg[3]/NET0131  & n3754 ;
  assign n3793 = ~n3791 & ~n3792 ;
  assign n3794 = n3790 & n3793 ;
  assign n3795 = \rf_conf15_reg[15]/NET0131  & n3760 ;
  assign n3796 = \rf_conf15_reg[13]/NET0131  & n3758 ;
  assign n3797 = ~n3795 & ~n3796 ;
  assign n3798 = \rf_conf15_reg[9]/NET0131  & n3765 ;
  assign n3799 = \rf_conf15_reg[11]/NET0131  & n3763 ;
  assign n3800 = ~n3798 & ~n3799 ;
  assign n3801 = n3797 & n3800 ;
  assign n3802 = n3794 & n3801 ;
  assign n3803 = \s15_next_reg/P0001  & ~n3802 ;
  assign n3804 = ~n3787 & ~n3803 ;
  assign n3805 = ~n3786 & n3804 ;
  assign n3806 = ~rst_i_pad & ~n3805 ;
  assign n3807 = ~\s15_msel_arb3_state_reg[0]/NET0131  & ~\s15_msel_arb3_state_reg[1]/NET0131  ;
  assign n3808 = n3794 & n3807 ;
  assign n3809 = \rf_conf15_reg[3]/NET0131  & ~\s15_msel_arb3_state_reg[1]/NET0131  ;
  assign n3810 = n3754 & n3809 ;
  assign n3811 = ~n3807 & ~n3810 ;
  assign n3812 = \s15_msel_arb3_state_reg[0]/NET0131  & \s15_msel_arb3_state_reg[1]/NET0131  ;
  assign n3813 = n3789 & ~n3812 ;
  assign n3814 = ~\s15_msel_arb3_state_reg[2]/NET0131  & ~n3788 ;
  assign n3815 = ~n3813 & n3814 ;
  assign n3816 = n3811 & n3815 ;
  assign n3817 = ~n3808 & ~n3816 ;
  assign n3818 = ~n3801 & ~n3817 ;
  assign n3819 = ~\s15_msel_arb3_state_reg[1]/NET0131  & n3799 ;
  assign n3820 = n3798 & n3807 ;
  assign n3821 = ~n3819 & ~n3820 ;
  assign n3822 = n3796 & ~n3812 ;
  assign n3823 = ~n3795 & ~n3822 ;
  assign n3824 = ~n3794 & n3823 ;
  assign n3825 = n3821 & n3824 ;
  assign n3826 = \s15_msel_arb3_state_reg[2]/NET0131  & ~n3825 ;
  assign n3827 = ~n3818 & ~n3826 ;
  assign n3828 = ~\s15_msel_arb1_state_reg[1]/NET0131  & n3755 ;
  assign n3829 = ~\s15_msel_arb1_state_reg[0]/NET0131  & ~\s15_msel_arb1_state_reg[1]/NET0131  ;
  assign n3830 = n3753 & n3829 ;
  assign n3831 = ~n3828 & ~n3830 ;
  assign n3832 = \s15_msel_arb1_state_reg[0]/NET0131  & \s15_msel_arb1_state_reg[1]/NET0131  ;
  assign n3833 = n3750 & ~n3832 ;
  assign n3834 = ~n3748 & ~n3833 ;
  assign n3835 = ~n3768 & n3834 ;
  assign n3836 = n3831 & n3835 ;
  assign n3837 = ~\s15_msel_arb1_state_reg[2]/NET0131  & ~n3836 ;
  assign n3838 = ~\rf_conf15_reg[9]/NET0131  & ~\s15_msel_arb1_state_reg[0]/NET0131  ;
  assign n3839 = n3765 & n3838 ;
  assign n3840 = ~n3764 & ~n3839 ;
  assign n3841 = ~\s15_msel_arb1_state_reg[1]/NET0131  & ~n3840 ;
  assign n3842 = \s15_msel_arb1_state_reg[2]/NET0131  & ~n3761 ;
  assign n3843 = n3759 & ~n3832 ;
  assign n3844 = n3842 & ~n3843 ;
  assign n3845 = ~n3757 & n3844 ;
  assign n3846 = ~n3841 & n3845 ;
  assign n3847 = ~n3837 & ~n3846 ;
  assign n3848 = \m5_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[10]/NET0131  ;
  assign n3849 = \rf_conf13_reg[11]/NET0131  & n3848 ;
  assign n3850 = \m4_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[8]/NET0131  ;
  assign n3851 = \rf_conf13_reg[9]/NET0131  & n3850 ;
  assign n3852 = ~n3849 & ~n3851 ;
  assign n3853 = ~\s13_msel_arb3_state_reg[0]/NET0131  & n3852 ;
  assign n3854 = \s13_msel_arb3_state_reg[0]/NET0131  & \s13_msel_arb3_state_reg[2]/NET0131  ;
  assign n3855 = ~\s13_msel_arb3_state_reg[1]/NET0131  & ~n3854 ;
  assign n3856 = \rf_conf13_reg[11]/NET0131  & ~\s13_msel_arb3_state_reg[1]/NET0131  ;
  assign n3857 = n3848 & n3856 ;
  assign n3858 = ~n3855 & ~n3857 ;
  assign n3859 = ~n3853 & ~n3858 ;
  assign n3860 = \m7_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[14]/NET0131  ;
  assign n3861 = \rf_conf13_reg[15]/NET0131  & n3860 ;
  assign n3862 = \m6_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[12]/NET0131  ;
  assign n3863 = \rf_conf13_reg[13]/NET0131  & n3862 ;
  assign n3864 = ~n3861 & ~n3863 ;
  assign n3865 = \m3_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[6]/NET0131  ;
  assign n3866 = \rf_conf13_reg[7]/NET0131  & n3865 ;
  assign n3867 = \m2_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[4]/NET0131  ;
  assign n3868 = \rf_conf13_reg[5]/NET0131  & n3867 ;
  assign n3869 = ~n3866 & ~n3868 ;
  assign n3870 = \m1_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[2]/NET0131  ;
  assign n3871 = \rf_conf13_reg[3]/NET0131  & n3870 ;
  assign n3872 = \m0_s13_cyc_o_reg/NET0131  & \rf_conf13_reg[0]/NET0131  ;
  assign n3873 = \rf_conf13_reg[1]/NET0131  & n3872 ;
  assign n3874 = ~n3871 & ~n3873 ;
  assign n3875 = n3869 & n3874 ;
  assign n3876 = n3864 & ~n3875 ;
  assign n3877 = ~n3859 & n3876 ;
  assign n3878 = ~\s13_msel_arb3_state_reg[0]/NET0131  & n3874 ;
  assign n3879 = ~\s13_msel_arb3_state_reg[1]/NET0131  & ~n3878 ;
  assign n3880 = n3852 & n3864 ;
  assign n3881 = \rf_conf13_reg[5]/NET0131  & ~\s13_msel_arb3_state_reg[0]/NET0131  ;
  assign n3882 = n3867 & n3881 ;
  assign n3883 = ~\s13_msel_arb3_state_reg[2]/NET0131  & ~n3882 ;
  assign n3884 = ~n3866 & n3883 ;
  assign n3885 = ~n3880 & n3884 ;
  assign n3886 = ~n3879 & n3885 ;
  assign n3887 = n3877 & ~n3886 ;
  assign n3888 = \s13_msel_arb3_state_reg[0]/NET0131  & \s13_msel_arb3_state_reg[1]/NET0131  ;
  assign n3889 = \s13_msel_arb3_state_reg[0]/NET0131  & ~n3868 ;
  assign n3890 = ~n3866 & ~n3871 ;
  assign n3891 = n3889 & n3890 ;
  assign n3892 = ~n3880 & n3891 ;
  assign n3893 = ~\s13_msel_arb3_state_reg[2]/NET0131  & ~n3892 ;
  assign n3894 = ~n3888 & ~n3893 ;
  assign n3895 = ~n3861 & ~n3875 ;
  assign n3896 = \s13_msel_arb3_state_reg[1]/NET0131  & \s13_msel_arb3_state_reg[2]/NET0131  ;
  assign n3897 = \s13_msel_arb3_state_reg[0]/NET0131  & n3896 ;
  assign n3898 = ~n3895 & n3897 ;
  assign n3899 = ~n3886 & ~n3898 ;
  assign n3900 = ~n3894 & n3899 ;
  assign n3901 = ~n3887 & ~n3900 ;
  assign n3902 = \rf_conf14_reg[11]/NET0131  & n2926 ;
  assign n3903 = \rf_conf14_reg[9]/NET0131  & n2928 ;
  assign n3904 = ~n3902 & ~n3903 ;
  assign n3905 = ~\s14_msel_arb2_state_reg[0]/NET0131  & n3904 ;
  assign n3906 = \s14_msel_arb2_state_reg[0]/NET0131  & \s14_msel_arb2_state_reg[2]/NET0131  ;
  assign n3907 = ~\s14_msel_arb2_state_reg[1]/NET0131  & ~n3906 ;
  assign n3908 = \rf_conf14_reg[11]/NET0131  & ~\s14_msel_arb2_state_reg[1]/NET0131  ;
  assign n3909 = n2926 & n3908 ;
  assign n3910 = ~n3907 & ~n3909 ;
  assign n3911 = ~n3905 & ~n3910 ;
  assign n3912 = \rf_conf14_reg[15]/NET0131  & n2931 ;
  assign n3913 = \rf_conf14_reg[13]/NET0131  & n2933 ;
  assign n3914 = ~n3912 & ~n3913 ;
  assign n3915 = \rf_conf14_reg[7]/NET0131  & n2943 ;
  assign n3916 = \rf_conf14_reg[5]/NET0131  & n2949 ;
  assign n3917 = ~n3915 & ~n3916 ;
  assign n3918 = \rf_conf14_reg[3]/NET0131  & n2936 ;
  assign n3919 = \rf_conf14_reg[1]/NET0131  & n2938 ;
  assign n3920 = ~n3918 & ~n3919 ;
  assign n3921 = n3917 & n3920 ;
  assign n3922 = n3914 & ~n3921 ;
  assign n3923 = ~n3911 & n3922 ;
  assign n3924 = ~\s14_msel_arb2_state_reg[0]/NET0131  & n3920 ;
  assign n3925 = ~\s14_msel_arb2_state_reg[1]/NET0131  & ~n3924 ;
  assign n3926 = n3904 & n3914 ;
  assign n3927 = \rf_conf14_reg[5]/NET0131  & ~\s14_msel_arb2_state_reg[0]/NET0131  ;
  assign n3928 = n2949 & n3927 ;
  assign n3929 = ~\s14_msel_arb2_state_reg[2]/NET0131  & ~n3928 ;
  assign n3930 = ~n3915 & n3929 ;
  assign n3931 = ~n3926 & n3930 ;
  assign n3932 = ~n3925 & n3931 ;
  assign n3933 = n3923 & ~n3932 ;
  assign n3934 = \s14_msel_arb2_state_reg[0]/NET0131  & \s14_msel_arb2_state_reg[1]/NET0131  ;
  assign n3935 = \s14_msel_arb2_state_reg[0]/NET0131  & ~n3916 ;
  assign n3936 = ~n3915 & ~n3918 ;
  assign n3937 = n3935 & n3936 ;
  assign n3938 = ~n3926 & n3937 ;
  assign n3939 = ~\s14_msel_arb2_state_reg[2]/NET0131  & ~n3938 ;
  assign n3940 = ~n3934 & ~n3939 ;
  assign n3941 = ~n3912 & ~n3921 ;
  assign n3942 = \s14_msel_arb2_state_reg[1]/NET0131  & \s14_msel_arb2_state_reg[2]/NET0131  ;
  assign n3943 = \s14_msel_arb2_state_reg[0]/NET0131  & n3942 ;
  assign n3944 = ~n3941 & n3943 ;
  assign n3945 = ~n3932 & ~n3944 ;
  assign n3946 = ~n3940 & n3945 ;
  assign n3947 = ~n3933 & ~n3946 ;
  assign n3948 = \m5_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[10]/NET0131  ;
  assign n3949 = \rf_conf2_reg[11]/NET0131  & n3948 ;
  assign n3950 = \m4_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[8]/NET0131  ;
  assign n3951 = \rf_conf2_reg[9]/NET0131  & n3950 ;
  assign n3952 = ~n3949 & ~n3951 ;
  assign n3953 = ~\s2_msel_arb3_state_reg[0]/NET0131  & n3952 ;
  assign n3954 = \s2_msel_arb3_state_reg[0]/NET0131  & \s2_msel_arb3_state_reg[2]/NET0131  ;
  assign n3955 = ~\s2_msel_arb3_state_reg[1]/NET0131  & ~n3954 ;
  assign n3956 = \rf_conf2_reg[11]/NET0131  & ~\s2_msel_arb3_state_reg[1]/NET0131  ;
  assign n3957 = n3948 & n3956 ;
  assign n3958 = ~n3955 & ~n3957 ;
  assign n3959 = ~n3953 & ~n3958 ;
  assign n3960 = \m7_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[14]/NET0131  ;
  assign n3961 = \rf_conf2_reg[15]/NET0131  & n3960 ;
  assign n3962 = \m6_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[12]/NET0131  ;
  assign n3963 = \rf_conf2_reg[13]/NET0131  & n3962 ;
  assign n3964 = ~n3961 & ~n3963 ;
  assign n3965 = \m3_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[6]/NET0131  ;
  assign n3966 = \rf_conf2_reg[7]/NET0131  & n3965 ;
  assign n3967 = \m2_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[4]/NET0131  ;
  assign n3968 = \rf_conf2_reg[5]/NET0131  & n3967 ;
  assign n3969 = ~n3966 & ~n3968 ;
  assign n3970 = \m1_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[2]/NET0131  ;
  assign n3971 = \rf_conf2_reg[3]/NET0131  & n3970 ;
  assign n3972 = \m0_s2_cyc_o_reg/NET0131  & \rf_conf2_reg[0]/NET0131  ;
  assign n3973 = \rf_conf2_reg[1]/NET0131  & n3972 ;
  assign n3974 = ~n3971 & ~n3973 ;
  assign n3975 = n3969 & n3974 ;
  assign n3976 = n3964 & ~n3975 ;
  assign n3977 = ~n3959 & n3976 ;
  assign n3978 = ~\s2_msel_arb3_state_reg[0]/NET0131  & n3974 ;
  assign n3979 = ~\s2_msel_arb3_state_reg[1]/NET0131  & ~n3978 ;
  assign n3980 = n3952 & n3964 ;
  assign n3981 = \rf_conf2_reg[5]/NET0131  & ~\s2_msel_arb3_state_reg[0]/NET0131  ;
  assign n3982 = n3967 & n3981 ;
  assign n3983 = ~\s2_msel_arb3_state_reg[2]/NET0131  & ~n3982 ;
  assign n3984 = ~n3966 & n3983 ;
  assign n3985 = ~n3980 & n3984 ;
  assign n3986 = ~n3979 & n3985 ;
  assign n3987 = n3977 & ~n3986 ;
  assign n3988 = \s2_msel_arb3_state_reg[0]/NET0131  & \s2_msel_arb3_state_reg[1]/NET0131  ;
  assign n3989 = \s2_msel_arb3_state_reg[0]/NET0131  & ~n3968 ;
  assign n3990 = ~n3966 & ~n3971 ;
  assign n3991 = n3989 & n3990 ;
  assign n3992 = ~n3980 & n3991 ;
  assign n3993 = ~\s2_msel_arb3_state_reg[2]/NET0131  & ~n3992 ;
  assign n3994 = ~n3988 & ~n3993 ;
  assign n3995 = ~n3961 & ~n3975 ;
  assign n3996 = \s2_msel_arb3_state_reg[1]/NET0131  & \s2_msel_arb3_state_reg[2]/NET0131  ;
  assign n3997 = \s2_msel_arb3_state_reg[0]/NET0131  & n3996 ;
  assign n3998 = ~n3995 & n3997 ;
  assign n3999 = ~n3986 & ~n3998 ;
  assign n4000 = ~n3994 & n3999 ;
  assign n4001 = ~n3987 & ~n4000 ;
  assign n4002 = \rf_conf3_reg[11]/NET0131  & n3059 ;
  assign n4003 = \rf_conf3_reg[9]/NET0131  & n3061 ;
  assign n4004 = ~n4002 & ~n4003 ;
  assign n4005 = \rf_conf3_reg[13]/NET0131  & n3066 ;
  assign n4006 = \rf_conf3_reg[15]/NET0131  & n3064 ;
  assign n4007 = ~n4005 & ~n4006 ;
  assign n4008 = n4004 & n4007 ;
  assign n4009 = \rf_conf3_reg[7]/NET0131  & n3076 ;
  assign n4010 = ~\s3_msel_arb2_state_reg[2]/NET0131  & ~n4009 ;
  assign n4011 = ~n4008 & n4010 ;
  assign n4012 = \rf_conf3_reg[5]/NET0131  & n3082 ;
  assign n4013 = \rf_conf3_reg[1]/NET0131  & ~\s3_msel_arb2_state_reg[1]/NET0131  ;
  assign n4014 = n3071 & n4013 ;
  assign n4015 = ~n4012 & ~n4014 ;
  assign n4016 = ~\s3_msel_arb2_state_reg[0]/NET0131  & ~n4015 ;
  assign n4017 = \rf_conf3_reg[3]/NET0131  & n3069 ;
  assign n4018 = ~n4012 & ~n4017 ;
  assign n4019 = ~\s3_msel_arb2_state_reg[1]/NET0131  & ~n4018 ;
  assign n4020 = ~n4016 & ~n4019 ;
  assign n4021 = n4011 & n4020 ;
  assign n4022 = ~n4009 & ~n4012 ;
  assign n4023 = \rf_conf3_reg[1]/NET0131  & n3071 ;
  assign n4024 = ~n4017 & ~n4023 ;
  assign n4025 = n4022 & n4024 ;
  assign n4026 = ~n4006 & ~n4025 ;
  assign n4027 = \rf_conf3_reg[9]/NET0131  & ~\s3_msel_arb2_state_reg[1]/NET0131  ;
  assign n4028 = n3061 & n4027 ;
  assign n4029 = ~n4005 & ~n4028 ;
  assign n4030 = ~\s3_msel_arb2_state_reg[0]/NET0131  & ~n4029 ;
  assign n4031 = ~n4002 & ~n4005 ;
  assign n4032 = ~\s3_msel_arb2_state_reg[1]/NET0131  & ~n4031 ;
  assign n4033 = ~n4030 & ~n4032 ;
  assign n4034 = n4026 & n4033 ;
  assign n4035 = \s3_msel_arb2_state_reg[2]/NET0131  & ~n4034 ;
  assign n4036 = ~n4021 & ~n4035 ;
  assign n4037 = ~\s4_msel_arb3_state_reg[1]/NET0131  & \s4_msel_arb3_state_reg[2]/NET0131  ;
  assign n4038 = \m1_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[2]/NET0131  ;
  assign n4039 = \rf_conf4_reg[3]/NET0131  & n4038 ;
  assign n4040 = \m0_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[0]/NET0131  ;
  assign n4041 = \rf_conf4_reg[1]/NET0131  & n4040 ;
  assign n4042 = ~n4039 & ~n4041 ;
  assign n4043 = \m3_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[6]/NET0131  ;
  assign n4044 = \rf_conf4_reg[7]/NET0131  & n4043 ;
  assign n4045 = \m2_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[4]/NET0131  ;
  assign n4046 = \rf_conf4_reg[5]/NET0131  & n4045 ;
  assign n4047 = ~n4044 & ~n4046 ;
  assign n4048 = n4042 & n4047 ;
  assign n4049 = \m5_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[10]/NET0131  ;
  assign n4050 = \rf_conf4_reg[11]/NET0131  & n4049 ;
  assign n4051 = \m7_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[14]/NET0131  ;
  assign n4052 = \rf_conf4_reg[15]/NET0131  & n4051 ;
  assign n4053 = \m6_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[12]/NET0131  ;
  assign n4054 = \rf_conf4_reg[13]/NET0131  & n4053 ;
  assign n4055 = ~n4052 & ~n4054 ;
  assign n4056 = ~n4050 & n4055 ;
  assign n4057 = ~n4048 & n4056 ;
  assign n4058 = n4037 & ~n4057 ;
  assign n4059 = ~n4048 & ~n4052 ;
  assign n4060 = \s4_msel_arb3_state_reg[1]/NET0131  & \s4_msel_arb3_state_reg[2]/NET0131  ;
  assign n4061 = ~n4059 & n4060 ;
  assign n4062 = \m4_s4_cyc_o_reg/NET0131  & \rf_conf4_reg[8]/NET0131  ;
  assign n4063 = \rf_conf4_reg[9]/NET0131  & n4062 ;
  assign n4064 = ~n4050 & ~n4063 ;
  assign n4065 = n4055 & n4064 ;
  assign n4066 = ~n4044 & ~n4065 ;
  assign n4067 = ~\s4_msel_arb3_state_reg[2]/NET0131  & ~n4039 ;
  assign n4068 = ~\s4_msel_arb3_state_reg[1]/NET0131  & ~n4046 ;
  assign n4069 = n4067 & n4068 ;
  assign n4070 = n4066 & n4069 ;
  assign n4071 = ~n4061 & ~n4070 ;
  assign n4072 = ~n4058 & n4071 ;
  assign n4073 = \s4_msel_arb3_state_reg[0]/NET0131  & ~n4072 ;
  assign n4074 = \rf_conf4_reg[5]/NET0131  & ~\s4_msel_arb3_state_reg[0]/NET0131  ;
  assign n4075 = n4045 & n4074 ;
  assign n4076 = ~\s4_msel_arb3_state_reg[1]/NET0131  & ~n4042 ;
  assign n4077 = ~n4075 & ~n4076 ;
  assign n4078 = n4066 & n4077 ;
  assign n4079 = ~\s4_msel_arb3_state_reg[2]/NET0131  & ~n4078 ;
  assign n4080 = \s4_msel_arb3_state_reg[1]/NET0131  & ~\s4_msel_arb3_state_reg[2]/NET0131  ;
  assign n4081 = \s4_msel_arb3_state_reg[0]/NET0131  & ~n4080 ;
  assign n4082 = ~n4048 & n4055 ;
  assign n4083 = ~n4060 & ~n4064 ;
  assign n4084 = n4082 & ~n4083 ;
  assign n4085 = ~n4081 & ~n4084 ;
  assign n4086 = ~n4079 & n4085 ;
  assign n4087 = ~n4073 & ~n4086 ;
  assign n4088 = \rf_conf6_reg[11]/NET0131  & n3245 ;
  assign n4089 = \rf_conf6_reg[9]/NET0131  & n3247 ;
  assign n4090 = ~n4088 & ~n4089 ;
  assign n4091 = \rf_conf6_reg[13]/NET0131  & n3252 ;
  assign n4092 = \rf_conf6_reg[15]/NET0131  & n3250 ;
  assign n4093 = ~n4091 & ~n4092 ;
  assign n4094 = n4090 & n4093 ;
  assign n4095 = \rf_conf6_reg[7]/NET0131  & n3262 ;
  assign n4096 = ~\s6_msel_arb2_state_reg[2]/NET0131  & ~n4095 ;
  assign n4097 = ~n4094 & n4096 ;
  assign n4098 = \rf_conf6_reg[5]/NET0131  & n3268 ;
  assign n4099 = \rf_conf6_reg[1]/NET0131  & ~\s6_msel_arb2_state_reg[1]/NET0131  ;
  assign n4100 = n3257 & n4099 ;
  assign n4101 = ~n4098 & ~n4100 ;
  assign n4102 = ~\s6_msel_arb2_state_reg[0]/NET0131  & ~n4101 ;
  assign n4103 = \rf_conf6_reg[3]/NET0131  & n3255 ;
  assign n4104 = ~n4098 & ~n4103 ;
  assign n4105 = ~\s6_msel_arb2_state_reg[1]/NET0131  & ~n4104 ;
  assign n4106 = ~n4102 & ~n4105 ;
  assign n4107 = n4097 & n4106 ;
  assign n4108 = ~n4095 & ~n4098 ;
  assign n4109 = \rf_conf6_reg[1]/NET0131  & n3257 ;
  assign n4110 = ~n4103 & ~n4109 ;
  assign n4111 = n4108 & n4110 ;
  assign n4112 = ~n4092 & ~n4111 ;
  assign n4113 = \rf_conf6_reg[9]/NET0131  & ~\s6_msel_arb2_state_reg[1]/NET0131  ;
  assign n4114 = n3247 & n4113 ;
  assign n4115 = ~n4091 & ~n4114 ;
  assign n4116 = ~\s6_msel_arb2_state_reg[0]/NET0131  & ~n4115 ;
  assign n4117 = ~n4088 & ~n4091 ;
  assign n4118 = ~\s6_msel_arb2_state_reg[1]/NET0131  & ~n4117 ;
  assign n4119 = ~n4116 & ~n4118 ;
  assign n4120 = n4112 & n4119 ;
  assign n4121 = \s6_msel_arb2_state_reg[2]/NET0131  & ~n4120 ;
  assign n4122 = ~n4107 & ~n4121 ;
  assign n4123 = \rf_conf8_reg[11]/NET0131  & n3307 ;
  assign n4124 = \rf_conf8_reg[9]/NET0131  & n3309 ;
  assign n4125 = ~n4123 & ~n4124 ;
  assign n4126 = \rf_conf8_reg[13]/NET0131  & n3314 ;
  assign n4127 = \rf_conf8_reg[15]/NET0131  & n3312 ;
  assign n4128 = ~n4126 & ~n4127 ;
  assign n4129 = n4125 & n4128 ;
  assign n4130 = \rf_conf8_reg[7]/NET0131  & n3324 ;
  assign n4131 = ~\s8_msel_arb2_state_reg[2]/NET0131  & ~n4130 ;
  assign n4132 = ~n4129 & n4131 ;
  assign n4133 = \rf_conf8_reg[5]/NET0131  & n3330 ;
  assign n4134 = \rf_conf8_reg[1]/NET0131  & ~\s8_msel_arb2_state_reg[1]/NET0131  ;
  assign n4135 = n3319 & n4134 ;
  assign n4136 = ~n4133 & ~n4135 ;
  assign n4137 = ~\s8_msel_arb2_state_reg[0]/NET0131  & ~n4136 ;
  assign n4138 = \rf_conf8_reg[3]/NET0131  & n3317 ;
  assign n4139 = ~n4133 & ~n4138 ;
  assign n4140 = ~\s8_msel_arb2_state_reg[1]/NET0131  & ~n4139 ;
  assign n4141 = ~n4137 & ~n4140 ;
  assign n4142 = n4132 & n4141 ;
  assign n4143 = ~n4130 & ~n4133 ;
  assign n4144 = \rf_conf8_reg[1]/NET0131  & n3319 ;
  assign n4145 = ~n4138 & ~n4144 ;
  assign n4146 = n4143 & n4145 ;
  assign n4147 = ~n4127 & ~n4146 ;
  assign n4148 = \rf_conf8_reg[9]/NET0131  & ~\s8_msel_arb2_state_reg[1]/NET0131  ;
  assign n4149 = n3309 & n4148 ;
  assign n4150 = ~n4126 & ~n4149 ;
  assign n4151 = ~\s8_msel_arb2_state_reg[0]/NET0131  & ~n4150 ;
  assign n4152 = ~n4123 & ~n4126 ;
  assign n4153 = ~\s8_msel_arb2_state_reg[1]/NET0131  & ~n4152 ;
  assign n4154 = ~n4151 & ~n4153 ;
  assign n4155 = n4147 & n4154 ;
  assign n4156 = \s8_msel_arb2_state_reg[2]/NET0131  & ~n4155 ;
  assign n4157 = ~n4142 & ~n4156 ;
  assign n4158 = \rf_conf0_reg[11]/NET0131  & n3628 ;
  assign n4159 = \rf_conf0_reg[9]/NET0131  & n3626 ;
  assign n4160 = ~n4158 & ~n4159 ;
  assign n4161 = \rf_conf0_reg[13]/NET0131  & n3633 ;
  assign n4162 = \rf_conf0_reg[15]/NET0131  & n3631 ;
  assign n4163 = ~n4161 & ~n4162 ;
  assign n4164 = n4160 & n4163 ;
  assign n4165 = \rf_conf0_reg[7]/NET0131  & n3621 ;
  assign n4166 = ~\s0_msel_arb2_state_reg[2]/NET0131  & ~n4165 ;
  assign n4167 = ~n4164 & n4166 ;
  assign n4168 = \rf_conf0_reg[5]/NET0131  & n3623 ;
  assign n4169 = \rf_conf0_reg[1]/NET0131  & ~\s0_msel_arb2_state_reg[1]/NET0131  ;
  assign n4170 = n3640 & n4169 ;
  assign n4171 = ~n4168 & ~n4170 ;
  assign n4172 = ~\s0_msel_arb2_state_reg[0]/NET0131  & ~n4171 ;
  assign n4173 = \rf_conf0_reg[3]/NET0131  & n3638 ;
  assign n4174 = ~n4168 & ~n4173 ;
  assign n4175 = ~\s0_msel_arb2_state_reg[1]/NET0131  & ~n4174 ;
  assign n4176 = ~n4172 & ~n4175 ;
  assign n4177 = n4167 & n4176 ;
  assign n4178 = ~n4165 & ~n4168 ;
  assign n4179 = \rf_conf0_reg[1]/NET0131  & n3640 ;
  assign n4180 = ~n4173 & ~n4179 ;
  assign n4181 = n4178 & n4180 ;
  assign n4182 = ~n4162 & ~n4181 ;
  assign n4183 = \rf_conf0_reg[9]/NET0131  & ~\s0_msel_arb2_state_reg[1]/NET0131  ;
  assign n4184 = n3626 & n4183 ;
  assign n4185 = ~n4161 & ~n4184 ;
  assign n4186 = ~\s0_msel_arb2_state_reg[0]/NET0131  & ~n4185 ;
  assign n4187 = ~n4158 & ~n4161 ;
  assign n4188 = ~\s0_msel_arb2_state_reg[1]/NET0131  & ~n4187 ;
  assign n4189 = ~n4186 & ~n4188 ;
  assign n4190 = n4182 & n4189 ;
  assign n4191 = \s0_msel_arb2_state_reg[2]/NET0131  & ~n4190 ;
  assign n4192 = ~n4177 & ~n4191 ;
  assign n4193 = \m5_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[10]/NET0131  ;
  assign n4194 = \rf_conf10_reg[11]/NET0131  & n4193 ;
  assign n4195 = \m4_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[8]/NET0131  ;
  assign n4196 = \rf_conf10_reg[9]/NET0131  & n4195 ;
  assign n4197 = ~n4194 & ~n4196 ;
  assign n4198 = ~\s10_msel_arb3_state_reg[0]/NET0131  & n4197 ;
  assign n4199 = \s10_msel_arb3_state_reg[0]/NET0131  & \s10_msel_arb3_state_reg[2]/NET0131  ;
  assign n4200 = ~\s10_msel_arb3_state_reg[1]/NET0131  & ~n4199 ;
  assign n4201 = \rf_conf10_reg[11]/NET0131  & ~\s10_msel_arb3_state_reg[1]/NET0131  ;
  assign n4202 = n4193 & n4201 ;
  assign n4203 = ~n4200 & ~n4202 ;
  assign n4204 = ~n4198 & ~n4203 ;
  assign n4205 = \m7_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[14]/NET0131  ;
  assign n4206 = \rf_conf10_reg[15]/NET0131  & n4205 ;
  assign n4207 = \m6_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[12]/NET0131  ;
  assign n4208 = \rf_conf10_reg[13]/NET0131  & n4207 ;
  assign n4209 = ~n4206 & ~n4208 ;
  assign n4210 = \m3_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[6]/NET0131  ;
  assign n4211 = \rf_conf10_reg[7]/NET0131  & n4210 ;
  assign n4212 = \m2_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[4]/NET0131  ;
  assign n4213 = \rf_conf10_reg[5]/NET0131  & n4212 ;
  assign n4214 = ~n4211 & ~n4213 ;
  assign n4215 = \m1_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[2]/NET0131  ;
  assign n4216 = \rf_conf10_reg[3]/NET0131  & n4215 ;
  assign n4217 = \m0_s10_cyc_o_reg/NET0131  & \rf_conf10_reg[0]/NET0131  ;
  assign n4218 = \rf_conf10_reg[1]/NET0131  & n4217 ;
  assign n4219 = ~n4216 & ~n4218 ;
  assign n4220 = n4214 & n4219 ;
  assign n4221 = n4209 & ~n4220 ;
  assign n4222 = ~n4204 & n4221 ;
  assign n4223 = ~\s10_msel_arb3_state_reg[0]/NET0131  & n4219 ;
  assign n4224 = ~\s10_msel_arb3_state_reg[1]/NET0131  & ~n4223 ;
  assign n4225 = n4197 & n4209 ;
  assign n4226 = \rf_conf10_reg[5]/NET0131  & ~\s10_msel_arb3_state_reg[0]/NET0131  ;
  assign n4227 = n4212 & n4226 ;
  assign n4228 = ~\s10_msel_arb3_state_reg[2]/NET0131  & ~n4227 ;
  assign n4229 = ~n4211 & n4228 ;
  assign n4230 = ~n4225 & n4229 ;
  assign n4231 = ~n4224 & n4230 ;
  assign n4232 = n4222 & ~n4231 ;
  assign n4233 = \s10_msel_arb3_state_reg[0]/NET0131  & \s10_msel_arb3_state_reg[1]/NET0131  ;
  assign n4234 = \s10_msel_arb3_state_reg[0]/NET0131  & ~n4213 ;
  assign n4235 = ~n4211 & ~n4216 ;
  assign n4236 = n4234 & n4235 ;
  assign n4237 = ~n4225 & n4236 ;
  assign n4238 = ~\s10_msel_arb3_state_reg[2]/NET0131  & ~n4237 ;
  assign n4239 = ~n4233 & ~n4238 ;
  assign n4240 = ~n4206 & ~n4220 ;
  assign n4241 = \s10_msel_arb3_state_reg[1]/NET0131  & \s10_msel_arb3_state_reg[2]/NET0131  ;
  assign n4242 = \s10_msel_arb3_state_reg[0]/NET0131  & n4241 ;
  assign n4243 = ~n4240 & n4242 ;
  assign n4244 = ~n4231 & ~n4243 ;
  assign n4245 = ~n4239 & n4244 ;
  assign n4246 = ~n4232 & ~n4245 ;
  assign n4247 = \rf_conf11_reg[11]/NET0131  & n2740 ;
  assign n4248 = \rf_conf11_reg[9]/NET0131  & n2742 ;
  assign n4249 = ~n4247 & ~n4248 ;
  assign n4250 = \rf_conf11_reg[13]/NET0131  & n2747 ;
  assign n4251 = \rf_conf11_reg[15]/NET0131  & n2745 ;
  assign n4252 = ~n4250 & ~n4251 ;
  assign n4253 = n4249 & n4252 ;
  assign n4254 = \rf_conf11_reg[7]/NET0131  & n2757 ;
  assign n4255 = ~\s11_msel_arb2_state_reg[2]/NET0131  & ~n4254 ;
  assign n4256 = ~n4253 & n4255 ;
  assign n4257 = \rf_conf11_reg[5]/NET0131  & n2763 ;
  assign n4258 = \rf_conf11_reg[1]/NET0131  & ~\s11_msel_arb2_state_reg[1]/NET0131  ;
  assign n4259 = n2752 & n4258 ;
  assign n4260 = ~n4257 & ~n4259 ;
  assign n4261 = ~\s11_msel_arb2_state_reg[0]/NET0131  & ~n4260 ;
  assign n4262 = \rf_conf11_reg[3]/NET0131  & n2750 ;
  assign n4263 = ~n4257 & ~n4262 ;
  assign n4264 = ~\s11_msel_arb2_state_reg[1]/NET0131  & ~n4263 ;
  assign n4265 = ~n4261 & ~n4264 ;
  assign n4266 = n4256 & n4265 ;
  assign n4267 = ~n4254 & ~n4257 ;
  assign n4268 = \rf_conf11_reg[1]/NET0131  & n2752 ;
  assign n4269 = ~n4262 & ~n4268 ;
  assign n4270 = n4267 & n4269 ;
  assign n4271 = ~n4251 & ~n4270 ;
  assign n4272 = \rf_conf11_reg[9]/NET0131  & ~\s11_msel_arb2_state_reg[1]/NET0131  ;
  assign n4273 = n2742 & n4272 ;
  assign n4274 = ~n4250 & ~n4273 ;
  assign n4275 = ~\s11_msel_arb2_state_reg[0]/NET0131  & ~n4274 ;
  assign n4276 = ~n4247 & ~n4250 ;
  assign n4277 = ~\s11_msel_arb2_state_reg[1]/NET0131  & ~n4276 ;
  assign n4278 = ~n4275 & ~n4277 ;
  assign n4279 = n4271 & n4278 ;
  assign n4280 = \s11_msel_arb2_state_reg[2]/NET0131  & ~n4279 ;
  assign n4281 = ~n4266 & ~n4280 ;
  assign n4282 = ~\s11_msel_arb3_state_reg[1]/NET0131  & \s11_msel_arb3_state_reg[2]/NET0131  ;
  assign n4283 = \m1_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[2]/NET0131  ;
  assign n4284 = \rf_conf11_reg[3]/NET0131  & n4283 ;
  assign n4285 = \m0_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[0]/NET0131  ;
  assign n4286 = \rf_conf11_reg[1]/NET0131  & n4285 ;
  assign n4287 = ~n4284 & ~n4286 ;
  assign n4288 = \m3_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[6]/NET0131  ;
  assign n4289 = \rf_conf11_reg[7]/NET0131  & n4288 ;
  assign n4290 = \m2_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[4]/NET0131  ;
  assign n4291 = \rf_conf11_reg[5]/NET0131  & n4290 ;
  assign n4292 = ~n4289 & ~n4291 ;
  assign n4293 = n4287 & n4292 ;
  assign n4294 = \m5_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[10]/NET0131  ;
  assign n4295 = \rf_conf11_reg[11]/NET0131  & n4294 ;
  assign n4296 = \m7_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[14]/NET0131  ;
  assign n4297 = \rf_conf11_reg[15]/NET0131  & n4296 ;
  assign n4298 = \m6_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[12]/NET0131  ;
  assign n4299 = \rf_conf11_reg[13]/NET0131  & n4298 ;
  assign n4300 = ~n4297 & ~n4299 ;
  assign n4301 = ~n4295 & n4300 ;
  assign n4302 = ~n4293 & n4301 ;
  assign n4303 = n4282 & ~n4302 ;
  assign n4304 = ~n4293 & ~n4297 ;
  assign n4305 = \s11_msel_arb3_state_reg[1]/NET0131  & \s11_msel_arb3_state_reg[2]/NET0131  ;
  assign n4306 = ~n4304 & n4305 ;
  assign n4307 = \m4_s11_cyc_o_reg/NET0131  & \rf_conf11_reg[8]/NET0131  ;
  assign n4308 = \rf_conf11_reg[9]/NET0131  & n4307 ;
  assign n4309 = ~n4295 & ~n4308 ;
  assign n4310 = n4300 & n4309 ;
  assign n4311 = ~n4289 & ~n4310 ;
  assign n4312 = ~\s11_msel_arb3_state_reg[2]/NET0131  & ~n4284 ;
  assign n4313 = ~\s11_msel_arb3_state_reg[1]/NET0131  & ~n4291 ;
  assign n4314 = n4312 & n4313 ;
  assign n4315 = n4311 & n4314 ;
  assign n4316 = ~n4306 & ~n4315 ;
  assign n4317 = ~n4303 & n4316 ;
  assign n4318 = \s11_msel_arb3_state_reg[0]/NET0131  & ~n4317 ;
  assign n4319 = \rf_conf11_reg[5]/NET0131  & ~\s11_msel_arb3_state_reg[0]/NET0131  ;
  assign n4320 = n4290 & n4319 ;
  assign n4321 = ~\s11_msel_arb3_state_reg[1]/NET0131  & ~n4287 ;
  assign n4322 = ~n4320 & ~n4321 ;
  assign n4323 = n4311 & n4322 ;
  assign n4324 = ~\s11_msel_arb3_state_reg[2]/NET0131  & ~n4323 ;
  assign n4325 = \s11_msel_arb3_state_reg[1]/NET0131  & ~\s11_msel_arb3_state_reg[2]/NET0131  ;
  assign n4326 = \s11_msel_arb3_state_reg[0]/NET0131  & ~n4325 ;
  assign n4327 = ~n4293 & n4300 ;
  assign n4328 = ~n4305 & ~n4309 ;
  assign n4329 = n4327 & ~n4328 ;
  assign n4330 = ~n4326 & ~n4329 ;
  assign n4331 = ~n4324 & n4330 ;
  assign n4332 = ~n4318 & ~n4331 ;
  assign n4333 = \m5_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[10]/NET0131  ;
  assign n4334 = \rf_conf12_reg[11]/NET0131  & n4333 ;
  assign n4335 = \m4_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[8]/NET0131  ;
  assign n4336 = \rf_conf12_reg[9]/NET0131  & n4335 ;
  assign n4337 = ~n4334 & ~n4336 ;
  assign n4338 = ~\s12_msel_arb3_state_reg[0]/NET0131  & n4337 ;
  assign n4339 = \s12_msel_arb3_state_reg[0]/NET0131  & \s12_msel_arb3_state_reg[2]/NET0131  ;
  assign n4340 = ~\s12_msel_arb3_state_reg[1]/NET0131  & ~n4339 ;
  assign n4341 = \rf_conf12_reg[11]/NET0131  & ~\s12_msel_arb3_state_reg[1]/NET0131  ;
  assign n4342 = n4333 & n4341 ;
  assign n4343 = ~n4340 & ~n4342 ;
  assign n4344 = ~n4338 & ~n4343 ;
  assign n4345 = \m7_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[14]/NET0131  ;
  assign n4346 = \rf_conf12_reg[15]/NET0131  & n4345 ;
  assign n4347 = \m6_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[12]/NET0131  ;
  assign n4348 = \rf_conf12_reg[13]/NET0131  & n4347 ;
  assign n4349 = ~n4346 & ~n4348 ;
  assign n4350 = \m3_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[6]/NET0131  ;
  assign n4351 = \rf_conf12_reg[7]/NET0131  & n4350 ;
  assign n4352 = \m2_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[4]/NET0131  ;
  assign n4353 = \rf_conf12_reg[5]/NET0131  & n4352 ;
  assign n4354 = ~n4351 & ~n4353 ;
  assign n4355 = \m1_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[2]/NET0131  ;
  assign n4356 = \rf_conf12_reg[3]/NET0131  & n4355 ;
  assign n4357 = \m0_s12_cyc_o_reg/NET0131  & \rf_conf12_reg[0]/NET0131  ;
  assign n4358 = \rf_conf12_reg[1]/NET0131  & n4357 ;
  assign n4359 = ~n4356 & ~n4358 ;
  assign n4360 = n4354 & n4359 ;
  assign n4361 = n4349 & ~n4360 ;
  assign n4362 = ~n4344 & n4361 ;
  assign n4363 = ~\s12_msel_arb3_state_reg[0]/NET0131  & n4359 ;
  assign n4364 = ~\s12_msel_arb3_state_reg[1]/NET0131  & ~n4363 ;
  assign n4365 = n4337 & n4349 ;
  assign n4366 = \rf_conf12_reg[5]/NET0131  & ~\s12_msel_arb3_state_reg[0]/NET0131  ;
  assign n4367 = n4352 & n4366 ;
  assign n4368 = ~\s12_msel_arb3_state_reg[2]/NET0131  & ~n4367 ;
  assign n4369 = ~n4351 & n4368 ;
  assign n4370 = ~n4365 & n4369 ;
  assign n4371 = ~n4364 & n4370 ;
  assign n4372 = n4362 & ~n4371 ;
  assign n4373 = \s12_msel_arb3_state_reg[0]/NET0131  & \s12_msel_arb3_state_reg[1]/NET0131  ;
  assign n4374 = \s12_msel_arb3_state_reg[0]/NET0131  & ~n4353 ;
  assign n4375 = ~n4351 & ~n4356 ;
  assign n4376 = n4374 & n4375 ;
  assign n4377 = ~n4365 & n4376 ;
  assign n4378 = ~\s12_msel_arb3_state_reg[2]/NET0131  & ~n4377 ;
  assign n4379 = ~n4373 & ~n4378 ;
  assign n4380 = ~n4346 & ~n4360 ;
  assign n4381 = \s12_msel_arb3_state_reg[1]/NET0131  & \s12_msel_arb3_state_reg[2]/NET0131  ;
  assign n4382 = \s12_msel_arb3_state_reg[0]/NET0131  & n4381 ;
  assign n4383 = ~n4380 & n4382 ;
  assign n4384 = ~n4371 & ~n4383 ;
  assign n4385 = ~n4379 & n4384 ;
  assign n4386 = ~n4372 & ~n4385 ;
  assign n4387 = ~\s14_msel_arb3_state_reg[1]/NET0131  & \s14_msel_arb3_state_reg[2]/NET0131  ;
  assign n4388 = \m1_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[2]/NET0131  ;
  assign n4389 = \rf_conf14_reg[3]/NET0131  & n4388 ;
  assign n4390 = \m0_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[0]/NET0131  ;
  assign n4391 = \rf_conf14_reg[1]/NET0131  & n4390 ;
  assign n4392 = ~n4389 & ~n4391 ;
  assign n4393 = \m3_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[6]/NET0131  ;
  assign n4394 = \rf_conf14_reg[7]/NET0131  & n4393 ;
  assign n4395 = \m2_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[4]/NET0131  ;
  assign n4396 = \rf_conf14_reg[5]/NET0131  & n4395 ;
  assign n4397 = ~n4394 & ~n4396 ;
  assign n4398 = n4392 & n4397 ;
  assign n4399 = \m5_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[10]/NET0131  ;
  assign n4400 = \rf_conf14_reg[11]/NET0131  & n4399 ;
  assign n4401 = \m7_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[14]/NET0131  ;
  assign n4402 = \rf_conf14_reg[15]/NET0131  & n4401 ;
  assign n4403 = \m6_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[12]/NET0131  ;
  assign n4404 = \rf_conf14_reg[13]/NET0131  & n4403 ;
  assign n4405 = ~n4402 & ~n4404 ;
  assign n4406 = ~n4400 & n4405 ;
  assign n4407 = ~n4398 & n4406 ;
  assign n4408 = n4387 & ~n4407 ;
  assign n4409 = ~n4398 & ~n4402 ;
  assign n4410 = \s14_msel_arb3_state_reg[1]/NET0131  & \s14_msel_arb3_state_reg[2]/NET0131  ;
  assign n4411 = ~n4409 & n4410 ;
  assign n4412 = \m4_s14_cyc_o_reg/NET0131  & \rf_conf14_reg[8]/NET0131  ;
  assign n4413 = \rf_conf14_reg[9]/NET0131  & n4412 ;
  assign n4414 = ~n4400 & ~n4413 ;
  assign n4415 = n4405 & n4414 ;
  assign n4416 = ~n4394 & ~n4415 ;
  assign n4417 = ~\s14_msel_arb3_state_reg[2]/NET0131  & ~n4389 ;
  assign n4418 = ~\s14_msel_arb3_state_reg[1]/NET0131  & ~n4396 ;
  assign n4419 = n4417 & n4418 ;
  assign n4420 = n4416 & n4419 ;
  assign n4421 = ~n4411 & ~n4420 ;
  assign n4422 = ~n4408 & n4421 ;
  assign n4423 = \s14_msel_arb3_state_reg[0]/NET0131  & ~n4422 ;
  assign n4424 = \rf_conf14_reg[5]/NET0131  & ~\s14_msel_arb3_state_reg[0]/NET0131  ;
  assign n4425 = n4395 & n4424 ;
  assign n4426 = ~\s14_msel_arb3_state_reg[1]/NET0131  & ~n4392 ;
  assign n4427 = ~n4425 & ~n4426 ;
  assign n4428 = n4416 & n4427 ;
  assign n4429 = ~\s14_msel_arb3_state_reg[2]/NET0131  & ~n4428 ;
  assign n4430 = \s14_msel_arb3_state_reg[1]/NET0131  & ~\s14_msel_arb3_state_reg[2]/NET0131  ;
  assign n4431 = \s14_msel_arb3_state_reg[0]/NET0131  & ~n4430 ;
  assign n4432 = ~n4398 & n4405 ;
  assign n4433 = ~n4410 & ~n4414 ;
  assign n4434 = n4432 & ~n4433 ;
  assign n4435 = ~n4431 & ~n4434 ;
  assign n4436 = ~n4429 & n4435 ;
  assign n4437 = ~n4423 & ~n4436 ;
  assign n4438 = \rf_conf1_reg[11]/NET0131  & n3376 ;
  assign n4439 = \rf_conf1_reg[9]/NET0131  & n3374 ;
  assign n4440 = ~n4438 & ~n4439 ;
  assign n4441 = \rf_conf1_reg[13]/NET0131  & n3381 ;
  assign n4442 = \rf_conf1_reg[15]/NET0131  & n3379 ;
  assign n4443 = ~n4441 & ~n4442 ;
  assign n4444 = n4440 & n4443 ;
  assign n4445 = \rf_conf1_reg[7]/NET0131  & n3369 ;
  assign n4446 = ~\s1_msel_arb2_state_reg[2]/NET0131  & ~n4445 ;
  assign n4447 = ~n4444 & n4446 ;
  assign n4448 = \rf_conf1_reg[5]/NET0131  & n3371 ;
  assign n4449 = \rf_conf1_reg[1]/NET0131  & ~\s1_msel_arb2_state_reg[1]/NET0131  ;
  assign n4450 = n3388 & n4449 ;
  assign n4451 = ~n4448 & ~n4450 ;
  assign n4452 = ~\s1_msel_arb2_state_reg[0]/NET0131  & ~n4451 ;
  assign n4453 = \rf_conf1_reg[3]/NET0131  & n3386 ;
  assign n4454 = ~n4448 & ~n4453 ;
  assign n4455 = ~\s1_msel_arb2_state_reg[1]/NET0131  & ~n4454 ;
  assign n4456 = ~n4452 & ~n4455 ;
  assign n4457 = n4447 & n4456 ;
  assign n4458 = ~n4445 & ~n4448 ;
  assign n4459 = \rf_conf1_reg[1]/NET0131  & n3388 ;
  assign n4460 = ~n4453 & ~n4459 ;
  assign n4461 = n4458 & n4460 ;
  assign n4462 = ~n4442 & ~n4461 ;
  assign n4463 = \rf_conf1_reg[9]/NET0131  & ~\s1_msel_arb2_state_reg[1]/NET0131  ;
  assign n4464 = n3374 & n4463 ;
  assign n4465 = ~n4441 & ~n4464 ;
  assign n4466 = ~\s1_msel_arb2_state_reg[0]/NET0131  & ~n4465 ;
  assign n4467 = ~n4438 & ~n4441 ;
  assign n4468 = ~\s1_msel_arb2_state_reg[1]/NET0131  & ~n4467 ;
  assign n4469 = ~n4466 & ~n4468 ;
  assign n4470 = n4462 & n4469 ;
  assign n4471 = \s1_msel_arb2_state_reg[2]/NET0131  & ~n4470 ;
  assign n4472 = ~n4457 & ~n4471 ;
  assign n4473 = ~\s1_msel_arb3_state_reg[1]/NET0131  & \s1_msel_arb3_state_reg[2]/NET0131  ;
  assign n4474 = \m1_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[2]/NET0131  ;
  assign n4475 = \rf_conf1_reg[3]/NET0131  & n4474 ;
  assign n4476 = \m0_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[0]/NET0131  ;
  assign n4477 = \rf_conf1_reg[1]/NET0131  & n4476 ;
  assign n4478 = ~n4475 & ~n4477 ;
  assign n4479 = \m3_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[6]/NET0131  ;
  assign n4480 = \rf_conf1_reg[7]/NET0131  & n4479 ;
  assign n4481 = \m2_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[4]/NET0131  ;
  assign n4482 = \rf_conf1_reg[5]/NET0131  & n4481 ;
  assign n4483 = ~n4480 & ~n4482 ;
  assign n4484 = n4478 & n4483 ;
  assign n4485 = \m5_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[10]/NET0131  ;
  assign n4486 = \rf_conf1_reg[11]/NET0131  & n4485 ;
  assign n4487 = \m7_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[14]/NET0131  ;
  assign n4488 = \rf_conf1_reg[15]/NET0131  & n4487 ;
  assign n4489 = \m6_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[12]/NET0131  ;
  assign n4490 = \rf_conf1_reg[13]/NET0131  & n4489 ;
  assign n4491 = ~n4488 & ~n4490 ;
  assign n4492 = ~n4486 & n4491 ;
  assign n4493 = ~n4484 & n4492 ;
  assign n4494 = n4473 & ~n4493 ;
  assign n4495 = ~n4484 & ~n4488 ;
  assign n4496 = \s1_msel_arb3_state_reg[1]/NET0131  & \s1_msel_arb3_state_reg[2]/NET0131  ;
  assign n4497 = ~n4495 & n4496 ;
  assign n4498 = \m4_s1_cyc_o_reg/NET0131  & \rf_conf1_reg[8]/NET0131  ;
  assign n4499 = \rf_conf1_reg[9]/NET0131  & n4498 ;
  assign n4500 = ~n4486 & ~n4499 ;
  assign n4501 = n4491 & n4500 ;
  assign n4502 = ~n4480 & ~n4501 ;
  assign n4503 = ~\s1_msel_arb3_state_reg[2]/NET0131  & ~n4475 ;
  assign n4504 = ~\s1_msel_arb3_state_reg[1]/NET0131  & ~n4482 ;
  assign n4505 = n4503 & n4504 ;
  assign n4506 = n4502 & n4505 ;
  assign n4507 = ~n4497 & ~n4506 ;
  assign n4508 = ~n4494 & n4507 ;
  assign n4509 = \s1_msel_arb3_state_reg[0]/NET0131  & ~n4508 ;
  assign n4510 = \rf_conf1_reg[5]/NET0131  & ~\s1_msel_arb3_state_reg[0]/NET0131  ;
  assign n4511 = n4481 & n4510 ;
  assign n4512 = ~\s1_msel_arb3_state_reg[1]/NET0131  & ~n4478 ;
  assign n4513 = ~n4511 & ~n4512 ;
  assign n4514 = n4502 & n4513 ;
  assign n4515 = ~\s1_msel_arb3_state_reg[2]/NET0131  & ~n4514 ;
  assign n4516 = \s1_msel_arb3_state_reg[1]/NET0131  & ~\s1_msel_arb3_state_reg[2]/NET0131  ;
  assign n4517 = \s1_msel_arb3_state_reg[0]/NET0131  & ~n4516 ;
  assign n4518 = ~n4484 & n4491 ;
  assign n4519 = ~n4496 & ~n4500 ;
  assign n4520 = n4518 & ~n4519 ;
  assign n4521 = ~n4517 & ~n4520 ;
  assign n4522 = ~n4515 & n4521 ;
  assign n4523 = ~n4509 & ~n4522 ;
  assign n4524 = ~\s3_msel_arb3_state_reg[1]/NET0131  & \s3_msel_arb3_state_reg[2]/NET0131  ;
  assign n4525 = \m1_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[2]/NET0131  ;
  assign n4526 = \rf_conf3_reg[3]/NET0131  & n4525 ;
  assign n4527 = \m0_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[0]/NET0131  ;
  assign n4528 = \rf_conf3_reg[1]/NET0131  & n4527 ;
  assign n4529 = ~n4526 & ~n4528 ;
  assign n4530 = \m3_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[6]/NET0131  ;
  assign n4531 = \rf_conf3_reg[7]/NET0131  & n4530 ;
  assign n4532 = \m2_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[4]/NET0131  ;
  assign n4533 = \rf_conf3_reg[5]/NET0131  & n4532 ;
  assign n4534 = ~n4531 & ~n4533 ;
  assign n4535 = n4529 & n4534 ;
  assign n4536 = \m5_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[10]/NET0131  ;
  assign n4537 = \rf_conf3_reg[11]/NET0131  & n4536 ;
  assign n4538 = \m7_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[14]/NET0131  ;
  assign n4539 = \rf_conf3_reg[15]/NET0131  & n4538 ;
  assign n4540 = \m6_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[12]/NET0131  ;
  assign n4541 = \rf_conf3_reg[13]/NET0131  & n4540 ;
  assign n4542 = ~n4539 & ~n4541 ;
  assign n4543 = ~n4537 & n4542 ;
  assign n4544 = ~n4535 & n4543 ;
  assign n4545 = n4524 & ~n4544 ;
  assign n4546 = ~n4535 & ~n4539 ;
  assign n4547 = \s3_msel_arb3_state_reg[1]/NET0131  & \s3_msel_arb3_state_reg[2]/NET0131  ;
  assign n4548 = ~n4546 & n4547 ;
  assign n4549 = \m4_s3_cyc_o_reg/NET0131  & \rf_conf3_reg[8]/NET0131  ;
  assign n4550 = \rf_conf3_reg[9]/NET0131  & n4549 ;
  assign n4551 = ~n4537 & ~n4550 ;
  assign n4552 = n4542 & n4551 ;
  assign n4553 = ~n4531 & ~n4552 ;
  assign n4554 = ~\s3_msel_arb3_state_reg[2]/NET0131  & ~n4526 ;
  assign n4555 = ~\s3_msel_arb3_state_reg[1]/NET0131  & ~n4533 ;
  assign n4556 = n4554 & n4555 ;
  assign n4557 = n4553 & n4556 ;
  assign n4558 = ~n4548 & ~n4557 ;
  assign n4559 = ~n4545 & n4558 ;
  assign n4560 = \s3_msel_arb3_state_reg[0]/NET0131  & ~n4559 ;
  assign n4561 = \rf_conf3_reg[5]/NET0131  & ~\s3_msel_arb3_state_reg[0]/NET0131  ;
  assign n4562 = n4532 & n4561 ;
  assign n4563 = ~\s3_msel_arb3_state_reg[1]/NET0131  & ~n4529 ;
  assign n4564 = ~n4562 & ~n4563 ;
  assign n4565 = n4553 & n4564 ;
  assign n4566 = ~\s3_msel_arb3_state_reg[2]/NET0131  & ~n4565 ;
  assign n4567 = \s3_msel_arb3_state_reg[1]/NET0131  & ~\s3_msel_arb3_state_reg[2]/NET0131  ;
  assign n4568 = \s3_msel_arb3_state_reg[0]/NET0131  & ~n4567 ;
  assign n4569 = ~n4535 & n4542 ;
  assign n4570 = ~n4547 & ~n4551 ;
  assign n4571 = n4569 & ~n4570 ;
  assign n4572 = ~n4568 & ~n4571 ;
  assign n4573 = ~n4566 & n4572 ;
  assign n4574 = ~n4560 & ~n4573 ;
  assign n4575 = \rf_conf5_reg[11]/NET0131  & n3183 ;
  assign n4576 = \rf_conf5_reg[9]/NET0131  & n3185 ;
  assign n4577 = ~n4575 & ~n4576 ;
  assign n4578 = \rf_conf5_reg[13]/NET0131  & n3190 ;
  assign n4579 = \rf_conf5_reg[15]/NET0131  & n3188 ;
  assign n4580 = ~n4578 & ~n4579 ;
  assign n4581 = n4577 & n4580 ;
  assign n4582 = \rf_conf5_reg[7]/NET0131  & n3200 ;
  assign n4583 = ~\s5_msel_arb2_state_reg[2]/NET0131  & ~n4582 ;
  assign n4584 = ~n4581 & n4583 ;
  assign n4585 = \rf_conf5_reg[5]/NET0131  & n3206 ;
  assign n4586 = \rf_conf5_reg[1]/NET0131  & ~\s5_msel_arb2_state_reg[1]/NET0131  ;
  assign n4587 = n3195 & n4586 ;
  assign n4588 = ~n4585 & ~n4587 ;
  assign n4589 = ~\s5_msel_arb2_state_reg[0]/NET0131  & ~n4588 ;
  assign n4590 = \rf_conf5_reg[3]/NET0131  & n3193 ;
  assign n4591 = ~n4585 & ~n4590 ;
  assign n4592 = ~\s5_msel_arb2_state_reg[1]/NET0131  & ~n4591 ;
  assign n4593 = ~n4589 & ~n4592 ;
  assign n4594 = n4584 & n4593 ;
  assign n4595 = ~n4582 & ~n4585 ;
  assign n4596 = \rf_conf5_reg[1]/NET0131  & n3195 ;
  assign n4597 = ~n4590 & ~n4596 ;
  assign n4598 = n4595 & n4597 ;
  assign n4599 = ~n4579 & ~n4598 ;
  assign n4600 = \rf_conf5_reg[9]/NET0131  & ~\s5_msel_arb2_state_reg[1]/NET0131  ;
  assign n4601 = n3185 & n4600 ;
  assign n4602 = ~n4578 & ~n4601 ;
  assign n4603 = ~\s5_msel_arb2_state_reg[0]/NET0131  & ~n4602 ;
  assign n4604 = ~n4575 & ~n4578 ;
  assign n4605 = ~\s5_msel_arb2_state_reg[1]/NET0131  & ~n4604 ;
  assign n4606 = ~n4603 & ~n4605 ;
  assign n4607 = n4599 & n4606 ;
  assign n4608 = \s5_msel_arb2_state_reg[2]/NET0131  & ~n4607 ;
  assign n4609 = ~n4594 & ~n4608 ;
  assign n4610 = \m5_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[10]/NET0131  ;
  assign n4611 = \rf_conf5_reg[11]/NET0131  & n4610 ;
  assign n4612 = \m4_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[8]/NET0131  ;
  assign n4613 = \rf_conf5_reg[9]/NET0131  & n4612 ;
  assign n4614 = ~n4611 & ~n4613 ;
  assign n4615 = ~\s5_msel_arb3_state_reg[0]/NET0131  & n4614 ;
  assign n4616 = \s5_msel_arb3_state_reg[0]/NET0131  & \s5_msel_arb3_state_reg[2]/NET0131  ;
  assign n4617 = ~\s5_msel_arb3_state_reg[1]/NET0131  & ~n4616 ;
  assign n4618 = \rf_conf5_reg[11]/NET0131  & ~\s5_msel_arb3_state_reg[1]/NET0131  ;
  assign n4619 = n4610 & n4618 ;
  assign n4620 = ~n4617 & ~n4619 ;
  assign n4621 = ~n4615 & ~n4620 ;
  assign n4622 = \m7_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[14]/NET0131  ;
  assign n4623 = \rf_conf5_reg[15]/NET0131  & n4622 ;
  assign n4624 = \m6_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[12]/NET0131  ;
  assign n4625 = \rf_conf5_reg[13]/NET0131  & n4624 ;
  assign n4626 = ~n4623 & ~n4625 ;
  assign n4627 = \m3_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[6]/NET0131  ;
  assign n4628 = \rf_conf5_reg[7]/NET0131  & n4627 ;
  assign n4629 = \m2_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[4]/NET0131  ;
  assign n4630 = \rf_conf5_reg[5]/NET0131  & n4629 ;
  assign n4631 = ~n4628 & ~n4630 ;
  assign n4632 = \m1_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[2]/NET0131  ;
  assign n4633 = \rf_conf5_reg[3]/NET0131  & n4632 ;
  assign n4634 = \m0_s5_cyc_o_reg/NET0131  & \rf_conf5_reg[0]/NET0131  ;
  assign n4635 = \rf_conf5_reg[1]/NET0131  & n4634 ;
  assign n4636 = ~n4633 & ~n4635 ;
  assign n4637 = n4631 & n4636 ;
  assign n4638 = n4626 & ~n4637 ;
  assign n4639 = ~n4621 & n4638 ;
  assign n4640 = ~\s5_msel_arb3_state_reg[0]/NET0131  & n4636 ;
  assign n4641 = ~\s5_msel_arb3_state_reg[1]/NET0131  & ~n4640 ;
  assign n4642 = n4614 & n4626 ;
  assign n4643 = \rf_conf5_reg[5]/NET0131  & ~\s5_msel_arb3_state_reg[0]/NET0131  ;
  assign n4644 = n4629 & n4643 ;
  assign n4645 = ~\s5_msel_arb3_state_reg[2]/NET0131  & ~n4644 ;
  assign n4646 = ~n4628 & n4645 ;
  assign n4647 = ~n4642 & n4646 ;
  assign n4648 = ~n4641 & n4647 ;
  assign n4649 = n4639 & ~n4648 ;
  assign n4650 = \s5_msel_arb3_state_reg[0]/NET0131  & \s5_msel_arb3_state_reg[1]/NET0131  ;
  assign n4651 = \s5_msel_arb3_state_reg[0]/NET0131  & ~n4630 ;
  assign n4652 = ~n4628 & ~n4633 ;
  assign n4653 = n4651 & n4652 ;
  assign n4654 = ~n4642 & n4653 ;
  assign n4655 = ~\s5_msel_arb3_state_reg[2]/NET0131  & ~n4654 ;
  assign n4656 = ~n4650 & ~n4655 ;
  assign n4657 = ~n4623 & ~n4637 ;
  assign n4658 = \s5_msel_arb3_state_reg[1]/NET0131  & \s5_msel_arb3_state_reg[2]/NET0131  ;
  assign n4659 = \s5_msel_arb3_state_reg[0]/NET0131  & n4658 ;
  assign n4660 = ~n4657 & n4659 ;
  assign n4661 = ~n4648 & ~n4660 ;
  assign n4662 = ~n4656 & n4661 ;
  assign n4663 = ~n4649 & ~n4662 ;
  assign n4664 = \m5_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[10]/NET0131  ;
  assign n4665 = \rf_conf6_reg[11]/NET0131  & n4664 ;
  assign n4666 = \m4_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[8]/NET0131  ;
  assign n4667 = \rf_conf6_reg[9]/NET0131  & n4666 ;
  assign n4668 = ~n4665 & ~n4667 ;
  assign n4669 = ~\s6_msel_arb3_state_reg[0]/NET0131  & n4668 ;
  assign n4670 = \s6_msel_arb3_state_reg[0]/NET0131  & \s6_msel_arb3_state_reg[2]/NET0131  ;
  assign n4671 = ~\s6_msel_arb3_state_reg[1]/NET0131  & ~n4670 ;
  assign n4672 = \rf_conf6_reg[11]/NET0131  & ~\s6_msel_arb3_state_reg[1]/NET0131  ;
  assign n4673 = n4664 & n4672 ;
  assign n4674 = ~n4671 & ~n4673 ;
  assign n4675 = ~n4669 & ~n4674 ;
  assign n4676 = \m7_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[14]/NET0131  ;
  assign n4677 = \rf_conf6_reg[15]/NET0131  & n4676 ;
  assign n4678 = \m6_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[12]/NET0131  ;
  assign n4679 = \rf_conf6_reg[13]/NET0131  & n4678 ;
  assign n4680 = ~n4677 & ~n4679 ;
  assign n4681 = \m3_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[6]/NET0131  ;
  assign n4682 = \rf_conf6_reg[7]/NET0131  & n4681 ;
  assign n4683 = \m2_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[4]/NET0131  ;
  assign n4684 = \rf_conf6_reg[5]/NET0131  & n4683 ;
  assign n4685 = ~n4682 & ~n4684 ;
  assign n4686 = \m1_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[2]/NET0131  ;
  assign n4687 = \rf_conf6_reg[3]/NET0131  & n4686 ;
  assign n4688 = \m0_s6_cyc_o_reg/NET0131  & \rf_conf6_reg[0]/NET0131  ;
  assign n4689 = \rf_conf6_reg[1]/NET0131  & n4688 ;
  assign n4690 = ~n4687 & ~n4689 ;
  assign n4691 = n4685 & n4690 ;
  assign n4692 = n4680 & ~n4691 ;
  assign n4693 = ~n4675 & n4692 ;
  assign n4694 = ~\s6_msel_arb3_state_reg[0]/NET0131  & n4690 ;
  assign n4695 = ~\s6_msel_arb3_state_reg[1]/NET0131  & ~n4694 ;
  assign n4696 = n4668 & n4680 ;
  assign n4697 = \rf_conf6_reg[5]/NET0131  & ~\s6_msel_arb3_state_reg[0]/NET0131  ;
  assign n4698 = n4683 & n4697 ;
  assign n4699 = ~\s6_msel_arb3_state_reg[2]/NET0131  & ~n4698 ;
  assign n4700 = ~n4682 & n4699 ;
  assign n4701 = ~n4696 & n4700 ;
  assign n4702 = ~n4695 & n4701 ;
  assign n4703 = n4693 & ~n4702 ;
  assign n4704 = \s6_msel_arb3_state_reg[0]/NET0131  & \s6_msel_arb3_state_reg[1]/NET0131  ;
  assign n4705 = \s6_msel_arb3_state_reg[0]/NET0131  & ~n4684 ;
  assign n4706 = ~n4682 & ~n4687 ;
  assign n4707 = n4705 & n4706 ;
  assign n4708 = ~n4696 & n4707 ;
  assign n4709 = ~\s6_msel_arb3_state_reg[2]/NET0131  & ~n4708 ;
  assign n4710 = ~n4704 & ~n4709 ;
  assign n4711 = ~n4677 & ~n4691 ;
  assign n4712 = \s6_msel_arb3_state_reg[1]/NET0131  & \s6_msel_arb3_state_reg[2]/NET0131  ;
  assign n4713 = \s6_msel_arb3_state_reg[0]/NET0131  & n4712 ;
  assign n4714 = ~n4711 & n4713 ;
  assign n4715 = ~n4702 & ~n4714 ;
  assign n4716 = ~n4710 & n4715 ;
  assign n4717 = ~n4703 & ~n4716 ;
  assign n4718 = \m5_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[10]/NET0131  ;
  assign n4719 = \rf_conf7_reg[11]/NET0131  & n4718 ;
  assign n4720 = \m4_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[8]/NET0131  ;
  assign n4721 = \rf_conf7_reg[9]/NET0131  & n4720 ;
  assign n4722 = ~n4719 & ~n4721 ;
  assign n4723 = ~\s7_msel_arb3_state_reg[0]/NET0131  & n4722 ;
  assign n4724 = \s7_msel_arb3_state_reg[0]/NET0131  & \s7_msel_arb3_state_reg[2]/NET0131  ;
  assign n4725 = ~\s7_msel_arb3_state_reg[1]/NET0131  & ~n4724 ;
  assign n4726 = \rf_conf7_reg[11]/NET0131  & ~\s7_msel_arb3_state_reg[1]/NET0131  ;
  assign n4727 = n4718 & n4726 ;
  assign n4728 = ~n4725 & ~n4727 ;
  assign n4729 = ~n4723 & ~n4728 ;
  assign n4730 = \m7_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[14]/NET0131  ;
  assign n4731 = \rf_conf7_reg[15]/NET0131  & n4730 ;
  assign n4732 = \m6_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[12]/NET0131  ;
  assign n4733 = \rf_conf7_reg[13]/NET0131  & n4732 ;
  assign n4734 = ~n4731 & ~n4733 ;
  assign n4735 = \m3_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[6]/NET0131  ;
  assign n4736 = \rf_conf7_reg[7]/NET0131  & n4735 ;
  assign n4737 = \m2_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[4]/NET0131  ;
  assign n4738 = \rf_conf7_reg[5]/NET0131  & n4737 ;
  assign n4739 = ~n4736 & ~n4738 ;
  assign n4740 = \m1_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[2]/NET0131  ;
  assign n4741 = \rf_conf7_reg[3]/NET0131  & n4740 ;
  assign n4742 = \m0_s7_cyc_o_reg/NET0131  & \rf_conf7_reg[0]/NET0131  ;
  assign n4743 = \rf_conf7_reg[1]/NET0131  & n4742 ;
  assign n4744 = ~n4741 & ~n4743 ;
  assign n4745 = n4739 & n4744 ;
  assign n4746 = n4734 & ~n4745 ;
  assign n4747 = ~n4729 & n4746 ;
  assign n4748 = ~\s7_msel_arb3_state_reg[0]/NET0131  & n4744 ;
  assign n4749 = ~\s7_msel_arb3_state_reg[1]/NET0131  & ~n4748 ;
  assign n4750 = n4722 & n4734 ;
  assign n4751 = \rf_conf7_reg[5]/NET0131  & ~\s7_msel_arb3_state_reg[0]/NET0131  ;
  assign n4752 = n4737 & n4751 ;
  assign n4753 = ~\s7_msel_arb3_state_reg[2]/NET0131  & ~n4752 ;
  assign n4754 = ~n4736 & n4753 ;
  assign n4755 = ~n4750 & n4754 ;
  assign n4756 = ~n4749 & n4755 ;
  assign n4757 = n4747 & ~n4756 ;
  assign n4758 = \s7_msel_arb3_state_reg[0]/NET0131  & \s7_msel_arb3_state_reg[1]/NET0131  ;
  assign n4759 = \s7_msel_arb3_state_reg[0]/NET0131  & ~n4738 ;
  assign n4760 = ~n4736 & ~n4741 ;
  assign n4761 = n4759 & n4760 ;
  assign n4762 = ~n4750 & n4761 ;
  assign n4763 = ~\s7_msel_arb3_state_reg[2]/NET0131  & ~n4762 ;
  assign n4764 = ~n4758 & ~n4763 ;
  assign n4765 = ~n4731 & ~n4745 ;
  assign n4766 = \s7_msel_arb3_state_reg[1]/NET0131  & \s7_msel_arb3_state_reg[2]/NET0131  ;
  assign n4767 = \s7_msel_arb3_state_reg[0]/NET0131  & n4766 ;
  assign n4768 = ~n4765 & n4767 ;
  assign n4769 = ~n4756 & ~n4768 ;
  assign n4770 = ~n4764 & n4769 ;
  assign n4771 = ~n4757 & ~n4770 ;
  assign n4772 = ~\s8_msel_arb3_state_reg[1]/NET0131  & \s8_msel_arb3_state_reg[2]/NET0131  ;
  assign n4773 = \m1_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[2]/NET0131  ;
  assign n4774 = \rf_conf8_reg[3]/NET0131  & n4773 ;
  assign n4775 = \m0_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[0]/NET0131  ;
  assign n4776 = \rf_conf8_reg[1]/NET0131  & n4775 ;
  assign n4777 = ~n4774 & ~n4776 ;
  assign n4778 = \m3_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[6]/NET0131  ;
  assign n4779 = \rf_conf8_reg[7]/NET0131  & n4778 ;
  assign n4780 = \m2_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[4]/NET0131  ;
  assign n4781 = \rf_conf8_reg[5]/NET0131  & n4780 ;
  assign n4782 = ~n4779 & ~n4781 ;
  assign n4783 = n4777 & n4782 ;
  assign n4784 = \m5_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[10]/NET0131  ;
  assign n4785 = \rf_conf8_reg[11]/NET0131  & n4784 ;
  assign n4786 = \m7_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[14]/NET0131  ;
  assign n4787 = \rf_conf8_reg[15]/NET0131  & n4786 ;
  assign n4788 = \m6_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[12]/NET0131  ;
  assign n4789 = \rf_conf8_reg[13]/NET0131  & n4788 ;
  assign n4790 = ~n4787 & ~n4789 ;
  assign n4791 = ~n4785 & n4790 ;
  assign n4792 = ~n4783 & n4791 ;
  assign n4793 = n4772 & ~n4792 ;
  assign n4794 = ~n4783 & ~n4787 ;
  assign n4795 = \s8_msel_arb3_state_reg[1]/NET0131  & \s8_msel_arb3_state_reg[2]/NET0131  ;
  assign n4796 = ~n4794 & n4795 ;
  assign n4797 = \m4_s8_cyc_o_reg/NET0131  & \rf_conf8_reg[8]/NET0131  ;
  assign n4798 = \rf_conf8_reg[9]/NET0131  & n4797 ;
  assign n4799 = ~n4785 & ~n4798 ;
  assign n4800 = n4790 & n4799 ;
  assign n4801 = ~n4779 & ~n4800 ;
  assign n4802 = ~\s8_msel_arb3_state_reg[2]/NET0131  & ~n4774 ;
  assign n4803 = ~\s8_msel_arb3_state_reg[1]/NET0131  & ~n4781 ;
  assign n4804 = n4802 & n4803 ;
  assign n4805 = n4801 & n4804 ;
  assign n4806 = ~n4796 & ~n4805 ;
  assign n4807 = ~n4793 & n4806 ;
  assign n4808 = \s8_msel_arb3_state_reg[0]/NET0131  & ~n4807 ;
  assign n4809 = \rf_conf8_reg[5]/NET0131  & ~\s8_msel_arb3_state_reg[0]/NET0131  ;
  assign n4810 = n4780 & n4809 ;
  assign n4811 = ~\s8_msel_arb3_state_reg[1]/NET0131  & ~n4777 ;
  assign n4812 = ~n4810 & ~n4811 ;
  assign n4813 = n4801 & n4812 ;
  assign n4814 = ~\s8_msel_arb3_state_reg[2]/NET0131  & ~n4813 ;
  assign n4815 = \s8_msel_arb3_state_reg[1]/NET0131  & ~\s8_msel_arb3_state_reg[2]/NET0131  ;
  assign n4816 = \s8_msel_arb3_state_reg[0]/NET0131  & ~n4815 ;
  assign n4817 = ~n4783 & n4790 ;
  assign n4818 = ~n4795 & ~n4799 ;
  assign n4819 = n4817 & ~n4818 ;
  assign n4820 = ~n4816 & ~n4819 ;
  assign n4821 = ~n4814 & n4820 ;
  assign n4822 = ~n4808 & ~n4821 ;
  assign n4823 = \m5_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[10]/NET0131  ;
  assign n4824 = \rf_conf0_reg[11]/NET0131  & n4823 ;
  assign n4825 = \m4_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[8]/NET0131  ;
  assign n4826 = \rf_conf0_reg[9]/NET0131  & n4825 ;
  assign n4827 = ~n4824 & ~n4826 ;
  assign n4828 = ~\s0_msel_arb3_state_reg[0]/NET0131  & n4827 ;
  assign n4829 = \s0_msel_arb3_state_reg[0]/NET0131  & \s0_msel_arb3_state_reg[2]/NET0131  ;
  assign n4830 = ~\s0_msel_arb3_state_reg[1]/NET0131  & ~n4829 ;
  assign n4831 = \rf_conf0_reg[11]/NET0131  & ~\s0_msel_arb3_state_reg[1]/NET0131  ;
  assign n4832 = n4823 & n4831 ;
  assign n4833 = ~n4830 & ~n4832 ;
  assign n4834 = ~n4828 & ~n4833 ;
  assign n4835 = \m7_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[14]/NET0131  ;
  assign n4836 = \rf_conf0_reg[15]/NET0131  & n4835 ;
  assign n4837 = \m6_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[12]/NET0131  ;
  assign n4838 = \rf_conf0_reg[13]/NET0131  & n4837 ;
  assign n4839 = ~n4836 & ~n4838 ;
  assign n4840 = \m3_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[6]/NET0131  ;
  assign n4841 = \rf_conf0_reg[7]/NET0131  & n4840 ;
  assign n4842 = \m2_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[4]/NET0131  ;
  assign n4843 = \rf_conf0_reg[5]/NET0131  & n4842 ;
  assign n4844 = ~n4841 & ~n4843 ;
  assign n4845 = \m1_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[2]/NET0131  ;
  assign n4846 = \rf_conf0_reg[3]/NET0131  & n4845 ;
  assign n4847 = \m0_s0_cyc_o_reg/NET0131  & \rf_conf0_reg[0]/NET0131  ;
  assign n4848 = \rf_conf0_reg[1]/NET0131  & n4847 ;
  assign n4849 = ~n4846 & ~n4848 ;
  assign n4850 = n4844 & n4849 ;
  assign n4851 = n4839 & ~n4850 ;
  assign n4852 = ~n4834 & n4851 ;
  assign n4853 = ~\s0_msel_arb3_state_reg[0]/NET0131  & n4849 ;
  assign n4854 = ~\s0_msel_arb3_state_reg[1]/NET0131  & ~n4853 ;
  assign n4855 = n4827 & n4839 ;
  assign n4856 = \rf_conf0_reg[5]/NET0131  & ~\s0_msel_arb3_state_reg[0]/NET0131  ;
  assign n4857 = n4842 & n4856 ;
  assign n4858 = ~\s0_msel_arb3_state_reg[2]/NET0131  & ~n4857 ;
  assign n4859 = ~n4841 & n4858 ;
  assign n4860 = ~n4855 & n4859 ;
  assign n4861 = ~n4854 & n4860 ;
  assign n4862 = n4852 & ~n4861 ;
  assign n4863 = \s0_msel_arb3_state_reg[0]/NET0131  & \s0_msel_arb3_state_reg[1]/NET0131  ;
  assign n4864 = \s0_msel_arb3_state_reg[0]/NET0131  & ~n4843 ;
  assign n4865 = ~n4841 & ~n4846 ;
  assign n4866 = n4864 & n4865 ;
  assign n4867 = ~n4855 & n4866 ;
  assign n4868 = ~\s0_msel_arb3_state_reg[2]/NET0131  & ~n4867 ;
  assign n4869 = ~n4863 & ~n4868 ;
  assign n4870 = ~n4836 & ~n4850 ;
  assign n4871 = \s0_msel_arb3_state_reg[1]/NET0131  & \s0_msel_arb3_state_reg[2]/NET0131  ;
  assign n4872 = \s0_msel_arb3_state_reg[0]/NET0131  & n4871 ;
  assign n4873 = ~n4870 & n4872 ;
  assign n4874 = ~n4861 & ~n4873 ;
  assign n4875 = ~n4869 & n4874 ;
  assign n4876 = ~n4862 & ~n4875 ;
  assign n4877 = ~\rf_conf10_reg[11]/NET0131  & n4193 ;
  assign n4878 = ~\s10_msel_arb1_state_reg[1]/NET0131  & n4877 ;
  assign n4879 = ~\rf_conf10_reg[9]/NET0131  & n4195 ;
  assign n4880 = ~\s10_msel_arb1_state_reg[0]/NET0131  & ~\s10_msel_arb1_state_reg[1]/NET0131  ;
  assign n4881 = n4879 & n4880 ;
  assign n4882 = ~n4878 & ~n4881 ;
  assign n4883 = ~\rf_conf10_reg[5]/NET0131  & n4212 ;
  assign n4884 = ~\rf_conf10_reg[7]/NET0131  & n4210 ;
  assign n4885 = ~n4883 & ~n4884 ;
  assign n4886 = ~\rf_conf10_reg[3]/NET0131  & n4215 ;
  assign n4887 = ~\rf_conf10_reg[1]/NET0131  & n4217 ;
  assign n4888 = ~n4886 & ~n4887 ;
  assign n4889 = n4885 & n4888 ;
  assign n4890 = ~\rf_conf10_reg[15]/NET0131  & n4205 ;
  assign n4891 = ~\rf_conf10_reg[13]/NET0131  & n4207 ;
  assign n4892 = \s10_msel_arb1_state_reg[0]/NET0131  & \s10_msel_arb1_state_reg[1]/NET0131  ;
  assign n4893 = n4891 & ~n4892 ;
  assign n4894 = ~n4890 & ~n4893 ;
  assign n4895 = ~n4889 & n4894 ;
  assign n4896 = n4882 & n4895 ;
  assign n4897 = \s10_msel_arb1_state_reg[2]/NET0131  & ~n4896 ;
  assign n4898 = ~\rf_conf10_reg[1]/NET0131  & ~\s10_msel_arb1_state_reg[0]/NET0131  ;
  assign n4899 = n4217 & n4898 ;
  assign n4900 = ~n4886 & ~n4899 ;
  assign n4901 = ~\s10_msel_arb1_state_reg[1]/NET0131  & ~n4900 ;
  assign n4902 = ~n4877 & ~n4879 ;
  assign n4903 = ~n4890 & ~n4891 ;
  assign n4904 = n4902 & n4903 ;
  assign n4905 = n4883 & ~n4892 ;
  assign n4906 = ~\s10_msel_arb1_state_reg[2]/NET0131  & ~n4884 ;
  assign n4907 = ~n4905 & n4906 ;
  assign n4908 = ~n4904 & n4907 ;
  assign n4909 = ~n4901 & n4908 ;
  assign n4910 = ~n4897 & ~n4909 ;
  assign n4911 = ~\rf_conf11_reg[7]/NET0131  & n4288 ;
  assign n4912 = \s11_msel_arb1_state_reg[1]/NET0131  & ~\s11_msel_arb1_state_reg[2]/NET0131  ;
  assign n4913 = \s11_msel_arb1_state_reg[0]/NET0131  & n4912 ;
  assign n4914 = ~\rf_conf11_reg[15]/NET0131  & n4296 ;
  assign n4915 = ~\rf_conf11_reg[13]/NET0131  & n4298 ;
  assign n4916 = ~n4914 & ~n4915 ;
  assign n4917 = ~\rf_conf11_reg[9]/NET0131  & n4307 ;
  assign n4918 = ~\rf_conf11_reg[11]/NET0131  & n4294 ;
  assign n4919 = ~n4917 & ~n4918 ;
  assign n4920 = n4916 & n4919 ;
  assign n4921 = n4913 & ~n4920 ;
  assign n4922 = ~n4911 & n4921 ;
  assign n4923 = ~\rf_conf11_reg[1]/NET0131  & n4285 ;
  assign n4924 = \s11_msel_arb1_state_reg[1]/NET0131  & \s11_msel_arb1_state_reg[2]/NET0131  ;
  assign n4925 = ~n4923 & n4924 ;
  assign n4926 = ~\s11_msel_arb1_state_reg[0]/NET0131  & \s11_msel_arb1_state_reg[1]/NET0131  ;
  assign n4927 = ~\rf_conf11_reg[1]/NET0131  & ~\s11_msel_arb1_state_reg[0]/NET0131  ;
  assign n4928 = n4285 & n4927 ;
  assign n4929 = ~n4926 & ~n4928 ;
  assign n4930 = ~\s11_msel_arb1_state_reg[2]/NET0131  & n4929 ;
  assign n4931 = ~n4920 & n4930 ;
  assign n4932 = ~n4925 & ~n4931 ;
  assign n4933 = ~\rf_conf11_reg[5]/NET0131  & n4290 ;
  assign n4934 = ~\rf_conf11_reg[3]/NET0131  & n4283 ;
  assign n4935 = ~n4933 & ~n4934 ;
  assign n4936 = ~n4911 & n4935 ;
  assign n4937 = ~n4932 & n4936 ;
  assign n4938 = ~n4922 & ~n4937 ;
  assign n4939 = ~n4911 & ~n4933 ;
  assign n4940 = n4912 & n4939 ;
  assign n4941 = ~n4920 & n4940 ;
  assign n4942 = ~\s11_msel_arb1_state_reg[0]/NET0131  & n4941 ;
  assign n4943 = ~n4923 & ~n4934 ;
  assign n4944 = n4939 & n4943 ;
  assign n4945 = n4920 & ~n4944 ;
  assign n4946 = ~\s11_msel_arb1_state_reg[1]/NET0131  & \s11_msel_arb1_state_reg[2]/NET0131  ;
  assign n4947 = ~\s11_msel_arb1_state_reg[0]/NET0131  & n4946 ;
  assign n4948 = ~n4945 & n4947 ;
  assign n4949 = ~n4942 & ~n4948 ;
  assign n4950 = ~\rf_conf11_reg[13]/NET0131  & ~\s11_msel_arb1_state_reg[0]/NET0131  ;
  assign n4951 = n4298 & n4950 ;
  assign n4952 = ~n4914 & ~n4951 ;
  assign n4953 = \s11_msel_arb1_state_reg[1]/NET0131  & ~n4952 ;
  assign n4954 = \s11_msel_arb1_state_reg[2]/NET0131  & n4953 ;
  assign n4955 = n4916 & ~n4918 ;
  assign n4956 = ~n4944 & n4955 ;
  assign n4957 = \s11_msel_arb1_state_reg[0]/NET0131  & ~\s11_msel_arb1_state_reg[1]/NET0131  ;
  assign n4958 = \s11_msel_arb1_state_reg[2]/NET0131  & n4957 ;
  assign n4959 = ~n4956 & n4958 ;
  assign n4960 = ~n4954 & ~n4959 ;
  assign n4961 = n4949 & n4960 ;
  assign n4962 = n4938 & n4961 ;
  assign n4963 = ~\rf_conf12_reg[3]/NET0131  & n4355 ;
  assign n4964 = ~\rf_conf12_reg[1]/NET0131  & ~\s12_msel_arb1_state_reg[0]/NET0131  ;
  assign n4965 = n4357 & n4964 ;
  assign n4966 = ~n4963 & ~n4965 ;
  assign n4967 = ~\s12_msel_arb1_state_reg[1]/NET0131  & ~n4966 ;
  assign n4968 = ~\rf_conf12_reg[15]/NET0131  & n4345 ;
  assign n4969 = ~\rf_conf12_reg[13]/NET0131  & n4347 ;
  assign n4970 = ~n4968 & ~n4969 ;
  assign n4971 = ~\rf_conf12_reg[9]/NET0131  & n4335 ;
  assign n4972 = ~\rf_conf12_reg[11]/NET0131  & n4333 ;
  assign n4973 = ~n4971 & ~n4972 ;
  assign n4974 = n4970 & n4973 ;
  assign n4975 = \s12_msel_arb1_state_reg[0]/NET0131  & \s12_msel_arb1_state_reg[1]/NET0131  ;
  assign n4976 = ~\rf_conf12_reg[5]/NET0131  & n4352 ;
  assign n4977 = ~n4975 & n4976 ;
  assign n4978 = ~\rf_conf12_reg[7]/NET0131  & n4350 ;
  assign n4979 = ~n4977 & ~n4978 ;
  assign n4980 = ~n4974 & n4979 ;
  assign n4981 = ~n4967 & n4980 ;
  assign n4982 = ~\s12_msel_arb1_state_reg[2]/NET0131  & ~n4981 ;
  assign n4983 = ~\rf_conf12_reg[13]/NET0131  & ~\s12_msel_arb1_state_reg[0]/NET0131  ;
  assign n4984 = n4347 & n4983 ;
  assign n4985 = \s12_msel_arb1_state_reg[1]/NET0131  & ~n4984 ;
  assign n4986 = ~\rf_conf12_reg[9]/NET0131  & ~\s12_msel_arb1_state_reg[0]/NET0131  ;
  assign n4987 = n4335 & n4986 ;
  assign n4988 = ~n4972 & ~n4987 ;
  assign n4989 = ~n4969 & n4988 ;
  assign n4990 = ~n4985 & ~n4989 ;
  assign n4991 = \s12_msel_arb1_state_reg[2]/NET0131  & ~n4968 ;
  assign n4992 = ~\rf_conf12_reg[1]/NET0131  & n4357 ;
  assign n4993 = ~n4963 & ~n4992 ;
  assign n4994 = ~n4976 & ~n4978 ;
  assign n4995 = n4993 & n4994 ;
  assign n4996 = n4991 & ~n4995 ;
  assign n4997 = ~n4990 & n4996 ;
  assign n4998 = ~n4982 & ~n4997 ;
  assign n4999 = ~\rf_conf13_reg[11]/NET0131  & n3848 ;
  assign n5000 = ~\s13_msel_arb1_state_reg[1]/NET0131  & n4999 ;
  assign n5001 = ~\rf_conf13_reg[9]/NET0131  & n3850 ;
  assign n5002 = ~\s13_msel_arb1_state_reg[0]/NET0131  & ~\s13_msel_arb1_state_reg[1]/NET0131  ;
  assign n5003 = n5001 & n5002 ;
  assign n5004 = ~n5000 & ~n5003 ;
  assign n5005 = ~\rf_conf13_reg[5]/NET0131  & n3867 ;
  assign n5006 = ~\rf_conf13_reg[7]/NET0131  & n3865 ;
  assign n5007 = ~n5005 & ~n5006 ;
  assign n5008 = ~\rf_conf13_reg[3]/NET0131  & n3870 ;
  assign n5009 = ~\rf_conf13_reg[1]/NET0131  & n3872 ;
  assign n5010 = ~n5008 & ~n5009 ;
  assign n5011 = n5007 & n5010 ;
  assign n5012 = ~\rf_conf13_reg[15]/NET0131  & n3860 ;
  assign n5013 = ~\rf_conf13_reg[13]/NET0131  & n3862 ;
  assign n5014 = \s13_msel_arb1_state_reg[0]/NET0131  & \s13_msel_arb1_state_reg[1]/NET0131  ;
  assign n5015 = n5013 & ~n5014 ;
  assign n5016 = ~n5012 & ~n5015 ;
  assign n5017 = ~n5011 & n5016 ;
  assign n5018 = n5004 & n5017 ;
  assign n5019 = \s13_msel_arb1_state_reg[2]/NET0131  & ~n5018 ;
  assign n5020 = ~\rf_conf13_reg[1]/NET0131  & ~\s13_msel_arb1_state_reg[0]/NET0131  ;
  assign n5021 = n3872 & n5020 ;
  assign n5022 = ~n5008 & ~n5021 ;
  assign n5023 = ~\s13_msel_arb1_state_reg[1]/NET0131  & ~n5022 ;
  assign n5024 = ~n4999 & ~n5001 ;
  assign n5025 = ~n5012 & ~n5013 ;
  assign n5026 = n5024 & n5025 ;
  assign n5027 = n5005 & ~n5014 ;
  assign n5028 = ~\s13_msel_arb1_state_reg[2]/NET0131  & ~n5006 ;
  assign n5029 = ~n5027 & n5028 ;
  assign n5030 = ~n5026 & n5029 ;
  assign n5031 = ~n5023 & n5030 ;
  assign n5032 = ~n5019 & ~n5031 ;
  assign n5033 = ~\rf_conf14_reg[13]/NET0131  & n4403 ;
  assign n5034 = ~\rf_conf14_reg[15]/NET0131  & n4401 ;
  assign n5035 = ~n5033 & ~n5034 ;
  assign n5036 = ~\rf_conf14_reg[9]/NET0131  & n4412 ;
  assign n5037 = ~\rf_conf14_reg[11]/NET0131  & n4399 ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5039 = n5035 & n5038 ;
  assign n5040 = ~\s14_msel_arb1_state_reg[1]/NET0131  & \s14_msel_arb1_state_reg[2]/NET0131  ;
  assign n5041 = ~\s14_msel_arb1_state_reg[0]/NET0131  & n5040 ;
  assign n5042 = ~\rf_conf14_reg[7]/NET0131  & n4393 ;
  assign n5043 = ~\s14_msel_arb1_state_reg[2]/NET0131  & ~n5042 ;
  assign n5044 = ~n5041 & ~n5043 ;
  assign n5045 = ~\rf_conf14_reg[1]/NET0131  & ~\s14_msel_arb1_state_reg[0]/NET0131  ;
  assign n5046 = n4390 & n5045 ;
  assign n5047 = ~\rf_conf14_reg[5]/NET0131  & n4395 ;
  assign n5048 = ~\rf_conf14_reg[3]/NET0131  & n4388 ;
  assign n5049 = ~n5047 & ~n5048 ;
  assign n5050 = ~n5046 & n5049 ;
  assign n5051 = ~\rf_conf14_reg[5]/NET0131  & ~\s14_msel_arb1_state_reg[0]/NET0131  ;
  assign n5052 = n4395 & n5051 ;
  assign n5053 = \s14_msel_arb1_state_reg[1]/NET0131  & ~n5052 ;
  assign n5054 = ~n5041 & ~n5053 ;
  assign n5055 = ~n5050 & n5054 ;
  assign n5056 = ~n5044 & ~n5055 ;
  assign n5057 = ~n5039 & n5056 ;
  assign n5058 = ~\rf_conf14_reg[1]/NET0131  & n4390 ;
  assign n5059 = ~n5048 & ~n5058 ;
  assign n5060 = ~n5042 & ~n5047 ;
  assign n5061 = n5059 & n5060 ;
  assign n5062 = \s14_msel_arb1_state_reg[1]/NET0131  & ~n5035 ;
  assign n5063 = ~\s14_msel_arb1_state_reg[0]/NET0131  & ~n5062 ;
  assign n5064 = ~n5033 & ~n5037 ;
  assign n5065 = \s14_msel_arb1_state_reg[0]/NET0131  & \s14_msel_arb1_state_reg[1]/NET0131  ;
  assign n5066 = ~n5064 & ~n5065 ;
  assign n5067 = ~n5034 & ~n5066 ;
  assign n5068 = ~n5063 & ~n5067 ;
  assign n5069 = ~n5061 & ~n5068 ;
  assign n5070 = \s14_msel_arb1_state_reg[2]/NET0131  & ~n5069 ;
  assign n5071 = ~n5057 & ~n5070 ;
  assign n5072 = ~\rf_conf1_reg[13]/NET0131  & n4489 ;
  assign n5073 = ~\rf_conf1_reg[15]/NET0131  & n4487 ;
  assign n5074 = ~n5072 & ~n5073 ;
  assign n5075 = ~\rf_conf1_reg[9]/NET0131  & n4498 ;
  assign n5076 = ~\rf_conf1_reg[11]/NET0131  & n4485 ;
  assign n5077 = ~n5075 & ~n5076 ;
  assign n5078 = n5074 & n5077 ;
  assign n5079 = ~\s1_msel_arb1_state_reg[1]/NET0131  & \s1_msel_arb1_state_reg[2]/NET0131  ;
  assign n5080 = ~\s1_msel_arb1_state_reg[0]/NET0131  & n5079 ;
  assign n5081 = ~\rf_conf1_reg[7]/NET0131  & n4479 ;
  assign n5082 = ~\s1_msel_arb1_state_reg[2]/NET0131  & ~n5081 ;
  assign n5083 = ~n5080 & ~n5082 ;
  assign n5084 = ~\rf_conf1_reg[1]/NET0131  & ~\s1_msel_arb1_state_reg[0]/NET0131  ;
  assign n5085 = n4476 & n5084 ;
  assign n5086 = ~\rf_conf1_reg[5]/NET0131  & n4481 ;
  assign n5087 = ~\rf_conf1_reg[3]/NET0131  & n4474 ;
  assign n5088 = ~n5086 & ~n5087 ;
  assign n5089 = ~n5085 & n5088 ;
  assign n5090 = ~\rf_conf1_reg[5]/NET0131  & ~\s1_msel_arb1_state_reg[0]/NET0131  ;
  assign n5091 = n4481 & n5090 ;
  assign n5092 = \s1_msel_arb1_state_reg[1]/NET0131  & ~n5091 ;
  assign n5093 = ~n5080 & ~n5092 ;
  assign n5094 = ~n5089 & n5093 ;
  assign n5095 = ~n5083 & ~n5094 ;
  assign n5096 = ~n5078 & n5095 ;
  assign n5097 = ~\rf_conf1_reg[1]/NET0131  & n4476 ;
  assign n5098 = ~n5087 & ~n5097 ;
  assign n5099 = ~n5081 & ~n5086 ;
  assign n5100 = n5098 & n5099 ;
  assign n5101 = \s1_msel_arb1_state_reg[1]/NET0131  & ~n5074 ;
  assign n5102 = ~\s1_msel_arb1_state_reg[0]/NET0131  & ~n5101 ;
  assign n5103 = ~n5072 & ~n5076 ;
  assign n5104 = \s1_msel_arb1_state_reg[0]/NET0131  & \s1_msel_arb1_state_reg[1]/NET0131  ;
  assign n5105 = ~n5103 & ~n5104 ;
  assign n5106 = ~n5073 & ~n5105 ;
  assign n5107 = ~n5102 & ~n5106 ;
  assign n5108 = ~n5100 & ~n5107 ;
  assign n5109 = \s1_msel_arb1_state_reg[2]/NET0131  & ~n5108 ;
  assign n5110 = ~n5096 & ~n5109 ;
  assign n5111 = ~\rf_conf2_reg[11]/NET0131  & n3948 ;
  assign n5112 = ~\s2_msel_arb1_state_reg[1]/NET0131  & n5111 ;
  assign n5113 = ~\rf_conf2_reg[9]/NET0131  & n3950 ;
  assign n5114 = ~\s2_msel_arb1_state_reg[0]/NET0131  & ~\s2_msel_arb1_state_reg[1]/NET0131  ;
  assign n5115 = n5113 & n5114 ;
  assign n5116 = ~n5112 & ~n5115 ;
  assign n5117 = ~\rf_conf2_reg[5]/NET0131  & n3967 ;
  assign n5118 = ~\rf_conf2_reg[7]/NET0131  & n3965 ;
  assign n5119 = ~n5117 & ~n5118 ;
  assign n5120 = ~\rf_conf2_reg[3]/NET0131  & n3970 ;
  assign n5121 = ~\rf_conf2_reg[1]/NET0131  & n3972 ;
  assign n5122 = ~n5120 & ~n5121 ;
  assign n5123 = n5119 & n5122 ;
  assign n5124 = ~\rf_conf2_reg[15]/NET0131  & n3960 ;
  assign n5125 = ~\rf_conf2_reg[13]/NET0131  & n3962 ;
  assign n5126 = \s2_msel_arb1_state_reg[0]/NET0131  & \s2_msel_arb1_state_reg[1]/NET0131  ;
  assign n5127 = n5125 & ~n5126 ;
  assign n5128 = ~n5124 & ~n5127 ;
  assign n5129 = ~n5123 & n5128 ;
  assign n5130 = n5116 & n5129 ;
  assign n5131 = \s2_msel_arb1_state_reg[2]/NET0131  & ~n5130 ;
  assign n5132 = ~\rf_conf2_reg[1]/NET0131  & ~\s2_msel_arb1_state_reg[0]/NET0131  ;
  assign n5133 = n3972 & n5132 ;
  assign n5134 = ~n5120 & ~n5133 ;
  assign n5135 = ~\s2_msel_arb1_state_reg[1]/NET0131  & ~n5134 ;
  assign n5136 = ~n5111 & ~n5113 ;
  assign n5137 = ~n5124 & ~n5125 ;
  assign n5138 = n5136 & n5137 ;
  assign n5139 = n5117 & ~n5126 ;
  assign n5140 = ~\s2_msel_arb1_state_reg[2]/NET0131  & ~n5118 ;
  assign n5141 = ~n5139 & n5140 ;
  assign n5142 = ~n5138 & n5141 ;
  assign n5143 = ~n5135 & n5142 ;
  assign n5144 = ~n5131 & ~n5143 ;
  assign n5145 = ~\s3_msel_arb1_state_reg[0]/NET0131  & \s3_msel_arb1_state_reg[1]/NET0131  ;
  assign n5146 = ~\rf_conf3_reg[15]/NET0131  & n4538 ;
  assign n5147 = ~\rf_conf3_reg[13]/NET0131  & n4540 ;
  assign n5148 = ~n5146 & ~n5147 ;
  assign n5149 = \s3_msel_arb1_state_reg[2]/NET0131  & ~n5148 ;
  assign n5150 = ~\rf_conf3_reg[9]/NET0131  & n4549 ;
  assign n5151 = ~\rf_conf3_reg[11]/NET0131  & n4536 ;
  assign n5152 = ~n5150 & ~n5151 ;
  assign n5153 = n5148 & n5152 ;
  assign n5154 = ~\s3_msel_arb1_state_reg[2]/NET0131  & n5153 ;
  assign n5155 = ~\rf_conf3_reg[5]/NET0131  & n4532 ;
  assign n5156 = ~\rf_conf3_reg[7]/NET0131  & n4530 ;
  assign n5157 = ~n5155 & ~n5156 ;
  assign n5158 = ~\rf_conf3_reg[3]/NET0131  & n4525 ;
  assign n5159 = ~\rf_conf3_reg[1]/NET0131  & n4527 ;
  assign n5160 = ~n5158 & ~n5159 ;
  assign n5161 = \s3_msel_arb1_state_reg[2]/NET0131  & ~n5160 ;
  assign n5162 = n5157 & ~n5161 ;
  assign n5163 = ~n5154 & n5162 ;
  assign n5164 = ~n5149 & ~n5163 ;
  assign n5165 = n5145 & ~n5164 ;
  assign n5166 = ~\s3_msel_arb1_state_reg[2]/NET0131  & ~n5156 ;
  assign n5167 = ~n5153 & n5166 ;
  assign n5168 = ~\rf_conf3_reg[1]/NET0131  & ~\s3_msel_arb1_state_reg[0]/NET0131  ;
  assign n5169 = n4527 & n5168 ;
  assign n5170 = ~n5145 & ~n5169 ;
  assign n5171 = ~n5155 & ~n5158 ;
  assign n5172 = ~\s3_msel_arb1_state_reg[1]/NET0131  & ~n5171 ;
  assign n5173 = n5170 & ~n5172 ;
  assign n5174 = n5167 & n5173 ;
  assign n5175 = ~\rf_conf3_reg[9]/NET0131  & ~\s3_msel_arb1_state_reg[0]/NET0131  ;
  assign n5176 = n4549 & n5175 ;
  assign n5177 = ~n5147 & ~n5151 ;
  assign n5178 = ~n5176 & n5177 ;
  assign n5179 = ~\s3_msel_arb1_state_reg[1]/NET0131  & ~n5178 ;
  assign n5180 = n5157 & n5160 ;
  assign n5181 = ~n5146 & ~n5180 ;
  assign n5182 = ~n5179 & n5181 ;
  assign n5183 = \s3_msel_arb1_state_reg[2]/NET0131  & ~n5145 ;
  assign n5184 = ~n5182 & n5183 ;
  assign n5185 = ~n5174 & ~n5184 ;
  assign n5186 = ~n5165 & n5185 ;
  assign n5187 = ~\rf_conf4_reg[13]/NET0131  & n4053 ;
  assign n5188 = ~\rf_conf4_reg[15]/NET0131  & n4051 ;
  assign n5189 = ~n5187 & ~n5188 ;
  assign n5190 = ~\rf_conf4_reg[9]/NET0131  & n4062 ;
  assign n5191 = ~\rf_conf4_reg[11]/NET0131  & n4049 ;
  assign n5192 = ~n5190 & ~n5191 ;
  assign n5193 = n5189 & n5192 ;
  assign n5194 = ~\s4_msel_arb1_state_reg[1]/NET0131  & \s4_msel_arb1_state_reg[2]/NET0131  ;
  assign n5195 = ~\s4_msel_arb1_state_reg[0]/NET0131  & n5194 ;
  assign n5196 = ~\rf_conf4_reg[7]/NET0131  & n4043 ;
  assign n5197 = ~\s4_msel_arb1_state_reg[2]/NET0131  & ~n5196 ;
  assign n5198 = ~n5195 & ~n5197 ;
  assign n5199 = ~\rf_conf4_reg[1]/NET0131  & ~\s4_msel_arb1_state_reg[0]/NET0131  ;
  assign n5200 = n4040 & n5199 ;
  assign n5201 = ~\rf_conf4_reg[5]/NET0131  & n4045 ;
  assign n5202 = ~\rf_conf4_reg[3]/NET0131  & n4038 ;
  assign n5203 = ~n5201 & ~n5202 ;
  assign n5204 = ~n5200 & n5203 ;
  assign n5205 = ~\rf_conf4_reg[5]/NET0131  & ~\s4_msel_arb1_state_reg[0]/NET0131  ;
  assign n5206 = n4045 & n5205 ;
  assign n5207 = \s4_msel_arb1_state_reg[1]/NET0131  & ~n5206 ;
  assign n5208 = ~n5195 & ~n5207 ;
  assign n5209 = ~n5204 & n5208 ;
  assign n5210 = ~n5198 & ~n5209 ;
  assign n5211 = ~n5193 & n5210 ;
  assign n5212 = ~\rf_conf4_reg[1]/NET0131  & n4040 ;
  assign n5213 = ~n5202 & ~n5212 ;
  assign n5214 = ~n5196 & ~n5201 ;
  assign n5215 = n5213 & n5214 ;
  assign n5216 = \s4_msel_arb1_state_reg[1]/NET0131  & ~n5189 ;
  assign n5217 = ~\s4_msel_arb1_state_reg[0]/NET0131  & ~n5216 ;
  assign n5218 = ~n5187 & ~n5191 ;
  assign n5219 = \s4_msel_arb1_state_reg[0]/NET0131  & \s4_msel_arb1_state_reg[1]/NET0131  ;
  assign n5220 = ~n5218 & ~n5219 ;
  assign n5221 = ~n5188 & ~n5220 ;
  assign n5222 = ~n5217 & ~n5221 ;
  assign n5223 = ~n5215 & ~n5222 ;
  assign n5224 = \s4_msel_arb1_state_reg[2]/NET0131  & ~n5223 ;
  assign n5225 = ~n5211 & ~n5224 ;
  assign n5226 = ~\rf_conf5_reg[7]/NET0131  & n4627 ;
  assign n5227 = ~\rf_conf5_reg[5]/NET0131  & n4629 ;
  assign n5228 = ~n5226 & ~n5227 ;
  assign n5229 = ~\rf_conf5_reg[1]/NET0131  & n4634 ;
  assign n5230 = ~\rf_conf5_reg[3]/NET0131  & n4632 ;
  assign n5231 = ~n5229 & ~n5230 ;
  assign n5232 = \s5_msel_arb1_state_reg[2]/NET0131  & n5231 ;
  assign n5233 = n5228 & n5232 ;
  assign n5234 = ~\rf_conf5_reg[15]/NET0131  & n4622 ;
  assign n5235 = ~\rf_conf5_reg[13]/NET0131  & n4624 ;
  assign n5236 = ~n5234 & ~n5235 ;
  assign n5237 = ~\rf_conf5_reg[9]/NET0131  & n4612 ;
  assign n5238 = ~\rf_conf5_reg[11]/NET0131  & n4610 ;
  assign n5239 = ~n5237 & ~n5238 ;
  assign n5240 = n5236 & n5239 ;
  assign n5241 = ~\s5_msel_arb1_state_reg[1]/NET0131  & ~\s5_msel_arb1_state_reg[2]/NET0131  ;
  assign n5242 = ~n5230 & n5241 ;
  assign n5243 = n5228 & n5242 ;
  assign n5244 = ~n5240 & n5243 ;
  assign n5245 = ~n5233 & ~n5244 ;
  assign n5246 = \s5_msel_arb1_state_reg[2]/NET0131  & n5234 ;
  assign n5247 = ~n5235 & ~n5238 ;
  assign n5248 = ~\s5_msel_arb1_state_reg[1]/NET0131  & \s5_msel_arb1_state_reg[2]/NET0131  ;
  assign n5249 = ~n5247 & n5248 ;
  assign n5250 = ~n5246 & ~n5249 ;
  assign n5251 = n5245 & n5250 ;
  assign n5252 = \s5_msel_arb1_state_reg[0]/NET0131  & ~n5251 ;
  assign n5253 = ~\s5_msel_arb1_state_reg[2]/NET0131  & n5240 ;
  assign n5254 = \s5_msel_arb1_state_reg[1]/NET0131  & ~\s5_msel_arb1_state_reg[2]/NET0131  ;
  assign n5255 = ~\s5_msel_arb1_state_reg[0]/NET0131  & n5231 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = ~\rf_conf5_reg[5]/NET0131  & ~\s5_msel_arb1_state_reg[0]/NET0131  ;
  assign n5258 = n4629 & n5257 ;
  assign n5259 = ~n5226 & ~n5258 ;
  assign n5260 = ~n5256 & n5259 ;
  assign n5261 = ~n5253 & n5260 ;
  assign n5262 = ~\s5_msel_arb1_state_reg[0]/NET0131  & \s5_msel_arb1_state_reg[2]/NET0131  ;
  assign n5263 = ~n5236 & n5262 ;
  assign n5264 = ~\s5_msel_arb1_state_reg[1]/NET0131  & n5262 ;
  assign n5265 = ~n5239 & n5264 ;
  assign n5266 = ~n5263 & ~n5265 ;
  assign n5267 = ~n5261 & n5266 ;
  assign n5268 = ~n5252 & n5267 ;
  assign n5269 = ~\rf_conf6_reg[7]/NET0131  & n4681 ;
  assign n5270 = ~\rf_conf6_reg[5]/NET0131  & n4683 ;
  assign n5271 = ~n5269 & ~n5270 ;
  assign n5272 = ~\rf_conf6_reg[1]/NET0131  & n4688 ;
  assign n5273 = ~\rf_conf6_reg[3]/NET0131  & n4686 ;
  assign n5274 = ~n5272 & ~n5273 ;
  assign n5275 = \s6_msel_arb1_state_reg[2]/NET0131  & n5274 ;
  assign n5276 = n5271 & n5275 ;
  assign n5277 = ~\rf_conf6_reg[15]/NET0131  & n4676 ;
  assign n5278 = ~\rf_conf6_reg[13]/NET0131  & n4678 ;
  assign n5279 = ~n5277 & ~n5278 ;
  assign n5280 = ~\rf_conf6_reg[9]/NET0131  & n4666 ;
  assign n5281 = ~\rf_conf6_reg[11]/NET0131  & n4664 ;
  assign n5282 = ~n5280 & ~n5281 ;
  assign n5283 = n5279 & n5282 ;
  assign n5284 = ~\s6_msel_arb1_state_reg[1]/NET0131  & ~\s6_msel_arb1_state_reg[2]/NET0131  ;
  assign n5285 = ~n5273 & n5284 ;
  assign n5286 = n5271 & n5285 ;
  assign n5287 = ~n5283 & n5286 ;
  assign n5288 = ~n5276 & ~n5287 ;
  assign n5289 = \s6_msel_arb1_state_reg[2]/NET0131  & n5277 ;
  assign n5290 = ~n5278 & ~n5281 ;
  assign n5291 = ~\s6_msel_arb1_state_reg[1]/NET0131  & \s6_msel_arb1_state_reg[2]/NET0131  ;
  assign n5292 = ~n5290 & n5291 ;
  assign n5293 = ~n5289 & ~n5292 ;
  assign n5294 = n5288 & n5293 ;
  assign n5295 = \s6_msel_arb1_state_reg[0]/NET0131  & ~n5294 ;
  assign n5296 = ~\s6_msel_arb1_state_reg[2]/NET0131  & n5283 ;
  assign n5297 = \s6_msel_arb1_state_reg[1]/NET0131  & ~\s6_msel_arb1_state_reg[2]/NET0131  ;
  assign n5298 = ~\s6_msel_arb1_state_reg[0]/NET0131  & n5274 ;
  assign n5299 = ~n5297 & ~n5298 ;
  assign n5300 = ~\rf_conf6_reg[5]/NET0131  & ~\s6_msel_arb1_state_reg[0]/NET0131  ;
  assign n5301 = n4683 & n5300 ;
  assign n5302 = ~n5269 & ~n5301 ;
  assign n5303 = ~n5299 & n5302 ;
  assign n5304 = ~n5296 & n5303 ;
  assign n5305 = ~\s6_msel_arb1_state_reg[0]/NET0131  & \s6_msel_arb1_state_reg[2]/NET0131  ;
  assign n5306 = ~n5279 & n5305 ;
  assign n5307 = ~\s6_msel_arb1_state_reg[1]/NET0131  & n5305 ;
  assign n5308 = ~n5282 & n5307 ;
  assign n5309 = ~n5306 & ~n5308 ;
  assign n5310 = ~n5304 & n5309 ;
  assign n5311 = ~n5295 & n5310 ;
  assign n5312 = ~\rf_conf7_reg[3]/NET0131  & n4740 ;
  assign n5313 = ~\rf_conf7_reg[1]/NET0131  & n4742 ;
  assign n5314 = ~n5312 & ~n5313 ;
  assign n5315 = ~\rf_conf7_reg[7]/NET0131  & n4735 ;
  assign n5316 = ~\rf_conf7_reg[5]/NET0131  & n4737 ;
  assign n5317 = ~n5315 & ~n5316 ;
  assign n5318 = n5314 & n5317 ;
  assign n5319 = ~\rf_conf7_reg[11]/NET0131  & n4718 ;
  assign n5320 = ~\rf_conf7_reg[9]/NET0131  & n4720 ;
  assign n5321 = ~n5319 & ~n5320 ;
  assign n5322 = ~\rf_conf7_reg[15]/NET0131  & n4730 ;
  assign n5323 = ~\rf_conf7_reg[13]/NET0131  & n4732 ;
  assign n5324 = ~n5322 & ~n5323 ;
  assign n5325 = n5321 & n5324 ;
  assign n5326 = ~\s7_msel_arb1_state_reg[0]/NET0131  & ~\s7_msel_arb1_state_reg[1]/NET0131  ;
  assign n5327 = n5325 & n5326 ;
  assign n5328 = ~n5318 & n5327 ;
  assign n5329 = ~\rf_conf7_reg[13]/NET0131  & ~\s7_msel_arb1_state_reg[0]/NET0131  ;
  assign n5330 = n4732 & n5329 ;
  assign n5331 = \s7_msel_arb1_state_reg[1]/NET0131  & ~n5330 ;
  assign n5332 = \s7_msel_arb1_state_reg[0]/NET0131  & ~n5323 ;
  assign n5333 = ~n5319 & n5332 ;
  assign n5334 = ~n5331 & ~n5333 ;
  assign n5335 = \s7_msel_arb1_state_reg[2]/NET0131  & ~n5322 ;
  assign n5336 = ~n5318 & n5335 ;
  assign n5337 = ~n5334 & n5336 ;
  assign n5338 = ~n5328 & ~n5337 ;
  assign n5339 = ~\rf_conf7_reg[1]/NET0131  & ~\s7_msel_arb1_state_reg[0]/NET0131  ;
  assign n5340 = n4742 & n5339 ;
  assign n5341 = ~n5312 & ~n5340 ;
  assign n5342 = ~\s7_msel_arb1_state_reg[1]/NET0131  & ~n5341 ;
  assign n5343 = \s7_msel_arb1_state_reg[0]/NET0131  & \s7_msel_arb1_state_reg[1]/NET0131  ;
  assign n5344 = n5316 & ~n5343 ;
  assign n5345 = ~n5315 & ~n5344 ;
  assign n5346 = ~n5325 & n5345 ;
  assign n5347 = ~n5342 & n5346 ;
  assign n5348 = ~\s7_msel_arb1_state_reg[2]/NET0131  & ~n5347 ;
  assign n5349 = n5338 & ~n5348 ;
  assign n5350 = ~\rf_conf8_reg[7]/NET0131  & n4778 ;
  assign n5351 = ~\rf_conf8_reg[5]/NET0131  & n4780 ;
  assign n5352 = ~n5350 & ~n5351 ;
  assign n5353 = ~\rf_conf8_reg[1]/NET0131  & n4775 ;
  assign n5354 = ~\rf_conf8_reg[3]/NET0131  & n4773 ;
  assign n5355 = ~n5353 & ~n5354 ;
  assign n5356 = \s8_msel_arb1_state_reg[2]/NET0131  & n5355 ;
  assign n5357 = n5352 & n5356 ;
  assign n5358 = ~\rf_conf8_reg[15]/NET0131  & n4786 ;
  assign n5359 = ~\rf_conf8_reg[13]/NET0131  & n4788 ;
  assign n5360 = ~n5358 & ~n5359 ;
  assign n5361 = ~\rf_conf8_reg[9]/NET0131  & n4797 ;
  assign n5362 = ~\rf_conf8_reg[11]/NET0131  & n4784 ;
  assign n5363 = ~n5361 & ~n5362 ;
  assign n5364 = n5360 & n5363 ;
  assign n5365 = ~\s8_msel_arb1_state_reg[1]/NET0131  & ~\s8_msel_arb1_state_reg[2]/NET0131  ;
  assign n5366 = ~n5354 & n5365 ;
  assign n5367 = n5352 & n5366 ;
  assign n5368 = ~n5364 & n5367 ;
  assign n5369 = ~n5357 & ~n5368 ;
  assign n5370 = \s8_msel_arb1_state_reg[2]/NET0131  & n5358 ;
  assign n5371 = ~n5359 & ~n5362 ;
  assign n5372 = ~\s8_msel_arb1_state_reg[1]/NET0131  & \s8_msel_arb1_state_reg[2]/NET0131  ;
  assign n5373 = ~n5371 & n5372 ;
  assign n5374 = ~n5370 & ~n5373 ;
  assign n5375 = n5369 & n5374 ;
  assign n5376 = \s8_msel_arb1_state_reg[0]/NET0131  & ~n5375 ;
  assign n5377 = ~\s8_msel_arb1_state_reg[2]/NET0131  & n5364 ;
  assign n5378 = \s8_msel_arb1_state_reg[1]/NET0131  & ~\s8_msel_arb1_state_reg[2]/NET0131  ;
  assign n5379 = ~\s8_msel_arb1_state_reg[0]/NET0131  & n5355 ;
  assign n5380 = ~n5378 & ~n5379 ;
  assign n5381 = ~\rf_conf8_reg[5]/NET0131  & ~\s8_msel_arb1_state_reg[0]/NET0131  ;
  assign n5382 = n4780 & n5381 ;
  assign n5383 = ~n5350 & ~n5382 ;
  assign n5384 = ~n5380 & n5383 ;
  assign n5385 = ~n5377 & n5384 ;
  assign n5386 = ~\s8_msel_arb1_state_reg[0]/NET0131  & \s8_msel_arb1_state_reg[2]/NET0131  ;
  assign n5387 = ~n5360 & n5386 ;
  assign n5388 = ~\s8_msel_arb1_state_reg[1]/NET0131  & n5386 ;
  assign n5389 = ~n5363 & n5388 ;
  assign n5390 = ~n5387 & ~n5389 ;
  assign n5391 = ~n5385 & n5390 ;
  assign n5392 = ~n5376 & n5391 ;
  assign n5393 = \m3_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[6]/NET0131  ;
  assign n5394 = ~\rf_conf9_reg[7]/NET0131  & n5393 ;
  assign n5395 = \m2_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[4]/NET0131  ;
  assign n5396 = ~\rf_conf9_reg[5]/NET0131  & n5395 ;
  assign n5397 = ~n5394 & ~n5396 ;
  assign n5398 = \m0_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[0]/NET0131  ;
  assign n5399 = ~\rf_conf9_reg[1]/NET0131  & n5398 ;
  assign n5400 = \m1_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[2]/NET0131  ;
  assign n5401 = ~\rf_conf9_reg[3]/NET0131  & n5400 ;
  assign n5402 = ~n5399 & ~n5401 ;
  assign n5403 = \s9_msel_arb1_state_reg[2]/NET0131  & n5402 ;
  assign n5404 = n5397 & n5403 ;
  assign n5405 = \m7_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[14]/NET0131  ;
  assign n5406 = ~\rf_conf9_reg[15]/NET0131  & n5405 ;
  assign n5407 = \m6_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[12]/NET0131  ;
  assign n5408 = ~\rf_conf9_reg[13]/NET0131  & n5407 ;
  assign n5409 = ~n5406 & ~n5408 ;
  assign n5410 = \m4_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[8]/NET0131  ;
  assign n5411 = ~\rf_conf9_reg[9]/NET0131  & n5410 ;
  assign n5412 = \m5_s9_cyc_o_reg/NET0131  & \rf_conf9_reg[10]/NET0131  ;
  assign n5413 = ~\rf_conf9_reg[11]/NET0131  & n5412 ;
  assign n5414 = ~n5411 & ~n5413 ;
  assign n5415 = n5409 & n5414 ;
  assign n5416 = ~\s9_msel_arb1_state_reg[1]/NET0131  & ~\s9_msel_arb1_state_reg[2]/NET0131  ;
  assign n5417 = ~n5401 & n5416 ;
  assign n5418 = n5397 & n5417 ;
  assign n5419 = ~n5415 & n5418 ;
  assign n5420 = ~n5404 & ~n5419 ;
  assign n5421 = \s9_msel_arb1_state_reg[2]/NET0131  & n5406 ;
  assign n5422 = ~n5408 & ~n5413 ;
  assign n5423 = ~\s9_msel_arb1_state_reg[1]/NET0131  & \s9_msel_arb1_state_reg[2]/NET0131  ;
  assign n5424 = ~n5422 & n5423 ;
  assign n5425 = ~n5421 & ~n5424 ;
  assign n5426 = n5420 & n5425 ;
  assign n5427 = \s9_msel_arb1_state_reg[0]/NET0131  & ~n5426 ;
  assign n5428 = ~\s9_msel_arb1_state_reg[2]/NET0131  & n5415 ;
  assign n5429 = \s9_msel_arb1_state_reg[1]/NET0131  & ~\s9_msel_arb1_state_reg[2]/NET0131  ;
  assign n5430 = ~\s9_msel_arb1_state_reg[0]/NET0131  & n5402 ;
  assign n5431 = ~n5429 & ~n5430 ;
  assign n5432 = ~\rf_conf9_reg[5]/NET0131  & ~\s9_msel_arb1_state_reg[0]/NET0131  ;
  assign n5433 = n5395 & n5432 ;
  assign n5434 = ~n5394 & ~n5433 ;
  assign n5435 = ~n5431 & n5434 ;
  assign n5436 = ~n5428 & n5435 ;
  assign n5437 = ~\s9_msel_arb1_state_reg[0]/NET0131  & \s9_msel_arb1_state_reg[2]/NET0131  ;
  assign n5438 = ~n5409 & n5437 ;
  assign n5439 = ~\s9_msel_arb1_state_reg[1]/NET0131  & n5437 ;
  assign n5440 = ~n5414 & n5439 ;
  assign n5441 = ~n5438 & ~n5440 ;
  assign n5442 = ~n5436 & n5441 ;
  assign n5443 = ~n5427 & n5442 ;
  assign n5444 = ~\rf_conf0_reg[7]/NET0131  & n4840 ;
  assign n5445 = ~\rf_conf0_reg[5]/NET0131  & n4842 ;
  assign n5446 = ~n5444 & ~n5445 ;
  assign n5447 = ~\rf_conf0_reg[1]/NET0131  & n4847 ;
  assign n5448 = ~\rf_conf0_reg[3]/NET0131  & n4845 ;
  assign n5449 = ~n5447 & ~n5448 ;
  assign n5450 = \s0_msel_arb1_state_reg[2]/NET0131  & n5449 ;
  assign n5451 = n5446 & n5450 ;
  assign n5452 = ~\rf_conf0_reg[15]/NET0131  & n4835 ;
  assign n5453 = ~\rf_conf0_reg[13]/NET0131  & n4837 ;
  assign n5454 = ~n5452 & ~n5453 ;
  assign n5455 = ~\rf_conf0_reg[9]/NET0131  & n4825 ;
  assign n5456 = ~\rf_conf0_reg[11]/NET0131  & n4823 ;
  assign n5457 = ~n5455 & ~n5456 ;
  assign n5458 = n5454 & n5457 ;
  assign n5459 = ~\s0_msel_arb1_state_reg[1]/NET0131  & ~\s0_msel_arb1_state_reg[2]/NET0131  ;
  assign n5460 = ~n5448 & n5459 ;
  assign n5461 = n5446 & n5460 ;
  assign n5462 = ~n5458 & n5461 ;
  assign n5463 = ~n5451 & ~n5462 ;
  assign n5464 = \s0_msel_arb1_state_reg[2]/NET0131  & n5452 ;
  assign n5465 = ~n5453 & ~n5456 ;
  assign n5466 = ~\s0_msel_arb1_state_reg[1]/NET0131  & \s0_msel_arb1_state_reg[2]/NET0131  ;
  assign n5467 = ~n5465 & n5466 ;
  assign n5468 = ~n5464 & ~n5467 ;
  assign n5469 = n5463 & n5468 ;
  assign n5470 = \s0_msel_arb1_state_reg[0]/NET0131  & ~n5469 ;
  assign n5471 = ~\s0_msel_arb1_state_reg[2]/NET0131  & n5458 ;
  assign n5472 = \s0_msel_arb1_state_reg[1]/NET0131  & ~\s0_msel_arb1_state_reg[2]/NET0131  ;
  assign n5473 = ~\s0_msel_arb1_state_reg[0]/NET0131  & n5449 ;
  assign n5474 = ~n5472 & ~n5473 ;
  assign n5475 = ~\rf_conf0_reg[5]/NET0131  & ~\s0_msel_arb1_state_reg[0]/NET0131  ;
  assign n5476 = n4842 & n5475 ;
  assign n5477 = ~n5444 & ~n5476 ;
  assign n5478 = ~n5474 & n5477 ;
  assign n5479 = ~n5471 & n5478 ;
  assign n5480 = ~\s0_msel_arb1_state_reg[0]/NET0131  & \s0_msel_arb1_state_reg[2]/NET0131  ;
  assign n5481 = ~n5454 & n5480 ;
  assign n5482 = ~\s0_msel_arb1_state_reg[1]/NET0131  & n5480 ;
  assign n5483 = ~n5457 & n5482 ;
  assign n5484 = ~n5481 & ~n5483 ;
  assign n5485 = ~n5479 & n5484 ;
  assign n5486 = ~n5470 & n5485 ;
  assign n5487 = ~n4877 & ~n4890 ;
  assign n5488 = ~n4877 & n4891 ;
  assign n5489 = ~n4879 & ~n5488 ;
  assign n5490 = ~n5487 & n5489 ;
  assign n5491 = ~n4879 & ~n4891 ;
  assign n5492 = n4886 & ~n4887 ;
  assign n5493 = n5491 & n5492 ;
  assign n5494 = ~n4884 & ~n5493 ;
  assign n5495 = ~n5490 & n5494 ;
  assign n5496 = \s10_msel_arb1_state_reg[1]/NET0131  & ~\s10_msel_arb1_state_reg[2]/NET0131  ;
  assign n5497 = ~n4883 & n5496 ;
  assign n5498 = ~n5495 & n5497 ;
  assign n5499 = ~\s10_msel_arb1_state_reg[0]/NET0131  & n5498 ;
  assign n5500 = n4877 & ~n4879 ;
  assign n5501 = ~n5491 & ~n5500 ;
  assign n5502 = n4887 & ~n4890 ;
  assign n5503 = ~n4883 & n4884 ;
  assign n5504 = ~n4886 & ~n4890 ;
  assign n5505 = ~n5503 & n5504 ;
  assign n5506 = ~n5502 & ~n5505 ;
  assign n5507 = \s10_msel_arb1_state_reg[0]/NET0131  & ~n4887 ;
  assign n5508 = ~n4883 & n5507 ;
  assign n5509 = ~n5500 & ~n5508 ;
  assign n5510 = ~n5506 & n5509 ;
  assign n5511 = ~n5501 & ~n5510 ;
  assign n5512 = ~\s10_msel_arb1_state_reg[1]/NET0131  & \s10_msel_arb1_state_reg[2]/NET0131  ;
  assign n5513 = ~\s10_msel_arb1_state_reg[0]/NET0131  & n5512 ;
  assign n5514 = n5511 & n5513 ;
  assign n5515 = ~n5499 & ~n5514 ;
  assign n5516 = ~n4884 & ~n5490 ;
  assign n5517 = ~n5492 & ~n5508 ;
  assign n5518 = n5491 & ~n5517 ;
  assign n5519 = n5516 & ~n5518 ;
  assign n5520 = n5496 & ~n5519 ;
  assign n5521 = ~\s10_msel_arb1_state_reg[1]/NET0131  & ~\s10_msel_arb1_state_reg[2]/NET0131  ;
  assign n5522 = ~n4886 & ~n5503 ;
  assign n5523 = ~n4883 & n5500 ;
  assign n5524 = n5522 & ~n5523 ;
  assign n5525 = ~n4883 & n5491 ;
  assign n5526 = ~n4890 & ~n5507 ;
  assign n5527 = n5525 & ~n5526 ;
  assign n5528 = n5524 & ~n5527 ;
  assign n5529 = n5521 & ~n5528 ;
  assign n5530 = ~n4879 & ~n4883 ;
  assign n5531 = n5507 & n5530 ;
  assign n5532 = ~n4877 & ~n5531 ;
  assign n5533 = ~n5506 & n5532 ;
  assign n5534 = ~n5488 & n5512 ;
  assign n5535 = ~n5533 & n5534 ;
  assign n5536 = ~n5529 & ~n5535 ;
  assign n5537 = ~n5520 & n5536 ;
  assign n5538 = \s10_msel_arb1_state_reg[0]/NET0131  & ~n5537 ;
  assign n5539 = ~\rf_conf10_reg[13]/NET0131  & ~\s10_msel_arb1_state_reg[0]/NET0131  ;
  assign n5540 = n4207 & n5539 ;
  assign n5541 = \s10_msel_arb1_state_reg[1]/NET0131  & \s10_msel_arb1_state_reg[2]/NET0131  ;
  assign n5542 = ~n5540 & n5541 ;
  assign n5543 = n4890 & n5542 ;
  assign n5544 = \s10_msel_arb1_state_reg[0]/NET0131  & ~n4883 ;
  assign n5545 = n5491 & n5544 ;
  assign n5546 = n5524 & ~n5545 ;
  assign n5547 = n5542 & ~n5546 ;
  assign n5548 = ~n4887 & n5547 ;
  assign n5549 = ~n4883 & ~n5487 ;
  assign n5550 = n5489 & n5549 ;
  assign n5551 = ~n5503 & ~n5550 ;
  assign n5552 = ~n4886 & n5551 ;
  assign n5553 = ~\s10_msel_arb1_state_reg[0]/NET0131  & n5521 ;
  assign n5554 = ~n4887 & n5553 ;
  assign n5555 = ~n5552 & n5554 ;
  assign n5556 = ~n5548 & ~n5555 ;
  assign n5557 = ~n5543 & n5556 ;
  assign n5558 = ~n5538 & n5557 ;
  assign n5559 = n5515 & n5558 ;
  assign n5560 = \rf_conf10_reg[5]/NET0131  & n3686 ;
  assign n5561 = \rf_conf10_reg[7]/NET0131  & n3684 ;
  assign n5562 = ~n5560 & n5561 ;
  assign n5563 = \s10_msel_arb2_state_reg[1]/NET0131  & ~\s10_msel_arb2_state_reg[2]/NET0131  ;
  assign n5564 = n5562 & n5563 ;
  assign n5565 = \rf_conf10_reg[11]/NET0131  & n3691 ;
  assign n5566 = \rf_conf10_reg[15]/NET0131  & n3694 ;
  assign n5567 = \rf_conf10_reg[13]/NET0131  & n3696 ;
  assign n5568 = n5566 & ~n5567 ;
  assign n5569 = ~n5565 & ~n5568 ;
  assign n5570 = \rf_conf10_reg[3]/NET0131  & n3701 ;
  assign n5571 = \rf_conf10_reg[1]/NET0131  & n3703 ;
  assign n5572 = ~n5567 & ~n5571 ;
  assign n5573 = n5570 & n5572 ;
  assign n5574 = n5569 & ~n5573 ;
  assign n5575 = \rf_conf10_reg[9]/NET0131  & n3689 ;
  assign n5576 = ~n5560 & ~n5575 ;
  assign n5577 = n5563 & n5576 ;
  assign n5578 = ~n5574 & n5577 ;
  assign n5579 = ~n5564 & ~n5578 ;
  assign n5580 = ~n5562 & ~n5570 ;
  assign n5581 = ~\s10_msel_arb2_state_reg[1]/NET0131  & ~\s10_msel_arb2_state_reg[2]/NET0131  ;
  assign n5582 = ~n5571 & n5581 ;
  assign n5583 = ~n5580 & n5582 ;
  assign n5584 = n5576 & n5582 ;
  assign n5585 = ~n5569 & n5584 ;
  assign n5586 = ~n5583 & ~n5585 ;
  assign n5587 = ~\s10_msel_arb2_state_reg[0]/NET0131  & n5586 ;
  assign n5588 = n5579 & n5587 ;
  assign n5589 = \s10_msel_arb2_state_reg[1]/NET0131  & \s10_msel_arb2_state_reg[2]/NET0131  ;
  assign n5590 = n5568 & n5589 ;
  assign n5591 = n5565 & n5576 ;
  assign n5592 = n5580 & ~n5591 ;
  assign n5593 = n5572 & n5589 ;
  assign n5594 = ~n5592 & n5593 ;
  assign n5595 = ~n5590 & ~n5594 ;
  assign n5596 = ~\s10_msel_arb2_state_reg[1]/NET0131  & \s10_msel_arb2_state_reg[2]/NET0131  ;
  assign n5597 = ~n5575 & n5596 ;
  assign n5598 = n5565 & n5597 ;
  assign n5599 = ~n5566 & n5571 ;
  assign n5600 = ~n5566 & ~n5570 ;
  assign n5601 = ~n5562 & n5600 ;
  assign n5602 = ~n5599 & ~n5601 ;
  assign n5603 = ~n5567 & n5597 ;
  assign n5604 = n5602 & n5603 ;
  assign n5605 = ~n5598 & ~n5604 ;
  assign n5606 = n5595 & n5605 ;
  assign n5607 = n5588 & n5606 ;
  assign n5608 = \s10_msel_arb2_state_reg[0]/NET0131  & ~n5571 ;
  assign n5609 = n5576 & n5608 ;
  assign n5610 = ~n5602 & ~n5609 ;
  assign n5611 = \s10_msel_arb2_state_reg[0]/NET0131  & n5596 ;
  assign n5612 = ~n5565 & n5611 ;
  assign n5613 = ~n5567 & n5612 ;
  assign n5614 = ~n5610 & n5613 ;
  assign n5615 = n5607 & ~n5614 ;
  assign n5616 = ~n5569 & n5576 ;
  assign n5617 = n5580 & ~n5616 ;
  assign n5618 = \s10_msel_arb2_state_reg[0]/NET0131  & n5576 ;
  assign n5619 = n5572 & n5618 ;
  assign n5620 = n5617 & ~n5619 ;
  assign n5621 = n5581 & ~n5620 ;
  assign n5622 = n5561 & n5563 ;
  assign n5623 = n5560 & ~n5570 ;
  assign n5624 = n5572 & ~n5623 ;
  assign n5625 = n5569 & ~n5624 ;
  assign n5626 = n5563 & ~n5575 ;
  assign n5627 = ~n5625 & n5626 ;
  assign n5628 = ~n5622 & ~n5627 ;
  assign n5629 = n5565 & n5596 ;
  assign n5630 = \s10_msel_arb2_state_reg[0]/NET0131  & ~n5629 ;
  assign n5631 = n5628 & n5630 ;
  assign n5632 = ~n5621 & n5631 ;
  assign n5633 = \s10_msel_arb2_state_reg[0]/NET0131  & ~n5567 ;
  assign n5634 = n5576 & n5633 ;
  assign n5635 = ~n5566 & ~n5634 ;
  assign n5636 = n5592 & n5635 ;
  assign n5637 = ~n5599 & ~n5636 ;
  assign n5638 = n5589 & n5637 ;
  assign n5639 = ~n5614 & ~n5638 ;
  assign n5640 = n5632 & n5639 ;
  assign n5641 = ~n5615 & ~n5640 ;
  assign n5642 = \s10_msel_arb3_state_reg[1]/NET0131  & ~\s10_msel_arb3_state_reg[2]/NET0131  ;
  assign n5643 = ~n4227 & n5642 ;
  assign n5644 = ~n4194 & ~n4206 ;
  assign n5645 = ~n4194 & n4208 ;
  assign n5646 = ~n5644 & ~n5645 ;
  assign n5647 = n5643 & n5646 ;
  assign n5648 = ~n4216 & ~n4234 ;
  assign n5649 = ~n4208 & ~n4218 ;
  assign n5650 = n5643 & n5649 ;
  assign n5651 = ~n5648 & n5650 ;
  assign n5652 = ~n5647 & ~n5651 ;
  assign n5653 = ~n4196 & ~n5652 ;
  assign n5654 = n4211 & ~n4213 ;
  assign n5655 = ~n4216 & ~n5654 ;
  assign n5656 = ~n4218 & ~n5655 ;
  assign n5657 = n5644 & ~n5656 ;
  assign n5658 = ~\s10_msel_arb3_state_reg[0]/NET0131  & \s10_msel_arb3_state_reg[2]/NET0131  ;
  assign n5659 = ~\s10_msel_arb3_state_reg[1]/NET0131  & n5658 ;
  assign n5660 = ~n5645 & n5659 ;
  assign n5661 = ~n4196 & n5660 ;
  assign n5662 = ~n5657 & n5661 ;
  assign n5663 = ~n5653 & ~n5662 ;
  assign n5664 = ~\s10_msel_arb3_state_reg[1]/NET0131  & ~\s10_msel_arb3_state_reg[2]/NET0131  ;
  assign n5665 = \rf_conf10_reg[1]/NET0131  & ~\s10_msel_arb3_state_reg[0]/NET0131  ;
  assign n5666 = n4217 & n5665 ;
  assign n5667 = n5664 & ~n5666 ;
  assign n5668 = ~n5655 & n5667 ;
  assign n5669 = ~n4196 & ~n4213 ;
  assign n5670 = n5667 & n5669 ;
  assign n5671 = n5646 & n5670 ;
  assign n5672 = ~n5668 & ~n5671 ;
  assign n5673 = n4211 & n5643 ;
  assign n5674 = ~\s10_msel_arb3_state_reg[1]/NET0131  & n4199 ;
  assign n5675 = n4194 & n5674 ;
  assign n5676 = ~n5673 & ~n5675 ;
  assign n5677 = n5672 & n5676 ;
  assign n5678 = n5663 & n5677 ;
  assign n5679 = \s10_msel_arb3_state_reg[0]/NET0131  & n5664 ;
  assign n5680 = ~n4218 & n5679 ;
  assign n5681 = n5669 & n5680 ;
  assign n5682 = ~n4194 & n5674 ;
  assign n5683 = ~n5681 & ~n5682 ;
  assign n5684 = ~n4206 & n4218 ;
  assign n5685 = ~n4206 & ~n4216 ;
  assign n5686 = ~n5654 & n5685 ;
  assign n5687 = ~n5684 & ~n5686 ;
  assign n5688 = \s10_msel_arb3_state_reg[0]/NET0131  & ~n4218 ;
  assign n5689 = n5669 & n5688 ;
  assign n5690 = ~n5681 & ~n5689 ;
  assign n5691 = ~n5687 & n5690 ;
  assign n5692 = ~n5683 & ~n5691 ;
  assign n5693 = ~n4208 & n5692 ;
  assign n5694 = ~n4218 & n5669 ;
  assign n5695 = ~\s10_msel_arb3_state_reg[0]/NET0131  & ~n4194 ;
  assign n5696 = n5694 & ~n5695 ;
  assign n5697 = ~n5687 & ~n5696 ;
  assign n5698 = ~\s10_msel_arb3_state_reg[0]/NET0131  & n4208 ;
  assign n5699 = n4208 & n5644 ;
  assign n5700 = n5655 & n5699 ;
  assign n5701 = ~n5698 & ~n5700 ;
  assign n5702 = n4241 & n5701 ;
  assign n5703 = ~n5697 & n5702 ;
  assign n5704 = ~n5693 & ~n5703 ;
  assign n5705 = n5678 & n5704 ;
  assign n5706 = ~n2751 & n2764 ;
  assign n5707 = n2746 & ~n2748 ;
  assign n5708 = ~n2743 & n5707 ;
  assign n5709 = ~n2748 & ~n2753 ;
  assign n5710 = \s11_msel_arb0_state_reg[0]/NET0131  & ~n2743 ;
  assign n5711 = n5709 & n5710 ;
  assign n5712 = ~n5708 & ~n5711 ;
  assign n5713 = n2743 & ~n2758 ;
  assign n5714 = ~n2741 & ~n2758 ;
  assign n5715 = ~n5713 & ~n5714 ;
  assign n5716 = ~n2751 & ~n5715 ;
  assign n5717 = n5712 & n5716 ;
  assign n5718 = ~n5706 & ~n5717 ;
  assign n5719 = n2787 & n5718 ;
  assign n5720 = \s11_msel_arb0_state_reg[1]/NET0131  & \s11_msel_arb0_state_reg[2]/NET0131  ;
  assign n5721 = n2758 & ~n2764 ;
  assign n5722 = ~n2751 & ~n5721 ;
  assign n5723 = ~n2753 & ~n5722 ;
  assign n5724 = ~n2743 & ~n2764 ;
  assign n5725 = ~\s11_msel_arb0_state_reg[0]/NET0131  & ~n2741 ;
  assign n5726 = n5724 & ~n5725 ;
  assign n5727 = ~n2741 & n2748 ;
  assign n5728 = ~n2753 & ~n5727 ;
  assign n5729 = n5726 & n5728 ;
  assign n5730 = ~n5723 & ~n5729 ;
  assign n5731 = ~n2746 & n5730 ;
  assign n5732 = n5720 & ~n5731 ;
  assign n5733 = n2751 & ~n2753 ;
  assign n5734 = ~n2741 & ~n2746 ;
  assign n5735 = ~n5733 & n5734 ;
  assign n5736 = ~n5727 & ~n5735 ;
  assign n5737 = \s11_msel_arb0_state_reg[0]/NET0131  & ~n2764 ;
  assign n5738 = n5709 & n5737 ;
  assign n5739 = ~n2758 & ~n5738 ;
  assign n5740 = ~n5736 & n5739 ;
  assign n5741 = \s11_msel_arb0_state_reg[1]/NET0131  & ~\s11_msel_arb0_state_reg[2]/NET0131  ;
  assign n5742 = ~n5713 & n5741 ;
  assign n5743 = ~n5740 & n5742 ;
  assign n5744 = ~n5732 & ~n5743 ;
  assign n5745 = ~n5719 & n5744 ;
  assign n5746 = \s11_msel_arb0_state_reg[0]/NET0131  & ~n5745 ;
  assign n5747 = \s11_msel_arb0_state_reg[0]/NET0131  & n5709 ;
  assign n5748 = n5724 & n5747 ;
  assign n5749 = n5724 & ~n5727 ;
  assign n5750 = ~n5735 & n5749 ;
  assign n5751 = ~n5748 & ~n5750 ;
  assign n5752 = ~n5721 & n5751 ;
  assign n5753 = n5741 & ~n5752 ;
  assign n5754 = n5707 & n5720 ;
  assign n5755 = n5722 & ~n5726 ;
  assign n5756 = n5709 & n5720 ;
  assign n5757 = ~n5755 & n5756 ;
  assign n5758 = ~n5754 & ~n5757 ;
  assign n5759 = n2787 & n5733 ;
  assign n5760 = ~n2743 & ~n2748 ;
  assign n5761 = ~\s11_msel_arb0_state_reg[0]/NET0131  & ~n2746 ;
  assign n5762 = n5760 & ~n5761 ;
  assign n5763 = ~n5715 & ~n5762 ;
  assign n5764 = ~n2753 & ~n2764 ;
  assign n5765 = n2787 & n5764 ;
  assign n5766 = ~n5763 & n5765 ;
  assign n5767 = ~n5759 & ~n5766 ;
  assign n5768 = n5758 & n5767 ;
  assign n5769 = ~n5753 & n5768 ;
  assign n5770 = ~\s11_msel_arb0_state_reg[0]/NET0131  & ~n5769 ;
  assign n5771 = \s11_msel_arb0_state_reg[0]/NET0131  & n5764 ;
  assign n5772 = n5760 & n5771 ;
  assign n5773 = n2791 & n5772 ;
  assign n5774 = n2758 & n5764 ;
  assign n5775 = n5735 & ~n5774 ;
  assign n5776 = ~\rf_conf11_reg[9]/NET0131  & ~\s11_msel_arb0_state_reg[0]/NET0131  ;
  assign n5777 = n2742 & n5776 ;
  assign n5778 = ~n5727 & ~n5777 ;
  assign n5779 = n2791 & n5778 ;
  assign n5780 = ~n5775 & n5779 ;
  assign n5781 = ~n5773 & ~n5780 ;
  assign n5782 = ~n5770 & n5781 ;
  assign n5783 = ~n5746 & n5782 ;
  assign n5784 = ~\rf_conf11_reg[9]/NET0131  & ~\s11_msel_arb1_state_reg[0]/NET0131  ;
  assign n5785 = n4307 & n5784 ;
  assign n5786 = n4946 & ~n5785 ;
  assign n5787 = ~n4914 & n4923 ;
  assign n5788 = n4911 & ~n4933 ;
  assign n5789 = ~n4914 & ~n4934 ;
  assign n5790 = ~n5788 & n5789 ;
  assign n5791 = ~n5787 & ~n5790 ;
  assign n5792 = ~n4915 & n5791 ;
  assign n5793 = ~n4915 & ~n4923 ;
  assign n5794 = ~n4917 & ~n4933 ;
  assign n5795 = \s11_msel_arb1_state_reg[0]/NET0131  & n5794 ;
  assign n5796 = n5793 & n5795 ;
  assign n5797 = ~n4918 & ~n5796 ;
  assign n5798 = ~n5792 & n5797 ;
  assign n5799 = n5786 & ~n5798 ;
  assign n5800 = ~\s11_msel_arb1_state_reg[0]/NET0131  & n4912 ;
  assign n5801 = n5788 & n5800 ;
  assign n5802 = n4914 & ~n4915 ;
  assign n5803 = ~n4918 & ~n5802 ;
  assign n5804 = ~\s11_msel_arb1_state_reg[0]/NET0131  & ~n4934 ;
  assign n5805 = n5793 & ~n5804 ;
  assign n5806 = n5803 & ~n5805 ;
  assign n5807 = n5794 & n5800 ;
  assign n5808 = ~n5806 & n5807 ;
  assign n5809 = ~n5801 & ~n5808 ;
  assign n5810 = n4918 & ~n4923 ;
  assign n5811 = n5794 & n5810 ;
  assign n5812 = ~n5796 & ~n5811 ;
  assign n5813 = ~n5791 & n5812 ;
  assign n5814 = n4924 & ~n4951 ;
  assign n5815 = ~n5813 & n5814 ;
  assign n5816 = n5809 & ~n5815 ;
  assign n5817 = ~n5799 & n5816 ;
  assign n5818 = ~n4917 & ~n5803 ;
  assign n5819 = n4933 & ~n4934 ;
  assign n5820 = ~n4917 & ~n5819 ;
  assign n5821 = n5805 & n5820 ;
  assign n5822 = ~n5818 & ~n5821 ;
  assign n5823 = ~n4911 & n5822 ;
  assign n5824 = n4913 & ~n5823 ;
  assign n5825 = ~n4934 & ~n5788 ;
  assign n5826 = ~n4928 & ~n5825 ;
  assign n5827 = ~n4928 & n5794 ;
  assign n5828 = ~n5803 & n5827 ;
  assign n5829 = ~n5826 & ~n5828 ;
  assign n5830 = ~n5796 & n5829 ;
  assign n5831 = ~\s11_msel_arb1_state_reg[1]/NET0131  & ~\s11_msel_arb1_state_reg[2]/NET0131  ;
  assign n5832 = ~n5830 & n5831 ;
  assign n5833 = ~n5824 & ~n5832 ;
  assign n5834 = n5817 & n5833 ;
  assign n5835 = ~\s11_msel_arb2_state_reg[1]/NET0131  & \s11_msel_arb2_state_reg[2]/NET0131  ;
  assign n5836 = ~n4248 & n5835 ;
  assign n5837 = n4247 & n5836 ;
  assign n5838 = ~n4251 & n4268 ;
  assign n5839 = n4254 & ~n4257 ;
  assign n5840 = ~n4251 & ~n4262 ;
  assign n5841 = ~n5839 & n5840 ;
  assign n5842 = ~n5838 & ~n5841 ;
  assign n5843 = ~n4250 & n5836 ;
  assign n5844 = n5842 & n5843 ;
  assign n5845 = ~n5837 & ~n5844 ;
  assign n5846 = ~\s11_msel_arb2_state_reg[0]/NET0131  & ~n5845 ;
  assign n5847 = ~n4248 & ~n4257 ;
  assign n5848 = ~n5839 & ~n5847 ;
  assign n5849 = ~n4250 & n4251 ;
  assign n5850 = ~n4247 & ~n5849 ;
  assign n5851 = ~n4250 & ~n4268 ;
  assign n5852 = n4262 & n5851 ;
  assign n5853 = n5850 & ~n5852 ;
  assign n5854 = \s11_msel_arb2_state_reg[0]/NET0131  & n5851 ;
  assign n5855 = ~n5839 & ~n5854 ;
  assign n5856 = n5853 & n5855 ;
  assign n5857 = ~n5848 & ~n5856 ;
  assign n5858 = \s11_msel_arb2_state_reg[1]/NET0131  & ~\s11_msel_arb2_state_reg[2]/NET0131  ;
  assign n5859 = ~\s11_msel_arb2_state_reg[0]/NET0131  & n5858 ;
  assign n5860 = n5857 & n5859 ;
  assign n5861 = ~n5846 & ~n5860 ;
  assign n5862 = \s11_msel_arb2_state_reg[0]/NET0131  & ~n4250 ;
  assign n5863 = ~n4247 & ~n5862 ;
  assign n5864 = ~n4268 & n5847 ;
  assign n5865 = ~n5863 & n5864 ;
  assign n5866 = ~n5842 & ~n5865 ;
  assign n5867 = \rf_conf11_reg[13]/NET0131  & ~\s11_msel_arb2_state_reg[0]/NET0131  ;
  assign n5868 = n2747 & n5867 ;
  assign n5869 = \s11_msel_arb2_state_reg[1]/NET0131  & \s11_msel_arb2_state_reg[2]/NET0131  ;
  assign n5870 = ~n5868 & n5869 ;
  assign n5871 = ~n5866 & n5870 ;
  assign n5872 = ~n4248 & ~n5853 ;
  assign n5873 = n5847 & n5854 ;
  assign n5874 = ~n4254 & ~n5873 ;
  assign n5875 = ~n5872 & n5874 ;
  assign n5876 = \s11_msel_arb2_state_reg[0]/NET0131  & n5858 ;
  assign n5877 = ~n5875 & n5876 ;
  assign n5878 = ~n5871 & ~n5877 ;
  assign n5879 = \s11_msel_arb2_state_reg[0]/NET0131  & ~\s11_msel_arb2_state_reg[1]/NET0131  ;
  assign n5880 = \s11_msel_arb2_state_reg[2]/NET0131  & n5879 ;
  assign n5881 = ~n4250 & n5842 ;
  assign n5882 = ~n4247 & ~n5873 ;
  assign n5883 = ~n5881 & n5882 ;
  assign n5884 = n5880 & ~n5883 ;
  assign n5885 = ~n4262 & ~n5839 ;
  assign n5886 = \rf_conf11_reg[1]/NET0131  & ~\s11_msel_arb2_state_reg[0]/NET0131  ;
  assign n5887 = n2752 & n5886 ;
  assign n5888 = ~n5885 & ~n5887 ;
  assign n5889 = n5847 & ~n5887 ;
  assign n5890 = ~n5850 & n5889 ;
  assign n5891 = ~n5888 & ~n5890 ;
  assign n5892 = ~n5873 & n5891 ;
  assign n5893 = ~\s11_msel_arb2_state_reg[1]/NET0131  & ~\s11_msel_arb2_state_reg[2]/NET0131  ;
  assign n5894 = ~n5892 & n5893 ;
  assign n5895 = ~n5884 & ~n5894 ;
  assign n5896 = n5878 & n5895 ;
  assign n5897 = n5861 & n5896 ;
  assign n5898 = ~n4291 & ~n4308 ;
  assign n5899 = n4289 & ~n4291 ;
  assign n5900 = ~n5898 & ~n5899 ;
  assign n5901 = ~n4295 & n4299 ;
  assign n5902 = n4284 & ~n4286 ;
  assign n5903 = ~n4295 & ~n4297 ;
  assign n5904 = ~n5902 & n5903 ;
  assign n5905 = ~n5901 & ~n5904 ;
  assign n5906 = \s11_msel_arb3_state_reg[0]/NET0131  & ~n4299 ;
  assign n5907 = ~n4286 & n5906 ;
  assign n5908 = ~n5899 & ~n5907 ;
  assign n5909 = ~n5905 & n5908 ;
  assign n5910 = ~n5900 & ~n5909 ;
  assign n5911 = n4325 & n5910 ;
  assign n5912 = ~\s11_msel_arb3_state_reg[1]/NET0131  & ~\s11_msel_arb3_state_reg[2]/NET0131  ;
  assign n5913 = n5902 & n5912 ;
  assign n5914 = ~n4289 & n4308 ;
  assign n5915 = n4297 & ~n4299 ;
  assign n5916 = ~n4289 & ~n4295 ;
  assign n5917 = ~n5915 & n5916 ;
  assign n5918 = ~n5914 & ~n5917 ;
  assign n5919 = ~n4286 & ~n4291 ;
  assign n5920 = n5912 & n5919 ;
  assign n5921 = n5918 & n5920 ;
  assign n5922 = ~n5913 & ~n5921 ;
  assign n5923 = n4282 & ~n4308 ;
  assign n5924 = n4295 & n5923 ;
  assign n5925 = ~n4297 & ~n5902 ;
  assign n5926 = ~n4286 & n5899 ;
  assign n5927 = n5925 & ~n5926 ;
  assign n5928 = ~n4299 & n5923 ;
  assign n5929 = ~n5927 & n5928 ;
  assign n5930 = ~n5924 & ~n5929 ;
  assign n5931 = ~\s11_msel_arb3_state_reg[0]/NET0131  & n5930 ;
  assign n5932 = n5922 & n5931 ;
  assign n5933 = ~n5911 & n5932 ;
  assign n5934 = ~n4299 & ~n5927 ;
  assign n5935 = ~n4286 & ~n4299 ;
  assign n5936 = n5898 & n5935 ;
  assign n5937 = ~n4295 & ~n5936 ;
  assign n5938 = ~n5934 & n5937 ;
  assign n5939 = n4282 & ~n5938 ;
  assign n5940 = n4289 & n4325 ;
  assign n5941 = \s11_msel_arb3_state_reg[0]/NET0131  & ~n5940 ;
  assign n5942 = ~n5939 & n5941 ;
  assign n5943 = ~n5933 & ~n5942 ;
  assign n5944 = ~n4284 & n4291 ;
  assign n5945 = ~n4286 & ~n4308 ;
  assign n5946 = n5906 & n5945 ;
  assign n5947 = ~n4284 & ~n5946 ;
  assign n5948 = ~n5918 & n5947 ;
  assign n5949 = ~n5944 & ~n5948 ;
  assign n5950 = \s11_msel_arb3_state_reg[0]/NET0131  & n5912 ;
  assign n5951 = n5949 & n5950 ;
  assign n5952 = ~n4295 & ~n5906 ;
  assign n5953 = ~n4286 & n5898 ;
  assign n5954 = ~n5952 & n5953 ;
  assign n5955 = n5927 & ~n5954 ;
  assign n5956 = \rf_conf11_reg[13]/NET0131  & ~\s11_msel_arb3_state_reg[0]/NET0131  ;
  assign n5957 = n4298 & n5956 ;
  assign n5958 = n4305 & ~n5957 ;
  assign n5959 = ~n5955 & n5958 ;
  assign n5960 = n5906 & n5919 ;
  assign n5961 = ~n5905 & ~n5960 ;
  assign n5962 = \s11_msel_arb3_state_reg[0]/NET0131  & n4325 ;
  assign n5963 = ~n4289 & n5962 ;
  assign n5964 = ~n4308 & n5963 ;
  assign n5965 = ~n5961 & n5964 ;
  assign n5966 = ~n5959 & ~n5965 ;
  assign n5967 = ~n5951 & n5966 ;
  assign n5968 = ~n5943 & n5967 ;
  assign n5969 = ~n2813 & n2826 ;
  assign n5970 = n2808 & ~n2810 ;
  assign n5971 = ~n2805 & n5970 ;
  assign n5972 = ~n2810 & ~n2815 ;
  assign n5973 = \s12_msel_arb0_state_reg[0]/NET0131  & ~n2805 ;
  assign n5974 = n5972 & n5973 ;
  assign n5975 = ~n5971 & ~n5974 ;
  assign n5976 = n2805 & ~n2820 ;
  assign n5977 = ~n2803 & ~n2820 ;
  assign n5978 = ~n5976 & ~n5977 ;
  assign n5979 = ~n2813 & ~n5978 ;
  assign n5980 = n5975 & n5979 ;
  assign n5981 = ~n5969 & ~n5980 ;
  assign n5982 = n2849 & n5981 ;
  assign n5983 = \s12_msel_arb0_state_reg[1]/NET0131  & \s12_msel_arb0_state_reg[2]/NET0131  ;
  assign n5984 = n2820 & ~n2826 ;
  assign n5985 = ~n2813 & ~n5984 ;
  assign n5986 = ~n2815 & ~n5985 ;
  assign n5987 = ~n2805 & ~n2826 ;
  assign n5988 = ~\s12_msel_arb0_state_reg[0]/NET0131  & ~n2803 ;
  assign n5989 = n5987 & ~n5988 ;
  assign n5990 = ~n2803 & n2810 ;
  assign n5991 = ~n2815 & ~n5990 ;
  assign n5992 = n5989 & n5991 ;
  assign n5993 = ~n5986 & ~n5992 ;
  assign n5994 = ~n2808 & n5993 ;
  assign n5995 = n5983 & ~n5994 ;
  assign n5996 = n2813 & ~n2815 ;
  assign n5997 = ~n2803 & ~n2808 ;
  assign n5998 = ~n5996 & n5997 ;
  assign n5999 = ~n5990 & ~n5998 ;
  assign n6000 = \s12_msel_arb0_state_reg[0]/NET0131  & ~n2826 ;
  assign n6001 = n5972 & n6000 ;
  assign n6002 = ~n2820 & ~n6001 ;
  assign n6003 = ~n5999 & n6002 ;
  assign n6004 = \s12_msel_arb0_state_reg[1]/NET0131  & ~\s12_msel_arb0_state_reg[2]/NET0131  ;
  assign n6005 = ~n5976 & n6004 ;
  assign n6006 = ~n6003 & n6005 ;
  assign n6007 = ~n5995 & ~n6006 ;
  assign n6008 = ~n5982 & n6007 ;
  assign n6009 = \s12_msel_arb0_state_reg[0]/NET0131  & ~n6008 ;
  assign n6010 = \s12_msel_arb0_state_reg[0]/NET0131  & n5972 ;
  assign n6011 = n5987 & n6010 ;
  assign n6012 = n5987 & ~n5990 ;
  assign n6013 = ~n5998 & n6012 ;
  assign n6014 = ~n6011 & ~n6013 ;
  assign n6015 = ~n5984 & n6014 ;
  assign n6016 = n6004 & ~n6015 ;
  assign n6017 = n5970 & n5983 ;
  assign n6018 = n5985 & ~n5989 ;
  assign n6019 = n5972 & n5983 ;
  assign n6020 = ~n6018 & n6019 ;
  assign n6021 = ~n6017 & ~n6020 ;
  assign n6022 = n2849 & n5996 ;
  assign n6023 = ~n2805 & ~n2810 ;
  assign n6024 = ~\s12_msel_arb0_state_reg[0]/NET0131  & ~n2808 ;
  assign n6025 = n6023 & ~n6024 ;
  assign n6026 = ~n5978 & ~n6025 ;
  assign n6027 = ~n2815 & ~n2826 ;
  assign n6028 = n2849 & n6027 ;
  assign n6029 = ~n6026 & n6028 ;
  assign n6030 = ~n6022 & ~n6029 ;
  assign n6031 = n6021 & n6030 ;
  assign n6032 = ~n6016 & n6031 ;
  assign n6033 = ~\s12_msel_arb0_state_reg[0]/NET0131  & ~n6032 ;
  assign n6034 = \s12_msel_arb0_state_reg[0]/NET0131  & n6027 ;
  assign n6035 = n6023 & n6034 ;
  assign n6036 = n2853 & n6035 ;
  assign n6037 = n2820 & n6027 ;
  assign n6038 = n5998 & ~n6037 ;
  assign n6039 = ~\rf_conf12_reg[9]/NET0131  & ~\s12_msel_arb0_state_reg[0]/NET0131  ;
  assign n6040 = n2804 & n6039 ;
  assign n6041 = ~n5990 & ~n6040 ;
  assign n6042 = n2853 & n6041 ;
  assign n6043 = ~n6038 & n6042 ;
  assign n6044 = ~n6036 & ~n6043 ;
  assign n6045 = ~n6033 & n6044 ;
  assign n6046 = ~n6009 & n6045 ;
  assign n6047 = ~n4971 & n4972 ;
  assign n6048 = ~n4978 & ~n6047 ;
  assign n6049 = ~n4976 & ~n6048 ;
  assign n6050 = ~n4969 & ~n4971 ;
  assign n6051 = n4968 & ~n4976 ;
  assign n6052 = n6050 & n6051 ;
  assign n6053 = ~n4963 & ~n6052 ;
  assign n6054 = ~n6049 & n6053 ;
  assign n6055 = ~n4965 & ~n6054 ;
  assign n6056 = \s12_msel_arb1_state_reg[0]/NET0131  & ~n4976 ;
  assign n6057 = ~n4992 & n6056 ;
  assign n6058 = n6050 & n6057 ;
  assign n6059 = ~\s12_msel_arb1_state_reg[1]/NET0131  & ~n6058 ;
  assign n6060 = ~n6055 & n6059 ;
  assign n6061 = ~\s12_msel_arb1_state_reg[2]/NET0131  & n6060 ;
  assign n6062 = n4963 & ~n4992 ;
  assign n6063 = ~n4968 & ~n6062 ;
  assign n6064 = ~n6057 & n6063 ;
  assign n6065 = n6050 & ~n6064 ;
  assign n6066 = \s12_msel_arb1_state_reg[0]/NET0131  & ~n4978 ;
  assign n6067 = ~n6047 & n6066 ;
  assign n6068 = ~n6065 & n6067 ;
  assign n6069 = n4969 & ~n4972 ;
  assign n6070 = ~n4968 & ~n4972 ;
  assign n6071 = ~n6062 & n6070 ;
  assign n6072 = ~n6069 & ~n6071 ;
  assign n6073 = ~n4971 & ~n4976 ;
  assign n6074 = n6072 & n6073 ;
  assign n6075 = ~n4976 & n4978 ;
  assign n6076 = ~\s12_msel_arb1_state_reg[0]/NET0131  & ~n6075 ;
  assign n6077 = ~n6074 & n6076 ;
  assign n6078 = ~n6068 & ~n6077 ;
  assign n6079 = \s12_msel_arb1_state_reg[1]/NET0131  & ~\s12_msel_arb1_state_reg[2]/NET0131  ;
  assign n6080 = ~n6078 & n6079 ;
  assign n6081 = ~n6061 & ~n6080 ;
  assign n6082 = ~n4969 & ~n4992 ;
  assign n6083 = n6075 & n6082 ;
  assign n6084 = ~n6072 & ~n6083 ;
  assign n6085 = ~\s12_msel_arb1_state_reg[1]/NET0131  & ~n4987 ;
  assign n6086 = ~n6084 & n6085 ;
  assign n6087 = ~n4976 & ~n4992 ;
  assign n6088 = ~n6048 & n6087 ;
  assign n6089 = n6063 & ~n6088 ;
  assign n6090 = n4985 & ~n6089 ;
  assign n6091 = \s12_msel_arb1_state_reg[2]/NET0131  & ~n6058 ;
  assign n6092 = ~n6090 & n6091 ;
  assign n6093 = ~n6086 & n6092 ;
  assign n6094 = n6081 & ~n6093 ;
  assign n6095 = \rf_conf12_reg[5]/NET0131  & n2825 ;
  assign n6096 = \rf_conf12_reg[7]/NET0131  & n2819 ;
  assign n6097 = ~n6095 & n6096 ;
  assign n6098 = \s12_msel_arb2_state_reg[1]/NET0131  & ~\s12_msel_arb2_state_reg[2]/NET0131  ;
  assign n6099 = n6097 & n6098 ;
  assign n6100 = \rf_conf12_reg[11]/NET0131  & n2802 ;
  assign n6101 = \rf_conf12_reg[15]/NET0131  & n2807 ;
  assign n6102 = \rf_conf12_reg[13]/NET0131  & n2809 ;
  assign n6103 = n6101 & ~n6102 ;
  assign n6104 = ~n6100 & ~n6103 ;
  assign n6105 = \rf_conf12_reg[3]/NET0131  & n2812 ;
  assign n6106 = \rf_conf12_reg[1]/NET0131  & n2814 ;
  assign n6107 = ~n6102 & ~n6106 ;
  assign n6108 = n6105 & n6107 ;
  assign n6109 = n6104 & ~n6108 ;
  assign n6110 = \rf_conf12_reg[9]/NET0131  & n2804 ;
  assign n6111 = ~n6095 & ~n6110 ;
  assign n6112 = n6098 & n6111 ;
  assign n6113 = ~n6109 & n6112 ;
  assign n6114 = ~n6099 & ~n6113 ;
  assign n6115 = ~n6097 & ~n6105 ;
  assign n6116 = ~\s12_msel_arb2_state_reg[1]/NET0131  & ~\s12_msel_arb2_state_reg[2]/NET0131  ;
  assign n6117 = ~n6106 & n6116 ;
  assign n6118 = ~n6115 & n6117 ;
  assign n6119 = n6111 & n6117 ;
  assign n6120 = ~n6104 & n6119 ;
  assign n6121 = ~n6118 & ~n6120 ;
  assign n6122 = ~\s12_msel_arb2_state_reg[0]/NET0131  & n6121 ;
  assign n6123 = n6114 & n6122 ;
  assign n6124 = \s12_msel_arb2_state_reg[1]/NET0131  & \s12_msel_arb2_state_reg[2]/NET0131  ;
  assign n6125 = n6103 & n6124 ;
  assign n6126 = n6100 & n6111 ;
  assign n6127 = n6115 & ~n6126 ;
  assign n6128 = n6107 & n6124 ;
  assign n6129 = ~n6127 & n6128 ;
  assign n6130 = ~n6125 & ~n6129 ;
  assign n6131 = ~\s12_msel_arb2_state_reg[1]/NET0131  & \s12_msel_arb2_state_reg[2]/NET0131  ;
  assign n6132 = ~n6110 & n6131 ;
  assign n6133 = n6100 & n6132 ;
  assign n6134 = ~n6101 & n6106 ;
  assign n6135 = ~n6101 & ~n6105 ;
  assign n6136 = ~n6097 & n6135 ;
  assign n6137 = ~n6134 & ~n6136 ;
  assign n6138 = ~n6102 & n6132 ;
  assign n6139 = n6137 & n6138 ;
  assign n6140 = ~n6133 & ~n6139 ;
  assign n6141 = n6130 & n6140 ;
  assign n6142 = n6123 & n6141 ;
  assign n6143 = \s12_msel_arb2_state_reg[0]/NET0131  & ~n6106 ;
  assign n6144 = n6111 & n6143 ;
  assign n6145 = ~n6137 & ~n6144 ;
  assign n6146 = \s12_msel_arb2_state_reg[0]/NET0131  & n6131 ;
  assign n6147 = ~n6100 & n6146 ;
  assign n6148 = ~n6102 & n6147 ;
  assign n6149 = ~n6145 & n6148 ;
  assign n6150 = n6142 & ~n6149 ;
  assign n6151 = ~n6104 & n6111 ;
  assign n6152 = n6115 & ~n6151 ;
  assign n6153 = \s12_msel_arb2_state_reg[0]/NET0131  & n6111 ;
  assign n6154 = n6107 & n6153 ;
  assign n6155 = n6152 & ~n6154 ;
  assign n6156 = n6116 & ~n6155 ;
  assign n6157 = n6096 & n6098 ;
  assign n6158 = n6095 & ~n6105 ;
  assign n6159 = n6107 & ~n6158 ;
  assign n6160 = n6104 & ~n6159 ;
  assign n6161 = n6098 & ~n6110 ;
  assign n6162 = ~n6160 & n6161 ;
  assign n6163 = ~n6157 & ~n6162 ;
  assign n6164 = n6100 & n6131 ;
  assign n6165 = \s12_msel_arb2_state_reg[0]/NET0131  & ~n6164 ;
  assign n6166 = n6163 & n6165 ;
  assign n6167 = ~n6156 & n6166 ;
  assign n6168 = \s12_msel_arb2_state_reg[0]/NET0131  & ~n6102 ;
  assign n6169 = n6111 & n6168 ;
  assign n6170 = ~n6101 & ~n6169 ;
  assign n6171 = n6127 & n6170 ;
  assign n6172 = ~n6134 & ~n6171 ;
  assign n6173 = n6124 & n6172 ;
  assign n6174 = ~n6149 & ~n6173 ;
  assign n6175 = n6167 & n6174 ;
  assign n6176 = ~n6150 & ~n6175 ;
  assign n6177 = \s12_msel_arb3_state_reg[1]/NET0131  & ~\s12_msel_arb3_state_reg[2]/NET0131  ;
  assign n6178 = ~n4367 & n6177 ;
  assign n6179 = ~n4334 & ~n4346 ;
  assign n6180 = ~n4334 & n4348 ;
  assign n6181 = ~n6179 & ~n6180 ;
  assign n6182 = n6178 & n6181 ;
  assign n6183 = ~n4356 & ~n4374 ;
  assign n6184 = ~n4348 & ~n4358 ;
  assign n6185 = n6178 & n6184 ;
  assign n6186 = ~n6183 & n6185 ;
  assign n6187 = ~n6182 & ~n6186 ;
  assign n6188 = ~n4336 & ~n6187 ;
  assign n6189 = n4351 & ~n4353 ;
  assign n6190 = ~n4356 & ~n6189 ;
  assign n6191 = ~n4358 & ~n6190 ;
  assign n6192 = n6179 & ~n6191 ;
  assign n6193 = ~\s12_msel_arb3_state_reg[0]/NET0131  & \s12_msel_arb3_state_reg[2]/NET0131  ;
  assign n6194 = ~\s12_msel_arb3_state_reg[1]/NET0131  & n6193 ;
  assign n6195 = ~n6180 & n6194 ;
  assign n6196 = ~n4336 & n6195 ;
  assign n6197 = ~n6192 & n6196 ;
  assign n6198 = ~n6188 & ~n6197 ;
  assign n6199 = ~\s12_msel_arb3_state_reg[1]/NET0131  & ~\s12_msel_arb3_state_reg[2]/NET0131  ;
  assign n6200 = \rf_conf12_reg[1]/NET0131  & ~\s12_msel_arb3_state_reg[0]/NET0131  ;
  assign n6201 = n4357 & n6200 ;
  assign n6202 = n6199 & ~n6201 ;
  assign n6203 = ~n6190 & n6202 ;
  assign n6204 = ~n4336 & ~n4353 ;
  assign n6205 = n6202 & n6204 ;
  assign n6206 = n6181 & n6205 ;
  assign n6207 = ~n6203 & ~n6206 ;
  assign n6208 = n4351 & n6178 ;
  assign n6209 = ~\s12_msel_arb3_state_reg[1]/NET0131  & n4339 ;
  assign n6210 = n4334 & n6209 ;
  assign n6211 = ~n6208 & ~n6210 ;
  assign n6212 = n6207 & n6211 ;
  assign n6213 = n6198 & n6212 ;
  assign n6214 = \s12_msel_arb3_state_reg[0]/NET0131  & n6199 ;
  assign n6215 = ~n4358 & n6214 ;
  assign n6216 = n6204 & n6215 ;
  assign n6217 = ~n4334 & n6209 ;
  assign n6218 = ~n6216 & ~n6217 ;
  assign n6219 = ~n4346 & n4358 ;
  assign n6220 = ~n4346 & ~n4356 ;
  assign n6221 = ~n6189 & n6220 ;
  assign n6222 = ~n6219 & ~n6221 ;
  assign n6223 = \s12_msel_arb3_state_reg[0]/NET0131  & ~n4358 ;
  assign n6224 = n6204 & n6223 ;
  assign n6225 = ~n6216 & ~n6224 ;
  assign n6226 = ~n6222 & n6225 ;
  assign n6227 = ~n6218 & ~n6226 ;
  assign n6228 = ~n4348 & n6227 ;
  assign n6229 = ~n4358 & n6204 ;
  assign n6230 = ~\s12_msel_arb3_state_reg[0]/NET0131  & ~n4334 ;
  assign n6231 = n6229 & ~n6230 ;
  assign n6232 = ~n6222 & ~n6231 ;
  assign n6233 = ~\s12_msel_arb3_state_reg[0]/NET0131  & n4348 ;
  assign n6234 = n4348 & n6179 ;
  assign n6235 = n6190 & n6234 ;
  assign n6236 = ~n6233 & ~n6235 ;
  assign n6237 = n4381 & n6236 ;
  assign n6238 = ~n6232 & n6237 ;
  assign n6239 = ~n6228 & ~n6238 ;
  assign n6240 = n6213 & n6239 ;
  assign n6241 = ~n2875 & n2888 ;
  assign n6242 = n2870 & ~n2872 ;
  assign n6243 = ~n2867 & n6242 ;
  assign n6244 = ~n2872 & ~n2877 ;
  assign n6245 = \s13_msel_arb0_state_reg[0]/NET0131  & ~n2867 ;
  assign n6246 = n6244 & n6245 ;
  assign n6247 = ~n6243 & ~n6246 ;
  assign n6248 = n2867 & ~n2882 ;
  assign n6249 = ~n2865 & ~n2882 ;
  assign n6250 = ~n6248 & ~n6249 ;
  assign n6251 = ~n2875 & ~n6250 ;
  assign n6252 = n6247 & n6251 ;
  assign n6253 = ~n6241 & ~n6252 ;
  assign n6254 = n2911 & n6253 ;
  assign n6255 = \s13_msel_arb0_state_reg[1]/NET0131  & \s13_msel_arb0_state_reg[2]/NET0131  ;
  assign n6256 = n2882 & ~n2888 ;
  assign n6257 = ~n2875 & ~n6256 ;
  assign n6258 = ~n2877 & ~n6257 ;
  assign n6259 = ~n2867 & ~n2888 ;
  assign n6260 = ~\s13_msel_arb0_state_reg[0]/NET0131  & ~n2865 ;
  assign n6261 = n6259 & ~n6260 ;
  assign n6262 = ~n2865 & n2872 ;
  assign n6263 = ~n2877 & ~n6262 ;
  assign n6264 = n6261 & n6263 ;
  assign n6265 = ~n6258 & ~n6264 ;
  assign n6266 = ~n2870 & n6265 ;
  assign n6267 = n6255 & ~n6266 ;
  assign n6268 = n2875 & ~n2877 ;
  assign n6269 = ~n2865 & ~n2870 ;
  assign n6270 = ~n6268 & n6269 ;
  assign n6271 = ~n6262 & ~n6270 ;
  assign n6272 = \s13_msel_arb0_state_reg[0]/NET0131  & ~n2888 ;
  assign n6273 = n6244 & n6272 ;
  assign n6274 = ~n2882 & ~n6273 ;
  assign n6275 = ~n6271 & n6274 ;
  assign n6276 = \s13_msel_arb0_state_reg[1]/NET0131  & ~\s13_msel_arb0_state_reg[2]/NET0131  ;
  assign n6277 = ~n6248 & n6276 ;
  assign n6278 = ~n6275 & n6277 ;
  assign n6279 = ~n6267 & ~n6278 ;
  assign n6280 = ~n6254 & n6279 ;
  assign n6281 = \s13_msel_arb0_state_reg[0]/NET0131  & ~n6280 ;
  assign n6282 = \s13_msel_arb0_state_reg[0]/NET0131  & n6244 ;
  assign n6283 = n6259 & n6282 ;
  assign n6284 = n6259 & ~n6262 ;
  assign n6285 = ~n6270 & n6284 ;
  assign n6286 = ~n6283 & ~n6285 ;
  assign n6287 = ~n6256 & n6286 ;
  assign n6288 = n6276 & ~n6287 ;
  assign n6289 = n6242 & n6255 ;
  assign n6290 = n6257 & ~n6261 ;
  assign n6291 = n6244 & n6255 ;
  assign n6292 = ~n6290 & n6291 ;
  assign n6293 = ~n6289 & ~n6292 ;
  assign n6294 = n2911 & n6268 ;
  assign n6295 = ~n2867 & ~n2872 ;
  assign n6296 = ~\s13_msel_arb0_state_reg[0]/NET0131  & ~n2870 ;
  assign n6297 = n6295 & ~n6296 ;
  assign n6298 = ~n6250 & ~n6297 ;
  assign n6299 = ~n2877 & ~n2888 ;
  assign n6300 = n2911 & n6299 ;
  assign n6301 = ~n6298 & n6300 ;
  assign n6302 = ~n6294 & ~n6301 ;
  assign n6303 = n6293 & n6302 ;
  assign n6304 = ~n6288 & n6303 ;
  assign n6305 = ~\s13_msel_arb0_state_reg[0]/NET0131  & ~n6304 ;
  assign n6306 = \s13_msel_arb0_state_reg[0]/NET0131  & n6299 ;
  assign n6307 = n6295 & n6306 ;
  assign n6308 = n2915 & n6307 ;
  assign n6309 = n2882 & n6299 ;
  assign n6310 = n6270 & ~n6309 ;
  assign n6311 = ~\rf_conf13_reg[9]/NET0131  & ~\s13_msel_arb0_state_reg[0]/NET0131  ;
  assign n6312 = n2866 & n6311 ;
  assign n6313 = ~n6262 & ~n6312 ;
  assign n6314 = n2915 & n6313 ;
  assign n6315 = ~n6310 & n6314 ;
  assign n6316 = ~n6308 & ~n6315 ;
  assign n6317 = ~n6305 & n6316 ;
  assign n6318 = ~n6281 & n6317 ;
  assign n6319 = ~n4999 & ~n5012 ;
  assign n6320 = ~n4999 & n5013 ;
  assign n6321 = ~n5001 & ~n6320 ;
  assign n6322 = ~n6319 & n6321 ;
  assign n6323 = ~n5001 & ~n5013 ;
  assign n6324 = n5008 & ~n5009 ;
  assign n6325 = n6323 & n6324 ;
  assign n6326 = ~n5006 & ~n6325 ;
  assign n6327 = ~n6322 & n6326 ;
  assign n6328 = \s13_msel_arb1_state_reg[1]/NET0131  & ~\s13_msel_arb1_state_reg[2]/NET0131  ;
  assign n6329 = ~n5005 & n6328 ;
  assign n6330 = ~n6327 & n6329 ;
  assign n6331 = ~\s13_msel_arb1_state_reg[0]/NET0131  & n6330 ;
  assign n6332 = n4999 & ~n5001 ;
  assign n6333 = ~n6323 & ~n6332 ;
  assign n6334 = n5009 & ~n5012 ;
  assign n6335 = ~n5005 & n5006 ;
  assign n6336 = ~n5008 & ~n5012 ;
  assign n6337 = ~n6335 & n6336 ;
  assign n6338 = ~n6334 & ~n6337 ;
  assign n6339 = \s13_msel_arb1_state_reg[0]/NET0131  & ~n5009 ;
  assign n6340 = ~n5005 & n6339 ;
  assign n6341 = ~n6332 & ~n6340 ;
  assign n6342 = ~n6338 & n6341 ;
  assign n6343 = ~n6333 & ~n6342 ;
  assign n6344 = ~\s13_msel_arb1_state_reg[1]/NET0131  & \s13_msel_arb1_state_reg[2]/NET0131  ;
  assign n6345 = ~\s13_msel_arb1_state_reg[0]/NET0131  & n6344 ;
  assign n6346 = n6343 & n6345 ;
  assign n6347 = ~n6331 & ~n6346 ;
  assign n6348 = ~n5006 & ~n6322 ;
  assign n6349 = ~n6324 & ~n6340 ;
  assign n6350 = n6323 & ~n6349 ;
  assign n6351 = n6348 & ~n6350 ;
  assign n6352 = n6328 & ~n6351 ;
  assign n6353 = ~\s13_msel_arb1_state_reg[1]/NET0131  & ~\s13_msel_arb1_state_reg[2]/NET0131  ;
  assign n6354 = ~n5008 & ~n6335 ;
  assign n6355 = ~n5005 & n6332 ;
  assign n6356 = n6354 & ~n6355 ;
  assign n6357 = ~n5005 & n6323 ;
  assign n6358 = ~n5012 & ~n6339 ;
  assign n6359 = n6357 & ~n6358 ;
  assign n6360 = n6356 & ~n6359 ;
  assign n6361 = n6353 & ~n6360 ;
  assign n6362 = ~n5001 & ~n5005 ;
  assign n6363 = n6339 & n6362 ;
  assign n6364 = ~n4999 & ~n6363 ;
  assign n6365 = ~n6338 & n6364 ;
  assign n6366 = ~n6320 & n6344 ;
  assign n6367 = ~n6365 & n6366 ;
  assign n6368 = ~n6361 & ~n6367 ;
  assign n6369 = ~n6352 & n6368 ;
  assign n6370 = \s13_msel_arb1_state_reg[0]/NET0131  & ~n6369 ;
  assign n6371 = ~\rf_conf13_reg[13]/NET0131  & ~\s13_msel_arb1_state_reg[0]/NET0131  ;
  assign n6372 = n3862 & n6371 ;
  assign n6373 = \s13_msel_arb1_state_reg[1]/NET0131  & \s13_msel_arb1_state_reg[2]/NET0131  ;
  assign n6374 = ~n6372 & n6373 ;
  assign n6375 = n5012 & n6374 ;
  assign n6376 = \s13_msel_arb1_state_reg[0]/NET0131  & ~n5005 ;
  assign n6377 = n6323 & n6376 ;
  assign n6378 = n6356 & ~n6377 ;
  assign n6379 = n6374 & ~n6378 ;
  assign n6380 = ~n5009 & n6379 ;
  assign n6381 = ~n5005 & ~n6319 ;
  assign n6382 = n6321 & n6381 ;
  assign n6383 = ~n6335 & ~n6382 ;
  assign n6384 = ~n5008 & n6383 ;
  assign n6385 = ~\s13_msel_arb1_state_reg[0]/NET0131  & n6353 ;
  assign n6386 = ~n5009 & n6385 ;
  assign n6387 = ~n6384 & n6386 ;
  assign n6388 = ~n6380 & ~n6387 ;
  assign n6389 = ~n6375 & n6388 ;
  assign n6390 = ~n6370 & n6389 ;
  assign n6391 = n6347 & n6390 ;
  assign n6392 = \rf_conf13_reg[9]/NET0131  & n2866 ;
  assign n6393 = \rf_conf13_reg[15]/NET0131  & n2869 ;
  assign n6394 = \rf_conf13_reg[1]/NET0131  & n2876 ;
  assign n6395 = ~n6393 & n6394 ;
  assign n6396 = \rf_conf13_reg[7]/NET0131  & n2881 ;
  assign n6397 = \rf_conf13_reg[5]/NET0131  & n2887 ;
  assign n6398 = n6396 & ~n6397 ;
  assign n6399 = \rf_conf13_reg[3]/NET0131  & n2874 ;
  assign n6400 = ~n6393 & ~n6399 ;
  assign n6401 = ~n6398 & n6400 ;
  assign n6402 = ~n6395 & ~n6401 ;
  assign n6403 = \rf_conf13_reg[11]/NET0131  & n2864 ;
  assign n6404 = ~n6402 & ~n6403 ;
  assign n6405 = \rf_conf13_reg[13]/NET0131  & n2871 ;
  assign n6406 = ~n6403 & n6405 ;
  assign n6407 = \s13_msel_arb2_state_reg[0]/NET0131  & ~n6406 ;
  assign n6408 = ~n6404 & n6407 ;
  assign n6409 = n6392 & ~n6408 ;
  assign n6410 = ~n6394 & ~n6405 ;
  assign n6411 = \s13_msel_arb2_state_reg[0]/NET0131  & ~n6397 ;
  assign n6412 = n6410 & n6411 ;
  assign n6413 = n6406 & ~n6412 ;
  assign n6414 = ~n6403 & ~n6412 ;
  assign n6415 = ~n6402 & n6414 ;
  assign n6416 = ~n6413 & ~n6415 ;
  assign n6417 = ~\s13_msel_arb2_state_reg[1]/NET0131  & \s13_msel_arb2_state_reg[2]/NET0131  ;
  assign n6418 = n6416 & n6417 ;
  assign n6419 = ~n6409 & n6418 ;
  assign n6420 = \s13_msel_arb2_state_reg[1]/NET0131  & \s13_msel_arb2_state_reg[2]/NET0131  ;
  assign n6421 = n6393 & ~n6405 ;
  assign n6422 = n6420 & n6421 ;
  assign n6423 = ~n6398 & ~n6399 ;
  assign n6424 = ~\s13_msel_arb2_state_reg[0]/NET0131  & ~n6403 ;
  assign n6425 = ~n6392 & ~n6397 ;
  assign n6426 = ~n6424 & n6425 ;
  assign n6427 = n6423 & ~n6426 ;
  assign n6428 = n6410 & n6420 ;
  assign n6429 = ~n6427 & n6428 ;
  assign n6430 = ~n6422 & ~n6429 ;
  assign n6431 = ~\s13_msel_arb2_state_reg[1]/NET0131  & ~\s13_msel_arb2_state_reg[2]/NET0131  ;
  assign n6432 = ~n6394 & n6399 ;
  assign n6433 = n6431 & n6432 ;
  assign n6434 = n6392 & ~n6396 ;
  assign n6435 = ~n6396 & ~n6403 ;
  assign n6436 = ~n6421 & n6435 ;
  assign n6437 = ~n6434 & ~n6436 ;
  assign n6438 = ~n6394 & ~n6397 ;
  assign n6439 = n6431 & n6438 ;
  assign n6440 = n6437 & n6439 ;
  assign n6441 = ~n6433 & ~n6440 ;
  assign n6442 = n6430 & n6441 ;
  assign n6443 = ~\s13_msel_arb2_state_reg[0]/NET0131  & ~n6442 ;
  assign n6444 = n6399 & n6431 ;
  assign n6445 = \s13_msel_arb2_state_reg[0]/NET0131  & n6444 ;
  assign n6446 = ~n6394 & ~n6406 ;
  assign n6447 = n6426 & n6446 ;
  assign n6448 = ~n6402 & ~n6447 ;
  assign n6449 = \s13_msel_arb2_state_reg[0]/NET0131  & n6420 ;
  assign n6450 = ~n6448 & n6449 ;
  assign n6451 = ~n6445 & ~n6450 ;
  assign n6452 = ~n6399 & n6431 ;
  assign n6453 = n6411 & n6452 ;
  assign n6454 = \rf_conf13_reg[5]/NET0131  & ~\s13_msel_arb2_state_reg[0]/NET0131  ;
  assign n6455 = n2887 & n6454 ;
  assign n6456 = \s13_msel_arb2_state_reg[1]/NET0131  & ~\s13_msel_arb2_state_reg[2]/NET0131  ;
  assign n6457 = ~n6455 & n6456 ;
  assign n6458 = ~n6453 & ~n6457 ;
  assign n6459 = n6437 & ~n6458 ;
  assign n6460 = n6410 & n6453 ;
  assign n6461 = ~n6392 & n6460 ;
  assign n6462 = ~n6405 & n6432 ;
  assign n6463 = ~n6412 & ~n6462 ;
  assign n6464 = ~n6392 & n6457 ;
  assign n6465 = ~n6463 & n6464 ;
  assign n6466 = ~n6461 & ~n6465 ;
  assign n6467 = ~n6459 & n6466 ;
  assign n6468 = n6451 & n6467 ;
  assign n6469 = ~n6443 & n6468 ;
  assign n6470 = ~n6419 & n6469 ;
  assign n6471 = \s13_msel_arb3_state_reg[1]/NET0131  & ~\s13_msel_arb3_state_reg[2]/NET0131  ;
  assign n6472 = ~n3882 & n6471 ;
  assign n6473 = ~n3849 & ~n3861 ;
  assign n6474 = ~n3849 & n3863 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = n6472 & n6475 ;
  assign n6477 = ~n3871 & ~n3889 ;
  assign n6478 = ~n3863 & ~n3873 ;
  assign n6479 = n6472 & n6478 ;
  assign n6480 = ~n6477 & n6479 ;
  assign n6481 = ~n6476 & ~n6480 ;
  assign n6482 = ~n3851 & ~n6481 ;
  assign n6483 = n3866 & ~n3868 ;
  assign n6484 = ~n3871 & ~n6483 ;
  assign n6485 = ~n3873 & ~n6484 ;
  assign n6486 = n6473 & ~n6485 ;
  assign n6487 = ~\s13_msel_arb3_state_reg[0]/NET0131  & \s13_msel_arb3_state_reg[2]/NET0131  ;
  assign n6488 = ~\s13_msel_arb3_state_reg[1]/NET0131  & n6487 ;
  assign n6489 = ~n6474 & n6488 ;
  assign n6490 = ~n3851 & n6489 ;
  assign n6491 = ~n6486 & n6490 ;
  assign n6492 = ~n6482 & ~n6491 ;
  assign n6493 = ~\s13_msel_arb3_state_reg[1]/NET0131  & ~\s13_msel_arb3_state_reg[2]/NET0131  ;
  assign n6494 = \rf_conf13_reg[1]/NET0131  & ~\s13_msel_arb3_state_reg[0]/NET0131  ;
  assign n6495 = n3872 & n6494 ;
  assign n6496 = n6493 & ~n6495 ;
  assign n6497 = ~n6484 & n6496 ;
  assign n6498 = ~n3851 & ~n3868 ;
  assign n6499 = n6496 & n6498 ;
  assign n6500 = n6475 & n6499 ;
  assign n6501 = ~n6497 & ~n6500 ;
  assign n6502 = n3866 & n6472 ;
  assign n6503 = ~\s13_msel_arb3_state_reg[1]/NET0131  & n3854 ;
  assign n6504 = n3849 & n6503 ;
  assign n6505 = ~n6502 & ~n6504 ;
  assign n6506 = n6501 & n6505 ;
  assign n6507 = n6492 & n6506 ;
  assign n6508 = \s13_msel_arb3_state_reg[0]/NET0131  & n6493 ;
  assign n6509 = ~n3873 & n6508 ;
  assign n6510 = n6498 & n6509 ;
  assign n6511 = ~n3849 & n6503 ;
  assign n6512 = ~n6510 & ~n6511 ;
  assign n6513 = ~n3861 & n3873 ;
  assign n6514 = ~n3861 & ~n3871 ;
  assign n6515 = ~n6483 & n6514 ;
  assign n6516 = ~n6513 & ~n6515 ;
  assign n6517 = \s13_msel_arb3_state_reg[0]/NET0131  & ~n3873 ;
  assign n6518 = n6498 & n6517 ;
  assign n6519 = ~n6510 & ~n6518 ;
  assign n6520 = ~n6516 & n6519 ;
  assign n6521 = ~n6512 & ~n6520 ;
  assign n6522 = ~n3863 & n6521 ;
  assign n6523 = ~n3873 & n6498 ;
  assign n6524 = ~\s13_msel_arb3_state_reg[0]/NET0131  & ~n3849 ;
  assign n6525 = n6523 & ~n6524 ;
  assign n6526 = ~n6516 & ~n6525 ;
  assign n6527 = ~\s13_msel_arb3_state_reg[0]/NET0131  & n3863 ;
  assign n6528 = n3863 & n6473 ;
  assign n6529 = n6484 & n6528 ;
  assign n6530 = ~n6527 & ~n6529 ;
  assign n6531 = n3896 & n6530 ;
  assign n6532 = ~n6526 & n6531 ;
  assign n6533 = ~n6522 & ~n6532 ;
  assign n6534 = n6507 & n6533 ;
  assign n6535 = ~n2937 & n2950 ;
  assign n6536 = n2932 & ~n2934 ;
  assign n6537 = ~n2929 & n6536 ;
  assign n6538 = ~n2934 & ~n2939 ;
  assign n6539 = \s14_msel_arb0_state_reg[0]/NET0131  & ~n2929 ;
  assign n6540 = n6538 & n6539 ;
  assign n6541 = ~n6537 & ~n6540 ;
  assign n6542 = n2929 & ~n2944 ;
  assign n6543 = ~n2927 & ~n2944 ;
  assign n6544 = ~n6542 & ~n6543 ;
  assign n6545 = ~n2937 & ~n6544 ;
  assign n6546 = n6541 & n6545 ;
  assign n6547 = ~n6535 & ~n6546 ;
  assign n6548 = n2973 & n6547 ;
  assign n6549 = \s14_msel_arb0_state_reg[1]/NET0131  & \s14_msel_arb0_state_reg[2]/NET0131  ;
  assign n6550 = n2944 & ~n2950 ;
  assign n6551 = ~n2937 & ~n6550 ;
  assign n6552 = ~n2939 & ~n6551 ;
  assign n6553 = ~n2929 & ~n2950 ;
  assign n6554 = ~\s14_msel_arb0_state_reg[0]/NET0131  & ~n2927 ;
  assign n6555 = n6553 & ~n6554 ;
  assign n6556 = ~n2927 & n2934 ;
  assign n6557 = ~n2939 & ~n6556 ;
  assign n6558 = n6555 & n6557 ;
  assign n6559 = ~n6552 & ~n6558 ;
  assign n6560 = ~n2932 & n6559 ;
  assign n6561 = n6549 & ~n6560 ;
  assign n6562 = n2937 & ~n2939 ;
  assign n6563 = ~n2927 & ~n2932 ;
  assign n6564 = ~n6562 & n6563 ;
  assign n6565 = ~n6556 & ~n6564 ;
  assign n6566 = \s14_msel_arb0_state_reg[0]/NET0131  & ~n2950 ;
  assign n6567 = n6538 & n6566 ;
  assign n6568 = ~n2944 & ~n6567 ;
  assign n6569 = ~n6565 & n6568 ;
  assign n6570 = \s14_msel_arb0_state_reg[1]/NET0131  & ~\s14_msel_arb0_state_reg[2]/NET0131  ;
  assign n6571 = ~n6542 & n6570 ;
  assign n6572 = ~n6569 & n6571 ;
  assign n6573 = ~n6561 & ~n6572 ;
  assign n6574 = ~n6548 & n6573 ;
  assign n6575 = \s14_msel_arb0_state_reg[0]/NET0131  & ~n6574 ;
  assign n6576 = \s14_msel_arb0_state_reg[0]/NET0131  & n6538 ;
  assign n6577 = n6553 & n6576 ;
  assign n6578 = n6553 & ~n6556 ;
  assign n6579 = ~n6564 & n6578 ;
  assign n6580 = ~n6577 & ~n6579 ;
  assign n6581 = ~n6550 & n6580 ;
  assign n6582 = n6570 & ~n6581 ;
  assign n6583 = n6536 & n6549 ;
  assign n6584 = n6551 & ~n6555 ;
  assign n6585 = n6538 & n6549 ;
  assign n6586 = ~n6584 & n6585 ;
  assign n6587 = ~n6583 & ~n6586 ;
  assign n6588 = n2973 & n6562 ;
  assign n6589 = ~n2929 & ~n2934 ;
  assign n6590 = ~\s14_msel_arb0_state_reg[0]/NET0131  & ~n2932 ;
  assign n6591 = n6589 & ~n6590 ;
  assign n6592 = ~n6544 & ~n6591 ;
  assign n6593 = ~n2939 & ~n2950 ;
  assign n6594 = n2973 & n6593 ;
  assign n6595 = ~n6592 & n6594 ;
  assign n6596 = ~n6588 & ~n6595 ;
  assign n6597 = n6587 & n6596 ;
  assign n6598 = ~n6582 & n6597 ;
  assign n6599 = ~\s14_msel_arb0_state_reg[0]/NET0131  & ~n6598 ;
  assign n6600 = \s14_msel_arb0_state_reg[0]/NET0131  & n6593 ;
  assign n6601 = n6589 & n6600 ;
  assign n6602 = n2977 & n6601 ;
  assign n6603 = n2944 & n6593 ;
  assign n6604 = n6564 & ~n6603 ;
  assign n6605 = ~\rf_conf14_reg[9]/NET0131  & ~\s14_msel_arb0_state_reg[0]/NET0131  ;
  assign n6606 = n2928 & n6605 ;
  assign n6607 = ~n6556 & ~n6606 ;
  assign n6608 = n2977 & n6607 ;
  assign n6609 = ~n6604 & n6608 ;
  assign n6610 = ~n6602 & ~n6609 ;
  assign n6611 = ~n6599 & n6610 ;
  assign n6612 = ~n6575 & n6611 ;
  assign n6613 = n5036 & ~n5042 ;
  assign n6614 = ~n5033 & n5034 ;
  assign n6615 = ~n5037 & ~n5042 ;
  assign n6616 = ~n6614 & n6615 ;
  assign n6617 = ~n6613 & ~n6616 ;
  assign n6618 = ~n5048 & ~n6617 ;
  assign n6619 = n5047 & ~n5048 ;
  assign n6620 = ~\s14_msel_arb1_state_reg[1]/NET0131  & ~\s14_msel_arb1_state_reg[2]/NET0131  ;
  assign n6621 = ~n5058 & n6620 ;
  assign n6622 = ~n6619 & n6621 ;
  assign n6623 = ~n6618 & n6622 ;
  assign n6624 = n5042 & ~n5047 ;
  assign n6625 = \s14_msel_arb1_state_reg[1]/NET0131  & ~\s14_msel_arb1_state_reg[2]/NET0131  ;
  assign n6626 = n6624 & n6625 ;
  assign n6627 = ~n5037 & ~n6614 ;
  assign n6628 = ~n5033 & ~n5058 ;
  assign n6629 = ~\s14_msel_arb1_state_reg[0]/NET0131  & ~n5048 ;
  assign n6630 = n6628 & ~n6629 ;
  assign n6631 = n6627 & ~n6630 ;
  assign n6632 = ~n5036 & ~n5047 ;
  assign n6633 = n6625 & n6632 ;
  assign n6634 = ~n6631 & n6633 ;
  assign n6635 = ~n6626 & ~n6634 ;
  assign n6636 = ~n5036 & n5040 ;
  assign n6637 = ~n6627 & n6636 ;
  assign n6638 = ~n5048 & ~n6624 ;
  assign n6639 = n6628 & n6636 ;
  assign n6640 = ~n6638 & n6639 ;
  assign n6641 = ~n6637 & ~n6640 ;
  assign n6642 = n6635 & n6641 ;
  assign n6643 = ~n6623 & n6642 ;
  assign n6644 = ~\s14_msel_arb1_state_reg[0]/NET0131  & ~n6643 ;
  assign n6645 = \s14_msel_arb1_state_reg[0]/NET0131  & ~n5058 ;
  assign n6646 = ~n5033 & n6632 ;
  assign n6647 = n6645 & n6646 ;
  assign n6648 = ~\rf_conf14_reg[13]/NET0131  & ~\s14_msel_arb1_state_reg[0]/NET0131  ;
  assign n6649 = n4403 & n6648 ;
  assign n6650 = n5034 & ~n6649 ;
  assign n6651 = n5037 & n6632 ;
  assign n6652 = n6638 & ~n6651 ;
  assign n6653 = ~n5058 & ~n6649 ;
  assign n6654 = ~n6652 & n6653 ;
  assign n6655 = ~n6650 & ~n6654 ;
  assign n6656 = ~n6647 & n6655 ;
  assign n6657 = \s14_msel_arb1_state_reg[1]/NET0131  & \s14_msel_arb1_state_reg[2]/NET0131  ;
  assign n6658 = ~n6656 & n6657 ;
  assign n6659 = \s14_msel_arb1_state_reg[0]/NET0131  & ~\s14_msel_arb1_state_reg[1]/NET0131  ;
  assign n6660 = \s14_msel_arb1_state_reg[2]/NET0131  & n6659 ;
  assign n6661 = n6628 & ~n6638 ;
  assign n6662 = n6627 & ~n6661 ;
  assign n6663 = ~n6647 & n6662 ;
  assign n6664 = n6660 & ~n6663 ;
  assign n6665 = ~n5034 & ~n6645 ;
  assign n6666 = n6646 & ~n6665 ;
  assign n6667 = n6652 & ~n6666 ;
  assign n6668 = \s14_msel_arb1_state_reg[0]/NET0131  & n6620 ;
  assign n6669 = ~n6667 & n6668 ;
  assign n6670 = ~n5036 & ~n6619 ;
  assign n6671 = n6630 & n6670 ;
  assign n6672 = ~n6617 & ~n6671 ;
  assign n6673 = \s14_msel_arb1_state_reg[0]/NET0131  & n6625 ;
  assign n6674 = ~n6672 & n6673 ;
  assign n6675 = ~n6669 & ~n6674 ;
  assign n6676 = ~n6664 & n6675 ;
  assign n6677 = ~n6658 & n6676 ;
  assign n6678 = ~n6644 & n6677 ;
  assign n6679 = \s14_msel_arb2_state_reg[1]/NET0131  & ~\s14_msel_arb2_state_reg[2]/NET0131  ;
  assign n6680 = ~n3928 & n6679 ;
  assign n6681 = ~n3902 & ~n3912 ;
  assign n6682 = ~n3902 & n3913 ;
  assign n6683 = ~n6681 & ~n6682 ;
  assign n6684 = n6680 & n6683 ;
  assign n6685 = ~n3918 & ~n3935 ;
  assign n6686 = ~n3913 & ~n3919 ;
  assign n6687 = n6680 & n6686 ;
  assign n6688 = ~n6685 & n6687 ;
  assign n6689 = ~n6684 & ~n6688 ;
  assign n6690 = ~n3903 & ~n6689 ;
  assign n6691 = n3915 & ~n3916 ;
  assign n6692 = ~n3918 & ~n6691 ;
  assign n6693 = ~n3919 & ~n6692 ;
  assign n6694 = n6681 & ~n6693 ;
  assign n6695 = ~\s14_msel_arb2_state_reg[0]/NET0131  & \s14_msel_arb2_state_reg[2]/NET0131  ;
  assign n6696 = ~\s14_msel_arb2_state_reg[1]/NET0131  & n6695 ;
  assign n6697 = ~n6682 & n6696 ;
  assign n6698 = ~n3903 & n6697 ;
  assign n6699 = ~n6694 & n6698 ;
  assign n6700 = ~n6690 & ~n6699 ;
  assign n6701 = ~\s14_msel_arb2_state_reg[1]/NET0131  & ~\s14_msel_arb2_state_reg[2]/NET0131  ;
  assign n6702 = \rf_conf14_reg[1]/NET0131  & ~\s14_msel_arb2_state_reg[0]/NET0131  ;
  assign n6703 = n2938 & n6702 ;
  assign n6704 = n6701 & ~n6703 ;
  assign n6705 = ~n6692 & n6704 ;
  assign n6706 = ~n3903 & ~n3916 ;
  assign n6707 = n6704 & n6706 ;
  assign n6708 = n6683 & n6707 ;
  assign n6709 = ~n6705 & ~n6708 ;
  assign n6710 = n3915 & n6680 ;
  assign n6711 = ~\s14_msel_arb2_state_reg[1]/NET0131  & n3906 ;
  assign n6712 = n3902 & n6711 ;
  assign n6713 = ~n6710 & ~n6712 ;
  assign n6714 = n6709 & n6713 ;
  assign n6715 = n6700 & n6714 ;
  assign n6716 = \s14_msel_arb2_state_reg[0]/NET0131  & n6701 ;
  assign n6717 = ~n3919 & n6716 ;
  assign n6718 = n6706 & n6717 ;
  assign n6719 = ~n3902 & n6711 ;
  assign n6720 = ~n6718 & ~n6719 ;
  assign n6721 = ~n3912 & n3919 ;
  assign n6722 = ~n3912 & ~n3918 ;
  assign n6723 = ~n6691 & n6722 ;
  assign n6724 = ~n6721 & ~n6723 ;
  assign n6725 = \s14_msel_arb2_state_reg[0]/NET0131  & ~n3919 ;
  assign n6726 = n6706 & n6725 ;
  assign n6727 = ~n6718 & ~n6726 ;
  assign n6728 = ~n6724 & n6727 ;
  assign n6729 = ~n6720 & ~n6728 ;
  assign n6730 = ~n3913 & n6729 ;
  assign n6731 = ~n3919 & n6706 ;
  assign n6732 = ~\s14_msel_arb2_state_reg[0]/NET0131  & ~n3902 ;
  assign n6733 = n6731 & ~n6732 ;
  assign n6734 = ~n6724 & ~n6733 ;
  assign n6735 = ~\s14_msel_arb2_state_reg[0]/NET0131  & n3913 ;
  assign n6736 = n3913 & n6681 ;
  assign n6737 = n6692 & n6736 ;
  assign n6738 = ~n6735 & ~n6737 ;
  assign n6739 = n3942 & n6738 ;
  assign n6740 = ~n6734 & n6739 ;
  assign n6741 = ~n6730 & ~n6740 ;
  assign n6742 = n6715 & n6741 ;
  assign n6743 = ~n4396 & ~n4413 ;
  assign n6744 = n4394 & ~n4396 ;
  assign n6745 = ~n6743 & ~n6744 ;
  assign n6746 = ~n4400 & n4404 ;
  assign n6747 = n4389 & ~n4391 ;
  assign n6748 = ~n4400 & ~n4402 ;
  assign n6749 = ~n6747 & n6748 ;
  assign n6750 = ~n6746 & ~n6749 ;
  assign n6751 = \s14_msel_arb3_state_reg[0]/NET0131  & ~n4404 ;
  assign n6752 = ~n4391 & n6751 ;
  assign n6753 = ~n6744 & ~n6752 ;
  assign n6754 = ~n6750 & n6753 ;
  assign n6755 = ~n6745 & ~n6754 ;
  assign n6756 = n4430 & n6755 ;
  assign n6757 = ~\s14_msel_arb3_state_reg[1]/NET0131  & ~\s14_msel_arb3_state_reg[2]/NET0131  ;
  assign n6758 = n6747 & n6757 ;
  assign n6759 = ~n4394 & n4413 ;
  assign n6760 = n4402 & ~n4404 ;
  assign n6761 = ~n4394 & ~n4400 ;
  assign n6762 = ~n6760 & n6761 ;
  assign n6763 = ~n6759 & ~n6762 ;
  assign n6764 = ~n4391 & ~n4396 ;
  assign n6765 = n6757 & n6764 ;
  assign n6766 = n6763 & n6765 ;
  assign n6767 = ~n6758 & ~n6766 ;
  assign n6768 = n4387 & ~n4413 ;
  assign n6769 = n4400 & n6768 ;
  assign n6770 = ~n4402 & ~n6747 ;
  assign n6771 = ~n4391 & n6744 ;
  assign n6772 = n6770 & ~n6771 ;
  assign n6773 = ~n4404 & n6768 ;
  assign n6774 = ~n6772 & n6773 ;
  assign n6775 = ~n6769 & ~n6774 ;
  assign n6776 = ~\s14_msel_arb3_state_reg[0]/NET0131  & n6775 ;
  assign n6777 = n6767 & n6776 ;
  assign n6778 = ~n6756 & n6777 ;
  assign n6779 = ~n4404 & ~n6772 ;
  assign n6780 = ~n4391 & ~n4404 ;
  assign n6781 = n6743 & n6780 ;
  assign n6782 = ~n4400 & ~n6781 ;
  assign n6783 = ~n6779 & n6782 ;
  assign n6784 = n4387 & ~n6783 ;
  assign n6785 = n4394 & n4430 ;
  assign n6786 = \s14_msel_arb3_state_reg[0]/NET0131  & ~n6785 ;
  assign n6787 = ~n6784 & n6786 ;
  assign n6788 = ~n6778 & ~n6787 ;
  assign n6789 = ~n4389 & n4396 ;
  assign n6790 = ~n4391 & ~n4413 ;
  assign n6791 = n6751 & n6790 ;
  assign n6792 = ~n4389 & ~n6791 ;
  assign n6793 = ~n6763 & n6792 ;
  assign n6794 = ~n6789 & ~n6793 ;
  assign n6795 = \s14_msel_arb3_state_reg[0]/NET0131  & n6757 ;
  assign n6796 = n6794 & n6795 ;
  assign n6797 = ~n4400 & ~n6751 ;
  assign n6798 = ~n4391 & n6743 ;
  assign n6799 = ~n6797 & n6798 ;
  assign n6800 = n6772 & ~n6799 ;
  assign n6801 = \rf_conf14_reg[13]/NET0131  & ~\s14_msel_arb3_state_reg[0]/NET0131  ;
  assign n6802 = n4403 & n6801 ;
  assign n6803 = n4410 & ~n6802 ;
  assign n6804 = ~n6800 & n6803 ;
  assign n6805 = n6751 & n6764 ;
  assign n6806 = ~n6750 & ~n6805 ;
  assign n6807 = \s14_msel_arb3_state_reg[0]/NET0131  & n4430 ;
  assign n6808 = ~n4394 & n6807 ;
  assign n6809 = ~n4413 & n6808 ;
  assign n6810 = ~n6806 & n6809 ;
  assign n6811 = ~n6804 & ~n6810 ;
  assign n6812 = ~n6796 & n6811 ;
  assign n6813 = ~n6788 & n6812 ;
  assign n6814 = ~n3755 & ~n3761 ;
  assign n6815 = n3753 & ~n3761 ;
  assign n6816 = ~n6814 & ~n6815 ;
  assign n6817 = ~n3764 & ~n6816 ;
  assign n6818 = ~n3750 & ~n3753 ;
  assign n6819 = \s15_msel_arb1_state_reg[0]/NET0131  & ~n3766 ;
  assign n6820 = ~n3748 & ~n6819 ;
  assign n6821 = n6818 & ~n6820 ;
  assign n6822 = n6817 & ~n6821 ;
  assign n6823 = n3759 & ~n3764 ;
  assign n6824 = \s15_msel_arb1_state_reg[2]/NET0131  & ~n3839 ;
  assign n6825 = ~n6823 & n6824 ;
  assign n6826 = ~n6822 & n6825 ;
  assign n6827 = ~\s15_msel_arb1_state_reg[1]/NET0131  & n6826 ;
  assign n6828 = ~\s15_msel_arb1_state_reg[2]/NET0131  & n3755 ;
  assign n6829 = n3764 & ~n3766 ;
  assign n6830 = ~n3748 & ~n6829 ;
  assign n6831 = ~\s15_msel_arb1_state_reg[0]/NET0131  & ~n3761 ;
  assign n6832 = ~n3759 & ~n3766 ;
  assign n6833 = ~n6831 & n6832 ;
  assign n6834 = n6830 & ~n6833 ;
  assign n6835 = ~\s15_msel_arb1_state_reg[2]/NET0131  & ~n3750 ;
  assign n6836 = ~n6834 & n6835 ;
  assign n6837 = ~n6828 & ~n6836 ;
  assign n6838 = ~\s15_msel_arb1_state_reg[0]/NET0131  & n3753 ;
  assign n6839 = n3753 & n6814 ;
  assign n6840 = n6830 & n6839 ;
  assign n6841 = ~n6838 & ~n6840 ;
  assign n6842 = ~\s15_msel_arb1_state_reg[1]/NET0131  & n6841 ;
  assign n6843 = ~n6837 & n6842 ;
  assign n6844 = ~n6827 & ~n6843 ;
  assign n6845 = ~n3766 & ~n6823 ;
  assign n6846 = ~n3748 & ~n6845 ;
  assign n6847 = ~n3748 & ~n3764 ;
  assign n6848 = ~n6816 & n6847 ;
  assign n6849 = ~n6846 & ~n6848 ;
  assign n6850 = ~\rf_conf15_reg[5]/NET0131  & ~\s15_msel_arb1_state_reg[0]/NET0131  ;
  assign n6851 = n3749 & n6850 ;
  assign n6852 = ~\s15_msel_arb1_state_reg[2]/NET0131  & ~n6851 ;
  assign n6853 = n6849 & n6852 ;
  assign n6854 = ~\rf_conf15_reg[13]/NET0131  & ~\s15_msel_arb1_state_reg[0]/NET0131  ;
  assign n6855 = n3758 & n6854 ;
  assign n6856 = \s15_msel_arb1_state_reg[2]/NET0131  & ~n6855 ;
  assign n6857 = n6816 & n6856 ;
  assign n6858 = n6818 & n6856 ;
  assign n6859 = ~n6830 & n6858 ;
  assign n6860 = ~n6857 & ~n6859 ;
  assign n6861 = ~n3759 & n6818 ;
  assign n6862 = n6819 & n6861 ;
  assign n6863 = n6860 & ~n6862 ;
  assign n6864 = ~n6853 & n6863 ;
  assign n6865 = \s15_msel_arb1_state_reg[1]/NET0131  & ~n6864 ;
  assign n6866 = n6844 & ~n6865 ;
  assign n6867 = ~n3773 & n3774 ;
  assign n6868 = ~n3780 & ~n6867 ;
  assign n6869 = \s15_msel_arb2_state_reg[2]/NET0131  & ~n6868 ;
  assign n6870 = ~n3777 & n3778 ;
  assign n6871 = ~n3770 & ~n6870 ;
  assign n6872 = ~n3771 & ~n3773 ;
  assign n6873 = \s15_msel_arb2_state_reg[2]/NET0131  & n6872 ;
  assign n6874 = ~n6871 & n6873 ;
  assign n6875 = ~n6869 & ~n6874 ;
  assign n6876 = ~n3781 & ~n6875 ;
  assign n6877 = ~\s15_msel_arb2_state_reg[2]/NET0131  & ~n6871 ;
  assign n6878 = ~n3777 & ~n3781 ;
  assign n6879 = ~\s15_msel_arb2_state_reg[2]/NET0131  & n6878 ;
  assign n6880 = ~n6868 & n6879 ;
  assign n6881 = ~n6877 & ~n6880 ;
  assign n6882 = ~n3771 & ~n6881 ;
  assign n6883 = ~\s15_msel_arb2_state_reg[0]/NET0131  & ~n6882 ;
  assign n6884 = ~n6876 & n6883 ;
  assign n6885 = n6872 & n6878 ;
  assign n6886 = \s15_msel_arb2_state_reg[0]/NET0131  & ~n6885 ;
  assign n6887 = n6875 & n6886 ;
  assign n6888 = n6881 & n6887 ;
  assign n6889 = \s15_msel_arb2_state_reg[1]/NET0131  & ~n6888 ;
  assign n6890 = ~n6884 & n6889 ;
  assign n6891 = n3780 & n6878 ;
  assign n6892 = n6871 & ~n6891 ;
  assign n6893 = \s15_msel_arb2_state_reg[0]/NET0131  & n6878 ;
  assign n6894 = n6892 & ~n6893 ;
  assign n6895 = ~n3770 & n3773 ;
  assign n6896 = ~n6870 & n6895 ;
  assign n6897 = ~n6891 & n6896 ;
  assign n6898 = ~n3771 & ~n3774 ;
  assign n6899 = ~\s15_msel_arb2_state_reg[2]/NET0131  & n6898 ;
  assign n6900 = ~n6897 & n6899 ;
  assign n6901 = ~n6894 & n6900 ;
  assign n6902 = ~\s15_msel_arb2_state_reg[2]/NET0131  & ~n3774 ;
  assign n6903 = \s15_msel_arb2_state_reg[2]/NET0131  & ~n3778 ;
  assign n6904 = ~n6902 & ~n6903 ;
  assign n6905 = ~n3778 & ~n3781 ;
  assign n6906 = \s15_msel_arb2_state_reg[2]/NET0131  & n6905 ;
  assign n6907 = ~n6904 & ~n6906 ;
  assign n6908 = n3770 & n6872 ;
  assign n6909 = n6868 & ~n6908 ;
  assign n6910 = \s15_msel_arb2_state_reg[0]/NET0131  & ~n3777 ;
  assign n6911 = n6872 & n6910 ;
  assign n6912 = ~n6904 & ~n6911 ;
  assign n6913 = n6909 & n6912 ;
  assign n6914 = ~n6907 & ~n6913 ;
  assign n6915 = ~n6901 & ~n6914 ;
  assign n6916 = \s15_msel_arb2_state_reg[0]/NET0131  & ~\s15_msel_arb2_state_reg[1]/NET0131  ;
  assign n6917 = ~n6915 & n6916 ;
  assign n6918 = ~\s15_msel_arb2_state_reg[0]/NET0131  & ~\s15_msel_arb2_state_reg[1]/NET0131  ;
  assign n6919 = \s15_msel_arb2_state_reg[2]/NET0131  & n6918 ;
  assign n6920 = \rf_conf15_reg[9]/NET0131  & ~\s15_msel_arb2_state_reg[0]/NET0131  ;
  assign n6921 = n2990 & n6920 ;
  assign n6922 = ~n3779 & ~n6921 ;
  assign n6923 = ~n6878 & ~n6922 ;
  assign n6924 = \s15_msel_arb2_state_reg[0]/NET0131  & n6872 ;
  assign n6925 = ~n6922 & ~n6924 ;
  assign n6926 = n6909 & n6925 ;
  assign n6927 = ~n6923 & ~n6926 ;
  assign n6928 = n6919 & n6927 ;
  assign n6929 = \rf_conf15_reg[1]/NET0131  & ~\s15_msel_arb2_state_reg[0]/NET0131  ;
  assign n6930 = n3009 & n6929 ;
  assign n6931 = ~n3775 & ~n6930 ;
  assign n6932 = ~n6872 & ~n6931 ;
  assign n6933 = ~n6893 & ~n6931 ;
  assign n6934 = n6892 & n6933 ;
  assign n6935 = ~n6932 & ~n6934 ;
  assign n6936 = ~\s15_msel_arb2_state_reg[2]/NET0131  & n6918 ;
  assign n6937 = n6935 & n6936 ;
  assign n6938 = ~n6928 & ~n6937 ;
  assign n6939 = ~n6917 & n6938 ;
  assign n6940 = ~n6890 & n6939 ;
  assign n6941 = \rf_conf15_reg[13]/NET0131  & ~\s15_msel_arb2_state_reg[0]/NET0131  ;
  assign n6942 = n2993 & n6941 ;
  assign n6943 = ~n3780 & ~n6942 ;
  assign n6944 = ~n6918 & ~n6943 ;
  assign n6945 = ~\s15_msel_arb2_state_reg[1]/NET0131  & ~n6918 ;
  assign n6946 = ~n6905 & n6945 ;
  assign n6947 = ~n6944 & ~n6946 ;
  assign n6948 = ~n3776 & n6947 ;
  assign n6949 = \s15_msel_arb2_state_reg[2]/NET0131  & ~n6948 ;
  assign n6950 = ~\s15_msel_arb2_state_reg[2]/NET0131  & ~n3770 ;
  assign n6951 = ~n6919 & ~n6950 ;
  assign n6952 = n6898 & ~n6930 ;
  assign n6953 = \rf_conf15_reg[5]/NET0131  & ~\s15_msel_arb2_state_reg[0]/NET0131  ;
  assign n6954 = n3003 & n6953 ;
  assign n6955 = \s15_msel_arb2_state_reg[1]/NET0131  & ~n6954 ;
  assign n6956 = ~n6919 & ~n6955 ;
  assign n6957 = ~n6952 & n6956 ;
  assign n6958 = ~n6951 & ~n6957 ;
  assign n6959 = ~n3783 & n6958 ;
  assign n6960 = ~n6949 & ~n6959 ;
  assign n6961 = n3791 & ~n3795 ;
  assign n6962 = n3788 & ~n3789 ;
  assign n6963 = ~n3792 & ~n3795 ;
  assign n6964 = ~n6962 & n6963 ;
  assign n6965 = ~n6961 & ~n6964 ;
  assign n6966 = ~n3799 & ~n6965 ;
  assign n6967 = n3796 & ~n3799 ;
  assign n6968 = \s15_msel_arb3_state_reg[2]/NET0131  & ~n6967 ;
  assign n6969 = ~n3798 & n6968 ;
  assign n6970 = ~n6966 & n6969 ;
  assign n6971 = ~\s15_msel_arb3_state_reg[1]/NET0131  & n6970 ;
  assign n6972 = ~n6966 & n6968 ;
  assign n6973 = ~n3792 & ~n6962 ;
  assign n6974 = ~\s15_msel_arb3_state_reg[2]/NET0131  & ~n6973 ;
  assign n6975 = ~n3795 & ~n3799 ;
  assign n6976 = ~n6967 & ~n6975 ;
  assign n6977 = ~n3789 & ~n3798 ;
  assign n6978 = ~\s15_msel_arb3_state_reg[2]/NET0131  & n6977 ;
  assign n6979 = n6976 & n6978 ;
  assign n6980 = ~n6974 & ~n6979 ;
  assign n6981 = ~n3791 & ~n3796 ;
  assign n6982 = \s15_msel_arb3_state_reg[0]/NET0131  & n6981 ;
  assign n6983 = n6977 & n6982 ;
  assign n6984 = n6980 & ~n6983 ;
  assign n6985 = ~n6972 & n6984 ;
  assign n6986 = \s15_msel_arb3_state_reg[0]/NET0131  & ~\s15_msel_arb3_state_reg[1]/NET0131  ;
  assign n6987 = ~n6985 & n6986 ;
  assign n6988 = ~n6971 & ~n6987 ;
  assign n6989 = ~\s15_msel_arb3_state_reg[1]/NET0131  & ~n3791 ;
  assign n6990 = ~n6980 & n6989 ;
  assign n6991 = ~\s15_msel_arb3_state_reg[0]/NET0131  & n6990 ;
  assign n6992 = n3792 & n6981 ;
  assign n6993 = ~n6976 & ~n6992 ;
  assign n6994 = ~n6982 & n6993 ;
  assign n6995 = n6977 & ~n6994 ;
  assign n6996 = \rf_conf15_reg[5]/NET0131  & ~\s15_msel_arb3_state_reg[0]/NET0131  ;
  assign n6997 = n3749 & n6996 ;
  assign n6998 = ~n3790 & ~n6997 ;
  assign n6999 = ~\s15_msel_arb3_state_reg[2]/NET0131  & ~n6998 ;
  assign n7000 = ~n6995 & n6999 ;
  assign n7001 = \rf_conf15_reg[13]/NET0131  & ~\s15_msel_arb3_state_reg[0]/NET0131  ;
  assign n7002 = n3758 & n7001 ;
  assign n7003 = ~n3797 & ~n7002 ;
  assign n7004 = \s15_msel_arb3_state_reg[2]/NET0131  & ~n7003 ;
  assign n7005 = \s15_msel_arb3_state_reg[1]/NET0131  & ~n7004 ;
  assign n7006 = ~\s15_msel_arb3_state_reg[0]/NET0131  & ~n3799 ;
  assign n7007 = n6977 & ~n7006 ;
  assign n7008 = n6973 & ~n7007 ;
  assign n7009 = \s15_msel_arb3_state_reg[1]/NET0131  & n6981 ;
  assign n7010 = ~n7008 & n7009 ;
  assign n7011 = ~n7005 & ~n7010 ;
  assign n7012 = ~\s15_msel_arb3_state_reg[0]/NET0131  & ~n7011 ;
  assign n7013 = ~n7000 & n7012 ;
  assign n7014 = ~n6991 & ~n7013 ;
  assign n7015 = ~n3791 & ~n6967 ;
  assign n7016 = n7007 & n7015 ;
  assign n7017 = \s15_msel_arb3_state_reg[2]/NET0131  & ~n7016 ;
  assign n7018 = ~n6965 & n7017 ;
  assign n7019 = ~n3798 & ~n6993 ;
  assign n7020 = n3814 & ~n6983 ;
  assign n7021 = ~n7019 & n7020 ;
  assign n7022 = n3812 & ~n7021 ;
  assign n7023 = ~n7018 & n7022 ;
  assign n7024 = n7014 & ~n7023 ;
  assign n7025 = n6988 & n7024 ;
  assign n7026 = ~n3380 & n3389 ;
  assign n7027 = n3370 & ~n3372 ;
  assign n7028 = ~n3380 & ~n3387 ;
  assign n7029 = ~n7027 & n7028 ;
  assign n7030 = ~n7026 & ~n7029 ;
  assign n7031 = ~n3372 & ~n3389 ;
  assign n7032 = ~n3375 & n7031 ;
  assign n7033 = ~n3377 & n3382 ;
  assign n7034 = ~\s1_msel_arb0_state_reg[0]/NET0131  & ~n3377 ;
  assign n7035 = ~n7033 & ~n7034 ;
  assign n7036 = n7032 & n7035 ;
  assign n7037 = ~n7030 & ~n7036 ;
  assign n7038 = n3423 & ~n7037 ;
  assign n7039 = ~n3377 & ~n3380 ;
  assign n7040 = ~n7033 & ~n7039 ;
  assign n7041 = ~\s1_msel_arb0_state_reg[1]/NET0131  & \s1_msel_arb0_state_reg[2]/NET0131  ;
  assign n7042 = ~\rf_conf1_reg[3]/NET0131  & ~\s1_msel_arb0_state_reg[1]/NET0131  ;
  assign n7043 = n3386 & n7042 ;
  assign n7044 = ~n7041 & ~n7043 ;
  assign n7045 = n7040 & ~n7044 ;
  assign n7046 = ~n3370 & n3375 ;
  assign n7047 = ~n3372 & ~n7046 ;
  assign n7048 = ~n3387 & ~n7047 ;
  assign n7049 = ~n3382 & ~n3389 ;
  assign n7050 = \s1_msel_arb0_state_reg[2]/NET0131  & ~n7049 ;
  assign n7051 = ~n7044 & ~n7050 ;
  assign n7052 = ~n7048 & n7051 ;
  assign n7053 = ~n7045 & ~n7052 ;
  assign n7054 = ~n7038 & n7053 ;
  assign n7055 = \s1_msel_arb0_state_reg[0]/NET0131  & ~n7054 ;
  assign n7056 = \s1_msel_arb0_state_reg[0]/NET0131  & n7049 ;
  assign n7057 = ~n3372 & ~n3375 ;
  assign n7058 = n7056 & n7057 ;
  assign n7059 = n3417 & n7058 ;
  assign n7060 = n3387 & n7049 ;
  assign n7061 = ~n3370 & ~n7040 ;
  assign n7062 = ~n7060 & n7061 ;
  assign n7063 = ~\rf_conf1_reg[5]/NET0131  & ~\s1_msel_arb0_state_reg[0]/NET0131  ;
  assign n7064 = n3371 & n7063 ;
  assign n7065 = ~n7046 & ~n7064 ;
  assign n7066 = n3417 & n7065 ;
  assign n7067 = ~n7062 & n7066 ;
  assign n7068 = ~n7059 & ~n7067 ;
  assign n7069 = ~n3387 & ~n7027 ;
  assign n7070 = ~n3389 & ~n7069 ;
  assign n7071 = ~n3375 & ~n3382 ;
  assign n7072 = \s1_msel_arb0_state_reg[2]/NET0131  & ~n7071 ;
  assign n7073 = n7070 & ~n7072 ;
  assign n7074 = ~\s1_msel_arb0_state_reg[2]/NET0131  & ~n7031 ;
  assign n7075 = ~n3375 & n7040 ;
  assign n7076 = ~n7074 & n7075 ;
  assign n7077 = ~n7073 & ~n7076 ;
  assign n7078 = ~\s1_msel_arb0_state_reg[0]/NET0131  & ~\s1_msel_arb0_state_reg[1]/NET0131  ;
  assign n7079 = ~n7077 & n7078 ;
  assign n7080 = ~n7056 & n7061 ;
  assign n7081 = ~\s1_msel_arb0_state_reg[1]/NET0131  & ~\s1_msel_arb0_state_reg[2]/NET0131  ;
  assign n7082 = \s1_msel_arb0_state_reg[0]/NET0131  & n7081 ;
  assign n7083 = ~n3387 & n7082 ;
  assign n7084 = n7047 & n7083 ;
  assign n7085 = ~n7080 & n7084 ;
  assign n7086 = n7032 & ~n7034 ;
  assign n7087 = ~n7030 & ~n7086 ;
  assign n7088 = \s1_msel_arb0_state_reg[2]/NET0131  & n3406 ;
  assign n7089 = ~n3382 & n7088 ;
  assign n7090 = ~n7087 & n7089 ;
  assign n7091 = ~n7085 & ~n7090 ;
  assign n7092 = ~n7079 & n7091 ;
  assign n7093 = n7068 & n7092 ;
  assign n7094 = ~n7055 & n7093 ;
  assign n7095 = n5075 & ~n5081 ;
  assign n7096 = ~n5072 & n5073 ;
  assign n7097 = ~n5076 & ~n5081 ;
  assign n7098 = ~n7096 & n7097 ;
  assign n7099 = ~n7095 & ~n7098 ;
  assign n7100 = ~n5087 & ~n7099 ;
  assign n7101 = n5086 & ~n5087 ;
  assign n7102 = ~\s1_msel_arb1_state_reg[1]/NET0131  & ~\s1_msel_arb1_state_reg[2]/NET0131  ;
  assign n7103 = ~n5097 & n7102 ;
  assign n7104 = ~n7101 & n7103 ;
  assign n7105 = ~n7100 & n7104 ;
  assign n7106 = n5081 & ~n5086 ;
  assign n7107 = \s1_msel_arb1_state_reg[1]/NET0131  & ~\s1_msel_arb1_state_reg[2]/NET0131  ;
  assign n7108 = n7106 & n7107 ;
  assign n7109 = ~n5076 & ~n7096 ;
  assign n7110 = ~n5072 & ~n5097 ;
  assign n7111 = ~\s1_msel_arb1_state_reg[0]/NET0131  & ~n5087 ;
  assign n7112 = n7110 & ~n7111 ;
  assign n7113 = n7109 & ~n7112 ;
  assign n7114 = ~n5075 & ~n5086 ;
  assign n7115 = n7107 & n7114 ;
  assign n7116 = ~n7113 & n7115 ;
  assign n7117 = ~n7108 & ~n7116 ;
  assign n7118 = ~n5075 & n5079 ;
  assign n7119 = ~n7109 & n7118 ;
  assign n7120 = ~n5087 & ~n7106 ;
  assign n7121 = n7110 & n7118 ;
  assign n7122 = ~n7120 & n7121 ;
  assign n7123 = ~n7119 & ~n7122 ;
  assign n7124 = n7117 & n7123 ;
  assign n7125 = ~n7105 & n7124 ;
  assign n7126 = ~\s1_msel_arb1_state_reg[0]/NET0131  & ~n7125 ;
  assign n7127 = \s1_msel_arb1_state_reg[0]/NET0131  & ~n5097 ;
  assign n7128 = ~n5072 & n7114 ;
  assign n7129 = n7127 & n7128 ;
  assign n7130 = ~\rf_conf1_reg[13]/NET0131  & ~\s1_msel_arb1_state_reg[0]/NET0131  ;
  assign n7131 = n4489 & n7130 ;
  assign n7132 = n5073 & ~n7131 ;
  assign n7133 = n5076 & n7114 ;
  assign n7134 = n7120 & ~n7133 ;
  assign n7135 = ~n5097 & ~n7131 ;
  assign n7136 = ~n7134 & n7135 ;
  assign n7137 = ~n7132 & ~n7136 ;
  assign n7138 = ~n7129 & n7137 ;
  assign n7139 = \s1_msel_arb1_state_reg[1]/NET0131  & \s1_msel_arb1_state_reg[2]/NET0131  ;
  assign n7140 = ~n7138 & n7139 ;
  assign n7141 = \s1_msel_arb1_state_reg[0]/NET0131  & ~\s1_msel_arb1_state_reg[1]/NET0131  ;
  assign n7142 = \s1_msel_arb1_state_reg[2]/NET0131  & n7141 ;
  assign n7143 = n7110 & ~n7120 ;
  assign n7144 = n7109 & ~n7143 ;
  assign n7145 = ~n7129 & n7144 ;
  assign n7146 = n7142 & ~n7145 ;
  assign n7147 = ~n5073 & ~n7127 ;
  assign n7148 = n7128 & ~n7147 ;
  assign n7149 = n7134 & ~n7148 ;
  assign n7150 = \s1_msel_arb1_state_reg[0]/NET0131  & n7102 ;
  assign n7151 = ~n7149 & n7150 ;
  assign n7152 = ~n5075 & ~n7101 ;
  assign n7153 = n7112 & n7152 ;
  assign n7154 = ~n7099 & ~n7153 ;
  assign n7155 = \s1_msel_arb1_state_reg[0]/NET0131  & n7107 ;
  assign n7156 = ~n7154 & n7155 ;
  assign n7157 = ~n7151 & ~n7156 ;
  assign n7158 = ~n7146 & n7157 ;
  assign n7159 = ~n7140 & n7158 ;
  assign n7160 = ~n7126 & n7159 ;
  assign n7161 = ~\s1_msel_arb2_state_reg[1]/NET0131  & \s1_msel_arb2_state_reg[2]/NET0131  ;
  assign n7162 = ~n4439 & n7161 ;
  assign n7163 = n4438 & n7162 ;
  assign n7164 = ~n4442 & n4459 ;
  assign n7165 = n4445 & ~n4448 ;
  assign n7166 = ~n4442 & ~n4453 ;
  assign n7167 = ~n7165 & n7166 ;
  assign n7168 = ~n7164 & ~n7167 ;
  assign n7169 = ~n4441 & n7162 ;
  assign n7170 = n7168 & n7169 ;
  assign n7171 = ~n7163 & ~n7170 ;
  assign n7172 = ~\s1_msel_arb2_state_reg[0]/NET0131  & ~n7171 ;
  assign n7173 = ~n4439 & ~n4448 ;
  assign n7174 = ~n7165 & ~n7173 ;
  assign n7175 = ~n4441 & n4442 ;
  assign n7176 = ~n4438 & ~n7175 ;
  assign n7177 = ~n4441 & ~n4459 ;
  assign n7178 = n4453 & n7177 ;
  assign n7179 = n7176 & ~n7178 ;
  assign n7180 = \s1_msel_arb2_state_reg[0]/NET0131  & n7177 ;
  assign n7181 = ~n7165 & ~n7180 ;
  assign n7182 = n7179 & n7181 ;
  assign n7183 = ~n7174 & ~n7182 ;
  assign n7184 = \s1_msel_arb2_state_reg[1]/NET0131  & ~\s1_msel_arb2_state_reg[2]/NET0131  ;
  assign n7185 = ~\s1_msel_arb2_state_reg[0]/NET0131  & n7184 ;
  assign n7186 = n7183 & n7185 ;
  assign n7187 = ~n7172 & ~n7186 ;
  assign n7188 = \s1_msel_arb2_state_reg[0]/NET0131  & ~n4441 ;
  assign n7189 = ~n4438 & ~n7188 ;
  assign n7190 = ~n4459 & n7173 ;
  assign n7191 = ~n7189 & n7190 ;
  assign n7192 = ~n7168 & ~n7191 ;
  assign n7193 = \rf_conf1_reg[13]/NET0131  & ~\s1_msel_arb2_state_reg[0]/NET0131  ;
  assign n7194 = n3381 & n7193 ;
  assign n7195 = \s1_msel_arb2_state_reg[1]/NET0131  & \s1_msel_arb2_state_reg[2]/NET0131  ;
  assign n7196 = ~n7194 & n7195 ;
  assign n7197 = ~n7192 & n7196 ;
  assign n7198 = ~n4439 & ~n7179 ;
  assign n7199 = n7173 & n7180 ;
  assign n7200 = ~n4445 & ~n7199 ;
  assign n7201 = ~n7198 & n7200 ;
  assign n7202 = \s1_msel_arb2_state_reg[0]/NET0131  & n7184 ;
  assign n7203 = ~n7201 & n7202 ;
  assign n7204 = ~n7197 & ~n7203 ;
  assign n7205 = \s1_msel_arb2_state_reg[0]/NET0131  & ~\s1_msel_arb2_state_reg[1]/NET0131  ;
  assign n7206 = \s1_msel_arb2_state_reg[2]/NET0131  & n7205 ;
  assign n7207 = ~n4441 & n7168 ;
  assign n7208 = ~n4438 & ~n7199 ;
  assign n7209 = ~n7207 & n7208 ;
  assign n7210 = n7206 & ~n7209 ;
  assign n7211 = ~n4453 & ~n7165 ;
  assign n7212 = \rf_conf1_reg[1]/NET0131  & ~\s1_msel_arb2_state_reg[0]/NET0131  ;
  assign n7213 = n3388 & n7212 ;
  assign n7214 = ~n7211 & ~n7213 ;
  assign n7215 = n7173 & ~n7213 ;
  assign n7216 = ~n7176 & n7215 ;
  assign n7217 = ~n7214 & ~n7216 ;
  assign n7218 = ~n7199 & n7217 ;
  assign n7219 = ~\s1_msel_arb2_state_reg[1]/NET0131  & ~\s1_msel_arb2_state_reg[2]/NET0131  ;
  assign n7220 = ~n7218 & n7219 ;
  assign n7221 = ~n7210 & ~n7220 ;
  assign n7222 = n7204 & n7221 ;
  assign n7223 = n7187 & n7222 ;
  assign n7224 = ~n4482 & ~n4499 ;
  assign n7225 = n4480 & ~n4482 ;
  assign n7226 = ~n7224 & ~n7225 ;
  assign n7227 = ~n4486 & n4490 ;
  assign n7228 = n4475 & ~n4477 ;
  assign n7229 = ~n4486 & ~n4488 ;
  assign n7230 = ~n7228 & n7229 ;
  assign n7231 = ~n7227 & ~n7230 ;
  assign n7232 = \s1_msel_arb3_state_reg[0]/NET0131  & ~n4490 ;
  assign n7233 = ~n4477 & n7232 ;
  assign n7234 = ~n7225 & ~n7233 ;
  assign n7235 = ~n7231 & n7234 ;
  assign n7236 = ~n7226 & ~n7235 ;
  assign n7237 = n4516 & n7236 ;
  assign n7238 = ~\s1_msel_arb3_state_reg[1]/NET0131  & ~\s1_msel_arb3_state_reg[2]/NET0131  ;
  assign n7239 = n7228 & n7238 ;
  assign n7240 = ~n4480 & n4499 ;
  assign n7241 = n4488 & ~n4490 ;
  assign n7242 = ~n4480 & ~n4486 ;
  assign n7243 = ~n7241 & n7242 ;
  assign n7244 = ~n7240 & ~n7243 ;
  assign n7245 = ~n4477 & ~n4482 ;
  assign n7246 = n7238 & n7245 ;
  assign n7247 = n7244 & n7246 ;
  assign n7248 = ~n7239 & ~n7247 ;
  assign n7249 = n4473 & ~n4499 ;
  assign n7250 = n4486 & n7249 ;
  assign n7251 = ~n4488 & ~n7228 ;
  assign n7252 = ~n4477 & n7225 ;
  assign n7253 = n7251 & ~n7252 ;
  assign n7254 = ~n4490 & n7249 ;
  assign n7255 = ~n7253 & n7254 ;
  assign n7256 = ~n7250 & ~n7255 ;
  assign n7257 = ~\s1_msel_arb3_state_reg[0]/NET0131  & n7256 ;
  assign n7258 = n7248 & n7257 ;
  assign n7259 = ~n7237 & n7258 ;
  assign n7260 = ~n4490 & ~n7253 ;
  assign n7261 = ~n4477 & ~n4490 ;
  assign n7262 = n7224 & n7261 ;
  assign n7263 = ~n4486 & ~n7262 ;
  assign n7264 = ~n7260 & n7263 ;
  assign n7265 = n4473 & ~n7264 ;
  assign n7266 = n4480 & n4516 ;
  assign n7267 = \s1_msel_arb3_state_reg[0]/NET0131  & ~n7266 ;
  assign n7268 = ~n7265 & n7267 ;
  assign n7269 = ~n7259 & ~n7268 ;
  assign n7270 = ~n4475 & n4482 ;
  assign n7271 = ~n4477 & ~n4499 ;
  assign n7272 = n7232 & n7271 ;
  assign n7273 = ~n4475 & ~n7272 ;
  assign n7274 = ~n7244 & n7273 ;
  assign n7275 = ~n7270 & ~n7274 ;
  assign n7276 = \s1_msel_arb3_state_reg[0]/NET0131  & n7238 ;
  assign n7277 = n7275 & n7276 ;
  assign n7278 = ~n4486 & ~n7232 ;
  assign n7279 = ~n4477 & n7224 ;
  assign n7280 = ~n7278 & n7279 ;
  assign n7281 = n7253 & ~n7280 ;
  assign n7282 = \rf_conf1_reg[13]/NET0131  & ~\s1_msel_arb3_state_reg[0]/NET0131  ;
  assign n7283 = n4489 & n7282 ;
  assign n7284 = n4496 & ~n7283 ;
  assign n7285 = ~n7281 & n7284 ;
  assign n7286 = n7232 & n7245 ;
  assign n7287 = ~n7231 & ~n7286 ;
  assign n7288 = \s1_msel_arb3_state_reg[0]/NET0131  & n4516 ;
  assign n7289 = ~n4480 & n7288 ;
  assign n7290 = ~n4499 & n7289 ;
  assign n7291 = ~n7287 & n7290 ;
  assign n7292 = ~n7285 & ~n7291 ;
  assign n7293 = ~n7277 & n7292 ;
  assign n7294 = ~n7269 & n7293 ;
  assign n7295 = ~n3443 & n3452 ;
  assign n7296 = n3433 & ~n3435 ;
  assign n7297 = ~n3443 & ~n3450 ;
  assign n7298 = ~n7296 & n7297 ;
  assign n7299 = ~n7295 & ~n7298 ;
  assign n7300 = ~n3435 & ~n3452 ;
  assign n7301 = ~n3438 & n7300 ;
  assign n7302 = ~n3440 & n3445 ;
  assign n7303 = ~\s2_msel_arb0_state_reg[0]/NET0131  & ~n3440 ;
  assign n7304 = ~n7302 & ~n7303 ;
  assign n7305 = n7301 & n7304 ;
  assign n7306 = ~n7299 & ~n7305 ;
  assign n7307 = n3486 & ~n7306 ;
  assign n7308 = ~n3440 & ~n3443 ;
  assign n7309 = ~n7302 & ~n7308 ;
  assign n7310 = ~\s2_msel_arb0_state_reg[1]/NET0131  & \s2_msel_arb0_state_reg[2]/NET0131  ;
  assign n7311 = ~\rf_conf2_reg[3]/NET0131  & ~\s2_msel_arb0_state_reg[1]/NET0131  ;
  assign n7312 = n3449 & n7311 ;
  assign n7313 = ~n7310 & ~n7312 ;
  assign n7314 = n7309 & ~n7313 ;
  assign n7315 = ~n3433 & n3438 ;
  assign n7316 = ~n3435 & ~n7315 ;
  assign n7317 = ~n3450 & ~n7316 ;
  assign n7318 = ~n3445 & ~n3452 ;
  assign n7319 = \s2_msel_arb0_state_reg[2]/NET0131  & ~n7318 ;
  assign n7320 = ~n7313 & ~n7319 ;
  assign n7321 = ~n7317 & n7320 ;
  assign n7322 = ~n7314 & ~n7321 ;
  assign n7323 = ~n7307 & n7322 ;
  assign n7324 = \s2_msel_arb0_state_reg[0]/NET0131  & ~n7323 ;
  assign n7325 = \s2_msel_arb0_state_reg[0]/NET0131  & n7318 ;
  assign n7326 = ~n3435 & ~n3438 ;
  assign n7327 = n7325 & n7326 ;
  assign n7328 = n3480 & n7327 ;
  assign n7329 = n3450 & n7318 ;
  assign n7330 = ~n3433 & ~n7309 ;
  assign n7331 = ~n7329 & n7330 ;
  assign n7332 = ~\rf_conf2_reg[5]/NET0131  & ~\s2_msel_arb0_state_reg[0]/NET0131  ;
  assign n7333 = n3434 & n7332 ;
  assign n7334 = ~n7315 & ~n7333 ;
  assign n7335 = n3480 & n7334 ;
  assign n7336 = ~n7331 & n7335 ;
  assign n7337 = ~n7328 & ~n7336 ;
  assign n7338 = ~n3450 & ~n7296 ;
  assign n7339 = ~n3452 & ~n7338 ;
  assign n7340 = ~n3438 & ~n3445 ;
  assign n7341 = \s2_msel_arb0_state_reg[2]/NET0131  & ~n7340 ;
  assign n7342 = n7339 & ~n7341 ;
  assign n7343 = ~\s2_msel_arb0_state_reg[2]/NET0131  & ~n7300 ;
  assign n7344 = ~n3438 & n7309 ;
  assign n7345 = ~n7343 & n7344 ;
  assign n7346 = ~n7342 & ~n7345 ;
  assign n7347 = ~\s2_msel_arb0_state_reg[0]/NET0131  & ~\s2_msel_arb0_state_reg[1]/NET0131  ;
  assign n7348 = ~n7346 & n7347 ;
  assign n7349 = ~n7325 & n7330 ;
  assign n7350 = ~\s2_msel_arb0_state_reg[1]/NET0131  & ~\s2_msel_arb0_state_reg[2]/NET0131  ;
  assign n7351 = \s2_msel_arb0_state_reg[0]/NET0131  & n7350 ;
  assign n7352 = ~n3450 & n7351 ;
  assign n7353 = n7316 & n7352 ;
  assign n7354 = ~n7349 & n7353 ;
  assign n7355 = n7301 & ~n7303 ;
  assign n7356 = ~n7299 & ~n7355 ;
  assign n7357 = \s2_msel_arb0_state_reg[2]/NET0131  & n3469 ;
  assign n7358 = ~n3445 & n7357 ;
  assign n7359 = ~n7356 & n7358 ;
  assign n7360 = ~n7354 & ~n7359 ;
  assign n7361 = ~n7348 & n7360 ;
  assign n7362 = n7337 & n7361 ;
  assign n7363 = ~n7324 & n7362 ;
  assign n7364 = ~n5111 & ~n5124 ;
  assign n7365 = ~n5111 & n5125 ;
  assign n7366 = ~n5113 & ~n7365 ;
  assign n7367 = ~n7364 & n7366 ;
  assign n7368 = ~n5113 & ~n5125 ;
  assign n7369 = n5120 & ~n5121 ;
  assign n7370 = n7368 & n7369 ;
  assign n7371 = ~n5118 & ~n7370 ;
  assign n7372 = ~n7367 & n7371 ;
  assign n7373 = \s2_msel_arb1_state_reg[1]/NET0131  & ~\s2_msel_arb1_state_reg[2]/NET0131  ;
  assign n7374 = ~n5117 & n7373 ;
  assign n7375 = ~n7372 & n7374 ;
  assign n7376 = ~\s2_msel_arb1_state_reg[0]/NET0131  & n7375 ;
  assign n7377 = n5111 & ~n5113 ;
  assign n7378 = ~n7368 & ~n7377 ;
  assign n7379 = n5121 & ~n5124 ;
  assign n7380 = ~n5117 & n5118 ;
  assign n7381 = ~n5120 & ~n5124 ;
  assign n7382 = ~n7380 & n7381 ;
  assign n7383 = ~n7379 & ~n7382 ;
  assign n7384 = \s2_msel_arb1_state_reg[0]/NET0131  & ~n5121 ;
  assign n7385 = ~n5117 & n7384 ;
  assign n7386 = ~n7377 & ~n7385 ;
  assign n7387 = ~n7383 & n7386 ;
  assign n7388 = ~n7378 & ~n7387 ;
  assign n7389 = ~\s2_msel_arb1_state_reg[1]/NET0131  & \s2_msel_arb1_state_reg[2]/NET0131  ;
  assign n7390 = ~\s2_msel_arb1_state_reg[0]/NET0131  & n7389 ;
  assign n7391 = n7388 & n7390 ;
  assign n7392 = ~n7376 & ~n7391 ;
  assign n7393 = ~n5118 & ~n7367 ;
  assign n7394 = ~n7369 & ~n7385 ;
  assign n7395 = n7368 & ~n7394 ;
  assign n7396 = n7393 & ~n7395 ;
  assign n7397 = n7373 & ~n7396 ;
  assign n7398 = ~\s2_msel_arb1_state_reg[1]/NET0131  & ~\s2_msel_arb1_state_reg[2]/NET0131  ;
  assign n7399 = ~n5120 & ~n7380 ;
  assign n7400 = ~n5117 & n7377 ;
  assign n7401 = n7399 & ~n7400 ;
  assign n7402 = ~n5117 & n7368 ;
  assign n7403 = ~n5124 & ~n7384 ;
  assign n7404 = n7402 & ~n7403 ;
  assign n7405 = n7401 & ~n7404 ;
  assign n7406 = n7398 & ~n7405 ;
  assign n7407 = ~n5113 & ~n5117 ;
  assign n7408 = n7384 & n7407 ;
  assign n7409 = ~n5111 & ~n7408 ;
  assign n7410 = ~n7383 & n7409 ;
  assign n7411 = ~n7365 & n7389 ;
  assign n7412 = ~n7410 & n7411 ;
  assign n7413 = ~n7406 & ~n7412 ;
  assign n7414 = ~n7397 & n7413 ;
  assign n7415 = \s2_msel_arb1_state_reg[0]/NET0131  & ~n7414 ;
  assign n7416 = ~\rf_conf2_reg[13]/NET0131  & ~\s2_msel_arb1_state_reg[0]/NET0131  ;
  assign n7417 = n3962 & n7416 ;
  assign n7418 = \s2_msel_arb1_state_reg[1]/NET0131  & \s2_msel_arb1_state_reg[2]/NET0131  ;
  assign n7419 = ~n7417 & n7418 ;
  assign n7420 = n5124 & n7419 ;
  assign n7421 = \s2_msel_arb1_state_reg[0]/NET0131  & ~n5117 ;
  assign n7422 = n7368 & n7421 ;
  assign n7423 = n7401 & ~n7422 ;
  assign n7424 = n7419 & ~n7423 ;
  assign n7425 = ~n5121 & n7424 ;
  assign n7426 = ~n5117 & ~n7364 ;
  assign n7427 = n7366 & n7426 ;
  assign n7428 = ~n7380 & ~n7427 ;
  assign n7429 = ~n5120 & n7428 ;
  assign n7430 = ~\s2_msel_arb1_state_reg[0]/NET0131  & n7398 ;
  assign n7431 = ~n5121 & n7430 ;
  assign n7432 = ~n7429 & n7431 ;
  assign n7433 = ~n7425 & ~n7432 ;
  assign n7434 = ~n7420 & n7433 ;
  assign n7435 = ~n7415 & n7434 ;
  assign n7436 = n7392 & n7435 ;
  assign n7437 = \rf_conf2_reg[9]/NET0131  & n3437 ;
  assign n7438 = \rf_conf2_reg[15]/NET0131  & n3442 ;
  assign n7439 = \rf_conf2_reg[1]/NET0131  & n3451 ;
  assign n7440 = ~n7438 & n7439 ;
  assign n7441 = \rf_conf2_reg[7]/NET0131  & n3432 ;
  assign n7442 = \rf_conf2_reg[5]/NET0131  & n3434 ;
  assign n7443 = n7441 & ~n7442 ;
  assign n7444 = \rf_conf2_reg[3]/NET0131  & n3449 ;
  assign n7445 = ~n7438 & ~n7444 ;
  assign n7446 = ~n7443 & n7445 ;
  assign n7447 = ~n7440 & ~n7446 ;
  assign n7448 = \rf_conf2_reg[11]/NET0131  & n3439 ;
  assign n7449 = ~n7447 & ~n7448 ;
  assign n7450 = \rf_conf2_reg[13]/NET0131  & n3444 ;
  assign n7451 = ~n7448 & n7450 ;
  assign n7452 = \s2_msel_arb2_state_reg[0]/NET0131  & ~n7451 ;
  assign n7453 = ~n7449 & n7452 ;
  assign n7454 = n7437 & ~n7453 ;
  assign n7455 = ~n7439 & ~n7450 ;
  assign n7456 = \s2_msel_arb2_state_reg[0]/NET0131  & ~n7442 ;
  assign n7457 = n7455 & n7456 ;
  assign n7458 = n7451 & ~n7457 ;
  assign n7459 = ~n7448 & ~n7457 ;
  assign n7460 = ~n7447 & n7459 ;
  assign n7461 = ~n7458 & ~n7460 ;
  assign n7462 = ~\s2_msel_arb2_state_reg[1]/NET0131  & \s2_msel_arb2_state_reg[2]/NET0131  ;
  assign n7463 = n7461 & n7462 ;
  assign n7464 = ~n7454 & n7463 ;
  assign n7465 = \s2_msel_arb2_state_reg[1]/NET0131  & \s2_msel_arb2_state_reg[2]/NET0131  ;
  assign n7466 = n7438 & ~n7450 ;
  assign n7467 = n7465 & n7466 ;
  assign n7468 = ~n7443 & ~n7444 ;
  assign n7469 = ~\s2_msel_arb2_state_reg[0]/NET0131  & ~n7448 ;
  assign n7470 = ~n7437 & ~n7442 ;
  assign n7471 = ~n7469 & n7470 ;
  assign n7472 = n7468 & ~n7471 ;
  assign n7473 = n7455 & n7465 ;
  assign n7474 = ~n7472 & n7473 ;
  assign n7475 = ~n7467 & ~n7474 ;
  assign n7476 = ~\s2_msel_arb2_state_reg[1]/NET0131  & ~\s2_msel_arb2_state_reg[2]/NET0131  ;
  assign n7477 = ~n7439 & n7444 ;
  assign n7478 = n7476 & n7477 ;
  assign n7479 = n7437 & ~n7441 ;
  assign n7480 = ~n7441 & ~n7448 ;
  assign n7481 = ~n7466 & n7480 ;
  assign n7482 = ~n7479 & ~n7481 ;
  assign n7483 = ~n7439 & ~n7442 ;
  assign n7484 = n7476 & n7483 ;
  assign n7485 = n7482 & n7484 ;
  assign n7486 = ~n7478 & ~n7485 ;
  assign n7487 = n7475 & n7486 ;
  assign n7488 = ~\s2_msel_arb2_state_reg[0]/NET0131  & ~n7487 ;
  assign n7489 = n7444 & n7476 ;
  assign n7490 = \s2_msel_arb2_state_reg[0]/NET0131  & n7489 ;
  assign n7491 = ~n7439 & ~n7451 ;
  assign n7492 = n7471 & n7491 ;
  assign n7493 = ~n7447 & ~n7492 ;
  assign n7494 = \s2_msel_arb2_state_reg[0]/NET0131  & n7465 ;
  assign n7495 = ~n7493 & n7494 ;
  assign n7496 = ~n7490 & ~n7495 ;
  assign n7497 = ~n7444 & n7476 ;
  assign n7498 = n7456 & n7497 ;
  assign n7499 = \rf_conf2_reg[5]/NET0131  & ~\s2_msel_arb2_state_reg[0]/NET0131  ;
  assign n7500 = n3434 & n7499 ;
  assign n7501 = \s2_msel_arb2_state_reg[1]/NET0131  & ~\s2_msel_arb2_state_reg[2]/NET0131  ;
  assign n7502 = ~n7500 & n7501 ;
  assign n7503 = ~n7498 & ~n7502 ;
  assign n7504 = n7482 & ~n7503 ;
  assign n7505 = n7455 & n7498 ;
  assign n7506 = ~n7437 & n7505 ;
  assign n7507 = ~n7450 & n7477 ;
  assign n7508 = ~n7457 & ~n7507 ;
  assign n7509 = ~n7437 & n7502 ;
  assign n7510 = ~n7508 & n7509 ;
  assign n7511 = ~n7506 & ~n7510 ;
  assign n7512 = ~n7504 & n7511 ;
  assign n7513 = n7496 & n7512 ;
  assign n7514 = ~n7488 & n7513 ;
  assign n7515 = ~n7464 & n7514 ;
  assign n7516 = \s2_msel_arb3_state_reg[1]/NET0131  & ~\s2_msel_arb3_state_reg[2]/NET0131  ;
  assign n7517 = ~n3982 & n7516 ;
  assign n7518 = ~n3949 & ~n3961 ;
  assign n7519 = ~n3949 & n3963 ;
  assign n7520 = ~n7518 & ~n7519 ;
  assign n7521 = n7517 & n7520 ;
  assign n7522 = ~n3971 & ~n3989 ;
  assign n7523 = ~n3963 & ~n3973 ;
  assign n7524 = n7517 & n7523 ;
  assign n7525 = ~n7522 & n7524 ;
  assign n7526 = ~n7521 & ~n7525 ;
  assign n7527 = ~n3951 & ~n7526 ;
  assign n7528 = n3966 & ~n3968 ;
  assign n7529 = ~n3971 & ~n7528 ;
  assign n7530 = ~n3973 & ~n7529 ;
  assign n7531 = n7518 & ~n7530 ;
  assign n7532 = ~\s2_msel_arb3_state_reg[0]/NET0131  & \s2_msel_arb3_state_reg[2]/NET0131  ;
  assign n7533 = ~\s2_msel_arb3_state_reg[1]/NET0131  & n7532 ;
  assign n7534 = ~n7519 & n7533 ;
  assign n7535 = ~n3951 & n7534 ;
  assign n7536 = ~n7531 & n7535 ;
  assign n7537 = ~n7527 & ~n7536 ;
  assign n7538 = ~\s2_msel_arb3_state_reg[1]/NET0131  & ~\s2_msel_arb3_state_reg[2]/NET0131  ;
  assign n7539 = \rf_conf2_reg[1]/NET0131  & ~\s2_msel_arb3_state_reg[0]/NET0131  ;
  assign n7540 = n3972 & n7539 ;
  assign n7541 = n7538 & ~n7540 ;
  assign n7542 = ~n7529 & n7541 ;
  assign n7543 = ~n3951 & ~n3968 ;
  assign n7544 = n7541 & n7543 ;
  assign n7545 = n7520 & n7544 ;
  assign n7546 = ~n7542 & ~n7545 ;
  assign n7547 = n3966 & n7517 ;
  assign n7548 = ~\s2_msel_arb3_state_reg[1]/NET0131  & n3954 ;
  assign n7549 = n3949 & n7548 ;
  assign n7550 = ~n7547 & ~n7549 ;
  assign n7551 = n7546 & n7550 ;
  assign n7552 = n7537 & n7551 ;
  assign n7553 = \s2_msel_arb3_state_reg[0]/NET0131  & n7538 ;
  assign n7554 = ~n3973 & n7553 ;
  assign n7555 = n7543 & n7554 ;
  assign n7556 = ~n3949 & n7548 ;
  assign n7557 = ~n7555 & ~n7556 ;
  assign n7558 = ~n3961 & n3973 ;
  assign n7559 = ~n3961 & ~n3971 ;
  assign n7560 = ~n7528 & n7559 ;
  assign n7561 = ~n7558 & ~n7560 ;
  assign n7562 = \s2_msel_arb3_state_reg[0]/NET0131  & ~n3973 ;
  assign n7563 = n7543 & n7562 ;
  assign n7564 = ~n7555 & ~n7563 ;
  assign n7565 = ~n7561 & n7564 ;
  assign n7566 = ~n7557 & ~n7565 ;
  assign n7567 = ~n3963 & n7566 ;
  assign n7568 = ~n3973 & n7543 ;
  assign n7569 = ~\s2_msel_arb3_state_reg[0]/NET0131  & ~n3949 ;
  assign n7570 = n7568 & ~n7569 ;
  assign n7571 = ~n7561 & ~n7570 ;
  assign n7572 = ~\s2_msel_arb3_state_reg[0]/NET0131  & n3963 ;
  assign n7573 = n3963 & n7518 ;
  assign n7574 = n7529 & n7573 ;
  assign n7575 = ~n7572 & ~n7574 ;
  assign n7576 = n3996 & n7575 ;
  assign n7577 = ~n7571 & n7576 ;
  assign n7578 = ~n7567 & ~n7577 ;
  assign n7579 = n7552 & n7578 ;
  assign n7580 = ~n3070 & n3083 ;
  assign n7581 = n3065 & ~n3067 ;
  assign n7582 = ~n3062 & n7581 ;
  assign n7583 = ~n3067 & ~n3072 ;
  assign n7584 = \s3_msel_arb0_state_reg[0]/NET0131  & ~n3062 ;
  assign n7585 = n7583 & n7584 ;
  assign n7586 = ~n7582 & ~n7585 ;
  assign n7587 = n3062 & ~n3077 ;
  assign n7588 = ~n3060 & ~n3077 ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = ~n3070 & ~n7589 ;
  assign n7591 = n7586 & n7590 ;
  assign n7592 = ~n7580 & ~n7591 ;
  assign n7593 = n3106 & n7592 ;
  assign n7594 = \s3_msel_arb0_state_reg[1]/NET0131  & \s3_msel_arb0_state_reg[2]/NET0131  ;
  assign n7595 = n3077 & ~n3083 ;
  assign n7596 = ~n3070 & ~n7595 ;
  assign n7597 = ~n3072 & ~n7596 ;
  assign n7598 = ~n3062 & ~n3083 ;
  assign n7599 = ~\s3_msel_arb0_state_reg[0]/NET0131  & ~n3060 ;
  assign n7600 = n7598 & ~n7599 ;
  assign n7601 = ~n3060 & n3067 ;
  assign n7602 = ~n3072 & ~n7601 ;
  assign n7603 = n7600 & n7602 ;
  assign n7604 = ~n7597 & ~n7603 ;
  assign n7605 = ~n3065 & n7604 ;
  assign n7606 = n7594 & ~n7605 ;
  assign n7607 = n3070 & ~n3072 ;
  assign n7608 = ~n3060 & ~n3065 ;
  assign n7609 = ~n7607 & n7608 ;
  assign n7610 = ~n7601 & ~n7609 ;
  assign n7611 = \s3_msel_arb0_state_reg[0]/NET0131  & ~n3083 ;
  assign n7612 = n7583 & n7611 ;
  assign n7613 = ~n3077 & ~n7612 ;
  assign n7614 = ~n7610 & n7613 ;
  assign n7615 = \s3_msel_arb0_state_reg[1]/NET0131  & ~\s3_msel_arb0_state_reg[2]/NET0131  ;
  assign n7616 = ~n7587 & n7615 ;
  assign n7617 = ~n7614 & n7616 ;
  assign n7618 = ~n7606 & ~n7617 ;
  assign n7619 = ~n7593 & n7618 ;
  assign n7620 = \s3_msel_arb0_state_reg[0]/NET0131  & ~n7619 ;
  assign n7621 = \s3_msel_arb0_state_reg[0]/NET0131  & n7583 ;
  assign n7622 = n7598 & n7621 ;
  assign n7623 = n7598 & ~n7601 ;
  assign n7624 = ~n7609 & n7623 ;
  assign n7625 = ~n7622 & ~n7624 ;
  assign n7626 = ~n7595 & n7625 ;
  assign n7627 = n7615 & ~n7626 ;
  assign n7628 = n7581 & n7594 ;
  assign n7629 = n7596 & ~n7600 ;
  assign n7630 = n7583 & n7594 ;
  assign n7631 = ~n7629 & n7630 ;
  assign n7632 = ~n7628 & ~n7631 ;
  assign n7633 = n3106 & n7607 ;
  assign n7634 = ~n3062 & ~n3067 ;
  assign n7635 = ~\s3_msel_arb0_state_reg[0]/NET0131  & ~n3065 ;
  assign n7636 = n7634 & ~n7635 ;
  assign n7637 = ~n7589 & ~n7636 ;
  assign n7638 = ~n3072 & ~n3083 ;
  assign n7639 = n3106 & n7638 ;
  assign n7640 = ~n7637 & n7639 ;
  assign n7641 = ~n7633 & ~n7640 ;
  assign n7642 = n7632 & n7641 ;
  assign n7643 = ~n7627 & n7642 ;
  assign n7644 = ~\s3_msel_arb0_state_reg[0]/NET0131  & ~n7643 ;
  assign n7645 = \s3_msel_arb0_state_reg[0]/NET0131  & n7638 ;
  assign n7646 = n7634 & n7645 ;
  assign n7647 = n3110 & n7646 ;
  assign n7648 = n3077 & n7638 ;
  assign n7649 = n7609 & ~n7648 ;
  assign n7650 = ~\rf_conf3_reg[9]/NET0131  & ~\s3_msel_arb0_state_reg[0]/NET0131  ;
  assign n7651 = n3061 & n7650 ;
  assign n7652 = ~n7601 & ~n7651 ;
  assign n7653 = n3110 & n7652 ;
  assign n7654 = ~n7649 & n7653 ;
  assign n7655 = ~n7647 & ~n7654 ;
  assign n7656 = ~n7644 & n7655 ;
  assign n7657 = ~n7620 & n7656 ;
  assign n7658 = ~n5155 & n5156 ;
  assign n7659 = ~n5158 & ~n7658 ;
  assign n7660 = ~n5150 & ~n5155 ;
  assign n7661 = n5151 & n7660 ;
  assign n7662 = n7659 & ~n7661 ;
  assign n7663 = ~n5159 & ~n7662 ;
  assign n7664 = \s3_msel_arb1_state_reg[0]/NET0131  & ~n5159 ;
  assign n7665 = n7660 & n7664 ;
  assign n7666 = ~n5146 & ~n7665 ;
  assign n7667 = ~n7663 & n7666 ;
  assign n7668 = \s3_msel_arb1_state_reg[1]/NET0131  & \s3_msel_arb1_state_reg[2]/NET0131  ;
  assign n7669 = ~n5147 & n7668 ;
  assign n7670 = ~n7667 & n7669 ;
  assign n7671 = ~n5159 & ~n7659 ;
  assign n7672 = ~n5146 & ~n5151 ;
  assign n7673 = ~n5155 & n7664 ;
  assign n7674 = n7672 & ~n7673 ;
  assign n7675 = ~n7671 & n7674 ;
  assign n7676 = n5147 & ~n5151 ;
  assign n7677 = ~\s3_msel_arb1_state_reg[1]/NET0131  & \s3_msel_arb1_state_reg[2]/NET0131  ;
  assign n7678 = ~n5150 & n7677 ;
  assign n7679 = ~n7676 & n7678 ;
  assign n7680 = ~n7675 & n7679 ;
  assign n7681 = ~\s3_msel_arb1_state_reg[1]/NET0131  & ~\s3_msel_arb1_state_reg[2]/NET0131  ;
  assign n7682 = ~n5159 & n7681 ;
  assign n7683 = ~n7659 & n7682 ;
  assign n7684 = n7660 & ~n7676 ;
  assign n7685 = ~n7672 & n7682 ;
  assign n7686 = n7684 & n7685 ;
  assign n7687 = ~n7683 & ~n7686 ;
  assign n7688 = ~n7680 & n7687 ;
  assign n7689 = ~n7670 & n7688 ;
  assign n7690 = ~\s3_msel_arb1_state_reg[0]/NET0131  & ~n7689 ;
  assign n7691 = n5158 & ~n5159 ;
  assign n7692 = n7672 & ~n7691 ;
  assign n7693 = n7684 & ~n7692 ;
  assign n7694 = ~n7658 & ~n7693 ;
  assign n7695 = n5145 & ~n7694 ;
  assign n7696 = ~\s3_msel_arb1_state_reg[2]/NET0131  & n7695 ;
  assign n7697 = \s3_msel_arb1_state_reg[1]/NET0131  & ~n5156 ;
  assign n7698 = \s3_msel_arb1_state_reg[0]/NET0131  & ~n7697 ;
  assign n7699 = ~n7673 & n7692 ;
  assign n7700 = ~n5150 & ~n7676 ;
  assign n7701 = \s3_msel_arb1_state_reg[0]/NET0131  & n7700 ;
  assign n7702 = ~n7699 & n7701 ;
  assign n7703 = ~n7698 & ~n7702 ;
  assign n7704 = ~n5146 & ~n7664 ;
  assign n7705 = ~n5147 & n7660 ;
  assign n7706 = ~n7704 & n7705 ;
  assign n7707 = ~\s3_msel_arb1_state_reg[1]/NET0131  & ~n5158 ;
  assign n7708 = ~n7658 & n7707 ;
  assign n7709 = ~n7661 & n7708 ;
  assign n7710 = ~n7706 & n7709 ;
  assign n7711 = ~\s3_msel_arb1_state_reg[2]/NET0131  & ~n7710 ;
  assign n7712 = ~n7703 & n7711 ;
  assign n7713 = ~n7696 & ~n7712 ;
  assign n7714 = ~n5147 & ~n5159 ;
  assign n7715 = n7660 & n7714 ;
  assign n7716 = ~n5146 & ~n7715 ;
  assign n7717 = ~n7663 & n7716 ;
  assign n7718 = \s3_msel_arb1_state_reg[0]/NET0131  & n7668 ;
  assign n7719 = ~n7717 & n7718 ;
  assign n7720 = ~n7665 & n7672 ;
  assign n7721 = ~n7671 & n7720 ;
  assign n7722 = \s3_msel_arb1_state_reg[0]/NET0131  & n7677 ;
  assign n7723 = ~n7676 & n7722 ;
  assign n7724 = ~n7721 & n7723 ;
  assign n7725 = ~n7719 & ~n7724 ;
  assign n7726 = n7713 & n7725 ;
  assign n7727 = ~n7690 & n7726 ;
  assign n7728 = ~\s3_msel_arb2_state_reg[1]/NET0131  & \s3_msel_arb2_state_reg[2]/NET0131  ;
  assign n7729 = ~n4003 & n7728 ;
  assign n7730 = n4002 & n7729 ;
  assign n7731 = ~n4006 & n4023 ;
  assign n7732 = n4009 & ~n4012 ;
  assign n7733 = ~n4006 & ~n4017 ;
  assign n7734 = ~n7732 & n7733 ;
  assign n7735 = ~n7731 & ~n7734 ;
  assign n7736 = ~n4005 & n7729 ;
  assign n7737 = n7735 & n7736 ;
  assign n7738 = ~n7730 & ~n7737 ;
  assign n7739 = ~\s3_msel_arb2_state_reg[0]/NET0131  & ~n7738 ;
  assign n7740 = ~n4003 & ~n4012 ;
  assign n7741 = ~n7732 & ~n7740 ;
  assign n7742 = ~n4005 & n4006 ;
  assign n7743 = ~n4002 & ~n7742 ;
  assign n7744 = ~n4005 & ~n4023 ;
  assign n7745 = n4017 & n7744 ;
  assign n7746 = n7743 & ~n7745 ;
  assign n7747 = \s3_msel_arb2_state_reg[0]/NET0131  & n7744 ;
  assign n7748 = ~n7732 & ~n7747 ;
  assign n7749 = n7746 & n7748 ;
  assign n7750 = ~n7741 & ~n7749 ;
  assign n7751 = \s3_msel_arb2_state_reg[1]/NET0131  & ~\s3_msel_arb2_state_reg[2]/NET0131  ;
  assign n7752 = ~\s3_msel_arb2_state_reg[0]/NET0131  & n7751 ;
  assign n7753 = n7750 & n7752 ;
  assign n7754 = ~n7739 & ~n7753 ;
  assign n7755 = \s3_msel_arb2_state_reg[0]/NET0131  & ~n4005 ;
  assign n7756 = ~n4002 & ~n7755 ;
  assign n7757 = ~n4023 & n7740 ;
  assign n7758 = ~n7756 & n7757 ;
  assign n7759 = ~n7735 & ~n7758 ;
  assign n7760 = \rf_conf3_reg[13]/NET0131  & ~\s3_msel_arb2_state_reg[0]/NET0131  ;
  assign n7761 = n3066 & n7760 ;
  assign n7762 = \s3_msel_arb2_state_reg[1]/NET0131  & \s3_msel_arb2_state_reg[2]/NET0131  ;
  assign n7763 = ~n7761 & n7762 ;
  assign n7764 = ~n7759 & n7763 ;
  assign n7765 = ~n4003 & ~n7746 ;
  assign n7766 = n7740 & n7747 ;
  assign n7767 = ~n4009 & ~n7766 ;
  assign n7768 = ~n7765 & n7767 ;
  assign n7769 = \s3_msel_arb2_state_reg[0]/NET0131  & n7751 ;
  assign n7770 = ~n7768 & n7769 ;
  assign n7771 = ~n7764 & ~n7770 ;
  assign n7772 = \s3_msel_arb2_state_reg[0]/NET0131  & ~\s3_msel_arb2_state_reg[1]/NET0131  ;
  assign n7773 = \s3_msel_arb2_state_reg[2]/NET0131  & n7772 ;
  assign n7774 = ~n4005 & n7735 ;
  assign n7775 = ~n4002 & ~n7766 ;
  assign n7776 = ~n7774 & n7775 ;
  assign n7777 = n7773 & ~n7776 ;
  assign n7778 = ~n4017 & ~n7732 ;
  assign n7779 = \rf_conf3_reg[1]/NET0131  & ~\s3_msel_arb2_state_reg[0]/NET0131  ;
  assign n7780 = n3071 & n7779 ;
  assign n7781 = ~n7778 & ~n7780 ;
  assign n7782 = n7740 & ~n7780 ;
  assign n7783 = ~n7743 & n7782 ;
  assign n7784 = ~n7781 & ~n7783 ;
  assign n7785 = ~n7766 & n7784 ;
  assign n7786 = ~\s3_msel_arb2_state_reg[1]/NET0131  & ~\s3_msel_arb2_state_reg[2]/NET0131  ;
  assign n7787 = ~n7785 & n7786 ;
  assign n7788 = ~n7777 & ~n7787 ;
  assign n7789 = n7771 & n7788 ;
  assign n7790 = n7754 & n7789 ;
  assign n7791 = ~n4533 & ~n4550 ;
  assign n7792 = n4531 & ~n4533 ;
  assign n7793 = ~n7791 & ~n7792 ;
  assign n7794 = ~n4537 & n4541 ;
  assign n7795 = n4526 & ~n4528 ;
  assign n7796 = ~n4537 & ~n4539 ;
  assign n7797 = ~n7795 & n7796 ;
  assign n7798 = ~n7794 & ~n7797 ;
  assign n7799 = \s3_msel_arb3_state_reg[0]/NET0131  & ~n4541 ;
  assign n7800 = ~n4528 & n7799 ;
  assign n7801 = ~n7792 & ~n7800 ;
  assign n7802 = ~n7798 & n7801 ;
  assign n7803 = ~n7793 & ~n7802 ;
  assign n7804 = n4567 & n7803 ;
  assign n7805 = ~\s3_msel_arb3_state_reg[1]/NET0131  & ~\s3_msel_arb3_state_reg[2]/NET0131  ;
  assign n7806 = n7795 & n7805 ;
  assign n7807 = ~n4531 & n4550 ;
  assign n7808 = n4539 & ~n4541 ;
  assign n7809 = ~n4531 & ~n4537 ;
  assign n7810 = ~n7808 & n7809 ;
  assign n7811 = ~n7807 & ~n7810 ;
  assign n7812 = ~n4528 & ~n4533 ;
  assign n7813 = n7805 & n7812 ;
  assign n7814 = n7811 & n7813 ;
  assign n7815 = ~n7806 & ~n7814 ;
  assign n7816 = n4524 & ~n4550 ;
  assign n7817 = n4537 & n7816 ;
  assign n7818 = ~n4539 & ~n7795 ;
  assign n7819 = ~n4528 & n7792 ;
  assign n7820 = n7818 & ~n7819 ;
  assign n7821 = ~n4541 & n7816 ;
  assign n7822 = ~n7820 & n7821 ;
  assign n7823 = ~n7817 & ~n7822 ;
  assign n7824 = ~\s3_msel_arb3_state_reg[0]/NET0131  & n7823 ;
  assign n7825 = n7815 & n7824 ;
  assign n7826 = ~n7804 & n7825 ;
  assign n7827 = ~n4541 & ~n7820 ;
  assign n7828 = ~n4528 & ~n4541 ;
  assign n7829 = n7791 & n7828 ;
  assign n7830 = ~n4537 & ~n7829 ;
  assign n7831 = ~n7827 & n7830 ;
  assign n7832 = n4524 & ~n7831 ;
  assign n7833 = n4531 & n4567 ;
  assign n7834 = \s3_msel_arb3_state_reg[0]/NET0131  & ~n7833 ;
  assign n7835 = ~n7832 & n7834 ;
  assign n7836 = ~n7826 & ~n7835 ;
  assign n7837 = ~n4526 & n4533 ;
  assign n7838 = ~n4528 & ~n4550 ;
  assign n7839 = n7799 & n7838 ;
  assign n7840 = ~n4526 & ~n7839 ;
  assign n7841 = ~n7811 & n7840 ;
  assign n7842 = ~n7837 & ~n7841 ;
  assign n7843 = \s3_msel_arb3_state_reg[0]/NET0131  & n7805 ;
  assign n7844 = n7842 & n7843 ;
  assign n7845 = ~n4537 & ~n7799 ;
  assign n7846 = ~n4528 & n7791 ;
  assign n7847 = ~n7845 & n7846 ;
  assign n7848 = n7820 & ~n7847 ;
  assign n7849 = \rf_conf3_reg[13]/NET0131  & ~\s3_msel_arb3_state_reg[0]/NET0131  ;
  assign n7850 = n4540 & n7849 ;
  assign n7851 = n4547 & ~n7850 ;
  assign n7852 = ~n7848 & n7851 ;
  assign n7853 = n7799 & n7812 ;
  assign n7854 = ~n7798 & ~n7853 ;
  assign n7855 = \s3_msel_arb3_state_reg[0]/NET0131  & n4567 ;
  assign n7856 = ~n4531 & n7855 ;
  assign n7857 = ~n4550 & n7856 ;
  assign n7858 = ~n7854 & n7857 ;
  assign n7859 = ~n7852 & ~n7858 ;
  assign n7860 = ~n7844 & n7859 ;
  assign n7861 = ~n7836 & n7860 ;
  assign n7862 = ~n3132 & n3145 ;
  assign n7863 = n3127 & ~n3129 ;
  assign n7864 = ~n3124 & n7863 ;
  assign n7865 = ~n3129 & ~n3134 ;
  assign n7866 = \s4_msel_arb0_state_reg[0]/NET0131  & ~n3124 ;
  assign n7867 = n7865 & n7866 ;
  assign n7868 = ~n7864 & ~n7867 ;
  assign n7869 = n3124 & ~n3139 ;
  assign n7870 = ~n3122 & ~n3139 ;
  assign n7871 = ~n7869 & ~n7870 ;
  assign n7872 = ~n3132 & ~n7871 ;
  assign n7873 = n7868 & n7872 ;
  assign n7874 = ~n7862 & ~n7873 ;
  assign n7875 = n3168 & n7874 ;
  assign n7876 = \s4_msel_arb0_state_reg[1]/NET0131  & \s4_msel_arb0_state_reg[2]/NET0131  ;
  assign n7877 = n3139 & ~n3145 ;
  assign n7878 = ~n3132 & ~n7877 ;
  assign n7879 = ~n3134 & ~n7878 ;
  assign n7880 = ~n3124 & ~n3145 ;
  assign n7881 = ~\s4_msel_arb0_state_reg[0]/NET0131  & ~n3122 ;
  assign n7882 = n7880 & ~n7881 ;
  assign n7883 = ~n3122 & n3129 ;
  assign n7884 = ~n3134 & ~n7883 ;
  assign n7885 = n7882 & n7884 ;
  assign n7886 = ~n7879 & ~n7885 ;
  assign n7887 = ~n3127 & n7886 ;
  assign n7888 = n7876 & ~n7887 ;
  assign n7889 = n3132 & ~n3134 ;
  assign n7890 = ~n3122 & ~n3127 ;
  assign n7891 = ~n7889 & n7890 ;
  assign n7892 = ~n7883 & ~n7891 ;
  assign n7893 = \s4_msel_arb0_state_reg[0]/NET0131  & ~n3145 ;
  assign n7894 = n7865 & n7893 ;
  assign n7895 = ~n3139 & ~n7894 ;
  assign n7896 = ~n7892 & n7895 ;
  assign n7897 = \s4_msel_arb0_state_reg[1]/NET0131  & ~\s4_msel_arb0_state_reg[2]/NET0131  ;
  assign n7898 = ~n7869 & n7897 ;
  assign n7899 = ~n7896 & n7898 ;
  assign n7900 = ~n7888 & ~n7899 ;
  assign n7901 = ~n7875 & n7900 ;
  assign n7902 = \s4_msel_arb0_state_reg[0]/NET0131  & ~n7901 ;
  assign n7903 = \s4_msel_arb0_state_reg[0]/NET0131  & n7865 ;
  assign n7904 = n7880 & n7903 ;
  assign n7905 = n7880 & ~n7883 ;
  assign n7906 = ~n7891 & n7905 ;
  assign n7907 = ~n7904 & ~n7906 ;
  assign n7908 = ~n7877 & n7907 ;
  assign n7909 = n7897 & ~n7908 ;
  assign n7910 = n7863 & n7876 ;
  assign n7911 = n7878 & ~n7882 ;
  assign n7912 = n7865 & n7876 ;
  assign n7913 = ~n7911 & n7912 ;
  assign n7914 = ~n7910 & ~n7913 ;
  assign n7915 = n3168 & n7889 ;
  assign n7916 = ~n3124 & ~n3129 ;
  assign n7917 = ~\s4_msel_arb0_state_reg[0]/NET0131  & ~n3127 ;
  assign n7918 = n7916 & ~n7917 ;
  assign n7919 = ~n7871 & ~n7918 ;
  assign n7920 = ~n3134 & ~n3145 ;
  assign n7921 = n3168 & n7920 ;
  assign n7922 = ~n7919 & n7921 ;
  assign n7923 = ~n7915 & ~n7922 ;
  assign n7924 = n7914 & n7923 ;
  assign n7925 = ~n7909 & n7924 ;
  assign n7926 = ~\s4_msel_arb0_state_reg[0]/NET0131  & ~n7925 ;
  assign n7927 = \s4_msel_arb0_state_reg[0]/NET0131  & n7920 ;
  assign n7928 = n7916 & n7927 ;
  assign n7929 = n3172 & n7928 ;
  assign n7930 = n3139 & n7920 ;
  assign n7931 = n7891 & ~n7930 ;
  assign n7932 = ~\rf_conf4_reg[9]/NET0131  & ~\s4_msel_arb0_state_reg[0]/NET0131  ;
  assign n7933 = n3123 & n7932 ;
  assign n7934 = ~n7883 & ~n7933 ;
  assign n7935 = n3172 & n7934 ;
  assign n7936 = ~n7931 & n7935 ;
  assign n7937 = ~n7929 & ~n7936 ;
  assign n7938 = ~n7926 & n7937 ;
  assign n7939 = ~n7902 & n7938 ;
  assign n7940 = n5190 & ~n5196 ;
  assign n7941 = ~n5187 & n5188 ;
  assign n7942 = ~n5191 & ~n5196 ;
  assign n7943 = ~n7941 & n7942 ;
  assign n7944 = ~n7940 & ~n7943 ;
  assign n7945 = ~n5202 & ~n7944 ;
  assign n7946 = n5201 & ~n5202 ;
  assign n7947 = ~\s4_msel_arb1_state_reg[1]/NET0131  & ~\s4_msel_arb1_state_reg[2]/NET0131  ;
  assign n7948 = ~n5212 & n7947 ;
  assign n7949 = ~n7946 & n7948 ;
  assign n7950 = ~n7945 & n7949 ;
  assign n7951 = n5196 & ~n5201 ;
  assign n7952 = \s4_msel_arb1_state_reg[1]/NET0131  & ~\s4_msel_arb1_state_reg[2]/NET0131  ;
  assign n7953 = n7951 & n7952 ;
  assign n7954 = ~n5191 & ~n7941 ;
  assign n7955 = ~n5187 & ~n5212 ;
  assign n7956 = ~\s4_msel_arb1_state_reg[0]/NET0131  & ~n5202 ;
  assign n7957 = n7955 & ~n7956 ;
  assign n7958 = n7954 & ~n7957 ;
  assign n7959 = ~n5190 & ~n5201 ;
  assign n7960 = n7952 & n7959 ;
  assign n7961 = ~n7958 & n7960 ;
  assign n7962 = ~n7953 & ~n7961 ;
  assign n7963 = ~n5190 & n5194 ;
  assign n7964 = ~n7954 & n7963 ;
  assign n7965 = ~n5202 & ~n7951 ;
  assign n7966 = n7955 & n7963 ;
  assign n7967 = ~n7965 & n7966 ;
  assign n7968 = ~n7964 & ~n7967 ;
  assign n7969 = n7962 & n7968 ;
  assign n7970 = ~n7950 & n7969 ;
  assign n7971 = ~\s4_msel_arb1_state_reg[0]/NET0131  & ~n7970 ;
  assign n7972 = \s4_msel_arb1_state_reg[0]/NET0131  & ~n5212 ;
  assign n7973 = ~n5187 & n7959 ;
  assign n7974 = n7972 & n7973 ;
  assign n7975 = ~\rf_conf4_reg[13]/NET0131  & ~\s4_msel_arb1_state_reg[0]/NET0131  ;
  assign n7976 = n4053 & n7975 ;
  assign n7977 = n5188 & ~n7976 ;
  assign n7978 = n5191 & n7959 ;
  assign n7979 = n7965 & ~n7978 ;
  assign n7980 = ~n5212 & ~n7976 ;
  assign n7981 = ~n7979 & n7980 ;
  assign n7982 = ~n7977 & ~n7981 ;
  assign n7983 = ~n7974 & n7982 ;
  assign n7984 = \s4_msel_arb1_state_reg[1]/NET0131  & \s4_msel_arb1_state_reg[2]/NET0131  ;
  assign n7985 = ~n7983 & n7984 ;
  assign n7986 = \s4_msel_arb1_state_reg[0]/NET0131  & ~\s4_msel_arb1_state_reg[1]/NET0131  ;
  assign n7987 = \s4_msel_arb1_state_reg[2]/NET0131  & n7986 ;
  assign n7988 = n7955 & ~n7965 ;
  assign n7989 = n7954 & ~n7988 ;
  assign n7990 = ~n7974 & n7989 ;
  assign n7991 = n7987 & ~n7990 ;
  assign n7992 = ~n5188 & ~n7972 ;
  assign n7993 = n7973 & ~n7992 ;
  assign n7994 = n7979 & ~n7993 ;
  assign n7995 = \s4_msel_arb1_state_reg[0]/NET0131  & n7947 ;
  assign n7996 = ~n7994 & n7995 ;
  assign n7997 = ~n5190 & ~n7946 ;
  assign n7998 = n7957 & n7997 ;
  assign n7999 = ~n7944 & ~n7998 ;
  assign n8000 = \s4_msel_arb1_state_reg[0]/NET0131  & n7952 ;
  assign n8001 = ~n7999 & n8000 ;
  assign n8002 = ~n7996 & ~n8001 ;
  assign n8003 = ~n7991 & n8002 ;
  assign n8004 = ~n7985 & n8003 ;
  assign n8005 = ~n7971 & n8004 ;
  assign n8006 = \rf_conf4_reg[9]/NET0131  & n3123 ;
  assign n8007 = \rf_conf4_reg[15]/NET0131  & n3126 ;
  assign n8008 = \rf_conf4_reg[1]/NET0131  & n3133 ;
  assign n8009 = ~n8007 & n8008 ;
  assign n8010 = \rf_conf4_reg[7]/NET0131  & n3138 ;
  assign n8011 = \rf_conf4_reg[5]/NET0131  & n3144 ;
  assign n8012 = n8010 & ~n8011 ;
  assign n8013 = \rf_conf4_reg[3]/NET0131  & n3131 ;
  assign n8014 = ~n8007 & ~n8013 ;
  assign n8015 = ~n8012 & n8014 ;
  assign n8016 = ~n8009 & ~n8015 ;
  assign n8017 = \rf_conf4_reg[11]/NET0131  & n3121 ;
  assign n8018 = ~n8016 & ~n8017 ;
  assign n8019 = \rf_conf4_reg[13]/NET0131  & n3128 ;
  assign n8020 = ~n8017 & n8019 ;
  assign n8021 = \s4_msel_arb2_state_reg[0]/NET0131  & ~n8020 ;
  assign n8022 = ~n8018 & n8021 ;
  assign n8023 = n8006 & ~n8022 ;
  assign n8024 = ~n8008 & ~n8019 ;
  assign n8025 = \s4_msel_arb2_state_reg[0]/NET0131  & ~n8011 ;
  assign n8026 = n8024 & n8025 ;
  assign n8027 = n8020 & ~n8026 ;
  assign n8028 = ~n8017 & ~n8026 ;
  assign n8029 = ~n8016 & n8028 ;
  assign n8030 = ~n8027 & ~n8029 ;
  assign n8031 = ~\s4_msel_arb2_state_reg[1]/NET0131  & \s4_msel_arb2_state_reg[2]/NET0131  ;
  assign n8032 = n8030 & n8031 ;
  assign n8033 = ~n8023 & n8032 ;
  assign n8034 = \s4_msel_arb2_state_reg[1]/NET0131  & \s4_msel_arb2_state_reg[2]/NET0131  ;
  assign n8035 = n8007 & ~n8019 ;
  assign n8036 = n8034 & n8035 ;
  assign n8037 = ~n8012 & ~n8013 ;
  assign n8038 = ~\s4_msel_arb2_state_reg[0]/NET0131  & ~n8017 ;
  assign n8039 = ~n8006 & ~n8011 ;
  assign n8040 = ~n8038 & n8039 ;
  assign n8041 = n8037 & ~n8040 ;
  assign n8042 = n8024 & n8034 ;
  assign n8043 = ~n8041 & n8042 ;
  assign n8044 = ~n8036 & ~n8043 ;
  assign n8045 = ~\s4_msel_arb2_state_reg[1]/NET0131  & ~\s4_msel_arb2_state_reg[2]/NET0131  ;
  assign n8046 = ~n8008 & n8013 ;
  assign n8047 = n8045 & n8046 ;
  assign n8048 = n8006 & ~n8010 ;
  assign n8049 = ~n8010 & ~n8017 ;
  assign n8050 = ~n8035 & n8049 ;
  assign n8051 = ~n8048 & ~n8050 ;
  assign n8052 = ~n8008 & ~n8011 ;
  assign n8053 = n8045 & n8052 ;
  assign n8054 = n8051 & n8053 ;
  assign n8055 = ~n8047 & ~n8054 ;
  assign n8056 = n8044 & n8055 ;
  assign n8057 = ~\s4_msel_arb2_state_reg[0]/NET0131  & ~n8056 ;
  assign n8058 = n8013 & n8045 ;
  assign n8059 = \s4_msel_arb2_state_reg[0]/NET0131  & n8058 ;
  assign n8060 = ~n8008 & ~n8020 ;
  assign n8061 = n8040 & n8060 ;
  assign n8062 = ~n8016 & ~n8061 ;
  assign n8063 = \s4_msel_arb2_state_reg[0]/NET0131  & n8034 ;
  assign n8064 = ~n8062 & n8063 ;
  assign n8065 = ~n8059 & ~n8064 ;
  assign n8066 = ~n8013 & n8045 ;
  assign n8067 = n8025 & n8066 ;
  assign n8068 = \rf_conf4_reg[5]/NET0131  & ~\s4_msel_arb2_state_reg[0]/NET0131  ;
  assign n8069 = n3144 & n8068 ;
  assign n8070 = \s4_msel_arb2_state_reg[1]/NET0131  & ~\s4_msel_arb2_state_reg[2]/NET0131  ;
  assign n8071 = ~n8069 & n8070 ;
  assign n8072 = ~n8067 & ~n8071 ;
  assign n8073 = n8051 & ~n8072 ;
  assign n8074 = n8024 & n8067 ;
  assign n8075 = ~n8006 & n8074 ;
  assign n8076 = ~n8019 & n8046 ;
  assign n8077 = ~n8026 & ~n8076 ;
  assign n8078 = ~n8006 & n8071 ;
  assign n8079 = ~n8077 & n8078 ;
  assign n8080 = ~n8075 & ~n8079 ;
  assign n8081 = ~n8073 & n8080 ;
  assign n8082 = n8065 & n8081 ;
  assign n8083 = ~n8057 & n8082 ;
  assign n8084 = ~n8033 & n8083 ;
  assign n8085 = ~n4046 & ~n4063 ;
  assign n8086 = n4044 & ~n4046 ;
  assign n8087 = ~n8085 & ~n8086 ;
  assign n8088 = ~n4050 & n4054 ;
  assign n8089 = n4039 & ~n4041 ;
  assign n8090 = ~n4050 & ~n4052 ;
  assign n8091 = ~n8089 & n8090 ;
  assign n8092 = ~n8088 & ~n8091 ;
  assign n8093 = \s4_msel_arb3_state_reg[0]/NET0131  & ~n4054 ;
  assign n8094 = ~n4041 & n8093 ;
  assign n8095 = ~n8086 & ~n8094 ;
  assign n8096 = ~n8092 & n8095 ;
  assign n8097 = ~n8087 & ~n8096 ;
  assign n8098 = n4080 & n8097 ;
  assign n8099 = ~\s4_msel_arb3_state_reg[1]/NET0131  & ~\s4_msel_arb3_state_reg[2]/NET0131  ;
  assign n8100 = n8089 & n8099 ;
  assign n8101 = ~n4044 & n4063 ;
  assign n8102 = n4052 & ~n4054 ;
  assign n8103 = ~n4044 & ~n4050 ;
  assign n8104 = ~n8102 & n8103 ;
  assign n8105 = ~n8101 & ~n8104 ;
  assign n8106 = ~n4041 & ~n4046 ;
  assign n8107 = n8099 & n8106 ;
  assign n8108 = n8105 & n8107 ;
  assign n8109 = ~n8100 & ~n8108 ;
  assign n8110 = n4037 & ~n4063 ;
  assign n8111 = n4050 & n8110 ;
  assign n8112 = ~n4052 & ~n8089 ;
  assign n8113 = ~n4041 & n8086 ;
  assign n8114 = n8112 & ~n8113 ;
  assign n8115 = ~n4054 & n8110 ;
  assign n8116 = ~n8114 & n8115 ;
  assign n8117 = ~n8111 & ~n8116 ;
  assign n8118 = ~\s4_msel_arb3_state_reg[0]/NET0131  & n8117 ;
  assign n8119 = n8109 & n8118 ;
  assign n8120 = ~n8098 & n8119 ;
  assign n8121 = ~n4054 & ~n8114 ;
  assign n8122 = ~n4041 & ~n4054 ;
  assign n8123 = n8085 & n8122 ;
  assign n8124 = ~n4050 & ~n8123 ;
  assign n8125 = ~n8121 & n8124 ;
  assign n8126 = n4037 & ~n8125 ;
  assign n8127 = n4044 & n4080 ;
  assign n8128 = \s4_msel_arb3_state_reg[0]/NET0131  & ~n8127 ;
  assign n8129 = ~n8126 & n8128 ;
  assign n8130 = ~n8120 & ~n8129 ;
  assign n8131 = ~n4039 & n4046 ;
  assign n8132 = ~n4041 & ~n4063 ;
  assign n8133 = n8093 & n8132 ;
  assign n8134 = ~n4039 & ~n8133 ;
  assign n8135 = ~n8105 & n8134 ;
  assign n8136 = ~n8131 & ~n8135 ;
  assign n8137 = \s4_msel_arb3_state_reg[0]/NET0131  & n8099 ;
  assign n8138 = n8136 & n8137 ;
  assign n8139 = ~n4050 & ~n8093 ;
  assign n8140 = ~n4041 & n8085 ;
  assign n8141 = ~n8139 & n8140 ;
  assign n8142 = n8114 & ~n8141 ;
  assign n8143 = \rf_conf4_reg[13]/NET0131  & ~\s4_msel_arb3_state_reg[0]/NET0131  ;
  assign n8144 = n4053 & n8143 ;
  assign n8145 = n4060 & ~n8144 ;
  assign n8146 = ~n8142 & n8145 ;
  assign n8147 = n8093 & n8106 ;
  assign n8148 = ~n8092 & ~n8147 ;
  assign n8149 = \s4_msel_arb3_state_reg[0]/NET0131  & n4080 ;
  assign n8150 = ~n4044 & n8149 ;
  assign n8151 = ~n4063 & n8150 ;
  assign n8152 = ~n8148 & n8151 ;
  assign n8153 = ~n8146 & ~n8152 ;
  assign n8154 = ~n8138 & n8153 ;
  assign n8155 = ~n8130 & n8154 ;
  assign n8156 = ~n3194 & n3207 ;
  assign n8157 = n3189 & ~n3191 ;
  assign n8158 = ~n3186 & n8157 ;
  assign n8159 = ~n3191 & ~n3196 ;
  assign n8160 = \s5_msel_arb0_state_reg[0]/NET0131  & ~n3186 ;
  assign n8161 = n8159 & n8160 ;
  assign n8162 = ~n8158 & ~n8161 ;
  assign n8163 = n3186 & ~n3201 ;
  assign n8164 = ~n3184 & ~n3201 ;
  assign n8165 = ~n8163 & ~n8164 ;
  assign n8166 = ~n3194 & ~n8165 ;
  assign n8167 = n8162 & n8166 ;
  assign n8168 = ~n8156 & ~n8167 ;
  assign n8169 = n3230 & n8168 ;
  assign n8170 = \s5_msel_arb0_state_reg[1]/NET0131  & \s5_msel_arb0_state_reg[2]/NET0131  ;
  assign n8171 = n3201 & ~n3207 ;
  assign n8172 = ~n3194 & ~n8171 ;
  assign n8173 = ~n3196 & ~n8172 ;
  assign n8174 = ~n3186 & ~n3207 ;
  assign n8175 = ~\s5_msel_arb0_state_reg[0]/NET0131  & ~n3184 ;
  assign n8176 = n8174 & ~n8175 ;
  assign n8177 = ~n3184 & n3191 ;
  assign n8178 = ~n3196 & ~n8177 ;
  assign n8179 = n8176 & n8178 ;
  assign n8180 = ~n8173 & ~n8179 ;
  assign n8181 = ~n3189 & n8180 ;
  assign n8182 = n8170 & ~n8181 ;
  assign n8183 = n3194 & ~n3196 ;
  assign n8184 = ~n3184 & ~n3189 ;
  assign n8185 = ~n8183 & n8184 ;
  assign n8186 = ~n8177 & ~n8185 ;
  assign n8187 = \s5_msel_arb0_state_reg[0]/NET0131  & ~n3207 ;
  assign n8188 = n8159 & n8187 ;
  assign n8189 = ~n3201 & ~n8188 ;
  assign n8190 = ~n8186 & n8189 ;
  assign n8191 = \s5_msel_arb0_state_reg[1]/NET0131  & ~\s5_msel_arb0_state_reg[2]/NET0131  ;
  assign n8192 = ~n8163 & n8191 ;
  assign n8193 = ~n8190 & n8192 ;
  assign n8194 = ~n8182 & ~n8193 ;
  assign n8195 = ~n8169 & n8194 ;
  assign n8196 = \s5_msel_arb0_state_reg[0]/NET0131  & ~n8195 ;
  assign n8197 = \s5_msel_arb0_state_reg[0]/NET0131  & n8159 ;
  assign n8198 = n8174 & n8197 ;
  assign n8199 = n8174 & ~n8177 ;
  assign n8200 = ~n8185 & n8199 ;
  assign n8201 = ~n8198 & ~n8200 ;
  assign n8202 = ~n8171 & n8201 ;
  assign n8203 = n8191 & ~n8202 ;
  assign n8204 = n8157 & n8170 ;
  assign n8205 = n8172 & ~n8176 ;
  assign n8206 = n8159 & n8170 ;
  assign n8207 = ~n8205 & n8206 ;
  assign n8208 = ~n8204 & ~n8207 ;
  assign n8209 = n3230 & n8183 ;
  assign n8210 = ~n3186 & ~n3191 ;
  assign n8211 = ~\s5_msel_arb0_state_reg[0]/NET0131  & ~n3189 ;
  assign n8212 = n8210 & ~n8211 ;
  assign n8213 = ~n8165 & ~n8212 ;
  assign n8214 = ~n3196 & ~n3207 ;
  assign n8215 = n3230 & n8214 ;
  assign n8216 = ~n8213 & n8215 ;
  assign n8217 = ~n8209 & ~n8216 ;
  assign n8218 = n8208 & n8217 ;
  assign n8219 = ~n8203 & n8218 ;
  assign n8220 = ~\s5_msel_arb0_state_reg[0]/NET0131  & ~n8219 ;
  assign n8221 = \s5_msel_arb0_state_reg[0]/NET0131  & n8214 ;
  assign n8222 = n8210 & n8221 ;
  assign n8223 = n3234 & n8222 ;
  assign n8224 = n3201 & n8214 ;
  assign n8225 = n8185 & ~n8224 ;
  assign n8226 = ~\rf_conf5_reg[9]/NET0131  & ~\s5_msel_arb0_state_reg[0]/NET0131  ;
  assign n8227 = n3185 & n8226 ;
  assign n8228 = ~n8177 & ~n8227 ;
  assign n8229 = n3234 & n8228 ;
  assign n8230 = ~n8225 & n8229 ;
  assign n8231 = ~n8223 & ~n8230 ;
  assign n8232 = ~n8220 & n8231 ;
  assign n8233 = ~n8196 & n8232 ;
  assign n8234 = ~n5234 & ~n5238 ;
  assign n8235 = n5235 & ~n5238 ;
  assign n8236 = ~n8234 & ~n8235 ;
  assign n8237 = ~\rf_conf5_reg[9]/NET0131  & ~\s5_msel_arb1_state_reg[0]/NET0131  ;
  assign n8238 = n4612 & n8237 ;
  assign n8239 = ~\s5_msel_arb1_state_reg[1]/NET0131  & \s5_msel_arb1_state_reg[2]/NET0131  ;
  assign n8240 = ~n8238 & n8239 ;
  assign n8241 = n8236 & n8240 ;
  assign n8242 = n5227 & ~n5230 ;
  assign n8243 = ~n5226 & ~n5230 ;
  assign n8244 = ~n8242 & ~n8243 ;
  assign n8245 = ~n5227 & ~n5237 ;
  assign n8246 = \s5_msel_arb1_state_reg[0]/NET0131  & n8245 ;
  assign n8247 = ~n8244 & ~n8246 ;
  assign n8248 = ~n5229 & ~n5235 ;
  assign n8249 = n8240 & n8248 ;
  assign n8250 = ~n8247 & n8249 ;
  assign n8251 = ~n8241 & ~n8250 ;
  assign n8252 = ~n8242 & n8248 ;
  assign n8253 = ~n8236 & ~n8252 ;
  assign n8254 = ~n5237 & ~n8253 ;
  assign n8255 = ~n5226 & ~n8254 ;
  assign n8256 = \s5_msel_arb1_state_reg[0]/NET0131  & n5254 ;
  assign n8257 = n8234 & n8243 ;
  assign n8258 = ~n5227 & n5254 ;
  assign n8259 = ~n8257 & n8258 ;
  assign n8260 = ~n8256 & ~n8259 ;
  assign n8261 = ~n8255 & ~n8260 ;
  assign n8262 = n8251 & ~n8261 ;
  assign n8263 = ~\rf_conf5_reg[1]/NET0131  & ~\s5_msel_arb1_state_reg[0]/NET0131  ;
  assign n8264 = n4634 & n8263 ;
  assign n8265 = n8244 & ~n8264 ;
  assign n8266 = n8245 & ~n8264 ;
  assign n8267 = n8236 & n8266 ;
  assign n8268 = ~n8265 & ~n8267 ;
  assign n8269 = n8246 & n8248 ;
  assign n8270 = n8268 & ~n8269 ;
  assign n8271 = n5241 & ~n8270 ;
  assign n8272 = n5238 & n8245 ;
  assign n8273 = ~n8244 & ~n8272 ;
  assign n8274 = ~n5229 & ~n8273 ;
  assign n8275 = ~n5234 & ~n8269 ;
  assign n8276 = ~n8274 & n8275 ;
  assign n8277 = ~\rf_conf5_reg[13]/NET0131  & ~\s5_msel_arb1_state_reg[0]/NET0131  ;
  assign n8278 = n4624 & n8277 ;
  assign n8279 = \s5_msel_arb1_state_reg[1]/NET0131  & \s5_msel_arb1_state_reg[2]/NET0131  ;
  assign n8280 = ~n8278 & n8279 ;
  assign n8281 = ~n8276 & n8280 ;
  assign n8282 = ~n8271 & ~n8281 ;
  assign n8283 = n8262 & n8282 ;
  assign n8284 = ~\s5_msel_arb2_state_reg[1]/NET0131  & \s5_msel_arb2_state_reg[2]/NET0131  ;
  assign n8285 = ~n4576 & n8284 ;
  assign n8286 = n4575 & n8285 ;
  assign n8287 = ~n4579 & n4596 ;
  assign n8288 = n4582 & ~n4585 ;
  assign n8289 = ~n4579 & ~n4590 ;
  assign n8290 = ~n8288 & n8289 ;
  assign n8291 = ~n8287 & ~n8290 ;
  assign n8292 = ~n4578 & n8285 ;
  assign n8293 = n8291 & n8292 ;
  assign n8294 = ~n8286 & ~n8293 ;
  assign n8295 = ~\s5_msel_arb2_state_reg[0]/NET0131  & ~n8294 ;
  assign n8296 = ~n4576 & ~n4585 ;
  assign n8297 = ~n8288 & ~n8296 ;
  assign n8298 = ~n4578 & n4579 ;
  assign n8299 = ~n4575 & ~n8298 ;
  assign n8300 = ~n4578 & ~n4596 ;
  assign n8301 = n4590 & n8300 ;
  assign n8302 = n8299 & ~n8301 ;
  assign n8303 = \s5_msel_arb2_state_reg[0]/NET0131  & n8300 ;
  assign n8304 = ~n8288 & ~n8303 ;
  assign n8305 = n8302 & n8304 ;
  assign n8306 = ~n8297 & ~n8305 ;
  assign n8307 = \s5_msel_arb2_state_reg[1]/NET0131  & ~\s5_msel_arb2_state_reg[2]/NET0131  ;
  assign n8308 = ~\s5_msel_arb2_state_reg[0]/NET0131  & n8307 ;
  assign n8309 = n8306 & n8308 ;
  assign n8310 = ~n8295 & ~n8309 ;
  assign n8311 = \s5_msel_arb2_state_reg[0]/NET0131  & ~n4578 ;
  assign n8312 = ~n4575 & ~n8311 ;
  assign n8313 = ~n4596 & n8296 ;
  assign n8314 = ~n8312 & n8313 ;
  assign n8315 = ~n8291 & ~n8314 ;
  assign n8316 = \rf_conf5_reg[13]/NET0131  & ~\s5_msel_arb2_state_reg[0]/NET0131  ;
  assign n8317 = n3190 & n8316 ;
  assign n8318 = \s5_msel_arb2_state_reg[1]/NET0131  & \s5_msel_arb2_state_reg[2]/NET0131  ;
  assign n8319 = ~n8317 & n8318 ;
  assign n8320 = ~n8315 & n8319 ;
  assign n8321 = ~n4576 & ~n8302 ;
  assign n8322 = n8296 & n8303 ;
  assign n8323 = ~n4582 & ~n8322 ;
  assign n8324 = ~n8321 & n8323 ;
  assign n8325 = \s5_msel_arb2_state_reg[0]/NET0131  & n8307 ;
  assign n8326 = ~n8324 & n8325 ;
  assign n8327 = ~n8320 & ~n8326 ;
  assign n8328 = \s5_msel_arb2_state_reg[0]/NET0131  & ~\s5_msel_arb2_state_reg[1]/NET0131  ;
  assign n8329 = \s5_msel_arb2_state_reg[2]/NET0131  & n8328 ;
  assign n8330 = ~n4578 & n8291 ;
  assign n8331 = ~n4575 & ~n8322 ;
  assign n8332 = ~n8330 & n8331 ;
  assign n8333 = n8329 & ~n8332 ;
  assign n8334 = ~n4590 & ~n8288 ;
  assign n8335 = \rf_conf5_reg[1]/NET0131  & ~\s5_msel_arb2_state_reg[0]/NET0131  ;
  assign n8336 = n3195 & n8335 ;
  assign n8337 = ~n8334 & ~n8336 ;
  assign n8338 = n8296 & ~n8336 ;
  assign n8339 = ~n8299 & n8338 ;
  assign n8340 = ~n8337 & ~n8339 ;
  assign n8341 = ~n8322 & n8340 ;
  assign n8342 = ~\s5_msel_arb2_state_reg[1]/NET0131  & ~\s5_msel_arb2_state_reg[2]/NET0131  ;
  assign n8343 = ~n8341 & n8342 ;
  assign n8344 = ~n8333 & ~n8343 ;
  assign n8345 = n8327 & n8344 ;
  assign n8346 = n8310 & n8345 ;
  assign n8347 = \s5_msel_arb3_state_reg[1]/NET0131  & ~\s5_msel_arb3_state_reg[2]/NET0131  ;
  assign n8348 = ~n4644 & n8347 ;
  assign n8349 = ~n4611 & ~n4623 ;
  assign n8350 = ~n4611 & n4625 ;
  assign n8351 = ~n8349 & ~n8350 ;
  assign n8352 = n8348 & n8351 ;
  assign n8353 = ~n4633 & ~n4651 ;
  assign n8354 = ~n4625 & ~n4635 ;
  assign n8355 = n8348 & n8354 ;
  assign n8356 = ~n8353 & n8355 ;
  assign n8357 = ~n8352 & ~n8356 ;
  assign n8358 = ~n4613 & ~n8357 ;
  assign n8359 = n4628 & ~n4630 ;
  assign n8360 = ~n4633 & ~n8359 ;
  assign n8361 = ~n4635 & ~n8360 ;
  assign n8362 = n8349 & ~n8361 ;
  assign n8363 = ~\s5_msel_arb3_state_reg[0]/NET0131  & \s5_msel_arb3_state_reg[2]/NET0131  ;
  assign n8364 = ~\s5_msel_arb3_state_reg[1]/NET0131  & n8363 ;
  assign n8365 = ~n8350 & n8364 ;
  assign n8366 = ~n4613 & n8365 ;
  assign n8367 = ~n8362 & n8366 ;
  assign n8368 = ~n8358 & ~n8367 ;
  assign n8369 = ~\s5_msel_arb3_state_reg[1]/NET0131  & ~\s5_msel_arb3_state_reg[2]/NET0131  ;
  assign n8370 = \rf_conf5_reg[1]/NET0131  & ~\s5_msel_arb3_state_reg[0]/NET0131  ;
  assign n8371 = n4634 & n8370 ;
  assign n8372 = n8369 & ~n8371 ;
  assign n8373 = ~n8360 & n8372 ;
  assign n8374 = ~n4613 & ~n4630 ;
  assign n8375 = n8372 & n8374 ;
  assign n8376 = n8351 & n8375 ;
  assign n8377 = ~n8373 & ~n8376 ;
  assign n8378 = n4628 & n8348 ;
  assign n8379 = ~\s5_msel_arb3_state_reg[1]/NET0131  & n4616 ;
  assign n8380 = n4611 & n8379 ;
  assign n8381 = ~n8378 & ~n8380 ;
  assign n8382 = n8377 & n8381 ;
  assign n8383 = n8368 & n8382 ;
  assign n8384 = \s5_msel_arb3_state_reg[0]/NET0131  & n8369 ;
  assign n8385 = ~n4635 & n8384 ;
  assign n8386 = n8374 & n8385 ;
  assign n8387 = ~n4611 & n8379 ;
  assign n8388 = ~n8386 & ~n8387 ;
  assign n8389 = ~n4623 & n4635 ;
  assign n8390 = ~n4623 & ~n4633 ;
  assign n8391 = ~n8359 & n8390 ;
  assign n8392 = ~n8389 & ~n8391 ;
  assign n8393 = \s5_msel_arb3_state_reg[0]/NET0131  & ~n4635 ;
  assign n8394 = n8374 & n8393 ;
  assign n8395 = ~n8386 & ~n8394 ;
  assign n8396 = ~n8392 & n8395 ;
  assign n8397 = ~n8388 & ~n8396 ;
  assign n8398 = ~n4625 & n8397 ;
  assign n8399 = ~n4635 & n8374 ;
  assign n8400 = ~\s5_msel_arb3_state_reg[0]/NET0131  & ~n4611 ;
  assign n8401 = n8399 & ~n8400 ;
  assign n8402 = ~n8392 & ~n8401 ;
  assign n8403 = ~\s5_msel_arb3_state_reg[0]/NET0131  & n4625 ;
  assign n8404 = n4625 & n8349 ;
  assign n8405 = n8360 & n8404 ;
  assign n8406 = ~n8403 & ~n8405 ;
  assign n8407 = n4658 & n8406 ;
  assign n8408 = ~n8402 & n8407 ;
  assign n8409 = ~n8398 & ~n8408 ;
  assign n8410 = n8383 & n8409 ;
  assign n8411 = ~n3256 & n3269 ;
  assign n8412 = n3251 & ~n3253 ;
  assign n8413 = ~n3248 & n8412 ;
  assign n8414 = ~n3253 & ~n3258 ;
  assign n8415 = \s6_msel_arb0_state_reg[0]/NET0131  & ~n3248 ;
  assign n8416 = n8414 & n8415 ;
  assign n8417 = ~n8413 & ~n8416 ;
  assign n8418 = n3248 & ~n3263 ;
  assign n8419 = ~n3246 & ~n3263 ;
  assign n8420 = ~n8418 & ~n8419 ;
  assign n8421 = ~n3256 & ~n8420 ;
  assign n8422 = n8417 & n8421 ;
  assign n8423 = ~n8411 & ~n8422 ;
  assign n8424 = n3292 & n8423 ;
  assign n8425 = \s6_msel_arb0_state_reg[1]/NET0131  & \s6_msel_arb0_state_reg[2]/NET0131  ;
  assign n8426 = n3263 & ~n3269 ;
  assign n8427 = ~n3256 & ~n8426 ;
  assign n8428 = ~n3258 & ~n8427 ;
  assign n8429 = ~n3248 & ~n3269 ;
  assign n8430 = ~\s6_msel_arb0_state_reg[0]/NET0131  & ~n3246 ;
  assign n8431 = n8429 & ~n8430 ;
  assign n8432 = ~n3246 & n3253 ;
  assign n8433 = ~n3258 & ~n8432 ;
  assign n8434 = n8431 & n8433 ;
  assign n8435 = ~n8428 & ~n8434 ;
  assign n8436 = ~n3251 & n8435 ;
  assign n8437 = n8425 & ~n8436 ;
  assign n8438 = n3256 & ~n3258 ;
  assign n8439 = ~n3246 & ~n3251 ;
  assign n8440 = ~n8438 & n8439 ;
  assign n8441 = ~n8432 & ~n8440 ;
  assign n8442 = \s6_msel_arb0_state_reg[0]/NET0131  & ~n3269 ;
  assign n8443 = n8414 & n8442 ;
  assign n8444 = ~n3263 & ~n8443 ;
  assign n8445 = ~n8441 & n8444 ;
  assign n8446 = \s6_msel_arb0_state_reg[1]/NET0131  & ~\s6_msel_arb0_state_reg[2]/NET0131  ;
  assign n8447 = ~n8418 & n8446 ;
  assign n8448 = ~n8445 & n8447 ;
  assign n8449 = ~n8437 & ~n8448 ;
  assign n8450 = ~n8424 & n8449 ;
  assign n8451 = \s6_msel_arb0_state_reg[0]/NET0131  & ~n8450 ;
  assign n8452 = \s6_msel_arb0_state_reg[0]/NET0131  & n8414 ;
  assign n8453 = n8429 & n8452 ;
  assign n8454 = n8429 & ~n8432 ;
  assign n8455 = ~n8440 & n8454 ;
  assign n8456 = ~n8453 & ~n8455 ;
  assign n8457 = ~n8426 & n8456 ;
  assign n8458 = n8446 & ~n8457 ;
  assign n8459 = n8412 & n8425 ;
  assign n8460 = n8427 & ~n8431 ;
  assign n8461 = n8414 & n8425 ;
  assign n8462 = ~n8460 & n8461 ;
  assign n8463 = ~n8459 & ~n8462 ;
  assign n8464 = n3292 & n8438 ;
  assign n8465 = ~n3248 & ~n3253 ;
  assign n8466 = ~\s6_msel_arb0_state_reg[0]/NET0131  & ~n3251 ;
  assign n8467 = n8465 & ~n8466 ;
  assign n8468 = ~n8420 & ~n8467 ;
  assign n8469 = ~n3258 & ~n3269 ;
  assign n8470 = n3292 & n8469 ;
  assign n8471 = ~n8468 & n8470 ;
  assign n8472 = ~n8464 & ~n8471 ;
  assign n8473 = n8463 & n8472 ;
  assign n8474 = ~n8458 & n8473 ;
  assign n8475 = ~\s6_msel_arb0_state_reg[0]/NET0131  & ~n8474 ;
  assign n8476 = \s6_msel_arb0_state_reg[0]/NET0131  & n8469 ;
  assign n8477 = n8465 & n8476 ;
  assign n8478 = n3296 & n8477 ;
  assign n8479 = n3263 & n8469 ;
  assign n8480 = n8440 & ~n8479 ;
  assign n8481 = ~\rf_conf6_reg[9]/NET0131  & ~\s6_msel_arb0_state_reg[0]/NET0131  ;
  assign n8482 = n3247 & n8481 ;
  assign n8483 = ~n8432 & ~n8482 ;
  assign n8484 = n3296 & n8483 ;
  assign n8485 = ~n8480 & n8484 ;
  assign n8486 = ~n8478 & ~n8485 ;
  assign n8487 = ~n8475 & n8486 ;
  assign n8488 = ~n8451 & n8487 ;
  assign n8489 = ~n5277 & ~n5281 ;
  assign n8490 = n5278 & ~n5281 ;
  assign n8491 = ~n8489 & ~n8490 ;
  assign n8492 = ~\rf_conf6_reg[9]/NET0131  & ~\s6_msel_arb1_state_reg[0]/NET0131  ;
  assign n8493 = n4666 & n8492 ;
  assign n8494 = n5291 & ~n8493 ;
  assign n8495 = n8491 & n8494 ;
  assign n8496 = n5270 & ~n5273 ;
  assign n8497 = ~n5269 & ~n5273 ;
  assign n8498 = ~n8496 & ~n8497 ;
  assign n8499 = ~n5270 & ~n5280 ;
  assign n8500 = \s6_msel_arb1_state_reg[0]/NET0131  & n8499 ;
  assign n8501 = ~n8498 & ~n8500 ;
  assign n8502 = ~n5272 & ~n5278 ;
  assign n8503 = n8494 & n8502 ;
  assign n8504 = ~n8501 & n8503 ;
  assign n8505 = ~n8495 & ~n8504 ;
  assign n8506 = ~n8496 & n8502 ;
  assign n8507 = ~n8491 & ~n8506 ;
  assign n8508 = ~n5280 & ~n8507 ;
  assign n8509 = ~n5269 & ~n8508 ;
  assign n8510 = \s6_msel_arb1_state_reg[0]/NET0131  & n5297 ;
  assign n8511 = n8489 & n8497 ;
  assign n8512 = ~n5270 & n5297 ;
  assign n8513 = ~n8511 & n8512 ;
  assign n8514 = ~n8510 & ~n8513 ;
  assign n8515 = ~n8509 & ~n8514 ;
  assign n8516 = n8505 & ~n8515 ;
  assign n8517 = ~\rf_conf6_reg[1]/NET0131  & ~\s6_msel_arb1_state_reg[0]/NET0131  ;
  assign n8518 = n4688 & n8517 ;
  assign n8519 = n8498 & ~n8518 ;
  assign n8520 = n8499 & ~n8518 ;
  assign n8521 = n8491 & n8520 ;
  assign n8522 = ~n8519 & ~n8521 ;
  assign n8523 = n8500 & n8502 ;
  assign n8524 = n8522 & ~n8523 ;
  assign n8525 = n5284 & ~n8524 ;
  assign n8526 = n5281 & n8499 ;
  assign n8527 = ~n8498 & ~n8526 ;
  assign n8528 = ~n5272 & ~n8527 ;
  assign n8529 = ~n5277 & ~n8523 ;
  assign n8530 = ~n8528 & n8529 ;
  assign n8531 = ~\rf_conf6_reg[13]/NET0131  & ~\s6_msel_arb1_state_reg[0]/NET0131  ;
  assign n8532 = n4678 & n8531 ;
  assign n8533 = \s6_msel_arb1_state_reg[1]/NET0131  & \s6_msel_arb1_state_reg[2]/NET0131  ;
  assign n8534 = ~n8532 & n8533 ;
  assign n8535 = ~n8530 & n8534 ;
  assign n8536 = ~n8525 & ~n8535 ;
  assign n8537 = n8516 & n8536 ;
  assign n8538 = ~\s6_msel_arb2_state_reg[1]/NET0131  & \s6_msel_arb2_state_reg[2]/NET0131  ;
  assign n8539 = ~n4089 & n8538 ;
  assign n8540 = n4088 & n8539 ;
  assign n8541 = ~n4092 & n4109 ;
  assign n8542 = n4095 & ~n4098 ;
  assign n8543 = ~n4092 & ~n4103 ;
  assign n8544 = ~n8542 & n8543 ;
  assign n8545 = ~n8541 & ~n8544 ;
  assign n8546 = ~n4091 & n8539 ;
  assign n8547 = n8545 & n8546 ;
  assign n8548 = ~n8540 & ~n8547 ;
  assign n8549 = ~\s6_msel_arb2_state_reg[0]/NET0131  & ~n8548 ;
  assign n8550 = ~n4089 & ~n4098 ;
  assign n8551 = ~n8542 & ~n8550 ;
  assign n8552 = ~n4091 & n4092 ;
  assign n8553 = ~n4088 & ~n8552 ;
  assign n8554 = ~n4091 & ~n4109 ;
  assign n8555 = n4103 & n8554 ;
  assign n8556 = n8553 & ~n8555 ;
  assign n8557 = \s6_msel_arb2_state_reg[0]/NET0131  & n8554 ;
  assign n8558 = ~n8542 & ~n8557 ;
  assign n8559 = n8556 & n8558 ;
  assign n8560 = ~n8551 & ~n8559 ;
  assign n8561 = \s6_msel_arb2_state_reg[1]/NET0131  & ~\s6_msel_arb2_state_reg[2]/NET0131  ;
  assign n8562 = ~\s6_msel_arb2_state_reg[0]/NET0131  & n8561 ;
  assign n8563 = n8560 & n8562 ;
  assign n8564 = ~n8549 & ~n8563 ;
  assign n8565 = \s6_msel_arb2_state_reg[0]/NET0131  & ~n4091 ;
  assign n8566 = ~n4088 & ~n8565 ;
  assign n8567 = ~n4109 & n8550 ;
  assign n8568 = ~n8566 & n8567 ;
  assign n8569 = ~n8545 & ~n8568 ;
  assign n8570 = \rf_conf6_reg[13]/NET0131  & ~\s6_msel_arb2_state_reg[0]/NET0131  ;
  assign n8571 = n3252 & n8570 ;
  assign n8572 = \s6_msel_arb2_state_reg[1]/NET0131  & \s6_msel_arb2_state_reg[2]/NET0131  ;
  assign n8573 = ~n8571 & n8572 ;
  assign n8574 = ~n8569 & n8573 ;
  assign n8575 = ~n4089 & ~n8556 ;
  assign n8576 = n8550 & n8557 ;
  assign n8577 = ~n4095 & ~n8576 ;
  assign n8578 = ~n8575 & n8577 ;
  assign n8579 = \s6_msel_arb2_state_reg[0]/NET0131  & n8561 ;
  assign n8580 = ~n8578 & n8579 ;
  assign n8581 = ~n8574 & ~n8580 ;
  assign n8582 = \s6_msel_arb2_state_reg[0]/NET0131  & ~\s6_msel_arb2_state_reg[1]/NET0131  ;
  assign n8583 = \s6_msel_arb2_state_reg[2]/NET0131  & n8582 ;
  assign n8584 = ~n4091 & n8545 ;
  assign n8585 = ~n4088 & ~n8576 ;
  assign n8586 = ~n8584 & n8585 ;
  assign n8587 = n8583 & ~n8586 ;
  assign n8588 = ~n4103 & ~n8542 ;
  assign n8589 = \rf_conf6_reg[1]/NET0131  & ~\s6_msel_arb2_state_reg[0]/NET0131  ;
  assign n8590 = n3257 & n8589 ;
  assign n8591 = ~n8588 & ~n8590 ;
  assign n8592 = n8550 & ~n8590 ;
  assign n8593 = ~n8553 & n8592 ;
  assign n8594 = ~n8591 & ~n8593 ;
  assign n8595 = ~n8576 & n8594 ;
  assign n8596 = ~\s6_msel_arb2_state_reg[1]/NET0131  & ~\s6_msel_arb2_state_reg[2]/NET0131  ;
  assign n8597 = ~n8595 & n8596 ;
  assign n8598 = ~n8587 & ~n8597 ;
  assign n8599 = n8581 & n8598 ;
  assign n8600 = n8564 & n8599 ;
  assign n8601 = \s6_msel_arb3_state_reg[1]/NET0131  & ~\s6_msel_arb3_state_reg[2]/NET0131  ;
  assign n8602 = ~n4698 & n8601 ;
  assign n8603 = ~n4665 & ~n4677 ;
  assign n8604 = ~n4665 & n4679 ;
  assign n8605 = ~n8603 & ~n8604 ;
  assign n8606 = n8602 & n8605 ;
  assign n8607 = ~n4687 & ~n4705 ;
  assign n8608 = ~n4679 & ~n4689 ;
  assign n8609 = n8602 & n8608 ;
  assign n8610 = ~n8607 & n8609 ;
  assign n8611 = ~n8606 & ~n8610 ;
  assign n8612 = ~n4667 & ~n8611 ;
  assign n8613 = n4682 & ~n4684 ;
  assign n8614 = ~n4687 & ~n8613 ;
  assign n8615 = ~n4689 & ~n8614 ;
  assign n8616 = n8603 & ~n8615 ;
  assign n8617 = ~\s6_msel_arb3_state_reg[0]/NET0131  & \s6_msel_arb3_state_reg[2]/NET0131  ;
  assign n8618 = ~\s6_msel_arb3_state_reg[1]/NET0131  & n8617 ;
  assign n8619 = ~n8604 & n8618 ;
  assign n8620 = ~n4667 & n8619 ;
  assign n8621 = ~n8616 & n8620 ;
  assign n8622 = ~n8612 & ~n8621 ;
  assign n8623 = ~\s6_msel_arb3_state_reg[1]/NET0131  & ~\s6_msel_arb3_state_reg[2]/NET0131  ;
  assign n8624 = \rf_conf6_reg[1]/NET0131  & ~\s6_msel_arb3_state_reg[0]/NET0131  ;
  assign n8625 = n4688 & n8624 ;
  assign n8626 = n8623 & ~n8625 ;
  assign n8627 = ~n8614 & n8626 ;
  assign n8628 = ~n4667 & ~n4684 ;
  assign n8629 = n8626 & n8628 ;
  assign n8630 = n8605 & n8629 ;
  assign n8631 = ~n8627 & ~n8630 ;
  assign n8632 = n4682 & n8602 ;
  assign n8633 = ~\s6_msel_arb3_state_reg[1]/NET0131  & n4670 ;
  assign n8634 = n4665 & n8633 ;
  assign n8635 = ~n8632 & ~n8634 ;
  assign n8636 = n8631 & n8635 ;
  assign n8637 = n8622 & n8636 ;
  assign n8638 = \s6_msel_arb3_state_reg[0]/NET0131  & n8623 ;
  assign n8639 = ~n4689 & n8638 ;
  assign n8640 = n8628 & n8639 ;
  assign n8641 = ~n4665 & n8633 ;
  assign n8642 = ~n8640 & ~n8641 ;
  assign n8643 = ~n4677 & n4689 ;
  assign n8644 = ~n4677 & ~n4687 ;
  assign n8645 = ~n8613 & n8644 ;
  assign n8646 = ~n8643 & ~n8645 ;
  assign n8647 = \s6_msel_arb3_state_reg[0]/NET0131  & ~n4689 ;
  assign n8648 = n8628 & n8647 ;
  assign n8649 = ~n8640 & ~n8648 ;
  assign n8650 = ~n8646 & n8649 ;
  assign n8651 = ~n8642 & ~n8650 ;
  assign n8652 = ~n4679 & n8651 ;
  assign n8653 = ~n4689 & n8628 ;
  assign n8654 = ~\s6_msel_arb3_state_reg[0]/NET0131  & ~n4665 ;
  assign n8655 = n8653 & ~n8654 ;
  assign n8656 = ~n8646 & ~n8655 ;
  assign n8657 = ~\s6_msel_arb3_state_reg[0]/NET0131  & n4679 ;
  assign n8658 = n4679 & n8603 ;
  assign n8659 = n8614 & n8658 ;
  assign n8660 = ~n8657 & ~n8659 ;
  assign n8661 = n4712 & n8660 ;
  assign n8662 = ~n8656 & n8661 ;
  assign n8663 = ~n8652 & ~n8662 ;
  assign n8664 = n8637 & n8663 ;
  assign n8665 = ~n3506 & n3515 ;
  assign n8666 = n3496 & ~n3498 ;
  assign n8667 = ~n3506 & ~n3513 ;
  assign n8668 = ~n8666 & n8667 ;
  assign n8669 = ~n8665 & ~n8668 ;
  assign n8670 = ~n3498 & ~n3515 ;
  assign n8671 = ~n3501 & n8670 ;
  assign n8672 = ~n3503 & n3508 ;
  assign n8673 = ~\s7_msel_arb0_state_reg[0]/NET0131  & ~n3503 ;
  assign n8674 = ~n8672 & ~n8673 ;
  assign n8675 = n8671 & n8674 ;
  assign n8676 = ~n8669 & ~n8675 ;
  assign n8677 = n3549 & ~n8676 ;
  assign n8678 = ~n3503 & ~n3506 ;
  assign n8679 = ~n8672 & ~n8678 ;
  assign n8680 = ~\s7_msel_arb0_state_reg[1]/NET0131  & \s7_msel_arb0_state_reg[2]/NET0131  ;
  assign n8681 = ~\rf_conf7_reg[3]/NET0131  & ~\s7_msel_arb0_state_reg[1]/NET0131  ;
  assign n8682 = n3512 & n8681 ;
  assign n8683 = ~n8680 & ~n8682 ;
  assign n8684 = n8679 & ~n8683 ;
  assign n8685 = ~n3496 & n3501 ;
  assign n8686 = ~n3498 & ~n8685 ;
  assign n8687 = ~n3513 & ~n8686 ;
  assign n8688 = ~n3508 & ~n3515 ;
  assign n8689 = \s7_msel_arb0_state_reg[2]/NET0131  & ~n8688 ;
  assign n8690 = ~n8683 & ~n8689 ;
  assign n8691 = ~n8687 & n8690 ;
  assign n8692 = ~n8684 & ~n8691 ;
  assign n8693 = ~n8677 & n8692 ;
  assign n8694 = \s7_msel_arb0_state_reg[0]/NET0131  & ~n8693 ;
  assign n8695 = \s7_msel_arb0_state_reg[0]/NET0131  & n8688 ;
  assign n8696 = ~n3498 & ~n3501 ;
  assign n8697 = n8695 & n8696 ;
  assign n8698 = n3543 & n8697 ;
  assign n8699 = n3513 & n8688 ;
  assign n8700 = ~n3496 & ~n8679 ;
  assign n8701 = ~n8699 & n8700 ;
  assign n8702 = ~\rf_conf7_reg[5]/NET0131  & ~\s7_msel_arb0_state_reg[0]/NET0131  ;
  assign n8703 = n3497 & n8702 ;
  assign n8704 = ~n8685 & ~n8703 ;
  assign n8705 = n3543 & n8704 ;
  assign n8706 = ~n8701 & n8705 ;
  assign n8707 = ~n8698 & ~n8706 ;
  assign n8708 = ~n3513 & ~n8666 ;
  assign n8709 = ~n3515 & ~n8708 ;
  assign n8710 = ~n3501 & ~n3508 ;
  assign n8711 = \s7_msel_arb0_state_reg[2]/NET0131  & ~n8710 ;
  assign n8712 = n8709 & ~n8711 ;
  assign n8713 = ~\s7_msel_arb0_state_reg[2]/NET0131  & ~n8670 ;
  assign n8714 = ~n3501 & n8679 ;
  assign n8715 = ~n8713 & n8714 ;
  assign n8716 = ~n8712 & ~n8715 ;
  assign n8717 = ~\s7_msel_arb0_state_reg[0]/NET0131  & ~\s7_msel_arb0_state_reg[1]/NET0131  ;
  assign n8718 = ~n8716 & n8717 ;
  assign n8719 = ~n8695 & n8700 ;
  assign n8720 = ~\s7_msel_arb0_state_reg[1]/NET0131  & ~\s7_msel_arb0_state_reg[2]/NET0131  ;
  assign n8721 = \s7_msel_arb0_state_reg[0]/NET0131  & n8720 ;
  assign n8722 = ~n3513 & n8721 ;
  assign n8723 = n8686 & n8722 ;
  assign n8724 = ~n8719 & n8723 ;
  assign n8725 = n8671 & ~n8673 ;
  assign n8726 = ~n8669 & ~n8725 ;
  assign n8727 = \s7_msel_arb0_state_reg[2]/NET0131  & n3532 ;
  assign n8728 = ~n3508 & n8727 ;
  assign n8729 = ~n8726 & n8728 ;
  assign n8730 = ~n8724 & ~n8729 ;
  assign n8731 = ~n8718 & n8730 ;
  assign n8732 = n8707 & n8731 ;
  assign n8733 = ~n8694 & n8732 ;
  assign n8734 = n5315 & ~n5316 ;
  assign n8735 = ~n5312 & ~n8734 ;
  assign n8736 = ~n5316 & ~n5320 ;
  assign n8737 = n5319 & n8736 ;
  assign n8738 = n8735 & ~n8737 ;
  assign n8739 = ~n5313 & ~n8738 ;
  assign n8740 = ~n5313 & ~n5323 ;
  assign n8741 = n8736 & n8740 ;
  assign n8742 = \s7_msel_arb1_state_reg[2]/NET0131  & ~n8741 ;
  assign n8743 = ~n5322 & n8742 ;
  assign n8744 = ~n8739 & n8743 ;
  assign n8745 = ~\s7_msel_arb1_state_reg[2]/NET0131  & ~n5315 ;
  assign n8746 = n5343 & ~n8745 ;
  assign n8747 = \s7_msel_arb1_state_reg[0]/NET0131  & ~n5313 ;
  assign n8748 = ~n5316 & n8747 ;
  assign n8749 = ~n5319 & ~n5322 ;
  assign n8750 = n5312 & ~n5313 ;
  assign n8751 = n8749 & ~n8750 ;
  assign n8752 = ~n8748 & n8751 ;
  assign n8753 = ~n5319 & n5323 ;
  assign n8754 = ~n5320 & ~n8753 ;
  assign n8755 = n5343 & n8754 ;
  assign n8756 = ~n8752 & n8755 ;
  assign n8757 = ~n8746 & ~n8756 ;
  assign n8758 = ~n8744 & ~n8757 ;
  assign n8759 = ~n5323 & n8736 ;
  assign n8760 = ~n5322 & ~n8747 ;
  assign n8761 = n8759 & ~n8760 ;
  assign n8762 = n8738 & ~n8761 ;
  assign n8763 = ~\s7_msel_arb1_state_reg[1]/NET0131  & ~\s7_msel_arb1_state_reg[2]/NET0131  ;
  assign n8764 = \s7_msel_arb1_state_reg[0]/NET0131  & n8763 ;
  assign n8765 = ~n8762 & n8764 ;
  assign n8766 = ~n5313 & ~n8735 ;
  assign n8767 = n8736 & n8747 ;
  assign n8768 = n8749 & ~n8767 ;
  assign n8769 = ~n8766 & n8768 ;
  assign n8770 = ~\s7_msel_arb1_state_reg[1]/NET0131  & \s7_msel_arb1_state_reg[2]/NET0131  ;
  assign n8771 = \s7_msel_arb1_state_reg[0]/NET0131  & n8770 ;
  assign n8772 = ~n8753 & n8771 ;
  assign n8773 = ~n8769 & n8772 ;
  assign n8774 = ~n8765 & ~n8773 ;
  assign n8775 = ~n8758 & n8774 ;
  assign n8776 = \s7_msel_arb1_state_reg[0]/NET0131  & n8775 ;
  assign n8777 = ~n5316 & ~n8749 ;
  assign n8778 = n8754 & n8777 ;
  assign n8779 = ~n8734 & ~n8778 ;
  assign n8780 = ~\s7_msel_arb1_state_reg[2]/NET0131  & ~n8779 ;
  assign n8781 = \s7_msel_arb1_state_reg[1]/NET0131  & n8780 ;
  assign n8782 = \s7_msel_arb1_state_reg[2]/NET0131  & n5322 ;
  assign n8783 = \s7_msel_arb1_state_reg[2]/NET0131  & ~n5313 ;
  assign n8784 = ~n8738 & n8783 ;
  assign n8785 = ~n8782 & ~n8784 ;
  assign n8786 = ~n8747 & ~n8750 ;
  assign n8787 = ~\s7_msel_arb1_state_reg[2]/NET0131  & n8736 ;
  assign n8788 = ~n8786 & n8787 ;
  assign n8789 = n8785 & ~n8788 ;
  assign n8790 = \s7_msel_arb1_state_reg[1]/NET0131  & ~n5323 ;
  assign n8791 = ~n8789 & n8790 ;
  assign n8792 = ~n8781 & ~n8791 ;
  assign n8793 = ~n8748 & n8749 ;
  assign n8794 = ~n8766 & n8793 ;
  assign n8795 = ~n5320 & n8770 ;
  assign n8796 = ~n8753 & n8795 ;
  assign n8797 = ~n8794 & n8796 ;
  assign n8798 = n8735 & ~n8778 ;
  assign n8799 = ~n5313 & n8763 ;
  assign n8800 = ~n8798 & n8799 ;
  assign n8801 = ~n8797 & ~n8800 ;
  assign n8802 = n8775 & n8801 ;
  assign n8803 = n8792 & n8802 ;
  assign n8804 = ~n8776 & ~n8803 ;
  assign n8805 = \rf_conf7_reg[5]/NET0131  & n3497 ;
  assign n8806 = \rf_conf7_reg[7]/NET0131  & n3495 ;
  assign n8807 = ~n8805 & n8806 ;
  assign n8808 = \s7_msel_arb2_state_reg[1]/NET0131  & ~\s7_msel_arb2_state_reg[2]/NET0131  ;
  assign n8809 = n8807 & n8808 ;
  assign n8810 = \rf_conf7_reg[11]/NET0131  & n3502 ;
  assign n8811 = \rf_conf7_reg[15]/NET0131  & n3505 ;
  assign n8812 = \rf_conf7_reg[13]/NET0131  & n3507 ;
  assign n8813 = n8811 & ~n8812 ;
  assign n8814 = ~n8810 & ~n8813 ;
  assign n8815 = \rf_conf7_reg[3]/NET0131  & n3512 ;
  assign n8816 = \rf_conf7_reg[1]/NET0131  & n3514 ;
  assign n8817 = ~n8812 & ~n8816 ;
  assign n8818 = n8815 & n8817 ;
  assign n8819 = n8814 & ~n8818 ;
  assign n8820 = \rf_conf7_reg[9]/NET0131  & n3500 ;
  assign n8821 = ~n8805 & ~n8820 ;
  assign n8822 = n8808 & n8821 ;
  assign n8823 = ~n8819 & n8822 ;
  assign n8824 = ~n8809 & ~n8823 ;
  assign n8825 = ~n8807 & ~n8815 ;
  assign n8826 = ~\s7_msel_arb2_state_reg[1]/NET0131  & ~\s7_msel_arb2_state_reg[2]/NET0131  ;
  assign n8827 = ~n8816 & n8826 ;
  assign n8828 = ~n8825 & n8827 ;
  assign n8829 = n8821 & n8827 ;
  assign n8830 = ~n8814 & n8829 ;
  assign n8831 = ~n8828 & ~n8830 ;
  assign n8832 = ~\s7_msel_arb2_state_reg[0]/NET0131  & n8831 ;
  assign n8833 = n8824 & n8832 ;
  assign n8834 = \s7_msel_arb2_state_reg[1]/NET0131  & \s7_msel_arb2_state_reg[2]/NET0131  ;
  assign n8835 = n8813 & n8834 ;
  assign n8836 = n8810 & n8821 ;
  assign n8837 = n8825 & ~n8836 ;
  assign n8838 = n8817 & n8834 ;
  assign n8839 = ~n8837 & n8838 ;
  assign n8840 = ~n8835 & ~n8839 ;
  assign n8841 = ~\s7_msel_arb2_state_reg[1]/NET0131  & \s7_msel_arb2_state_reg[2]/NET0131  ;
  assign n8842 = ~n8820 & n8841 ;
  assign n8843 = n8810 & n8842 ;
  assign n8844 = ~n8811 & n8816 ;
  assign n8845 = ~n8811 & ~n8815 ;
  assign n8846 = ~n8807 & n8845 ;
  assign n8847 = ~n8844 & ~n8846 ;
  assign n8848 = ~n8812 & n8842 ;
  assign n8849 = n8847 & n8848 ;
  assign n8850 = ~n8843 & ~n8849 ;
  assign n8851 = n8840 & n8850 ;
  assign n8852 = n8833 & n8851 ;
  assign n8853 = \s7_msel_arb2_state_reg[0]/NET0131  & ~n8816 ;
  assign n8854 = n8821 & n8853 ;
  assign n8855 = ~n8847 & ~n8854 ;
  assign n8856 = \s7_msel_arb2_state_reg[0]/NET0131  & n8841 ;
  assign n8857 = ~n8810 & n8856 ;
  assign n8858 = ~n8812 & n8857 ;
  assign n8859 = ~n8855 & n8858 ;
  assign n8860 = n8852 & ~n8859 ;
  assign n8861 = ~n8814 & n8821 ;
  assign n8862 = n8825 & ~n8861 ;
  assign n8863 = \s7_msel_arb2_state_reg[0]/NET0131  & n8821 ;
  assign n8864 = n8817 & n8863 ;
  assign n8865 = n8862 & ~n8864 ;
  assign n8866 = n8826 & ~n8865 ;
  assign n8867 = n8806 & n8808 ;
  assign n8868 = n8805 & ~n8815 ;
  assign n8869 = n8817 & ~n8868 ;
  assign n8870 = n8814 & ~n8869 ;
  assign n8871 = n8808 & ~n8820 ;
  assign n8872 = ~n8870 & n8871 ;
  assign n8873 = ~n8867 & ~n8872 ;
  assign n8874 = n8810 & n8841 ;
  assign n8875 = \s7_msel_arb2_state_reg[0]/NET0131  & ~n8874 ;
  assign n8876 = n8873 & n8875 ;
  assign n8877 = ~n8866 & n8876 ;
  assign n8878 = \s7_msel_arb2_state_reg[0]/NET0131  & ~n8812 ;
  assign n8879 = n8821 & n8878 ;
  assign n8880 = ~n8811 & ~n8879 ;
  assign n8881 = n8837 & n8880 ;
  assign n8882 = ~n8844 & ~n8881 ;
  assign n8883 = n8834 & n8882 ;
  assign n8884 = ~n8859 & ~n8883 ;
  assign n8885 = n8877 & n8884 ;
  assign n8886 = ~n8860 & ~n8885 ;
  assign n8887 = \s7_msel_arb3_state_reg[1]/NET0131  & ~\s7_msel_arb3_state_reg[2]/NET0131  ;
  assign n8888 = ~n4752 & n8887 ;
  assign n8889 = ~n4719 & ~n4731 ;
  assign n8890 = ~n4719 & n4733 ;
  assign n8891 = ~n8889 & ~n8890 ;
  assign n8892 = n8888 & n8891 ;
  assign n8893 = ~n4741 & ~n4759 ;
  assign n8894 = ~n4733 & ~n4743 ;
  assign n8895 = n8888 & n8894 ;
  assign n8896 = ~n8893 & n8895 ;
  assign n8897 = ~n8892 & ~n8896 ;
  assign n8898 = ~n4721 & ~n8897 ;
  assign n8899 = n4736 & ~n4738 ;
  assign n8900 = ~n4741 & ~n8899 ;
  assign n8901 = ~n4743 & ~n8900 ;
  assign n8902 = n8889 & ~n8901 ;
  assign n8903 = ~\s7_msel_arb3_state_reg[0]/NET0131  & \s7_msel_arb3_state_reg[2]/NET0131  ;
  assign n8904 = ~\s7_msel_arb3_state_reg[1]/NET0131  & n8903 ;
  assign n8905 = ~n8890 & n8904 ;
  assign n8906 = ~n4721 & n8905 ;
  assign n8907 = ~n8902 & n8906 ;
  assign n8908 = ~n8898 & ~n8907 ;
  assign n8909 = ~\s7_msel_arb3_state_reg[1]/NET0131  & ~\s7_msel_arb3_state_reg[2]/NET0131  ;
  assign n8910 = \rf_conf7_reg[1]/NET0131  & ~\s7_msel_arb3_state_reg[0]/NET0131  ;
  assign n8911 = n4742 & n8910 ;
  assign n8912 = n8909 & ~n8911 ;
  assign n8913 = ~n8900 & n8912 ;
  assign n8914 = ~n4721 & ~n4738 ;
  assign n8915 = n8912 & n8914 ;
  assign n8916 = n8891 & n8915 ;
  assign n8917 = ~n8913 & ~n8916 ;
  assign n8918 = n4736 & n8888 ;
  assign n8919 = ~\s7_msel_arb3_state_reg[1]/NET0131  & n4724 ;
  assign n8920 = n4719 & n8919 ;
  assign n8921 = ~n8918 & ~n8920 ;
  assign n8922 = n8917 & n8921 ;
  assign n8923 = n8908 & n8922 ;
  assign n8924 = \s7_msel_arb3_state_reg[0]/NET0131  & n8909 ;
  assign n8925 = ~n4743 & n8924 ;
  assign n8926 = n8914 & n8925 ;
  assign n8927 = ~n4719 & n8919 ;
  assign n8928 = ~n8926 & ~n8927 ;
  assign n8929 = ~n4731 & n4743 ;
  assign n8930 = ~n4731 & ~n4741 ;
  assign n8931 = ~n8899 & n8930 ;
  assign n8932 = ~n8929 & ~n8931 ;
  assign n8933 = \s7_msel_arb3_state_reg[0]/NET0131  & ~n4743 ;
  assign n8934 = n8914 & n8933 ;
  assign n8935 = ~n8926 & ~n8934 ;
  assign n8936 = ~n8932 & n8935 ;
  assign n8937 = ~n8928 & ~n8936 ;
  assign n8938 = ~n4733 & n8937 ;
  assign n8939 = ~n4743 & n8914 ;
  assign n8940 = ~\s7_msel_arb3_state_reg[0]/NET0131  & ~n4719 ;
  assign n8941 = n8939 & ~n8940 ;
  assign n8942 = ~n8932 & ~n8941 ;
  assign n8943 = ~\s7_msel_arb3_state_reg[0]/NET0131  & n4733 ;
  assign n8944 = n4733 & n8889 ;
  assign n8945 = n8900 & n8944 ;
  assign n8946 = ~n8943 & ~n8945 ;
  assign n8947 = n4766 & n8946 ;
  assign n8948 = ~n8942 & n8947 ;
  assign n8949 = ~n8938 & ~n8948 ;
  assign n8950 = n8923 & n8949 ;
  assign n8951 = ~n3318 & n3331 ;
  assign n8952 = n3313 & ~n3315 ;
  assign n8953 = ~n3310 & n8952 ;
  assign n8954 = ~n3315 & ~n3320 ;
  assign n8955 = \s8_msel_arb0_state_reg[0]/NET0131  & ~n3310 ;
  assign n8956 = n8954 & n8955 ;
  assign n8957 = ~n8953 & ~n8956 ;
  assign n8958 = n3310 & ~n3325 ;
  assign n8959 = ~n3308 & ~n3325 ;
  assign n8960 = ~n8958 & ~n8959 ;
  assign n8961 = ~n3318 & ~n8960 ;
  assign n8962 = n8957 & n8961 ;
  assign n8963 = ~n8951 & ~n8962 ;
  assign n8964 = n3354 & n8963 ;
  assign n8965 = \s8_msel_arb0_state_reg[1]/NET0131  & \s8_msel_arb0_state_reg[2]/NET0131  ;
  assign n8966 = n3325 & ~n3331 ;
  assign n8967 = ~n3318 & ~n8966 ;
  assign n8968 = ~n3320 & ~n8967 ;
  assign n8969 = ~n3310 & ~n3331 ;
  assign n8970 = ~\s8_msel_arb0_state_reg[0]/NET0131  & ~n3308 ;
  assign n8971 = n8969 & ~n8970 ;
  assign n8972 = ~n3308 & n3315 ;
  assign n8973 = ~n3320 & ~n8972 ;
  assign n8974 = n8971 & n8973 ;
  assign n8975 = ~n8968 & ~n8974 ;
  assign n8976 = ~n3313 & n8975 ;
  assign n8977 = n8965 & ~n8976 ;
  assign n8978 = n3318 & ~n3320 ;
  assign n8979 = ~n3308 & ~n3313 ;
  assign n8980 = ~n8978 & n8979 ;
  assign n8981 = ~n8972 & ~n8980 ;
  assign n8982 = \s8_msel_arb0_state_reg[0]/NET0131  & ~n3331 ;
  assign n8983 = n8954 & n8982 ;
  assign n8984 = ~n3325 & ~n8983 ;
  assign n8985 = ~n8981 & n8984 ;
  assign n8986 = \s8_msel_arb0_state_reg[1]/NET0131  & ~\s8_msel_arb0_state_reg[2]/NET0131  ;
  assign n8987 = ~n8958 & n8986 ;
  assign n8988 = ~n8985 & n8987 ;
  assign n8989 = ~n8977 & ~n8988 ;
  assign n8990 = ~n8964 & n8989 ;
  assign n8991 = \s8_msel_arb0_state_reg[0]/NET0131  & ~n8990 ;
  assign n8992 = \s8_msel_arb0_state_reg[0]/NET0131  & n8954 ;
  assign n8993 = n8969 & n8992 ;
  assign n8994 = n8969 & ~n8972 ;
  assign n8995 = ~n8980 & n8994 ;
  assign n8996 = ~n8993 & ~n8995 ;
  assign n8997 = ~n8966 & n8996 ;
  assign n8998 = n8986 & ~n8997 ;
  assign n8999 = n8952 & n8965 ;
  assign n9000 = n8967 & ~n8971 ;
  assign n9001 = n8954 & n8965 ;
  assign n9002 = ~n9000 & n9001 ;
  assign n9003 = ~n8999 & ~n9002 ;
  assign n9004 = n3354 & n8978 ;
  assign n9005 = ~n3310 & ~n3315 ;
  assign n9006 = ~\s8_msel_arb0_state_reg[0]/NET0131  & ~n3313 ;
  assign n9007 = n9005 & ~n9006 ;
  assign n9008 = ~n8960 & ~n9007 ;
  assign n9009 = ~n3320 & ~n3331 ;
  assign n9010 = n3354 & n9009 ;
  assign n9011 = ~n9008 & n9010 ;
  assign n9012 = ~n9004 & ~n9011 ;
  assign n9013 = n9003 & n9012 ;
  assign n9014 = ~n8998 & n9013 ;
  assign n9015 = ~\s8_msel_arb0_state_reg[0]/NET0131  & ~n9014 ;
  assign n9016 = \s8_msel_arb0_state_reg[0]/NET0131  & n9009 ;
  assign n9017 = n9005 & n9016 ;
  assign n9018 = n3358 & n9017 ;
  assign n9019 = n3325 & n9009 ;
  assign n9020 = n8980 & ~n9019 ;
  assign n9021 = ~\rf_conf8_reg[9]/NET0131  & ~\s8_msel_arb0_state_reg[0]/NET0131  ;
  assign n9022 = n3309 & n9021 ;
  assign n9023 = ~n8972 & ~n9022 ;
  assign n9024 = n3358 & n9023 ;
  assign n9025 = ~n9020 & n9024 ;
  assign n9026 = ~n9018 & ~n9025 ;
  assign n9027 = ~n9015 & n9026 ;
  assign n9028 = ~n8991 & n9027 ;
  assign n9029 = ~n5358 & ~n5362 ;
  assign n9030 = n5359 & ~n5362 ;
  assign n9031 = ~n9029 & ~n9030 ;
  assign n9032 = ~\rf_conf8_reg[9]/NET0131  & ~\s8_msel_arb1_state_reg[0]/NET0131  ;
  assign n9033 = n4797 & n9032 ;
  assign n9034 = n5372 & ~n9033 ;
  assign n9035 = n9031 & n9034 ;
  assign n9036 = n5351 & ~n5354 ;
  assign n9037 = ~n5350 & ~n5354 ;
  assign n9038 = ~n9036 & ~n9037 ;
  assign n9039 = ~n5351 & ~n5361 ;
  assign n9040 = \s8_msel_arb1_state_reg[0]/NET0131  & n9039 ;
  assign n9041 = ~n9038 & ~n9040 ;
  assign n9042 = ~n5353 & ~n5359 ;
  assign n9043 = n9034 & n9042 ;
  assign n9044 = ~n9041 & n9043 ;
  assign n9045 = ~n9035 & ~n9044 ;
  assign n9046 = ~n9036 & n9042 ;
  assign n9047 = ~n9031 & ~n9046 ;
  assign n9048 = ~n5361 & ~n9047 ;
  assign n9049 = ~n5350 & ~n9048 ;
  assign n9050 = \s8_msel_arb1_state_reg[0]/NET0131  & n5378 ;
  assign n9051 = n9029 & n9037 ;
  assign n9052 = ~n5351 & n5378 ;
  assign n9053 = ~n9051 & n9052 ;
  assign n9054 = ~n9050 & ~n9053 ;
  assign n9055 = ~n9049 & ~n9054 ;
  assign n9056 = n9045 & ~n9055 ;
  assign n9057 = ~\rf_conf8_reg[1]/NET0131  & ~\s8_msel_arb1_state_reg[0]/NET0131  ;
  assign n9058 = n4775 & n9057 ;
  assign n9059 = n9038 & ~n9058 ;
  assign n9060 = n9039 & ~n9058 ;
  assign n9061 = n9031 & n9060 ;
  assign n9062 = ~n9059 & ~n9061 ;
  assign n9063 = n9040 & n9042 ;
  assign n9064 = n9062 & ~n9063 ;
  assign n9065 = n5365 & ~n9064 ;
  assign n9066 = n5362 & n9039 ;
  assign n9067 = ~n9038 & ~n9066 ;
  assign n9068 = ~n5353 & ~n9067 ;
  assign n9069 = ~n5358 & ~n9063 ;
  assign n9070 = ~n9068 & n9069 ;
  assign n9071 = ~\rf_conf8_reg[13]/NET0131  & ~\s8_msel_arb1_state_reg[0]/NET0131  ;
  assign n9072 = n4788 & n9071 ;
  assign n9073 = \s8_msel_arb1_state_reg[1]/NET0131  & \s8_msel_arb1_state_reg[2]/NET0131  ;
  assign n9074 = ~n9072 & n9073 ;
  assign n9075 = ~n9070 & n9074 ;
  assign n9076 = ~n9065 & ~n9075 ;
  assign n9077 = n9056 & n9076 ;
  assign n9078 = ~\s8_msel_arb2_state_reg[1]/NET0131  & \s8_msel_arb2_state_reg[2]/NET0131  ;
  assign n9079 = ~n4124 & n9078 ;
  assign n9080 = n4123 & n9079 ;
  assign n9081 = ~n4127 & n4144 ;
  assign n9082 = n4130 & ~n4133 ;
  assign n9083 = ~n4127 & ~n4138 ;
  assign n9084 = ~n9082 & n9083 ;
  assign n9085 = ~n9081 & ~n9084 ;
  assign n9086 = ~n4126 & n9079 ;
  assign n9087 = n9085 & n9086 ;
  assign n9088 = ~n9080 & ~n9087 ;
  assign n9089 = ~\s8_msel_arb2_state_reg[0]/NET0131  & ~n9088 ;
  assign n9090 = ~n4124 & ~n4133 ;
  assign n9091 = ~n9082 & ~n9090 ;
  assign n9092 = ~n4126 & n4127 ;
  assign n9093 = ~n4123 & ~n9092 ;
  assign n9094 = ~n4126 & ~n4144 ;
  assign n9095 = n4138 & n9094 ;
  assign n9096 = n9093 & ~n9095 ;
  assign n9097 = \s8_msel_arb2_state_reg[0]/NET0131  & n9094 ;
  assign n9098 = ~n9082 & ~n9097 ;
  assign n9099 = n9096 & n9098 ;
  assign n9100 = ~n9091 & ~n9099 ;
  assign n9101 = \s8_msel_arb2_state_reg[1]/NET0131  & ~\s8_msel_arb2_state_reg[2]/NET0131  ;
  assign n9102 = ~\s8_msel_arb2_state_reg[0]/NET0131  & n9101 ;
  assign n9103 = n9100 & n9102 ;
  assign n9104 = ~n9089 & ~n9103 ;
  assign n9105 = \s8_msel_arb2_state_reg[0]/NET0131  & ~n4126 ;
  assign n9106 = ~n4123 & ~n9105 ;
  assign n9107 = ~n4144 & n9090 ;
  assign n9108 = ~n9106 & n9107 ;
  assign n9109 = ~n9085 & ~n9108 ;
  assign n9110 = \rf_conf8_reg[13]/NET0131  & ~\s8_msel_arb2_state_reg[0]/NET0131  ;
  assign n9111 = n3314 & n9110 ;
  assign n9112 = \s8_msel_arb2_state_reg[1]/NET0131  & \s8_msel_arb2_state_reg[2]/NET0131  ;
  assign n9113 = ~n9111 & n9112 ;
  assign n9114 = ~n9109 & n9113 ;
  assign n9115 = ~n4124 & ~n9096 ;
  assign n9116 = n9090 & n9097 ;
  assign n9117 = ~n4130 & ~n9116 ;
  assign n9118 = ~n9115 & n9117 ;
  assign n9119 = \s8_msel_arb2_state_reg[0]/NET0131  & n9101 ;
  assign n9120 = ~n9118 & n9119 ;
  assign n9121 = ~n9114 & ~n9120 ;
  assign n9122 = \s8_msel_arb2_state_reg[0]/NET0131  & ~\s8_msel_arb2_state_reg[1]/NET0131  ;
  assign n9123 = \s8_msel_arb2_state_reg[2]/NET0131  & n9122 ;
  assign n9124 = ~n4126 & n9085 ;
  assign n9125 = ~n4123 & ~n9116 ;
  assign n9126 = ~n9124 & n9125 ;
  assign n9127 = n9123 & ~n9126 ;
  assign n9128 = ~n4138 & ~n9082 ;
  assign n9129 = \rf_conf8_reg[1]/NET0131  & ~\s8_msel_arb2_state_reg[0]/NET0131  ;
  assign n9130 = n3319 & n9129 ;
  assign n9131 = ~n9128 & ~n9130 ;
  assign n9132 = n9090 & ~n9130 ;
  assign n9133 = ~n9093 & n9132 ;
  assign n9134 = ~n9131 & ~n9133 ;
  assign n9135 = ~n9116 & n9134 ;
  assign n9136 = ~\s8_msel_arb2_state_reg[1]/NET0131  & ~\s8_msel_arb2_state_reg[2]/NET0131  ;
  assign n9137 = ~n9135 & n9136 ;
  assign n9138 = ~n9127 & ~n9137 ;
  assign n9139 = n9121 & n9138 ;
  assign n9140 = n9104 & n9139 ;
  assign n9141 = ~n4781 & ~n4798 ;
  assign n9142 = n4779 & ~n4781 ;
  assign n9143 = ~n9141 & ~n9142 ;
  assign n9144 = ~n4785 & n4789 ;
  assign n9145 = n4774 & ~n4776 ;
  assign n9146 = ~n4785 & ~n4787 ;
  assign n9147 = ~n9145 & n9146 ;
  assign n9148 = ~n9144 & ~n9147 ;
  assign n9149 = \s8_msel_arb3_state_reg[0]/NET0131  & ~n4789 ;
  assign n9150 = ~n4776 & n9149 ;
  assign n9151 = ~n9142 & ~n9150 ;
  assign n9152 = ~n9148 & n9151 ;
  assign n9153 = ~n9143 & ~n9152 ;
  assign n9154 = n4815 & n9153 ;
  assign n9155 = ~\s8_msel_arb3_state_reg[1]/NET0131  & ~\s8_msel_arb3_state_reg[2]/NET0131  ;
  assign n9156 = n9145 & n9155 ;
  assign n9157 = ~n4779 & n4798 ;
  assign n9158 = n4787 & ~n4789 ;
  assign n9159 = ~n4779 & ~n4785 ;
  assign n9160 = ~n9158 & n9159 ;
  assign n9161 = ~n9157 & ~n9160 ;
  assign n9162 = ~n4776 & ~n4781 ;
  assign n9163 = n9155 & n9162 ;
  assign n9164 = n9161 & n9163 ;
  assign n9165 = ~n9156 & ~n9164 ;
  assign n9166 = n4772 & ~n4798 ;
  assign n9167 = n4785 & n9166 ;
  assign n9168 = ~n4787 & ~n9145 ;
  assign n9169 = ~n4776 & n9142 ;
  assign n9170 = n9168 & ~n9169 ;
  assign n9171 = ~n4789 & n9166 ;
  assign n9172 = ~n9170 & n9171 ;
  assign n9173 = ~n9167 & ~n9172 ;
  assign n9174 = ~\s8_msel_arb3_state_reg[0]/NET0131  & n9173 ;
  assign n9175 = n9165 & n9174 ;
  assign n9176 = ~n9154 & n9175 ;
  assign n9177 = ~n4789 & ~n9170 ;
  assign n9178 = ~n4776 & ~n4789 ;
  assign n9179 = n9141 & n9178 ;
  assign n9180 = ~n4785 & ~n9179 ;
  assign n9181 = ~n9177 & n9180 ;
  assign n9182 = n4772 & ~n9181 ;
  assign n9183 = n4779 & n4815 ;
  assign n9184 = \s8_msel_arb3_state_reg[0]/NET0131  & ~n9183 ;
  assign n9185 = ~n9182 & n9184 ;
  assign n9186 = ~n9176 & ~n9185 ;
  assign n9187 = ~n4774 & n4781 ;
  assign n9188 = ~n4776 & ~n4798 ;
  assign n9189 = n9149 & n9188 ;
  assign n9190 = ~n4774 & ~n9189 ;
  assign n9191 = ~n9161 & n9190 ;
  assign n9192 = ~n9187 & ~n9191 ;
  assign n9193 = \s8_msel_arb3_state_reg[0]/NET0131  & n9155 ;
  assign n9194 = n9192 & n9193 ;
  assign n9195 = ~n4785 & ~n9149 ;
  assign n9196 = ~n4776 & n9141 ;
  assign n9197 = ~n9195 & n9196 ;
  assign n9198 = n9170 & ~n9197 ;
  assign n9199 = \rf_conf8_reg[13]/NET0131  & ~\s8_msel_arb3_state_reg[0]/NET0131  ;
  assign n9200 = n4788 & n9199 ;
  assign n9201 = n4795 & ~n9200 ;
  assign n9202 = ~n9198 & n9201 ;
  assign n9203 = n9149 & n9162 ;
  assign n9204 = ~n9148 & ~n9203 ;
  assign n9205 = \s8_msel_arb3_state_reg[0]/NET0131  & n4815 ;
  assign n9206 = ~n4779 & n9205 ;
  assign n9207 = ~n4798 & n9206 ;
  assign n9208 = ~n9204 & n9207 ;
  assign n9209 = ~n9202 & ~n9208 ;
  assign n9210 = ~n9194 & n9209 ;
  assign n9211 = ~n9186 & n9210 ;
  assign n9212 = ~n3569 & n3578 ;
  assign n9213 = n3559 & ~n3561 ;
  assign n9214 = ~n3569 & ~n3576 ;
  assign n9215 = ~n9213 & n9214 ;
  assign n9216 = ~n9212 & ~n9215 ;
  assign n9217 = ~n3561 & ~n3578 ;
  assign n9218 = ~n3564 & n9217 ;
  assign n9219 = ~n3566 & n3571 ;
  assign n9220 = ~\s9_msel_arb0_state_reg[0]/NET0131  & ~n3566 ;
  assign n9221 = ~n9219 & ~n9220 ;
  assign n9222 = n9218 & n9221 ;
  assign n9223 = ~n9216 & ~n9222 ;
  assign n9224 = n3612 & ~n9223 ;
  assign n9225 = ~n3566 & ~n3569 ;
  assign n9226 = ~n9219 & ~n9225 ;
  assign n9227 = ~\s9_msel_arb0_state_reg[1]/NET0131  & \s9_msel_arb0_state_reg[2]/NET0131  ;
  assign n9228 = ~\rf_conf9_reg[3]/NET0131  & ~\s9_msel_arb0_state_reg[1]/NET0131  ;
  assign n9229 = n3575 & n9228 ;
  assign n9230 = ~n9227 & ~n9229 ;
  assign n9231 = n9226 & ~n9230 ;
  assign n9232 = ~n3559 & n3564 ;
  assign n9233 = ~n3561 & ~n9232 ;
  assign n9234 = ~n3576 & ~n9233 ;
  assign n9235 = ~n3571 & ~n3578 ;
  assign n9236 = \s9_msel_arb0_state_reg[2]/NET0131  & ~n9235 ;
  assign n9237 = ~n9230 & ~n9236 ;
  assign n9238 = ~n9234 & n9237 ;
  assign n9239 = ~n9231 & ~n9238 ;
  assign n9240 = ~n9224 & n9239 ;
  assign n9241 = \s9_msel_arb0_state_reg[0]/NET0131  & ~n9240 ;
  assign n9242 = \s9_msel_arb0_state_reg[0]/NET0131  & n9235 ;
  assign n9243 = ~n3561 & ~n3564 ;
  assign n9244 = n9242 & n9243 ;
  assign n9245 = n3606 & n9244 ;
  assign n9246 = n3576 & n9235 ;
  assign n9247 = ~n3559 & ~n9226 ;
  assign n9248 = ~n9246 & n9247 ;
  assign n9249 = ~\rf_conf9_reg[5]/NET0131  & ~\s9_msel_arb0_state_reg[0]/NET0131  ;
  assign n9250 = n3560 & n9249 ;
  assign n9251 = ~n9232 & ~n9250 ;
  assign n9252 = n3606 & n9251 ;
  assign n9253 = ~n9248 & n9252 ;
  assign n9254 = ~n9245 & ~n9253 ;
  assign n9255 = ~n3576 & ~n9213 ;
  assign n9256 = ~n3578 & ~n9255 ;
  assign n9257 = ~n3564 & ~n3571 ;
  assign n9258 = \s9_msel_arb0_state_reg[2]/NET0131  & ~n9257 ;
  assign n9259 = n9256 & ~n9258 ;
  assign n9260 = ~\s9_msel_arb0_state_reg[2]/NET0131  & ~n9217 ;
  assign n9261 = ~n3564 & n9226 ;
  assign n9262 = ~n9260 & n9261 ;
  assign n9263 = ~n9259 & ~n9262 ;
  assign n9264 = ~\s9_msel_arb0_state_reg[0]/NET0131  & ~\s9_msel_arb0_state_reg[1]/NET0131  ;
  assign n9265 = ~n9263 & n9264 ;
  assign n9266 = ~n9242 & n9247 ;
  assign n9267 = ~\s9_msel_arb0_state_reg[1]/NET0131  & ~\s9_msel_arb0_state_reg[2]/NET0131  ;
  assign n9268 = \s9_msel_arb0_state_reg[0]/NET0131  & n9267 ;
  assign n9269 = ~n3576 & n9268 ;
  assign n9270 = n9233 & n9269 ;
  assign n9271 = ~n9266 & n9270 ;
  assign n9272 = n9218 & ~n9220 ;
  assign n9273 = ~n9216 & ~n9272 ;
  assign n9274 = \s9_msel_arb0_state_reg[2]/NET0131  & n3595 ;
  assign n9275 = ~n3571 & n9274 ;
  assign n9276 = ~n9273 & n9275 ;
  assign n9277 = ~n9271 & ~n9276 ;
  assign n9278 = ~n9265 & n9277 ;
  assign n9279 = n9254 & n9278 ;
  assign n9280 = ~n9241 & n9279 ;
  assign n9281 = ~n5406 & ~n5413 ;
  assign n9282 = n5408 & ~n5413 ;
  assign n9283 = ~n9281 & ~n9282 ;
  assign n9284 = ~\rf_conf9_reg[9]/NET0131  & ~\s9_msel_arb1_state_reg[0]/NET0131  ;
  assign n9285 = n5410 & n9284 ;
  assign n9286 = n5423 & ~n9285 ;
  assign n9287 = n9283 & n9286 ;
  assign n9288 = n5396 & ~n5401 ;
  assign n9289 = ~n5394 & ~n5401 ;
  assign n9290 = ~n9288 & ~n9289 ;
  assign n9291 = ~n5396 & ~n5411 ;
  assign n9292 = \s9_msel_arb1_state_reg[0]/NET0131  & n9291 ;
  assign n9293 = ~n9290 & ~n9292 ;
  assign n9294 = ~n5399 & ~n5408 ;
  assign n9295 = n9286 & n9294 ;
  assign n9296 = ~n9293 & n9295 ;
  assign n9297 = ~n9287 & ~n9296 ;
  assign n9298 = ~n9288 & n9294 ;
  assign n9299 = ~n9283 & ~n9298 ;
  assign n9300 = ~n5411 & ~n9299 ;
  assign n9301 = ~n5394 & ~n9300 ;
  assign n9302 = \s9_msel_arb1_state_reg[0]/NET0131  & n5429 ;
  assign n9303 = n9281 & n9289 ;
  assign n9304 = ~n5396 & n5429 ;
  assign n9305 = ~n9303 & n9304 ;
  assign n9306 = ~n9302 & ~n9305 ;
  assign n9307 = ~n9301 & ~n9306 ;
  assign n9308 = n9297 & ~n9307 ;
  assign n9309 = ~\rf_conf9_reg[1]/NET0131  & ~\s9_msel_arb1_state_reg[0]/NET0131  ;
  assign n9310 = n5398 & n9309 ;
  assign n9311 = n9290 & ~n9310 ;
  assign n9312 = n9291 & ~n9310 ;
  assign n9313 = n9283 & n9312 ;
  assign n9314 = ~n9311 & ~n9313 ;
  assign n9315 = n9292 & n9294 ;
  assign n9316 = n9314 & ~n9315 ;
  assign n9317 = n5416 & ~n9316 ;
  assign n9318 = n5413 & n9291 ;
  assign n9319 = ~n9290 & ~n9318 ;
  assign n9320 = ~n5399 & ~n9319 ;
  assign n9321 = ~n5406 & ~n9315 ;
  assign n9322 = ~n9320 & n9321 ;
  assign n9323 = ~\rf_conf9_reg[13]/NET0131  & ~\s9_msel_arb1_state_reg[0]/NET0131  ;
  assign n9324 = n5407 & n9323 ;
  assign n9325 = \s9_msel_arb1_state_reg[1]/NET0131  & \s9_msel_arb1_state_reg[2]/NET0131  ;
  assign n9326 = ~n9324 & n9325 ;
  assign n9327 = ~n9322 & n9326 ;
  assign n9328 = ~n9317 & ~n9327 ;
  assign n9329 = n9308 & n9328 ;
  assign n9330 = \rf_conf9_reg[5]/NET0131  & n3560 ;
  assign n9331 = \rf_conf9_reg[7]/NET0131  & n3558 ;
  assign n9332 = ~n9330 & n9331 ;
  assign n9333 = \s9_msel_arb2_state_reg[1]/NET0131  & ~\s9_msel_arb2_state_reg[2]/NET0131  ;
  assign n9334 = n9332 & n9333 ;
  assign n9335 = \rf_conf9_reg[11]/NET0131  & n3565 ;
  assign n9336 = \rf_conf9_reg[15]/NET0131  & n3568 ;
  assign n9337 = \rf_conf9_reg[13]/NET0131  & n3570 ;
  assign n9338 = n9336 & ~n9337 ;
  assign n9339 = ~n9335 & ~n9338 ;
  assign n9340 = \rf_conf9_reg[3]/NET0131  & n3575 ;
  assign n9341 = \rf_conf9_reg[1]/NET0131  & n3577 ;
  assign n9342 = ~n9337 & ~n9341 ;
  assign n9343 = n9340 & n9342 ;
  assign n9344 = n9339 & ~n9343 ;
  assign n9345 = \rf_conf9_reg[9]/NET0131  & n3563 ;
  assign n9346 = ~n9330 & ~n9345 ;
  assign n9347 = n9333 & n9346 ;
  assign n9348 = ~n9344 & n9347 ;
  assign n9349 = ~n9334 & ~n9348 ;
  assign n9350 = ~n9332 & ~n9340 ;
  assign n9351 = ~\s9_msel_arb2_state_reg[1]/NET0131  & ~\s9_msel_arb2_state_reg[2]/NET0131  ;
  assign n9352 = ~n9341 & n9351 ;
  assign n9353 = ~n9350 & n9352 ;
  assign n9354 = n9346 & n9352 ;
  assign n9355 = ~n9339 & n9354 ;
  assign n9356 = ~n9353 & ~n9355 ;
  assign n9357 = ~\s9_msel_arb2_state_reg[0]/NET0131  & n9356 ;
  assign n9358 = n9349 & n9357 ;
  assign n9359 = \s9_msel_arb2_state_reg[1]/NET0131  & \s9_msel_arb2_state_reg[2]/NET0131  ;
  assign n9360 = n9338 & n9359 ;
  assign n9361 = n9335 & n9346 ;
  assign n9362 = n9350 & ~n9361 ;
  assign n9363 = n9342 & n9359 ;
  assign n9364 = ~n9362 & n9363 ;
  assign n9365 = ~n9360 & ~n9364 ;
  assign n9366 = ~\s9_msel_arb2_state_reg[1]/NET0131  & \s9_msel_arb2_state_reg[2]/NET0131  ;
  assign n9367 = ~n9345 & n9366 ;
  assign n9368 = n9335 & n9367 ;
  assign n9369 = ~n9336 & n9341 ;
  assign n9370 = ~n9336 & ~n9340 ;
  assign n9371 = ~n9332 & n9370 ;
  assign n9372 = ~n9369 & ~n9371 ;
  assign n9373 = ~n9337 & n9367 ;
  assign n9374 = n9372 & n9373 ;
  assign n9375 = ~n9368 & ~n9374 ;
  assign n9376 = n9365 & n9375 ;
  assign n9377 = n9358 & n9376 ;
  assign n9378 = \s9_msel_arb2_state_reg[0]/NET0131  & ~n9341 ;
  assign n9379 = n9346 & n9378 ;
  assign n9380 = ~n9372 & ~n9379 ;
  assign n9381 = \s9_msel_arb2_state_reg[0]/NET0131  & n9366 ;
  assign n9382 = ~n9335 & n9381 ;
  assign n9383 = ~n9337 & n9382 ;
  assign n9384 = ~n9380 & n9383 ;
  assign n9385 = n9377 & ~n9384 ;
  assign n9386 = ~n9339 & n9346 ;
  assign n9387 = n9350 & ~n9386 ;
  assign n9388 = \s9_msel_arb2_state_reg[0]/NET0131  & n9346 ;
  assign n9389 = n9342 & n9388 ;
  assign n9390 = n9387 & ~n9389 ;
  assign n9391 = n9351 & ~n9390 ;
  assign n9392 = n9331 & n9333 ;
  assign n9393 = n9330 & ~n9340 ;
  assign n9394 = n9342 & ~n9393 ;
  assign n9395 = n9339 & ~n9394 ;
  assign n9396 = n9333 & ~n9345 ;
  assign n9397 = ~n9395 & n9396 ;
  assign n9398 = ~n9392 & ~n9397 ;
  assign n9399 = n9335 & n9366 ;
  assign n9400 = \s9_msel_arb2_state_reg[0]/NET0131  & ~n9399 ;
  assign n9401 = n9398 & n9400 ;
  assign n9402 = ~n9391 & n9401 ;
  assign n9403 = \s9_msel_arb2_state_reg[0]/NET0131  & ~n9337 ;
  assign n9404 = n9346 & n9403 ;
  assign n9405 = ~n9336 & ~n9404 ;
  assign n9406 = n9362 & n9405 ;
  assign n9407 = ~n9369 & ~n9406 ;
  assign n9408 = n9359 & n9407 ;
  assign n9409 = ~n9384 & ~n9408 ;
  assign n9410 = n9402 & n9409 ;
  assign n9411 = ~n9385 & ~n9410 ;
  assign n9412 = \rf_conf9_reg[9]/NET0131  & n5410 ;
  assign n9413 = \rf_conf9_reg[15]/NET0131  & n5405 ;
  assign n9414 = \rf_conf9_reg[1]/NET0131  & n5398 ;
  assign n9415 = ~n9413 & n9414 ;
  assign n9416 = \rf_conf9_reg[7]/NET0131  & n5393 ;
  assign n9417 = \rf_conf9_reg[5]/NET0131  & n5395 ;
  assign n9418 = n9416 & ~n9417 ;
  assign n9419 = \rf_conf9_reg[3]/NET0131  & n5400 ;
  assign n9420 = ~n9413 & ~n9419 ;
  assign n9421 = ~n9418 & n9420 ;
  assign n9422 = ~n9415 & ~n9421 ;
  assign n9423 = \rf_conf9_reg[11]/NET0131  & n5412 ;
  assign n9424 = ~n9422 & ~n9423 ;
  assign n9425 = \rf_conf9_reg[13]/NET0131  & n5407 ;
  assign n9426 = ~n9423 & n9425 ;
  assign n9427 = \s9_msel_arb3_state_reg[0]/NET0131  & ~n9426 ;
  assign n9428 = ~n9424 & n9427 ;
  assign n9429 = n9412 & ~n9428 ;
  assign n9430 = ~n9414 & ~n9425 ;
  assign n9431 = \s9_msel_arb3_state_reg[0]/NET0131  & ~n9417 ;
  assign n9432 = n9430 & n9431 ;
  assign n9433 = n9426 & ~n9432 ;
  assign n9434 = ~n9423 & ~n9432 ;
  assign n9435 = ~n9422 & n9434 ;
  assign n9436 = ~n9433 & ~n9435 ;
  assign n9437 = ~\s9_msel_arb3_state_reg[1]/NET0131  & \s9_msel_arb3_state_reg[2]/NET0131  ;
  assign n9438 = n9436 & n9437 ;
  assign n9439 = ~n9429 & n9438 ;
  assign n9440 = \s9_msel_arb3_state_reg[1]/NET0131  & \s9_msel_arb3_state_reg[2]/NET0131  ;
  assign n9441 = n9413 & ~n9425 ;
  assign n9442 = n9440 & n9441 ;
  assign n9443 = ~n9418 & ~n9419 ;
  assign n9444 = ~\s9_msel_arb3_state_reg[0]/NET0131  & ~n9423 ;
  assign n9445 = ~n9412 & ~n9417 ;
  assign n9446 = ~n9444 & n9445 ;
  assign n9447 = n9443 & ~n9446 ;
  assign n9448 = n9430 & n9440 ;
  assign n9449 = ~n9447 & n9448 ;
  assign n9450 = ~n9442 & ~n9449 ;
  assign n9451 = ~\s9_msel_arb3_state_reg[1]/NET0131  & ~\s9_msel_arb3_state_reg[2]/NET0131  ;
  assign n9452 = ~n9414 & n9419 ;
  assign n9453 = n9451 & n9452 ;
  assign n9454 = n9412 & ~n9416 ;
  assign n9455 = ~n9416 & ~n9423 ;
  assign n9456 = ~n9441 & n9455 ;
  assign n9457 = ~n9454 & ~n9456 ;
  assign n9458 = ~n9414 & ~n9417 ;
  assign n9459 = n9451 & n9458 ;
  assign n9460 = n9457 & n9459 ;
  assign n9461 = ~n9453 & ~n9460 ;
  assign n9462 = n9450 & n9461 ;
  assign n9463 = ~\s9_msel_arb3_state_reg[0]/NET0131  & ~n9462 ;
  assign n9464 = n9419 & n9451 ;
  assign n9465 = \s9_msel_arb3_state_reg[0]/NET0131  & n9464 ;
  assign n9466 = ~n9414 & ~n9426 ;
  assign n9467 = n9446 & n9466 ;
  assign n9468 = ~n9422 & ~n9467 ;
  assign n9469 = \s9_msel_arb3_state_reg[0]/NET0131  & n9440 ;
  assign n9470 = ~n9468 & n9469 ;
  assign n9471 = ~n9465 & ~n9470 ;
  assign n9472 = ~n9419 & n9451 ;
  assign n9473 = n9431 & n9472 ;
  assign n9474 = \rf_conf9_reg[5]/NET0131  & ~\s9_msel_arb3_state_reg[0]/NET0131  ;
  assign n9475 = n5395 & n9474 ;
  assign n9476 = \s9_msel_arb3_state_reg[1]/NET0131  & ~\s9_msel_arb3_state_reg[2]/NET0131  ;
  assign n9477 = ~n9475 & n9476 ;
  assign n9478 = ~n9473 & ~n9477 ;
  assign n9479 = n9457 & ~n9478 ;
  assign n9480 = n9430 & n9473 ;
  assign n9481 = ~n9412 & n9480 ;
  assign n9482 = ~n9425 & n9452 ;
  assign n9483 = ~n9432 & ~n9482 ;
  assign n9484 = ~n9412 & n9477 ;
  assign n9485 = ~n9483 & n9484 ;
  assign n9486 = ~n9481 & ~n9485 ;
  assign n9487 = ~n9479 & n9486 ;
  assign n9488 = n9471 & n9487 ;
  assign n9489 = ~n9463 & n9488 ;
  assign n9490 = ~n9439 & n9489 ;
  assign n9491 = ~n3632 & n3641 ;
  assign n9492 = n3622 & ~n3624 ;
  assign n9493 = ~n3632 & ~n3639 ;
  assign n9494 = ~n9492 & n9493 ;
  assign n9495 = ~n9491 & ~n9494 ;
  assign n9496 = ~n3624 & ~n3641 ;
  assign n9497 = ~n3627 & n9496 ;
  assign n9498 = ~n3629 & n3634 ;
  assign n9499 = ~\s0_msel_arb0_state_reg[0]/NET0131  & ~n3629 ;
  assign n9500 = ~n9498 & ~n9499 ;
  assign n9501 = n9497 & n9500 ;
  assign n9502 = ~n9495 & ~n9501 ;
  assign n9503 = n3675 & ~n9502 ;
  assign n9504 = ~n3629 & ~n3632 ;
  assign n9505 = ~n9498 & ~n9504 ;
  assign n9506 = ~\s0_msel_arb0_state_reg[1]/NET0131  & \s0_msel_arb0_state_reg[2]/NET0131  ;
  assign n9507 = ~\rf_conf0_reg[3]/NET0131  & ~\s0_msel_arb0_state_reg[1]/NET0131  ;
  assign n9508 = n3638 & n9507 ;
  assign n9509 = ~n9506 & ~n9508 ;
  assign n9510 = n9505 & ~n9509 ;
  assign n9511 = ~n3622 & n3627 ;
  assign n9512 = ~n3624 & ~n9511 ;
  assign n9513 = ~n3639 & ~n9512 ;
  assign n9514 = ~n3634 & ~n3641 ;
  assign n9515 = \s0_msel_arb0_state_reg[2]/NET0131  & ~n9514 ;
  assign n9516 = ~n9509 & ~n9515 ;
  assign n9517 = ~n9513 & n9516 ;
  assign n9518 = ~n9510 & ~n9517 ;
  assign n9519 = ~n9503 & n9518 ;
  assign n9520 = \s0_msel_arb0_state_reg[0]/NET0131  & ~n9519 ;
  assign n9521 = \s0_msel_arb0_state_reg[0]/NET0131  & n9514 ;
  assign n9522 = ~n3624 & ~n3627 ;
  assign n9523 = n9521 & n9522 ;
  assign n9524 = n3669 & n9523 ;
  assign n9525 = n3639 & n9514 ;
  assign n9526 = ~n3622 & ~n9505 ;
  assign n9527 = ~n9525 & n9526 ;
  assign n9528 = ~\rf_conf0_reg[5]/NET0131  & ~\s0_msel_arb0_state_reg[0]/NET0131  ;
  assign n9529 = n3623 & n9528 ;
  assign n9530 = ~n9511 & ~n9529 ;
  assign n9531 = n3669 & n9530 ;
  assign n9532 = ~n9527 & n9531 ;
  assign n9533 = ~n9524 & ~n9532 ;
  assign n9534 = ~n3639 & ~n9492 ;
  assign n9535 = ~n3641 & ~n9534 ;
  assign n9536 = ~n3627 & ~n3634 ;
  assign n9537 = \s0_msel_arb0_state_reg[2]/NET0131  & ~n9536 ;
  assign n9538 = n9535 & ~n9537 ;
  assign n9539 = ~\s0_msel_arb0_state_reg[2]/NET0131  & ~n9496 ;
  assign n9540 = ~n3627 & n9505 ;
  assign n9541 = ~n9539 & n9540 ;
  assign n9542 = ~n9538 & ~n9541 ;
  assign n9543 = ~\s0_msel_arb0_state_reg[0]/NET0131  & ~\s0_msel_arb0_state_reg[1]/NET0131  ;
  assign n9544 = ~n9542 & n9543 ;
  assign n9545 = ~n9521 & n9526 ;
  assign n9546 = ~\s0_msel_arb0_state_reg[1]/NET0131  & ~\s0_msel_arb0_state_reg[2]/NET0131  ;
  assign n9547 = \s0_msel_arb0_state_reg[0]/NET0131  & n9546 ;
  assign n9548 = ~n3639 & n9547 ;
  assign n9549 = n9512 & n9548 ;
  assign n9550 = ~n9545 & n9549 ;
  assign n9551 = n9497 & ~n9499 ;
  assign n9552 = ~n9495 & ~n9551 ;
  assign n9553 = \s0_msel_arb0_state_reg[2]/NET0131  & n3658 ;
  assign n9554 = ~n3634 & n9553 ;
  assign n9555 = ~n9552 & n9554 ;
  assign n9556 = ~n9550 & ~n9555 ;
  assign n9557 = ~n9544 & n9556 ;
  assign n9558 = n9533 & n9557 ;
  assign n9559 = ~n9520 & n9558 ;
  assign n9560 = ~n5452 & ~n5456 ;
  assign n9561 = n5453 & ~n5456 ;
  assign n9562 = ~n9560 & ~n9561 ;
  assign n9563 = ~\rf_conf0_reg[9]/NET0131  & ~\s0_msel_arb1_state_reg[0]/NET0131  ;
  assign n9564 = n4825 & n9563 ;
  assign n9565 = n5466 & ~n9564 ;
  assign n9566 = n9562 & n9565 ;
  assign n9567 = n5445 & ~n5448 ;
  assign n9568 = ~n5444 & ~n5448 ;
  assign n9569 = ~n9567 & ~n9568 ;
  assign n9570 = ~n5445 & ~n5455 ;
  assign n9571 = \s0_msel_arb1_state_reg[0]/NET0131  & n9570 ;
  assign n9572 = ~n9569 & ~n9571 ;
  assign n9573 = ~n5447 & ~n5453 ;
  assign n9574 = n9565 & n9573 ;
  assign n9575 = ~n9572 & n9574 ;
  assign n9576 = ~n9566 & ~n9575 ;
  assign n9577 = ~n9567 & n9573 ;
  assign n9578 = ~n9562 & ~n9577 ;
  assign n9579 = ~n5455 & ~n9578 ;
  assign n9580 = ~n5444 & ~n9579 ;
  assign n9581 = \s0_msel_arb1_state_reg[0]/NET0131  & n5472 ;
  assign n9582 = n9560 & n9568 ;
  assign n9583 = ~n5445 & n5472 ;
  assign n9584 = ~n9582 & n9583 ;
  assign n9585 = ~n9581 & ~n9584 ;
  assign n9586 = ~n9580 & ~n9585 ;
  assign n9587 = n9576 & ~n9586 ;
  assign n9588 = ~\rf_conf0_reg[1]/NET0131  & ~\s0_msel_arb1_state_reg[0]/NET0131  ;
  assign n9589 = n4847 & n9588 ;
  assign n9590 = n9569 & ~n9589 ;
  assign n9591 = n9570 & ~n9589 ;
  assign n9592 = n9562 & n9591 ;
  assign n9593 = ~n9590 & ~n9592 ;
  assign n9594 = n9571 & n9573 ;
  assign n9595 = n9593 & ~n9594 ;
  assign n9596 = n5459 & ~n9595 ;
  assign n9597 = n5456 & n9570 ;
  assign n9598 = ~n9569 & ~n9597 ;
  assign n9599 = ~n5447 & ~n9598 ;
  assign n9600 = ~n5452 & ~n9594 ;
  assign n9601 = ~n9599 & n9600 ;
  assign n9602 = ~\rf_conf0_reg[13]/NET0131  & ~\s0_msel_arb1_state_reg[0]/NET0131  ;
  assign n9603 = n4837 & n9602 ;
  assign n9604 = \s0_msel_arb1_state_reg[1]/NET0131  & \s0_msel_arb1_state_reg[2]/NET0131  ;
  assign n9605 = ~n9603 & n9604 ;
  assign n9606 = ~n9601 & n9605 ;
  assign n9607 = ~n9596 & ~n9606 ;
  assign n9608 = n9587 & n9607 ;
  assign n9609 = ~\s0_msel_arb2_state_reg[1]/NET0131  & \s0_msel_arb2_state_reg[2]/NET0131  ;
  assign n9610 = ~n4159 & n9609 ;
  assign n9611 = n4158 & n9610 ;
  assign n9612 = ~n4162 & n4179 ;
  assign n9613 = n4165 & ~n4168 ;
  assign n9614 = ~n4162 & ~n4173 ;
  assign n9615 = ~n9613 & n9614 ;
  assign n9616 = ~n9612 & ~n9615 ;
  assign n9617 = ~n4161 & n9610 ;
  assign n9618 = n9616 & n9617 ;
  assign n9619 = ~n9611 & ~n9618 ;
  assign n9620 = ~\s0_msel_arb2_state_reg[0]/NET0131  & ~n9619 ;
  assign n9621 = ~n4159 & ~n4168 ;
  assign n9622 = ~n9613 & ~n9621 ;
  assign n9623 = ~n4161 & n4162 ;
  assign n9624 = ~n4158 & ~n9623 ;
  assign n9625 = ~n4161 & ~n4179 ;
  assign n9626 = n4173 & n9625 ;
  assign n9627 = n9624 & ~n9626 ;
  assign n9628 = \s0_msel_arb2_state_reg[0]/NET0131  & n9625 ;
  assign n9629 = ~n9613 & ~n9628 ;
  assign n9630 = n9627 & n9629 ;
  assign n9631 = ~n9622 & ~n9630 ;
  assign n9632 = \s0_msel_arb2_state_reg[1]/NET0131  & ~\s0_msel_arb2_state_reg[2]/NET0131  ;
  assign n9633 = ~\s0_msel_arb2_state_reg[0]/NET0131  & n9632 ;
  assign n9634 = n9631 & n9633 ;
  assign n9635 = ~n9620 & ~n9634 ;
  assign n9636 = \s0_msel_arb2_state_reg[0]/NET0131  & ~n4161 ;
  assign n9637 = ~n4158 & ~n9636 ;
  assign n9638 = ~n4179 & n9621 ;
  assign n9639 = ~n9637 & n9638 ;
  assign n9640 = ~n9616 & ~n9639 ;
  assign n9641 = \rf_conf0_reg[13]/NET0131  & ~\s0_msel_arb2_state_reg[0]/NET0131  ;
  assign n9642 = n3633 & n9641 ;
  assign n9643 = \s0_msel_arb2_state_reg[1]/NET0131  & \s0_msel_arb2_state_reg[2]/NET0131  ;
  assign n9644 = ~n9642 & n9643 ;
  assign n9645 = ~n9640 & n9644 ;
  assign n9646 = ~n4159 & ~n9627 ;
  assign n9647 = n9621 & n9628 ;
  assign n9648 = ~n4165 & ~n9647 ;
  assign n9649 = ~n9646 & n9648 ;
  assign n9650 = \s0_msel_arb2_state_reg[0]/NET0131  & n9632 ;
  assign n9651 = ~n9649 & n9650 ;
  assign n9652 = ~n9645 & ~n9651 ;
  assign n9653 = \s0_msel_arb2_state_reg[0]/NET0131  & ~\s0_msel_arb2_state_reg[1]/NET0131  ;
  assign n9654 = \s0_msel_arb2_state_reg[2]/NET0131  & n9653 ;
  assign n9655 = ~n4161 & n9616 ;
  assign n9656 = ~n4158 & ~n9647 ;
  assign n9657 = ~n9655 & n9656 ;
  assign n9658 = n9654 & ~n9657 ;
  assign n9659 = ~n4173 & ~n9613 ;
  assign n9660 = \rf_conf0_reg[1]/NET0131  & ~\s0_msel_arb2_state_reg[0]/NET0131  ;
  assign n9661 = n3640 & n9660 ;
  assign n9662 = ~n9659 & ~n9661 ;
  assign n9663 = n9621 & ~n9661 ;
  assign n9664 = ~n9624 & n9663 ;
  assign n9665 = ~n9662 & ~n9664 ;
  assign n9666 = ~n9647 & n9665 ;
  assign n9667 = ~\s0_msel_arb2_state_reg[1]/NET0131  & ~\s0_msel_arb2_state_reg[2]/NET0131  ;
  assign n9668 = ~n9666 & n9667 ;
  assign n9669 = ~n9658 & ~n9668 ;
  assign n9670 = n9652 & n9669 ;
  assign n9671 = n9635 & n9670 ;
  assign n9672 = \s0_msel_arb3_state_reg[1]/NET0131  & ~\s0_msel_arb3_state_reg[2]/NET0131  ;
  assign n9673 = ~n4857 & n9672 ;
  assign n9674 = ~n4824 & ~n4836 ;
  assign n9675 = ~n4824 & n4838 ;
  assign n9676 = ~n9674 & ~n9675 ;
  assign n9677 = n9673 & n9676 ;
  assign n9678 = ~n4846 & ~n4864 ;
  assign n9679 = ~n4838 & ~n4848 ;
  assign n9680 = n9673 & n9679 ;
  assign n9681 = ~n9678 & n9680 ;
  assign n9682 = ~n9677 & ~n9681 ;
  assign n9683 = ~n4826 & ~n9682 ;
  assign n9684 = n4841 & ~n4843 ;
  assign n9685 = ~n4846 & ~n9684 ;
  assign n9686 = ~n4848 & ~n9685 ;
  assign n9687 = n9674 & ~n9686 ;
  assign n9688 = ~\s0_msel_arb3_state_reg[0]/NET0131  & \s0_msel_arb3_state_reg[2]/NET0131  ;
  assign n9689 = ~\s0_msel_arb3_state_reg[1]/NET0131  & n9688 ;
  assign n9690 = ~n9675 & n9689 ;
  assign n9691 = ~n4826 & n9690 ;
  assign n9692 = ~n9687 & n9691 ;
  assign n9693 = ~n9683 & ~n9692 ;
  assign n9694 = ~\s0_msel_arb3_state_reg[1]/NET0131  & ~\s0_msel_arb3_state_reg[2]/NET0131  ;
  assign n9695 = \rf_conf0_reg[1]/NET0131  & ~\s0_msel_arb3_state_reg[0]/NET0131  ;
  assign n9696 = n4847 & n9695 ;
  assign n9697 = n9694 & ~n9696 ;
  assign n9698 = ~n9685 & n9697 ;
  assign n9699 = ~n4826 & ~n4843 ;
  assign n9700 = n9697 & n9699 ;
  assign n9701 = n9676 & n9700 ;
  assign n9702 = ~n9698 & ~n9701 ;
  assign n9703 = n4841 & n9673 ;
  assign n9704 = ~\s0_msel_arb3_state_reg[1]/NET0131  & n4829 ;
  assign n9705 = n4824 & n9704 ;
  assign n9706 = ~n9703 & ~n9705 ;
  assign n9707 = n9702 & n9706 ;
  assign n9708 = n9693 & n9707 ;
  assign n9709 = \s0_msel_arb3_state_reg[0]/NET0131  & n9694 ;
  assign n9710 = ~n4848 & n9709 ;
  assign n9711 = n9699 & n9710 ;
  assign n9712 = ~n4824 & n9704 ;
  assign n9713 = ~n9711 & ~n9712 ;
  assign n9714 = ~n4836 & n4848 ;
  assign n9715 = ~n4836 & ~n4846 ;
  assign n9716 = ~n9684 & n9715 ;
  assign n9717 = ~n9714 & ~n9716 ;
  assign n9718 = \s0_msel_arb3_state_reg[0]/NET0131  & ~n4848 ;
  assign n9719 = n9699 & n9718 ;
  assign n9720 = ~n9711 & ~n9719 ;
  assign n9721 = ~n9717 & n9720 ;
  assign n9722 = ~n9713 & ~n9721 ;
  assign n9723 = ~n4838 & n9722 ;
  assign n9724 = ~n4848 & n9699 ;
  assign n9725 = ~\s0_msel_arb3_state_reg[0]/NET0131  & ~n4824 ;
  assign n9726 = n9724 & ~n9725 ;
  assign n9727 = ~n9717 & ~n9726 ;
  assign n9728 = ~\s0_msel_arb3_state_reg[0]/NET0131  & n4838 ;
  assign n9729 = n4838 & n9674 ;
  assign n9730 = n9685 & n9729 ;
  assign n9731 = ~n9728 & ~n9730 ;
  assign n9732 = n4871 & n9731 ;
  assign n9733 = ~n9727 & n9732 ;
  assign n9734 = ~n9723 & ~n9733 ;
  assign n9735 = n9708 & n9734 ;
  assign n9736 = ~n3695 & n3704 ;
  assign n9737 = n3685 & ~n3687 ;
  assign n9738 = ~n3695 & ~n3702 ;
  assign n9739 = ~n9737 & n9738 ;
  assign n9740 = ~n9736 & ~n9739 ;
  assign n9741 = ~n3687 & ~n3704 ;
  assign n9742 = ~n3690 & n9741 ;
  assign n9743 = ~n3692 & n3697 ;
  assign n9744 = ~\s10_msel_arb0_state_reg[0]/NET0131  & ~n3692 ;
  assign n9745 = ~n9743 & ~n9744 ;
  assign n9746 = n9742 & n9745 ;
  assign n9747 = ~n9740 & ~n9746 ;
  assign n9748 = n3738 & ~n9747 ;
  assign n9749 = ~n3692 & ~n3695 ;
  assign n9750 = ~n9743 & ~n9749 ;
  assign n9751 = ~\s10_msel_arb0_state_reg[1]/NET0131  & \s10_msel_arb0_state_reg[2]/NET0131  ;
  assign n9752 = ~\rf_conf10_reg[3]/NET0131  & ~\s10_msel_arb0_state_reg[1]/NET0131  ;
  assign n9753 = n3701 & n9752 ;
  assign n9754 = ~n9751 & ~n9753 ;
  assign n9755 = n9750 & ~n9754 ;
  assign n9756 = ~n3685 & n3690 ;
  assign n9757 = ~n3687 & ~n9756 ;
  assign n9758 = ~n3702 & ~n9757 ;
  assign n9759 = ~n3697 & ~n3704 ;
  assign n9760 = \s10_msel_arb0_state_reg[2]/NET0131  & ~n9759 ;
  assign n9761 = ~n9754 & ~n9760 ;
  assign n9762 = ~n9758 & n9761 ;
  assign n9763 = ~n9755 & ~n9762 ;
  assign n9764 = ~n9748 & n9763 ;
  assign n9765 = \s10_msel_arb0_state_reg[0]/NET0131  & ~n9764 ;
  assign n9766 = \s10_msel_arb0_state_reg[0]/NET0131  & n9759 ;
  assign n9767 = ~n3687 & ~n3690 ;
  assign n9768 = n9766 & n9767 ;
  assign n9769 = n3732 & n9768 ;
  assign n9770 = n3702 & n9759 ;
  assign n9771 = ~n3685 & ~n9750 ;
  assign n9772 = ~n9770 & n9771 ;
  assign n9773 = ~\rf_conf10_reg[5]/NET0131  & ~\s10_msel_arb0_state_reg[0]/NET0131  ;
  assign n9774 = n3686 & n9773 ;
  assign n9775 = ~n9756 & ~n9774 ;
  assign n9776 = n3732 & n9775 ;
  assign n9777 = ~n9772 & n9776 ;
  assign n9778 = ~n9769 & ~n9777 ;
  assign n9779 = ~n3702 & ~n9737 ;
  assign n9780 = ~n3704 & ~n9779 ;
  assign n9781 = ~n3690 & ~n3697 ;
  assign n9782 = \s10_msel_arb0_state_reg[2]/NET0131  & ~n9781 ;
  assign n9783 = n9780 & ~n9782 ;
  assign n9784 = ~\s10_msel_arb0_state_reg[2]/NET0131  & ~n9741 ;
  assign n9785 = ~n3690 & n9750 ;
  assign n9786 = ~n9784 & n9785 ;
  assign n9787 = ~n9783 & ~n9786 ;
  assign n9788 = ~\s10_msel_arb0_state_reg[0]/NET0131  & ~\s10_msel_arb0_state_reg[1]/NET0131  ;
  assign n9789 = ~n9787 & n9788 ;
  assign n9790 = ~n9766 & n9771 ;
  assign n9791 = ~\s10_msel_arb0_state_reg[1]/NET0131  & ~\s10_msel_arb0_state_reg[2]/NET0131  ;
  assign n9792 = \s10_msel_arb0_state_reg[0]/NET0131  & n9791 ;
  assign n9793 = ~n3702 & n9792 ;
  assign n9794 = n9757 & n9793 ;
  assign n9795 = ~n9790 & n9794 ;
  assign n9796 = n9742 & ~n9744 ;
  assign n9797 = ~n9740 & ~n9796 ;
  assign n9798 = \s10_msel_arb0_state_reg[2]/NET0131  & n3721 ;
  assign n9799 = ~n3697 & n9798 ;
  assign n9800 = ~n9797 & n9799 ;
  assign n9801 = ~n9795 & ~n9800 ;
  assign n9802 = ~n9789 & n9801 ;
  assign n9803 = n9778 & n9802 ;
  assign n9804 = ~n9765 & n9803 ;
  assign n9805 = ~n5570 & ~n5571 ;
  assign n9806 = ~n5560 & n5596 ;
  assign n9807 = n9805 & n9806 ;
  assign n9808 = ~n5561 & n9807 ;
  assign n9809 = ~n5560 & ~n5570 ;
  assign n9810 = ~\s10_msel_arb2_state_reg[1]/NET0131  & ~n9809 ;
  assign n9811 = ~\s10_msel_arb2_state_reg[2]/NET0131  & ~n9810 ;
  assign n9812 = ~n5566 & ~n5567 ;
  assign n9813 = ~n5565 & ~n5575 ;
  assign n9814 = n9812 & n9813 ;
  assign n9815 = ~n5561 & ~n9814 ;
  assign n9816 = n9811 & n9815 ;
  assign n9817 = ~n9808 & ~n9816 ;
  assign n9818 = ~n5565 & n9812 ;
  assign n9819 = n5596 & ~n9818 ;
  assign n9820 = n9817 & ~n9819 ;
  assign n9821 = \s10_msel_arb2_state_reg[0]/NET0131  & ~n9820 ;
  assign n9822 = \s10_msel_arb2_state_reg[0]/NET0131  & ~\s10_msel_arb2_state_reg[1]/NET0131  ;
  assign n9823 = ~n5560 & ~n5561 ;
  assign n9824 = n9805 & n9823 ;
  assign n9825 = \s10_msel_arb2_state_reg[0]/NET0131  & ~n5566 ;
  assign n9826 = ~n9824 & n9825 ;
  assign n9827 = ~n9822 & ~n9826 ;
  assign n9828 = ~\s10_msel_arb2_state_reg[1]/NET0131  & ~n9813 ;
  assign n9829 = n9812 & ~n9828 ;
  assign n9830 = ~n9824 & n9829 ;
  assign n9831 = n9827 & ~n9830 ;
  assign n9832 = \s10_msel_arb2_state_reg[2]/NET0131  & ~n9831 ;
  assign n9833 = ~\s10_msel_arb2_state_reg[0]/NET0131  & ~n9814 ;
  assign n9834 = ~\s10_msel_arb2_state_reg[1]/NET0131  & ~n9805 ;
  assign n9835 = n9823 & ~n9834 ;
  assign n9836 = n9833 & n9835 ;
  assign n9837 = ~\s10_msel_arb2_state_reg[2]/NET0131  & ~n9836 ;
  assign n9838 = ~n9832 & ~n9837 ;
  assign n9839 = ~n9821 & ~n9838 ;
  assign n9840 = ~n6105 & ~n6106 ;
  assign n9841 = ~n6095 & n6131 ;
  assign n9842 = n9840 & n9841 ;
  assign n9843 = ~n6096 & n9842 ;
  assign n9844 = ~n6095 & ~n6105 ;
  assign n9845 = ~\s12_msel_arb2_state_reg[1]/NET0131  & ~n9844 ;
  assign n9846 = ~\s12_msel_arb2_state_reg[2]/NET0131  & ~n9845 ;
  assign n9847 = ~n6101 & ~n6102 ;
  assign n9848 = ~n6100 & ~n6110 ;
  assign n9849 = n9847 & n9848 ;
  assign n9850 = ~n6096 & ~n9849 ;
  assign n9851 = n9846 & n9850 ;
  assign n9852 = ~n9843 & ~n9851 ;
  assign n9853 = ~n6100 & n9847 ;
  assign n9854 = n6131 & ~n9853 ;
  assign n9855 = n9852 & ~n9854 ;
  assign n9856 = \s12_msel_arb2_state_reg[0]/NET0131  & ~n9855 ;
  assign n9857 = \s12_msel_arb2_state_reg[0]/NET0131  & ~\s12_msel_arb2_state_reg[1]/NET0131  ;
  assign n9858 = ~n6095 & ~n6096 ;
  assign n9859 = n9840 & n9858 ;
  assign n9860 = \s12_msel_arb2_state_reg[0]/NET0131  & ~n6101 ;
  assign n9861 = ~n9859 & n9860 ;
  assign n9862 = ~n9857 & ~n9861 ;
  assign n9863 = ~\s12_msel_arb2_state_reg[1]/NET0131  & ~n9848 ;
  assign n9864 = n9847 & ~n9863 ;
  assign n9865 = ~n9859 & n9864 ;
  assign n9866 = n9862 & ~n9865 ;
  assign n9867 = \s12_msel_arb2_state_reg[2]/NET0131  & ~n9866 ;
  assign n9868 = ~\s12_msel_arb2_state_reg[0]/NET0131  & ~n9849 ;
  assign n9869 = ~\s12_msel_arb2_state_reg[1]/NET0131  & ~n9840 ;
  assign n9870 = n9858 & ~n9869 ;
  assign n9871 = n9868 & n9870 ;
  assign n9872 = ~\s12_msel_arb2_state_reg[2]/NET0131  & ~n9871 ;
  assign n9873 = ~n9867 & ~n9872 ;
  assign n9874 = ~n9856 & ~n9873 ;
  assign n9875 = ~n6394 & ~n6399 ;
  assign n9876 = ~n6396 & ~n6397 ;
  assign n9877 = n9875 & n9876 ;
  assign n9878 = ~n6393 & ~n9877 ;
  assign n9879 = \rf_conf13_reg[9]/NET0131  & ~\s13_msel_arb2_state_reg[1]/NET0131  ;
  assign n9880 = n2866 & n9879 ;
  assign n9881 = ~n6405 & ~n9880 ;
  assign n9882 = ~\s13_msel_arb2_state_reg[0]/NET0131  & ~n9881 ;
  assign n9883 = ~n6403 & ~n6405 ;
  assign n9884 = ~\s13_msel_arb2_state_reg[1]/NET0131  & ~n9883 ;
  assign n9885 = ~n9882 & ~n9884 ;
  assign n9886 = n9878 & n9885 ;
  assign n9887 = \s13_msel_arb2_state_reg[2]/NET0131  & ~n9886 ;
  assign n9888 = ~\s13_msel_arb2_state_reg[2]/NET0131  & ~n6396 ;
  assign n9889 = ~n6397 & ~n6399 ;
  assign n9890 = ~\s13_msel_arb2_state_reg[1]/NET0131  & ~n9889 ;
  assign n9891 = n9888 & ~n9890 ;
  assign n9892 = ~n6393 & ~n6405 ;
  assign n9893 = ~n6392 & ~n6403 ;
  assign n9894 = n9892 & n9893 ;
  assign n9895 = ~\s13_msel_arb2_state_reg[0]/NET0131  & n6397 ;
  assign n9896 = ~\s13_msel_arb2_state_reg[0]/NET0131  & ~\s13_msel_arb2_state_reg[1]/NET0131  ;
  assign n9897 = n6394 & n9896 ;
  assign n9898 = ~n9895 & ~n9897 ;
  assign n9899 = ~n9894 & n9898 ;
  assign n9900 = n9891 & n9899 ;
  assign n9901 = ~n9887 & ~n9900 ;
  assign n9902 = ~n7439 & ~n7444 ;
  assign n9903 = ~n7441 & ~n7442 ;
  assign n9904 = n9902 & n9903 ;
  assign n9905 = ~n7438 & ~n9904 ;
  assign n9906 = \rf_conf2_reg[9]/NET0131  & ~\s2_msel_arb2_state_reg[1]/NET0131  ;
  assign n9907 = n3437 & n9906 ;
  assign n9908 = ~n7450 & ~n9907 ;
  assign n9909 = ~\s2_msel_arb2_state_reg[0]/NET0131  & ~n9908 ;
  assign n9910 = ~n7448 & ~n7450 ;
  assign n9911 = ~\s2_msel_arb2_state_reg[1]/NET0131  & ~n9910 ;
  assign n9912 = ~n9909 & ~n9911 ;
  assign n9913 = n9905 & n9912 ;
  assign n9914 = \s2_msel_arb2_state_reg[2]/NET0131  & ~n9913 ;
  assign n9915 = ~\s2_msel_arb2_state_reg[2]/NET0131  & ~n7441 ;
  assign n9916 = ~n7442 & ~n7444 ;
  assign n9917 = ~\s2_msel_arb2_state_reg[1]/NET0131  & ~n9916 ;
  assign n9918 = n9915 & ~n9917 ;
  assign n9919 = ~n7438 & ~n7450 ;
  assign n9920 = ~n7437 & ~n7448 ;
  assign n9921 = n9919 & n9920 ;
  assign n9922 = ~\s2_msel_arb2_state_reg[0]/NET0131  & n7442 ;
  assign n9923 = ~\s2_msel_arb2_state_reg[0]/NET0131  & ~\s2_msel_arb2_state_reg[1]/NET0131  ;
  assign n9924 = n7439 & n9923 ;
  assign n9925 = ~n9922 & ~n9924 ;
  assign n9926 = ~n9921 & n9925 ;
  assign n9927 = n9918 & n9926 ;
  assign n9928 = ~n9914 & ~n9927 ;
  assign n9929 = ~n8008 & ~n8013 ;
  assign n9930 = ~n8010 & ~n8011 ;
  assign n9931 = n9929 & n9930 ;
  assign n9932 = ~n8007 & ~n9931 ;
  assign n9933 = \rf_conf4_reg[9]/NET0131  & ~\s4_msel_arb2_state_reg[1]/NET0131  ;
  assign n9934 = n3123 & n9933 ;
  assign n9935 = ~n8019 & ~n9934 ;
  assign n9936 = ~\s4_msel_arb2_state_reg[0]/NET0131  & ~n9935 ;
  assign n9937 = ~n8017 & ~n8019 ;
  assign n9938 = ~\s4_msel_arb2_state_reg[1]/NET0131  & ~n9937 ;
  assign n9939 = ~n9936 & ~n9938 ;
  assign n9940 = n9932 & n9939 ;
  assign n9941 = \s4_msel_arb2_state_reg[2]/NET0131  & ~n9940 ;
  assign n9942 = ~\s4_msel_arb2_state_reg[2]/NET0131  & ~n8010 ;
  assign n9943 = ~n8011 & ~n8013 ;
  assign n9944 = ~\s4_msel_arb2_state_reg[1]/NET0131  & ~n9943 ;
  assign n9945 = n9942 & ~n9944 ;
  assign n9946 = ~n8007 & ~n8019 ;
  assign n9947 = ~n8006 & ~n8017 ;
  assign n9948 = n9946 & n9947 ;
  assign n9949 = ~\s4_msel_arb2_state_reg[0]/NET0131  & n8011 ;
  assign n9950 = ~\s4_msel_arb2_state_reg[0]/NET0131  & ~\s4_msel_arb2_state_reg[1]/NET0131  ;
  assign n9951 = n8008 & n9950 ;
  assign n9952 = ~n9949 & ~n9951 ;
  assign n9953 = ~n9948 & n9952 ;
  assign n9954 = n9945 & n9953 ;
  assign n9955 = ~n9941 & ~n9954 ;
  assign n9956 = ~n8815 & ~n8816 ;
  assign n9957 = ~n8805 & n8841 ;
  assign n9958 = n9956 & n9957 ;
  assign n9959 = ~n8806 & n9958 ;
  assign n9960 = ~n8805 & ~n8815 ;
  assign n9961 = ~\s7_msel_arb2_state_reg[1]/NET0131  & ~n9960 ;
  assign n9962 = ~\s7_msel_arb2_state_reg[2]/NET0131  & ~n9961 ;
  assign n9963 = ~n8811 & ~n8812 ;
  assign n9964 = ~n8810 & ~n8820 ;
  assign n9965 = n9963 & n9964 ;
  assign n9966 = ~n8806 & ~n9965 ;
  assign n9967 = n9962 & n9966 ;
  assign n9968 = ~n9959 & ~n9967 ;
  assign n9969 = ~n8810 & n9963 ;
  assign n9970 = n8841 & ~n9969 ;
  assign n9971 = n9968 & ~n9970 ;
  assign n9972 = \s7_msel_arb2_state_reg[0]/NET0131  & ~n9971 ;
  assign n9973 = \s7_msel_arb2_state_reg[0]/NET0131  & ~\s7_msel_arb2_state_reg[1]/NET0131  ;
  assign n9974 = ~n8805 & ~n8806 ;
  assign n9975 = n9956 & n9974 ;
  assign n9976 = \s7_msel_arb2_state_reg[0]/NET0131  & ~n8811 ;
  assign n9977 = ~n9975 & n9976 ;
  assign n9978 = ~n9973 & ~n9977 ;
  assign n9979 = ~\s7_msel_arb2_state_reg[1]/NET0131  & ~n9964 ;
  assign n9980 = n9963 & ~n9979 ;
  assign n9981 = ~n9975 & n9980 ;
  assign n9982 = n9978 & ~n9981 ;
  assign n9983 = \s7_msel_arb2_state_reg[2]/NET0131  & ~n9982 ;
  assign n9984 = ~\s7_msel_arb2_state_reg[0]/NET0131  & ~n9965 ;
  assign n9985 = ~\s7_msel_arb2_state_reg[1]/NET0131  & ~n9956 ;
  assign n9986 = n9974 & ~n9985 ;
  assign n9987 = n9984 & n9986 ;
  assign n9988 = ~\s7_msel_arb2_state_reg[2]/NET0131  & ~n9987 ;
  assign n9989 = ~n9983 & ~n9988 ;
  assign n9990 = ~n9972 & ~n9989 ;
  assign n9991 = ~n9340 & ~n9341 ;
  assign n9992 = ~n9330 & n9366 ;
  assign n9993 = n9991 & n9992 ;
  assign n9994 = ~n9331 & n9993 ;
  assign n9995 = ~n9330 & ~n9340 ;
  assign n9996 = ~\s9_msel_arb2_state_reg[1]/NET0131  & ~n9995 ;
  assign n9997 = ~\s9_msel_arb2_state_reg[2]/NET0131  & ~n9996 ;
  assign n9998 = ~n9336 & ~n9337 ;
  assign n9999 = ~n9335 & ~n9345 ;
  assign n10000 = n9998 & n9999 ;
  assign n10001 = ~n9331 & ~n10000 ;
  assign n10002 = n9997 & n10001 ;
  assign n10003 = ~n9994 & ~n10002 ;
  assign n10004 = ~n9335 & n9998 ;
  assign n10005 = n9366 & ~n10004 ;
  assign n10006 = n10003 & ~n10005 ;
  assign n10007 = \s9_msel_arb2_state_reg[0]/NET0131  & ~n10006 ;
  assign n10008 = \s9_msel_arb2_state_reg[0]/NET0131  & ~\s9_msel_arb2_state_reg[1]/NET0131  ;
  assign n10009 = ~n9330 & ~n9331 ;
  assign n10010 = n9991 & n10009 ;
  assign n10011 = \s9_msel_arb2_state_reg[0]/NET0131  & ~n9336 ;
  assign n10012 = ~n10010 & n10011 ;
  assign n10013 = ~n10008 & ~n10012 ;
  assign n10014 = ~\s9_msel_arb2_state_reg[1]/NET0131  & ~n9999 ;
  assign n10015 = n9998 & ~n10014 ;
  assign n10016 = ~n10010 & n10015 ;
  assign n10017 = n10013 & ~n10016 ;
  assign n10018 = \s9_msel_arb2_state_reg[2]/NET0131  & ~n10017 ;
  assign n10019 = ~\s9_msel_arb2_state_reg[0]/NET0131  & ~n10000 ;
  assign n10020 = ~\s9_msel_arb2_state_reg[1]/NET0131  & ~n9991 ;
  assign n10021 = n10009 & ~n10020 ;
  assign n10022 = n10019 & n10021 ;
  assign n10023 = ~\s9_msel_arb2_state_reg[2]/NET0131  & ~n10022 ;
  assign n10024 = ~n10018 & ~n10023 ;
  assign n10025 = ~n10007 & ~n10024 ;
  assign n10026 = ~n9414 & ~n9419 ;
  assign n10027 = ~n9416 & ~n9417 ;
  assign n10028 = n10026 & n10027 ;
  assign n10029 = ~n9413 & ~n10028 ;
  assign n10030 = \rf_conf9_reg[9]/NET0131  & ~\s9_msel_arb3_state_reg[1]/NET0131  ;
  assign n10031 = n5410 & n10030 ;
  assign n10032 = ~n9425 & ~n10031 ;
  assign n10033 = ~\s9_msel_arb3_state_reg[0]/NET0131  & ~n10032 ;
  assign n10034 = ~n9423 & ~n9425 ;
  assign n10035 = ~\s9_msel_arb3_state_reg[1]/NET0131  & ~n10034 ;
  assign n10036 = ~n10033 & ~n10035 ;
  assign n10037 = n10029 & n10036 ;
  assign n10038 = \s9_msel_arb3_state_reg[2]/NET0131  & ~n10037 ;
  assign n10039 = ~\s9_msel_arb3_state_reg[2]/NET0131  & ~n9416 ;
  assign n10040 = ~n9417 & ~n9419 ;
  assign n10041 = ~\s9_msel_arb3_state_reg[1]/NET0131  & ~n10040 ;
  assign n10042 = n10039 & ~n10041 ;
  assign n10043 = ~n9413 & ~n9425 ;
  assign n10044 = ~n9412 & ~n9423 ;
  assign n10045 = n10043 & n10044 ;
  assign n10046 = ~\s9_msel_arb3_state_reg[0]/NET0131  & n9417 ;
  assign n10047 = ~\s9_msel_arb3_state_reg[0]/NET0131  & ~\s9_msel_arb3_state_reg[1]/NET0131  ;
  assign n10048 = n9414 & n10047 ;
  assign n10049 = ~n10046 & ~n10048 ;
  assign n10050 = ~n10045 & n10049 ;
  assign n10051 = n10042 & n10050 ;
  assign n10052 = ~n10038 & ~n10051 ;
  assign n10053 = ~\s10_msel_arb0_state_reg[1]/NET0131  & ~n3727 ;
  assign n10054 = n3688 & n3705 ;
  assign n10055 = \s10_msel_arb0_state_reg[0]/NET0131  & \s10_msel_arb0_state_reg[1]/NET0131  ;
  assign n10056 = n3697 & ~n10055 ;
  assign n10057 = ~n3695 & ~n10056 ;
  assign n10058 = ~n10054 & n10057 ;
  assign n10059 = ~n10053 & n10058 ;
  assign n10060 = \s10_msel_arb0_state_reg[2]/NET0131  & ~n10059 ;
  assign n10061 = ~\s10_msel_arb0_state_reg[1]/NET0131  & n3702 ;
  assign n10062 = n3704 & n9788 ;
  assign n10063 = ~n10061 & ~n10062 ;
  assign n10064 = ~n3687 & n10063 ;
  assign n10065 = ~n10055 & ~n10064 ;
  assign n10066 = n9749 & n9781 ;
  assign n10067 = ~\s10_msel_arb0_state_reg[2]/NET0131  & ~n3685 ;
  assign n10068 = ~n10066 & n10067 ;
  assign n10069 = ~n10065 & n10068 ;
  assign n10070 = ~n10060 & ~n10069 ;
  assign n10071 = ~\s11_msel_arb0_state_reg[0]/NET0131  & n5741 ;
  assign n10072 = ~n2743 & ~n2748 ;
  assign n10073 = n5734 & n10072 ;
  assign n10074 = ~n2758 & n5741 ;
  assign n10075 = ~n10073 & n10074 ;
  assign n10076 = ~n10071 & ~n10075 ;
  assign n10077 = ~\rf_conf11_reg[9]/NET0131  & ~\s11_msel_arb0_state_reg[2]/NET0131  ;
  assign n10078 = n2742 & n10077 ;
  assign n10079 = ~n2748 & ~n10078 ;
  assign n10080 = n5734 & n10079 ;
  assign n10081 = ~n2751 & n2765 ;
  assign n10082 = ~n10080 & n10081 ;
  assign n10083 = ~\s11_msel_arb0_state_reg[1]/NET0131  & n10082 ;
  assign n10084 = ~n2748 & n5734 ;
  assign n10085 = n2754 & n2765 ;
  assign n10086 = n10084 & ~n10085 ;
  assign n10087 = n2791 & ~n10086 ;
  assign n10088 = ~n10083 & ~n10087 ;
  assign n10089 = n10076 & n10088 ;
  assign n10090 = n2765 & n5741 ;
  assign n10091 = ~n10073 & n10090 ;
  assign n10092 = ~\s11_msel_arb0_state_reg[0]/NET0131  & ~n10091 ;
  assign n10093 = ~n10089 & ~n10092 ;
  assign n10094 = ~\rf_conf11_reg[13]/NET0131  & \s11_msel_arb0_state_reg[1]/NET0131  ;
  assign n10095 = n2747 & n10094 ;
  assign n10096 = ~n10085 & ~n10095 ;
  assign n10097 = \s11_msel_arb0_state_reg[2]/NET0131  & ~n10096 ;
  assign n10098 = ~\s11_msel_arb0_state_reg[2]/NET0131  & ~n10085 ;
  assign n10099 = ~\s11_msel_arb0_state_reg[1]/NET0131  & ~n10073 ;
  assign n10100 = ~n10098 & n10099 ;
  assign n10101 = ~n10097 & ~n10100 ;
  assign n10102 = ~\s11_msel_arb0_state_reg[0]/NET0131  & ~n10101 ;
  assign n10103 = ~n2746 & ~n10085 ;
  assign n10104 = n5720 & ~n10103 ;
  assign n10105 = ~n10102 & ~n10104 ;
  assign n10106 = ~n10093 & n10105 ;
  assign n10107 = ~\s12_msel_arb0_state_reg[0]/NET0131  & n6004 ;
  assign n10108 = n5997 & n6023 ;
  assign n10109 = ~n2820 & n6004 ;
  assign n10110 = ~n10108 & n10109 ;
  assign n10111 = ~n10107 & ~n10110 ;
  assign n10112 = ~\rf_conf12_reg[9]/NET0131  & ~\s12_msel_arb0_state_reg[2]/NET0131  ;
  assign n10113 = n2804 & n10112 ;
  assign n10114 = ~n2810 & ~n10113 ;
  assign n10115 = n5997 & n10114 ;
  assign n10116 = ~n2813 & n2827 ;
  assign n10117 = ~n10115 & n10116 ;
  assign n10118 = ~\s12_msel_arb0_state_reg[1]/NET0131  & n10117 ;
  assign n10119 = ~n2810 & n5997 ;
  assign n10120 = n2816 & n2827 ;
  assign n10121 = n10119 & ~n10120 ;
  assign n10122 = n2853 & ~n10121 ;
  assign n10123 = ~n10118 & ~n10122 ;
  assign n10124 = n10111 & n10123 ;
  assign n10125 = n2827 & n6004 ;
  assign n10126 = ~n10108 & n10125 ;
  assign n10127 = ~\s12_msel_arb0_state_reg[0]/NET0131  & ~n10126 ;
  assign n10128 = ~n10124 & ~n10127 ;
  assign n10129 = ~\rf_conf12_reg[13]/NET0131  & \s12_msel_arb0_state_reg[1]/NET0131  ;
  assign n10130 = n2809 & n10129 ;
  assign n10131 = ~n10120 & ~n10130 ;
  assign n10132 = \s12_msel_arb0_state_reg[2]/NET0131  & ~n10131 ;
  assign n10133 = ~\s12_msel_arb0_state_reg[2]/NET0131  & ~n10120 ;
  assign n10134 = ~\s12_msel_arb0_state_reg[1]/NET0131  & ~n10108 ;
  assign n10135 = ~n10133 & n10134 ;
  assign n10136 = ~n10132 & ~n10135 ;
  assign n10137 = ~\s12_msel_arb0_state_reg[0]/NET0131  & ~n10136 ;
  assign n10138 = ~n2808 & ~n10120 ;
  assign n10139 = n5983 & ~n10138 ;
  assign n10140 = ~n10137 & ~n10139 ;
  assign n10141 = ~n10128 & n10140 ;
  assign n10142 = ~\s13_msel_arb0_state_reg[0]/NET0131  & n6276 ;
  assign n10143 = n6269 & n6295 ;
  assign n10144 = ~n2882 & n6276 ;
  assign n10145 = ~n10143 & n10144 ;
  assign n10146 = ~n10142 & ~n10145 ;
  assign n10147 = ~\rf_conf13_reg[9]/NET0131  & ~\s13_msel_arb0_state_reg[2]/NET0131  ;
  assign n10148 = n2866 & n10147 ;
  assign n10149 = ~n2872 & ~n10148 ;
  assign n10150 = n6269 & n10149 ;
  assign n10151 = ~n2875 & n2889 ;
  assign n10152 = ~n10150 & n10151 ;
  assign n10153 = ~\s13_msel_arb0_state_reg[1]/NET0131  & n10152 ;
  assign n10154 = ~n2872 & n6269 ;
  assign n10155 = n2878 & n2889 ;
  assign n10156 = n10154 & ~n10155 ;
  assign n10157 = n2915 & ~n10156 ;
  assign n10158 = ~n10153 & ~n10157 ;
  assign n10159 = n10146 & n10158 ;
  assign n10160 = n2889 & n6276 ;
  assign n10161 = ~n10143 & n10160 ;
  assign n10162 = ~\s13_msel_arb0_state_reg[0]/NET0131  & ~n10161 ;
  assign n10163 = ~n10159 & ~n10162 ;
  assign n10164 = ~\rf_conf13_reg[13]/NET0131  & \s13_msel_arb0_state_reg[1]/NET0131  ;
  assign n10165 = n2871 & n10164 ;
  assign n10166 = ~n10155 & ~n10165 ;
  assign n10167 = \s13_msel_arb0_state_reg[2]/NET0131  & ~n10166 ;
  assign n10168 = ~\s13_msel_arb0_state_reg[2]/NET0131  & ~n10155 ;
  assign n10169 = ~\s13_msel_arb0_state_reg[1]/NET0131  & ~n10143 ;
  assign n10170 = ~n10168 & n10169 ;
  assign n10171 = ~n10167 & ~n10170 ;
  assign n10172 = ~\s13_msel_arb0_state_reg[0]/NET0131  & ~n10171 ;
  assign n10173 = ~n2870 & ~n10155 ;
  assign n10174 = n6255 & ~n10173 ;
  assign n10175 = ~n10172 & ~n10174 ;
  assign n10176 = ~n10163 & n10175 ;
  assign n10177 = ~\s14_msel_arb0_state_reg[0]/NET0131  & n6570 ;
  assign n10178 = n6563 & n6589 ;
  assign n10179 = ~n2944 & n6570 ;
  assign n10180 = ~n10178 & n10179 ;
  assign n10181 = ~n10177 & ~n10180 ;
  assign n10182 = ~\rf_conf14_reg[9]/NET0131  & ~\s14_msel_arb0_state_reg[2]/NET0131  ;
  assign n10183 = n2928 & n10182 ;
  assign n10184 = ~n2934 & ~n10183 ;
  assign n10185 = n6563 & n10184 ;
  assign n10186 = ~n2937 & n2951 ;
  assign n10187 = ~n10185 & n10186 ;
  assign n10188 = ~\s14_msel_arb0_state_reg[1]/NET0131  & n10187 ;
  assign n10189 = ~n2934 & n6563 ;
  assign n10190 = n2940 & n2951 ;
  assign n10191 = n10189 & ~n10190 ;
  assign n10192 = n2977 & ~n10191 ;
  assign n10193 = ~n10188 & ~n10192 ;
  assign n10194 = n10181 & n10193 ;
  assign n10195 = n2951 & n6570 ;
  assign n10196 = ~n10178 & n10195 ;
  assign n10197 = ~\s14_msel_arb0_state_reg[0]/NET0131  & ~n10196 ;
  assign n10198 = ~n10194 & ~n10197 ;
  assign n10199 = ~\rf_conf14_reg[13]/NET0131  & \s14_msel_arb0_state_reg[1]/NET0131  ;
  assign n10200 = n2933 & n10199 ;
  assign n10201 = ~n10190 & ~n10200 ;
  assign n10202 = \s14_msel_arb0_state_reg[2]/NET0131  & ~n10201 ;
  assign n10203 = ~\s14_msel_arb0_state_reg[2]/NET0131  & ~n10190 ;
  assign n10204 = ~\s14_msel_arb0_state_reg[1]/NET0131  & ~n10178 ;
  assign n10205 = ~n10203 & n10204 ;
  assign n10206 = ~n10202 & ~n10205 ;
  assign n10207 = ~\s14_msel_arb0_state_reg[0]/NET0131  & ~n10206 ;
  assign n10208 = ~n2932 & ~n10190 ;
  assign n10209 = n6549 & ~n10208 ;
  assign n10210 = ~n10207 & ~n10209 ;
  assign n10211 = ~n10198 & n10210 ;
  assign n10212 = n3008 & ~n3010 ;
  assign n10213 = ~n2996 & ~n10212 ;
  assign n10214 = ~n3004 & ~n3010 ;
  assign n10215 = n3002 & n10214 ;
  assign n10216 = n10213 & ~n10215 ;
  assign n10217 = \s15_msel_arb0_state_reg[0]/NET0131  & ~n2991 ;
  assign n10218 = n10214 & n10217 ;
  assign n10219 = n10216 & ~n10218 ;
  assign n10220 = ~n2994 & n3048 ;
  assign n10221 = ~n10219 & n10220 ;
  assign n10222 = n2989 & ~n2991 ;
  assign n10223 = ~n3002 & ~n10222 ;
  assign n10224 = ~n2991 & ~n2994 ;
  assign n10225 = n2996 & n10224 ;
  assign n10226 = n10223 & ~n10225 ;
  assign n10227 = \s15_msel_arb0_state_reg[0]/NET0131  & ~n3010 ;
  assign n10228 = n10224 & n10227 ;
  assign n10229 = n10226 & ~n10228 ;
  assign n10230 = ~n3004 & n3042 ;
  assign n10231 = ~n10229 & n10230 ;
  assign n10232 = ~\s15_msel_arb0_state_reg[2]/NET0131  & n3040 ;
  assign n10233 = n3008 & n10232 ;
  assign n10234 = n2989 & n3047 ;
  assign n10235 = ~n10233 & ~n10234 ;
  assign n10236 = n3053 & n10235 ;
  assign n10237 = ~n10231 & n10236 ;
  assign n10238 = ~n10221 & n10237 ;
  assign n10239 = ~n2989 & n2994 ;
  assign n10240 = ~n2989 & ~n2996 ;
  assign n10241 = ~n10212 & n10240 ;
  assign n10242 = ~n10239 & ~n10241 ;
  assign n10243 = \s15_msel_arb0_state_reg[0]/NET0131  & ~n2994 ;
  assign n10244 = n10214 & n10243 ;
  assign n10245 = ~n10242 & ~n10244 ;
  assign n10246 = ~n2991 & n3018 ;
  assign n10247 = ~n10245 & n10246 ;
  assign n10248 = n3004 & ~n3008 ;
  assign n10249 = ~n3002 & ~n3008 ;
  assign n10250 = ~n10222 & n10249 ;
  assign n10251 = ~n10248 & ~n10250 ;
  assign n10252 = \s15_msel_arb0_state_reg[0]/NET0131  & ~n3004 ;
  assign n10253 = n10224 & n10252 ;
  assign n10254 = ~n10251 & ~n10253 ;
  assign n10255 = ~n2996 & ~n3010 ;
  assign n10256 = n3051 & n10255 ;
  assign n10257 = ~n10254 & n10256 ;
  assign n10258 = ~n10247 & ~n10257 ;
  assign n10259 = n10238 & n10258 ;
  assign n10260 = n3002 & ~n3004 ;
  assign n10261 = ~n2991 & ~n3004 ;
  assign n10262 = n10242 & n10261 ;
  assign n10263 = ~n10260 & ~n10262 ;
  assign n10264 = ~\s15_msel_arb0_state_reg[2]/NET0131  & n3035 ;
  assign n10265 = ~n10263 & n10264 ;
  assign n10266 = ~n2994 & n2996 ;
  assign n10267 = ~n2994 & ~n3010 ;
  assign n10268 = n10251 & n10267 ;
  assign n10269 = ~n10266 & ~n10268 ;
  assign n10270 = \s15_msel_arb0_state_reg[2]/NET0131  & n3035 ;
  assign n10271 = ~n10269 & n10270 ;
  assign n10272 = ~n10265 & ~n10271 ;
  assign n10273 = ~\rf_conf15_reg[1]/NET0131  & ~\s15_msel_arb0_state_reg[0]/NET0131  ;
  assign n10274 = n3009 & n10273 ;
  assign n10275 = ~n3011 & ~n10274 ;
  assign n10276 = ~n10214 & ~n10275 ;
  assign n10277 = \s15_msel_arb0_state_reg[0]/NET0131  & n10224 ;
  assign n10278 = ~n10275 & ~n10277 ;
  assign n10279 = n10226 & n10278 ;
  assign n10280 = ~n10276 & ~n10279 ;
  assign n10281 = n3043 & n10280 ;
  assign n10282 = ~\rf_conf15_reg[9]/NET0131  & \s15_msel_arb0_state_reg[0]/NET0131  ;
  assign n10283 = n2990 & n10282 ;
  assign n10284 = ~n10222 & ~n10283 ;
  assign n10285 = ~n10224 & n10284 ;
  assign n10286 = \s15_msel_arb0_state_reg[0]/NET0131  & n10214 ;
  assign n10287 = n10284 & ~n10286 ;
  assign n10288 = n10216 & n10287 ;
  assign n10289 = ~n10285 & ~n10288 ;
  assign n10290 = n2999 & n10289 ;
  assign n10291 = ~n10281 & ~n10290 ;
  assign n10292 = n10272 & n10291 ;
  assign n10293 = n10259 & n10292 ;
  assign n10294 = n2992 & n2997 ;
  assign n10295 = ~\s15_msel_arb0_state_reg[2]/NET0131  & ~n3008 ;
  assign n10296 = n3005 & n10295 ;
  assign n10297 = ~n10274 & n10296 ;
  assign n10298 = ~n10294 & n10297 ;
  assign n10299 = n3005 & n3011 ;
  assign n10300 = n10294 & ~n10299 ;
  assign n10301 = ~\s15_msel_arb0_state_reg[0]/NET0131  & \s15_msel_arb0_state_reg[2]/NET0131  ;
  assign n10302 = ~n10300 & n10301 ;
  assign n10303 = ~n10298 & ~n10302 ;
  assign n10304 = ~\s15_msel_arb0_state_reg[1]/NET0131  & ~n10303 ;
  assign n10305 = ~n3004 & n3047 ;
  assign n10306 = n3011 & n10305 ;
  assign n10307 = ~n3002 & n10306 ;
  assign n10308 = ~\rf_conf15_reg[5]/NET0131  & ~\s15_msel_arb0_state_reg[0]/NET0131  ;
  assign n10309 = n3003 & n10308 ;
  assign n10310 = \s15_msel_arb0_state_reg[1]/NET0131  & ~\s15_msel_arb0_state_reg[2]/NET0131  ;
  assign n10311 = ~n10309 & n10310 ;
  assign n10312 = ~n3002 & n10311 ;
  assign n10313 = ~n10294 & n10312 ;
  assign n10314 = ~n10307 & ~n10313 ;
  assign n10315 = ~n2989 & n2997 ;
  assign n10316 = n3047 & ~n10315 ;
  assign n10317 = ~\rf_conf15_reg[13]/NET0131  & ~\s15_msel_arb0_state_reg[0]/NET0131  ;
  assign n10318 = n2993 & n10317 ;
  assign n10319 = ~n2996 & ~n10318 ;
  assign n10320 = ~n10299 & n10319 ;
  assign n10321 = \s15_msel_arb0_state_reg[1]/NET0131  & \s15_msel_arb0_state_reg[2]/NET0131  ;
  assign n10322 = ~n10320 & n10321 ;
  assign n10323 = ~n10316 & ~n10322 ;
  assign n10324 = n10314 & n10323 ;
  assign n10325 = ~n10304 & n10324 ;
  assign n10326 = n3772 & ~n3779 ;
  assign n10327 = n3775 & ~n10326 ;
  assign n10328 = \s15_msel_arb2_state_reg[2]/NET0131  & n6943 ;
  assign n10329 = ~n10327 & n10328 ;
  assign n10330 = n6950 & ~n6954 ;
  assign n10331 = \s15_msel_arb2_state_reg[1]/NET0131  & ~n10330 ;
  assign n10332 = ~n3775 & n3782 ;
  assign n10333 = \s15_msel_arb2_state_reg[1]/NET0131  & n3779 ;
  assign n10334 = ~n10332 & n10333 ;
  assign n10335 = ~n10331 & ~n10334 ;
  assign n10336 = ~n10329 & ~n10335 ;
  assign n10337 = ~n3772 & n3775 ;
  assign n10338 = n3782 & ~n10337 ;
  assign n10339 = ~\s15_msel_arb2_state_reg[1]/NET0131  & ~n6921 ;
  assign n10340 = n6903 & n10339 ;
  assign n10341 = ~n10338 & n10340 ;
  assign n10342 = n3779 & ~n3782 ;
  assign n10343 = n3772 & ~n10342 ;
  assign n10344 = ~\s15_msel_arb2_state_reg[1]/NET0131  & ~n6930 ;
  assign n10345 = n6902 & n10344 ;
  assign n10346 = ~n10343 & n10345 ;
  assign n10347 = ~n10341 & ~n10346 ;
  assign n10348 = ~n10336 & n10347 ;
  assign n10349 = ~n3800 & ~n3813 ;
  assign n10350 = ~n3788 & n10349 ;
  assign n10351 = n3792 & ~n6997 ;
  assign n10352 = \s15_msel_arb3_state_reg[1]/NET0131  & ~n3791 ;
  assign n10353 = ~n3813 & ~n10352 ;
  assign n10354 = ~n10351 & ~n10353 ;
  assign n10355 = ~n3788 & n3797 ;
  assign n10356 = ~n10354 & n10355 ;
  assign n10357 = ~n10350 & ~n10356 ;
  assign n10358 = ~n3793 & ~n3811 ;
  assign n10359 = ~\s15_msel_arb3_state_reg[2]/NET0131  & ~n10358 ;
  assign n10360 = n10357 & n10359 ;
  assign n10361 = ~\s15_msel_arb3_state_reg[1]/NET0131  & ~n3796 ;
  assign n10362 = n3799 & ~n7002 ;
  assign n10363 = ~n10361 & ~n10362 ;
  assign n10364 = n3790 & ~n10363 ;
  assign n10365 = ~n3795 & n10364 ;
  assign n10366 = n3790 & n3798 ;
  assign n10367 = n3793 & ~n10366 ;
  assign n10368 = n3823 & ~n10367 ;
  assign n10369 = ~n10365 & ~n10368 ;
  assign n10370 = \s15_msel_arb3_state_reg[2]/NET0131  & n3821 ;
  assign n10371 = n10369 & n10370 ;
  assign n10372 = ~n10360 & ~n10371 ;
  assign n10373 = ~\s1_msel_arb0_state_reg[1]/NET0131  & ~n3412 ;
  assign n10374 = n3373 & n3390 ;
  assign n10375 = \s1_msel_arb0_state_reg[0]/NET0131  & \s1_msel_arb0_state_reg[1]/NET0131  ;
  assign n10376 = n3382 & ~n10375 ;
  assign n10377 = ~n3380 & ~n10376 ;
  assign n10378 = ~n10374 & n10377 ;
  assign n10379 = ~n10373 & n10378 ;
  assign n10380 = \s1_msel_arb0_state_reg[2]/NET0131  & ~n10379 ;
  assign n10381 = ~\s1_msel_arb0_state_reg[1]/NET0131  & n3387 ;
  assign n10382 = n3389 & n7078 ;
  assign n10383 = ~n10381 & ~n10382 ;
  assign n10384 = ~n3372 & n10383 ;
  assign n10385 = ~n10375 & ~n10384 ;
  assign n10386 = n7039 & n7071 ;
  assign n10387 = ~\s1_msel_arb0_state_reg[2]/NET0131  & ~n3370 ;
  assign n10388 = ~n10386 & n10387 ;
  assign n10389 = ~n10385 & n10388 ;
  assign n10390 = ~n10380 & ~n10389 ;
  assign n10391 = ~\s2_msel_arb0_state_reg[1]/NET0131  & ~n3475 ;
  assign n10392 = n3436 & n3453 ;
  assign n10393 = \s2_msel_arb0_state_reg[0]/NET0131  & \s2_msel_arb0_state_reg[1]/NET0131  ;
  assign n10394 = n3445 & ~n10393 ;
  assign n10395 = ~n3443 & ~n10394 ;
  assign n10396 = ~n10392 & n10395 ;
  assign n10397 = ~n10391 & n10396 ;
  assign n10398 = \s2_msel_arb0_state_reg[2]/NET0131  & ~n10397 ;
  assign n10399 = ~\s2_msel_arb0_state_reg[1]/NET0131  & n3450 ;
  assign n10400 = n3452 & n7347 ;
  assign n10401 = ~n10399 & ~n10400 ;
  assign n10402 = ~n3435 & n10401 ;
  assign n10403 = ~n10393 & ~n10402 ;
  assign n10404 = n7308 & n7340 ;
  assign n10405 = ~\s2_msel_arb0_state_reg[2]/NET0131  & ~n3433 ;
  assign n10406 = ~n10404 & n10405 ;
  assign n10407 = ~n10403 & n10406 ;
  assign n10408 = ~n10398 & ~n10407 ;
  assign n10409 = ~\s3_msel_arb0_state_reg[0]/NET0131  & n7615 ;
  assign n10410 = n7608 & n7634 ;
  assign n10411 = ~n3077 & n7615 ;
  assign n10412 = ~n10410 & n10411 ;
  assign n10413 = ~n10409 & ~n10412 ;
  assign n10414 = ~\rf_conf3_reg[9]/NET0131  & ~\s3_msel_arb0_state_reg[2]/NET0131  ;
  assign n10415 = n3061 & n10414 ;
  assign n10416 = ~n3067 & ~n10415 ;
  assign n10417 = n7608 & n10416 ;
  assign n10418 = ~n3070 & n3084 ;
  assign n10419 = ~n10417 & n10418 ;
  assign n10420 = ~\s3_msel_arb0_state_reg[1]/NET0131  & n10419 ;
  assign n10421 = ~n3067 & n7608 ;
  assign n10422 = n3073 & n3084 ;
  assign n10423 = n10421 & ~n10422 ;
  assign n10424 = n3110 & ~n10423 ;
  assign n10425 = ~n10420 & ~n10424 ;
  assign n10426 = n10413 & n10425 ;
  assign n10427 = n3084 & n7615 ;
  assign n10428 = ~n10410 & n10427 ;
  assign n10429 = ~\s3_msel_arb0_state_reg[0]/NET0131  & ~n10428 ;
  assign n10430 = ~n10426 & ~n10429 ;
  assign n10431 = ~\rf_conf3_reg[13]/NET0131  & \s3_msel_arb0_state_reg[1]/NET0131  ;
  assign n10432 = n3066 & n10431 ;
  assign n10433 = ~n10422 & ~n10432 ;
  assign n10434 = \s3_msel_arb0_state_reg[2]/NET0131  & ~n10433 ;
  assign n10435 = ~\s3_msel_arb0_state_reg[2]/NET0131  & ~n10422 ;
  assign n10436 = ~\s3_msel_arb0_state_reg[1]/NET0131  & ~n10410 ;
  assign n10437 = ~n10435 & n10436 ;
  assign n10438 = ~n10434 & ~n10437 ;
  assign n10439 = ~\s3_msel_arb0_state_reg[0]/NET0131  & ~n10438 ;
  assign n10440 = ~n3065 & ~n10422 ;
  assign n10441 = n7594 & ~n10440 ;
  assign n10442 = ~n10439 & ~n10441 ;
  assign n10443 = ~n10430 & n10442 ;
  assign n10444 = ~\s4_msel_arb0_state_reg[0]/NET0131  & n7897 ;
  assign n10445 = n7890 & n7916 ;
  assign n10446 = ~n3139 & n7897 ;
  assign n10447 = ~n10445 & n10446 ;
  assign n10448 = ~n10444 & ~n10447 ;
  assign n10449 = ~\rf_conf4_reg[9]/NET0131  & ~\s4_msel_arb0_state_reg[2]/NET0131  ;
  assign n10450 = n3123 & n10449 ;
  assign n10451 = ~n3129 & ~n10450 ;
  assign n10452 = n7890 & n10451 ;
  assign n10453 = ~n3132 & n3146 ;
  assign n10454 = ~n10452 & n10453 ;
  assign n10455 = ~\s4_msel_arb0_state_reg[1]/NET0131  & n10454 ;
  assign n10456 = ~n3129 & n7890 ;
  assign n10457 = n3135 & n3146 ;
  assign n10458 = n10456 & ~n10457 ;
  assign n10459 = n3172 & ~n10458 ;
  assign n10460 = ~n10455 & ~n10459 ;
  assign n10461 = n10448 & n10460 ;
  assign n10462 = n3146 & n7897 ;
  assign n10463 = ~n10445 & n10462 ;
  assign n10464 = ~\s4_msel_arb0_state_reg[0]/NET0131  & ~n10463 ;
  assign n10465 = ~n10461 & ~n10464 ;
  assign n10466 = ~\rf_conf4_reg[13]/NET0131  & \s4_msel_arb0_state_reg[1]/NET0131  ;
  assign n10467 = n3128 & n10466 ;
  assign n10468 = ~n10457 & ~n10467 ;
  assign n10469 = \s4_msel_arb0_state_reg[2]/NET0131  & ~n10468 ;
  assign n10470 = ~\s4_msel_arb0_state_reg[2]/NET0131  & ~n10457 ;
  assign n10471 = ~\s4_msel_arb0_state_reg[1]/NET0131  & ~n10445 ;
  assign n10472 = ~n10470 & n10471 ;
  assign n10473 = ~n10469 & ~n10472 ;
  assign n10474 = ~\s4_msel_arb0_state_reg[0]/NET0131  & ~n10473 ;
  assign n10475 = ~n3127 & ~n10457 ;
  assign n10476 = n7876 & ~n10475 ;
  assign n10477 = ~n10474 & ~n10476 ;
  assign n10478 = ~n10465 & n10477 ;
  assign n10479 = ~\s5_msel_arb0_state_reg[0]/NET0131  & n8191 ;
  assign n10480 = n8184 & n8210 ;
  assign n10481 = ~n3201 & n8191 ;
  assign n10482 = ~n10480 & n10481 ;
  assign n10483 = ~n10479 & ~n10482 ;
  assign n10484 = ~\rf_conf5_reg[9]/NET0131  & ~\s5_msel_arb0_state_reg[2]/NET0131  ;
  assign n10485 = n3185 & n10484 ;
  assign n10486 = ~n3191 & ~n10485 ;
  assign n10487 = n8184 & n10486 ;
  assign n10488 = ~n3194 & n3208 ;
  assign n10489 = ~n10487 & n10488 ;
  assign n10490 = ~\s5_msel_arb0_state_reg[1]/NET0131  & n10489 ;
  assign n10491 = ~n3191 & n8184 ;
  assign n10492 = n3197 & n3208 ;
  assign n10493 = n10491 & ~n10492 ;
  assign n10494 = n3234 & ~n10493 ;
  assign n10495 = ~n10490 & ~n10494 ;
  assign n10496 = n10483 & n10495 ;
  assign n10497 = n3208 & n8191 ;
  assign n10498 = ~n10480 & n10497 ;
  assign n10499 = ~\s5_msel_arb0_state_reg[0]/NET0131  & ~n10498 ;
  assign n10500 = ~n10496 & ~n10499 ;
  assign n10501 = ~\rf_conf5_reg[13]/NET0131  & \s5_msel_arb0_state_reg[1]/NET0131  ;
  assign n10502 = n3190 & n10501 ;
  assign n10503 = ~n10492 & ~n10502 ;
  assign n10504 = \s5_msel_arb0_state_reg[2]/NET0131  & ~n10503 ;
  assign n10505 = ~\s5_msel_arb0_state_reg[2]/NET0131  & ~n10492 ;
  assign n10506 = ~\s5_msel_arb0_state_reg[1]/NET0131  & ~n10480 ;
  assign n10507 = ~n10505 & n10506 ;
  assign n10508 = ~n10504 & ~n10507 ;
  assign n10509 = ~\s5_msel_arb0_state_reg[0]/NET0131  & ~n10508 ;
  assign n10510 = ~n3189 & ~n10492 ;
  assign n10511 = n8170 & ~n10510 ;
  assign n10512 = ~n10509 & ~n10511 ;
  assign n10513 = ~n10500 & n10512 ;
  assign n10514 = ~\s6_msel_arb0_state_reg[0]/NET0131  & n8446 ;
  assign n10515 = n8439 & n8465 ;
  assign n10516 = ~n3263 & n8446 ;
  assign n10517 = ~n10515 & n10516 ;
  assign n10518 = ~n10514 & ~n10517 ;
  assign n10519 = ~\rf_conf6_reg[9]/NET0131  & ~\s6_msel_arb0_state_reg[2]/NET0131  ;
  assign n10520 = n3247 & n10519 ;
  assign n10521 = ~n3253 & ~n10520 ;
  assign n10522 = n8439 & n10521 ;
  assign n10523 = ~n3256 & n3270 ;
  assign n10524 = ~n10522 & n10523 ;
  assign n10525 = ~\s6_msel_arb0_state_reg[1]/NET0131  & n10524 ;
  assign n10526 = ~n3253 & n8439 ;
  assign n10527 = n3259 & n3270 ;
  assign n10528 = n10526 & ~n10527 ;
  assign n10529 = n3296 & ~n10528 ;
  assign n10530 = ~n10525 & ~n10529 ;
  assign n10531 = n10518 & n10530 ;
  assign n10532 = n3270 & n8446 ;
  assign n10533 = ~n10515 & n10532 ;
  assign n10534 = ~\s6_msel_arb0_state_reg[0]/NET0131  & ~n10533 ;
  assign n10535 = ~n10531 & ~n10534 ;
  assign n10536 = ~\rf_conf6_reg[13]/NET0131  & \s6_msel_arb0_state_reg[1]/NET0131  ;
  assign n10537 = n3252 & n10536 ;
  assign n10538 = ~n10527 & ~n10537 ;
  assign n10539 = \s6_msel_arb0_state_reg[2]/NET0131  & ~n10538 ;
  assign n10540 = ~\s6_msel_arb0_state_reg[2]/NET0131  & ~n10527 ;
  assign n10541 = ~\s6_msel_arb0_state_reg[1]/NET0131  & ~n10515 ;
  assign n10542 = ~n10540 & n10541 ;
  assign n10543 = ~n10539 & ~n10542 ;
  assign n10544 = ~\s6_msel_arb0_state_reg[0]/NET0131  & ~n10543 ;
  assign n10545 = ~n3251 & ~n10527 ;
  assign n10546 = n8425 & ~n10545 ;
  assign n10547 = ~n10544 & ~n10546 ;
  assign n10548 = ~n10535 & n10547 ;
  assign n10549 = ~\s7_msel_arb0_state_reg[1]/NET0131  & ~n3538 ;
  assign n10550 = n3499 & n3516 ;
  assign n10551 = \s7_msel_arb0_state_reg[0]/NET0131  & \s7_msel_arb0_state_reg[1]/NET0131  ;
  assign n10552 = n3508 & ~n10551 ;
  assign n10553 = ~n3506 & ~n10552 ;
  assign n10554 = ~n10550 & n10553 ;
  assign n10555 = ~n10549 & n10554 ;
  assign n10556 = \s7_msel_arb0_state_reg[2]/NET0131  & ~n10555 ;
  assign n10557 = ~\s7_msel_arb0_state_reg[1]/NET0131  & n3513 ;
  assign n10558 = n3515 & n8717 ;
  assign n10559 = ~n10557 & ~n10558 ;
  assign n10560 = ~n3498 & n10559 ;
  assign n10561 = ~n10551 & ~n10560 ;
  assign n10562 = n8678 & n8710 ;
  assign n10563 = ~\s7_msel_arb0_state_reg[2]/NET0131  & ~n3496 ;
  assign n10564 = ~n10562 & n10563 ;
  assign n10565 = ~n10561 & n10564 ;
  assign n10566 = ~n10556 & ~n10565 ;
  assign n10567 = ~\s8_msel_arb0_state_reg[0]/NET0131  & n8986 ;
  assign n10568 = n8979 & n9005 ;
  assign n10569 = ~n3325 & n8986 ;
  assign n10570 = ~n10568 & n10569 ;
  assign n10571 = ~n10567 & ~n10570 ;
  assign n10572 = ~\rf_conf8_reg[9]/NET0131  & ~\s8_msel_arb0_state_reg[2]/NET0131  ;
  assign n10573 = n3309 & n10572 ;
  assign n10574 = ~n3315 & ~n10573 ;
  assign n10575 = n8979 & n10574 ;
  assign n10576 = ~n3318 & n3332 ;
  assign n10577 = ~n10575 & n10576 ;
  assign n10578 = ~\s8_msel_arb0_state_reg[1]/NET0131  & n10577 ;
  assign n10579 = ~n3315 & n8979 ;
  assign n10580 = n3321 & n3332 ;
  assign n10581 = n10579 & ~n10580 ;
  assign n10582 = ~\s8_msel_arb0_state_reg[1]/NET0131  & \s8_msel_arb0_state_reg[2]/NET0131  ;
  assign n10583 = ~n10581 & n10582 ;
  assign n10584 = ~n10578 & ~n10583 ;
  assign n10585 = n10571 & n10584 ;
  assign n10586 = n3332 & n8986 ;
  assign n10587 = ~n10568 & n10586 ;
  assign n10588 = ~\s8_msel_arb0_state_reg[0]/NET0131  & ~n10587 ;
  assign n10589 = ~n10585 & ~n10588 ;
  assign n10590 = ~\rf_conf8_reg[13]/NET0131  & \s8_msel_arb0_state_reg[1]/NET0131  ;
  assign n10591 = n3314 & n10590 ;
  assign n10592 = ~n10580 & ~n10591 ;
  assign n10593 = \s8_msel_arb0_state_reg[2]/NET0131  & ~n10592 ;
  assign n10594 = ~\s8_msel_arb0_state_reg[2]/NET0131  & ~n10580 ;
  assign n10595 = ~\s8_msel_arb0_state_reg[1]/NET0131  & ~n10568 ;
  assign n10596 = ~n10594 & n10595 ;
  assign n10597 = ~n10593 & ~n10596 ;
  assign n10598 = ~\s8_msel_arb0_state_reg[0]/NET0131  & ~n10597 ;
  assign n10599 = ~n3313 & ~n10580 ;
  assign n10600 = n8965 & ~n10599 ;
  assign n10601 = ~n10598 & ~n10600 ;
  assign n10602 = ~n10589 & n10601 ;
  assign n10603 = ~\s9_msel_arb0_state_reg[1]/NET0131  & ~n3601 ;
  assign n10604 = n3562 & n3579 ;
  assign n10605 = \s9_msel_arb0_state_reg[0]/NET0131  & \s9_msel_arb0_state_reg[1]/NET0131  ;
  assign n10606 = n3571 & ~n10605 ;
  assign n10607 = ~n3569 & ~n10606 ;
  assign n10608 = ~n10604 & n10607 ;
  assign n10609 = ~n10603 & n10608 ;
  assign n10610 = \s9_msel_arb0_state_reg[2]/NET0131  & ~n10609 ;
  assign n10611 = ~\s9_msel_arb0_state_reg[1]/NET0131  & n3576 ;
  assign n10612 = n3578 & n9264 ;
  assign n10613 = ~n10611 & ~n10612 ;
  assign n10614 = ~n3561 & n10613 ;
  assign n10615 = ~n10605 & ~n10614 ;
  assign n10616 = n9225 & n9257 ;
  assign n10617 = ~\s9_msel_arb0_state_reg[2]/NET0131  & ~n3559 ;
  assign n10618 = ~n10616 & n10617 ;
  assign n10619 = ~n10615 & n10618 ;
  assign n10620 = ~n10610 & ~n10619 ;
  assign n10621 = ~\s0_msel_arb0_state_reg[1]/NET0131  & ~n3664 ;
  assign n10622 = n3625 & n3642 ;
  assign n10623 = \s0_msel_arb0_state_reg[0]/NET0131  & \s0_msel_arb0_state_reg[1]/NET0131  ;
  assign n10624 = n3634 & ~n10623 ;
  assign n10625 = ~n3632 & ~n10624 ;
  assign n10626 = ~n10622 & n10625 ;
  assign n10627 = ~n10621 & n10626 ;
  assign n10628 = \s0_msel_arb0_state_reg[2]/NET0131  & ~n10627 ;
  assign n10629 = ~\s0_msel_arb0_state_reg[1]/NET0131  & n3639 ;
  assign n10630 = n3641 & n9543 ;
  assign n10631 = ~n10629 & ~n10630 ;
  assign n10632 = ~n3624 & n10631 ;
  assign n10633 = ~n10623 & ~n10632 ;
  assign n10634 = n9504 & n9536 ;
  assign n10635 = ~\s0_msel_arb0_state_reg[2]/NET0131  & ~n3622 ;
  assign n10636 = ~n10634 & n10635 ;
  assign n10637 = ~n10633 & n10636 ;
  assign n10638 = ~n10628 & ~n10637 ;
  assign n10639 = ~\s10_msel_arb2_state_reg[2]/NET0131  & ~n9823 ;
  assign n10640 = ~n9805 & n9812 ;
  assign n10641 = ~\s10_msel_arb2_state_reg[0]/NET0131  & n10640 ;
  assign n10642 = ~n9828 & ~n10641 ;
  assign n10643 = ~n10639 & ~n10642 ;
  assign n10644 = ~\s10_msel_arb2_state_reg[1]/NET0131  & n9812 ;
  assign n10645 = n9823 & n10644 ;
  assign n10646 = ~n10643 & ~n10645 ;
  assign n10647 = \s10_msel_arb2_state_reg[2]/NET0131  & ~n9812 ;
  assign n10648 = ~n9813 & n9823 ;
  assign n10649 = ~\s10_msel_arb2_state_reg[0]/NET0131  & n10648 ;
  assign n10650 = ~n9834 & ~n10649 ;
  assign n10651 = ~n10647 & ~n10650 ;
  assign n10652 = n5566 & n5589 ;
  assign n10653 = n5589 & n9805 ;
  assign n10654 = ~n10648 & n10653 ;
  assign n10655 = ~n10652 & ~n10654 ;
  assign n10656 = \s10_msel_arb2_state_reg[0]/NET0131  & n10655 ;
  assign n10657 = ~n10651 & ~n10656 ;
  assign n10658 = n10646 & n10657 ;
  assign n10659 = n5612 & ~n9812 ;
  assign n10660 = \s10_msel_arb2_state_reg[1]/NET0131  & ~n5575 ;
  assign n10661 = n9823 & ~n10660 ;
  assign n10662 = n5612 & n9805 ;
  assign n10663 = ~n10661 & n10662 ;
  assign n10664 = ~n10659 & ~n10663 ;
  assign n10665 = \s10_msel_arb2_state_reg[1]/NET0131  & n5561 ;
  assign n10666 = \s10_msel_arb2_state_reg[1]/NET0131  & n9813 ;
  assign n10667 = ~n10640 & n10666 ;
  assign n10668 = ~n10665 & ~n10667 ;
  assign n10669 = ~n9812 & n9813 ;
  assign n10670 = n9823 & ~n10669 ;
  assign n10671 = ~\s10_msel_arb2_state_reg[1]/NET0131  & ~n5570 ;
  assign n10672 = ~n10670 & n10671 ;
  assign n10673 = n10668 & ~n10672 ;
  assign n10674 = \s10_msel_arb2_state_reg[0]/NET0131  & ~\s10_msel_arb2_state_reg[2]/NET0131  ;
  assign n10675 = ~n10673 & n10674 ;
  assign n10676 = n10664 & ~n10675 ;
  assign n10677 = ~n10658 & n10676 ;
  assign n10678 = ~n4216 & ~n5666 ;
  assign n10679 = ~\s10_msel_arb3_state_reg[2]/NET0131  & ~n10678 ;
  assign n10680 = ~n4199 & ~n10679 ;
  assign n10681 = n4197 & ~n4209 ;
  assign n10682 = n10680 & n10681 ;
  assign n10683 = \s10_msel_arb3_state_reg[2]/NET0131  & ~n4198 ;
  assign n10684 = ~n4214 & n10678 ;
  assign n10685 = ~n10683 & n10684 ;
  assign n10686 = ~n4194 & n4199 ;
  assign n10687 = ~n4214 & n4219 ;
  assign n10688 = n4209 & ~n10687 ;
  assign n10689 = n10686 & ~n10688 ;
  assign n10690 = ~n10685 & ~n10689 ;
  assign n10691 = ~n10682 & n10690 ;
  assign n10692 = ~\s10_msel_arb3_state_reg[1]/NET0131  & ~n10691 ;
  assign n10693 = \rf_conf10_reg[13]/NET0131  & ~\s10_msel_arb3_state_reg[0]/NET0131  ;
  assign n10694 = n4207 & n10693 ;
  assign n10695 = \s10_msel_arb3_state_reg[2]/NET0131  & ~n4219 ;
  assign n10696 = ~n4197 & n4214 ;
  assign n10697 = ~n10695 & ~n10696 ;
  assign n10698 = ~n10694 & ~n10697 ;
  assign n10699 = ~n4219 & ~n4227 ;
  assign n10700 = \s10_msel_arb3_state_reg[0]/NET0131  & n5664 ;
  assign n10701 = ~n4213 & n10700 ;
  assign n10702 = ~n10699 & ~n10701 ;
  assign n10703 = ~n4208 & ~n4211 ;
  assign n10704 = ~n10702 & n10703 ;
  assign n10705 = ~n10698 & ~n10704 ;
  assign n10706 = ~n4206 & ~n10705 ;
  assign n10707 = ~n4197 & ~n4211 ;
  assign n10708 = n4228 & n10707 ;
  assign n10709 = \s10_msel_arb3_state_reg[1]/NET0131  & ~n10708 ;
  assign n10710 = ~n10706 & n10709 ;
  assign n10711 = ~n10692 & ~n10710 ;
  assign n10712 = \rf_conf11_reg[5]/NET0131  & ~\s11_msel_arb2_state_reg[0]/NET0131  ;
  assign n10713 = n2763 & n10712 ;
  assign n10714 = n4249 & ~n10713 ;
  assign n10715 = \rf_conf11_reg[7]/NET0131  & \s11_msel_arb2_state_reg[0]/NET0131  ;
  assign n10716 = n2757 & n10715 ;
  assign n10717 = ~\s11_msel_arb2_state_reg[2]/NET0131  & ~n10716 ;
  assign n10718 = ~n10714 & n10717 ;
  assign n10719 = ~\s11_msel_arb2_state_reg[1]/NET0131  & ~n4257 ;
  assign n10720 = n4269 & ~n10719 ;
  assign n10721 = n4252 & n10717 ;
  assign n10722 = ~n10720 & n10721 ;
  assign n10723 = ~n10718 & ~n10722 ;
  assign n10724 = \s11_msel_arb2_state_reg[2]/NET0131  & ~n5868 ;
  assign n10725 = ~n4251 & n10724 ;
  assign n10726 = \s11_msel_arb2_state_reg[1]/NET0131  & ~n10725 ;
  assign n10727 = ~n4249 & n4267 ;
  assign n10728 = \s11_msel_arb2_state_reg[1]/NET0131  & n4269 ;
  assign n10729 = ~n10727 & n10728 ;
  assign n10730 = ~n10726 & ~n10729 ;
  assign n10731 = n10723 & ~n10730 ;
  assign n10732 = ~n4267 & n4269 ;
  assign n10733 = n4252 & ~n10732 ;
  assign n10734 = ~n4247 & n5880 ;
  assign n10735 = ~\s11_msel_arb2_state_reg[2]/NET0131  & ~n4269 ;
  assign n10736 = ~\s11_msel_arb2_state_reg[0]/NET0131  & ~\s11_msel_arb2_state_reg[1]/NET0131  ;
  assign n10737 = n4249 & n10736 ;
  assign n10738 = ~n10735 & n10737 ;
  assign n10739 = ~n10734 & ~n10738 ;
  assign n10740 = ~n10733 & ~n10739 ;
  assign n10741 = ~\s11_msel_arb2_state_reg[1]/NET0131  & ~n4269 ;
  assign n10742 = ~\s11_msel_arb2_state_reg[0]/NET0131  & ~n4267 ;
  assign n10743 = ~n10741 & n10742 ;
  assign n10744 = ~\s11_msel_arb2_state_reg[2]/NET0131  & n10743 ;
  assign n10745 = n4249 & ~n4252 ;
  assign n10746 = n4267 & ~n10745 ;
  assign n10747 = ~n4262 & n5879 ;
  assign n10748 = ~\s11_msel_arb2_state_reg[2]/NET0131  & n10747 ;
  assign n10749 = ~n10746 & n10748 ;
  assign n10750 = ~n10744 & ~n10749 ;
  assign n10751 = ~n10740 & n10750 ;
  assign n10752 = ~n10731 & n10751 ;
  assign n10753 = n4287 & ~n4292 ;
  assign n10754 = ~n4295 & n10753 ;
  assign n10755 = ~n4284 & ~n4308 ;
  assign n10756 = ~\s11_msel_arb3_state_reg[2]/NET0131  & ~n10755 ;
  assign n10757 = ~n4295 & ~n4300 ;
  assign n10758 = ~n10756 & n10757 ;
  assign n10759 = ~n10754 & ~n10758 ;
  assign n10760 = ~n4292 & n4312 ;
  assign n10761 = n10759 & ~n10760 ;
  assign n10762 = ~\s11_msel_arb3_state_reg[1]/NET0131  & ~n10761 ;
  assign n10763 = \s11_msel_arb3_state_reg[2]/NET0131  & ~n4287 ;
  assign n10764 = ~n4297 & n10763 ;
  assign n10765 = ~n4287 & ~n4299 ;
  assign n10766 = ~n4291 & ~n4309 ;
  assign n10767 = ~n10765 & ~n10766 ;
  assign n10768 = ~n4289 & ~n4297 ;
  assign n10769 = ~n10767 & n10768 ;
  assign n10770 = ~n10764 & ~n10769 ;
  assign n10771 = ~\s11_msel_arb3_state_reg[2]/NET0131  & ~n4289 ;
  assign n10772 = ~n4309 & n10771 ;
  assign n10773 = \s11_msel_arb3_state_reg[1]/NET0131  & ~n10772 ;
  assign n10774 = n10770 & n10773 ;
  assign n10775 = ~n10762 & ~n10774 ;
  assign n10776 = \s11_msel_arb3_state_reg[0]/NET0131  & ~n10775 ;
  assign n10777 = ~\s11_msel_arb3_state_reg[1]/NET0131  & ~n4309 ;
  assign n10778 = ~n4287 & n4300 ;
  assign n10779 = ~n10777 & ~n10778 ;
  assign n10780 = \s11_msel_arb3_state_reg[2]/NET0131  & ~n10779 ;
  assign n10781 = ~\s11_msel_arb3_state_reg[0]/NET0131  & ~n10780 ;
  assign n10782 = n4292 & ~n4309 ;
  assign n10783 = ~n4321 & ~n10782 ;
  assign n10784 = ~\s11_msel_arb3_state_reg[2]/NET0131  & ~n10783 ;
  assign n10785 = \s11_msel_arb3_state_reg[1]/NET0131  & n4287 ;
  assign n10786 = n4309 & n10785 ;
  assign n10787 = n4292 & n4300 ;
  assign n10788 = ~n10786 & n10787 ;
  assign n10789 = ~n10784 & ~n10788 ;
  assign n10790 = n10781 & n10789 ;
  assign n10791 = ~n10776 & ~n10790 ;
  assign n10792 = ~\s12_msel_arb2_state_reg[2]/NET0131  & ~n9858 ;
  assign n10793 = ~n9840 & n9847 ;
  assign n10794 = ~\s12_msel_arb2_state_reg[0]/NET0131  & n10793 ;
  assign n10795 = ~n9863 & ~n10794 ;
  assign n10796 = ~n10792 & ~n10795 ;
  assign n10797 = ~\s12_msel_arb2_state_reg[1]/NET0131  & n9847 ;
  assign n10798 = n9858 & n10797 ;
  assign n10799 = ~n10796 & ~n10798 ;
  assign n10800 = \s12_msel_arb2_state_reg[2]/NET0131  & ~n9847 ;
  assign n10801 = ~n9848 & n9858 ;
  assign n10802 = ~\s12_msel_arb2_state_reg[0]/NET0131  & n10801 ;
  assign n10803 = ~n9869 & ~n10802 ;
  assign n10804 = ~n10800 & ~n10803 ;
  assign n10805 = n6101 & n6124 ;
  assign n10806 = n6124 & n9840 ;
  assign n10807 = ~n10801 & n10806 ;
  assign n10808 = ~n10805 & ~n10807 ;
  assign n10809 = \s12_msel_arb2_state_reg[0]/NET0131  & n10808 ;
  assign n10810 = ~n10804 & ~n10809 ;
  assign n10811 = n10799 & n10810 ;
  assign n10812 = n6147 & ~n9847 ;
  assign n10813 = \s12_msel_arb2_state_reg[1]/NET0131  & ~n6110 ;
  assign n10814 = n9858 & ~n10813 ;
  assign n10815 = n6147 & n9840 ;
  assign n10816 = ~n10814 & n10815 ;
  assign n10817 = ~n10812 & ~n10816 ;
  assign n10818 = \s12_msel_arb2_state_reg[1]/NET0131  & n6096 ;
  assign n10819 = \s12_msel_arb2_state_reg[1]/NET0131  & n9848 ;
  assign n10820 = ~n10793 & n10819 ;
  assign n10821 = ~n10818 & ~n10820 ;
  assign n10822 = ~n9847 & n9848 ;
  assign n10823 = n9858 & ~n10822 ;
  assign n10824 = ~\s12_msel_arb2_state_reg[1]/NET0131  & ~n6105 ;
  assign n10825 = ~n10823 & n10824 ;
  assign n10826 = n10821 & ~n10825 ;
  assign n10827 = \s12_msel_arb2_state_reg[0]/NET0131  & ~\s12_msel_arb2_state_reg[2]/NET0131  ;
  assign n10828 = ~n10826 & n10827 ;
  assign n10829 = n10817 & ~n10828 ;
  assign n10830 = ~n10811 & n10829 ;
  assign n10831 = ~n4356 & ~n6201 ;
  assign n10832 = ~\s12_msel_arb3_state_reg[2]/NET0131  & ~n10831 ;
  assign n10833 = ~n4339 & ~n10832 ;
  assign n10834 = n4337 & ~n4349 ;
  assign n10835 = n10833 & n10834 ;
  assign n10836 = \s12_msel_arb3_state_reg[2]/NET0131  & ~n4338 ;
  assign n10837 = ~n4354 & n10831 ;
  assign n10838 = ~n10836 & n10837 ;
  assign n10839 = ~n4334 & n4339 ;
  assign n10840 = ~n4354 & n4359 ;
  assign n10841 = n4349 & ~n10840 ;
  assign n10842 = n10839 & ~n10841 ;
  assign n10843 = ~n10838 & ~n10842 ;
  assign n10844 = ~n10835 & n10843 ;
  assign n10845 = ~\s12_msel_arb3_state_reg[1]/NET0131  & ~n10844 ;
  assign n10846 = \rf_conf12_reg[13]/NET0131  & ~\s12_msel_arb3_state_reg[0]/NET0131  ;
  assign n10847 = n4347 & n10846 ;
  assign n10848 = \s12_msel_arb3_state_reg[2]/NET0131  & ~n4359 ;
  assign n10849 = ~n4337 & n4354 ;
  assign n10850 = ~n10848 & ~n10849 ;
  assign n10851 = ~n10847 & ~n10850 ;
  assign n10852 = ~n4359 & ~n4367 ;
  assign n10853 = ~n4353 & n6214 ;
  assign n10854 = ~n10852 & ~n10853 ;
  assign n10855 = ~n4348 & ~n4351 ;
  assign n10856 = ~n10854 & n10855 ;
  assign n10857 = ~n10851 & ~n10856 ;
  assign n10858 = ~n4346 & ~n10857 ;
  assign n10859 = ~n4337 & ~n4351 ;
  assign n10860 = n4368 & n10859 ;
  assign n10861 = \s12_msel_arb3_state_reg[1]/NET0131  & ~n10860 ;
  assign n10862 = ~n10858 & n10861 ;
  assign n10863 = ~n10845 & ~n10862 ;
  assign n10864 = n9876 & ~n9893 ;
  assign n10865 = \s13_msel_arb2_state_reg[1]/NET0131  & ~n10864 ;
  assign n10866 = ~\s13_msel_arb2_state_reg[1]/NET0131  & ~n9893 ;
  assign n10867 = \s13_msel_arb2_state_reg[2]/NET0131  & ~n10866 ;
  assign n10868 = ~n10865 & ~n10867 ;
  assign n10869 = ~\s13_msel_arb2_state_reg[0]/NET0131  & n10868 ;
  assign n10870 = \s13_msel_arb2_state_reg[1]/NET0131  & n9893 ;
  assign n10871 = n9876 & ~n10870 ;
  assign n10872 = n9875 & ~n10871 ;
  assign n10873 = ~\s13_msel_arb2_state_reg[2]/NET0131  & ~n9876 ;
  assign n10874 = n9892 & ~n10873 ;
  assign n10875 = ~\s13_msel_arb2_state_reg[0]/NET0131  & n10874 ;
  assign n10876 = ~n10872 & n10875 ;
  assign n10877 = ~n10869 & ~n10876 ;
  assign n10878 = ~n6393 & n10864 ;
  assign n10879 = ~n6396 & ~n6405 ;
  assign n10880 = ~\s13_msel_arb2_state_reg[2]/NET0131  & ~n10879 ;
  assign n10881 = ~n6393 & ~n9875 ;
  assign n10882 = ~n10880 & n10881 ;
  assign n10883 = ~n10878 & ~n10882 ;
  assign n10884 = n9888 & ~n9893 ;
  assign n10885 = \s13_msel_arb2_state_reg[1]/NET0131  & ~n10884 ;
  assign n10886 = n10883 & n10885 ;
  assign n10887 = ~n6403 & n6417 ;
  assign n10888 = \s13_msel_arb2_state_reg[0]/NET0131  & ~n10887 ;
  assign n10889 = n9875 & ~n9876 ;
  assign n10890 = \s13_msel_arb2_state_reg[0]/NET0131  & n9892 ;
  assign n10891 = ~n10889 & n10890 ;
  assign n10892 = ~n10888 & ~n10891 ;
  assign n10893 = ~n10886 & ~n10892 ;
  assign n10894 = n10877 & ~n10893 ;
  assign n10895 = ~n9892 & n9893 ;
  assign n10896 = n9876 & ~n10895 ;
  assign n10897 = \rf_conf13_reg[1]/NET0131  & ~\s13_msel_arb2_state_reg[0]/NET0131  ;
  assign n10898 = n2876 & n10897 ;
  assign n10899 = n6452 & ~n10898 ;
  assign n10900 = ~n10896 & n10899 ;
  assign n10901 = ~n10894 & ~n10900 ;
  assign n10902 = ~n3871 & ~n6495 ;
  assign n10903 = ~\s13_msel_arb3_state_reg[2]/NET0131  & ~n10902 ;
  assign n10904 = ~n3854 & ~n10903 ;
  assign n10905 = n3852 & ~n3864 ;
  assign n10906 = n10904 & n10905 ;
  assign n10907 = \s13_msel_arb3_state_reg[2]/NET0131  & ~n3853 ;
  assign n10908 = ~n3869 & n10902 ;
  assign n10909 = ~n10907 & n10908 ;
  assign n10910 = ~n3849 & n3854 ;
  assign n10911 = ~n3869 & n3874 ;
  assign n10912 = n3864 & ~n10911 ;
  assign n10913 = n10910 & ~n10912 ;
  assign n10914 = ~n10909 & ~n10913 ;
  assign n10915 = ~n10906 & n10914 ;
  assign n10916 = ~\s13_msel_arb3_state_reg[1]/NET0131  & ~n10915 ;
  assign n10917 = \rf_conf13_reg[13]/NET0131  & ~\s13_msel_arb3_state_reg[0]/NET0131  ;
  assign n10918 = n3862 & n10917 ;
  assign n10919 = \s13_msel_arb3_state_reg[2]/NET0131  & ~n3874 ;
  assign n10920 = ~n3852 & n3869 ;
  assign n10921 = ~n10919 & ~n10920 ;
  assign n10922 = ~n10918 & ~n10921 ;
  assign n10923 = ~n3874 & ~n3882 ;
  assign n10924 = ~n3868 & n6508 ;
  assign n10925 = ~n10923 & ~n10924 ;
  assign n10926 = ~n3863 & ~n3866 ;
  assign n10927 = ~n10925 & n10926 ;
  assign n10928 = ~n10922 & ~n10927 ;
  assign n10929 = ~n3861 & ~n10928 ;
  assign n10930 = ~n3852 & ~n3866 ;
  assign n10931 = n3883 & n10930 ;
  assign n10932 = \s13_msel_arb3_state_reg[1]/NET0131  & ~n10931 ;
  assign n10933 = ~n10929 & n10932 ;
  assign n10934 = ~n10916 & ~n10933 ;
  assign n10935 = ~n3918 & ~n6703 ;
  assign n10936 = ~\s14_msel_arb2_state_reg[2]/NET0131  & ~n10935 ;
  assign n10937 = ~n3906 & ~n10936 ;
  assign n10938 = n3904 & ~n3914 ;
  assign n10939 = n10937 & n10938 ;
  assign n10940 = \s14_msel_arb2_state_reg[2]/NET0131  & ~n3905 ;
  assign n10941 = ~n3917 & n10935 ;
  assign n10942 = ~n10940 & n10941 ;
  assign n10943 = ~n3902 & n3906 ;
  assign n10944 = ~n3917 & n3920 ;
  assign n10945 = n3914 & ~n10944 ;
  assign n10946 = n10943 & ~n10945 ;
  assign n10947 = ~n10942 & ~n10946 ;
  assign n10948 = ~n10939 & n10947 ;
  assign n10949 = ~\s14_msel_arb2_state_reg[1]/NET0131  & ~n10948 ;
  assign n10950 = \rf_conf14_reg[13]/NET0131  & ~\s14_msel_arb2_state_reg[0]/NET0131  ;
  assign n10951 = n2933 & n10950 ;
  assign n10952 = \s14_msel_arb2_state_reg[2]/NET0131  & ~n3920 ;
  assign n10953 = ~n3904 & n3917 ;
  assign n10954 = ~n10952 & ~n10953 ;
  assign n10955 = ~n10951 & ~n10954 ;
  assign n10956 = ~n3920 & ~n3928 ;
  assign n10957 = ~n3916 & n6716 ;
  assign n10958 = ~n10956 & ~n10957 ;
  assign n10959 = ~n3913 & ~n3915 ;
  assign n10960 = ~n10958 & n10959 ;
  assign n10961 = ~n10955 & ~n10960 ;
  assign n10962 = ~n3912 & ~n10961 ;
  assign n10963 = ~n3904 & ~n3915 ;
  assign n10964 = n3929 & n10963 ;
  assign n10965 = \s14_msel_arb2_state_reg[1]/NET0131  & ~n10964 ;
  assign n10966 = ~n10962 & n10965 ;
  assign n10967 = ~n10949 & ~n10966 ;
  assign n10968 = n4392 & ~n4397 ;
  assign n10969 = ~n4400 & n10968 ;
  assign n10970 = ~n4389 & ~n4413 ;
  assign n10971 = ~\s14_msel_arb3_state_reg[2]/NET0131  & ~n10970 ;
  assign n10972 = ~n4400 & ~n4405 ;
  assign n10973 = ~n10971 & n10972 ;
  assign n10974 = ~n10969 & ~n10973 ;
  assign n10975 = ~n4397 & n4417 ;
  assign n10976 = n10974 & ~n10975 ;
  assign n10977 = ~\s14_msel_arb3_state_reg[1]/NET0131  & ~n10976 ;
  assign n10978 = \s14_msel_arb3_state_reg[2]/NET0131  & ~n4392 ;
  assign n10979 = ~n4402 & n10978 ;
  assign n10980 = ~n4392 & ~n4404 ;
  assign n10981 = ~n4396 & ~n4414 ;
  assign n10982 = ~n10980 & ~n10981 ;
  assign n10983 = ~n4394 & ~n4402 ;
  assign n10984 = ~n10982 & n10983 ;
  assign n10985 = ~n10979 & ~n10984 ;
  assign n10986 = ~\s14_msel_arb3_state_reg[2]/NET0131  & ~n4394 ;
  assign n10987 = ~n4414 & n10986 ;
  assign n10988 = \s14_msel_arb3_state_reg[1]/NET0131  & ~n10987 ;
  assign n10989 = n10985 & n10988 ;
  assign n10990 = ~n10977 & ~n10989 ;
  assign n10991 = \s14_msel_arb3_state_reg[0]/NET0131  & ~n10990 ;
  assign n10992 = ~\s14_msel_arb3_state_reg[1]/NET0131  & ~n4414 ;
  assign n10993 = ~n4392 & n4405 ;
  assign n10994 = ~n10992 & ~n10993 ;
  assign n10995 = \s14_msel_arb3_state_reg[2]/NET0131  & ~n10994 ;
  assign n10996 = ~\s14_msel_arb3_state_reg[0]/NET0131  & ~n10995 ;
  assign n10997 = n4397 & ~n4414 ;
  assign n10998 = ~n4426 & ~n10997 ;
  assign n10999 = ~\s14_msel_arb3_state_reg[2]/NET0131  & ~n10998 ;
  assign n11000 = \s14_msel_arb3_state_reg[1]/NET0131  & n4392 ;
  assign n11001 = n4414 & n11000 ;
  assign n11002 = n4397 & n4405 ;
  assign n11003 = ~n11001 & n11002 ;
  assign n11004 = ~n10999 & ~n11003 ;
  assign n11005 = n10996 & n11004 ;
  assign n11006 = ~n10991 & ~n11005 ;
  assign n11007 = \rf_conf1_reg[5]/NET0131  & ~\s1_msel_arb2_state_reg[0]/NET0131  ;
  assign n11008 = n3371 & n11007 ;
  assign n11009 = n4440 & ~n11008 ;
  assign n11010 = \rf_conf1_reg[7]/NET0131  & \s1_msel_arb2_state_reg[0]/NET0131  ;
  assign n11011 = n3369 & n11010 ;
  assign n11012 = ~\s1_msel_arb2_state_reg[2]/NET0131  & ~n11011 ;
  assign n11013 = ~n11009 & n11012 ;
  assign n11014 = ~\s1_msel_arb2_state_reg[1]/NET0131  & ~n4448 ;
  assign n11015 = n4460 & ~n11014 ;
  assign n11016 = n4443 & n11012 ;
  assign n11017 = ~n11015 & n11016 ;
  assign n11018 = ~n11013 & ~n11017 ;
  assign n11019 = \s1_msel_arb2_state_reg[2]/NET0131  & ~n7194 ;
  assign n11020 = ~n4442 & n11019 ;
  assign n11021 = \s1_msel_arb2_state_reg[1]/NET0131  & ~n11020 ;
  assign n11022 = ~n4440 & n4458 ;
  assign n11023 = \s1_msel_arb2_state_reg[1]/NET0131  & n4460 ;
  assign n11024 = ~n11022 & n11023 ;
  assign n11025 = ~n11021 & ~n11024 ;
  assign n11026 = n11018 & ~n11025 ;
  assign n11027 = ~n4458 & n4460 ;
  assign n11028 = n4443 & ~n11027 ;
  assign n11029 = ~n4438 & n7206 ;
  assign n11030 = ~\s1_msel_arb2_state_reg[2]/NET0131  & ~n4460 ;
  assign n11031 = ~\s1_msel_arb2_state_reg[0]/NET0131  & ~\s1_msel_arb2_state_reg[1]/NET0131  ;
  assign n11032 = n4440 & n11031 ;
  assign n11033 = ~n11030 & n11032 ;
  assign n11034 = ~n11029 & ~n11033 ;
  assign n11035 = ~n11028 & ~n11034 ;
  assign n11036 = ~\s1_msel_arb2_state_reg[1]/NET0131  & ~n4460 ;
  assign n11037 = ~\s1_msel_arb2_state_reg[0]/NET0131  & ~n4458 ;
  assign n11038 = ~n11036 & n11037 ;
  assign n11039 = ~\s1_msel_arb2_state_reg[2]/NET0131  & n11038 ;
  assign n11040 = n4440 & ~n4443 ;
  assign n11041 = n4458 & ~n11040 ;
  assign n11042 = ~n4453 & n7205 ;
  assign n11043 = ~\s1_msel_arb2_state_reg[2]/NET0131  & n11042 ;
  assign n11044 = ~n11041 & n11043 ;
  assign n11045 = ~n11039 & ~n11044 ;
  assign n11046 = ~n11035 & n11045 ;
  assign n11047 = ~n11026 & n11046 ;
  assign n11048 = n4478 & ~n4483 ;
  assign n11049 = ~n4486 & n11048 ;
  assign n11050 = ~n4475 & ~n4499 ;
  assign n11051 = ~\s1_msel_arb3_state_reg[2]/NET0131  & ~n11050 ;
  assign n11052 = ~n4486 & ~n4491 ;
  assign n11053 = ~n11051 & n11052 ;
  assign n11054 = ~n11049 & ~n11053 ;
  assign n11055 = ~n4483 & n4503 ;
  assign n11056 = n11054 & ~n11055 ;
  assign n11057 = ~\s1_msel_arb3_state_reg[1]/NET0131  & ~n11056 ;
  assign n11058 = \s1_msel_arb3_state_reg[2]/NET0131  & ~n4478 ;
  assign n11059 = ~n4488 & n11058 ;
  assign n11060 = ~n4478 & ~n4490 ;
  assign n11061 = ~n4482 & ~n4500 ;
  assign n11062 = ~n11060 & ~n11061 ;
  assign n11063 = ~n4480 & ~n4488 ;
  assign n11064 = ~n11062 & n11063 ;
  assign n11065 = ~n11059 & ~n11064 ;
  assign n11066 = ~\s1_msel_arb3_state_reg[2]/NET0131  & ~n4480 ;
  assign n11067 = ~n4500 & n11066 ;
  assign n11068 = \s1_msel_arb3_state_reg[1]/NET0131  & ~n11067 ;
  assign n11069 = n11065 & n11068 ;
  assign n11070 = ~n11057 & ~n11069 ;
  assign n11071 = \s1_msel_arb3_state_reg[0]/NET0131  & ~n11070 ;
  assign n11072 = ~\s1_msel_arb3_state_reg[1]/NET0131  & ~n4500 ;
  assign n11073 = ~n4478 & n4491 ;
  assign n11074 = ~n11072 & ~n11073 ;
  assign n11075 = \s1_msel_arb3_state_reg[2]/NET0131  & ~n11074 ;
  assign n11076 = ~\s1_msel_arb3_state_reg[0]/NET0131  & ~n11075 ;
  assign n11077 = n4483 & ~n4500 ;
  assign n11078 = ~n4512 & ~n11077 ;
  assign n11079 = ~\s1_msel_arb3_state_reg[2]/NET0131  & ~n11078 ;
  assign n11080 = \s1_msel_arb3_state_reg[1]/NET0131  & n4478 ;
  assign n11081 = n4500 & n11080 ;
  assign n11082 = n4483 & n4491 ;
  assign n11083 = ~n11081 & n11082 ;
  assign n11084 = ~n11079 & ~n11083 ;
  assign n11085 = n11076 & n11084 ;
  assign n11086 = ~n11071 & ~n11085 ;
  assign n11087 = n9903 & ~n9920 ;
  assign n11088 = \s2_msel_arb2_state_reg[1]/NET0131  & ~n11087 ;
  assign n11089 = ~\s2_msel_arb2_state_reg[1]/NET0131  & ~n9920 ;
  assign n11090 = \s2_msel_arb2_state_reg[2]/NET0131  & ~n11089 ;
  assign n11091 = ~n11088 & ~n11090 ;
  assign n11092 = ~\s2_msel_arb2_state_reg[0]/NET0131  & n11091 ;
  assign n11093 = \s2_msel_arb2_state_reg[1]/NET0131  & n9920 ;
  assign n11094 = n9903 & ~n11093 ;
  assign n11095 = n9902 & ~n11094 ;
  assign n11096 = ~\s2_msel_arb2_state_reg[2]/NET0131  & ~n9903 ;
  assign n11097 = n9919 & ~n11096 ;
  assign n11098 = ~\s2_msel_arb2_state_reg[0]/NET0131  & n11097 ;
  assign n11099 = ~n11095 & n11098 ;
  assign n11100 = ~n11092 & ~n11099 ;
  assign n11101 = ~n7438 & n11087 ;
  assign n11102 = ~n7441 & ~n7450 ;
  assign n11103 = ~\s2_msel_arb2_state_reg[2]/NET0131  & ~n11102 ;
  assign n11104 = ~n7438 & ~n9902 ;
  assign n11105 = ~n11103 & n11104 ;
  assign n11106 = ~n11101 & ~n11105 ;
  assign n11107 = n9915 & ~n9920 ;
  assign n11108 = \s2_msel_arb2_state_reg[1]/NET0131  & ~n11107 ;
  assign n11109 = n11106 & n11108 ;
  assign n11110 = ~n7448 & n7462 ;
  assign n11111 = \s2_msel_arb2_state_reg[0]/NET0131  & ~n11110 ;
  assign n11112 = n9902 & ~n9903 ;
  assign n11113 = \s2_msel_arb2_state_reg[0]/NET0131  & n9919 ;
  assign n11114 = ~n11112 & n11113 ;
  assign n11115 = ~n11111 & ~n11114 ;
  assign n11116 = ~n11109 & ~n11115 ;
  assign n11117 = n11100 & ~n11116 ;
  assign n11118 = ~n9919 & n9920 ;
  assign n11119 = n9903 & ~n11118 ;
  assign n11120 = \rf_conf2_reg[1]/NET0131  & ~\s2_msel_arb2_state_reg[0]/NET0131  ;
  assign n11121 = n3451 & n11120 ;
  assign n11122 = n7497 & ~n11121 ;
  assign n11123 = ~n11119 & n11122 ;
  assign n11124 = ~n11117 & ~n11123 ;
  assign n11125 = ~n3971 & ~n7540 ;
  assign n11126 = ~\s2_msel_arb3_state_reg[2]/NET0131  & ~n11125 ;
  assign n11127 = ~n3954 & ~n11126 ;
  assign n11128 = n3952 & ~n3964 ;
  assign n11129 = n11127 & n11128 ;
  assign n11130 = \s2_msel_arb3_state_reg[2]/NET0131  & ~n3953 ;
  assign n11131 = ~n3969 & n11125 ;
  assign n11132 = ~n11130 & n11131 ;
  assign n11133 = ~n3949 & n3954 ;
  assign n11134 = ~n3969 & n3974 ;
  assign n11135 = n3964 & ~n11134 ;
  assign n11136 = n11133 & ~n11135 ;
  assign n11137 = ~n11132 & ~n11136 ;
  assign n11138 = ~n11129 & n11137 ;
  assign n11139 = ~\s2_msel_arb3_state_reg[1]/NET0131  & ~n11138 ;
  assign n11140 = \rf_conf2_reg[13]/NET0131  & ~\s2_msel_arb3_state_reg[0]/NET0131  ;
  assign n11141 = n3962 & n11140 ;
  assign n11142 = \s2_msel_arb3_state_reg[2]/NET0131  & ~n3974 ;
  assign n11143 = ~n3952 & n3969 ;
  assign n11144 = ~n11142 & ~n11143 ;
  assign n11145 = ~n11141 & ~n11144 ;
  assign n11146 = ~n3974 & ~n3982 ;
  assign n11147 = ~n3968 & n7553 ;
  assign n11148 = ~n11146 & ~n11147 ;
  assign n11149 = ~n3963 & ~n3966 ;
  assign n11150 = ~n11148 & n11149 ;
  assign n11151 = ~n11145 & ~n11150 ;
  assign n11152 = ~n3961 & ~n11151 ;
  assign n11153 = ~n3952 & ~n3966 ;
  assign n11154 = n3983 & n11153 ;
  assign n11155 = \s2_msel_arb3_state_reg[1]/NET0131  & ~n11154 ;
  assign n11156 = ~n11152 & n11155 ;
  assign n11157 = ~n11139 & ~n11156 ;
  assign n11158 = \rf_conf3_reg[5]/NET0131  & ~\s3_msel_arb2_state_reg[0]/NET0131  ;
  assign n11159 = n3082 & n11158 ;
  assign n11160 = n4004 & ~n11159 ;
  assign n11161 = \rf_conf3_reg[7]/NET0131  & \s3_msel_arb2_state_reg[0]/NET0131  ;
  assign n11162 = n3076 & n11161 ;
  assign n11163 = ~\s3_msel_arb2_state_reg[2]/NET0131  & ~n11162 ;
  assign n11164 = ~n11160 & n11163 ;
  assign n11165 = ~\s3_msel_arb2_state_reg[1]/NET0131  & ~n4012 ;
  assign n11166 = n4024 & ~n11165 ;
  assign n11167 = n4007 & n11163 ;
  assign n11168 = ~n11166 & n11167 ;
  assign n11169 = ~n11164 & ~n11168 ;
  assign n11170 = \s3_msel_arb2_state_reg[2]/NET0131  & ~n7761 ;
  assign n11171 = ~n4006 & n11170 ;
  assign n11172 = \s3_msel_arb2_state_reg[1]/NET0131  & ~n11171 ;
  assign n11173 = ~n4004 & n4022 ;
  assign n11174 = \s3_msel_arb2_state_reg[1]/NET0131  & n4024 ;
  assign n11175 = ~n11173 & n11174 ;
  assign n11176 = ~n11172 & ~n11175 ;
  assign n11177 = n11169 & ~n11176 ;
  assign n11178 = ~n4022 & n4024 ;
  assign n11179 = n4007 & ~n11178 ;
  assign n11180 = ~n4002 & n7773 ;
  assign n11181 = ~\s3_msel_arb2_state_reg[2]/NET0131  & ~n4024 ;
  assign n11182 = ~\s3_msel_arb2_state_reg[0]/NET0131  & ~\s3_msel_arb2_state_reg[1]/NET0131  ;
  assign n11183 = n4004 & n11182 ;
  assign n11184 = ~n11181 & n11183 ;
  assign n11185 = ~n11180 & ~n11184 ;
  assign n11186 = ~n11179 & ~n11185 ;
  assign n11187 = ~\s3_msel_arb2_state_reg[1]/NET0131  & ~n4024 ;
  assign n11188 = ~\s3_msel_arb2_state_reg[0]/NET0131  & ~n4022 ;
  assign n11189 = ~n11187 & n11188 ;
  assign n11190 = ~\s3_msel_arb2_state_reg[2]/NET0131  & n11189 ;
  assign n11191 = n4004 & ~n4007 ;
  assign n11192 = n4022 & ~n11191 ;
  assign n11193 = ~n4017 & n7772 ;
  assign n11194 = ~\s3_msel_arb2_state_reg[2]/NET0131  & n11193 ;
  assign n11195 = ~n11192 & n11194 ;
  assign n11196 = ~n11190 & ~n11195 ;
  assign n11197 = ~n11186 & n11196 ;
  assign n11198 = ~n11177 & n11197 ;
  assign n11199 = n4529 & ~n4534 ;
  assign n11200 = ~n4537 & n11199 ;
  assign n11201 = ~n4526 & ~n4550 ;
  assign n11202 = ~\s3_msel_arb3_state_reg[2]/NET0131  & ~n11201 ;
  assign n11203 = ~n4537 & ~n4542 ;
  assign n11204 = ~n11202 & n11203 ;
  assign n11205 = ~n11200 & ~n11204 ;
  assign n11206 = ~n4534 & n4554 ;
  assign n11207 = n11205 & ~n11206 ;
  assign n11208 = ~\s3_msel_arb3_state_reg[1]/NET0131  & ~n11207 ;
  assign n11209 = \s3_msel_arb3_state_reg[2]/NET0131  & ~n4529 ;
  assign n11210 = ~n4539 & n11209 ;
  assign n11211 = ~n4529 & ~n4541 ;
  assign n11212 = ~n4533 & ~n4551 ;
  assign n11213 = ~n11211 & ~n11212 ;
  assign n11214 = ~n4531 & ~n4539 ;
  assign n11215 = ~n11213 & n11214 ;
  assign n11216 = ~n11210 & ~n11215 ;
  assign n11217 = ~\s3_msel_arb3_state_reg[2]/NET0131  & ~n4531 ;
  assign n11218 = ~n4551 & n11217 ;
  assign n11219 = \s3_msel_arb3_state_reg[1]/NET0131  & ~n11218 ;
  assign n11220 = n11216 & n11219 ;
  assign n11221 = ~n11208 & ~n11220 ;
  assign n11222 = \s3_msel_arb3_state_reg[0]/NET0131  & ~n11221 ;
  assign n11223 = ~\s3_msel_arb3_state_reg[1]/NET0131  & ~n4551 ;
  assign n11224 = ~n4529 & n4542 ;
  assign n11225 = ~n11223 & ~n11224 ;
  assign n11226 = \s3_msel_arb3_state_reg[2]/NET0131  & ~n11225 ;
  assign n11227 = ~\s3_msel_arb3_state_reg[0]/NET0131  & ~n11226 ;
  assign n11228 = n4534 & ~n4551 ;
  assign n11229 = ~n4563 & ~n11228 ;
  assign n11230 = ~\s3_msel_arb3_state_reg[2]/NET0131  & ~n11229 ;
  assign n11231 = \s3_msel_arb3_state_reg[1]/NET0131  & n4529 ;
  assign n11232 = n4551 & n11231 ;
  assign n11233 = n4534 & n4542 ;
  assign n11234 = ~n11232 & n11233 ;
  assign n11235 = ~n11230 & ~n11234 ;
  assign n11236 = n11227 & n11235 ;
  assign n11237 = ~n11222 & ~n11236 ;
  assign n11238 = n9930 & ~n9947 ;
  assign n11239 = \s4_msel_arb2_state_reg[1]/NET0131  & ~n11238 ;
  assign n11240 = ~\s4_msel_arb2_state_reg[1]/NET0131  & ~n9947 ;
  assign n11241 = \s4_msel_arb2_state_reg[2]/NET0131  & ~n11240 ;
  assign n11242 = ~n11239 & ~n11241 ;
  assign n11243 = ~\s4_msel_arb2_state_reg[0]/NET0131  & n11242 ;
  assign n11244 = \s4_msel_arb2_state_reg[1]/NET0131  & n9947 ;
  assign n11245 = n9930 & ~n11244 ;
  assign n11246 = n9929 & ~n11245 ;
  assign n11247 = ~\s4_msel_arb2_state_reg[2]/NET0131  & ~n9930 ;
  assign n11248 = n9946 & ~n11247 ;
  assign n11249 = ~\s4_msel_arb2_state_reg[0]/NET0131  & n11248 ;
  assign n11250 = ~n11246 & n11249 ;
  assign n11251 = ~n11243 & ~n11250 ;
  assign n11252 = ~n8007 & n11238 ;
  assign n11253 = ~n8010 & ~n8019 ;
  assign n11254 = ~\s4_msel_arb2_state_reg[2]/NET0131  & ~n11253 ;
  assign n11255 = ~n8007 & ~n9929 ;
  assign n11256 = ~n11254 & n11255 ;
  assign n11257 = ~n11252 & ~n11256 ;
  assign n11258 = n9942 & ~n9947 ;
  assign n11259 = \s4_msel_arb2_state_reg[1]/NET0131  & ~n11258 ;
  assign n11260 = n11257 & n11259 ;
  assign n11261 = ~n8017 & n8031 ;
  assign n11262 = \s4_msel_arb2_state_reg[0]/NET0131  & ~n11261 ;
  assign n11263 = n9929 & ~n9930 ;
  assign n11264 = \s4_msel_arb2_state_reg[0]/NET0131  & n9946 ;
  assign n11265 = ~n11263 & n11264 ;
  assign n11266 = ~n11262 & ~n11265 ;
  assign n11267 = ~n11260 & ~n11266 ;
  assign n11268 = n11251 & ~n11267 ;
  assign n11269 = ~n9946 & n9947 ;
  assign n11270 = n9930 & ~n11269 ;
  assign n11271 = \rf_conf4_reg[1]/NET0131  & ~\s4_msel_arb2_state_reg[0]/NET0131  ;
  assign n11272 = n3133 & n11271 ;
  assign n11273 = n8066 & ~n11272 ;
  assign n11274 = ~n11270 & n11273 ;
  assign n11275 = ~n11268 & ~n11274 ;
  assign n11276 = n4042 & ~n4047 ;
  assign n11277 = ~n4050 & n11276 ;
  assign n11278 = ~n4039 & ~n4063 ;
  assign n11279 = ~\s4_msel_arb3_state_reg[2]/NET0131  & ~n11278 ;
  assign n11280 = ~n4050 & ~n4055 ;
  assign n11281 = ~n11279 & n11280 ;
  assign n11282 = ~n11277 & ~n11281 ;
  assign n11283 = ~n4047 & n4067 ;
  assign n11284 = n11282 & ~n11283 ;
  assign n11285 = ~\s4_msel_arb3_state_reg[1]/NET0131  & ~n11284 ;
  assign n11286 = \s4_msel_arb3_state_reg[2]/NET0131  & ~n4042 ;
  assign n11287 = ~n4052 & n11286 ;
  assign n11288 = ~n4042 & ~n4054 ;
  assign n11289 = ~n4046 & ~n4064 ;
  assign n11290 = ~n11288 & ~n11289 ;
  assign n11291 = ~n4044 & ~n4052 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = ~n11287 & ~n11292 ;
  assign n11294 = ~\s4_msel_arb3_state_reg[2]/NET0131  & ~n4044 ;
  assign n11295 = ~n4064 & n11294 ;
  assign n11296 = \s4_msel_arb3_state_reg[1]/NET0131  & ~n11295 ;
  assign n11297 = n11293 & n11296 ;
  assign n11298 = ~n11285 & ~n11297 ;
  assign n11299 = \s4_msel_arb3_state_reg[0]/NET0131  & ~n11298 ;
  assign n11300 = ~\s4_msel_arb3_state_reg[1]/NET0131  & ~n4064 ;
  assign n11301 = ~n4042 & n4055 ;
  assign n11302 = ~n11300 & ~n11301 ;
  assign n11303 = \s4_msel_arb3_state_reg[2]/NET0131  & ~n11302 ;
  assign n11304 = ~\s4_msel_arb3_state_reg[0]/NET0131  & ~n11303 ;
  assign n11305 = n4047 & ~n4064 ;
  assign n11306 = ~n4076 & ~n11305 ;
  assign n11307 = ~\s4_msel_arb3_state_reg[2]/NET0131  & ~n11306 ;
  assign n11308 = \s4_msel_arb3_state_reg[1]/NET0131  & n4042 ;
  assign n11309 = n4064 & n11308 ;
  assign n11310 = n4047 & n4055 ;
  assign n11311 = ~n11309 & n11310 ;
  assign n11312 = ~n11307 & ~n11311 ;
  assign n11313 = n11304 & n11312 ;
  assign n11314 = ~n11299 & ~n11313 ;
  assign n11315 = \rf_conf5_reg[5]/NET0131  & ~\s5_msel_arb2_state_reg[0]/NET0131  ;
  assign n11316 = n3206 & n11315 ;
  assign n11317 = n4577 & ~n11316 ;
  assign n11318 = \rf_conf5_reg[7]/NET0131  & \s5_msel_arb2_state_reg[0]/NET0131  ;
  assign n11319 = n3200 & n11318 ;
  assign n11320 = ~\s5_msel_arb2_state_reg[2]/NET0131  & ~n11319 ;
  assign n11321 = ~n11317 & n11320 ;
  assign n11322 = ~\s5_msel_arb2_state_reg[1]/NET0131  & ~n4585 ;
  assign n11323 = n4597 & ~n11322 ;
  assign n11324 = n4580 & n11320 ;
  assign n11325 = ~n11323 & n11324 ;
  assign n11326 = ~n11321 & ~n11325 ;
  assign n11327 = \s5_msel_arb2_state_reg[2]/NET0131  & ~n8317 ;
  assign n11328 = ~n4579 & n11327 ;
  assign n11329 = \s5_msel_arb2_state_reg[1]/NET0131  & ~n11328 ;
  assign n11330 = ~n4577 & n4595 ;
  assign n11331 = \s5_msel_arb2_state_reg[1]/NET0131  & n4597 ;
  assign n11332 = ~n11330 & n11331 ;
  assign n11333 = ~n11329 & ~n11332 ;
  assign n11334 = n11326 & ~n11333 ;
  assign n11335 = ~n4595 & n4597 ;
  assign n11336 = n4580 & ~n11335 ;
  assign n11337 = ~n4575 & n8329 ;
  assign n11338 = ~\s5_msel_arb2_state_reg[2]/NET0131  & ~n4597 ;
  assign n11339 = ~\s5_msel_arb2_state_reg[0]/NET0131  & ~\s5_msel_arb2_state_reg[1]/NET0131  ;
  assign n11340 = n4577 & n11339 ;
  assign n11341 = ~n11338 & n11340 ;
  assign n11342 = ~n11337 & ~n11341 ;
  assign n11343 = ~n11336 & ~n11342 ;
  assign n11344 = ~\s5_msel_arb2_state_reg[1]/NET0131  & ~n4597 ;
  assign n11345 = ~\s5_msel_arb2_state_reg[0]/NET0131  & ~n4595 ;
  assign n11346 = ~n11344 & n11345 ;
  assign n11347 = ~\s5_msel_arb2_state_reg[2]/NET0131  & n11346 ;
  assign n11348 = n4577 & ~n4580 ;
  assign n11349 = n4595 & ~n11348 ;
  assign n11350 = ~n4590 & n8328 ;
  assign n11351 = ~\s5_msel_arb2_state_reg[2]/NET0131  & n11350 ;
  assign n11352 = ~n11349 & n11351 ;
  assign n11353 = ~n11347 & ~n11352 ;
  assign n11354 = ~n11343 & n11353 ;
  assign n11355 = ~n11334 & n11354 ;
  assign n11356 = ~n4633 & ~n8371 ;
  assign n11357 = ~\s5_msel_arb3_state_reg[2]/NET0131  & ~n11356 ;
  assign n11358 = ~n4616 & ~n11357 ;
  assign n11359 = n4614 & ~n4626 ;
  assign n11360 = n11358 & n11359 ;
  assign n11361 = \s5_msel_arb3_state_reg[2]/NET0131  & ~n4615 ;
  assign n11362 = ~n4631 & n11356 ;
  assign n11363 = ~n11361 & n11362 ;
  assign n11364 = ~n4611 & n4616 ;
  assign n11365 = ~n4631 & n4636 ;
  assign n11366 = n4626 & ~n11365 ;
  assign n11367 = n11364 & ~n11366 ;
  assign n11368 = ~n11363 & ~n11367 ;
  assign n11369 = ~n11360 & n11368 ;
  assign n11370 = ~\s5_msel_arb3_state_reg[1]/NET0131  & ~n11369 ;
  assign n11371 = \rf_conf5_reg[13]/NET0131  & ~\s5_msel_arb3_state_reg[0]/NET0131  ;
  assign n11372 = n4624 & n11371 ;
  assign n11373 = \s5_msel_arb3_state_reg[2]/NET0131  & ~n4636 ;
  assign n11374 = ~n4614 & n4631 ;
  assign n11375 = ~n11373 & ~n11374 ;
  assign n11376 = ~n11372 & ~n11375 ;
  assign n11377 = ~n4636 & ~n4644 ;
  assign n11378 = ~n4630 & n8384 ;
  assign n11379 = ~n11377 & ~n11378 ;
  assign n11380 = ~n4625 & ~n4628 ;
  assign n11381 = ~n11379 & n11380 ;
  assign n11382 = ~n11376 & ~n11381 ;
  assign n11383 = ~n4623 & ~n11382 ;
  assign n11384 = ~n4614 & ~n4628 ;
  assign n11385 = n4645 & n11384 ;
  assign n11386 = \s5_msel_arb3_state_reg[1]/NET0131  & ~n11385 ;
  assign n11387 = ~n11383 & n11386 ;
  assign n11388 = ~n11370 & ~n11387 ;
  assign n11389 = \rf_conf6_reg[5]/NET0131  & ~\s6_msel_arb2_state_reg[0]/NET0131  ;
  assign n11390 = n3268 & n11389 ;
  assign n11391 = n4090 & ~n11390 ;
  assign n11392 = \rf_conf6_reg[7]/NET0131  & \s6_msel_arb2_state_reg[0]/NET0131  ;
  assign n11393 = n3262 & n11392 ;
  assign n11394 = ~\s6_msel_arb2_state_reg[2]/NET0131  & ~n11393 ;
  assign n11395 = ~n11391 & n11394 ;
  assign n11396 = ~\s6_msel_arb2_state_reg[1]/NET0131  & ~n4098 ;
  assign n11397 = n4110 & ~n11396 ;
  assign n11398 = n4093 & n11394 ;
  assign n11399 = ~n11397 & n11398 ;
  assign n11400 = ~n11395 & ~n11399 ;
  assign n11401 = \s6_msel_arb2_state_reg[2]/NET0131  & ~n8571 ;
  assign n11402 = ~n4092 & n11401 ;
  assign n11403 = \s6_msel_arb2_state_reg[1]/NET0131  & ~n11402 ;
  assign n11404 = ~n4090 & n4108 ;
  assign n11405 = \s6_msel_arb2_state_reg[1]/NET0131  & n4110 ;
  assign n11406 = ~n11404 & n11405 ;
  assign n11407 = ~n11403 & ~n11406 ;
  assign n11408 = n11400 & ~n11407 ;
  assign n11409 = ~n4108 & n4110 ;
  assign n11410 = n4093 & ~n11409 ;
  assign n11411 = ~n4088 & n8583 ;
  assign n11412 = ~\s6_msel_arb2_state_reg[2]/NET0131  & ~n4110 ;
  assign n11413 = ~\s6_msel_arb2_state_reg[0]/NET0131  & ~\s6_msel_arb2_state_reg[1]/NET0131  ;
  assign n11414 = n4090 & n11413 ;
  assign n11415 = ~n11412 & n11414 ;
  assign n11416 = ~n11411 & ~n11415 ;
  assign n11417 = ~n11410 & ~n11416 ;
  assign n11418 = ~\s6_msel_arb2_state_reg[1]/NET0131  & ~n4110 ;
  assign n11419 = ~\s6_msel_arb2_state_reg[0]/NET0131  & ~n4108 ;
  assign n11420 = ~n11418 & n11419 ;
  assign n11421 = ~\s6_msel_arb2_state_reg[2]/NET0131  & n11420 ;
  assign n11422 = n4090 & ~n4093 ;
  assign n11423 = n4108 & ~n11422 ;
  assign n11424 = ~n4103 & n8582 ;
  assign n11425 = ~\s6_msel_arb2_state_reg[2]/NET0131  & n11424 ;
  assign n11426 = ~n11423 & n11425 ;
  assign n11427 = ~n11421 & ~n11426 ;
  assign n11428 = ~n11417 & n11427 ;
  assign n11429 = ~n11408 & n11428 ;
  assign n11430 = \s6_msel_arb3_state_reg[0]/NET0131  & \s6_msel_arb3_state_reg[2]/NET0131  ;
  assign n11431 = ~n4687 & ~n8625 ;
  assign n11432 = ~\s6_msel_arb3_state_reg[2]/NET0131  & ~n11431 ;
  assign n11433 = ~n11430 & ~n11432 ;
  assign n11434 = n4668 & ~n4680 ;
  assign n11435 = n11433 & n11434 ;
  assign n11436 = \s6_msel_arb3_state_reg[2]/NET0131  & ~n4669 ;
  assign n11437 = ~n4685 & n11431 ;
  assign n11438 = ~n11436 & n11437 ;
  assign n11439 = ~n4665 & n4670 ;
  assign n11440 = ~n4685 & n4690 ;
  assign n11441 = n4680 & ~n11440 ;
  assign n11442 = n11439 & ~n11441 ;
  assign n11443 = ~n11438 & ~n11442 ;
  assign n11444 = ~n11435 & n11443 ;
  assign n11445 = ~\s6_msel_arb3_state_reg[1]/NET0131  & ~n11444 ;
  assign n11446 = \rf_conf6_reg[13]/NET0131  & ~\s6_msel_arb3_state_reg[0]/NET0131  ;
  assign n11447 = n4678 & n11446 ;
  assign n11448 = \s6_msel_arb3_state_reg[2]/NET0131  & ~n4690 ;
  assign n11449 = ~n4668 & n4685 ;
  assign n11450 = ~n11448 & ~n11449 ;
  assign n11451 = ~n11447 & ~n11450 ;
  assign n11452 = ~n4690 & ~n4698 ;
  assign n11453 = ~n4684 & n8638 ;
  assign n11454 = ~n11452 & ~n11453 ;
  assign n11455 = ~n4679 & ~n4682 ;
  assign n11456 = ~n11454 & n11455 ;
  assign n11457 = ~n11451 & ~n11456 ;
  assign n11458 = ~n4677 & ~n11457 ;
  assign n11459 = ~n4668 & ~n4682 ;
  assign n11460 = n4699 & n11459 ;
  assign n11461 = \s6_msel_arb3_state_reg[1]/NET0131  & ~n11460 ;
  assign n11462 = ~n11458 & n11461 ;
  assign n11463 = ~n11445 & ~n11462 ;
  assign n11464 = ~\s7_msel_arb2_state_reg[2]/NET0131  & ~n9974 ;
  assign n11465 = ~n9956 & n9963 ;
  assign n11466 = ~\s7_msel_arb2_state_reg[0]/NET0131  & n11465 ;
  assign n11467 = ~n9979 & ~n11466 ;
  assign n11468 = ~n11464 & ~n11467 ;
  assign n11469 = ~\s7_msel_arb2_state_reg[1]/NET0131  & n9963 ;
  assign n11470 = n9974 & n11469 ;
  assign n11471 = ~n11468 & ~n11470 ;
  assign n11472 = \s7_msel_arb2_state_reg[2]/NET0131  & ~n9963 ;
  assign n11473 = ~n9964 & n9974 ;
  assign n11474 = ~\s7_msel_arb2_state_reg[0]/NET0131  & n11473 ;
  assign n11475 = ~n9985 & ~n11474 ;
  assign n11476 = ~n11472 & ~n11475 ;
  assign n11477 = n8811 & n8834 ;
  assign n11478 = n8834 & n9956 ;
  assign n11479 = ~n11473 & n11478 ;
  assign n11480 = ~n11477 & ~n11479 ;
  assign n11481 = \s7_msel_arb2_state_reg[0]/NET0131  & n11480 ;
  assign n11482 = ~n11476 & ~n11481 ;
  assign n11483 = n11471 & n11482 ;
  assign n11484 = n8857 & ~n9963 ;
  assign n11485 = \s7_msel_arb2_state_reg[1]/NET0131  & ~n8820 ;
  assign n11486 = n9974 & ~n11485 ;
  assign n11487 = n8857 & n9956 ;
  assign n11488 = ~n11486 & n11487 ;
  assign n11489 = ~n11484 & ~n11488 ;
  assign n11490 = \s7_msel_arb2_state_reg[1]/NET0131  & n8806 ;
  assign n11491 = \s7_msel_arb2_state_reg[1]/NET0131  & n9964 ;
  assign n11492 = ~n11465 & n11491 ;
  assign n11493 = ~n11490 & ~n11492 ;
  assign n11494 = ~n9963 & n9964 ;
  assign n11495 = n9974 & ~n11494 ;
  assign n11496 = ~\s7_msel_arb2_state_reg[1]/NET0131  & ~n8815 ;
  assign n11497 = ~n11495 & n11496 ;
  assign n11498 = n11493 & ~n11497 ;
  assign n11499 = \s7_msel_arb2_state_reg[0]/NET0131  & ~\s7_msel_arb2_state_reg[2]/NET0131  ;
  assign n11500 = ~n11498 & n11499 ;
  assign n11501 = n11489 & ~n11500 ;
  assign n11502 = ~n11483 & n11501 ;
  assign n11503 = ~n4741 & ~n8911 ;
  assign n11504 = ~\s7_msel_arb3_state_reg[2]/NET0131  & ~n11503 ;
  assign n11505 = ~n4724 & ~n11504 ;
  assign n11506 = n4722 & ~n4734 ;
  assign n11507 = n11505 & n11506 ;
  assign n11508 = \s7_msel_arb3_state_reg[2]/NET0131  & ~n4723 ;
  assign n11509 = ~n4739 & n11503 ;
  assign n11510 = ~n11508 & n11509 ;
  assign n11511 = ~n4719 & n4724 ;
  assign n11512 = ~n4739 & n4744 ;
  assign n11513 = n4734 & ~n11512 ;
  assign n11514 = n11511 & ~n11513 ;
  assign n11515 = ~n11510 & ~n11514 ;
  assign n11516 = ~n11507 & n11515 ;
  assign n11517 = ~\s7_msel_arb3_state_reg[1]/NET0131  & ~n11516 ;
  assign n11518 = \rf_conf7_reg[13]/NET0131  & ~\s7_msel_arb3_state_reg[0]/NET0131  ;
  assign n11519 = n4732 & n11518 ;
  assign n11520 = \s7_msel_arb3_state_reg[2]/NET0131  & ~n4744 ;
  assign n11521 = ~n4722 & n4739 ;
  assign n11522 = ~n11520 & ~n11521 ;
  assign n11523 = ~n11519 & ~n11522 ;
  assign n11524 = ~n4744 & ~n4752 ;
  assign n11525 = ~n4738 & n8924 ;
  assign n11526 = ~n11524 & ~n11525 ;
  assign n11527 = ~n4733 & ~n4736 ;
  assign n11528 = ~n11526 & n11527 ;
  assign n11529 = ~n11523 & ~n11528 ;
  assign n11530 = ~n4731 & ~n11529 ;
  assign n11531 = ~n4722 & ~n4736 ;
  assign n11532 = n4753 & n11531 ;
  assign n11533 = \s7_msel_arb3_state_reg[1]/NET0131  & ~n11532 ;
  assign n11534 = ~n11530 & n11533 ;
  assign n11535 = ~n11517 & ~n11534 ;
  assign n11536 = \rf_conf8_reg[5]/NET0131  & ~\s8_msel_arb2_state_reg[0]/NET0131  ;
  assign n11537 = n3330 & n11536 ;
  assign n11538 = n4125 & ~n11537 ;
  assign n11539 = \rf_conf8_reg[7]/NET0131  & \s8_msel_arb2_state_reg[0]/NET0131  ;
  assign n11540 = n3324 & n11539 ;
  assign n11541 = ~\s8_msel_arb2_state_reg[2]/NET0131  & ~n11540 ;
  assign n11542 = ~n11538 & n11541 ;
  assign n11543 = ~\s8_msel_arb2_state_reg[1]/NET0131  & ~n4133 ;
  assign n11544 = n4145 & ~n11543 ;
  assign n11545 = n4128 & n11541 ;
  assign n11546 = ~n11544 & n11545 ;
  assign n11547 = ~n11542 & ~n11546 ;
  assign n11548 = \s8_msel_arb2_state_reg[2]/NET0131  & ~n9111 ;
  assign n11549 = ~n4127 & n11548 ;
  assign n11550 = \s8_msel_arb2_state_reg[1]/NET0131  & ~n11549 ;
  assign n11551 = ~n4125 & n4143 ;
  assign n11552 = \s8_msel_arb2_state_reg[1]/NET0131  & n4145 ;
  assign n11553 = ~n11551 & n11552 ;
  assign n11554 = ~n11550 & ~n11553 ;
  assign n11555 = n11547 & ~n11554 ;
  assign n11556 = ~n4143 & n4145 ;
  assign n11557 = n4128 & ~n11556 ;
  assign n11558 = ~n4123 & n9123 ;
  assign n11559 = ~\s8_msel_arb2_state_reg[2]/NET0131  & ~n4145 ;
  assign n11560 = ~\s8_msel_arb2_state_reg[0]/NET0131  & ~\s8_msel_arb2_state_reg[1]/NET0131  ;
  assign n11561 = n4125 & n11560 ;
  assign n11562 = ~n11559 & n11561 ;
  assign n11563 = ~n11558 & ~n11562 ;
  assign n11564 = ~n11557 & ~n11563 ;
  assign n11565 = ~\s8_msel_arb2_state_reg[1]/NET0131  & ~n4145 ;
  assign n11566 = ~\s8_msel_arb2_state_reg[0]/NET0131  & ~n4143 ;
  assign n11567 = ~n11565 & n11566 ;
  assign n11568 = ~\s8_msel_arb2_state_reg[2]/NET0131  & n11567 ;
  assign n11569 = n4125 & ~n4128 ;
  assign n11570 = n4143 & ~n11569 ;
  assign n11571 = ~n4138 & n9122 ;
  assign n11572 = ~\s8_msel_arb2_state_reg[2]/NET0131  & n11571 ;
  assign n11573 = ~n11570 & n11572 ;
  assign n11574 = ~n11568 & ~n11573 ;
  assign n11575 = ~n11564 & n11574 ;
  assign n11576 = ~n11555 & n11575 ;
  assign n11577 = n4777 & ~n4782 ;
  assign n11578 = ~n4785 & n11577 ;
  assign n11579 = ~n4774 & ~n4798 ;
  assign n11580 = ~\s8_msel_arb3_state_reg[2]/NET0131  & ~n11579 ;
  assign n11581 = ~n4785 & ~n4790 ;
  assign n11582 = ~n11580 & n11581 ;
  assign n11583 = ~n11578 & ~n11582 ;
  assign n11584 = ~n4782 & n4802 ;
  assign n11585 = n11583 & ~n11584 ;
  assign n11586 = ~\s8_msel_arb3_state_reg[1]/NET0131  & ~n11585 ;
  assign n11587 = \s8_msel_arb3_state_reg[2]/NET0131  & ~n4777 ;
  assign n11588 = ~n4787 & n11587 ;
  assign n11589 = ~n4777 & ~n4789 ;
  assign n11590 = ~n4781 & ~n4799 ;
  assign n11591 = ~n11589 & ~n11590 ;
  assign n11592 = ~n4779 & ~n4787 ;
  assign n11593 = ~n11591 & n11592 ;
  assign n11594 = ~n11588 & ~n11593 ;
  assign n11595 = ~\s8_msel_arb3_state_reg[2]/NET0131  & ~n4779 ;
  assign n11596 = ~n4799 & n11595 ;
  assign n11597 = \s8_msel_arb3_state_reg[1]/NET0131  & ~n11596 ;
  assign n11598 = n11594 & n11597 ;
  assign n11599 = ~n11586 & ~n11598 ;
  assign n11600 = \s8_msel_arb3_state_reg[0]/NET0131  & ~n11599 ;
  assign n11601 = ~\s8_msel_arb3_state_reg[1]/NET0131  & ~n4799 ;
  assign n11602 = ~n4777 & n4790 ;
  assign n11603 = ~n11601 & ~n11602 ;
  assign n11604 = \s8_msel_arb3_state_reg[2]/NET0131  & ~n11603 ;
  assign n11605 = ~\s8_msel_arb3_state_reg[0]/NET0131  & ~n11604 ;
  assign n11606 = n4782 & ~n4799 ;
  assign n11607 = ~n4811 & ~n11606 ;
  assign n11608 = ~\s8_msel_arb3_state_reg[2]/NET0131  & ~n11607 ;
  assign n11609 = \s8_msel_arb3_state_reg[1]/NET0131  & n4777 ;
  assign n11610 = n4799 & n11609 ;
  assign n11611 = n4782 & n4790 ;
  assign n11612 = ~n11610 & n11611 ;
  assign n11613 = ~n11608 & ~n11612 ;
  assign n11614 = n11605 & n11613 ;
  assign n11615 = ~n11600 & ~n11614 ;
  assign n11616 = ~\s9_msel_arb2_state_reg[2]/NET0131  & ~n10009 ;
  assign n11617 = ~n9991 & n9998 ;
  assign n11618 = ~\s9_msel_arb2_state_reg[0]/NET0131  & n11617 ;
  assign n11619 = ~n10014 & ~n11618 ;
  assign n11620 = ~n11616 & ~n11619 ;
  assign n11621 = ~\s9_msel_arb2_state_reg[1]/NET0131  & n9998 ;
  assign n11622 = n10009 & n11621 ;
  assign n11623 = ~n11620 & ~n11622 ;
  assign n11624 = \s9_msel_arb2_state_reg[2]/NET0131  & ~n9998 ;
  assign n11625 = ~n9999 & n10009 ;
  assign n11626 = ~\s9_msel_arb2_state_reg[0]/NET0131  & n11625 ;
  assign n11627 = ~n10020 & ~n11626 ;
  assign n11628 = ~n11624 & ~n11627 ;
  assign n11629 = n9336 & n9359 ;
  assign n11630 = n9359 & n9991 ;
  assign n11631 = ~n11625 & n11630 ;
  assign n11632 = ~n11629 & ~n11631 ;
  assign n11633 = \s9_msel_arb2_state_reg[0]/NET0131  & n11632 ;
  assign n11634 = ~n11628 & ~n11633 ;
  assign n11635 = n11623 & n11634 ;
  assign n11636 = n9382 & ~n9998 ;
  assign n11637 = \s9_msel_arb2_state_reg[1]/NET0131  & ~n9345 ;
  assign n11638 = n10009 & ~n11637 ;
  assign n11639 = n9382 & n9991 ;
  assign n11640 = ~n11638 & n11639 ;
  assign n11641 = ~n11636 & ~n11640 ;
  assign n11642 = \s9_msel_arb2_state_reg[1]/NET0131  & n9331 ;
  assign n11643 = \s9_msel_arb2_state_reg[1]/NET0131  & n9999 ;
  assign n11644 = ~n11617 & n11643 ;
  assign n11645 = ~n11642 & ~n11644 ;
  assign n11646 = ~n9998 & n9999 ;
  assign n11647 = n10009 & ~n11646 ;
  assign n11648 = ~\s9_msel_arb2_state_reg[1]/NET0131  & ~n9340 ;
  assign n11649 = ~n11647 & n11648 ;
  assign n11650 = n11645 & ~n11649 ;
  assign n11651 = \s9_msel_arb2_state_reg[0]/NET0131  & ~\s9_msel_arb2_state_reg[2]/NET0131  ;
  assign n11652 = ~n11650 & n11651 ;
  assign n11653 = n11641 & ~n11652 ;
  assign n11654 = ~n11635 & n11653 ;
  assign n11655 = n10027 & ~n10044 ;
  assign n11656 = \s9_msel_arb3_state_reg[1]/NET0131  & ~n11655 ;
  assign n11657 = ~\s9_msel_arb3_state_reg[1]/NET0131  & ~n10044 ;
  assign n11658 = \s9_msel_arb3_state_reg[2]/NET0131  & ~n11657 ;
  assign n11659 = ~n11656 & ~n11658 ;
  assign n11660 = ~\s9_msel_arb3_state_reg[0]/NET0131  & n11659 ;
  assign n11661 = \s9_msel_arb3_state_reg[1]/NET0131  & n10044 ;
  assign n11662 = n10027 & ~n11661 ;
  assign n11663 = n10026 & ~n11662 ;
  assign n11664 = ~\s9_msel_arb3_state_reg[2]/NET0131  & ~n10027 ;
  assign n11665 = n10043 & ~n11664 ;
  assign n11666 = ~\s9_msel_arb3_state_reg[0]/NET0131  & n11665 ;
  assign n11667 = ~n11663 & n11666 ;
  assign n11668 = ~n11660 & ~n11667 ;
  assign n11669 = ~n9413 & n11655 ;
  assign n11670 = ~n9416 & ~n9425 ;
  assign n11671 = ~\s9_msel_arb3_state_reg[2]/NET0131  & ~n11670 ;
  assign n11672 = ~n9413 & ~n10026 ;
  assign n11673 = ~n11671 & n11672 ;
  assign n11674 = ~n11669 & ~n11673 ;
  assign n11675 = n10039 & ~n10044 ;
  assign n11676 = \s9_msel_arb3_state_reg[1]/NET0131  & ~n11675 ;
  assign n11677 = n11674 & n11676 ;
  assign n11678 = ~n9423 & n9437 ;
  assign n11679 = \s9_msel_arb3_state_reg[0]/NET0131  & ~n11678 ;
  assign n11680 = n10026 & ~n10027 ;
  assign n11681 = \s9_msel_arb3_state_reg[0]/NET0131  & n10043 ;
  assign n11682 = ~n11680 & n11681 ;
  assign n11683 = ~n11679 & ~n11682 ;
  assign n11684 = ~n11677 & ~n11683 ;
  assign n11685 = n11668 & ~n11684 ;
  assign n11686 = ~n10043 & n10044 ;
  assign n11687 = n10027 & ~n11686 ;
  assign n11688 = \rf_conf9_reg[1]/NET0131  & ~\s9_msel_arb3_state_reg[0]/NET0131  ;
  assign n11689 = n5398 & n11688 ;
  assign n11690 = n9472 & ~n11689 ;
  assign n11691 = ~n11687 & n11690 ;
  assign n11692 = ~n11685 & ~n11691 ;
  assign n11693 = \rf_conf0_reg[5]/NET0131  & ~\s0_msel_arb2_state_reg[0]/NET0131  ;
  assign n11694 = n3623 & n11693 ;
  assign n11695 = n4160 & ~n11694 ;
  assign n11696 = \rf_conf0_reg[7]/NET0131  & \s0_msel_arb2_state_reg[0]/NET0131  ;
  assign n11697 = n3621 & n11696 ;
  assign n11698 = ~\s0_msel_arb2_state_reg[2]/NET0131  & ~n11697 ;
  assign n11699 = ~n11695 & n11698 ;
  assign n11700 = ~\s0_msel_arb2_state_reg[1]/NET0131  & ~n4168 ;
  assign n11701 = n4180 & ~n11700 ;
  assign n11702 = n4163 & n11698 ;
  assign n11703 = ~n11701 & n11702 ;
  assign n11704 = ~n11699 & ~n11703 ;
  assign n11705 = \s0_msel_arb2_state_reg[2]/NET0131  & ~n9642 ;
  assign n11706 = ~n4162 & n11705 ;
  assign n11707 = \s0_msel_arb2_state_reg[1]/NET0131  & ~n11706 ;
  assign n11708 = ~n4160 & n4178 ;
  assign n11709 = \s0_msel_arb2_state_reg[1]/NET0131  & n4180 ;
  assign n11710 = ~n11708 & n11709 ;
  assign n11711 = ~n11707 & ~n11710 ;
  assign n11712 = n11704 & ~n11711 ;
  assign n11713 = ~n4178 & n4180 ;
  assign n11714 = n4163 & ~n11713 ;
  assign n11715 = ~n4158 & n9654 ;
  assign n11716 = ~\s0_msel_arb2_state_reg[2]/NET0131  & ~n4180 ;
  assign n11717 = ~\s0_msel_arb2_state_reg[0]/NET0131  & ~\s0_msel_arb2_state_reg[1]/NET0131  ;
  assign n11718 = n4160 & n11717 ;
  assign n11719 = ~n11716 & n11718 ;
  assign n11720 = ~n11715 & ~n11719 ;
  assign n11721 = ~n11714 & ~n11720 ;
  assign n11722 = ~\s0_msel_arb2_state_reg[1]/NET0131  & ~n4180 ;
  assign n11723 = ~\s0_msel_arb2_state_reg[0]/NET0131  & ~n4178 ;
  assign n11724 = ~n11722 & n11723 ;
  assign n11725 = ~\s0_msel_arb2_state_reg[2]/NET0131  & n11724 ;
  assign n11726 = n4160 & ~n4163 ;
  assign n11727 = n4178 & ~n11726 ;
  assign n11728 = ~n4173 & n9653 ;
  assign n11729 = ~\s0_msel_arb2_state_reg[2]/NET0131  & n11728 ;
  assign n11730 = ~n11727 & n11729 ;
  assign n11731 = ~n11725 & ~n11730 ;
  assign n11732 = ~n11721 & n11731 ;
  assign n11733 = ~n11712 & n11732 ;
  assign n11734 = ~n4846 & ~n9696 ;
  assign n11735 = ~\s0_msel_arb3_state_reg[2]/NET0131  & ~n11734 ;
  assign n11736 = ~n4829 & ~n11735 ;
  assign n11737 = n4827 & ~n4839 ;
  assign n11738 = n11736 & n11737 ;
  assign n11739 = \s0_msel_arb3_state_reg[2]/NET0131  & ~n4828 ;
  assign n11740 = ~n4844 & n11734 ;
  assign n11741 = ~n11739 & n11740 ;
  assign n11742 = ~n4824 & n4829 ;
  assign n11743 = ~n4844 & n4849 ;
  assign n11744 = n4839 & ~n11743 ;
  assign n11745 = n11742 & ~n11744 ;
  assign n11746 = ~n11741 & ~n11745 ;
  assign n11747 = ~n11738 & n11746 ;
  assign n11748 = ~\s0_msel_arb3_state_reg[1]/NET0131  & ~n11747 ;
  assign n11749 = \rf_conf0_reg[13]/NET0131  & ~\s0_msel_arb3_state_reg[0]/NET0131  ;
  assign n11750 = n4837 & n11749 ;
  assign n11751 = \s0_msel_arb3_state_reg[2]/NET0131  & ~n4849 ;
  assign n11752 = ~n4827 & n4844 ;
  assign n11753 = ~n11751 & ~n11752 ;
  assign n11754 = ~n11750 & ~n11753 ;
  assign n11755 = ~n4849 & ~n4857 ;
  assign n11756 = ~n4843 & n9709 ;
  assign n11757 = ~n11755 & ~n11756 ;
  assign n11758 = ~n4838 & ~n4841 ;
  assign n11759 = ~n11757 & n11758 ;
  assign n11760 = ~n11754 & ~n11759 ;
  assign n11761 = ~n4836 & ~n11760 ;
  assign n11762 = ~n4827 & ~n4841 ;
  assign n11763 = n4858 & n11762 ;
  assign n11764 = \s0_msel_arb3_state_reg[1]/NET0131  & ~n11763 ;
  assign n11765 = ~n11761 & n11764 ;
  assign n11766 = ~n11748 & ~n11765 ;
  assign n11767 = ~n4885 & n4888 ;
  assign n11768 = n4903 & ~n11767 ;
  assign n11769 = \s10_msel_arb1_state_reg[2]/NET0131  & n4902 ;
  assign n11770 = ~n11768 & n11769 ;
  assign n11771 = ~\s10_msel_arb1_state_reg[0]/NET0131  & n11770 ;
  assign n11772 = ~n4888 & n4903 ;
  assign n11773 = n4902 & ~n11772 ;
  assign n11774 = ~\s10_msel_arb1_state_reg[2]/NET0131  & ~n4885 ;
  assign n11775 = ~n11767 & ~n11774 ;
  assign n11776 = ~n11773 & n11775 ;
  assign n11777 = ~\s10_msel_arb1_state_reg[0]/NET0131  & \s10_msel_arb1_state_reg[1]/NET0131  ;
  assign n11778 = ~n11776 & n11777 ;
  assign n11779 = ~n11771 & ~n11778 ;
  assign n11780 = n4885 & ~n4902 ;
  assign n11781 = \s10_msel_arb1_state_reg[0]/NET0131  & n4888 ;
  assign n11782 = ~n11780 & n11781 ;
  assign n11783 = \s10_msel_arb1_state_reg[2]/NET0131  & ~n4890 ;
  assign n11784 = ~n5540 & n11783 ;
  assign n11785 = ~n11782 & n11784 ;
  assign n11786 = \s10_msel_arb1_state_reg[1]/NET0131  & n4902 ;
  assign n11787 = ~n11772 & n11786 ;
  assign n11788 = ~\rf_conf10_reg[7]/NET0131  & \s10_msel_arb1_state_reg[0]/NET0131  ;
  assign n11789 = n4210 & n11788 ;
  assign n11790 = ~\s10_msel_arb1_state_reg[2]/NET0131  & ~n11789 ;
  assign n11791 = \s10_msel_arb1_state_reg[1]/NET0131  & ~n11790 ;
  assign n11792 = ~n11787 & ~n11791 ;
  assign n11793 = ~n11785 & ~n11792 ;
  assign n11794 = n4902 & ~n4903 ;
  assign n11795 = n4885 & ~n11794 ;
  assign n11796 = n4900 & n5521 ;
  assign n11797 = ~n11795 & n11796 ;
  assign n11798 = \s10_msel_arb1_state_reg[0]/NET0131  & n5512 ;
  assign n11799 = ~n4877 & n11798 ;
  assign n11800 = ~n11768 & n11799 ;
  assign n11801 = ~n11797 & ~n11800 ;
  assign n11802 = ~n11793 & n11801 ;
  assign n11803 = n11779 & n11802 ;
  assign n11804 = ~n4916 & n4919 ;
  assign n11805 = n4939 & ~n11804 ;
  assign n11806 = ~\s11_msel_arb1_state_reg[1]/NET0131  & ~n4934 ;
  assign n11807 = ~n4928 & n11806 ;
  assign n11808 = ~n11805 & n11807 ;
  assign n11809 = ~\s11_msel_arb1_state_reg[2]/NET0131  & n11808 ;
  assign n11810 = n4916 & ~n4943 ;
  assign n11811 = \s11_msel_arb1_state_reg[0]/NET0131  & n4919 ;
  assign n11812 = ~n11810 & n11811 ;
  assign n11813 = ~\rf_conf11_reg[5]/NET0131  & ~\s11_msel_arb1_state_reg[0]/NET0131  ;
  assign n11814 = n4290 & n11813 ;
  assign n11815 = ~n4911 & ~n11814 ;
  assign n11816 = ~n11812 & n11815 ;
  assign n11817 = n4912 & ~n11816 ;
  assign n11818 = ~n11809 & ~n11817 ;
  assign n11819 = n5807 & ~n11810 ;
  assign n11820 = ~n4918 & n11819 ;
  assign n11821 = ~n4939 & n4943 ;
  assign n11822 = n4916 & ~n11821 ;
  assign n11823 = ~n4918 & n5786 ;
  assign n11824 = ~n11822 & n11823 ;
  assign n11825 = ~n11820 & ~n11824 ;
  assign n11826 = n4924 & ~n4952 ;
  assign n11827 = ~n4919 & n4939 ;
  assign n11828 = n4924 & n4943 ;
  assign n11829 = ~n11827 & n11828 ;
  assign n11830 = ~n11826 & ~n11829 ;
  assign n11831 = n11825 & n11830 ;
  assign n11832 = n11818 & n11831 ;
  assign n11833 = ~n4970 & n4973 ;
  assign n11834 = n4994 & ~n11833 ;
  assign n11835 = ~\s12_msel_arb1_state_reg[1]/NET0131  & n4966 ;
  assign n11836 = ~n11834 & n11835 ;
  assign n11837 = ~\s12_msel_arb1_state_reg[0]/NET0131  & \s12_msel_arb1_state_reg[1]/NET0131  ;
  assign n11838 = ~n4994 & n11837 ;
  assign n11839 = n4970 & ~n4993 ;
  assign n11840 = n4973 & n11837 ;
  assign n11841 = ~n11839 & n11840 ;
  assign n11842 = ~n11838 & ~n11841 ;
  assign n11843 = ~n11836 & n11842 ;
  assign n11844 = ~\s12_msel_arb1_state_reg[2]/NET0131  & ~n11843 ;
  assign n11845 = ~n4973 & n4994 ;
  assign n11846 = n4993 & ~n11845 ;
  assign n11847 = n4970 & ~n11846 ;
  assign n11848 = \s12_msel_arb1_state_reg[2]/NET0131  & ~n4975 ;
  assign n11849 = \s12_msel_arb1_state_reg[1]/NET0131  & n11848 ;
  assign n11850 = n4970 & n4994 ;
  assign n11851 = n4988 & n11848 ;
  assign n11852 = ~n11850 & n11851 ;
  assign n11853 = ~n11849 & ~n11852 ;
  assign n11854 = ~n11847 & ~n11853 ;
  assign n11855 = ~n4978 & n11839 ;
  assign n11856 = ~n4968 & ~n4976 ;
  assign n11857 = \s12_msel_arb1_state_reg[2]/NET0131  & ~n11856 ;
  assign n11858 = ~n4973 & ~n4978 ;
  assign n11859 = ~n11857 & n11858 ;
  assign n11860 = ~n11855 & ~n11859 ;
  assign n11861 = n4991 & ~n4993 ;
  assign n11862 = n4975 & ~n11861 ;
  assign n11863 = n11860 & n11862 ;
  assign n11864 = ~n11854 & ~n11863 ;
  assign n11865 = ~n11844 & n11864 ;
  assign n11866 = ~n5007 & n5010 ;
  assign n11867 = n5025 & ~n11866 ;
  assign n11868 = \s13_msel_arb1_state_reg[2]/NET0131  & n5024 ;
  assign n11869 = ~n11867 & n11868 ;
  assign n11870 = ~\s13_msel_arb1_state_reg[0]/NET0131  & n11869 ;
  assign n11871 = ~n5010 & n5025 ;
  assign n11872 = n5024 & ~n11871 ;
  assign n11873 = ~\s13_msel_arb1_state_reg[2]/NET0131  & ~n5007 ;
  assign n11874 = ~n11866 & ~n11873 ;
  assign n11875 = ~n11872 & n11874 ;
  assign n11876 = ~\s13_msel_arb1_state_reg[0]/NET0131  & \s13_msel_arb1_state_reg[1]/NET0131  ;
  assign n11877 = ~n11875 & n11876 ;
  assign n11878 = ~n11870 & ~n11877 ;
  assign n11879 = n5007 & ~n5024 ;
  assign n11880 = \s13_msel_arb1_state_reg[0]/NET0131  & n5010 ;
  assign n11881 = ~n11879 & n11880 ;
  assign n11882 = \s13_msel_arb1_state_reg[2]/NET0131  & ~n5012 ;
  assign n11883 = ~n6372 & n11882 ;
  assign n11884 = ~n11881 & n11883 ;
  assign n11885 = \s13_msel_arb1_state_reg[1]/NET0131  & n5024 ;
  assign n11886 = ~n11871 & n11885 ;
  assign n11887 = ~\rf_conf13_reg[7]/NET0131  & \s13_msel_arb1_state_reg[0]/NET0131  ;
  assign n11888 = n3865 & n11887 ;
  assign n11889 = ~\s13_msel_arb1_state_reg[2]/NET0131  & ~n11888 ;
  assign n11890 = \s13_msel_arb1_state_reg[1]/NET0131  & ~n11889 ;
  assign n11891 = ~n11886 & ~n11890 ;
  assign n11892 = ~n11884 & ~n11891 ;
  assign n11893 = n5024 & ~n5025 ;
  assign n11894 = n5007 & ~n11893 ;
  assign n11895 = n5022 & n6353 ;
  assign n11896 = ~n11894 & n11895 ;
  assign n11897 = \s13_msel_arb1_state_reg[0]/NET0131  & n6344 ;
  assign n11898 = ~n4999 & n11897 ;
  assign n11899 = ~n11867 & n11898 ;
  assign n11900 = ~n11896 & ~n11899 ;
  assign n11901 = ~n11892 & n11900 ;
  assign n11902 = n11878 & n11901 ;
  assign n11903 = n5038 & n5059 ;
  assign n11904 = ~n6649 & ~n11903 ;
  assign n11905 = \s14_msel_arb1_state_reg[1]/NET0131  & ~n11904 ;
  assign n11906 = ~\s14_msel_arb1_state_reg[0]/NET0131  & n5033 ;
  assign n11907 = n5038 & n11906 ;
  assign n11908 = ~\s14_msel_arb1_state_reg[0]/NET0131  & n5038 ;
  assign n11909 = ~\s14_msel_arb1_state_reg[1]/NET0131  & ~n11908 ;
  assign n11910 = n5059 & ~n5060 ;
  assign n11911 = ~n5034 & ~n11910 ;
  assign n11912 = ~n11909 & ~n11911 ;
  assign n11913 = ~n11907 & ~n11912 ;
  assign n11914 = ~n11905 & n11913 ;
  assign n11915 = \s14_msel_arb1_state_reg[2]/NET0131  & ~n11914 ;
  assign n11916 = ~n5058 & n6625 ;
  assign n11917 = n5038 & n11916 ;
  assign n11918 = ~n5048 & n11917 ;
  assign n11919 = ~n5035 & n5038 ;
  assign n11920 = n5060 & ~n11919 ;
  assign n11921 = ~n5046 & n6620 ;
  assign n11922 = ~n5048 & n11921 ;
  assign n11923 = ~n11920 & n11922 ;
  assign n11924 = ~n11918 & ~n11923 ;
  assign n11925 = ~n5042 & ~n5052 ;
  assign n11926 = ~n11919 & n11925 ;
  assign n11927 = n6625 & ~n11926 ;
  assign n11928 = n5035 & ~n11910 ;
  assign n11929 = ~n5037 & n6660 ;
  assign n11930 = ~n11928 & n11929 ;
  assign n11931 = ~n11927 & ~n11930 ;
  assign n11932 = n11924 & n11931 ;
  assign n11933 = ~n11915 & n11932 ;
  assign n11934 = n3751 & ~n3767 ;
  assign n11935 = n3756 & ~n11934 ;
  assign n11936 = n3842 & ~n11935 ;
  assign n11937 = ~\s15_msel_arb1_state_reg[2]/NET0131  & ~n3748 ;
  assign n11938 = \s15_msel_arb1_state_reg[1]/NET0131  & ~n11937 ;
  assign n11939 = ~n3756 & n3762 ;
  assign n11940 = \s15_msel_arb1_state_reg[1]/NET0131  & n3767 ;
  assign n11941 = ~n11939 & n11940 ;
  assign n11942 = ~n11938 & ~n11941 ;
  assign n11943 = ~n11936 & ~n11942 ;
  assign n11944 = \s15_msel_arb1_state_reg[0]/NET0131  & n11943 ;
  assign n11945 = \s15_msel_arb1_state_reg[2]/NET0131  & n3764 ;
  assign n11946 = ~n3751 & n3756 ;
  assign n11947 = \s15_msel_arb1_state_reg[2]/NET0131  & n3762 ;
  assign n11948 = ~n11946 & n11947 ;
  assign n11949 = ~n11945 & ~n11948 ;
  assign n11950 = ~\s15_msel_arb1_state_reg[1]/NET0131  & n11949 ;
  assign n11951 = ~\s15_msel_arb1_state_reg[2]/NET0131  & n3755 ;
  assign n11952 = ~n3762 & n3767 ;
  assign n11953 = ~\s15_msel_arb1_state_reg[2]/NET0131  & n3751 ;
  assign n11954 = ~n11952 & n11953 ;
  assign n11955 = ~n11951 & ~n11954 ;
  assign n11956 = \s15_msel_arb1_state_reg[0]/NET0131  & n11955 ;
  assign n11957 = n11950 & n11956 ;
  assign n11958 = ~n11944 & ~n11957 ;
  assign n11959 = ~\s15_msel_arb1_state_reg[1]/NET0131  & ~n3756 ;
  assign n11960 = ~n11934 & ~n11959 ;
  assign n11961 = ~\s15_msel_arb1_state_reg[2]/NET0131  & ~n11960 ;
  assign n11962 = ~\s15_msel_arb1_state_reg[0]/NET0131  & ~n11961 ;
  assign n11963 = \s15_msel_arb1_state_reg[2]/NET0131  & n11939 ;
  assign n11964 = ~\s15_msel_arb1_state_reg[1]/NET0131  & \s15_msel_arb1_state_reg[2]/NET0131  ;
  assign n11965 = ~n3767 & n11964 ;
  assign n11966 = ~n11963 & ~n11965 ;
  assign n11967 = \s15_msel_arb1_state_reg[1]/NET0131  & n3756 ;
  assign n11968 = n3767 & n11967 ;
  assign n11969 = n3751 & n3762 ;
  assign n11970 = ~n11968 & n11969 ;
  assign n11971 = n11966 & ~n11970 ;
  assign n11972 = n11962 & n11971 ;
  assign n11973 = n11958 & ~n11972 ;
  assign n11974 = n5077 & n5098 ;
  assign n11975 = ~n7131 & ~n11974 ;
  assign n11976 = \s1_msel_arb1_state_reg[1]/NET0131  & ~n11975 ;
  assign n11977 = ~\s1_msel_arb1_state_reg[0]/NET0131  & n5072 ;
  assign n11978 = n5077 & n11977 ;
  assign n11979 = ~\s1_msel_arb1_state_reg[0]/NET0131  & n5077 ;
  assign n11980 = ~\s1_msel_arb1_state_reg[1]/NET0131  & ~n11979 ;
  assign n11981 = n5098 & ~n5099 ;
  assign n11982 = ~n5073 & ~n11981 ;
  assign n11983 = ~n11980 & ~n11982 ;
  assign n11984 = ~n11978 & ~n11983 ;
  assign n11985 = ~n11976 & n11984 ;
  assign n11986 = \s1_msel_arb1_state_reg[2]/NET0131  & ~n11985 ;
  assign n11987 = ~n5097 & n7107 ;
  assign n11988 = n5077 & n11987 ;
  assign n11989 = ~n5087 & n11988 ;
  assign n11990 = ~n5074 & n5077 ;
  assign n11991 = n5099 & ~n11990 ;
  assign n11992 = ~n5085 & n7102 ;
  assign n11993 = ~n5087 & n11992 ;
  assign n11994 = ~n11991 & n11993 ;
  assign n11995 = ~n11989 & ~n11994 ;
  assign n11996 = ~n5081 & ~n5091 ;
  assign n11997 = ~n11990 & n11996 ;
  assign n11998 = n7107 & ~n11997 ;
  assign n11999 = n5074 & ~n11981 ;
  assign n12000 = ~n5076 & n7142 ;
  assign n12001 = ~n11999 & n12000 ;
  assign n12002 = ~n11998 & ~n12001 ;
  assign n12003 = n11995 & n12002 ;
  assign n12004 = ~n11986 & n12003 ;
  assign n12005 = ~n5119 & n5122 ;
  assign n12006 = n5137 & ~n12005 ;
  assign n12007 = \s2_msel_arb1_state_reg[2]/NET0131  & n5136 ;
  assign n12008 = ~n12006 & n12007 ;
  assign n12009 = ~\s2_msel_arb1_state_reg[0]/NET0131  & n12008 ;
  assign n12010 = ~n5122 & n5137 ;
  assign n12011 = n5136 & ~n12010 ;
  assign n12012 = ~\s2_msel_arb1_state_reg[2]/NET0131  & ~n5119 ;
  assign n12013 = ~n12005 & ~n12012 ;
  assign n12014 = ~n12011 & n12013 ;
  assign n12015 = ~\s2_msel_arb1_state_reg[0]/NET0131  & \s2_msel_arb1_state_reg[1]/NET0131  ;
  assign n12016 = ~n12014 & n12015 ;
  assign n12017 = ~n12009 & ~n12016 ;
  assign n12018 = n5119 & ~n5136 ;
  assign n12019 = \s2_msel_arb1_state_reg[0]/NET0131  & n5122 ;
  assign n12020 = ~n12018 & n12019 ;
  assign n12021 = \s2_msel_arb1_state_reg[2]/NET0131  & ~n5124 ;
  assign n12022 = ~n7417 & n12021 ;
  assign n12023 = ~n12020 & n12022 ;
  assign n12024 = \s2_msel_arb1_state_reg[1]/NET0131  & n5136 ;
  assign n12025 = ~n12010 & n12024 ;
  assign n12026 = ~\rf_conf2_reg[7]/NET0131  & \s2_msel_arb1_state_reg[0]/NET0131  ;
  assign n12027 = n3965 & n12026 ;
  assign n12028 = ~\s2_msel_arb1_state_reg[2]/NET0131  & ~n12027 ;
  assign n12029 = \s2_msel_arb1_state_reg[1]/NET0131  & ~n12028 ;
  assign n12030 = ~n12025 & ~n12029 ;
  assign n12031 = ~n12023 & ~n12030 ;
  assign n12032 = n5136 & ~n5137 ;
  assign n12033 = n5119 & ~n12032 ;
  assign n12034 = n5134 & n7398 ;
  assign n12035 = ~n12033 & n12034 ;
  assign n12036 = \s2_msel_arb1_state_reg[0]/NET0131  & n7389 ;
  assign n12037 = ~n5111 & n12036 ;
  assign n12038 = ~n12006 & n12037 ;
  assign n12039 = ~n12035 & ~n12038 ;
  assign n12040 = ~n12031 & n12039 ;
  assign n12041 = n12017 & n12040 ;
  assign n12042 = ~n5158 & ~n5169 ;
  assign n12043 = ~n5149 & ~n12042 ;
  assign n12044 = n5148 & n5157 ;
  assign n12045 = ~\s3_msel_arb1_state_reg[2]/NET0131  & ~n5157 ;
  assign n12046 = ~n5152 & ~n12045 ;
  assign n12047 = ~n12044 & ~n12046 ;
  assign n12048 = ~n12043 & n12047 ;
  assign n12049 = ~\s3_msel_arb1_state_reg[1]/NET0131  & ~n12048 ;
  assign n12050 = \s3_msel_arb1_state_reg[1]/NET0131  & ~n5146 ;
  assign n12051 = ~n7677 & ~n12050 ;
  assign n12052 = ~n5152 & n5157 ;
  assign n12053 = n5160 & ~n7677 ;
  assign n12054 = ~n12052 & n12053 ;
  assign n12055 = ~n12051 & ~n12054 ;
  assign n12056 = \s3_msel_arb1_state_reg[0]/NET0131  & n12055 ;
  assign n12057 = \s3_msel_arb1_state_reg[1]/NET0131  & ~\s3_msel_arb1_state_reg[2]/NET0131  ;
  assign n12058 = n5160 & ~n12052 ;
  assign n12059 = ~n5147 & n12050 ;
  assign n12060 = ~n12058 & n12059 ;
  assign n12061 = ~n12057 & ~n12060 ;
  assign n12062 = ~n12056 & n12061 ;
  assign n12063 = ~n12049 & n12062 ;
  assign n12064 = n5148 & ~n5160 ;
  assign n12065 = ~n5150 & n12057 ;
  assign n12066 = ~n12064 & n12065 ;
  assign n12067 = ~n5151 & n12066 ;
  assign n12068 = ~n5157 & n5160 ;
  assign n12069 = n5148 & ~n12068 ;
  assign n12070 = ~n5151 & n7722 ;
  assign n12071 = ~n12069 & n12070 ;
  assign n12072 = ~n12067 & ~n12071 ;
  assign n12073 = ~\rf_conf3_reg[7]/NET0131  & \s3_msel_arb1_state_reg[1]/NET0131  ;
  assign n12074 = n4530 & n12073 ;
  assign n12075 = ~n5145 & ~n12074 ;
  assign n12076 = n12045 & ~n12075 ;
  assign n12077 = n12072 & ~n12076 ;
  assign n12078 = ~n12063 & n12077 ;
  assign n12079 = n5192 & n5213 ;
  assign n12080 = ~n7976 & ~n12079 ;
  assign n12081 = \s4_msel_arb1_state_reg[1]/NET0131  & ~n12080 ;
  assign n12082 = ~\s4_msel_arb1_state_reg[0]/NET0131  & n5187 ;
  assign n12083 = n5192 & n12082 ;
  assign n12084 = ~\s4_msel_arb1_state_reg[0]/NET0131  & n5192 ;
  assign n12085 = ~\s4_msel_arb1_state_reg[1]/NET0131  & ~n12084 ;
  assign n12086 = n5213 & ~n5214 ;
  assign n12087 = ~n5188 & ~n12086 ;
  assign n12088 = ~n12085 & ~n12087 ;
  assign n12089 = ~n12083 & ~n12088 ;
  assign n12090 = ~n12081 & n12089 ;
  assign n12091 = \s4_msel_arb1_state_reg[2]/NET0131  & ~n12090 ;
  assign n12092 = ~n5212 & n7952 ;
  assign n12093 = n5192 & n12092 ;
  assign n12094 = ~n5202 & n12093 ;
  assign n12095 = ~n5189 & n5192 ;
  assign n12096 = n5214 & ~n12095 ;
  assign n12097 = ~n5200 & n7947 ;
  assign n12098 = ~n5202 & n12097 ;
  assign n12099 = ~n12096 & n12098 ;
  assign n12100 = ~n12094 & ~n12099 ;
  assign n12101 = ~n5196 & ~n5206 ;
  assign n12102 = ~n12095 & n12101 ;
  assign n12103 = n7952 & ~n12102 ;
  assign n12104 = n5189 & ~n12086 ;
  assign n12105 = ~n5191 & n7987 ;
  assign n12106 = ~n12104 & n12105 ;
  assign n12107 = ~n12103 & ~n12106 ;
  assign n12108 = n12100 & n12107 ;
  assign n12109 = ~n12091 & n12108 ;
  assign n12110 = ~\s5_msel_arb1_state_reg[2]/NET0131  & ~n5239 ;
  assign n12111 = ~n5231 & n5236 ;
  assign n12112 = ~n12110 & ~n12111 ;
  assign n12113 = n5259 & ~n12112 ;
  assign n12114 = \s5_msel_arb1_state_reg[2]/NET0131  & ~n5231 ;
  assign n12115 = n5228 & ~n5239 ;
  assign n12116 = ~n12114 & ~n12115 ;
  assign n12117 = ~n5234 & ~n8278 ;
  assign n12118 = ~n12116 & n12117 ;
  assign n12119 = \s5_msel_arb1_state_reg[1]/NET0131  & ~n12118 ;
  assign n12120 = ~n12113 & n12119 ;
  assign n12121 = ~n5236 & n5239 ;
  assign n12122 = n5228 & ~n12121 ;
  assign n12123 = n5242 & ~n8264 ;
  assign n12124 = ~n12122 & n12123 ;
  assign n12125 = ~n5228 & n5231 ;
  assign n12126 = n5236 & ~n12125 ;
  assign n12127 = ~n5238 & n8240 ;
  assign n12128 = ~n12126 & n12127 ;
  assign n12129 = ~n12124 & ~n12128 ;
  assign n12130 = ~n12120 & n12129 ;
  assign n12131 = ~\s6_msel_arb1_state_reg[2]/NET0131  & ~n5282 ;
  assign n12132 = ~n5274 & n5279 ;
  assign n12133 = ~n12131 & ~n12132 ;
  assign n12134 = n5302 & ~n12133 ;
  assign n12135 = \s6_msel_arb1_state_reg[2]/NET0131  & ~n5274 ;
  assign n12136 = n5271 & ~n5282 ;
  assign n12137 = ~n12135 & ~n12136 ;
  assign n12138 = ~n5277 & ~n8532 ;
  assign n12139 = ~n12137 & n12138 ;
  assign n12140 = \s6_msel_arb1_state_reg[1]/NET0131  & ~n12139 ;
  assign n12141 = ~n12134 & n12140 ;
  assign n12142 = ~n5279 & n5282 ;
  assign n12143 = n5271 & ~n12142 ;
  assign n12144 = n5285 & ~n8518 ;
  assign n12145 = ~n12143 & n12144 ;
  assign n12146 = ~n5271 & n5274 ;
  assign n12147 = n5279 & ~n12146 ;
  assign n12148 = ~n5281 & n8494 ;
  assign n12149 = ~n12147 & n12148 ;
  assign n12150 = ~n12145 & ~n12149 ;
  assign n12151 = ~n12141 & n12150 ;
  assign n12152 = ~n5314 & n5324 ;
  assign n12153 = n5321 & ~n12152 ;
  assign n12154 = ~\rf_conf7_reg[5]/NET0131  & ~\s7_msel_arb1_state_reg[0]/NET0131  ;
  assign n12155 = n4737 & n12154 ;
  assign n12156 = n8745 & ~n12155 ;
  assign n12157 = ~n12153 & n12156 ;
  assign n12158 = n5317 & ~n5321 ;
  assign n12159 = n5314 & ~n12158 ;
  assign n12160 = ~n5330 & n5335 ;
  assign n12161 = ~n12159 & n12160 ;
  assign n12162 = ~n12157 & ~n12161 ;
  assign n12163 = \s7_msel_arb1_state_reg[1]/NET0131  & ~n12162 ;
  assign n12164 = n5321 & ~n5324 ;
  assign n12165 = n5317 & ~n12164 ;
  assign n12166 = ~\s7_msel_arb1_state_reg[2]/NET0131  & n5341 ;
  assign n12167 = ~n12165 & n12166 ;
  assign n12168 = ~\rf_conf7_reg[9]/NET0131  & ~\s7_msel_arb1_state_reg[0]/NET0131  ;
  assign n12169 = n4720 & n12168 ;
  assign n12170 = \s7_msel_arb1_state_reg[2]/NET0131  & ~n5319 ;
  assign n12171 = ~n12169 & n12170 ;
  assign n12172 = ~\s7_msel_arb1_state_reg[1]/NET0131  & ~n12171 ;
  assign n12173 = n5314 & ~n5317 ;
  assign n12174 = ~\s7_msel_arb1_state_reg[1]/NET0131  & n5324 ;
  assign n12175 = ~n12173 & n12174 ;
  assign n12176 = ~n12172 & ~n12175 ;
  assign n12177 = ~n12167 & ~n12176 ;
  assign n12178 = ~n12163 & ~n12177 ;
  assign n12179 = ~\s8_msel_arb1_state_reg[2]/NET0131  & ~n5363 ;
  assign n12180 = ~n5355 & n5360 ;
  assign n12181 = ~n12179 & ~n12180 ;
  assign n12182 = n5383 & ~n12181 ;
  assign n12183 = \s8_msel_arb1_state_reg[2]/NET0131  & ~n5355 ;
  assign n12184 = n5352 & ~n5363 ;
  assign n12185 = ~n12183 & ~n12184 ;
  assign n12186 = ~n5358 & ~n9072 ;
  assign n12187 = ~n12185 & n12186 ;
  assign n12188 = \s8_msel_arb1_state_reg[1]/NET0131  & ~n12187 ;
  assign n12189 = ~n12182 & n12188 ;
  assign n12190 = ~n5360 & n5363 ;
  assign n12191 = n5352 & ~n12190 ;
  assign n12192 = n5366 & ~n9058 ;
  assign n12193 = ~n12191 & n12192 ;
  assign n12194 = ~n5352 & n5355 ;
  assign n12195 = n5360 & ~n12194 ;
  assign n12196 = ~n5362 & n9034 ;
  assign n12197 = ~n12195 & n12196 ;
  assign n12198 = ~n12193 & ~n12197 ;
  assign n12199 = ~n12189 & n12198 ;
  assign n12200 = ~\s9_msel_arb1_state_reg[2]/NET0131  & ~n5414 ;
  assign n12201 = ~n5402 & n5409 ;
  assign n12202 = ~n12200 & ~n12201 ;
  assign n12203 = n5434 & ~n12202 ;
  assign n12204 = \s9_msel_arb1_state_reg[2]/NET0131  & ~n5402 ;
  assign n12205 = n5397 & ~n5414 ;
  assign n12206 = ~n12204 & ~n12205 ;
  assign n12207 = ~n5406 & ~n9324 ;
  assign n12208 = ~n12206 & n12207 ;
  assign n12209 = \s9_msel_arb1_state_reg[1]/NET0131  & ~n12208 ;
  assign n12210 = ~n12203 & n12209 ;
  assign n12211 = ~n5409 & n5414 ;
  assign n12212 = n5397 & ~n12211 ;
  assign n12213 = n5417 & ~n9310 ;
  assign n12214 = ~n12212 & n12213 ;
  assign n12215 = ~n5397 & n5402 ;
  assign n12216 = n5409 & ~n12215 ;
  assign n12217 = ~n5413 & n9286 ;
  assign n12218 = ~n12216 & n12217 ;
  assign n12219 = ~n12214 & ~n12218 ;
  assign n12220 = ~n12210 & n12219 ;
  assign n12221 = ~\s0_msel_arb1_state_reg[2]/NET0131  & ~n5457 ;
  assign n12222 = ~n5449 & n5454 ;
  assign n12223 = ~n12221 & ~n12222 ;
  assign n12224 = n5477 & ~n12223 ;
  assign n12225 = \s0_msel_arb1_state_reg[2]/NET0131  & ~n5449 ;
  assign n12226 = n5446 & ~n5457 ;
  assign n12227 = ~n12225 & ~n12226 ;
  assign n12228 = ~n5452 & ~n9603 ;
  assign n12229 = ~n12227 & n12228 ;
  assign n12230 = \s0_msel_arb1_state_reg[1]/NET0131  & ~n12229 ;
  assign n12231 = ~n12224 & n12230 ;
  assign n12232 = ~n5454 & n5457 ;
  assign n12233 = n5446 & ~n12232 ;
  assign n12234 = n5460 & ~n9589 ;
  assign n12235 = ~n12233 & n12234 ;
  assign n12236 = ~n5446 & n5449 ;
  assign n12237 = n5454 & ~n12236 ;
  assign n12238 = ~n5456 & n9565 ;
  assign n12239 = ~n12237 & n12238 ;
  assign n12240 = ~n12235 & ~n12239 ;
  assign n12241 = ~n12231 & n12240 ;
  assign n12242 = n3785 & n3802 ;
  assign n12243 = ~\s15_msel_pri_out_reg[1]/NET0131  & ~\s15_next_reg/P0001  ;
  assign n12244 = ~rst_i_pad & ~n12243 ;
  assign n12245 = ~n12242 & n12244 ;
  assign n12246 = \m7_data_i[0]_pad  & ~n1910 ;
  assign n12247 = n1938 & n12246 ;
  assign n12248 = \m6_data_i[0]_pad  & ~n1925 ;
  assign n12249 = n1918 & n12248 ;
  assign n12250 = ~n12247 & ~n12249 ;
  assign n12251 = \m5_data_i[0]_pad  & ~n1910 ;
  assign n12252 = n1941 & n12251 ;
  assign n12253 = \m0_data_i[0]_pad  & n1925 ;
  assign n12254 = n1931 & n12253 ;
  assign n12255 = ~n12252 & ~n12254 ;
  assign n12256 = n12250 & n12255 ;
  assign n12257 = \m4_data_i[0]_pad  & n1925 ;
  assign n12258 = n1918 & n12257 ;
  assign n12259 = \m1_data_i[0]_pad  & n1910 ;
  assign n12260 = n1941 & n12259 ;
  assign n12261 = ~n12258 & ~n12260 ;
  assign n12262 = \m3_data_i[0]_pad  & n1910 ;
  assign n12263 = n1938 & n12262 ;
  assign n12264 = \m2_data_i[0]_pad  & ~n1925 ;
  assign n12265 = n1931 & n12264 ;
  assign n12266 = ~n12263 & ~n12265 ;
  assign n12267 = n12261 & n12266 ;
  assign n12268 = n12256 & n12267 ;
  assign n12269 = \rf_rf_we_reg/P0001  & ~n12268 ;
  assign n12270 = n2044 & n12269 ;
  assign n12271 = \rf_rf_we_reg/P0001  & n2044 ;
  assign n12272 = \rf_conf0_reg[0]/NET0131  & ~n12271 ;
  assign n12273 = ~n12270 & ~n12272 ;
  assign n12274 = \m7_data_i[10]_pad  & ~n1910 ;
  assign n12275 = n1938 & n12274 ;
  assign n12276 = \m6_data_i[10]_pad  & ~n1925 ;
  assign n12277 = n1918 & n12276 ;
  assign n12278 = ~n12275 & ~n12277 ;
  assign n12279 = \m5_data_i[10]_pad  & ~n1910 ;
  assign n12280 = n1941 & n12279 ;
  assign n12281 = \m2_data_i[10]_pad  & ~n1925 ;
  assign n12282 = n1931 & n12281 ;
  assign n12283 = ~n12280 & ~n12282 ;
  assign n12284 = n12278 & n12283 ;
  assign n12285 = \m4_data_i[10]_pad  & n1925 ;
  assign n12286 = n1918 & n12285 ;
  assign n12287 = \m3_data_i[10]_pad  & n1910 ;
  assign n12288 = n1938 & n12287 ;
  assign n12289 = ~n12286 & ~n12288 ;
  assign n12290 = \m1_data_i[10]_pad  & n1910 ;
  assign n12291 = n1941 & n12290 ;
  assign n12292 = \m0_data_i[10]_pad  & n1925 ;
  assign n12293 = n1931 & n12292 ;
  assign n12294 = ~n12291 & ~n12293 ;
  assign n12295 = n12289 & n12294 ;
  assign n12296 = n12284 & n12295 ;
  assign n12297 = \rf_rf_we_reg/P0001  & ~n12296 ;
  assign n12298 = n2044 & n12297 ;
  assign n12299 = \rf_conf0_reg[10]/NET0131  & ~n12271 ;
  assign n12300 = ~n12298 & ~n12299 ;
  assign n12301 = \m7_data_i[11]_pad  & ~n1910 ;
  assign n12302 = n1938 & n12301 ;
  assign n12303 = \m6_data_i[11]_pad  & ~n1925 ;
  assign n12304 = n1918 & n12303 ;
  assign n12305 = ~n12302 & ~n12304 ;
  assign n12306 = \m5_data_i[11]_pad  & ~n1910 ;
  assign n12307 = n1941 & n12306 ;
  assign n12308 = \m2_data_i[11]_pad  & ~n1925 ;
  assign n12309 = n1931 & n12308 ;
  assign n12310 = ~n12307 & ~n12309 ;
  assign n12311 = n12305 & n12310 ;
  assign n12312 = \m4_data_i[11]_pad  & n1925 ;
  assign n12313 = n1918 & n12312 ;
  assign n12314 = \m3_data_i[11]_pad  & n1910 ;
  assign n12315 = n1938 & n12314 ;
  assign n12316 = ~n12313 & ~n12315 ;
  assign n12317 = \m1_data_i[11]_pad  & n1910 ;
  assign n12318 = n1941 & n12317 ;
  assign n12319 = \m0_data_i[11]_pad  & n1925 ;
  assign n12320 = n1931 & n12319 ;
  assign n12321 = ~n12318 & ~n12320 ;
  assign n12322 = n12316 & n12321 ;
  assign n12323 = n12311 & n12322 ;
  assign n12324 = \rf_rf_we_reg/P0001  & ~n12323 ;
  assign n12325 = n2044 & n12324 ;
  assign n12326 = \rf_conf0_reg[11]/NET0131  & ~n12271 ;
  assign n12327 = ~n12325 & ~n12326 ;
  assign n12328 = \m7_data_i[12]_pad  & ~n1910 ;
  assign n12329 = n1938 & n12328 ;
  assign n12330 = \m6_data_i[12]_pad  & ~n1925 ;
  assign n12331 = n1918 & n12330 ;
  assign n12332 = ~n12329 & ~n12331 ;
  assign n12333 = \m5_data_i[12]_pad  & ~n1910 ;
  assign n12334 = n1941 & n12333 ;
  assign n12335 = \m2_data_i[12]_pad  & ~n1925 ;
  assign n12336 = n1931 & n12335 ;
  assign n12337 = ~n12334 & ~n12336 ;
  assign n12338 = n12332 & n12337 ;
  assign n12339 = \m4_data_i[12]_pad  & n1925 ;
  assign n12340 = n1918 & n12339 ;
  assign n12341 = \m3_data_i[12]_pad  & n1910 ;
  assign n12342 = n1938 & n12341 ;
  assign n12343 = ~n12340 & ~n12342 ;
  assign n12344 = \m1_data_i[12]_pad  & n1910 ;
  assign n12345 = n1941 & n12344 ;
  assign n12346 = \m0_data_i[12]_pad  & n1925 ;
  assign n12347 = n1931 & n12346 ;
  assign n12348 = ~n12345 & ~n12347 ;
  assign n12349 = n12343 & n12348 ;
  assign n12350 = n12338 & n12349 ;
  assign n12351 = \rf_rf_we_reg/P0001  & ~n12350 ;
  assign n12352 = n2044 & n12351 ;
  assign n12353 = \rf_conf0_reg[12]/NET0131  & ~n12271 ;
  assign n12354 = ~n12352 & ~n12353 ;
  assign n12355 = \m7_data_i[13]_pad  & ~n1910 ;
  assign n12356 = n1938 & n12355 ;
  assign n12357 = \m6_data_i[13]_pad  & ~n1925 ;
  assign n12358 = n1918 & n12357 ;
  assign n12359 = ~n12356 & ~n12358 ;
  assign n12360 = \m5_data_i[13]_pad  & ~n1910 ;
  assign n12361 = n1941 & n12360 ;
  assign n12362 = \m2_data_i[13]_pad  & ~n1925 ;
  assign n12363 = n1931 & n12362 ;
  assign n12364 = ~n12361 & ~n12363 ;
  assign n12365 = n12359 & n12364 ;
  assign n12366 = \m4_data_i[13]_pad  & n1925 ;
  assign n12367 = n1918 & n12366 ;
  assign n12368 = \m3_data_i[13]_pad  & n1910 ;
  assign n12369 = n1938 & n12368 ;
  assign n12370 = ~n12367 & ~n12369 ;
  assign n12371 = \m1_data_i[13]_pad  & n1910 ;
  assign n12372 = n1941 & n12371 ;
  assign n12373 = \m0_data_i[13]_pad  & n1925 ;
  assign n12374 = n1931 & n12373 ;
  assign n12375 = ~n12372 & ~n12374 ;
  assign n12376 = n12370 & n12375 ;
  assign n12377 = n12365 & n12376 ;
  assign n12378 = \rf_rf_we_reg/P0001  & ~n12377 ;
  assign n12379 = n2044 & n12378 ;
  assign n12380 = \rf_conf0_reg[13]/NET0131  & ~n12271 ;
  assign n12381 = ~n12379 & ~n12380 ;
  assign n12382 = \m7_data_i[14]_pad  & ~n1910 ;
  assign n12383 = n1938 & n12382 ;
  assign n12384 = \m6_data_i[14]_pad  & ~n1925 ;
  assign n12385 = n1918 & n12384 ;
  assign n12386 = ~n12383 & ~n12385 ;
  assign n12387 = \m5_data_i[14]_pad  & ~n1910 ;
  assign n12388 = n1941 & n12387 ;
  assign n12389 = \m2_data_i[14]_pad  & ~n1925 ;
  assign n12390 = n1931 & n12389 ;
  assign n12391 = ~n12388 & ~n12390 ;
  assign n12392 = n12386 & n12391 ;
  assign n12393 = \m4_data_i[14]_pad  & n1925 ;
  assign n12394 = n1918 & n12393 ;
  assign n12395 = \m3_data_i[14]_pad  & n1910 ;
  assign n12396 = n1938 & n12395 ;
  assign n12397 = ~n12394 & ~n12396 ;
  assign n12398 = \m1_data_i[14]_pad  & n1910 ;
  assign n12399 = n1941 & n12398 ;
  assign n12400 = \m0_data_i[14]_pad  & n1925 ;
  assign n12401 = n1931 & n12400 ;
  assign n12402 = ~n12399 & ~n12401 ;
  assign n12403 = n12397 & n12402 ;
  assign n12404 = n12392 & n12403 ;
  assign n12405 = \rf_rf_we_reg/P0001  & ~n12404 ;
  assign n12406 = n2044 & n12405 ;
  assign n12407 = \rf_conf0_reg[14]/NET0131  & ~n12271 ;
  assign n12408 = ~n12406 & ~n12407 ;
  assign n12409 = \m7_data_i[15]_pad  & ~n1910 ;
  assign n12410 = n1938 & n12409 ;
  assign n12411 = \m6_data_i[15]_pad  & ~n1925 ;
  assign n12412 = n1918 & n12411 ;
  assign n12413 = ~n12410 & ~n12412 ;
  assign n12414 = \m5_data_i[15]_pad  & ~n1910 ;
  assign n12415 = n1941 & n12414 ;
  assign n12416 = \m0_data_i[15]_pad  & n1925 ;
  assign n12417 = n1931 & n12416 ;
  assign n12418 = ~n12415 & ~n12417 ;
  assign n12419 = n12413 & n12418 ;
  assign n12420 = \m4_data_i[15]_pad  & n1925 ;
  assign n12421 = n1918 & n12420 ;
  assign n12422 = \m1_data_i[15]_pad  & n1910 ;
  assign n12423 = n1941 & n12422 ;
  assign n12424 = ~n12421 & ~n12423 ;
  assign n12425 = \m3_data_i[15]_pad  & n1910 ;
  assign n12426 = n1938 & n12425 ;
  assign n12427 = \m2_data_i[15]_pad  & ~n1925 ;
  assign n12428 = n1931 & n12427 ;
  assign n12429 = ~n12426 & ~n12428 ;
  assign n12430 = n12424 & n12429 ;
  assign n12431 = n12419 & n12430 ;
  assign n12432 = \rf_rf_we_reg/P0001  & ~n12431 ;
  assign n12433 = n2044 & n12432 ;
  assign n12434 = \rf_conf0_reg[15]/NET0131  & ~n12271 ;
  assign n12435 = ~n12433 & ~n12434 ;
  assign n12436 = \m7_data_i[1]_pad  & ~n1910 ;
  assign n12437 = n1938 & n12436 ;
  assign n12438 = \m6_data_i[1]_pad  & ~n1925 ;
  assign n12439 = n1918 & n12438 ;
  assign n12440 = ~n12437 & ~n12439 ;
  assign n12441 = \m5_data_i[1]_pad  & ~n1910 ;
  assign n12442 = n1941 & n12441 ;
  assign n12443 = \m0_data_i[1]_pad  & n1925 ;
  assign n12444 = n1931 & n12443 ;
  assign n12445 = ~n12442 & ~n12444 ;
  assign n12446 = n12440 & n12445 ;
  assign n12447 = \m4_data_i[1]_pad  & n1925 ;
  assign n12448 = n1918 & n12447 ;
  assign n12449 = \m1_data_i[1]_pad  & n1910 ;
  assign n12450 = n1941 & n12449 ;
  assign n12451 = ~n12448 & ~n12450 ;
  assign n12452 = \m3_data_i[1]_pad  & n1910 ;
  assign n12453 = n1938 & n12452 ;
  assign n12454 = \m2_data_i[1]_pad  & ~n1925 ;
  assign n12455 = n1931 & n12454 ;
  assign n12456 = ~n12453 & ~n12455 ;
  assign n12457 = n12451 & n12456 ;
  assign n12458 = n12446 & n12457 ;
  assign n12459 = \rf_rf_we_reg/P0001  & ~n12458 ;
  assign n12460 = n2044 & n12459 ;
  assign n12461 = \rf_conf0_reg[1]/NET0131  & ~n12271 ;
  assign n12462 = ~n12460 & ~n12461 ;
  assign n12463 = \m7_data_i[2]_pad  & ~n1910 ;
  assign n12464 = n1938 & n12463 ;
  assign n12465 = \m6_data_i[2]_pad  & ~n1925 ;
  assign n12466 = n1918 & n12465 ;
  assign n12467 = ~n12464 & ~n12466 ;
  assign n12468 = \m5_data_i[2]_pad  & ~n1910 ;
  assign n12469 = n1941 & n12468 ;
  assign n12470 = \m2_data_i[2]_pad  & ~n1925 ;
  assign n12471 = n1931 & n12470 ;
  assign n12472 = ~n12469 & ~n12471 ;
  assign n12473 = n12467 & n12472 ;
  assign n12474 = \m4_data_i[2]_pad  & n1925 ;
  assign n12475 = n1918 & n12474 ;
  assign n12476 = \m3_data_i[2]_pad  & n1910 ;
  assign n12477 = n1938 & n12476 ;
  assign n12478 = ~n12475 & ~n12477 ;
  assign n12479 = \m1_data_i[2]_pad  & n1910 ;
  assign n12480 = n1941 & n12479 ;
  assign n12481 = \m0_data_i[2]_pad  & n1925 ;
  assign n12482 = n1931 & n12481 ;
  assign n12483 = ~n12480 & ~n12482 ;
  assign n12484 = n12478 & n12483 ;
  assign n12485 = n12473 & n12484 ;
  assign n12486 = \rf_rf_we_reg/P0001  & ~n12485 ;
  assign n12487 = n2044 & n12486 ;
  assign n12488 = \rf_conf0_reg[2]/NET0131  & ~n12271 ;
  assign n12489 = ~n12487 & ~n12488 ;
  assign n12490 = \m7_data_i[3]_pad  & ~n1910 ;
  assign n12491 = n1938 & n12490 ;
  assign n12492 = \m6_data_i[3]_pad  & ~n1925 ;
  assign n12493 = n1918 & n12492 ;
  assign n12494 = ~n12491 & ~n12493 ;
  assign n12495 = \m5_data_i[3]_pad  & ~n1910 ;
  assign n12496 = n1941 & n12495 ;
  assign n12497 = \m2_data_i[3]_pad  & ~n1925 ;
  assign n12498 = n1931 & n12497 ;
  assign n12499 = ~n12496 & ~n12498 ;
  assign n12500 = n12494 & n12499 ;
  assign n12501 = \m4_data_i[3]_pad  & n1925 ;
  assign n12502 = n1918 & n12501 ;
  assign n12503 = \m3_data_i[3]_pad  & n1910 ;
  assign n12504 = n1938 & n12503 ;
  assign n12505 = ~n12502 & ~n12504 ;
  assign n12506 = \m1_data_i[3]_pad  & n1910 ;
  assign n12507 = n1941 & n12506 ;
  assign n12508 = \m0_data_i[3]_pad  & n1925 ;
  assign n12509 = n1931 & n12508 ;
  assign n12510 = ~n12507 & ~n12509 ;
  assign n12511 = n12505 & n12510 ;
  assign n12512 = n12500 & n12511 ;
  assign n12513 = \rf_rf_we_reg/P0001  & ~n12512 ;
  assign n12514 = n2044 & n12513 ;
  assign n12515 = \rf_conf0_reg[3]/NET0131  & ~n12271 ;
  assign n12516 = ~n12514 & ~n12515 ;
  assign n12517 = \m7_data_i[4]_pad  & ~n1910 ;
  assign n12518 = n1938 & n12517 ;
  assign n12519 = \m6_data_i[4]_pad  & ~n1925 ;
  assign n12520 = n1918 & n12519 ;
  assign n12521 = ~n12518 & ~n12520 ;
  assign n12522 = \m5_data_i[4]_pad  & ~n1910 ;
  assign n12523 = n1941 & n12522 ;
  assign n12524 = \m2_data_i[4]_pad  & ~n1925 ;
  assign n12525 = n1931 & n12524 ;
  assign n12526 = ~n12523 & ~n12525 ;
  assign n12527 = n12521 & n12526 ;
  assign n12528 = \m4_data_i[4]_pad  & n1925 ;
  assign n12529 = n1918 & n12528 ;
  assign n12530 = \m3_data_i[4]_pad  & n1910 ;
  assign n12531 = n1938 & n12530 ;
  assign n12532 = ~n12529 & ~n12531 ;
  assign n12533 = \m1_data_i[4]_pad  & n1910 ;
  assign n12534 = n1941 & n12533 ;
  assign n12535 = \m0_data_i[4]_pad  & n1925 ;
  assign n12536 = n1931 & n12535 ;
  assign n12537 = ~n12534 & ~n12536 ;
  assign n12538 = n12532 & n12537 ;
  assign n12539 = n12527 & n12538 ;
  assign n12540 = \rf_rf_we_reg/P0001  & ~n12539 ;
  assign n12541 = n2044 & n12540 ;
  assign n12542 = \rf_conf0_reg[4]/NET0131  & ~n12271 ;
  assign n12543 = ~n12541 & ~n12542 ;
  assign n12544 = \m3_data_i[5]_pad  & n1910 ;
  assign n12545 = n1938 & n12544 ;
  assign n12546 = \m2_data_i[5]_pad  & ~n1925 ;
  assign n12547 = n1931 & n12546 ;
  assign n12548 = ~n12545 & ~n12547 ;
  assign n12549 = \m5_data_i[5]_pad  & ~n1910 ;
  assign n12550 = n1941 & n12549 ;
  assign n12551 = \m0_data_i[5]_pad  & n1925 ;
  assign n12552 = n1931 & n12551 ;
  assign n12553 = ~n12550 & ~n12552 ;
  assign n12554 = n12548 & n12553 ;
  assign n12555 = \m4_data_i[5]_pad  & n1925 ;
  assign n12556 = n1918 & n12555 ;
  assign n12557 = \m1_data_i[5]_pad  & n1910 ;
  assign n12558 = n1941 & n12557 ;
  assign n12559 = ~n12556 & ~n12558 ;
  assign n12560 = \m7_data_i[5]_pad  & ~n1910 ;
  assign n12561 = n1938 & n12560 ;
  assign n12562 = \m6_data_i[5]_pad  & ~n1925 ;
  assign n12563 = n1918 & n12562 ;
  assign n12564 = ~n12561 & ~n12563 ;
  assign n12565 = n12559 & n12564 ;
  assign n12566 = n12554 & n12565 ;
  assign n12567 = \rf_rf_we_reg/P0001  & ~n12566 ;
  assign n12568 = n2044 & n12567 ;
  assign n12569 = \rf_conf0_reg[5]/NET0131  & ~n12271 ;
  assign n12570 = ~n12568 & ~n12569 ;
  assign n12571 = \m7_data_i[6]_pad  & ~n1910 ;
  assign n12572 = n1938 & n12571 ;
  assign n12573 = \m6_data_i[6]_pad  & ~n1925 ;
  assign n12574 = n1918 & n12573 ;
  assign n12575 = ~n12572 & ~n12574 ;
  assign n12576 = \m5_data_i[6]_pad  & ~n1910 ;
  assign n12577 = n1941 & n12576 ;
  assign n12578 = \m2_data_i[6]_pad  & ~n1925 ;
  assign n12579 = n1931 & n12578 ;
  assign n12580 = ~n12577 & ~n12579 ;
  assign n12581 = n12575 & n12580 ;
  assign n12582 = \m4_data_i[6]_pad  & n1925 ;
  assign n12583 = n1918 & n12582 ;
  assign n12584 = \m3_data_i[6]_pad  & n1910 ;
  assign n12585 = n1938 & n12584 ;
  assign n12586 = ~n12583 & ~n12585 ;
  assign n12587 = \m1_data_i[6]_pad  & n1910 ;
  assign n12588 = n1941 & n12587 ;
  assign n12589 = \m0_data_i[6]_pad  & n1925 ;
  assign n12590 = n1931 & n12589 ;
  assign n12591 = ~n12588 & ~n12590 ;
  assign n12592 = n12586 & n12591 ;
  assign n12593 = n12581 & n12592 ;
  assign n12594 = \rf_rf_we_reg/P0001  & ~n12593 ;
  assign n12595 = n2044 & n12594 ;
  assign n12596 = \rf_conf0_reg[6]/NET0131  & ~n12271 ;
  assign n12597 = ~n12595 & ~n12596 ;
  assign n12598 = \m7_data_i[7]_pad  & ~n1910 ;
  assign n12599 = n1938 & n12598 ;
  assign n12600 = \m6_data_i[7]_pad  & ~n1925 ;
  assign n12601 = n1918 & n12600 ;
  assign n12602 = ~n12599 & ~n12601 ;
  assign n12603 = \m5_data_i[7]_pad  & ~n1910 ;
  assign n12604 = n1941 & n12603 ;
  assign n12605 = \m2_data_i[7]_pad  & ~n1925 ;
  assign n12606 = n1931 & n12605 ;
  assign n12607 = ~n12604 & ~n12606 ;
  assign n12608 = n12602 & n12607 ;
  assign n12609 = \m4_data_i[7]_pad  & n1925 ;
  assign n12610 = n1918 & n12609 ;
  assign n12611 = \m3_data_i[7]_pad  & n1910 ;
  assign n12612 = n1938 & n12611 ;
  assign n12613 = ~n12610 & ~n12612 ;
  assign n12614 = \m1_data_i[7]_pad  & n1910 ;
  assign n12615 = n1941 & n12614 ;
  assign n12616 = \m0_data_i[7]_pad  & n1925 ;
  assign n12617 = n1931 & n12616 ;
  assign n12618 = ~n12615 & ~n12617 ;
  assign n12619 = n12613 & n12618 ;
  assign n12620 = n12608 & n12619 ;
  assign n12621 = \rf_rf_we_reg/P0001  & ~n12620 ;
  assign n12622 = n2044 & n12621 ;
  assign n12623 = \rf_conf0_reg[7]/NET0131  & ~n12271 ;
  assign n12624 = ~n12622 & ~n12623 ;
  assign n12625 = \m7_data_i[8]_pad  & ~n1910 ;
  assign n12626 = n1938 & n12625 ;
  assign n12627 = \m6_data_i[8]_pad  & ~n1925 ;
  assign n12628 = n1918 & n12627 ;
  assign n12629 = ~n12626 & ~n12628 ;
  assign n12630 = \m5_data_i[8]_pad  & ~n1910 ;
  assign n12631 = n1941 & n12630 ;
  assign n12632 = \m0_data_i[8]_pad  & n1925 ;
  assign n12633 = n1931 & n12632 ;
  assign n12634 = ~n12631 & ~n12633 ;
  assign n12635 = n12629 & n12634 ;
  assign n12636 = \m4_data_i[8]_pad  & n1925 ;
  assign n12637 = n1918 & n12636 ;
  assign n12638 = \m1_data_i[8]_pad  & n1910 ;
  assign n12639 = n1941 & n12638 ;
  assign n12640 = ~n12637 & ~n12639 ;
  assign n12641 = \m3_data_i[8]_pad  & n1910 ;
  assign n12642 = n1938 & n12641 ;
  assign n12643 = \m2_data_i[8]_pad  & ~n1925 ;
  assign n12644 = n1931 & n12643 ;
  assign n12645 = ~n12642 & ~n12644 ;
  assign n12646 = n12640 & n12645 ;
  assign n12647 = n12635 & n12646 ;
  assign n12648 = \rf_rf_we_reg/P0001  & ~n12647 ;
  assign n12649 = n2044 & n12648 ;
  assign n12650 = \rf_conf0_reg[8]/NET0131  & ~n12271 ;
  assign n12651 = ~n12649 & ~n12650 ;
  assign n12652 = \m5_data_i[9]_pad  & ~n1910 ;
  assign n12653 = n1941 & n12652 ;
  assign n12654 = \m4_data_i[9]_pad  & n1925 ;
  assign n12655 = n1918 & n12654 ;
  assign n12656 = ~n12653 & ~n12655 ;
  assign n12657 = \m7_data_i[9]_pad  & ~n1910 ;
  assign n12658 = n1938 & n12657 ;
  assign n12659 = \m0_data_i[9]_pad  & n1925 ;
  assign n12660 = n1931 & n12659 ;
  assign n12661 = ~n12658 & ~n12660 ;
  assign n12662 = n12656 & n12661 ;
  assign n12663 = \m6_data_i[9]_pad  & ~n1925 ;
  assign n12664 = n1918 & n12663 ;
  assign n12665 = \m1_data_i[9]_pad  & n1910 ;
  assign n12666 = n1941 & n12665 ;
  assign n12667 = ~n12664 & ~n12666 ;
  assign n12668 = \m3_data_i[9]_pad  & n1910 ;
  assign n12669 = n1938 & n12668 ;
  assign n12670 = \m2_data_i[9]_pad  & ~n1925 ;
  assign n12671 = n1931 & n12670 ;
  assign n12672 = ~n12669 & ~n12671 ;
  assign n12673 = n12667 & n12672 ;
  assign n12674 = n12662 & n12673 ;
  assign n12675 = \rf_rf_we_reg/P0001  & ~n12674 ;
  assign n12676 = n2044 & n12675 ;
  assign n12677 = \rf_conf0_reg[9]/NET0131  & ~n12271 ;
  assign n12678 = ~n12676 & ~n12677 ;
  assign n12679 = n2065 & n12269 ;
  assign n12680 = \rf_rf_we_reg/P0001  & n2065 ;
  assign n12681 = \rf_conf10_reg[0]/NET0131  & ~n12680 ;
  assign n12682 = ~n12679 & ~n12681 ;
  assign n12683 = n2065 & n12297 ;
  assign n12684 = \rf_conf10_reg[10]/NET0131  & ~n12680 ;
  assign n12685 = ~n12683 & ~n12684 ;
  assign n12686 = n2065 & n12324 ;
  assign n12687 = \rf_conf10_reg[11]/NET0131  & ~n12680 ;
  assign n12688 = ~n12686 & ~n12687 ;
  assign n12689 = n2065 & n12351 ;
  assign n12690 = \rf_conf10_reg[12]/NET0131  & ~n12680 ;
  assign n12691 = ~n12689 & ~n12690 ;
  assign n12692 = n2065 & n12378 ;
  assign n12693 = \rf_conf10_reg[13]/NET0131  & ~n12680 ;
  assign n12694 = ~n12692 & ~n12693 ;
  assign n12695 = n2065 & n12432 ;
  assign n12696 = \rf_conf10_reg[15]/NET0131  & ~n12680 ;
  assign n12697 = ~n12695 & ~n12696 ;
  assign n12698 = n2065 & n12459 ;
  assign n12699 = \rf_conf10_reg[1]/NET0131  & ~n12680 ;
  assign n12700 = ~n12698 & ~n12699 ;
  assign n12701 = n2065 & n12405 ;
  assign n12702 = \rf_conf10_reg[14]/NET0131  & ~n12680 ;
  assign n12703 = ~n12701 & ~n12702 ;
  assign n12704 = n2065 & n12486 ;
  assign n12705 = \rf_conf10_reg[2]/NET0131  & ~n12680 ;
  assign n12706 = ~n12704 & ~n12705 ;
  assign n12707 = n2065 & n12513 ;
  assign n12708 = \rf_conf10_reg[3]/NET0131  & ~n12680 ;
  assign n12709 = ~n12707 & ~n12708 ;
  assign n12710 = n2065 & n12540 ;
  assign n12711 = \rf_conf10_reg[4]/NET0131  & ~n12680 ;
  assign n12712 = ~n12710 & ~n12711 ;
  assign n12713 = n2065 & n12567 ;
  assign n12714 = \rf_conf10_reg[5]/NET0131  & ~n12680 ;
  assign n12715 = ~n12713 & ~n12714 ;
  assign n12716 = n2065 & n12594 ;
  assign n12717 = \rf_conf10_reg[6]/NET0131  & ~n12680 ;
  assign n12718 = ~n12716 & ~n12717 ;
  assign n12719 = n2065 & n12621 ;
  assign n12720 = \rf_conf10_reg[7]/NET0131  & ~n12680 ;
  assign n12721 = ~n12719 & ~n12720 ;
  assign n12722 = n2065 & n12648 ;
  assign n12723 = \rf_conf10_reg[8]/NET0131  & ~n12680 ;
  assign n12724 = ~n12722 & ~n12723 ;
  assign n12725 = n2065 & n12675 ;
  assign n12726 = \rf_conf10_reg[9]/NET0131  & ~n12680 ;
  assign n12727 = ~n12725 & ~n12726 ;
  assign n12728 = n2059 & n12269 ;
  assign n12729 = \rf_rf_we_reg/P0001  & n2059 ;
  assign n12730 = \rf_conf11_reg[0]/NET0131  & ~n12729 ;
  assign n12731 = ~n12728 & ~n12730 ;
  assign n12732 = n2059 & n12297 ;
  assign n12733 = \rf_conf11_reg[10]/NET0131  & ~n12729 ;
  assign n12734 = ~n12732 & ~n12733 ;
  assign n12735 = n2059 & n12351 ;
  assign n12736 = \rf_conf11_reg[12]/NET0131  & ~n12729 ;
  assign n12737 = ~n12735 & ~n12736 ;
  assign n12738 = n2059 & n12324 ;
  assign n12739 = \rf_conf11_reg[11]/NET0131  & ~n12729 ;
  assign n12740 = ~n12738 & ~n12739 ;
  assign n12741 = n2059 & n12378 ;
  assign n12742 = \rf_conf11_reg[13]/NET0131  & ~n12729 ;
  assign n12743 = ~n12741 & ~n12742 ;
  assign n12744 = n2059 & n12405 ;
  assign n12745 = \rf_conf11_reg[14]/NET0131  & ~n12729 ;
  assign n12746 = ~n12744 & ~n12745 ;
  assign n12747 = n2059 & n12432 ;
  assign n12748 = \rf_conf11_reg[15]/NET0131  & ~n12729 ;
  assign n12749 = ~n12747 & ~n12748 ;
  assign n12750 = n2059 & n12459 ;
  assign n12751 = \rf_conf11_reg[1]/NET0131  & ~n12729 ;
  assign n12752 = ~n12750 & ~n12751 ;
  assign n12753 = n2059 & n12486 ;
  assign n12754 = \rf_conf11_reg[2]/NET0131  & ~n12729 ;
  assign n12755 = ~n12753 & ~n12754 ;
  assign n12756 = n2059 & n12513 ;
  assign n12757 = \rf_conf11_reg[3]/NET0131  & ~n12729 ;
  assign n12758 = ~n12756 & ~n12757 ;
  assign n12759 = n2059 & n12540 ;
  assign n12760 = \rf_conf11_reg[4]/NET0131  & ~n12729 ;
  assign n12761 = ~n12759 & ~n12760 ;
  assign n12762 = n2059 & n12567 ;
  assign n12763 = \rf_conf11_reg[5]/NET0131  & ~n12729 ;
  assign n12764 = ~n12762 & ~n12763 ;
  assign n12765 = n2059 & n12594 ;
  assign n12766 = \rf_conf11_reg[6]/NET0131  & ~n12729 ;
  assign n12767 = ~n12765 & ~n12766 ;
  assign n12768 = n2059 & n12621 ;
  assign n12769 = \rf_conf11_reg[7]/NET0131  & ~n12729 ;
  assign n12770 = ~n12768 & ~n12769 ;
  assign n12771 = n2059 & n12648 ;
  assign n12772 = \rf_conf11_reg[8]/NET0131  & ~n12729 ;
  assign n12773 = ~n12771 & ~n12772 ;
  assign n12774 = n2059 & n12675 ;
  assign n12775 = \rf_conf11_reg[9]/NET0131  & ~n12729 ;
  assign n12776 = ~n12774 & ~n12775 ;
  assign n12777 = n2032 & n12269 ;
  assign n12778 = \rf_rf_we_reg/P0001  & n2032 ;
  assign n12779 = \rf_conf12_reg[0]/NET0131  & ~n12778 ;
  assign n12780 = ~n12777 & ~n12779 ;
  assign n12781 = n2032 & n12297 ;
  assign n12782 = \rf_conf12_reg[10]/NET0131  & ~n12778 ;
  assign n12783 = ~n12781 & ~n12782 ;
  assign n12784 = n2032 & n12324 ;
  assign n12785 = \rf_conf12_reg[11]/NET0131  & ~n12778 ;
  assign n12786 = ~n12784 & ~n12785 ;
  assign n12787 = n2032 & n12351 ;
  assign n12788 = \rf_conf12_reg[12]/NET0131  & ~n12778 ;
  assign n12789 = ~n12787 & ~n12788 ;
  assign n12790 = n2032 & n12378 ;
  assign n12791 = \rf_conf12_reg[13]/NET0131  & ~n12778 ;
  assign n12792 = ~n12790 & ~n12791 ;
  assign n12793 = n2032 & n12405 ;
  assign n12794 = \rf_conf12_reg[14]/NET0131  & ~n12778 ;
  assign n12795 = ~n12793 & ~n12794 ;
  assign n12796 = n2032 & n12432 ;
  assign n12797 = \rf_conf12_reg[15]/NET0131  & ~n12778 ;
  assign n12798 = ~n12796 & ~n12797 ;
  assign n12799 = n2032 & n12459 ;
  assign n12800 = \rf_conf12_reg[1]/NET0131  & ~n12778 ;
  assign n12801 = ~n12799 & ~n12800 ;
  assign n12802 = n2032 & n12486 ;
  assign n12803 = \rf_conf12_reg[2]/NET0131  & ~n12778 ;
  assign n12804 = ~n12802 & ~n12803 ;
  assign n12805 = n2032 & n12513 ;
  assign n12806 = \rf_conf12_reg[3]/NET0131  & ~n12778 ;
  assign n12807 = ~n12805 & ~n12806 ;
  assign n12808 = n2032 & n12540 ;
  assign n12809 = \rf_conf12_reg[4]/NET0131  & ~n12778 ;
  assign n12810 = ~n12808 & ~n12809 ;
  assign n12811 = n2032 & n12567 ;
  assign n12812 = \rf_conf12_reg[5]/NET0131  & ~n12778 ;
  assign n12813 = ~n12811 & ~n12812 ;
  assign n12814 = n2032 & n12594 ;
  assign n12815 = \rf_conf12_reg[6]/NET0131  & ~n12778 ;
  assign n12816 = ~n12814 & ~n12815 ;
  assign n12817 = n2032 & n12621 ;
  assign n12818 = \rf_conf12_reg[7]/NET0131  & ~n12778 ;
  assign n12819 = ~n12817 & ~n12818 ;
  assign n12820 = n2032 & n12648 ;
  assign n12821 = \rf_conf12_reg[8]/NET0131  & ~n12778 ;
  assign n12822 = ~n12820 & ~n12821 ;
  assign n12823 = n2032 & n12675 ;
  assign n12824 = \rf_conf12_reg[9]/NET0131  & ~n12778 ;
  assign n12825 = ~n12823 & ~n12824 ;
  assign n12826 = n2068 & n12269 ;
  assign n12827 = \rf_rf_we_reg/P0001  & n2068 ;
  assign n12828 = \rf_conf13_reg[0]/NET0131  & ~n12827 ;
  assign n12829 = ~n12826 & ~n12828 ;
  assign n12830 = n2068 & n12324 ;
  assign n12831 = \rf_conf13_reg[11]/NET0131  & ~n12827 ;
  assign n12832 = ~n12830 & ~n12831 ;
  assign n12833 = n2068 & n12297 ;
  assign n12834 = \rf_conf13_reg[10]/NET0131  & ~n12827 ;
  assign n12835 = ~n12833 & ~n12834 ;
  assign n12836 = n2068 & n12351 ;
  assign n12837 = \rf_conf13_reg[12]/NET0131  & ~n12827 ;
  assign n12838 = ~n12836 & ~n12837 ;
  assign n12839 = n2068 & n12378 ;
  assign n12840 = \rf_conf13_reg[13]/NET0131  & ~n12827 ;
  assign n12841 = ~n12839 & ~n12840 ;
  assign n12842 = n2068 & n12405 ;
  assign n12843 = \rf_conf13_reg[14]/NET0131  & ~n12827 ;
  assign n12844 = ~n12842 & ~n12843 ;
  assign n12845 = n2068 & n12432 ;
  assign n12846 = \rf_conf13_reg[15]/NET0131  & ~n12827 ;
  assign n12847 = ~n12845 & ~n12846 ;
  assign n12848 = n2068 & n12459 ;
  assign n12849 = \rf_conf13_reg[1]/NET0131  & ~n12827 ;
  assign n12850 = ~n12848 & ~n12849 ;
  assign n12851 = n2068 & n12486 ;
  assign n12852 = \rf_conf13_reg[2]/NET0131  & ~n12827 ;
  assign n12853 = ~n12851 & ~n12852 ;
  assign n12854 = n2068 & n12513 ;
  assign n12855 = \rf_conf13_reg[3]/NET0131  & ~n12827 ;
  assign n12856 = ~n12854 & ~n12855 ;
  assign n12857 = n2068 & n12540 ;
  assign n12858 = \rf_conf13_reg[4]/NET0131  & ~n12827 ;
  assign n12859 = ~n12857 & ~n12858 ;
  assign n12860 = n2068 & n12567 ;
  assign n12861 = \rf_conf13_reg[5]/NET0131  & ~n12827 ;
  assign n12862 = ~n12860 & ~n12861 ;
  assign n12863 = n2068 & n12594 ;
  assign n12864 = \rf_conf13_reg[6]/NET0131  & ~n12827 ;
  assign n12865 = ~n12863 & ~n12864 ;
  assign n12866 = n2068 & n12621 ;
  assign n12867 = \rf_conf13_reg[7]/NET0131  & ~n12827 ;
  assign n12868 = ~n12866 & ~n12867 ;
  assign n12869 = n2068 & n12648 ;
  assign n12870 = \rf_conf13_reg[8]/NET0131  & ~n12827 ;
  assign n12871 = ~n12869 & ~n12870 ;
  assign n12872 = n2068 & n12675 ;
  assign n12873 = \rf_conf13_reg[9]/NET0131  & ~n12827 ;
  assign n12874 = ~n12872 & ~n12873 ;
  assign n12875 = n2035 & n12269 ;
  assign n12876 = \rf_rf_we_reg/P0001  & n2035 ;
  assign n12877 = \rf_conf14_reg[0]/NET0131  & ~n12876 ;
  assign n12878 = ~n12875 & ~n12877 ;
  assign n12879 = n2035 & n12297 ;
  assign n12880 = \rf_conf14_reg[10]/NET0131  & ~n12876 ;
  assign n12881 = ~n12879 & ~n12880 ;
  assign n12882 = n2035 & n12324 ;
  assign n12883 = \rf_conf14_reg[11]/NET0131  & ~n12876 ;
  assign n12884 = ~n12882 & ~n12883 ;
  assign n12885 = n2035 & n12378 ;
  assign n12886 = \rf_conf14_reg[13]/NET0131  & ~n12876 ;
  assign n12887 = ~n12885 & ~n12886 ;
  assign n12888 = n2035 & n12405 ;
  assign n12889 = \rf_conf14_reg[14]/NET0131  & ~n12876 ;
  assign n12890 = ~n12888 & ~n12889 ;
  assign n12891 = n2035 & n12351 ;
  assign n12892 = \rf_conf14_reg[12]/NET0131  & ~n12876 ;
  assign n12893 = ~n12891 & ~n12892 ;
  assign n12894 = n2035 & n12432 ;
  assign n12895 = \rf_conf14_reg[15]/NET0131  & ~n12876 ;
  assign n12896 = ~n12894 & ~n12895 ;
  assign n12897 = n2035 & n12459 ;
  assign n12898 = \rf_conf14_reg[1]/NET0131  & ~n12876 ;
  assign n12899 = ~n12897 & ~n12898 ;
  assign n12900 = n2035 & n12486 ;
  assign n12901 = \rf_conf14_reg[2]/NET0131  & ~n12876 ;
  assign n12902 = ~n12900 & ~n12901 ;
  assign n12903 = n2035 & n12513 ;
  assign n12904 = \rf_conf14_reg[3]/NET0131  & ~n12876 ;
  assign n12905 = ~n12903 & ~n12904 ;
  assign n12906 = n2035 & n12567 ;
  assign n12907 = \rf_conf14_reg[5]/NET0131  & ~n12876 ;
  assign n12908 = ~n12906 & ~n12907 ;
  assign n12909 = n2035 & n12540 ;
  assign n12910 = \rf_conf14_reg[4]/NET0131  & ~n12876 ;
  assign n12911 = ~n12909 & ~n12910 ;
  assign n12912 = n2035 & n12594 ;
  assign n12913 = \rf_conf14_reg[6]/NET0131  & ~n12876 ;
  assign n12914 = ~n12912 & ~n12913 ;
  assign n12915 = n2035 & n12621 ;
  assign n12916 = \rf_conf14_reg[7]/NET0131  & ~n12876 ;
  assign n12917 = ~n12915 & ~n12916 ;
  assign n12918 = n2035 & n12648 ;
  assign n12919 = \rf_conf14_reg[8]/NET0131  & ~n12876 ;
  assign n12920 = ~n12918 & ~n12919 ;
  assign n12921 = n2035 & n12675 ;
  assign n12922 = \rf_conf14_reg[9]/NET0131  & ~n12876 ;
  assign n12923 = ~n12921 & ~n12922 ;
  assign n12924 = n2070 & n12269 ;
  assign n12925 = \rf_rf_we_reg/P0001  & n2070 ;
  assign n12926 = \rf_conf15_reg[0]/NET0131  & ~n12925 ;
  assign n12927 = ~n12924 & ~n12926 ;
  assign n12928 = n2070 & n12297 ;
  assign n12929 = \rf_conf15_reg[10]/NET0131  & ~n12925 ;
  assign n12930 = ~n12928 & ~n12929 ;
  assign n12931 = n2070 & n12324 ;
  assign n12932 = \rf_conf15_reg[11]/NET0131  & ~n12925 ;
  assign n12933 = ~n12931 & ~n12932 ;
  assign n12934 = n2070 & n12351 ;
  assign n12935 = \rf_conf15_reg[12]/NET0131  & ~n12925 ;
  assign n12936 = ~n12934 & ~n12935 ;
  assign n12937 = n2070 & n12378 ;
  assign n12938 = \rf_conf15_reg[13]/NET0131  & ~n12925 ;
  assign n12939 = ~n12937 & ~n12938 ;
  assign n12940 = n2070 & n12405 ;
  assign n12941 = \rf_conf15_reg[14]/NET0131  & ~n12925 ;
  assign n12942 = ~n12940 & ~n12941 ;
  assign n12943 = n2070 & n12432 ;
  assign n12944 = \rf_conf15_reg[15]/NET0131  & ~n12925 ;
  assign n12945 = ~n12943 & ~n12944 ;
  assign n12946 = n2070 & n12459 ;
  assign n12947 = \rf_conf15_reg[1]/NET0131  & ~n12925 ;
  assign n12948 = ~n12946 & ~n12947 ;
  assign n12949 = n2070 & n12486 ;
  assign n12950 = \rf_conf15_reg[2]/NET0131  & ~n12925 ;
  assign n12951 = ~n12949 & ~n12950 ;
  assign n12952 = n2070 & n12513 ;
  assign n12953 = \rf_conf15_reg[3]/NET0131  & ~n12925 ;
  assign n12954 = ~n12952 & ~n12953 ;
  assign n12955 = n2070 & n12540 ;
  assign n12956 = \rf_conf15_reg[4]/NET0131  & ~n12925 ;
  assign n12957 = ~n12955 & ~n12956 ;
  assign n12958 = n2070 & n12567 ;
  assign n12959 = \rf_conf15_reg[5]/NET0131  & ~n12925 ;
  assign n12960 = ~n12958 & ~n12959 ;
  assign n12961 = n2070 & n12594 ;
  assign n12962 = \rf_conf15_reg[6]/NET0131  & ~n12925 ;
  assign n12963 = ~n12961 & ~n12962 ;
  assign n12964 = n2070 & n12648 ;
  assign n12965 = \rf_conf15_reg[8]/NET0131  & ~n12925 ;
  assign n12966 = ~n12964 & ~n12965 ;
  assign n12967 = n2070 & n12621 ;
  assign n12968 = \rf_conf15_reg[7]/NET0131  & ~n12925 ;
  assign n12969 = ~n12967 & ~n12968 ;
  assign n12970 = n2070 & n12675 ;
  assign n12971 = \rf_conf15_reg[9]/NET0131  & ~n12925 ;
  assign n12972 = ~n12970 & ~n12971 ;
  assign n12973 = n2041 & n12269 ;
  assign n12974 = \rf_rf_we_reg/P0001  & n2041 ;
  assign n12975 = \rf_conf1_reg[0]/NET0131  & ~n12974 ;
  assign n12976 = ~n12973 & ~n12975 ;
  assign n12977 = n2041 & n12297 ;
  assign n12978 = \rf_conf1_reg[10]/NET0131  & ~n12974 ;
  assign n12979 = ~n12977 & ~n12978 ;
  assign n12980 = n2041 & n12324 ;
  assign n12981 = \rf_conf1_reg[11]/NET0131  & ~n12974 ;
  assign n12982 = ~n12980 & ~n12981 ;
  assign n12983 = n2041 & n12378 ;
  assign n12984 = \rf_conf1_reg[13]/NET0131  & ~n12974 ;
  assign n12985 = ~n12983 & ~n12984 ;
  assign n12986 = n2041 & n12351 ;
  assign n12987 = \rf_conf1_reg[12]/NET0131  & ~n12974 ;
  assign n12988 = ~n12986 & ~n12987 ;
  assign n12989 = n2041 & n12405 ;
  assign n12990 = \rf_conf1_reg[14]/NET0131  & ~n12974 ;
  assign n12991 = ~n12989 & ~n12990 ;
  assign n12992 = n2041 & n12432 ;
  assign n12993 = \rf_conf1_reg[15]/NET0131  & ~n12974 ;
  assign n12994 = ~n12992 & ~n12993 ;
  assign n12995 = n2041 & n12459 ;
  assign n12996 = \rf_conf1_reg[1]/NET0131  & ~n12974 ;
  assign n12997 = ~n12995 & ~n12996 ;
  assign n12998 = n2041 & n12486 ;
  assign n12999 = \rf_conf1_reg[2]/NET0131  & ~n12974 ;
  assign n13000 = ~n12998 & ~n12999 ;
  assign n13001 = n2041 & n12513 ;
  assign n13002 = \rf_conf1_reg[3]/NET0131  & ~n12974 ;
  assign n13003 = ~n13001 & ~n13002 ;
  assign n13004 = n2041 & n12540 ;
  assign n13005 = \rf_conf1_reg[4]/NET0131  & ~n12974 ;
  assign n13006 = ~n13004 & ~n13005 ;
  assign n13007 = n2041 & n12567 ;
  assign n13008 = \rf_conf1_reg[5]/NET0131  & ~n12974 ;
  assign n13009 = ~n13007 & ~n13008 ;
  assign n13010 = n2041 & n12594 ;
  assign n13011 = \rf_conf1_reg[6]/NET0131  & ~n12974 ;
  assign n13012 = ~n13010 & ~n13011 ;
  assign n13013 = n2041 & n12621 ;
  assign n13014 = \rf_conf1_reg[7]/NET0131  & ~n12974 ;
  assign n13015 = ~n13013 & ~n13014 ;
  assign n13016 = n2041 & n12648 ;
  assign n13017 = \rf_conf1_reg[8]/NET0131  & ~n12974 ;
  assign n13018 = ~n13016 & ~n13017 ;
  assign n13019 = n2041 & n12675 ;
  assign n13020 = \rf_conf1_reg[9]/NET0131  & ~n12974 ;
  assign n13021 = ~n13019 & ~n13020 ;
  assign n13022 = n2039 & n12269 ;
  assign n13023 = \rf_rf_we_reg/P0001  & n2039 ;
  assign n13024 = \rf_conf2_reg[0]/NET0131  & ~n13023 ;
  assign n13025 = ~n13022 & ~n13024 ;
  assign n13026 = n2039 & n12297 ;
  assign n13027 = \rf_conf2_reg[10]/NET0131  & ~n13023 ;
  assign n13028 = ~n13026 & ~n13027 ;
  assign n13029 = n2039 & n12324 ;
  assign n13030 = \rf_conf2_reg[11]/NET0131  & ~n13023 ;
  assign n13031 = ~n13029 & ~n13030 ;
  assign n13032 = n2039 & n12351 ;
  assign n13033 = \rf_conf2_reg[12]/NET0131  & ~n13023 ;
  assign n13034 = ~n13032 & ~n13033 ;
  assign n13035 = n2039 & n12378 ;
  assign n13036 = \rf_conf2_reg[13]/NET0131  & ~n13023 ;
  assign n13037 = ~n13035 & ~n13036 ;
  assign n13038 = n2039 & n12405 ;
  assign n13039 = \rf_conf2_reg[14]/NET0131  & ~n13023 ;
  assign n13040 = ~n13038 & ~n13039 ;
  assign n13041 = n2039 & n12459 ;
  assign n13042 = \rf_conf2_reg[1]/NET0131  & ~n13023 ;
  assign n13043 = ~n13041 & ~n13042 ;
  assign n13044 = n2039 & n12432 ;
  assign n13045 = \rf_conf2_reg[15]/NET0131  & ~n13023 ;
  assign n13046 = ~n13044 & ~n13045 ;
  assign n13047 = n2039 & n12486 ;
  assign n13048 = \rf_conf2_reg[2]/NET0131  & ~n13023 ;
  assign n13049 = ~n13047 & ~n13048 ;
  assign n13050 = n2039 & n12513 ;
  assign n13051 = \rf_conf2_reg[3]/NET0131  & ~n13023 ;
  assign n13052 = ~n13050 & ~n13051 ;
  assign n13053 = n2039 & n12540 ;
  assign n13054 = \rf_conf2_reg[4]/NET0131  & ~n13023 ;
  assign n13055 = ~n13053 & ~n13054 ;
  assign n13056 = n2039 & n12567 ;
  assign n13057 = \rf_conf2_reg[5]/NET0131  & ~n13023 ;
  assign n13058 = ~n13056 & ~n13057 ;
  assign n13059 = n2039 & n12594 ;
  assign n13060 = \rf_conf2_reg[6]/NET0131  & ~n13023 ;
  assign n13061 = ~n13059 & ~n13060 ;
  assign n13062 = n2039 & n12621 ;
  assign n13063 = \rf_conf2_reg[7]/NET0131  & ~n13023 ;
  assign n13064 = ~n13062 & ~n13063 ;
  assign n13065 = n2039 & n12648 ;
  assign n13066 = \rf_conf2_reg[8]/NET0131  & ~n13023 ;
  assign n13067 = ~n13065 & ~n13066 ;
  assign n13068 = n2039 & n12675 ;
  assign n13069 = \rf_conf2_reg[9]/NET0131  & ~n13023 ;
  assign n13070 = ~n13068 & ~n13069 ;
  assign n13071 = n2027 & n12269 ;
  assign n13072 = \rf_rf_we_reg/P0001  & n2027 ;
  assign n13073 = \rf_conf3_reg[0]/NET0131  & ~n13072 ;
  assign n13074 = ~n13071 & ~n13073 ;
  assign n13075 = n2027 & n12297 ;
  assign n13076 = \rf_conf3_reg[10]/NET0131  & ~n13072 ;
  assign n13077 = ~n13075 & ~n13076 ;
  assign n13078 = n2027 & n12324 ;
  assign n13079 = \rf_conf3_reg[11]/NET0131  & ~n13072 ;
  assign n13080 = ~n13078 & ~n13079 ;
  assign n13081 = n2027 & n12351 ;
  assign n13082 = \rf_conf3_reg[12]/NET0131  & ~n13072 ;
  assign n13083 = ~n13081 & ~n13082 ;
  assign n13084 = n2027 & n12378 ;
  assign n13085 = \rf_conf3_reg[13]/NET0131  & ~n13072 ;
  assign n13086 = ~n13084 & ~n13085 ;
  assign n13087 = n2027 & n12405 ;
  assign n13088 = \rf_conf3_reg[14]/NET0131  & ~n13072 ;
  assign n13089 = ~n13087 & ~n13088 ;
  assign n13090 = n2027 & n12432 ;
  assign n13091 = \rf_conf3_reg[15]/NET0131  & ~n13072 ;
  assign n13092 = ~n13090 & ~n13091 ;
  assign n13093 = n2027 & n12459 ;
  assign n13094 = \rf_conf3_reg[1]/NET0131  & ~n13072 ;
  assign n13095 = ~n13093 & ~n13094 ;
  assign n13096 = n2027 & n12486 ;
  assign n13097 = \rf_conf3_reg[2]/NET0131  & ~n13072 ;
  assign n13098 = ~n13096 & ~n13097 ;
  assign n13099 = n2027 & n12540 ;
  assign n13100 = \rf_conf3_reg[4]/NET0131  & ~n13072 ;
  assign n13101 = ~n13099 & ~n13100 ;
  assign n13102 = n2027 & n12513 ;
  assign n13103 = \rf_conf3_reg[3]/NET0131  & ~n13072 ;
  assign n13104 = ~n13102 & ~n13103 ;
  assign n13105 = n2027 & n12567 ;
  assign n13106 = \rf_conf3_reg[5]/NET0131  & ~n13072 ;
  assign n13107 = ~n13105 & ~n13106 ;
  assign n13108 = n2027 & n12594 ;
  assign n13109 = \rf_conf3_reg[6]/NET0131  & ~n13072 ;
  assign n13110 = ~n13108 & ~n13109 ;
  assign n13111 = n2027 & n12621 ;
  assign n13112 = \rf_conf3_reg[7]/NET0131  & ~n13072 ;
  assign n13113 = ~n13111 & ~n13112 ;
  assign n13114 = n2027 & n12648 ;
  assign n13115 = \rf_conf3_reg[8]/NET0131  & ~n13072 ;
  assign n13116 = ~n13114 & ~n13115 ;
  assign n13117 = n2027 & n12675 ;
  assign n13118 = \rf_conf3_reg[9]/NET0131  & ~n13072 ;
  assign n13119 = ~n13117 & ~n13118 ;
  assign n13120 = n2046 & n12269 ;
  assign n13121 = \rf_rf_we_reg/P0001  & n2046 ;
  assign n13122 = \rf_conf4_reg[0]/NET0131  & ~n13121 ;
  assign n13123 = ~n13120 & ~n13122 ;
  assign n13124 = n2046 & n12297 ;
  assign n13125 = \rf_conf4_reg[10]/NET0131  & ~n13121 ;
  assign n13126 = ~n13124 & ~n13125 ;
  assign n13127 = n2046 & n12324 ;
  assign n13128 = \rf_conf4_reg[11]/NET0131  & ~n13121 ;
  assign n13129 = ~n13127 & ~n13128 ;
  assign n13130 = n2046 & n12351 ;
  assign n13131 = \rf_conf4_reg[12]/NET0131  & ~n13121 ;
  assign n13132 = ~n13130 & ~n13131 ;
  assign n13133 = n2046 & n12378 ;
  assign n13134 = \rf_conf4_reg[13]/NET0131  & ~n13121 ;
  assign n13135 = ~n13133 & ~n13134 ;
  assign n13136 = n2046 & n12405 ;
  assign n13137 = \rf_conf4_reg[14]/NET0131  & ~n13121 ;
  assign n13138 = ~n13136 & ~n13137 ;
  assign n13139 = n2046 & n12432 ;
  assign n13140 = \rf_conf4_reg[15]/NET0131  & ~n13121 ;
  assign n13141 = ~n13139 & ~n13140 ;
  assign n13142 = n2046 & n12459 ;
  assign n13143 = \rf_conf4_reg[1]/NET0131  & ~n13121 ;
  assign n13144 = ~n13142 & ~n13143 ;
  assign n13145 = n2046 & n12486 ;
  assign n13146 = \rf_conf4_reg[2]/NET0131  & ~n13121 ;
  assign n13147 = ~n13145 & ~n13146 ;
  assign n13148 = n2046 & n12513 ;
  assign n13149 = \rf_conf4_reg[3]/NET0131  & ~n13121 ;
  assign n13150 = ~n13148 & ~n13149 ;
  assign n13151 = n2046 & n12540 ;
  assign n13152 = \rf_conf4_reg[4]/NET0131  & ~n13121 ;
  assign n13153 = ~n13151 & ~n13152 ;
  assign n13154 = n2046 & n12567 ;
  assign n13155 = \rf_conf4_reg[5]/NET0131  & ~n13121 ;
  assign n13156 = ~n13154 & ~n13155 ;
  assign n13157 = n2046 & n12594 ;
  assign n13158 = \rf_conf4_reg[6]/NET0131  & ~n13121 ;
  assign n13159 = ~n13157 & ~n13158 ;
  assign n13160 = n2046 & n12621 ;
  assign n13161 = \rf_conf4_reg[7]/NET0131  & ~n13121 ;
  assign n13162 = ~n13160 & ~n13161 ;
  assign n13163 = n2046 & n12648 ;
  assign n13164 = \rf_conf4_reg[8]/NET0131  & ~n13121 ;
  assign n13165 = ~n13163 & ~n13164 ;
  assign n13166 = n2046 & n12675 ;
  assign n13167 = \rf_conf4_reg[9]/NET0131  & ~n13121 ;
  assign n13168 = ~n13166 & ~n13167 ;
  assign n13169 = n2023 & n12269 ;
  assign n13170 = \rf_rf_we_reg/P0001  & n2023 ;
  assign n13171 = \rf_conf5_reg[0]/NET0131  & ~n13170 ;
  assign n13172 = ~n13169 & ~n13171 ;
  assign n13173 = n2023 & n12297 ;
  assign n13174 = \rf_conf5_reg[10]/NET0131  & ~n13170 ;
  assign n13175 = ~n13173 & ~n13174 ;
  assign n13176 = n2023 & n12324 ;
  assign n13177 = \rf_conf5_reg[11]/NET0131  & ~n13170 ;
  assign n13178 = ~n13176 & ~n13177 ;
  assign n13179 = n2023 & n12351 ;
  assign n13180 = \rf_conf5_reg[12]/NET0131  & ~n13170 ;
  assign n13181 = ~n13179 & ~n13180 ;
  assign n13182 = n2023 & n12378 ;
  assign n13183 = \rf_conf5_reg[13]/NET0131  & ~n13170 ;
  assign n13184 = ~n13182 & ~n13183 ;
  assign n13185 = n2023 & n12405 ;
  assign n13186 = \rf_conf5_reg[14]/NET0131  & ~n13170 ;
  assign n13187 = ~n13185 & ~n13186 ;
  assign n13188 = n2023 & n12432 ;
  assign n13189 = \rf_conf5_reg[15]/NET0131  & ~n13170 ;
  assign n13190 = ~n13188 & ~n13189 ;
  assign n13191 = n2023 & n12459 ;
  assign n13192 = \rf_conf5_reg[1]/NET0131  & ~n13170 ;
  assign n13193 = ~n13191 & ~n13192 ;
  assign n13194 = n2023 & n12513 ;
  assign n13195 = \rf_conf5_reg[3]/NET0131  & ~n13170 ;
  assign n13196 = ~n13194 & ~n13195 ;
  assign n13197 = n2023 & n12486 ;
  assign n13198 = \rf_conf5_reg[2]/NET0131  & ~n13170 ;
  assign n13199 = ~n13197 & ~n13198 ;
  assign n13200 = n2023 & n12540 ;
  assign n13201 = \rf_conf5_reg[4]/NET0131  & ~n13170 ;
  assign n13202 = ~n13200 & ~n13201 ;
  assign n13203 = n2023 & n12567 ;
  assign n13204 = \rf_conf5_reg[5]/NET0131  & ~n13170 ;
  assign n13205 = ~n13203 & ~n13204 ;
  assign n13206 = n2023 & n12594 ;
  assign n13207 = \rf_conf5_reg[6]/NET0131  & ~n13170 ;
  assign n13208 = ~n13206 & ~n13207 ;
  assign n13209 = n2023 & n12621 ;
  assign n13210 = \rf_conf5_reg[7]/NET0131  & ~n13170 ;
  assign n13211 = ~n13209 & ~n13210 ;
  assign n13212 = n2023 & n12648 ;
  assign n13213 = \rf_conf5_reg[8]/NET0131  & ~n13170 ;
  assign n13214 = ~n13212 & ~n13213 ;
  assign n13215 = n2023 & n12675 ;
  assign n13216 = \rf_conf5_reg[9]/NET0131  & ~n13170 ;
  assign n13217 = ~n13215 & ~n13216 ;
  assign n13218 = n2051 & n12269 ;
  assign n13219 = \rf_rf_we_reg/P0001  & n2051 ;
  assign n13220 = \rf_conf6_reg[0]/NET0131  & ~n13219 ;
  assign n13221 = ~n13218 & ~n13220 ;
  assign n13222 = n2051 & n12297 ;
  assign n13223 = \rf_conf6_reg[10]/NET0131  & ~n13219 ;
  assign n13224 = ~n13222 & ~n13223 ;
  assign n13225 = n2051 & n12324 ;
  assign n13226 = \rf_conf6_reg[11]/NET0131  & ~n13219 ;
  assign n13227 = ~n13225 & ~n13226 ;
  assign n13228 = n2051 & n12351 ;
  assign n13229 = \rf_conf6_reg[12]/NET0131  & ~n13219 ;
  assign n13230 = ~n13228 & ~n13229 ;
  assign n13231 = n2051 & n12378 ;
  assign n13232 = \rf_conf6_reg[13]/NET0131  & ~n13219 ;
  assign n13233 = ~n13231 & ~n13232 ;
  assign n13234 = n2051 & n12405 ;
  assign n13235 = \rf_conf6_reg[14]/NET0131  & ~n13219 ;
  assign n13236 = ~n13234 & ~n13235 ;
  assign n13237 = n2051 & n12432 ;
  assign n13238 = \rf_conf6_reg[15]/NET0131  & ~n13219 ;
  assign n13239 = ~n13237 & ~n13238 ;
  assign n13240 = n2051 & n12459 ;
  assign n13241 = \rf_conf6_reg[1]/NET0131  & ~n13219 ;
  assign n13242 = ~n13240 & ~n13241 ;
  assign n13243 = n2051 & n12486 ;
  assign n13244 = \rf_conf6_reg[2]/NET0131  & ~n13219 ;
  assign n13245 = ~n13243 & ~n13244 ;
  assign n13246 = n2051 & n12513 ;
  assign n13247 = \rf_conf6_reg[3]/NET0131  & ~n13219 ;
  assign n13248 = ~n13246 & ~n13247 ;
  assign n13249 = n2051 & n12540 ;
  assign n13250 = \rf_conf6_reg[4]/NET0131  & ~n13219 ;
  assign n13251 = ~n13249 & ~n13250 ;
  assign n13252 = n2051 & n12567 ;
  assign n13253 = \rf_conf6_reg[5]/NET0131  & ~n13219 ;
  assign n13254 = ~n13252 & ~n13253 ;
  assign n13255 = n2051 & n12594 ;
  assign n13256 = \rf_conf6_reg[6]/NET0131  & ~n13219 ;
  assign n13257 = ~n13255 & ~n13256 ;
  assign n13258 = n2051 & n12621 ;
  assign n13259 = \rf_conf6_reg[7]/NET0131  & ~n13219 ;
  assign n13260 = ~n13258 & ~n13259 ;
  assign n13261 = n2051 & n12648 ;
  assign n13262 = \rf_conf6_reg[8]/NET0131  & ~n13219 ;
  assign n13263 = ~n13261 & ~n13262 ;
  assign n13264 = n2051 & n12675 ;
  assign n13265 = \rf_conf6_reg[9]/NET0131  & ~n13219 ;
  assign n13266 = ~n13264 & ~n13265 ;
  assign n13267 = n2053 & n12269 ;
  assign n13268 = \rf_rf_we_reg/P0001  & n2053 ;
  assign n13269 = \rf_conf7_reg[0]/NET0131  & ~n13268 ;
  assign n13270 = ~n13267 & ~n13269 ;
  assign n13271 = n2053 & n12324 ;
  assign n13272 = \rf_conf7_reg[11]/NET0131  & ~n13268 ;
  assign n13273 = ~n13271 & ~n13272 ;
  assign n13274 = n2053 & n12297 ;
  assign n13275 = \rf_conf7_reg[10]/NET0131  & ~n13268 ;
  assign n13276 = ~n13274 & ~n13275 ;
  assign n13277 = n2053 & n12351 ;
  assign n13278 = \rf_conf7_reg[12]/NET0131  & ~n13268 ;
  assign n13279 = ~n13277 & ~n13278 ;
  assign n13280 = n2053 & n12378 ;
  assign n13281 = \rf_conf7_reg[13]/NET0131  & ~n13268 ;
  assign n13282 = ~n13280 & ~n13281 ;
  assign n13283 = n2053 & n12405 ;
  assign n13284 = \rf_conf7_reg[14]/NET0131  & ~n13268 ;
  assign n13285 = ~n13283 & ~n13284 ;
  assign n13286 = n2053 & n12432 ;
  assign n13287 = \rf_conf7_reg[15]/NET0131  & ~n13268 ;
  assign n13288 = ~n13286 & ~n13287 ;
  assign n13289 = n2053 & n12459 ;
  assign n13290 = \rf_conf7_reg[1]/NET0131  & ~n13268 ;
  assign n13291 = ~n13289 & ~n13290 ;
  assign n13292 = n2053 & n12486 ;
  assign n13293 = \rf_conf7_reg[2]/NET0131  & ~n13268 ;
  assign n13294 = ~n13292 & ~n13293 ;
  assign n13295 = n2053 & n12513 ;
  assign n13296 = \rf_conf7_reg[3]/NET0131  & ~n13268 ;
  assign n13297 = ~n13295 & ~n13296 ;
  assign n13298 = n2053 & n12540 ;
  assign n13299 = \rf_conf7_reg[4]/NET0131  & ~n13268 ;
  assign n13300 = ~n13298 & ~n13299 ;
  assign n13301 = n2053 & n12567 ;
  assign n13302 = \rf_conf7_reg[5]/NET0131  & ~n13268 ;
  assign n13303 = ~n13301 & ~n13302 ;
  assign n13304 = n2053 & n12594 ;
  assign n13305 = \rf_conf7_reg[6]/NET0131  & ~n13268 ;
  assign n13306 = ~n13304 & ~n13305 ;
  assign n13307 = n2053 & n12621 ;
  assign n13308 = \rf_conf7_reg[7]/NET0131  & ~n13268 ;
  assign n13309 = ~n13307 & ~n13308 ;
  assign n13310 = n2053 & n12648 ;
  assign n13311 = \rf_conf7_reg[8]/NET0131  & ~n13268 ;
  assign n13312 = ~n13310 & ~n13311 ;
  assign n13313 = n2053 & n12675 ;
  assign n13314 = \rf_conf7_reg[9]/NET0131  & ~n13268 ;
  assign n13315 = ~n13313 & ~n13314 ;
  assign n13316 = n2057 & n12269 ;
  assign n13317 = \rf_rf_we_reg/P0001  & n2057 ;
  assign n13318 = \rf_conf8_reg[0]/NET0131  & ~n13317 ;
  assign n13319 = ~n13316 & ~n13318 ;
  assign n13320 = n2057 & n12297 ;
  assign n13321 = \rf_conf8_reg[10]/NET0131  & ~n13317 ;
  assign n13322 = ~n13320 & ~n13321 ;
  assign n13323 = n2057 & n12324 ;
  assign n13324 = \rf_conf8_reg[11]/NET0131  & ~n13317 ;
  assign n13325 = ~n13323 & ~n13324 ;
  assign n13326 = n2057 & n12351 ;
  assign n13327 = \rf_conf8_reg[12]/NET0131  & ~n13317 ;
  assign n13328 = ~n13326 & ~n13327 ;
  assign n13329 = n2057 & n12378 ;
  assign n13330 = \rf_conf8_reg[13]/NET0131  & ~n13317 ;
  assign n13331 = ~n13329 & ~n13330 ;
  assign n13332 = n2057 & n12405 ;
  assign n13333 = \rf_conf8_reg[14]/NET0131  & ~n13317 ;
  assign n13334 = ~n13332 & ~n13333 ;
  assign n13335 = n2057 & n12432 ;
  assign n13336 = \rf_conf8_reg[15]/NET0131  & ~n13317 ;
  assign n13337 = ~n13335 & ~n13336 ;
  assign n13338 = n2057 & n12459 ;
  assign n13339 = \rf_conf8_reg[1]/NET0131  & ~n13317 ;
  assign n13340 = ~n13338 & ~n13339 ;
  assign n13341 = n2057 & n12486 ;
  assign n13342 = \rf_conf8_reg[2]/NET0131  & ~n13317 ;
  assign n13343 = ~n13341 & ~n13342 ;
  assign n13344 = n2057 & n12513 ;
  assign n13345 = \rf_conf8_reg[3]/NET0131  & ~n13317 ;
  assign n13346 = ~n13344 & ~n13345 ;
  assign n13347 = n2057 & n12567 ;
  assign n13348 = \rf_conf8_reg[5]/NET0131  & ~n13317 ;
  assign n13349 = ~n13347 & ~n13348 ;
  assign n13350 = n2057 & n12540 ;
  assign n13351 = \rf_conf8_reg[4]/NET0131  & ~n13317 ;
  assign n13352 = ~n13350 & ~n13351 ;
  assign n13353 = n2057 & n12594 ;
  assign n13354 = \rf_conf8_reg[6]/NET0131  & ~n13317 ;
  assign n13355 = ~n13353 & ~n13354 ;
  assign n13356 = n2057 & n12621 ;
  assign n13357 = \rf_conf8_reg[7]/NET0131  & ~n13317 ;
  assign n13358 = ~n13356 & ~n13357 ;
  assign n13359 = n2057 & n12648 ;
  assign n13360 = \rf_conf8_reg[8]/NET0131  & ~n13317 ;
  assign n13361 = ~n13359 & ~n13360 ;
  assign n13362 = n2057 & n12675 ;
  assign n13363 = \rf_conf8_reg[9]/NET0131  & ~n13317 ;
  assign n13364 = ~n13362 & ~n13363 ;
  assign n13365 = n2063 & n12269 ;
  assign n13366 = \rf_rf_we_reg/P0001  & n2063 ;
  assign n13367 = \rf_conf9_reg[0]/NET0131  & ~n13366 ;
  assign n13368 = ~n13365 & ~n13367 ;
  assign n13369 = n2063 & n12297 ;
  assign n13370 = \rf_conf9_reg[10]/NET0131  & ~n13366 ;
  assign n13371 = ~n13369 & ~n13370 ;
  assign n13372 = n2063 & n12324 ;
  assign n13373 = \rf_conf9_reg[11]/NET0131  & ~n13366 ;
  assign n13374 = ~n13372 & ~n13373 ;
  assign n13375 = n2063 & n12351 ;
  assign n13376 = \rf_conf9_reg[12]/NET0131  & ~n13366 ;
  assign n13377 = ~n13375 & ~n13376 ;
  assign n13378 = n2063 & n12378 ;
  assign n13379 = \rf_conf9_reg[13]/NET0131  & ~n13366 ;
  assign n13380 = ~n13378 & ~n13379 ;
  assign n13381 = n2063 & n12405 ;
  assign n13382 = \rf_conf9_reg[14]/NET0131  & ~n13366 ;
  assign n13383 = ~n13381 & ~n13382 ;
  assign n13384 = n2063 & n12432 ;
  assign n13385 = \rf_conf9_reg[15]/NET0131  & ~n13366 ;
  assign n13386 = ~n13384 & ~n13385 ;
  assign n13387 = n2063 & n12459 ;
  assign n13388 = \rf_conf9_reg[1]/NET0131  & ~n13366 ;
  assign n13389 = ~n13387 & ~n13388 ;
  assign n13390 = n2063 & n12486 ;
  assign n13391 = \rf_conf9_reg[2]/NET0131  & ~n13366 ;
  assign n13392 = ~n13390 & ~n13391 ;
  assign n13393 = n2063 & n12513 ;
  assign n13394 = \rf_conf9_reg[3]/NET0131  & ~n13366 ;
  assign n13395 = ~n13393 & ~n13394 ;
  assign n13396 = n2063 & n12540 ;
  assign n13397 = \rf_conf9_reg[4]/NET0131  & ~n13366 ;
  assign n13398 = ~n13396 & ~n13397 ;
  assign n13399 = n2063 & n12567 ;
  assign n13400 = \rf_conf9_reg[5]/NET0131  & ~n13366 ;
  assign n13401 = ~n13399 & ~n13400 ;
  assign n13402 = n2063 & n12594 ;
  assign n13403 = \rf_conf9_reg[6]/NET0131  & ~n13366 ;
  assign n13404 = ~n13402 & ~n13403 ;
  assign n13405 = n2063 & n12621 ;
  assign n13406 = \rf_conf9_reg[7]/NET0131  & ~n13366 ;
  assign n13407 = ~n13405 & ~n13406 ;
  assign n13408 = n2063 & n12648 ;
  assign n13409 = \rf_conf9_reg[8]/NET0131  & ~n13366 ;
  assign n13410 = ~n13408 & ~n13409 ;
  assign n13411 = n2063 & n12675 ;
  assign n13412 = \rf_conf9_reg[9]/NET0131  & ~n13366 ;
  assign n13413 = ~n13411 & ~n13412 ;
  assign n13414 = ~\rf_rf_ack_reg/P0001  & ~n2106 ;
  assign n13415 = n2153 & n13414 ;
  assign n13416 = n2257 & n13415 ;
  assign n13417 = \m7_we_i_pad  & ~n1910 ;
  assign n13418 = n1938 & n13417 ;
  assign n13419 = \m6_we_i_pad  & ~n1925 ;
  assign n13420 = n1918 & n13419 ;
  assign n13421 = ~n13418 & ~n13420 ;
  assign n13422 = \m5_we_i_pad  & ~n1910 ;
  assign n13423 = n1941 & n13422 ;
  assign n13424 = \m2_we_i_pad  & ~n1925 ;
  assign n13425 = n1931 & n13424 ;
  assign n13426 = ~n13423 & ~n13425 ;
  assign n13427 = n13421 & n13426 ;
  assign n13428 = \m4_we_i_pad  & n1925 ;
  assign n13429 = n1918 & n13428 ;
  assign n13430 = \m3_we_i_pad  & n1910 ;
  assign n13431 = n1938 & n13430 ;
  assign n13432 = ~n13429 & ~n13431 ;
  assign n13433 = \m1_we_i_pad  & n1910 ;
  assign n13434 = n1941 & n13433 ;
  assign n13435 = \m0_we_i_pad  & n1925 ;
  assign n13436 = n1931 & n13435 ;
  assign n13437 = ~n13434 & ~n13436 ;
  assign n13438 = n13432 & n13437 ;
  assign n13439 = n13427 & n13438 ;
  assign n13440 = ~\rf_rf_we_reg/P0001  & ~n13439 ;
  assign n13441 = n2258 & n13440 ;
  assign n13442 = ~\s4_msel_pri_out_reg[0]/NET0131  & \s4_msel_pri_out_reg[1]/NET0131  ;
  assign n13443 = \s4_msel_arb2_state_reg[1]/NET0131  & n13442 ;
  assign n13444 = \s4_msel_pri_out_reg[0]/NET0131  & ~\s4_msel_pri_out_reg[1]/NET0131  ;
  assign n13445 = \s4_msel_arb1_state_reg[1]/NET0131  & n13444 ;
  assign n13446 = ~n13443 & ~n13445 ;
  assign n13447 = \s4_msel_pri_out_reg[0]/NET0131  & \s4_msel_pri_out_reg[1]/NET0131  ;
  assign n13448 = \s4_msel_arb3_state_reg[1]/NET0131  & n13447 ;
  assign n13449 = ~\s4_msel_pri_out_reg[0]/NET0131  & ~\s4_msel_pri_out_reg[1]/NET0131  ;
  assign n13450 = \s4_msel_arb0_state_reg[1]/NET0131  & n13449 ;
  assign n13451 = ~n13448 & ~n13450 ;
  assign n13452 = n13446 & n13451 ;
  assign n13453 = \s4_msel_arb0_state_reg[2]/NET0131  & n13449 ;
  assign n13454 = \s4_msel_arb3_state_reg[2]/NET0131  & n13447 ;
  assign n13455 = ~n13453 & ~n13454 ;
  assign n13456 = \s4_msel_arb1_state_reg[2]/NET0131  & n13444 ;
  assign n13457 = \s4_msel_arb2_state_reg[2]/NET0131  & n13442 ;
  assign n13458 = ~n13456 & ~n13457 ;
  assign n13459 = n13455 & n13458 ;
  assign n13460 = n13452 & ~n13459 ;
  assign n13461 = \s4_msel_arb2_state_reg[0]/NET0131  & n13442 ;
  assign n13462 = \s4_msel_arb1_state_reg[0]/NET0131  & n13444 ;
  assign n13463 = ~n13461 & ~n13462 ;
  assign n13464 = \s4_msel_arb3_state_reg[0]/NET0131  & n13447 ;
  assign n13465 = \s4_msel_arb0_state_reg[0]/NET0131  & n13449 ;
  assign n13466 = ~n13464 & ~n13465 ;
  assign n13467 = n13463 & n13466 ;
  assign n13468 = \m5_s4_cyc_o_reg/NET0131  & \s4_m5_cyc_r_reg/P0001  ;
  assign n13469 = ~n13467 & n13468 ;
  assign n13470 = n13460 & n13469 ;
  assign n13471 = \m4_s4_cyc_o_reg/NET0131  & \s4_m4_cyc_r_reg/P0001  ;
  assign n13472 = n13467 & n13471 ;
  assign n13473 = n13460 & n13472 ;
  assign n13474 = ~n13470 & ~n13473 ;
  assign n13475 = n13452 & n13459 ;
  assign n13476 = \m1_s4_cyc_o_reg/NET0131  & \s4_m1_cyc_r_reg/P0001  ;
  assign n13477 = ~n13467 & n13476 ;
  assign n13478 = n13475 & n13477 ;
  assign n13479 = \m0_s4_cyc_o_reg/NET0131  & \s4_m0_cyc_r_reg/P0001  ;
  assign n13480 = n13467 & n13479 ;
  assign n13481 = n13475 & n13480 ;
  assign n13482 = ~n13478 & ~n13481 ;
  assign n13483 = n13474 & n13482 ;
  assign n13484 = ~n13452 & n13459 ;
  assign n13485 = \m3_s4_cyc_o_reg/NET0131  & \s4_m3_cyc_r_reg/P0001  ;
  assign n13486 = ~n13467 & n13485 ;
  assign n13487 = n13484 & n13486 ;
  assign n13488 = \m2_s4_cyc_o_reg/NET0131  & \s4_m2_cyc_r_reg/P0001  ;
  assign n13489 = n13467 & n13488 ;
  assign n13490 = n13484 & n13489 ;
  assign n13491 = ~n13487 & ~n13490 ;
  assign n13492 = ~n13452 & ~n13459 ;
  assign n13493 = \m7_s4_cyc_o_reg/NET0131  & \s4_m7_cyc_r_reg/P0001  ;
  assign n13494 = ~n13467 & n13493 ;
  assign n13495 = n13492 & n13494 ;
  assign n13496 = \m6_s4_cyc_o_reg/NET0131  & \s4_m6_cyc_r_reg/P0001  ;
  assign n13497 = n13467 & n13496 ;
  assign n13498 = n13492 & n13497 ;
  assign n13499 = ~n13495 & ~n13498 ;
  assign n13500 = n13491 & n13499 ;
  assign n13501 = n13483 & n13500 ;
  assign n13502 = n4889 & n4904 ;
  assign n13503 = \s10_next_reg/P0001  & n9814 ;
  assign n13504 = n9824 & n13503 ;
  assign n13505 = ~n13502 & n13504 ;
  assign n13506 = \s10_msel_pri_out_reg[0]/NET0131  & ~\s10_next_reg/P0001  ;
  assign n13507 = n4220 & n4225 ;
  assign n13508 = \s10_next_reg/P0001  & ~n13507 ;
  assign n13509 = ~n13506 & ~n13508 ;
  assign n13510 = ~n13505 & n13509 ;
  assign n13511 = ~rst_i_pad & ~n13510 ;
  assign n13512 = n4920 & n4944 ;
  assign n13513 = \s11_next_reg/P0001  & n4253 ;
  assign n13514 = n4270 & n13513 ;
  assign n13515 = ~n13512 & n13514 ;
  assign n13516 = \s11_msel_pri_out_reg[0]/NET0131  & ~\s11_next_reg/P0001  ;
  assign n13517 = n4293 & n4310 ;
  assign n13518 = \s11_next_reg/P0001  & ~n13517 ;
  assign n13519 = ~n13516 & ~n13518 ;
  assign n13520 = ~n13515 & n13519 ;
  assign n13521 = ~rst_i_pad & ~n13520 ;
  assign n13522 = ~\s5_msel_pri_out_reg[0]/NET0131  & \s5_msel_pri_out_reg[1]/NET0131  ;
  assign n13523 = \s5_msel_arb2_state_reg[1]/NET0131  & n13522 ;
  assign n13524 = \s5_msel_pri_out_reg[0]/NET0131  & ~\s5_msel_pri_out_reg[1]/NET0131  ;
  assign n13525 = \s5_msel_arb1_state_reg[1]/NET0131  & n13524 ;
  assign n13526 = ~n13523 & ~n13525 ;
  assign n13527 = \s5_msel_pri_out_reg[0]/NET0131  & \s5_msel_pri_out_reg[1]/NET0131  ;
  assign n13528 = \s5_msel_arb3_state_reg[1]/NET0131  & n13527 ;
  assign n13529 = ~\s5_msel_pri_out_reg[0]/NET0131  & ~\s5_msel_pri_out_reg[1]/NET0131  ;
  assign n13530 = \s5_msel_arb0_state_reg[1]/NET0131  & n13529 ;
  assign n13531 = ~n13528 & ~n13530 ;
  assign n13532 = n13526 & n13531 ;
  assign n13533 = \s5_msel_arb2_state_reg[2]/NET0131  & n13522 ;
  assign n13534 = \s5_msel_arb1_state_reg[2]/NET0131  & n13524 ;
  assign n13535 = ~n13533 & ~n13534 ;
  assign n13536 = \s5_msel_arb3_state_reg[2]/NET0131  & n13527 ;
  assign n13537 = \s5_msel_arb0_state_reg[2]/NET0131  & n13529 ;
  assign n13538 = ~n13536 & ~n13537 ;
  assign n13539 = n13535 & n13538 ;
  assign n13540 = ~n13532 & n13539 ;
  assign n13541 = \s5_msel_arb2_state_reg[0]/NET0131  & n13522 ;
  assign n13542 = \s5_msel_arb1_state_reg[0]/NET0131  & n13524 ;
  assign n13543 = ~n13541 & ~n13542 ;
  assign n13544 = \s5_msel_arb3_state_reg[0]/NET0131  & n13527 ;
  assign n13545 = \s5_msel_arb0_state_reg[0]/NET0131  & n13529 ;
  assign n13546 = ~n13544 & ~n13545 ;
  assign n13547 = n13543 & n13546 ;
  assign n13548 = \m3_s5_cyc_o_reg/NET0131  & \s5_m3_cyc_r_reg/P0001  ;
  assign n13549 = ~n13547 & n13548 ;
  assign n13550 = n13540 & n13549 ;
  assign n13551 = \m2_s5_cyc_o_reg/NET0131  & \s5_m2_cyc_r_reg/P0001  ;
  assign n13552 = n13547 & n13551 ;
  assign n13553 = n13540 & n13552 ;
  assign n13554 = ~n13550 & ~n13553 ;
  assign n13555 = n13532 & ~n13539 ;
  assign n13556 = \m5_s5_cyc_o_reg/NET0131  & \s5_m5_cyc_r_reg/P0001  ;
  assign n13557 = ~n13547 & n13556 ;
  assign n13558 = n13555 & n13557 ;
  assign n13559 = \m4_s5_cyc_o_reg/NET0131  & \s5_m4_cyc_r_reg/P0001  ;
  assign n13560 = n13547 & n13559 ;
  assign n13561 = n13555 & n13560 ;
  assign n13562 = ~n13558 & ~n13561 ;
  assign n13563 = n13554 & n13562 ;
  assign n13564 = ~n13532 & ~n13539 ;
  assign n13565 = \m7_s5_cyc_o_reg/NET0131  & \s5_m7_cyc_r_reg/P0001  ;
  assign n13566 = ~n13547 & n13565 ;
  assign n13567 = n13564 & n13566 ;
  assign n13568 = \m6_s5_cyc_o_reg/NET0131  & \s5_m6_cyc_r_reg/P0001  ;
  assign n13569 = n13547 & n13568 ;
  assign n13570 = n13564 & n13569 ;
  assign n13571 = ~n13567 & ~n13570 ;
  assign n13572 = n13532 & n13539 ;
  assign n13573 = \m1_s5_cyc_o_reg/NET0131  & \s5_m1_cyc_r_reg/P0001  ;
  assign n13574 = ~n13547 & n13573 ;
  assign n13575 = n13572 & n13574 ;
  assign n13576 = \m0_s5_cyc_o_reg/NET0131  & \s5_m0_cyc_r_reg/P0001  ;
  assign n13577 = n13547 & n13576 ;
  assign n13578 = n13572 & n13577 ;
  assign n13579 = ~n13575 & ~n13578 ;
  assign n13580 = n13571 & n13579 ;
  assign n13581 = n13563 & n13580 ;
  assign n13582 = n4974 & n4995 ;
  assign n13583 = \s12_next_reg/P0001  & n9849 ;
  assign n13584 = n9859 & n13583 ;
  assign n13585 = ~n13582 & n13584 ;
  assign n13586 = \s12_msel_pri_out_reg[0]/NET0131  & ~\s12_next_reg/P0001  ;
  assign n13587 = n4360 & n4365 ;
  assign n13588 = \s12_next_reg/P0001  & ~n13587 ;
  assign n13589 = ~n13586 & ~n13588 ;
  assign n13590 = ~n13585 & n13589 ;
  assign n13591 = ~rst_i_pad & ~n13590 ;
  assign n13592 = n5011 & n5026 ;
  assign n13593 = \s13_next_reg/P0001  & n9877 ;
  assign n13594 = n9894 & n13593 ;
  assign n13595 = ~n13592 & n13594 ;
  assign n13596 = \s13_msel_pri_out_reg[0]/NET0131  & ~\s13_next_reg/P0001  ;
  assign n13597 = n3875 & n3880 ;
  assign n13598 = \s13_next_reg/P0001  & ~n13597 ;
  assign n13599 = ~n13596 & ~n13598 ;
  assign n13600 = ~n13595 & n13599 ;
  assign n13601 = ~rst_i_pad & ~n13600 ;
  assign n13602 = ~\s6_msel_pri_out_reg[0]/NET0131  & ~\s6_msel_pri_out_reg[1]/NET0131  ;
  assign n13603 = \s6_msel_arb0_state_reg[1]/NET0131  & n13602 ;
  assign n13604 = \s6_msel_pri_out_reg[0]/NET0131  & \s6_msel_pri_out_reg[1]/NET0131  ;
  assign n13605 = \s6_msel_arb3_state_reg[1]/NET0131  & n13604 ;
  assign n13606 = ~n13603 & ~n13605 ;
  assign n13607 = ~\s6_msel_pri_out_reg[0]/NET0131  & \s6_msel_pri_out_reg[1]/NET0131  ;
  assign n13608 = \s6_msel_arb2_state_reg[1]/NET0131  & n13607 ;
  assign n13609 = \s6_msel_pri_out_reg[0]/NET0131  & ~\s6_msel_pri_out_reg[1]/NET0131  ;
  assign n13610 = \s6_msel_arb1_state_reg[1]/NET0131  & n13609 ;
  assign n13611 = ~n13608 & ~n13610 ;
  assign n13612 = n13606 & n13611 ;
  assign n13613 = \s6_msel_arb0_state_reg[2]/NET0131  & n13602 ;
  assign n13614 = \s6_msel_arb3_state_reg[2]/NET0131  & n13604 ;
  assign n13615 = ~n13613 & ~n13614 ;
  assign n13616 = \s6_msel_arb1_state_reg[2]/NET0131  & n13609 ;
  assign n13617 = \s6_msel_arb2_state_reg[2]/NET0131  & n13607 ;
  assign n13618 = ~n13616 & ~n13617 ;
  assign n13619 = n13615 & n13618 ;
  assign n13620 = n13612 & n13619 ;
  assign n13621 = \s6_msel_arb0_state_reg[0]/NET0131  & n13602 ;
  assign n13622 = \s6_msel_arb2_state_reg[0]/NET0131  & n13607 ;
  assign n13623 = ~n13621 & ~n13622 ;
  assign n13624 = \s6_msel_arb3_state_reg[0]/NET0131  & n13604 ;
  assign n13625 = \s6_msel_arb1_state_reg[0]/NET0131  & n13609 ;
  assign n13626 = ~n13624 & ~n13625 ;
  assign n13627 = n13623 & n13626 ;
  assign n13628 = \m1_s6_cyc_o_reg/NET0131  & \s6_m1_cyc_r_reg/P0001  ;
  assign n13629 = ~n13627 & n13628 ;
  assign n13630 = n13620 & n13629 ;
  assign n13631 = \m0_s6_cyc_o_reg/NET0131  & \s6_m0_cyc_r_reg/P0001  ;
  assign n13632 = n13627 & n13631 ;
  assign n13633 = n13620 & n13632 ;
  assign n13634 = ~n13630 & ~n13633 ;
  assign n13635 = ~n13612 & n13619 ;
  assign n13636 = \m3_s6_cyc_o_reg/NET0131  & \s6_m3_cyc_r_reg/P0001  ;
  assign n13637 = ~n13627 & n13636 ;
  assign n13638 = n13635 & n13637 ;
  assign n13639 = \m2_s6_cyc_o_reg/NET0131  & \s6_m2_cyc_r_reg/P0001  ;
  assign n13640 = n13627 & n13639 ;
  assign n13641 = n13635 & n13640 ;
  assign n13642 = ~n13638 & ~n13641 ;
  assign n13643 = n13634 & n13642 ;
  assign n13644 = ~n13612 & ~n13619 ;
  assign n13645 = \m7_s6_cyc_o_reg/NET0131  & \s6_m7_cyc_r_reg/P0001  ;
  assign n13646 = ~n13627 & n13645 ;
  assign n13647 = n13644 & n13646 ;
  assign n13648 = \m6_s6_cyc_o_reg/NET0131  & \s6_m6_cyc_r_reg/P0001  ;
  assign n13649 = n13627 & n13648 ;
  assign n13650 = n13644 & n13649 ;
  assign n13651 = ~n13647 & ~n13650 ;
  assign n13652 = n13612 & ~n13619 ;
  assign n13653 = \m5_s6_cyc_o_reg/NET0131  & \s6_m5_cyc_r_reg/P0001  ;
  assign n13654 = ~n13627 & n13653 ;
  assign n13655 = n13652 & n13654 ;
  assign n13656 = \m4_s6_cyc_o_reg/NET0131  & \s6_m4_cyc_r_reg/P0001  ;
  assign n13657 = n13627 & n13656 ;
  assign n13658 = n13652 & n13657 ;
  assign n13659 = ~n13655 & ~n13658 ;
  assign n13660 = n13651 & n13659 ;
  assign n13661 = n13643 & n13660 ;
  assign n13662 = n5039 & n5061 ;
  assign n13663 = \s14_next_reg/P0001  & n3926 ;
  assign n13664 = n3921 & n13663 ;
  assign n13665 = ~n13662 & n13664 ;
  assign n13666 = \s14_msel_pri_out_reg[0]/NET0131  & ~\s14_next_reg/P0001  ;
  assign n13667 = n4398 & n4415 ;
  assign n13668 = \s14_next_reg/P0001  & ~n13667 ;
  assign n13669 = ~n13666 & ~n13668 ;
  assign n13670 = ~n13665 & n13669 ;
  assign n13671 = ~rst_i_pad & ~n13670 ;
  assign n13672 = ~\s7_msel_pri_out_reg[0]/NET0131  & ~\s7_msel_pri_out_reg[1]/NET0131  ;
  assign n13673 = \s7_msel_arb0_state_reg[1]/NET0131  & n13672 ;
  assign n13674 = \s7_msel_pri_out_reg[0]/NET0131  & \s7_msel_pri_out_reg[1]/NET0131  ;
  assign n13675 = \s7_msel_arb3_state_reg[1]/NET0131  & n13674 ;
  assign n13676 = ~n13673 & ~n13675 ;
  assign n13677 = \s7_msel_pri_out_reg[0]/NET0131  & ~\s7_msel_pri_out_reg[1]/NET0131  ;
  assign n13678 = \s7_msel_arb1_state_reg[1]/NET0131  & n13677 ;
  assign n13679 = ~\s7_msel_pri_out_reg[0]/NET0131  & \s7_msel_pri_out_reg[1]/NET0131  ;
  assign n13680 = \s7_msel_arb2_state_reg[1]/NET0131  & n13679 ;
  assign n13681 = ~n13678 & ~n13680 ;
  assign n13682 = n13676 & n13681 ;
  assign n13683 = \s7_msel_arb2_state_reg[2]/NET0131  & n13679 ;
  assign n13684 = \s7_msel_arb1_state_reg[2]/NET0131  & n13677 ;
  assign n13685 = ~n13683 & ~n13684 ;
  assign n13686 = \s7_msel_arb3_state_reg[2]/NET0131  & n13674 ;
  assign n13687 = \s7_msel_arb0_state_reg[2]/NET0131  & n13672 ;
  assign n13688 = ~n13686 & ~n13687 ;
  assign n13689 = n13685 & n13688 ;
  assign n13690 = ~n13682 & ~n13689 ;
  assign n13691 = \s7_msel_arb2_state_reg[0]/NET0131  & n13679 ;
  assign n13692 = \s7_msel_arb1_state_reg[0]/NET0131  & n13677 ;
  assign n13693 = ~n13691 & ~n13692 ;
  assign n13694 = \s7_msel_arb3_state_reg[0]/NET0131  & n13674 ;
  assign n13695 = \s7_msel_arb0_state_reg[0]/NET0131  & n13672 ;
  assign n13696 = ~n13694 & ~n13695 ;
  assign n13697 = n13693 & n13696 ;
  assign n13698 = \m7_s7_cyc_o_reg/NET0131  & \s7_m7_cyc_r_reg/P0001  ;
  assign n13699 = ~n13697 & n13698 ;
  assign n13700 = n13690 & n13699 ;
  assign n13701 = \m6_s7_cyc_o_reg/NET0131  & \s7_m6_cyc_r_reg/P0001  ;
  assign n13702 = n13697 & n13701 ;
  assign n13703 = n13690 & n13702 ;
  assign n13704 = ~n13700 & ~n13703 ;
  assign n13705 = n13682 & n13689 ;
  assign n13706 = \m1_s7_cyc_o_reg/NET0131  & \s7_m1_cyc_r_reg/P0001  ;
  assign n13707 = ~n13697 & n13706 ;
  assign n13708 = n13705 & n13707 ;
  assign n13709 = \m0_s7_cyc_o_reg/NET0131  & \s7_m0_cyc_r_reg/P0001  ;
  assign n13710 = n13697 & n13709 ;
  assign n13711 = n13705 & n13710 ;
  assign n13712 = ~n13708 & ~n13711 ;
  assign n13713 = n13704 & n13712 ;
  assign n13714 = ~n13682 & n13689 ;
  assign n13715 = \m3_s7_cyc_o_reg/NET0131  & \s7_m3_cyc_r_reg/P0001  ;
  assign n13716 = ~n13697 & n13715 ;
  assign n13717 = n13714 & n13716 ;
  assign n13718 = \m2_s7_cyc_o_reg/NET0131  & \s7_m2_cyc_r_reg/P0001  ;
  assign n13719 = n13697 & n13718 ;
  assign n13720 = n13714 & n13719 ;
  assign n13721 = ~n13717 & ~n13720 ;
  assign n13722 = n13682 & ~n13689 ;
  assign n13723 = \m5_s7_cyc_o_reg/NET0131  & \s7_m5_cyc_r_reg/P0001  ;
  assign n13724 = ~n13697 & n13723 ;
  assign n13725 = n13722 & n13724 ;
  assign n13726 = \m4_s7_cyc_o_reg/NET0131  & \s7_m4_cyc_r_reg/P0001  ;
  assign n13727 = n13697 & n13726 ;
  assign n13728 = n13722 & n13727 ;
  assign n13729 = ~n13725 & ~n13728 ;
  assign n13730 = n13721 & n13729 ;
  assign n13731 = n13713 & n13730 ;
  assign n13732 = n5078 & n5100 ;
  assign n13733 = \s1_next_reg/P0001  & n4444 ;
  assign n13734 = n4461 & n13733 ;
  assign n13735 = ~n13732 & n13734 ;
  assign n13736 = \s1_msel_pri_out_reg[0]/NET0131  & ~\s1_next_reg/P0001  ;
  assign n13737 = n4484 & n4501 ;
  assign n13738 = \s1_next_reg/P0001  & ~n13737 ;
  assign n13739 = ~n13736 & ~n13738 ;
  assign n13740 = ~n13735 & n13739 ;
  assign n13741 = ~rst_i_pad & ~n13740 ;
  assign n13742 = ~\s8_msel_pri_out_reg[0]/NET0131  & \s8_msel_pri_out_reg[1]/NET0131  ;
  assign n13743 = \s8_msel_arb2_state_reg[1]/NET0131  & n13742 ;
  assign n13744 = \s8_msel_pri_out_reg[0]/NET0131  & ~\s8_msel_pri_out_reg[1]/NET0131  ;
  assign n13745 = \s8_msel_arb1_state_reg[1]/NET0131  & n13744 ;
  assign n13746 = ~n13743 & ~n13745 ;
  assign n13747 = \s8_msel_pri_out_reg[0]/NET0131  & \s8_msel_pri_out_reg[1]/NET0131  ;
  assign n13748 = \s8_msel_arb3_state_reg[1]/NET0131  & n13747 ;
  assign n13749 = ~\s8_msel_pri_out_reg[0]/NET0131  & ~\s8_msel_pri_out_reg[1]/NET0131  ;
  assign n13750 = \s8_msel_arb0_state_reg[1]/NET0131  & n13749 ;
  assign n13751 = ~n13748 & ~n13750 ;
  assign n13752 = n13746 & n13751 ;
  assign n13753 = \s8_msel_arb2_state_reg[2]/NET0131  & n13742 ;
  assign n13754 = \s8_msel_arb1_state_reg[2]/NET0131  & n13744 ;
  assign n13755 = ~n13753 & ~n13754 ;
  assign n13756 = \s8_msel_arb3_state_reg[2]/NET0131  & n13747 ;
  assign n13757 = \s8_msel_arb0_state_reg[2]/NET0131  & n13749 ;
  assign n13758 = ~n13756 & ~n13757 ;
  assign n13759 = n13755 & n13758 ;
  assign n13760 = n13752 & n13759 ;
  assign n13761 = \s8_msel_arb2_state_reg[0]/NET0131  & n13742 ;
  assign n13762 = \s8_msel_arb1_state_reg[0]/NET0131  & n13744 ;
  assign n13763 = ~n13761 & ~n13762 ;
  assign n13764 = \s8_msel_arb3_state_reg[0]/NET0131  & n13747 ;
  assign n13765 = \s8_msel_arb0_state_reg[0]/NET0131  & n13749 ;
  assign n13766 = ~n13764 & ~n13765 ;
  assign n13767 = n13763 & n13766 ;
  assign n13768 = \m1_s8_cyc_o_reg/NET0131  & \s8_m1_cyc_r_reg/P0001  ;
  assign n13769 = ~n13767 & n13768 ;
  assign n13770 = n13760 & n13769 ;
  assign n13771 = \m0_s8_cyc_o_reg/NET0131  & \s8_m0_cyc_r_reg/P0001  ;
  assign n13772 = n13767 & n13771 ;
  assign n13773 = n13760 & n13772 ;
  assign n13774 = ~n13770 & ~n13773 ;
  assign n13775 = ~n13752 & n13759 ;
  assign n13776 = \m3_s8_cyc_o_reg/NET0131  & \s8_m3_cyc_r_reg/P0001  ;
  assign n13777 = ~n13767 & n13776 ;
  assign n13778 = n13775 & n13777 ;
  assign n13779 = \m2_s8_cyc_o_reg/NET0131  & \s8_m2_cyc_r_reg/P0001  ;
  assign n13780 = n13767 & n13779 ;
  assign n13781 = n13775 & n13780 ;
  assign n13782 = ~n13778 & ~n13781 ;
  assign n13783 = n13774 & n13782 ;
  assign n13784 = ~n13752 & ~n13759 ;
  assign n13785 = \m7_s8_cyc_o_reg/NET0131  & \s8_m7_cyc_r_reg/P0001  ;
  assign n13786 = ~n13767 & n13785 ;
  assign n13787 = n13784 & n13786 ;
  assign n13788 = \m6_s8_cyc_o_reg/NET0131  & \s8_m6_cyc_r_reg/P0001  ;
  assign n13789 = n13767 & n13788 ;
  assign n13790 = n13784 & n13789 ;
  assign n13791 = ~n13787 & ~n13790 ;
  assign n13792 = n13752 & ~n13759 ;
  assign n13793 = \m5_s8_cyc_o_reg/NET0131  & \s8_m5_cyc_r_reg/P0001  ;
  assign n13794 = ~n13767 & n13793 ;
  assign n13795 = n13792 & n13794 ;
  assign n13796 = \m4_s8_cyc_o_reg/NET0131  & \s8_m4_cyc_r_reg/P0001  ;
  assign n13797 = n13767 & n13796 ;
  assign n13798 = n13792 & n13797 ;
  assign n13799 = ~n13795 & ~n13798 ;
  assign n13800 = n13791 & n13799 ;
  assign n13801 = n13783 & n13800 ;
  assign n13802 = n5123 & n5138 ;
  assign n13803 = \s2_next_reg/P0001  & n9904 ;
  assign n13804 = n9921 & n13803 ;
  assign n13805 = ~n13802 & n13804 ;
  assign n13806 = \s2_msel_pri_out_reg[0]/NET0131  & ~\s2_next_reg/P0001  ;
  assign n13807 = n3975 & n3980 ;
  assign n13808 = \s2_next_reg/P0001  & ~n13807 ;
  assign n13809 = ~n13806 & ~n13808 ;
  assign n13810 = ~n13805 & n13809 ;
  assign n13811 = ~rst_i_pad & ~n13810 ;
  assign n13812 = n5153 & n5180 ;
  assign n13813 = \s3_next_reg/P0001  & n4008 ;
  assign n13814 = n4025 & n13813 ;
  assign n13815 = ~n13812 & n13814 ;
  assign n13816 = \s3_msel_pri_out_reg[0]/NET0131  & ~\s3_next_reg/P0001  ;
  assign n13817 = n4535 & n4552 ;
  assign n13818 = \s3_next_reg/P0001  & ~n13817 ;
  assign n13819 = ~n13816 & ~n13818 ;
  assign n13820 = ~n13815 & n13819 ;
  assign n13821 = ~rst_i_pad & ~n13820 ;
  assign n13822 = ~\s9_msel_pri_out_reg[0]/NET0131  & \s9_msel_pri_out_reg[1]/NET0131  ;
  assign n13823 = \s9_msel_arb2_state_reg[1]/NET0131  & n13822 ;
  assign n13824 = \s9_msel_pri_out_reg[0]/NET0131  & ~\s9_msel_pri_out_reg[1]/NET0131  ;
  assign n13825 = \s9_msel_arb1_state_reg[1]/NET0131  & n13824 ;
  assign n13826 = ~n13823 & ~n13825 ;
  assign n13827 = \s9_msel_pri_out_reg[0]/NET0131  & \s9_msel_pri_out_reg[1]/NET0131  ;
  assign n13828 = \s9_msel_arb3_state_reg[1]/NET0131  & n13827 ;
  assign n13829 = ~\s9_msel_pri_out_reg[0]/NET0131  & ~\s9_msel_pri_out_reg[1]/NET0131  ;
  assign n13830 = \s9_msel_arb0_state_reg[1]/NET0131  & n13829 ;
  assign n13831 = ~n13828 & ~n13830 ;
  assign n13832 = n13826 & n13831 ;
  assign n13833 = \s9_msel_arb2_state_reg[2]/NET0131  & n13822 ;
  assign n13834 = \s9_msel_arb1_state_reg[2]/NET0131  & n13824 ;
  assign n13835 = ~n13833 & ~n13834 ;
  assign n13836 = \s9_msel_arb3_state_reg[2]/NET0131  & n13827 ;
  assign n13837 = \s9_msel_arb0_state_reg[2]/NET0131  & n13829 ;
  assign n13838 = ~n13836 & ~n13837 ;
  assign n13839 = n13835 & n13838 ;
  assign n13840 = ~n13832 & n13839 ;
  assign n13841 = \s9_msel_arb2_state_reg[0]/NET0131  & n13822 ;
  assign n13842 = \s9_msel_arb1_state_reg[0]/NET0131  & n13824 ;
  assign n13843 = ~n13841 & ~n13842 ;
  assign n13844 = \s9_msel_arb3_state_reg[0]/NET0131  & n13827 ;
  assign n13845 = \s9_msel_arb0_state_reg[0]/NET0131  & n13829 ;
  assign n13846 = ~n13844 & ~n13845 ;
  assign n13847 = n13843 & n13846 ;
  assign n13848 = \m3_s9_cyc_o_reg/NET0131  & \s9_m3_cyc_r_reg/P0001  ;
  assign n13849 = ~n13847 & n13848 ;
  assign n13850 = n13840 & n13849 ;
  assign n13851 = \m2_s9_cyc_o_reg/NET0131  & \s9_m2_cyc_r_reg/P0001  ;
  assign n13852 = n13847 & n13851 ;
  assign n13853 = n13840 & n13852 ;
  assign n13854 = ~n13850 & ~n13853 ;
  assign n13855 = n13832 & n13839 ;
  assign n13856 = \m1_s9_cyc_o_reg/NET0131  & \s9_m1_cyc_r_reg/P0001  ;
  assign n13857 = ~n13847 & n13856 ;
  assign n13858 = n13855 & n13857 ;
  assign n13859 = \m0_s9_cyc_o_reg/NET0131  & \s9_m0_cyc_r_reg/P0001  ;
  assign n13860 = n13847 & n13859 ;
  assign n13861 = n13855 & n13860 ;
  assign n13862 = ~n13858 & ~n13861 ;
  assign n13863 = n13854 & n13862 ;
  assign n13864 = ~n13832 & ~n13839 ;
  assign n13865 = \m7_s9_cyc_o_reg/NET0131  & \s9_m7_cyc_r_reg/P0001  ;
  assign n13866 = ~n13847 & n13865 ;
  assign n13867 = n13864 & n13866 ;
  assign n13868 = \m6_s9_cyc_o_reg/NET0131  & \s9_m6_cyc_r_reg/P0001  ;
  assign n13869 = n13847 & n13868 ;
  assign n13870 = n13864 & n13869 ;
  assign n13871 = ~n13867 & ~n13870 ;
  assign n13872 = n13832 & ~n13839 ;
  assign n13873 = \m5_s9_cyc_o_reg/NET0131  & \s9_m5_cyc_r_reg/P0001  ;
  assign n13874 = ~n13847 & n13873 ;
  assign n13875 = n13872 & n13874 ;
  assign n13876 = \m4_s9_cyc_o_reg/NET0131  & \s9_m4_cyc_r_reg/P0001  ;
  assign n13877 = n13847 & n13876 ;
  assign n13878 = n13872 & n13877 ;
  assign n13879 = ~n13875 & ~n13878 ;
  assign n13880 = n13871 & n13879 ;
  assign n13881 = n13863 & n13880 ;
  assign n13882 = n5193 & n5215 ;
  assign n13883 = \s4_next_reg/P0001  & n9931 ;
  assign n13884 = n9948 & n13883 ;
  assign n13885 = ~n13882 & n13884 ;
  assign n13886 = \s4_msel_pri_out_reg[0]/NET0131  & ~\s4_next_reg/P0001  ;
  assign n13887 = n4048 & n4065 ;
  assign n13888 = \s4_next_reg/P0001  & ~n13887 ;
  assign n13889 = ~n13886 & ~n13888 ;
  assign n13890 = ~n13885 & n13889 ;
  assign n13891 = ~rst_i_pad & ~n13890 ;
  assign n13892 = \s5_next_reg/P0001  & n4581 ;
  assign n13893 = n4598 & n13892 ;
  assign n13894 = n5228 & n5231 ;
  assign n13895 = n5240 & n13894 ;
  assign n13896 = n13893 & ~n13895 ;
  assign n13897 = \s5_msel_pri_out_reg[0]/NET0131  & ~\s5_next_reg/P0001  ;
  assign n13898 = n4637 & n4642 ;
  assign n13899 = \s5_next_reg/P0001  & ~n13898 ;
  assign n13900 = ~n13897 & ~n13899 ;
  assign n13901 = ~n13896 & n13900 ;
  assign n13902 = ~rst_i_pad & ~n13901 ;
  assign n13903 = ~\s10_msel_pri_out_reg[0]/NET0131  & ~\s10_msel_pri_out_reg[1]/NET0131  ;
  assign n13904 = \s10_msel_arb0_state_reg[1]/NET0131  & n13903 ;
  assign n13905 = \s10_msel_pri_out_reg[0]/NET0131  & \s10_msel_pri_out_reg[1]/NET0131  ;
  assign n13906 = \s10_msel_arb3_state_reg[1]/NET0131  & n13905 ;
  assign n13907 = ~n13904 & ~n13906 ;
  assign n13908 = \s10_msel_pri_out_reg[0]/NET0131  & ~\s10_msel_pri_out_reg[1]/NET0131  ;
  assign n13909 = \s10_msel_arb1_state_reg[1]/NET0131  & n13908 ;
  assign n13910 = ~\s10_msel_pri_out_reg[0]/NET0131  & \s10_msel_pri_out_reg[1]/NET0131  ;
  assign n13911 = \s10_msel_arb2_state_reg[1]/NET0131  & n13910 ;
  assign n13912 = ~n13909 & ~n13911 ;
  assign n13913 = n13907 & n13912 ;
  assign n13914 = \s10_msel_arb0_state_reg[2]/NET0131  & n13903 ;
  assign n13915 = \s10_msel_arb3_state_reg[2]/NET0131  & n13905 ;
  assign n13916 = ~n13914 & ~n13915 ;
  assign n13917 = \s10_msel_arb1_state_reg[2]/NET0131  & n13908 ;
  assign n13918 = \s10_msel_arb2_state_reg[2]/NET0131  & n13910 ;
  assign n13919 = ~n13917 & ~n13918 ;
  assign n13920 = n13916 & n13919 ;
  assign n13921 = ~n13913 & n13920 ;
  assign n13922 = \s10_msel_arb0_state_reg[0]/NET0131  & n13903 ;
  assign n13923 = \s10_msel_arb3_state_reg[0]/NET0131  & n13905 ;
  assign n13924 = ~n13922 & ~n13923 ;
  assign n13925 = \s10_msel_arb1_state_reg[0]/NET0131  & n13908 ;
  assign n13926 = \s10_msel_arb2_state_reg[0]/NET0131  & n13910 ;
  assign n13927 = ~n13925 & ~n13926 ;
  assign n13928 = n13924 & n13927 ;
  assign n13929 = \m3_s10_cyc_o_reg/NET0131  & \s10_m3_cyc_r_reg/P0001  ;
  assign n13930 = ~n13928 & n13929 ;
  assign n13931 = n13921 & n13930 ;
  assign n13932 = \m2_s10_cyc_o_reg/NET0131  & \s10_m2_cyc_r_reg/P0001  ;
  assign n13933 = n13928 & n13932 ;
  assign n13934 = n13921 & n13933 ;
  assign n13935 = ~n13931 & ~n13934 ;
  assign n13936 = ~n13913 & ~n13920 ;
  assign n13937 = \m7_s10_cyc_o_reg/NET0131  & \s10_m7_cyc_r_reg/P0001  ;
  assign n13938 = ~n13928 & n13937 ;
  assign n13939 = n13936 & n13938 ;
  assign n13940 = \m6_s10_cyc_o_reg/NET0131  & \s10_m6_cyc_r_reg/P0001  ;
  assign n13941 = n13928 & n13940 ;
  assign n13942 = n13936 & n13941 ;
  assign n13943 = ~n13939 & ~n13942 ;
  assign n13944 = n13935 & n13943 ;
  assign n13945 = n13913 & n13920 ;
  assign n13946 = \m1_s10_cyc_o_reg/NET0131  & \s10_m1_cyc_r_reg/P0001  ;
  assign n13947 = ~n13928 & n13946 ;
  assign n13948 = n13945 & n13947 ;
  assign n13949 = \m0_s10_cyc_o_reg/NET0131  & \s10_m0_cyc_r_reg/P0001  ;
  assign n13950 = n13928 & n13949 ;
  assign n13951 = n13945 & n13950 ;
  assign n13952 = ~n13948 & ~n13951 ;
  assign n13953 = n13913 & ~n13920 ;
  assign n13954 = \m5_s10_cyc_o_reg/NET0131  & \s10_m5_cyc_r_reg/P0001  ;
  assign n13955 = ~n13928 & n13954 ;
  assign n13956 = n13953 & n13955 ;
  assign n13957 = \m4_s10_cyc_o_reg/NET0131  & \s10_m4_cyc_r_reg/P0001  ;
  assign n13958 = n13928 & n13957 ;
  assign n13959 = n13953 & n13958 ;
  assign n13960 = ~n13956 & ~n13959 ;
  assign n13961 = n13952 & n13960 ;
  assign n13962 = n13944 & n13961 ;
  assign n13963 = \s6_next_reg/P0001  & n4094 ;
  assign n13964 = n4111 & n13963 ;
  assign n13965 = n5271 & n5274 ;
  assign n13966 = n5283 & n13965 ;
  assign n13967 = n13964 & ~n13966 ;
  assign n13968 = \s6_msel_pri_out_reg[0]/NET0131  & ~\s6_next_reg/P0001  ;
  assign n13969 = n4691 & n4696 ;
  assign n13970 = \s6_next_reg/P0001  & ~n13969 ;
  assign n13971 = ~n13968 & ~n13970 ;
  assign n13972 = ~n13967 & n13971 ;
  assign n13973 = ~rst_i_pad & ~n13972 ;
  assign n13974 = n5318 & n5325 ;
  assign n13975 = \s7_next_reg/P0001  & n9965 ;
  assign n13976 = n9975 & n13975 ;
  assign n13977 = ~n13974 & n13976 ;
  assign n13978 = \s7_msel_pri_out_reg[0]/NET0131  & ~\s7_next_reg/P0001  ;
  assign n13979 = n4745 & n4750 ;
  assign n13980 = \s7_next_reg/P0001  & ~n13979 ;
  assign n13981 = ~n13978 & ~n13980 ;
  assign n13982 = ~n13977 & n13981 ;
  assign n13983 = ~rst_i_pad & ~n13982 ;
  assign n13984 = ~\s11_msel_pri_out_reg[0]/NET0131  & \s11_msel_pri_out_reg[1]/NET0131  ;
  assign n13985 = \s11_msel_arb2_state_reg[1]/NET0131  & n13984 ;
  assign n13986 = \s11_msel_pri_out_reg[0]/NET0131  & ~\s11_msel_pri_out_reg[1]/NET0131  ;
  assign n13987 = \s11_msel_arb1_state_reg[1]/NET0131  & n13986 ;
  assign n13988 = ~n13985 & ~n13987 ;
  assign n13989 = \s11_msel_pri_out_reg[0]/NET0131  & \s11_msel_pri_out_reg[1]/NET0131  ;
  assign n13990 = \s11_msel_arb3_state_reg[1]/NET0131  & n13989 ;
  assign n13991 = ~\s11_msel_pri_out_reg[0]/NET0131  & ~\s11_msel_pri_out_reg[1]/NET0131  ;
  assign n13992 = \s11_msel_arb0_state_reg[1]/NET0131  & n13991 ;
  assign n13993 = ~n13990 & ~n13992 ;
  assign n13994 = n13988 & n13993 ;
  assign n13995 = \s11_msel_arb1_state_reg[2]/NET0131  & n13986 ;
  assign n13996 = \s11_msel_arb2_state_reg[2]/NET0131  & n13984 ;
  assign n13997 = ~n13995 & ~n13996 ;
  assign n13998 = \s11_msel_arb3_state_reg[2]/NET0131  & n13989 ;
  assign n13999 = \s11_msel_arb0_state_reg[2]/NET0131  & n13991 ;
  assign n14000 = ~n13998 & ~n13999 ;
  assign n14001 = n13997 & n14000 ;
  assign n14002 = n13994 & ~n14001 ;
  assign n14003 = \s11_msel_arb2_state_reg[0]/NET0131  & n13984 ;
  assign n14004 = \s11_msel_arb1_state_reg[0]/NET0131  & n13986 ;
  assign n14005 = ~n14003 & ~n14004 ;
  assign n14006 = \s11_msel_arb3_state_reg[0]/NET0131  & n13989 ;
  assign n14007 = \s11_msel_arb0_state_reg[0]/NET0131  & n13991 ;
  assign n14008 = ~n14006 & ~n14007 ;
  assign n14009 = n14005 & n14008 ;
  assign n14010 = \m5_s11_cyc_o_reg/NET0131  & \s11_m5_cyc_r_reg/P0001  ;
  assign n14011 = ~n14009 & n14010 ;
  assign n14012 = n14002 & n14011 ;
  assign n14013 = \m4_s11_cyc_o_reg/NET0131  & \s11_m4_cyc_r_reg/P0001  ;
  assign n14014 = n14009 & n14013 ;
  assign n14015 = n14002 & n14014 ;
  assign n14016 = ~n14012 & ~n14015 ;
  assign n14017 = n13994 & n14001 ;
  assign n14018 = \m1_s11_cyc_o_reg/NET0131  & \s11_m1_cyc_r_reg/P0001  ;
  assign n14019 = ~n14009 & n14018 ;
  assign n14020 = n14017 & n14019 ;
  assign n14021 = \m0_s11_cyc_o_reg/NET0131  & \s11_m0_cyc_r_reg/P0001  ;
  assign n14022 = n14009 & n14021 ;
  assign n14023 = n14017 & n14022 ;
  assign n14024 = ~n14020 & ~n14023 ;
  assign n14025 = n14016 & n14024 ;
  assign n14026 = ~n13994 & ~n14001 ;
  assign n14027 = \m7_s11_cyc_o_reg/NET0131  & \s11_m7_cyc_r_reg/P0001  ;
  assign n14028 = ~n14009 & n14027 ;
  assign n14029 = n14026 & n14028 ;
  assign n14030 = \m6_s11_cyc_o_reg/NET0131  & \s11_m6_cyc_r_reg/P0001  ;
  assign n14031 = n14009 & n14030 ;
  assign n14032 = n14026 & n14031 ;
  assign n14033 = ~n14029 & ~n14032 ;
  assign n14034 = ~n13994 & n14001 ;
  assign n14035 = \m3_s11_cyc_o_reg/NET0131  & \s11_m3_cyc_r_reg/P0001  ;
  assign n14036 = ~n14009 & n14035 ;
  assign n14037 = n14034 & n14036 ;
  assign n14038 = \m2_s11_cyc_o_reg/NET0131  & \s11_m2_cyc_r_reg/P0001  ;
  assign n14039 = n14009 & n14038 ;
  assign n14040 = n14034 & n14039 ;
  assign n14041 = ~n14037 & ~n14040 ;
  assign n14042 = n14033 & n14041 ;
  assign n14043 = n14025 & n14042 ;
  assign n14044 = ~\s0_msel_pri_out_reg[0]/NET0131  & \s0_msel_pri_out_reg[1]/NET0131  ;
  assign n14045 = \s0_msel_arb2_state_reg[1]/NET0131  & n14044 ;
  assign n14046 = \s0_msel_pri_out_reg[0]/NET0131  & ~\s0_msel_pri_out_reg[1]/NET0131  ;
  assign n14047 = \s0_msel_arb1_state_reg[1]/NET0131  & n14046 ;
  assign n14048 = ~n14045 & ~n14047 ;
  assign n14049 = \s0_msel_pri_out_reg[0]/NET0131  & \s0_msel_pri_out_reg[1]/NET0131  ;
  assign n14050 = \s0_msel_arb3_state_reg[1]/NET0131  & n14049 ;
  assign n14051 = ~\s0_msel_pri_out_reg[0]/NET0131  & ~\s0_msel_pri_out_reg[1]/NET0131  ;
  assign n14052 = \s0_msel_arb0_state_reg[1]/NET0131  & n14051 ;
  assign n14053 = ~n14050 & ~n14052 ;
  assign n14054 = n14048 & n14053 ;
  assign n14055 = \s0_msel_arb2_state_reg[2]/NET0131  & n14044 ;
  assign n14056 = \s0_msel_arb1_state_reg[2]/NET0131  & n14046 ;
  assign n14057 = ~n14055 & ~n14056 ;
  assign n14058 = \s0_msel_arb3_state_reg[2]/NET0131  & n14049 ;
  assign n14059 = \s0_msel_arb0_state_reg[2]/NET0131  & n14051 ;
  assign n14060 = ~n14058 & ~n14059 ;
  assign n14061 = n14057 & n14060 ;
  assign n14062 = ~n14054 & ~n14061 ;
  assign n14063 = \s0_msel_arb0_state_reg[0]/NET0131  & n14051 ;
  assign n14064 = \s0_msel_arb3_state_reg[0]/NET0131  & n14049 ;
  assign n14065 = ~n14063 & ~n14064 ;
  assign n14066 = \s0_msel_arb1_state_reg[0]/NET0131  & n14046 ;
  assign n14067 = \s0_msel_arb2_state_reg[0]/NET0131  & n14044 ;
  assign n14068 = ~n14066 & ~n14067 ;
  assign n14069 = n14065 & n14068 ;
  assign n14070 = \m7_s0_cyc_o_reg/NET0131  & \s0_m7_cyc_r_reg/P0001  ;
  assign n14071 = ~n14069 & n14070 ;
  assign n14072 = n14062 & n14071 ;
  assign n14073 = \m6_s0_cyc_o_reg/NET0131  & \s0_m6_cyc_r_reg/P0001  ;
  assign n14074 = n14069 & n14073 ;
  assign n14075 = n14062 & n14074 ;
  assign n14076 = ~n14072 & ~n14075 ;
  assign n14077 = n14054 & ~n14061 ;
  assign n14078 = \m5_s0_cyc_o_reg/NET0131  & \s0_m5_cyc_r_reg/P0001  ;
  assign n14079 = ~n14069 & n14078 ;
  assign n14080 = n14077 & n14079 ;
  assign n14081 = \m4_s0_cyc_o_reg/NET0131  & \s0_m4_cyc_r_reg/P0001  ;
  assign n14082 = n14069 & n14081 ;
  assign n14083 = n14077 & n14082 ;
  assign n14084 = ~n14080 & ~n14083 ;
  assign n14085 = n14076 & n14084 ;
  assign n14086 = ~n14054 & n14061 ;
  assign n14087 = \m3_s0_cyc_o_reg/NET0131  & \s0_m3_cyc_r_reg/P0001  ;
  assign n14088 = ~n14069 & n14087 ;
  assign n14089 = n14086 & n14088 ;
  assign n14090 = \m2_s0_cyc_o_reg/NET0131  & \s0_m2_cyc_r_reg/P0001  ;
  assign n14091 = n14069 & n14090 ;
  assign n14092 = n14086 & n14091 ;
  assign n14093 = ~n14089 & ~n14092 ;
  assign n14094 = n14054 & n14061 ;
  assign n14095 = \m1_s0_cyc_o_reg/NET0131  & \s0_m1_cyc_r_reg/P0001  ;
  assign n14096 = ~n14069 & n14095 ;
  assign n14097 = n14094 & n14096 ;
  assign n14098 = \m0_s0_cyc_o_reg/NET0131  & \s0_m0_cyc_r_reg/P0001  ;
  assign n14099 = n14069 & n14098 ;
  assign n14100 = n14094 & n14099 ;
  assign n14101 = ~n14097 & ~n14100 ;
  assign n14102 = n14093 & n14101 ;
  assign n14103 = n14085 & n14102 ;
  assign n14104 = \s8_next_reg/P0001  & n4129 ;
  assign n14105 = n4146 & n14104 ;
  assign n14106 = n5352 & n5355 ;
  assign n14107 = n5364 & n14106 ;
  assign n14108 = n14105 & ~n14107 ;
  assign n14109 = \s8_msel_pri_out_reg[0]/NET0131  & ~\s8_next_reg/P0001  ;
  assign n14110 = n4783 & n4800 ;
  assign n14111 = \s8_next_reg/P0001  & ~n14110 ;
  assign n14112 = ~n14109 & ~n14111 ;
  assign n14113 = ~n14108 & n14112 ;
  assign n14114 = ~rst_i_pad & ~n14113 ;
  assign n14115 = ~\s12_msel_pri_out_reg[0]/NET0131  & \s12_msel_pri_out_reg[1]/NET0131  ;
  assign n14116 = \s12_msel_arb2_state_reg[1]/NET0131  & n14115 ;
  assign n14117 = \s12_msel_pri_out_reg[0]/NET0131  & ~\s12_msel_pri_out_reg[1]/NET0131  ;
  assign n14118 = \s12_msel_arb1_state_reg[1]/NET0131  & n14117 ;
  assign n14119 = ~n14116 & ~n14118 ;
  assign n14120 = \s12_msel_pri_out_reg[0]/NET0131  & \s12_msel_pri_out_reg[1]/NET0131  ;
  assign n14121 = \s12_msel_arb3_state_reg[1]/NET0131  & n14120 ;
  assign n14122 = ~\s12_msel_pri_out_reg[0]/NET0131  & ~\s12_msel_pri_out_reg[1]/NET0131  ;
  assign n14123 = \s12_msel_arb0_state_reg[1]/NET0131  & n14122 ;
  assign n14124 = ~n14121 & ~n14123 ;
  assign n14125 = n14119 & n14124 ;
  assign n14126 = \s12_msel_arb0_state_reg[2]/NET0131  & n14122 ;
  assign n14127 = \s12_msel_arb2_state_reg[2]/NET0131  & n14115 ;
  assign n14128 = ~n14126 & ~n14127 ;
  assign n14129 = \s12_msel_arb3_state_reg[2]/NET0131  & n14120 ;
  assign n14130 = \s12_msel_arb1_state_reg[2]/NET0131  & n14117 ;
  assign n14131 = ~n14129 & ~n14130 ;
  assign n14132 = n14128 & n14131 ;
  assign n14133 = ~n14125 & n14132 ;
  assign n14134 = \s12_msel_arb2_state_reg[0]/NET0131  & n14115 ;
  assign n14135 = \s12_msel_arb1_state_reg[0]/NET0131  & n14117 ;
  assign n14136 = ~n14134 & ~n14135 ;
  assign n14137 = \s12_msel_arb3_state_reg[0]/NET0131  & n14120 ;
  assign n14138 = \s12_msel_arb0_state_reg[0]/NET0131  & n14122 ;
  assign n14139 = ~n14137 & ~n14138 ;
  assign n14140 = n14136 & n14139 ;
  assign n14141 = \m3_s12_cyc_o_reg/NET0131  & \s12_m3_cyc_r_reg/P0001  ;
  assign n14142 = ~n14140 & n14141 ;
  assign n14143 = n14133 & n14142 ;
  assign n14144 = \m2_s12_cyc_o_reg/NET0131  & \s12_m2_cyc_r_reg/P0001  ;
  assign n14145 = n14140 & n14144 ;
  assign n14146 = n14133 & n14145 ;
  assign n14147 = ~n14143 & ~n14146 ;
  assign n14148 = ~n14125 & ~n14132 ;
  assign n14149 = \m7_s12_cyc_o_reg/NET0131  & \s12_m7_cyc_r_reg/P0001  ;
  assign n14150 = ~n14140 & n14149 ;
  assign n14151 = n14148 & n14150 ;
  assign n14152 = \m6_s12_cyc_o_reg/NET0131  & \s12_m6_cyc_r_reg/P0001  ;
  assign n14153 = n14140 & n14152 ;
  assign n14154 = n14148 & n14153 ;
  assign n14155 = ~n14151 & ~n14154 ;
  assign n14156 = n14147 & n14155 ;
  assign n14157 = n14125 & ~n14132 ;
  assign n14158 = \m5_s12_cyc_o_reg/NET0131  & \s12_m5_cyc_r_reg/P0001  ;
  assign n14159 = ~n14140 & n14158 ;
  assign n14160 = n14157 & n14159 ;
  assign n14161 = \m4_s12_cyc_o_reg/NET0131  & \s12_m4_cyc_r_reg/P0001  ;
  assign n14162 = n14140 & n14161 ;
  assign n14163 = n14157 & n14162 ;
  assign n14164 = ~n14160 & ~n14163 ;
  assign n14165 = n14125 & n14132 ;
  assign n14166 = \m1_s12_cyc_o_reg/NET0131  & \s12_m1_cyc_r_reg/P0001  ;
  assign n14167 = ~n14140 & n14166 ;
  assign n14168 = n14165 & n14167 ;
  assign n14169 = \m0_s12_cyc_o_reg/NET0131  & \s12_m0_cyc_r_reg/P0001  ;
  assign n14170 = n14140 & n14169 ;
  assign n14171 = n14165 & n14170 ;
  assign n14172 = ~n14168 & ~n14171 ;
  assign n14173 = n14164 & n14172 ;
  assign n14174 = n14156 & n14173 ;
  assign n14175 = \s9_next_reg/P0001  & n10000 ;
  assign n14176 = n10010 & n14175 ;
  assign n14177 = n5397 & n5402 ;
  assign n14178 = n5415 & n14177 ;
  assign n14179 = n14176 & ~n14178 ;
  assign n14180 = n10028 & n10045 ;
  assign n14181 = \s9_next_reg/P0001  & ~n14180 ;
  assign n14182 = \s9_msel_pri_out_reg[0]/NET0131  & ~\s9_next_reg/P0001  ;
  assign n14183 = ~n14181 & ~n14182 ;
  assign n14184 = ~n14179 & n14183 ;
  assign n14185 = ~rst_i_pad & ~n14184 ;
  assign n14186 = \s13_msel_pri_out_reg[0]/NET0131  & ~\s13_msel_pri_out_reg[1]/NET0131  ;
  assign n14187 = \s13_msel_arb1_state_reg[1]/NET0131  & n14186 ;
  assign n14188 = ~\s13_msel_pri_out_reg[0]/NET0131  & \s13_msel_pri_out_reg[1]/NET0131  ;
  assign n14189 = \s13_msel_arb2_state_reg[1]/NET0131  & n14188 ;
  assign n14190 = ~n14187 & ~n14189 ;
  assign n14191 = \s13_msel_pri_out_reg[0]/NET0131  & \s13_msel_pri_out_reg[1]/NET0131  ;
  assign n14192 = \s13_msel_arb3_state_reg[1]/NET0131  & n14191 ;
  assign n14193 = ~\s13_msel_pri_out_reg[0]/NET0131  & ~\s13_msel_pri_out_reg[1]/NET0131  ;
  assign n14194 = \s13_msel_arb0_state_reg[1]/NET0131  & n14193 ;
  assign n14195 = ~n14192 & ~n14194 ;
  assign n14196 = n14190 & n14195 ;
  assign n14197 = \s13_msel_arb0_state_reg[2]/NET0131  & n14193 ;
  assign n14198 = \s13_msel_arb3_state_reg[2]/NET0131  & n14191 ;
  assign n14199 = ~n14197 & ~n14198 ;
  assign n14200 = \s13_msel_arb1_state_reg[2]/NET0131  & n14186 ;
  assign n14201 = \s13_msel_arb2_state_reg[2]/NET0131  & n14188 ;
  assign n14202 = ~n14200 & ~n14201 ;
  assign n14203 = n14199 & n14202 ;
  assign n14204 = ~n14196 & ~n14203 ;
  assign n14205 = \s13_msel_arb2_state_reg[0]/NET0131  & n14188 ;
  assign n14206 = \s13_msel_arb1_state_reg[0]/NET0131  & n14186 ;
  assign n14207 = ~n14205 & ~n14206 ;
  assign n14208 = \s13_msel_arb3_state_reg[0]/NET0131  & n14191 ;
  assign n14209 = \s13_msel_arb0_state_reg[0]/NET0131  & n14193 ;
  assign n14210 = ~n14208 & ~n14209 ;
  assign n14211 = n14207 & n14210 ;
  assign n14212 = \m7_s13_cyc_o_reg/NET0131  & \s13_m7_cyc_r_reg/P0001  ;
  assign n14213 = ~n14211 & n14212 ;
  assign n14214 = n14204 & n14213 ;
  assign n14215 = \m6_s13_cyc_o_reg/NET0131  & \s13_m6_cyc_r_reg/P0001  ;
  assign n14216 = n14211 & n14215 ;
  assign n14217 = n14204 & n14216 ;
  assign n14218 = ~n14214 & ~n14217 ;
  assign n14219 = n14196 & n14203 ;
  assign n14220 = \m1_s13_cyc_o_reg/NET0131  & \s13_m1_cyc_r_reg/P0001  ;
  assign n14221 = ~n14211 & n14220 ;
  assign n14222 = n14219 & n14221 ;
  assign n14223 = \m0_s13_cyc_o_reg/NET0131  & \s13_m0_cyc_r_reg/P0001  ;
  assign n14224 = n14211 & n14223 ;
  assign n14225 = n14219 & n14224 ;
  assign n14226 = ~n14222 & ~n14225 ;
  assign n14227 = n14218 & n14226 ;
  assign n14228 = ~n14196 & n14203 ;
  assign n14229 = \m3_s13_cyc_o_reg/NET0131  & \s13_m3_cyc_r_reg/P0001  ;
  assign n14230 = ~n14211 & n14229 ;
  assign n14231 = n14228 & n14230 ;
  assign n14232 = \m2_s13_cyc_o_reg/NET0131  & \s13_m2_cyc_r_reg/P0001  ;
  assign n14233 = n14211 & n14232 ;
  assign n14234 = n14228 & n14233 ;
  assign n14235 = ~n14231 & ~n14234 ;
  assign n14236 = n14196 & ~n14203 ;
  assign n14237 = \m5_s13_cyc_o_reg/NET0131  & \s13_m5_cyc_r_reg/P0001  ;
  assign n14238 = ~n14211 & n14237 ;
  assign n14239 = n14236 & n14238 ;
  assign n14240 = \m4_s13_cyc_o_reg/NET0131  & \s13_m4_cyc_r_reg/P0001  ;
  assign n14241 = n14211 & n14240 ;
  assign n14242 = n14236 & n14241 ;
  assign n14243 = ~n14239 & ~n14242 ;
  assign n14244 = n14235 & n14243 ;
  assign n14245 = n14227 & n14244 ;
  assign n14246 = ~\s1_msel_pri_out_reg[0]/NET0131  & \s1_msel_pri_out_reg[1]/NET0131  ;
  assign n14247 = \s1_msel_arb2_state_reg[1]/NET0131  & n14246 ;
  assign n14248 = \s1_msel_pri_out_reg[0]/NET0131  & ~\s1_msel_pri_out_reg[1]/NET0131  ;
  assign n14249 = \s1_msel_arb1_state_reg[1]/NET0131  & n14248 ;
  assign n14250 = ~n14247 & ~n14249 ;
  assign n14251 = \s1_msel_pri_out_reg[0]/NET0131  & \s1_msel_pri_out_reg[1]/NET0131  ;
  assign n14252 = \s1_msel_arb3_state_reg[1]/NET0131  & n14251 ;
  assign n14253 = ~\s1_msel_pri_out_reg[0]/NET0131  & ~\s1_msel_pri_out_reg[1]/NET0131  ;
  assign n14254 = \s1_msel_arb0_state_reg[1]/NET0131  & n14253 ;
  assign n14255 = ~n14252 & ~n14254 ;
  assign n14256 = n14250 & n14255 ;
  assign n14257 = \s1_msel_arb0_state_reg[2]/NET0131  & n14253 ;
  assign n14258 = \s1_msel_arb3_state_reg[2]/NET0131  & n14251 ;
  assign n14259 = ~n14257 & ~n14258 ;
  assign n14260 = \s1_msel_arb1_state_reg[2]/NET0131  & n14248 ;
  assign n14261 = \s1_msel_arb2_state_reg[2]/NET0131  & n14246 ;
  assign n14262 = ~n14260 & ~n14261 ;
  assign n14263 = n14259 & n14262 ;
  assign n14264 = ~n14256 & ~n14263 ;
  assign n14265 = \s1_msel_arb2_state_reg[0]/NET0131  & n14246 ;
  assign n14266 = \s1_msel_arb1_state_reg[0]/NET0131  & n14248 ;
  assign n14267 = ~n14265 & ~n14266 ;
  assign n14268 = \s1_msel_arb3_state_reg[0]/NET0131  & n14251 ;
  assign n14269 = \s1_msel_arb0_state_reg[0]/NET0131  & n14253 ;
  assign n14270 = ~n14268 & ~n14269 ;
  assign n14271 = n14267 & n14270 ;
  assign n14272 = \m7_s1_cyc_o_reg/NET0131  & \s1_m7_cyc_r_reg/P0001  ;
  assign n14273 = ~n14271 & n14272 ;
  assign n14274 = n14264 & n14273 ;
  assign n14275 = \m6_s1_cyc_o_reg/NET0131  & \s1_m6_cyc_r_reg/P0001  ;
  assign n14276 = n14271 & n14275 ;
  assign n14277 = n14264 & n14276 ;
  assign n14278 = ~n14274 & ~n14277 ;
  assign n14279 = ~n14256 & n14263 ;
  assign n14280 = \m3_s1_cyc_o_reg/NET0131  & \s1_m3_cyc_r_reg/P0001  ;
  assign n14281 = ~n14271 & n14280 ;
  assign n14282 = n14279 & n14281 ;
  assign n14283 = \m2_s1_cyc_o_reg/NET0131  & \s1_m2_cyc_r_reg/P0001  ;
  assign n14284 = n14271 & n14283 ;
  assign n14285 = n14279 & n14284 ;
  assign n14286 = ~n14282 & ~n14285 ;
  assign n14287 = n14278 & n14286 ;
  assign n14288 = n14256 & ~n14263 ;
  assign n14289 = \m5_s1_cyc_o_reg/NET0131  & \s1_m5_cyc_r_reg/P0001  ;
  assign n14290 = ~n14271 & n14289 ;
  assign n14291 = n14288 & n14290 ;
  assign n14292 = \m4_s1_cyc_o_reg/NET0131  & \s1_m4_cyc_r_reg/P0001  ;
  assign n14293 = n14271 & n14292 ;
  assign n14294 = n14288 & n14293 ;
  assign n14295 = ~n14291 & ~n14294 ;
  assign n14296 = n14256 & n14263 ;
  assign n14297 = \m1_s1_cyc_o_reg/NET0131  & \s1_m1_cyc_r_reg/P0001  ;
  assign n14298 = ~n14271 & n14297 ;
  assign n14299 = n14296 & n14298 ;
  assign n14300 = \m0_s1_cyc_o_reg/NET0131  & \s1_m0_cyc_r_reg/P0001  ;
  assign n14301 = n14271 & n14300 ;
  assign n14302 = n14296 & n14301 ;
  assign n14303 = ~n14299 & ~n14302 ;
  assign n14304 = n14295 & n14303 ;
  assign n14305 = n14287 & n14304 ;
  assign n14306 = \s14_msel_pri_out_reg[0]/NET0131  & ~\s14_msel_pri_out_reg[1]/NET0131  ;
  assign n14307 = \s14_msel_arb1_state_reg[2]/NET0131  & n14306 ;
  assign n14308 = ~\s14_msel_pri_out_reg[0]/NET0131  & \s14_msel_pri_out_reg[1]/NET0131  ;
  assign n14309 = \s14_msel_arb2_state_reg[2]/NET0131  & n14308 ;
  assign n14310 = ~n14307 & ~n14309 ;
  assign n14311 = \s14_msel_pri_out_reg[0]/NET0131  & \s14_msel_pri_out_reg[1]/NET0131  ;
  assign n14312 = \s14_msel_arb3_state_reg[2]/NET0131  & n14311 ;
  assign n14313 = ~\s14_msel_pri_out_reg[0]/NET0131  & ~\s14_msel_pri_out_reg[1]/NET0131  ;
  assign n14314 = \s14_msel_arb0_state_reg[2]/NET0131  & n14313 ;
  assign n14315 = ~n14312 & ~n14314 ;
  assign n14316 = n14310 & n14315 ;
  assign n14317 = \s14_msel_arb2_state_reg[1]/NET0131  & n14308 ;
  assign n14318 = \s14_msel_arb1_state_reg[1]/NET0131  & n14306 ;
  assign n14319 = ~n14317 & ~n14318 ;
  assign n14320 = \s14_msel_arb3_state_reg[1]/NET0131  & n14311 ;
  assign n14321 = \s14_msel_arb0_state_reg[1]/NET0131  & n14313 ;
  assign n14322 = ~n14320 & ~n14321 ;
  assign n14323 = n14319 & n14322 ;
  assign n14324 = n14316 & n14323 ;
  assign n14325 = \s14_msel_arb2_state_reg[0]/NET0131  & n14308 ;
  assign n14326 = \s14_msel_arb1_state_reg[0]/NET0131  & n14306 ;
  assign n14327 = ~n14325 & ~n14326 ;
  assign n14328 = \s14_msel_arb3_state_reg[0]/NET0131  & n14311 ;
  assign n14329 = \s14_msel_arb0_state_reg[0]/NET0131  & n14313 ;
  assign n14330 = ~n14328 & ~n14329 ;
  assign n14331 = n14327 & n14330 ;
  assign n14332 = \m1_s14_cyc_o_reg/NET0131  & \s14_m1_cyc_r_reg/P0001  ;
  assign n14333 = ~n14331 & n14332 ;
  assign n14334 = n14324 & n14333 ;
  assign n14335 = \m0_s14_cyc_o_reg/NET0131  & \s14_m0_cyc_r_reg/P0001  ;
  assign n14336 = n14331 & n14335 ;
  assign n14337 = n14324 & n14336 ;
  assign n14338 = ~n14334 & ~n14337 ;
  assign n14339 = n14316 & ~n14323 ;
  assign n14340 = \m3_s14_cyc_o_reg/NET0131  & \s14_m3_cyc_r_reg/P0001  ;
  assign n14341 = ~n14331 & n14340 ;
  assign n14342 = n14339 & n14341 ;
  assign n14343 = \m2_s14_cyc_o_reg/NET0131  & \s14_m2_cyc_r_reg/P0001  ;
  assign n14344 = n14331 & n14343 ;
  assign n14345 = n14339 & n14344 ;
  assign n14346 = ~n14342 & ~n14345 ;
  assign n14347 = n14338 & n14346 ;
  assign n14348 = ~n14316 & ~n14323 ;
  assign n14349 = \m7_s14_cyc_o_reg/NET0131  & \s14_m7_cyc_r_reg/P0001  ;
  assign n14350 = ~n14331 & n14349 ;
  assign n14351 = n14348 & n14350 ;
  assign n14352 = \m6_s14_cyc_o_reg/NET0131  & \s14_m6_cyc_r_reg/P0001  ;
  assign n14353 = n14331 & n14352 ;
  assign n14354 = n14348 & n14353 ;
  assign n14355 = ~n14351 & ~n14354 ;
  assign n14356 = ~n14316 & n14323 ;
  assign n14357 = \m5_s14_cyc_o_reg/NET0131  & \s14_m5_cyc_r_reg/P0001  ;
  assign n14358 = ~n14331 & n14357 ;
  assign n14359 = n14356 & n14358 ;
  assign n14360 = \m4_s14_cyc_o_reg/NET0131  & \s14_m4_cyc_r_reg/P0001  ;
  assign n14361 = n14331 & n14360 ;
  assign n14362 = n14356 & n14361 ;
  assign n14363 = ~n14359 & ~n14362 ;
  assign n14364 = n14355 & n14363 ;
  assign n14365 = n14347 & n14364 ;
  assign n14366 = ~\s2_msel_pri_out_reg[0]/NET0131  & \s2_msel_pri_out_reg[1]/NET0131  ;
  assign n14367 = \s2_msel_arb2_state_reg[1]/NET0131  & n14366 ;
  assign n14368 = \s2_msel_pri_out_reg[0]/NET0131  & ~\s2_msel_pri_out_reg[1]/NET0131  ;
  assign n14369 = \s2_msel_arb1_state_reg[1]/NET0131  & n14368 ;
  assign n14370 = ~n14367 & ~n14369 ;
  assign n14371 = \s2_msel_pri_out_reg[0]/NET0131  & \s2_msel_pri_out_reg[1]/NET0131  ;
  assign n14372 = \s2_msel_arb3_state_reg[1]/NET0131  & n14371 ;
  assign n14373 = ~\s2_msel_pri_out_reg[0]/NET0131  & ~\s2_msel_pri_out_reg[1]/NET0131  ;
  assign n14374 = \s2_msel_arb0_state_reg[1]/NET0131  & n14373 ;
  assign n14375 = ~n14372 & ~n14374 ;
  assign n14376 = n14370 & n14375 ;
  assign n14377 = \s2_msel_arb1_state_reg[2]/NET0131  & n14368 ;
  assign n14378 = \s2_msel_arb2_state_reg[2]/NET0131  & n14366 ;
  assign n14379 = ~n14377 & ~n14378 ;
  assign n14380 = \s2_msel_arb3_state_reg[2]/NET0131  & n14371 ;
  assign n14381 = \s2_msel_arb0_state_reg[2]/NET0131  & n14373 ;
  assign n14382 = ~n14380 & ~n14381 ;
  assign n14383 = n14379 & n14382 ;
  assign n14384 = n14376 & ~n14383 ;
  assign n14385 = \s2_msel_arb2_state_reg[0]/NET0131  & n14366 ;
  assign n14386 = \s2_msel_arb1_state_reg[0]/NET0131  & n14368 ;
  assign n14387 = ~n14385 & ~n14386 ;
  assign n14388 = \s2_msel_arb3_state_reg[0]/NET0131  & n14371 ;
  assign n14389 = \s2_msel_arb0_state_reg[0]/NET0131  & n14373 ;
  assign n14390 = ~n14388 & ~n14389 ;
  assign n14391 = n14387 & n14390 ;
  assign n14392 = \m5_s2_cyc_o_reg/NET0131  & \s2_m5_cyc_r_reg/P0001  ;
  assign n14393 = ~n14391 & n14392 ;
  assign n14394 = n14384 & n14393 ;
  assign n14395 = \m4_s2_cyc_o_reg/NET0131  & \s2_m4_cyc_r_reg/P0001  ;
  assign n14396 = n14391 & n14395 ;
  assign n14397 = n14384 & n14396 ;
  assign n14398 = ~n14394 & ~n14397 ;
  assign n14399 = n14376 & n14383 ;
  assign n14400 = \m1_s2_cyc_o_reg/NET0131  & \s2_m1_cyc_r_reg/P0001  ;
  assign n14401 = ~n14391 & n14400 ;
  assign n14402 = n14399 & n14401 ;
  assign n14403 = \m0_s2_cyc_o_reg/NET0131  & \s2_m0_cyc_r_reg/P0001  ;
  assign n14404 = n14391 & n14403 ;
  assign n14405 = n14399 & n14404 ;
  assign n14406 = ~n14402 & ~n14405 ;
  assign n14407 = n14398 & n14406 ;
  assign n14408 = ~n14376 & ~n14383 ;
  assign n14409 = \m7_s2_cyc_o_reg/NET0131  & \s2_m7_cyc_r_reg/P0001  ;
  assign n14410 = ~n14391 & n14409 ;
  assign n14411 = n14408 & n14410 ;
  assign n14412 = \m6_s2_cyc_o_reg/NET0131  & \s2_m6_cyc_r_reg/P0001  ;
  assign n14413 = n14391 & n14412 ;
  assign n14414 = n14408 & n14413 ;
  assign n14415 = ~n14411 & ~n14414 ;
  assign n14416 = ~n14376 & n14383 ;
  assign n14417 = \m3_s2_cyc_o_reg/NET0131  & \s2_m3_cyc_r_reg/P0001  ;
  assign n14418 = ~n14391 & n14417 ;
  assign n14419 = n14416 & n14418 ;
  assign n14420 = \m2_s2_cyc_o_reg/NET0131  & \s2_m2_cyc_r_reg/P0001  ;
  assign n14421 = n14391 & n14420 ;
  assign n14422 = n14416 & n14421 ;
  assign n14423 = ~n14419 & ~n14422 ;
  assign n14424 = n14415 & n14423 ;
  assign n14425 = n14407 & n14424 ;
  assign n14426 = ~\s3_msel_pri_out_reg[0]/NET0131  & \s3_msel_pri_out_reg[1]/NET0131  ;
  assign n14427 = \s3_msel_arb2_state_reg[1]/NET0131  & n14426 ;
  assign n14428 = \s3_msel_pri_out_reg[0]/NET0131  & ~\s3_msel_pri_out_reg[1]/NET0131  ;
  assign n14429 = \s3_msel_arb1_state_reg[1]/NET0131  & n14428 ;
  assign n14430 = ~n14427 & ~n14429 ;
  assign n14431 = \s3_msel_pri_out_reg[0]/NET0131  & \s3_msel_pri_out_reg[1]/NET0131  ;
  assign n14432 = \s3_msel_arb3_state_reg[1]/NET0131  & n14431 ;
  assign n14433 = ~\s3_msel_pri_out_reg[0]/NET0131  & ~\s3_msel_pri_out_reg[1]/NET0131  ;
  assign n14434 = \s3_msel_arb0_state_reg[1]/NET0131  & n14433 ;
  assign n14435 = ~n14432 & ~n14434 ;
  assign n14436 = n14430 & n14435 ;
  assign n14437 = \s3_msel_arb2_state_reg[2]/NET0131  & n14426 ;
  assign n14438 = \s3_msel_arb1_state_reg[2]/NET0131  & n14428 ;
  assign n14439 = ~n14437 & ~n14438 ;
  assign n14440 = \s3_msel_arb3_state_reg[2]/NET0131  & n14431 ;
  assign n14441 = \s3_msel_arb0_state_reg[2]/NET0131  & n14433 ;
  assign n14442 = ~n14440 & ~n14441 ;
  assign n14443 = n14439 & n14442 ;
  assign n14444 = n14436 & ~n14443 ;
  assign n14445 = \s3_msel_arb2_state_reg[0]/NET0131  & n14426 ;
  assign n14446 = \s3_msel_arb1_state_reg[0]/NET0131  & n14428 ;
  assign n14447 = ~n14445 & ~n14446 ;
  assign n14448 = \s3_msel_arb3_state_reg[0]/NET0131  & n14431 ;
  assign n14449 = \s3_msel_arb0_state_reg[0]/NET0131  & n14433 ;
  assign n14450 = ~n14448 & ~n14449 ;
  assign n14451 = n14447 & n14450 ;
  assign n14452 = \m5_s3_cyc_o_reg/NET0131  & \s3_m5_cyc_r_reg/P0001  ;
  assign n14453 = ~n14451 & n14452 ;
  assign n14454 = n14444 & n14453 ;
  assign n14455 = \m4_s3_cyc_o_reg/NET0131  & \s3_m4_cyc_r_reg/P0001  ;
  assign n14456 = n14451 & n14455 ;
  assign n14457 = n14444 & n14456 ;
  assign n14458 = ~n14454 & ~n14457 ;
  assign n14459 = ~n14436 & n14443 ;
  assign n14460 = \m3_s3_cyc_o_reg/NET0131  & \s3_m3_cyc_r_reg/P0001  ;
  assign n14461 = ~n14451 & n14460 ;
  assign n14462 = n14459 & n14461 ;
  assign n14463 = \m2_s3_cyc_o_reg/NET0131  & \s3_m2_cyc_r_reg/P0001  ;
  assign n14464 = n14451 & n14463 ;
  assign n14465 = n14459 & n14464 ;
  assign n14466 = ~n14462 & ~n14465 ;
  assign n14467 = n14458 & n14466 ;
  assign n14468 = ~n14436 & ~n14443 ;
  assign n14469 = \m7_s3_cyc_o_reg/NET0131  & \s3_m7_cyc_r_reg/P0001  ;
  assign n14470 = ~n14451 & n14469 ;
  assign n14471 = n14468 & n14470 ;
  assign n14472 = \m6_s3_cyc_o_reg/NET0131  & \s3_m6_cyc_r_reg/P0001  ;
  assign n14473 = n14451 & n14472 ;
  assign n14474 = n14468 & n14473 ;
  assign n14475 = ~n14471 & ~n14474 ;
  assign n14476 = n14436 & n14443 ;
  assign n14477 = \m1_s3_cyc_o_reg/NET0131  & \s3_m1_cyc_r_reg/P0001  ;
  assign n14478 = ~n14451 & n14477 ;
  assign n14479 = n14476 & n14478 ;
  assign n14480 = \m0_s3_cyc_o_reg/NET0131  & \s3_m0_cyc_r_reg/P0001  ;
  assign n14481 = n14451 & n14480 ;
  assign n14482 = n14476 & n14481 ;
  assign n14483 = ~n14479 & ~n14482 ;
  assign n14484 = n14475 & n14483 ;
  assign n14485 = n14467 & n14484 ;
  assign n14486 = \s0_next_reg/P0001  & n4164 ;
  assign n14487 = n4181 & n14486 ;
  assign n14488 = n5446 & n5449 ;
  assign n14489 = n5458 & n14488 ;
  assign n14490 = n14487 & ~n14489 ;
  assign n14491 = \s0_msel_pri_out_reg[0]/NET0131  & ~\s0_next_reg/P0001  ;
  assign n14492 = n4850 & n4855 ;
  assign n14493 = \s0_next_reg/P0001  & ~n14492 ;
  assign n14494 = ~n14491 & ~n14493 ;
  assign n14495 = ~n14490 & n14494 ;
  assign n14496 = ~rst_i_pad & ~n14495 ;
  assign n14497 = n13504 & n13507 ;
  assign n14498 = ~\s10_msel_pri_out_reg[1]/NET0131  & ~\s10_next_reg/P0001  ;
  assign n14499 = ~rst_i_pad & ~n14498 ;
  assign n14500 = ~n14497 & n14499 ;
  assign n14501 = n13514 & n13517 ;
  assign n14502 = ~\s11_msel_pri_out_reg[1]/NET0131  & ~\s11_next_reg/P0001  ;
  assign n14503 = ~rst_i_pad & ~n14502 ;
  assign n14504 = ~n14501 & n14503 ;
  assign n14505 = n13584 & n13587 ;
  assign n14506 = ~\s12_msel_pri_out_reg[1]/NET0131  & ~\s12_next_reg/P0001  ;
  assign n14507 = ~rst_i_pad & ~n14506 ;
  assign n14508 = ~n14505 & n14507 ;
  assign n14509 = n13594 & n13597 ;
  assign n14510 = ~\s13_msel_pri_out_reg[1]/NET0131  & ~\s13_next_reg/P0001  ;
  assign n14511 = ~rst_i_pad & ~n14510 ;
  assign n14512 = ~n14509 & n14511 ;
  assign n14513 = n13664 & n13667 ;
  assign n14514 = ~\s14_msel_pri_out_reg[1]/NET0131  & ~\s14_next_reg/P0001  ;
  assign n14515 = ~rst_i_pad & ~n14514 ;
  assign n14516 = ~n14513 & n14515 ;
  assign n14517 = n13734 & n13737 ;
  assign n14518 = ~\s1_msel_pri_out_reg[1]/NET0131  & ~\s1_next_reg/P0001  ;
  assign n14519 = ~rst_i_pad & ~n14518 ;
  assign n14520 = ~n14517 & n14519 ;
  assign n14521 = n13804 & n13807 ;
  assign n14522 = ~\s2_msel_pri_out_reg[1]/NET0131  & ~\s2_next_reg/P0001  ;
  assign n14523 = ~rst_i_pad & ~n14522 ;
  assign n14524 = ~n14521 & n14523 ;
  assign n14525 = n13814 & n13817 ;
  assign n14526 = ~\s3_msel_pri_out_reg[1]/NET0131  & ~\s3_next_reg/P0001  ;
  assign n14527 = ~rst_i_pad & ~n14526 ;
  assign n14528 = ~n14525 & n14527 ;
  assign n14529 = n13884 & n13887 ;
  assign n14530 = ~\s4_msel_pri_out_reg[1]/NET0131  & ~\s4_next_reg/P0001  ;
  assign n14531 = ~rst_i_pad & ~n14530 ;
  assign n14532 = ~n14529 & n14531 ;
  assign n14533 = n13893 & n13898 ;
  assign n14534 = ~\s5_msel_pri_out_reg[1]/NET0131  & ~\s5_next_reg/P0001  ;
  assign n14535 = ~rst_i_pad & ~n14534 ;
  assign n14536 = ~n14533 & n14535 ;
  assign n14537 = n13964 & n13969 ;
  assign n14538 = ~\s6_msel_pri_out_reg[1]/NET0131  & ~\s6_next_reg/P0001  ;
  assign n14539 = ~rst_i_pad & ~n14538 ;
  assign n14540 = ~n14537 & n14539 ;
  assign n14541 = n13976 & n13979 ;
  assign n14542 = ~\s7_msel_pri_out_reg[1]/NET0131  & ~\s7_next_reg/P0001  ;
  assign n14543 = ~rst_i_pad & ~n14542 ;
  assign n14544 = ~n14541 & n14543 ;
  assign n14545 = n14105 & n14110 ;
  assign n14546 = ~\s8_msel_pri_out_reg[1]/NET0131  & ~\s8_next_reg/P0001  ;
  assign n14547 = ~rst_i_pad & ~n14546 ;
  assign n14548 = ~n14545 & n14547 ;
  assign n14549 = n14176 & n14180 ;
  assign n14550 = ~\s9_msel_pri_out_reg[1]/NET0131  & ~\s9_next_reg/P0001  ;
  assign n14551 = ~rst_i_pad & ~n14550 ;
  assign n14552 = ~n14549 & n14551 ;
  assign n14553 = n14487 & n14492 ;
  assign n14554 = ~\s0_msel_pri_out_reg[1]/NET0131  & ~\s0_next_reg/P0001  ;
  assign n14555 = ~rst_i_pad & ~n14554 ;
  assign n14556 = ~n14553 & n14555 ;
  assign n14557 = \m5_cyc_i_pad  & ~\m5_stb_i_pad  ;
  assign n14558 = \m5_s1_cyc_o_reg/NET0131  & n14557 ;
  assign n14559 = ~\m5_addr_i[30]_pad  & ~\m5_addr_i[31]_pad  ;
  assign n14560 = \m5_addr_i[28]_pad  & ~\m5_addr_i[29]_pad  ;
  assign n14561 = n14559 & n14560 ;
  assign n14562 = \m5_cyc_i_pad  & \m5_stb_i_pad  ;
  assign n14563 = n14561 & n14562 ;
  assign n14564 = ~n14558 & ~n14563 ;
  assign n14565 = \m0_cyc_i_pad  & ~\m0_stb_i_pad  ;
  assign n14566 = \m0_s0_cyc_o_reg/NET0131  & n14565 ;
  assign n14567 = ~\m0_addr_i[29]_pad  & ~\m0_addr_i[31]_pad  ;
  assign n14568 = ~\m0_addr_i[28]_pad  & ~\m0_addr_i[30]_pad  ;
  assign n14569 = n14567 & n14568 ;
  assign n14570 = \m0_cyc_i_pad  & \m0_stb_i_pad  ;
  assign n14571 = n14569 & n14570 ;
  assign n14572 = ~n14566 & ~n14571 ;
  assign n14573 = \m0_s1_cyc_o_reg/NET0131  & n14565 ;
  assign n14574 = \m0_addr_i[28]_pad  & ~\m0_addr_i[30]_pad  ;
  assign n14575 = n14567 & n14574 ;
  assign n14576 = n14570 & n14575 ;
  assign n14577 = ~n14573 & ~n14576 ;
  assign n14578 = \m1_cyc_i_pad  & ~\m1_stb_i_pad  ;
  assign n14579 = \m1_s0_cyc_o_reg/NET0131  & n14578 ;
  assign n14580 = ~\m1_addr_i[30]_pad  & ~\m1_addr_i[31]_pad  ;
  assign n14581 = ~\m1_addr_i[28]_pad  & ~\m1_addr_i[29]_pad  ;
  assign n14582 = n14580 & n14581 ;
  assign n14583 = \m1_cyc_i_pad  & \m1_stb_i_pad  ;
  assign n14584 = n14582 & n14583 ;
  assign n14585 = ~n14579 & ~n14584 ;
  assign n14586 = \m2_cyc_i_pad  & ~\m2_stb_i_pad  ;
  assign n14587 = \m2_s0_cyc_o_reg/NET0131  & n14586 ;
  assign n14588 = ~\m2_addr_i[28]_pad  & ~\m2_addr_i[29]_pad  ;
  assign n14589 = ~\m2_addr_i[30]_pad  & ~\m2_addr_i[31]_pad  ;
  assign n14590 = n14588 & n14589 ;
  assign n14591 = \m2_cyc_i_pad  & \m2_stb_i_pad  ;
  assign n14592 = n14590 & n14591 ;
  assign n14593 = ~n14587 & ~n14592 ;
  assign n14594 = \m2_s1_cyc_o_reg/NET0131  & n14586 ;
  assign n14595 = \m2_addr_i[28]_pad  & ~\m2_addr_i[29]_pad  ;
  assign n14596 = n14589 & n14595 ;
  assign n14597 = n14591 & n14596 ;
  assign n14598 = ~n14594 & ~n14597 ;
  assign n14599 = \m3_cyc_i_pad  & ~\m3_stb_i_pad  ;
  assign n14600 = \m3_s0_cyc_o_reg/NET0131  & n14599 ;
  assign n14601 = ~\m3_addr_i[30]_pad  & ~\m3_addr_i[31]_pad  ;
  assign n14602 = ~\m3_addr_i[28]_pad  & ~\m3_addr_i[29]_pad  ;
  assign n14603 = n14601 & n14602 ;
  assign n14604 = \m3_cyc_i_pad  & \m3_stb_i_pad  ;
  assign n14605 = n14603 & n14604 ;
  assign n14606 = ~n14600 & ~n14605 ;
  assign n14607 = \m3_s1_cyc_o_reg/NET0131  & n14599 ;
  assign n14608 = \m3_addr_i[28]_pad  & ~\m3_addr_i[29]_pad  ;
  assign n14609 = n14601 & n14608 ;
  assign n14610 = n14604 & n14609 ;
  assign n14611 = ~n14607 & ~n14610 ;
  assign n14612 = \m4_cyc_i_pad  & ~\m4_stb_i_pad  ;
  assign n14613 = \m4_s0_cyc_o_reg/NET0131  & n14612 ;
  assign n14614 = ~\m4_addr_i[30]_pad  & ~\m4_addr_i[31]_pad  ;
  assign n14615 = ~\m4_addr_i[28]_pad  & ~\m4_addr_i[29]_pad  ;
  assign n14616 = n14614 & n14615 ;
  assign n14617 = \m4_cyc_i_pad  & \m4_stb_i_pad  ;
  assign n14618 = n14616 & n14617 ;
  assign n14619 = ~n14613 & ~n14618 ;
  assign n14620 = \m4_s1_cyc_o_reg/NET0131  & n14612 ;
  assign n14621 = \m4_addr_i[28]_pad  & ~\m4_addr_i[29]_pad  ;
  assign n14622 = n14614 & n14621 ;
  assign n14623 = n14617 & n14622 ;
  assign n14624 = ~n14620 & ~n14623 ;
  assign n14625 = \m5_s0_cyc_o_reg/NET0131  & n14557 ;
  assign n14626 = ~\m5_addr_i[28]_pad  & ~\m5_addr_i[29]_pad  ;
  assign n14627 = n14559 & n14626 ;
  assign n14628 = n14562 & n14627 ;
  assign n14629 = ~n14625 & ~n14628 ;
  assign n14630 = \m6_cyc_i_pad  & ~\m6_stb_i_pad  ;
  assign n14631 = \m6_s0_cyc_o_reg/NET0131  & n14630 ;
  assign n14632 = ~\m6_addr_i[30]_pad  & ~\m6_addr_i[31]_pad  ;
  assign n14633 = ~\m6_addr_i[28]_pad  & ~\m6_addr_i[29]_pad  ;
  assign n14634 = n14632 & n14633 ;
  assign n14635 = \m6_cyc_i_pad  & \m6_stb_i_pad  ;
  assign n14636 = n14634 & n14635 ;
  assign n14637 = ~n14631 & ~n14636 ;
  assign n14638 = \m6_s1_cyc_o_reg/NET0131  & n14630 ;
  assign n14639 = \m6_addr_i[28]_pad  & ~\m6_addr_i[29]_pad  ;
  assign n14640 = n14632 & n14639 ;
  assign n14641 = n14635 & n14640 ;
  assign n14642 = ~n14638 & ~n14641 ;
  assign n14643 = \m7_cyc_i_pad  & ~\m7_stb_i_pad  ;
  assign n14644 = \m7_s0_cyc_o_reg/NET0131  & n14643 ;
  assign n14645 = ~\m7_addr_i[30]_pad  & ~\m7_addr_i[31]_pad  ;
  assign n14646 = ~\m7_addr_i[28]_pad  & ~\m7_addr_i[29]_pad  ;
  assign n14647 = n14645 & n14646 ;
  assign n14648 = \m7_cyc_i_pad  & \m7_stb_i_pad  ;
  assign n14649 = n14647 & n14648 ;
  assign n14650 = ~n14644 & ~n14649 ;
  assign n14651 = \m7_s1_cyc_o_reg/NET0131  & n14643 ;
  assign n14652 = \m7_addr_i[28]_pad  & ~\m7_addr_i[29]_pad  ;
  assign n14653 = n14645 & n14652 ;
  assign n14654 = n14648 & n14653 ;
  assign n14655 = ~n14651 & ~n14654 ;
  assign n14656 = \m1_s1_cyc_o_reg/NET0131  & n14578 ;
  assign n14657 = \m1_addr_i[28]_pad  & ~\m1_addr_i[29]_pad  ;
  assign n14658 = n14580 & n14657 ;
  assign n14659 = n14583 & n14658 ;
  assign n14660 = ~n14656 & ~n14659 ;
  assign n14661 = \m5_s15_cyc_o_reg/NET0131  & n14557 ;
  assign n14662 = n2203 & n14562 ;
  assign n14663 = ~n14661 & ~n14662 ;
  assign n14664 = \m7_s9_cyc_o_reg/NET0131  & n14643 ;
  assign n14665 = ~\m7_addr_i[30]_pad  & \m7_addr_i[31]_pad  ;
  assign n14666 = n14652 & n14665 ;
  assign n14667 = n14648 & n14666 ;
  assign n14668 = ~n14664 & ~n14667 ;
  assign n14669 = \m7_s7_cyc_o_reg/NET0131  & n14643 ;
  assign n14670 = \m7_addr_i[30]_pad  & ~\m7_addr_i[31]_pad  ;
  assign n14671 = n2169 & n14670 ;
  assign n14672 = n14648 & n14671 ;
  assign n14673 = ~n14669 & ~n14672 ;
  assign n14674 = \m7_s5_cyc_o_reg/NET0131  & n14643 ;
  assign n14675 = n14652 & n14670 ;
  assign n14676 = n14648 & n14675 ;
  assign n14677 = ~n14674 & ~n14676 ;
  assign n14678 = \m6_s6_cyc_o_reg/NET0131  & n14630 ;
  assign n14679 = \m6_addr_i[30]_pad  & ~\m6_addr_i[31]_pad  ;
  assign n14680 = ~\m6_addr_i[28]_pad  & \m6_addr_i[29]_pad  ;
  assign n14681 = n14679 & n14680 ;
  assign n14682 = n14635 & n14681 ;
  assign n14683 = ~n14678 & ~n14682 ;
  assign n14684 = \m7_s12_cyc_o_reg/NET0131  & n14643 ;
  assign n14685 = n2168 & n14646 ;
  assign n14686 = n14648 & n14685 ;
  assign n14687 = ~n14684 & ~n14686 ;
  assign n14688 = \m6_s8_cyc_o_reg/NET0131  & n14630 ;
  assign n14689 = ~\m6_addr_i[30]_pad  & \m6_addr_i[31]_pad  ;
  assign n14690 = n14633 & n14689 ;
  assign n14691 = n14635 & n14690 ;
  assign n14692 = ~n14688 & ~n14691 ;
  assign n14693 = \m5_s7_cyc_o_reg/NET0131  & n14557 ;
  assign n14694 = \m5_addr_i[30]_pad  & ~\m5_addr_i[31]_pad  ;
  assign n14695 = n2201 & n14694 ;
  assign n14696 = n14562 & n14695 ;
  assign n14697 = ~n14693 & ~n14696 ;
  assign n14698 = \m5_s14_cyc_o_reg/NET0131  & n14557 ;
  assign n14699 = ~\m5_addr_i[28]_pad  & \m5_addr_i[29]_pad  ;
  assign n14700 = n2202 & n14699 ;
  assign n14701 = n14562 & n14700 ;
  assign n14702 = ~n14698 & ~n14701 ;
  assign n14703 = \m5_s3_cyc_o_reg/NET0131  & n14557 ;
  assign n14704 = n2201 & n14559 ;
  assign n14705 = n14562 & n14704 ;
  assign n14706 = ~n14703 & ~n14705 ;
  assign n14707 = \m5_s12_cyc_o_reg/NET0131  & n14557 ;
  assign n14708 = n2202 & n14626 ;
  assign n14709 = n14562 & n14708 ;
  assign n14710 = ~n14707 & ~n14709 ;
  assign n14711 = \m4_s9_cyc_o_reg/NET0131  & n14612 ;
  assign n14712 = ~\m4_addr_i[30]_pad  & \m4_addr_i[31]_pad  ;
  assign n14713 = n14621 & n14712 ;
  assign n14714 = n14617 & n14713 ;
  assign n14715 = ~n14711 & ~n14714 ;
  assign n14716 = \m4_s8_cyc_o_reg/NET0131  & n14612 ;
  assign n14717 = n14615 & n14712 ;
  assign n14718 = n14617 & n14717 ;
  assign n14719 = ~n14716 & ~n14718 ;
  assign n14720 = \m4_s6_cyc_o_reg/NET0131  & n14612 ;
  assign n14721 = \m4_addr_i[30]_pad  & ~\m4_addr_i[31]_pad  ;
  assign n14722 = ~\m4_addr_i[28]_pad  & \m4_addr_i[29]_pad  ;
  assign n14723 = n14721 & n14722 ;
  assign n14724 = n14617 & n14723 ;
  assign n14725 = ~n14720 & ~n14724 ;
  assign n14726 = \m4_s4_cyc_o_reg/NET0131  & n14612 ;
  assign n14727 = n14615 & n14721 ;
  assign n14728 = n14617 & n14727 ;
  assign n14729 = ~n14726 & ~n14728 ;
  assign n14730 = \m4_s13_cyc_o_reg/NET0131  & n14612 ;
  assign n14731 = n2196 & n14621 ;
  assign n14732 = n14617 & n14731 ;
  assign n14733 = ~n14730 & ~n14732 ;
  assign n14734 = \m4_s11_cyc_o_reg/NET0131  & n14612 ;
  assign n14735 = n2195 & n14712 ;
  assign n14736 = n14617 & n14735 ;
  assign n14737 = ~n14734 & ~n14736 ;
  assign n14738 = \m3_s7_cyc_o_reg/NET0131  & n14599 ;
  assign n14739 = \m3_addr_i[30]_pad  & ~\m3_addr_i[31]_pad  ;
  assign n14740 = n2188 & n14739 ;
  assign n14741 = n14604 & n14740 ;
  assign n14742 = ~n14738 & ~n14741 ;
  assign n14743 = \m3_s6_cyc_o_reg/NET0131  & n14599 ;
  assign n14744 = ~\m3_addr_i[28]_pad  & \m3_addr_i[29]_pad  ;
  assign n14745 = n14739 & n14744 ;
  assign n14746 = n14604 & n14745 ;
  assign n14747 = ~n14743 & ~n14746 ;
  assign n14748 = \m0_s10_cyc_o_reg/NET0131  & n14565 ;
  assign n14749 = n2161 & n14568 ;
  assign n14750 = n14570 & n14749 ;
  assign n14751 = ~n14748 & ~n14750 ;
  assign n14752 = \m0_s11_cyc_o_reg/NET0131  & n14565 ;
  assign n14753 = n2161 & n14574 ;
  assign n14754 = n14570 & n14753 ;
  assign n14755 = ~n14752 & ~n14754 ;
  assign n14756 = \m3_s5_cyc_o_reg/NET0131  & n14599 ;
  assign n14757 = n14608 & n14739 ;
  assign n14758 = n14604 & n14757 ;
  assign n14759 = ~n14756 & ~n14758 ;
  assign n14760 = \m0_s14_cyc_o_reg/NET0131  & n14565 ;
  assign n14761 = ~\m0_addr_i[28]_pad  & \m0_addr_i[30]_pad  ;
  assign n14762 = n2161 & n14761 ;
  assign n14763 = n14570 & n14762 ;
  assign n14764 = ~n14760 & ~n14763 ;
  assign n14765 = \m0_s15_cyc_o_reg/NET0131  & n14565 ;
  assign n14766 = n2163 & n14570 ;
  assign n14767 = ~n14765 & ~n14766 ;
  assign n14768 = \m0_s2_cyc_o_reg/NET0131  & n14565 ;
  assign n14769 = \m0_addr_i[29]_pad  & ~\m0_addr_i[31]_pad  ;
  assign n14770 = n14568 & n14769 ;
  assign n14771 = n14570 & n14770 ;
  assign n14772 = ~n14768 & ~n14771 ;
  assign n14773 = \m0_s3_cyc_o_reg/NET0131  & n14565 ;
  assign n14774 = n14574 & n14769 ;
  assign n14775 = n14570 & n14774 ;
  assign n14776 = ~n14773 & ~n14775 ;
  assign n14777 = \m0_s5_cyc_o_reg/NET0131  & n14565 ;
  assign n14778 = n2162 & n14567 ;
  assign n14779 = n14570 & n14778 ;
  assign n14780 = ~n14777 & ~n14779 ;
  assign n14781 = \m0_s6_cyc_o_reg/NET0131  & n14565 ;
  assign n14782 = n14761 & n14769 ;
  assign n14783 = n14570 & n14782 ;
  assign n14784 = ~n14781 & ~n14783 ;
  assign n14785 = \m0_s7_cyc_o_reg/NET0131  & n14565 ;
  assign n14786 = n2162 & n14769 ;
  assign n14787 = n14570 & n14786 ;
  assign n14788 = ~n14785 & ~n14787 ;
  assign n14789 = \m0_s8_cyc_o_reg/NET0131  & n14565 ;
  assign n14790 = ~\m0_addr_i[29]_pad  & \m0_addr_i[31]_pad  ;
  assign n14791 = n14568 & n14790 ;
  assign n14792 = n14570 & n14791 ;
  assign n14793 = ~n14789 & ~n14792 ;
  assign n14794 = \m1_s10_cyc_o_reg/NET0131  & n14578 ;
  assign n14795 = ~\m1_addr_i[30]_pad  & \m1_addr_i[31]_pad  ;
  assign n14796 = ~\m1_addr_i[28]_pad  & \m1_addr_i[29]_pad  ;
  assign n14797 = n14795 & n14796 ;
  assign n14798 = n14583 & n14797 ;
  assign n14799 = ~n14794 & ~n14798 ;
  assign n14800 = \m3_s3_cyc_o_reg/NET0131  & n14599 ;
  assign n14801 = n2188 & n14601 ;
  assign n14802 = n14604 & n14801 ;
  assign n14803 = ~n14800 & ~n14802 ;
  assign n14804 = \m1_s13_cyc_o_reg/NET0131  & n14578 ;
  assign n14805 = n2156 & n14657 ;
  assign n14806 = n14583 & n14805 ;
  assign n14807 = ~n14804 & ~n14806 ;
  assign n14808 = \m1_s14_cyc_o_reg/NET0131  & n14578 ;
  assign n14809 = n2156 & n14796 ;
  assign n14810 = n14583 & n14809 ;
  assign n14811 = ~n14808 & ~n14810 ;
  assign n14812 = \m1_s15_cyc_o_reg/NET0131  & n14578 ;
  assign n14813 = n2157 & n14583 ;
  assign n14814 = ~n14812 & ~n14813 ;
  assign n14815 = \m1_s2_cyc_o_reg/NET0131  & n14578 ;
  assign n14816 = n14580 & n14796 ;
  assign n14817 = n14583 & n14816 ;
  assign n14818 = ~n14815 & ~n14817 ;
  assign n14819 = \m1_s3_cyc_o_reg/NET0131  & n14578 ;
  assign n14820 = n2155 & n14580 ;
  assign n14821 = n14583 & n14820 ;
  assign n14822 = ~n14819 & ~n14821 ;
  assign n14823 = \m1_s4_cyc_o_reg/NET0131  & n14578 ;
  assign n14824 = \m1_addr_i[30]_pad  & ~\m1_addr_i[31]_pad  ;
  assign n14825 = n14581 & n14824 ;
  assign n14826 = n14583 & n14825 ;
  assign n14827 = ~n14823 & ~n14826 ;
  assign n14828 = \m1_s5_cyc_o_reg/NET0131  & n14578 ;
  assign n14829 = n14657 & n14824 ;
  assign n14830 = n14583 & n14829 ;
  assign n14831 = ~n14828 & ~n14830 ;
  assign n14832 = \m1_s6_cyc_o_reg/NET0131  & n14578 ;
  assign n14833 = n14796 & n14824 ;
  assign n14834 = n14583 & n14833 ;
  assign n14835 = ~n14832 & ~n14834 ;
  assign n14836 = \m1_s7_cyc_o_reg/NET0131  & n14578 ;
  assign n14837 = n2155 & n14824 ;
  assign n14838 = n14583 & n14837 ;
  assign n14839 = ~n14836 & ~n14838 ;
  assign n14840 = \m1_s8_cyc_o_reg/NET0131  & n14578 ;
  assign n14841 = n14581 & n14795 ;
  assign n14842 = n14583 & n14841 ;
  assign n14843 = ~n14840 & ~n14842 ;
  assign n14844 = \m1_s9_cyc_o_reg/NET0131  & n14578 ;
  assign n14845 = n14657 & n14795 ;
  assign n14846 = n14583 & n14845 ;
  assign n14847 = ~n14844 & ~n14846 ;
  assign n14848 = \m2_s10_cyc_o_reg/NET0131  & n14586 ;
  assign n14849 = ~\m2_addr_i[30]_pad  & \m2_addr_i[31]_pad  ;
  assign n14850 = ~\m2_addr_i[28]_pad  & \m2_addr_i[29]_pad  ;
  assign n14851 = n14849 & n14850 ;
  assign n14852 = n14591 & n14851 ;
  assign n14853 = ~n14848 & ~n14852 ;
  assign n14854 = \m2_s11_cyc_o_reg/NET0131  & n14586 ;
  assign n14855 = n2182 & n14849 ;
  assign n14856 = n14591 & n14855 ;
  assign n14857 = ~n14854 & ~n14856 ;
  assign n14858 = \m2_s12_cyc_o_reg/NET0131  & n14586 ;
  assign n14859 = n2183 & n14588 ;
  assign n14860 = n14591 & n14859 ;
  assign n14861 = ~n14858 & ~n14860 ;
  assign n14862 = \m2_s15_cyc_o_reg/NET0131  & n14586 ;
  assign n14863 = n2184 & n14591 ;
  assign n14864 = ~n14862 & ~n14863 ;
  assign n14865 = \m2_s2_cyc_o_reg/NET0131  & n14586 ;
  assign n14866 = n14589 & n14850 ;
  assign n14867 = n14591 & n14866 ;
  assign n14868 = ~n14865 & ~n14867 ;
  assign n14869 = \m2_s3_cyc_o_reg/NET0131  & n14586 ;
  assign n14870 = n2182 & n14589 ;
  assign n14871 = n14591 & n14870 ;
  assign n14872 = ~n14869 & ~n14871 ;
  assign n14873 = \m2_s4_cyc_o_reg/NET0131  & n14586 ;
  assign n14874 = \m2_addr_i[30]_pad  & ~\m2_addr_i[31]_pad  ;
  assign n14875 = n14588 & n14874 ;
  assign n14876 = n14591 & n14875 ;
  assign n14877 = ~n14873 & ~n14876 ;
  assign n14878 = \m2_s5_cyc_o_reg/NET0131  & n14586 ;
  assign n14879 = n14595 & n14874 ;
  assign n14880 = n14591 & n14879 ;
  assign n14881 = ~n14878 & ~n14880 ;
  assign n14882 = \m2_s6_cyc_o_reg/NET0131  & n14586 ;
  assign n14883 = n14850 & n14874 ;
  assign n14884 = n14591 & n14883 ;
  assign n14885 = ~n14882 & ~n14884 ;
  assign n14886 = \m2_s9_cyc_o_reg/NET0131  & n14586 ;
  assign n14887 = n14595 & n14849 ;
  assign n14888 = n14591 & n14887 ;
  assign n14889 = ~n14886 & ~n14888 ;
  assign n14890 = \m3_s10_cyc_o_reg/NET0131  & n14599 ;
  assign n14891 = ~\m3_addr_i[30]_pad  & \m3_addr_i[31]_pad  ;
  assign n14892 = n14744 & n14891 ;
  assign n14893 = n14604 & n14892 ;
  assign n14894 = ~n14890 & ~n14893 ;
  assign n14895 = \m3_s11_cyc_o_reg/NET0131  & n14599 ;
  assign n14896 = n2188 & n14891 ;
  assign n14897 = n14604 & n14896 ;
  assign n14898 = ~n14895 & ~n14897 ;
  assign n14899 = \m3_s12_cyc_o_reg/NET0131  & n14599 ;
  assign n14900 = n2189 & n14602 ;
  assign n14901 = n14604 & n14900 ;
  assign n14902 = ~n14899 & ~n14901 ;
  assign n14903 = \m3_s13_cyc_o_reg/NET0131  & n14599 ;
  assign n14904 = n2189 & n14608 ;
  assign n14905 = n14604 & n14904 ;
  assign n14906 = ~n14903 & ~n14905 ;
  assign n14907 = \m3_s15_cyc_o_reg/NET0131  & n14599 ;
  assign n14908 = n2190 & n14604 ;
  assign n14909 = ~n14907 & ~n14908 ;
  assign n14910 = \m3_s2_cyc_o_reg/NET0131  & n14599 ;
  assign n14911 = n14601 & n14744 ;
  assign n14912 = n14604 & n14911 ;
  assign n14913 = ~n14910 & ~n14912 ;
  assign n14914 = \m3_s14_cyc_o_reg/NET0131  & n14599 ;
  assign n14915 = n2189 & n14744 ;
  assign n14916 = n14604 & n14915 ;
  assign n14917 = ~n14914 & ~n14916 ;
  assign n14918 = \m3_s4_cyc_o_reg/NET0131  & n14599 ;
  assign n14919 = n14602 & n14739 ;
  assign n14920 = n14604 & n14919 ;
  assign n14921 = ~n14918 & ~n14920 ;
  assign n14922 = \m3_s8_cyc_o_reg/NET0131  & n14599 ;
  assign n14923 = n14602 & n14891 ;
  assign n14924 = n14604 & n14923 ;
  assign n14925 = ~n14922 & ~n14924 ;
  assign n14926 = \m3_s9_cyc_o_reg/NET0131  & n14599 ;
  assign n14927 = n14608 & n14891 ;
  assign n14928 = n14604 & n14927 ;
  assign n14929 = ~n14926 & ~n14928 ;
  assign n14930 = \m4_s10_cyc_o_reg/NET0131  & n14612 ;
  assign n14931 = n14712 & n14722 ;
  assign n14932 = n14617 & n14931 ;
  assign n14933 = ~n14930 & ~n14932 ;
  assign n14934 = \m4_s12_cyc_o_reg/NET0131  & n14612 ;
  assign n14935 = n2196 & n14615 ;
  assign n14936 = n14617 & n14935 ;
  assign n14937 = ~n14934 & ~n14936 ;
  assign n14938 = \m4_s14_cyc_o_reg/NET0131  & n14612 ;
  assign n14939 = n2196 & n14722 ;
  assign n14940 = n14617 & n14939 ;
  assign n14941 = ~n14938 & ~n14940 ;
  assign n14942 = \m4_s15_cyc_o_reg/NET0131  & n14612 ;
  assign n14943 = n2197 & n14617 ;
  assign n14944 = ~n14942 & ~n14943 ;
  assign n14945 = \m4_s2_cyc_o_reg/NET0131  & n14612 ;
  assign n14946 = n14614 & n14722 ;
  assign n14947 = n14617 & n14946 ;
  assign n14948 = ~n14945 & ~n14947 ;
  assign n14949 = \m4_s3_cyc_o_reg/NET0131  & n14612 ;
  assign n14950 = n2195 & n14614 ;
  assign n14951 = n14617 & n14950 ;
  assign n14952 = ~n14949 & ~n14951 ;
  assign n14953 = \m4_s5_cyc_o_reg/NET0131  & n14612 ;
  assign n14954 = n14621 & n14721 ;
  assign n14955 = n14617 & n14954 ;
  assign n14956 = ~n14953 & ~n14955 ;
  assign n14957 = \m4_s7_cyc_o_reg/NET0131  & n14612 ;
  assign n14958 = n2195 & n14721 ;
  assign n14959 = n14617 & n14958 ;
  assign n14960 = ~n14957 & ~n14959 ;
  assign n14961 = \m5_s10_cyc_o_reg/NET0131  & n14557 ;
  assign n14962 = ~\m5_addr_i[30]_pad  & \m5_addr_i[31]_pad  ;
  assign n14963 = n14699 & n14962 ;
  assign n14964 = n14562 & n14963 ;
  assign n14965 = ~n14961 & ~n14964 ;
  assign n14966 = \m5_s11_cyc_o_reg/NET0131  & n14557 ;
  assign n14967 = n2201 & n14962 ;
  assign n14968 = n14562 & n14967 ;
  assign n14969 = ~n14966 & ~n14968 ;
  assign n14970 = \m5_s13_cyc_o_reg/NET0131  & n14557 ;
  assign n14971 = n2202 & n14560 ;
  assign n14972 = n14562 & n14971 ;
  assign n14973 = ~n14970 & ~n14972 ;
  assign n14974 = \m5_s2_cyc_o_reg/NET0131  & n14557 ;
  assign n14975 = n14559 & n14699 ;
  assign n14976 = n14562 & n14975 ;
  assign n14977 = ~n14974 & ~n14976 ;
  assign n14978 = \m5_s4_cyc_o_reg/NET0131  & n14557 ;
  assign n14979 = n14626 & n14694 ;
  assign n14980 = n14562 & n14979 ;
  assign n14981 = ~n14978 & ~n14980 ;
  assign n14982 = \m5_s5_cyc_o_reg/NET0131  & n14557 ;
  assign n14983 = n14560 & n14694 ;
  assign n14984 = n14562 & n14983 ;
  assign n14985 = ~n14982 & ~n14984 ;
  assign n14986 = \m5_s6_cyc_o_reg/NET0131  & n14557 ;
  assign n14987 = n14694 & n14699 ;
  assign n14988 = n14562 & n14987 ;
  assign n14989 = ~n14986 & ~n14988 ;
  assign n14990 = \m5_s8_cyc_o_reg/NET0131  & n14557 ;
  assign n14991 = n14626 & n14962 ;
  assign n14992 = n14562 & n14991 ;
  assign n14993 = ~n14990 & ~n14992 ;
  assign n14994 = \m5_s9_cyc_o_reg/NET0131  & n14557 ;
  assign n14995 = n14560 & n14962 ;
  assign n14996 = n14562 & n14995 ;
  assign n14997 = ~n14994 & ~n14996 ;
  assign n14998 = \m6_s10_cyc_o_reg/NET0131  & n14630 ;
  assign n14999 = n14680 & n14689 ;
  assign n15000 = n14635 & n14999 ;
  assign n15001 = ~n14998 & ~n15000 ;
  assign n15002 = \m6_s11_cyc_o_reg/NET0131  & n14630 ;
  assign n15003 = n2174 & n14689 ;
  assign n15004 = n14635 & n15003 ;
  assign n15005 = ~n15002 & ~n15004 ;
  assign n15006 = \m6_s12_cyc_o_reg/NET0131  & n14630 ;
  assign n15007 = n2175 & n14633 ;
  assign n15008 = n14635 & n15007 ;
  assign n15009 = ~n15006 & ~n15008 ;
  assign n15010 = \m6_s13_cyc_o_reg/NET0131  & n14630 ;
  assign n15011 = n2175 & n14639 ;
  assign n15012 = n14635 & n15011 ;
  assign n15013 = ~n15010 & ~n15012 ;
  assign n15014 = \m6_s14_cyc_o_reg/NET0131  & n14630 ;
  assign n15015 = n2175 & n14680 ;
  assign n15016 = n14635 & n15015 ;
  assign n15017 = ~n15014 & ~n15016 ;
  assign n15018 = \m6_s15_cyc_o_reg/NET0131  & n14630 ;
  assign n15019 = n2176 & n14635 ;
  assign n15020 = ~n15018 & ~n15019 ;
  assign n15021 = \m6_s2_cyc_o_reg/NET0131  & n14630 ;
  assign n15022 = n14632 & n14680 ;
  assign n15023 = n14635 & n15022 ;
  assign n15024 = ~n15021 & ~n15023 ;
  assign n15025 = \m6_s3_cyc_o_reg/NET0131  & n14630 ;
  assign n15026 = n2174 & n14632 ;
  assign n15027 = n14635 & n15026 ;
  assign n15028 = ~n15025 & ~n15027 ;
  assign n15029 = \m6_s4_cyc_o_reg/NET0131  & n14630 ;
  assign n15030 = n14633 & n14679 ;
  assign n15031 = n14635 & n15030 ;
  assign n15032 = ~n15029 & ~n15031 ;
  assign n15033 = \m6_s5_cyc_o_reg/NET0131  & n14630 ;
  assign n15034 = n14639 & n14679 ;
  assign n15035 = n14635 & n15034 ;
  assign n15036 = ~n15033 & ~n15035 ;
  assign n15037 = \m6_s7_cyc_o_reg/NET0131  & n14630 ;
  assign n15038 = n2174 & n14679 ;
  assign n15039 = n14635 & n15038 ;
  assign n15040 = ~n15037 & ~n15039 ;
  assign n15041 = \m6_s9_cyc_o_reg/NET0131  & n14630 ;
  assign n15042 = n14639 & n14689 ;
  assign n15043 = n14635 & n15042 ;
  assign n15044 = ~n15041 & ~n15043 ;
  assign n15045 = \m7_s10_cyc_o_reg/NET0131  & n14643 ;
  assign n15046 = ~\m7_addr_i[28]_pad  & \m7_addr_i[29]_pad  ;
  assign n15047 = n14665 & n15046 ;
  assign n15048 = n14648 & n15047 ;
  assign n15049 = ~n15045 & ~n15048 ;
  assign n15050 = \m7_s11_cyc_o_reg/NET0131  & n14643 ;
  assign n15051 = n2169 & n14665 ;
  assign n15052 = n14648 & n15051 ;
  assign n15053 = ~n15050 & ~n15052 ;
  assign n15054 = \m7_s13_cyc_o_reg/NET0131  & n14643 ;
  assign n15055 = n2168 & n14652 ;
  assign n15056 = n14648 & n15055 ;
  assign n15057 = ~n15054 & ~n15056 ;
  assign n15058 = \m7_s14_cyc_o_reg/NET0131  & n14643 ;
  assign n15059 = n2168 & n15046 ;
  assign n15060 = n14648 & n15059 ;
  assign n15061 = ~n15058 & ~n15060 ;
  assign n15062 = \m7_s15_cyc_o_reg/NET0131  & n14643 ;
  assign n15063 = n2170 & n14648 ;
  assign n15064 = ~n15062 & ~n15063 ;
  assign n15065 = \m7_s2_cyc_o_reg/NET0131  & n14643 ;
  assign n15066 = n14645 & n15046 ;
  assign n15067 = n14648 & n15066 ;
  assign n15068 = ~n15065 & ~n15067 ;
  assign n15069 = \m7_s3_cyc_o_reg/NET0131  & n14643 ;
  assign n15070 = n2169 & n14645 ;
  assign n15071 = n14648 & n15070 ;
  assign n15072 = ~n15069 & ~n15071 ;
  assign n15073 = \m7_s4_cyc_o_reg/NET0131  & n14643 ;
  assign n15074 = n14646 & n14670 ;
  assign n15075 = n14648 & n15074 ;
  assign n15076 = ~n15073 & ~n15075 ;
  assign n15077 = \m7_s6_cyc_o_reg/NET0131  & n14643 ;
  assign n15078 = n14670 & n15046 ;
  assign n15079 = n14648 & n15078 ;
  assign n15080 = ~n15077 & ~n15079 ;
  assign n15081 = \m2_s8_cyc_o_reg/NET0131  & n14586 ;
  assign n15082 = n14588 & n14849 ;
  assign n15083 = n14591 & n15082 ;
  assign n15084 = ~n15081 & ~n15083 ;
  assign n15085 = \m7_s8_cyc_o_reg/NET0131  & n14643 ;
  assign n15086 = n14646 & n14665 ;
  assign n15087 = n14648 & n15086 ;
  assign n15088 = ~n15085 & ~n15087 ;
  assign n15089 = \m2_s7_cyc_o_reg/NET0131  & n14586 ;
  assign n15090 = n2182 & n14874 ;
  assign n15091 = n14591 & n15090 ;
  assign n15092 = ~n15089 & ~n15091 ;
  assign n15093 = \m2_s13_cyc_o_reg/NET0131  & n14586 ;
  assign n15094 = n2183 & n14595 ;
  assign n15095 = n14591 & n15094 ;
  assign n15096 = ~n15093 & ~n15095 ;
  assign n15097 = \m2_s14_cyc_o_reg/NET0131  & n14586 ;
  assign n15098 = n2183 & n14850 ;
  assign n15099 = n14591 & n15098 ;
  assign n15100 = ~n15097 & ~n15099 ;
  assign n15101 = \m1_s12_cyc_o_reg/NET0131  & n14578 ;
  assign n15102 = n2156 & n14581 ;
  assign n15103 = n14583 & n15102 ;
  assign n15104 = ~n15101 & ~n15103 ;
  assign n15105 = \m1_s11_cyc_o_reg/NET0131  & n14578 ;
  assign n15106 = n2155 & n14795 ;
  assign n15107 = n14583 & n15106 ;
  assign n15108 = ~n15105 & ~n15107 ;
  assign n15109 = \m0_s9_cyc_o_reg/NET0131  & n14565 ;
  assign n15110 = n14574 & n14790 ;
  assign n15111 = n14570 & n15110 ;
  assign n15112 = ~n15109 & ~n15111 ;
  assign n15113 = \m0_s4_cyc_o_reg/NET0131  & n14565 ;
  assign n15114 = n14567 & n14761 ;
  assign n15115 = n14570 & n15114 ;
  assign n15116 = ~n15113 & ~n15115 ;
  assign n15117 = \m0_s13_cyc_o_reg/NET0131  & n14565 ;
  assign n15118 = n2162 & n14790 ;
  assign n15119 = n14570 & n15118 ;
  assign n15120 = ~n15117 & ~n15119 ;
  assign n15121 = \m0_s12_cyc_o_reg/NET0131  & n14565 ;
  assign n15122 = n14761 & n14790 ;
  assign n15123 = n14570 & n15122 ;
  assign n15124 = ~n15121 & ~n15123 ;
  assign n15125 = ~\s15_ack_i_pad  & ~n2258 ;
  assign n15126 = n1925 & n2163 ;
  assign n15127 = n1931 & n15126 ;
  assign n15128 = ~n13416 & n15127 ;
  assign n15129 = ~n15125 & n15128 ;
  assign n15130 = \s14_ack_i_pad  & n14762 ;
  assign n15131 = n14331 & n15130 ;
  assign n15132 = n14324 & n15131 ;
  assign n15133 = \s3_ack_i_pad  & n14774 ;
  assign n15134 = n14451 & n15133 ;
  assign n15135 = n14476 & n15134 ;
  assign n15136 = ~n15132 & ~n15135 ;
  assign n15137 = \s1_ack_i_pad  & n14575 ;
  assign n15138 = n14271 & n15137 ;
  assign n15139 = n14296 & n15138 ;
  assign n15140 = \s4_ack_i_pad  & n15114 ;
  assign n15141 = n13467 & n15140 ;
  assign n15142 = n13475 & n15141 ;
  assign n15143 = ~n15139 & ~n15142 ;
  assign n15144 = n15136 & n15143 ;
  assign n15145 = \s10_ack_i_pad  & n14749 ;
  assign n15146 = n13928 & n15145 ;
  assign n15147 = n13945 & n15146 ;
  assign n15148 = \s2_ack_i_pad  & n14770 ;
  assign n15149 = n14391 & n15148 ;
  assign n15150 = n14399 & n15149 ;
  assign n15151 = ~n15147 & ~n15150 ;
  assign n15152 = \s13_ack_i_pad  & n15118 ;
  assign n15153 = n14211 & n15152 ;
  assign n15154 = n14219 & n15153 ;
  assign n15155 = \s0_ack_i_pad  & n14569 ;
  assign n15156 = n14069 & n15155 ;
  assign n15157 = n14094 & n15156 ;
  assign n15158 = ~n15154 & ~n15157 ;
  assign n15159 = n15151 & n15158 ;
  assign n15160 = n15144 & n15159 ;
  assign n15161 = \s6_ack_i_pad  & n14782 ;
  assign n15162 = n13627 & n15161 ;
  assign n15163 = n13620 & n15162 ;
  assign n15164 = \s11_ack_i_pad  & n14753 ;
  assign n15165 = n14009 & n15164 ;
  assign n15166 = n14017 & n15165 ;
  assign n15167 = \s9_ack_i_pad  & n15110 ;
  assign n15168 = n13847 & n15167 ;
  assign n15169 = n13855 & n15168 ;
  assign n15170 = ~n15166 & ~n15169 ;
  assign n15171 = ~n15163 & n15170 ;
  assign n15172 = \s7_ack_i_pad  & n14786 ;
  assign n15173 = n13697 & n15172 ;
  assign n15174 = n13705 & n15173 ;
  assign n15175 = \s12_ack_i_pad  & n15122 ;
  assign n15176 = n14140 & n15175 ;
  assign n15177 = n14165 & n15176 ;
  assign n15178 = ~n15174 & ~n15177 ;
  assign n15179 = \s5_ack_i_pad  & n14778 ;
  assign n15180 = n13547 & n15179 ;
  assign n15181 = n13572 & n15180 ;
  assign n15182 = \s8_ack_i_pad  & n14791 ;
  assign n15183 = n13767 & n15182 ;
  assign n15184 = n13760 & n15183 ;
  assign n15185 = ~n15181 & ~n15184 ;
  assign n15186 = n15178 & n15185 ;
  assign n15187 = n15171 & n15186 ;
  assign n15188 = n15160 & n15187 ;
  assign n15189 = ~n15129 & n15188 ;
  assign n15190 = \rf_rf_dout_reg[0]/P0001  & ~n2106 ;
  assign n15191 = n2153 & n15190 ;
  assign n15192 = n2257 & n15191 ;
  assign n15193 = n2163 & n15192 ;
  assign n15194 = \s15_data_i[0]_pad  & n2163 ;
  assign n15195 = ~n2258 & n15194 ;
  assign n15196 = ~n15193 & ~n15195 ;
  assign n15197 = \s8_data_i[0]_pad  & n14791 ;
  assign n15198 = \s1_data_i[0]_pad  & n14575 ;
  assign n15199 = ~n15197 & ~n15198 ;
  assign n15200 = \s4_data_i[0]_pad  & n15114 ;
  assign n15201 = \s6_data_i[0]_pad  & n14782 ;
  assign n15202 = ~n15200 & ~n15201 ;
  assign n15203 = n15199 & n15202 ;
  assign n15204 = \s5_data_i[0]_pad  & n14778 ;
  assign n15205 = \s9_data_i[0]_pad  & n15110 ;
  assign n15206 = ~n15204 & ~n15205 ;
  assign n15207 = \s10_data_i[0]_pad  & n14749 ;
  assign n15208 = \s7_data_i[0]_pad  & n14786 ;
  assign n15209 = ~n15207 & ~n15208 ;
  assign n15210 = n15206 & n15209 ;
  assign n15211 = n15203 & n15210 ;
  assign n15212 = \s11_data_i[0]_pad  & n14753 ;
  assign n15213 = \s14_data_i[0]_pad  & n14762 ;
  assign n15214 = \s3_data_i[0]_pad  & n14774 ;
  assign n15215 = ~n15213 & ~n15214 ;
  assign n15216 = ~n15212 & n15215 ;
  assign n15217 = \s2_data_i[0]_pad  & n14770 ;
  assign n15218 = \s12_data_i[0]_pad  & n15122 ;
  assign n15219 = ~n15217 & ~n15218 ;
  assign n15220 = \s13_data_i[0]_pad  & n15118 ;
  assign n15221 = \s0_data_i[0]_pad  & n14569 ;
  assign n15222 = ~n15220 & ~n15221 ;
  assign n15223 = n15219 & n15222 ;
  assign n15224 = n15216 & n15223 ;
  assign n15225 = n15211 & n15224 ;
  assign n15226 = n15196 & n15225 ;
  assign n15227 = \rf_rf_dout_reg[10]/P0001  & ~n2106 ;
  assign n15228 = n2153 & n15227 ;
  assign n15229 = n2257 & n15228 ;
  assign n15230 = n2163 & n15229 ;
  assign n15231 = \s15_data_i[10]_pad  & n2163 ;
  assign n15232 = ~n2258 & n15231 ;
  assign n15233 = ~n15230 & ~n15232 ;
  assign n15234 = \s8_data_i[10]_pad  & n14791 ;
  assign n15235 = \s1_data_i[10]_pad  & n14575 ;
  assign n15236 = ~n15234 & ~n15235 ;
  assign n15237 = \s4_data_i[10]_pad  & n15114 ;
  assign n15238 = \s6_data_i[10]_pad  & n14782 ;
  assign n15239 = ~n15237 & ~n15238 ;
  assign n15240 = n15236 & n15239 ;
  assign n15241 = \s5_data_i[10]_pad  & n14778 ;
  assign n15242 = \s9_data_i[10]_pad  & n15110 ;
  assign n15243 = ~n15241 & ~n15242 ;
  assign n15244 = \s10_data_i[10]_pad  & n14749 ;
  assign n15245 = \s7_data_i[10]_pad  & n14786 ;
  assign n15246 = ~n15244 & ~n15245 ;
  assign n15247 = n15243 & n15246 ;
  assign n15248 = n15240 & n15247 ;
  assign n15249 = \s11_data_i[10]_pad  & n14753 ;
  assign n15250 = \s14_data_i[10]_pad  & n14762 ;
  assign n15251 = \s3_data_i[10]_pad  & n14774 ;
  assign n15252 = ~n15250 & ~n15251 ;
  assign n15253 = ~n15249 & n15252 ;
  assign n15254 = \s2_data_i[10]_pad  & n14770 ;
  assign n15255 = \s12_data_i[10]_pad  & n15122 ;
  assign n15256 = ~n15254 & ~n15255 ;
  assign n15257 = \s13_data_i[10]_pad  & n15118 ;
  assign n15258 = \s0_data_i[10]_pad  & n14569 ;
  assign n15259 = ~n15257 & ~n15258 ;
  assign n15260 = n15256 & n15259 ;
  assign n15261 = n15253 & n15260 ;
  assign n15262 = n15248 & n15261 ;
  assign n15263 = n15233 & n15262 ;
  assign n15264 = \rf_rf_dout_reg[11]/P0001  & ~n2106 ;
  assign n15265 = n2153 & n15264 ;
  assign n15266 = n2257 & n15265 ;
  assign n15267 = n2163 & n15266 ;
  assign n15268 = \s15_data_i[11]_pad  & n2163 ;
  assign n15269 = ~n2258 & n15268 ;
  assign n15270 = ~n15267 & ~n15269 ;
  assign n15271 = \s8_data_i[11]_pad  & n14791 ;
  assign n15272 = \s1_data_i[11]_pad  & n14575 ;
  assign n15273 = ~n15271 & ~n15272 ;
  assign n15274 = \s4_data_i[11]_pad  & n15114 ;
  assign n15275 = \s6_data_i[11]_pad  & n14782 ;
  assign n15276 = ~n15274 & ~n15275 ;
  assign n15277 = n15273 & n15276 ;
  assign n15278 = \s5_data_i[11]_pad  & n14778 ;
  assign n15279 = \s9_data_i[11]_pad  & n15110 ;
  assign n15280 = ~n15278 & ~n15279 ;
  assign n15281 = \s10_data_i[11]_pad  & n14749 ;
  assign n15282 = \s7_data_i[11]_pad  & n14786 ;
  assign n15283 = ~n15281 & ~n15282 ;
  assign n15284 = n15280 & n15283 ;
  assign n15285 = n15277 & n15284 ;
  assign n15286 = \s11_data_i[11]_pad  & n14753 ;
  assign n15287 = \s14_data_i[11]_pad  & n14762 ;
  assign n15288 = \s3_data_i[11]_pad  & n14774 ;
  assign n15289 = ~n15287 & ~n15288 ;
  assign n15290 = ~n15286 & n15289 ;
  assign n15291 = \s2_data_i[11]_pad  & n14770 ;
  assign n15292 = \s12_data_i[11]_pad  & n15122 ;
  assign n15293 = ~n15291 & ~n15292 ;
  assign n15294 = \s13_data_i[11]_pad  & n15118 ;
  assign n15295 = \s0_data_i[11]_pad  & n14569 ;
  assign n15296 = ~n15294 & ~n15295 ;
  assign n15297 = n15293 & n15296 ;
  assign n15298 = n15290 & n15297 ;
  assign n15299 = n15285 & n15298 ;
  assign n15300 = n15270 & n15299 ;
  assign n15301 = \rf_rf_dout_reg[12]/P0001  & ~n2106 ;
  assign n15302 = n2153 & n15301 ;
  assign n15303 = n2257 & n15302 ;
  assign n15304 = n2163 & n15303 ;
  assign n15305 = \s15_data_i[12]_pad  & n2163 ;
  assign n15306 = ~n2258 & n15305 ;
  assign n15307 = ~n15304 & ~n15306 ;
  assign n15308 = \s8_data_i[12]_pad  & n14791 ;
  assign n15309 = \s1_data_i[12]_pad  & n14575 ;
  assign n15310 = ~n15308 & ~n15309 ;
  assign n15311 = \s4_data_i[12]_pad  & n15114 ;
  assign n15312 = \s6_data_i[12]_pad  & n14782 ;
  assign n15313 = ~n15311 & ~n15312 ;
  assign n15314 = n15310 & n15313 ;
  assign n15315 = \s5_data_i[12]_pad  & n14778 ;
  assign n15316 = \s9_data_i[12]_pad  & n15110 ;
  assign n15317 = ~n15315 & ~n15316 ;
  assign n15318 = \s10_data_i[12]_pad  & n14749 ;
  assign n15319 = \s7_data_i[12]_pad  & n14786 ;
  assign n15320 = ~n15318 & ~n15319 ;
  assign n15321 = n15317 & n15320 ;
  assign n15322 = n15314 & n15321 ;
  assign n15323 = \s11_data_i[12]_pad  & n14753 ;
  assign n15324 = \s14_data_i[12]_pad  & n14762 ;
  assign n15325 = \s3_data_i[12]_pad  & n14774 ;
  assign n15326 = ~n15324 & ~n15325 ;
  assign n15327 = ~n15323 & n15326 ;
  assign n15328 = \s2_data_i[12]_pad  & n14770 ;
  assign n15329 = \s12_data_i[12]_pad  & n15122 ;
  assign n15330 = ~n15328 & ~n15329 ;
  assign n15331 = \s13_data_i[12]_pad  & n15118 ;
  assign n15332 = \s0_data_i[12]_pad  & n14569 ;
  assign n15333 = ~n15331 & ~n15332 ;
  assign n15334 = n15330 & n15333 ;
  assign n15335 = n15327 & n15334 ;
  assign n15336 = n15322 & n15335 ;
  assign n15337 = n15307 & n15336 ;
  assign n15338 = \rf_rf_dout_reg[13]/P0001  & ~n2106 ;
  assign n15339 = n2153 & n15338 ;
  assign n15340 = n2257 & n15339 ;
  assign n15341 = n2163 & n15340 ;
  assign n15342 = \s15_data_i[13]_pad  & n2163 ;
  assign n15343 = ~n2258 & n15342 ;
  assign n15344 = ~n15341 & ~n15343 ;
  assign n15345 = \s8_data_i[13]_pad  & n14791 ;
  assign n15346 = \s1_data_i[13]_pad  & n14575 ;
  assign n15347 = ~n15345 & ~n15346 ;
  assign n15348 = \s4_data_i[13]_pad  & n15114 ;
  assign n15349 = \s6_data_i[13]_pad  & n14782 ;
  assign n15350 = ~n15348 & ~n15349 ;
  assign n15351 = n15347 & n15350 ;
  assign n15352 = \s5_data_i[13]_pad  & n14778 ;
  assign n15353 = \s9_data_i[13]_pad  & n15110 ;
  assign n15354 = ~n15352 & ~n15353 ;
  assign n15355 = \s10_data_i[13]_pad  & n14749 ;
  assign n15356 = \s7_data_i[13]_pad  & n14786 ;
  assign n15357 = ~n15355 & ~n15356 ;
  assign n15358 = n15354 & n15357 ;
  assign n15359 = n15351 & n15358 ;
  assign n15360 = \s11_data_i[13]_pad  & n14753 ;
  assign n15361 = \s14_data_i[13]_pad  & n14762 ;
  assign n15362 = \s3_data_i[13]_pad  & n14774 ;
  assign n15363 = ~n15361 & ~n15362 ;
  assign n15364 = ~n15360 & n15363 ;
  assign n15365 = \s2_data_i[13]_pad  & n14770 ;
  assign n15366 = \s12_data_i[13]_pad  & n15122 ;
  assign n15367 = ~n15365 & ~n15366 ;
  assign n15368 = \s13_data_i[13]_pad  & n15118 ;
  assign n15369 = \s0_data_i[13]_pad  & n14569 ;
  assign n15370 = ~n15368 & ~n15369 ;
  assign n15371 = n15367 & n15370 ;
  assign n15372 = n15364 & n15371 ;
  assign n15373 = n15359 & n15372 ;
  assign n15374 = n15344 & n15373 ;
  assign n15375 = \rf_rf_dout_reg[14]/P0001  & ~n2106 ;
  assign n15376 = n2153 & n15375 ;
  assign n15377 = n2257 & n15376 ;
  assign n15378 = n2163 & n15377 ;
  assign n15379 = \s15_data_i[14]_pad  & n2163 ;
  assign n15380 = ~n2258 & n15379 ;
  assign n15381 = ~n15378 & ~n15380 ;
  assign n15382 = \s8_data_i[14]_pad  & n14791 ;
  assign n15383 = \s1_data_i[14]_pad  & n14575 ;
  assign n15384 = ~n15382 & ~n15383 ;
  assign n15385 = \s4_data_i[14]_pad  & n15114 ;
  assign n15386 = \s6_data_i[14]_pad  & n14782 ;
  assign n15387 = ~n15385 & ~n15386 ;
  assign n15388 = n15384 & n15387 ;
  assign n15389 = \s5_data_i[14]_pad  & n14778 ;
  assign n15390 = \s9_data_i[14]_pad  & n15110 ;
  assign n15391 = ~n15389 & ~n15390 ;
  assign n15392 = \s10_data_i[14]_pad  & n14749 ;
  assign n15393 = \s7_data_i[14]_pad  & n14786 ;
  assign n15394 = ~n15392 & ~n15393 ;
  assign n15395 = n15391 & n15394 ;
  assign n15396 = n15388 & n15395 ;
  assign n15397 = \s11_data_i[14]_pad  & n14753 ;
  assign n15398 = \s14_data_i[14]_pad  & n14762 ;
  assign n15399 = \s3_data_i[14]_pad  & n14774 ;
  assign n15400 = ~n15398 & ~n15399 ;
  assign n15401 = ~n15397 & n15400 ;
  assign n15402 = \s2_data_i[14]_pad  & n14770 ;
  assign n15403 = \s12_data_i[14]_pad  & n15122 ;
  assign n15404 = ~n15402 & ~n15403 ;
  assign n15405 = \s13_data_i[14]_pad  & n15118 ;
  assign n15406 = \s0_data_i[14]_pad  & n14569 ;
  assign n15407 = ~n15405 & ~n15406 ;
  assign n15408 = n15404 & n15407 ;
  assign n15409 = n15401 & n15408 ;
  assign n15410 = n15396 & n15409 ;
  assign n15411 = n15381 & n15410 ;
  assign n15412 = \rf_rf_dout_reg[15]/P0001  & ~n2106 ;
  assign n15413 = n2153 & n15412 ;
  assign n15414 = n2257 & n15413 ;
  assign n15415 = n2163 & n15414 ;
  assign n15416 = \s15_data_i[15]_pad  & n2163 ;
  assign n15417 = ~n2258 & n15416 ;
  assign n15418 = ~n15415 & ~n15417 ;
  assign n15419 = \s8_data_i[15]_pad  & n14791 ;
  assign n15420 = \s1_data_i[15]_pad  & n14575 ;
  assign n15421 = ~n15419 & ~n15420 ;
  assign n15422 = \s4_data_i[15]_pad  & n15114 ;
  assign n15423 = \s6_data_i[15]_pad  & n14782 ;
  assign n15424 = ~n15422 & ~n15423 ;
  assign n15425 = n15421 & n15424 ;
  assign n15426 = \s5_data_i[15]_pad  & n14778 ;
  assign n15427 = \s9_data_i[15]_pad  & n15110 ;
  assign n15428 = ~n15426 & ~n15427 ;
  assign n15429 = \s10_data_i[15]_pad  & n14749 ;
  assign n15430 = \s7_data_i[15]_pad  & n14786 ;
  assign n15431 = ~n15429 & ~n15430 ;
  assign n15432 = n15428 & n15431 ;
  assign n15433 = n15425 & n15432 ;
  assign n15434 = \s11_data_i[15]_pad  & n14753 ;
  assign n15435 = \s14_data_i[15]_pad  & n14762 ;
  assign n15436 = \s3_data_i[15]_pad  & n14774 ;
  assign n15437 = ~n15435 & ~n15436 ;
  assign n15438 = ~n15434 & n15437 ;
  assign n15439 = \s2_data_i[15]_pad  & n14770 ;
  assign n15440 = \s12_data_i[15]_pad  & n15122 ;
  assign n15441 = ~n15439 & ~n15440 ;
  assign n15442 = \s13_data_i[15]_pad  & n15118 ;
  assign n15443 = \s0_data_i[15]_pad  & n14569 ;
  assign n15444 = ~n15442 & ~n15443 ;
  assign n15445 = n15441 & n15444 ;
  assign n15446 = n15438 & n15445 ;
  assign n15447 = n15433 & n15446 ;
  assign n15448 = n15418 & n15447 ;
  assign n15449 = \s15_data_i[16]_pad  & n2163 ;
  assign n15450 = ~n2258 & n15449 ;
  assign n15451 = \s8_data_i[16]_pad  & n14791 ;
  assign n15452 = \s1_data_i[16]_pad  & n14575 ;
  assign n15453 = ~n15451 & ~n15452 ;
  assign n15454 = \s4_data_i[16]_pad  & n15114 ;
  assign n15455 = \s6_data_i[16]_pad  & n14782 ;
  assign n15456 = ~n15454 & ~n15455 ;
  assign n15457 = n15453 & n15456 ;
  assign n15458 = \s5_data_i[16]_pad  & n14778 ;
  assign n15459 = \s9_data_i[16]_pad  & n15110 ;
  assign n15460 = ~n15458 & ~n15459 ;
  assign n15461 = \s10_data_i[16]_pad  & n14749 ;
  assign n15462 = \s7_data_i[16]_pad  & n14786 ;
  assign n15463 = ~n15461 & ~n15462 ;
  assign n15464 = n15460 & n15463 ;
  assign n15465 = n15457 & n15464 ;
  assign n15466 = \s11_data_i[16]_pad  & n14753 ;
  assign n15467 = \s14_data_i[16]_pad  & n14762 ;
  assign n15468 = \s3_data_i[16]_pad  & n14774 ;
  assign n15469 = ~n15467 & ~n15468 ;
  assign n15470 = ~n15466 & n15469 ;
  assign n15471 = \s2_data_i[16]_pad  & n14770 ;
  assign n15472 = \s12_data_i[16]_pad  & n15122 ;
  assign n15473 = ~n15471 & ~n15472 ;
  assign n15474 = \s13_data_i[16]_pad  & n15118 ;
  assign n15475 = \s0_data_i[16]_pad  & n14569 ;
  assign n15476 = ~n15474 & ~n15475 ;
  assign n15477 = n15473 & n15476 ;
  assign n15478 = n15470 & n15477 ;
  assign n15479 = n15465 & n15478 ;
  assign n15480 = ~n15450 & n15479 ;
  assign n15481 = \s15_data_i[17]_pad  & n2163 ;
  assign n15482 = ~n2258 & n15481 ;
  assign n15483 = \s8_data_i[17]_pad  & n14791 ;
  assign n15484 = \s1_data_i[17]_pad  & n14575 ;
  assign n15485 = ~n15483 & ~n15484 ;
  assign n15486 = \s4_data_i[17]_pad  & n15114 ;
  assign n15487 = \s6_data_i[17]_pad  & n14782 ;
  assign n15488 = ~n15486 & ~n15487 ;
  assign n15489 = n15485 & n15488 ;
  assign n15490 = \s5_data_i[17]_pad  & n14778 ;
  assign n15491 = \s9_data_i[17]_pad  & n15110 ;
  assign n15492 = ~n15490 & ~n15491 ;
  assign n15493 = \s10_data_i[17]_pad  & n14749 ;
  assign n15494 = \s7_data_i[17]_pad  & n14786 ;
  assign n15495 = ~n15493 & ~n15494 ;
  assign n15496 = n15492 & n15495 ;
  assign n15497 = n15489 & n15496 ;
  assign n15498 = \s11_data_i[17]_pad  & n14753 ;
  assign n15499 = \s14_data_i[17]_pad  & n14762 ;
  assign n15500 = \s3_data_i[17]_pad  & n14774 ;
  assign n15501 = ~n15499 & ~n15500 ;
  assign n15502 = ~n15498 & n15501 ;
  assign n15503 = \s2_data_i[17]_pad  & n14770 ;
  assign n15504 = \s12_data_i[17]_pad  & n15122 ;
  assign n15505 = ~n15503 & ~n15504 ;
  assign n15506 = \s13_data_i[17]_pad  & n15118 ;
  assign n15507 = \s0_data_i[17]_pad  & n14569 ;
  assign n15508 = ~n15506 & ~n15507 ;
  assign n15509 = n15505 & n15508 ;
  assign n15510 = n15502 & n15509 ;
  assign n15511 = n15497 & n15510 ;
  assign n15512 = ~n15482 & n15511 ;
  assign n15513 = \s15_data_i[18]_pad  & n2163 ;
  assign n15514 = ~n2258 & n15513 ;
  assign n15515 = \s8_data_i[18]_pad  & n14791 ;
  assign n15516 = \s1_data_i[18]_pad  & n14575 ;
  assign n15517 = ~n15515 & ~n15516 ;
  assign n15518 = \s4_data_i[18]_pad  & n15114 ;
  assign n15519 = \s6_data_i[18]_pad  & n14782 ;
  assign n15520 = ~n15518 & ~n15519 ;
  assign n15521 = n15517 & n15520 ;
  assign n15522 = \s5_data_i[18]_pad  & n14778 ;
  assign n15523 = \s9_data_i[18]_pad  & n15110 ;
  assign n15524 = ~n15522 & ~n15523 ;
  assign n15525 = \s10_data_i[18]_pad  & n14749 ;
  assign n15526 = \s7_data_i[18]_pad  & n14786 ;
  assign n15527 = ~n15525 & ~n15526 ;
  assign n15528 = n15524 & n15527 ;
  assign n15529 = n15521 & n15528 ;
  assign n15530 = \s11_data_i[18]_pad  & n14753 ;
  assign n15531 = \s14_data_i[18]_pad  & n14762 ;
  assign n15532 = \s3_data_i[18]_pad  & n14774 ;
  assign n15533 = ~n15531 & ~n15532 ;
  assign n15534 = ~n15530 & n15533 ;
  assign n15535 = \s2_data_i[18]_pad  & n14770 ;
  assign n15536 = \s12_data_i[18]_pad  & n15122 ;
  assign n15537 = ~n15535 & ~n15536 ;
  assign n15538 = \s13_data_i[18]_pad  & n15118 ;
  assign n15539 = \s0_data_i[18]_pad  & n14569 ;
  assign n15540 = ~n15538 & ~n15539 ;
  assign n15541 = n15537 & n15540 ;
  assign n15542 = n15534 & n15541 ;
  assign n15543 = n15529 & n15542 ;
  assign n15544 = ~n15514 & n15543 ;
  assign n15545 = \s15_data_i[19]_pad  & n2163 ;
  assign n15546 = ~n2258 & n15545 ;
  assign n15547 = \s8_data_i[19]_pad  & n14791 ;
  assign n15548 = \s1_data_i[19]_pad  & n14575 ;
  assign n15549 = ~n15547 & ~n15548 ;
  assign n15550 = \s4_data_i[19]_pad  & n15114 ;
  assign n15551 = \s6_data_i[19]_pad  & n14782 ;
  assign n15552 = ~n15550 & ~n15551 ;
  assign n15553 = n15549 & n15552 ;
  assign n15554 = \s5_data_i[19]_pad  & n14778 ;
  assign n15555 = \s9_data_i[19]_pad  & n15110 ;
  assign n15556 = ~n15554 & ~n15555 ;
  assign n15557 = \s10_data_i[19]_pad  & n14749 ;
  assign n15558 = \s7_data_i[19]_pad  & n14786 ;
  assign n15559 = ~n15557 & ~n15558 ;
  assign n15560 = n15556 & n15559 ;
  assign n15561 = n15553 & n15560 ;
  assign n15562 = \s11_data_i[19]_pad  & n14753 ;
  assign n15563 = \s14_data_i[19]_pad  & n14762 ;
  assign n15564 = \s3_data_i[19]_pad  & n14774 ;
  assign n15565 = ~n15563 & ~n15564 ;
  assign n15566 = ~n15562 & n15565 ;
  assign n15567 = \s2_data_i[19]_pad  & n14770 ;
  assign n15568 = \s12_data_i[19]_pad  & n15122 ;
  assign n15569 = ~n15567 & ~n15568 ;
  assign n15570 = \s13_data_i[19]_pad  & n15118 ;
  assign n15571 = \s0_data_i[19]_pad  & n14569 ;
  assign n15572 = ~n15570 & ~n15571 ;
  assign n15573 = n15569 & n15572 ;
  assign n15574 = n15566 & n15573 ;
  assign n15575 = n15561 & n15574 ;
  assign n15576 = ~n15546 & n15575 ;
  assign n15577 = \rf_rf_dout_reg[1]/P0001  & ~n2106 ;
  assign n15578 = n2153 & n15577 ;
  assign n15579 = n2257 & n15578 ;
  assign n15580 = n2163 & n15579 ;
  assign n15581 = \s15_data_i[1]_pad  & n2163 ;
  assign n15582 = ~n2258 & n15581 ;
  assign n15583 = ~n15580 & ~n15582 ;
  assign n15584 = \s8_data_i[1]_pad  & n14791 ;
  assign n15585 = \s1_data_i[1]_pad  & n14575 ;
  assign n15586 = ~n15584 & ~n15585 ;
  assign n15587 = \s4_data_i[1]_pad  & n15114 ;
  assign n15588 = \s6_data_i[1]_pad  & n14782 ;
  assign n15589 = ~n15587 & ~n15588 ;
  assign n15590 = n15586 & n15589 ;
  assign n15591 = \s5_data_i[1]_pad  & n14778 ;
  assign n15592 = \s9_data_i[1]_pad  & n15110 ;
  assign n15593 = ~n15591 & ~n15592 ;
  assign n15594 = \s10_data_i[1]_pad  & n14749 ;
  assign n15595 = \s7_data_i[1]_pad  & n14786 ;
  assign n15596 = ~n15594 & ~n15595 ;
  assign n15597 = n15593 & n15596 ;
  assign n15598 = n15590 & n15597 ;
  assign n15599 = \s11_data_i[1]_pad  & n14753 ;
  assign n15600 = \s14_data_i[1]_pad  & n14762 ;
  assign n15601 = \s3_data_i[1]_pad  & n14774 ;
  assign n15602 = ~n15600 & ~n15601 ;
  assign n15603 = ~n15599 & n15602 ;
  assign n15604 = \s2_data_i[1]_pad  & n14770 ;
  assign n15605 = \s12_data_i[1]_pad  & n15122 ;
  assign n15606 = ~n15604 & ~n15605 ;
  assign n15607 = \s13_data_i[1]_pad  & n15118 ;
  assign n15608 = \s0_data_i[1]_pad  & n14569 ;
  assign n15609 = ~n15607 & ~n15608 ;
  assign n15610 = n15606 & n15609 ;
  assign n15611 = n15603 & n15610 ;
  assign n15612 = n15598 & n15611 ;
  assign n15613 = n15583 & n15612 ;
  assign n15614 = \s15_data_i[20]_pad  & n2163 ;
  assign n15615 = ~n2258 & n15614 ;
  assign n15616 = \s8_data_i[20]_pad  & n14791 ;
  assign n15617 = \s1_data_i[20]_pad  & n14575 ;
  assign n15618 = ~n15616 & ~n15617 ;
  assign n15619 = \s4_data_i[20]_pad  & n15114 ;
  assign n15620 = \s6_data_i[20]_pad  & n14782 ;
  assign n15621 = ~n15619 & ~n15620 ;
  assign n15622 = n15618 & n15621 ;
  assign n15623 = \s5_data_i[20]_pad  & n14778 ;
  assign n15624 = \s9_data_i[20]_pad  & n15110 ;
  assign n15625 = ~n15623 & ~n15624 ;
  assign n15626 = \s10_data_i[20]_pad  & n14749 ;
  assign n15627 = \s7_data_i[20]_pad  & n14786 ;
  assign n15628 = ~n15626 & ~n15627 ;
  assign n15629 = n15625 & n15628 ;
  assign n15630 = n15622 & n15629 ;
  assign n15631 = \s11_data_i[20]_pad  & n14753 ;
  assign n15632 = \s14_data_i[20]_pad  & n14762 ;
  assign n15633 = \s3_data_i[20]_pad  & n14774 ;
  assign n15634 = ~n15632 & ~n15633 ;
  assign n15635 = ~n15631 & n15634 ;
  assign n15636 = \s2_data_i[20]_pad  & n14770 ;
  assign n15637 = \s12_data_i[20]_pad  & n15122 ;
  assign n15638 = ~n15636 & ~n15637 ;
  assign n15639 = \s13_data_i[20]_pad  & n15118 ;
  assign n15640 = \s0_data_i[20]_pad  & n14569 ;
  assign n15641 = ~n15639 & ~n15640 ;
  assign n15642 = n15638 & n15641 ;
  assign n15643 = n15635 & n15642 ;
  assign n15644 = n15630 & n15643 ;
  assign n15645 = ~n15615 & n15644 ;
  assign n15646 = \s15_data_i[21]_pad  & n2163 ;
  assign n15647 = ~n2258 & n15646 ;
  assign n15648 = \s8_data_i[21]_pad  & n14791 ;
  assign n15649 = \s1_data_i[21]_pad  & n14575 ;
  assign n15650 = ~n15648 & ~n15649 ;
  assign n15651 = \s4_data_i[21]_pad  & n15114 ;
  assign n15652 = \s6_data_i[21]_pad  & n14782 ;
  assign n15653 = ~n15651 & ~n15652 ;
  assign n15654 = n15650 & n15653 ;
  assign n15655 = \s5_data_i[21]_pad  & n14778 ;
  assign n15656 = \s9_data_i[21]_pad  & n15110 ;
  assign n15657 = ~n15655 & ~n15656 ;
  assign n15658 = \s10_data_i[21]_pad  & n14749 ;
  assign n15659 = \s7_data_i[21]_pad  & n14786 ;
  assign n15660 = ~n15658 & ~n15659 ;
  assign n15661 = n15657 & n15660 ;
  assign n15662 = n15654 & n15661 ;
  assign n15663 = \s11_data_i[21]_pad  & n14753 ;
  assign n15664 = \s14_data_i[21]_pad  & n14762 ;
  assign n15665 = \s3_data_i[21]_pad  & n14774 ;
  assign n15666 = ~n15664 & ~n15665 ;
  assign n15667 = ~n15663 & n15666 ;
  assign n15668 = \s2_data_i[21]_pad  & n14770 ;
  assign n15669 = \s12_data_i[21]_pad  & n15122 ;
  assign n15670 = ~n15668 & ~n15669 ;
  assign n15671 = \s13_data_i[21]_pad  & n15118 ;
  assign n15672 = \s0_data_i[21]_pad  & n14569 ;
  assign n15673 = ~n15671 & ~n15672 ;
  assign n15674 = n15670 & n15673 ;
  assign n15675 = n15667 & n15674 ;
  assign n15676 = n15662 & n15675 ;
  assign n15677 = ~n15647 & n15676 ;
  assign n15678 = \s15_data_i[22]_pad  & n2163 ;
  assign n15679 = ~n2258 & n15678 ;
  assign n15680 = \s8_data_i[22]_pad  & n14791 ;
  assign n15681 = \s1_data_i[22]_pad  & n14575 ;
  assign n15682 = ~n15680 & ~n15681 ;
  assign n15683 = \s4_data_i[22]_pad  & n15114 ;
  assign n15684 = \s6_data_i[22]_pad  & n14782 ;
  assign n15685 = ~n15683 & ~n15684 ;
  assign n15686 = n15682 & n15685 ;
  assign n15687 = \s5_data_i[22]_pad  & n14778 ;
  assign n15688 = \s9_data_i[22]_pad  & n15110 ;
  assign n15689 = ~n15687 & ~n15688 ;
  assign n15690 = \s10_data_i[22]_pad  & n14749 ;
  assign n15691 = \s7_data_i[22]_pad  & n14786 ;
  assign n15692 = ~n15690 & ~n15691 ;
  assign n15693 = n15689 & n15692 ;
  assign n15694 = n15686 & n15693 ;
  assign n15695 = \s11_data_i[22]_pad  & n14753 ;
  assign n15696 = \s14_data_i[22]_pad  & n14762 ;
  assign n15697 = \s3_data_i[22]_pad  & n14774 ;
  assign n15698 = ~n15696 & ~n15697 ;
  assign n15699 = ~n15695 & n15698 ;
  assign n15700 = \s2_data_i[22]_pad  & n14770 ;
  assign n15701 = \s12_data_i[22]_pad  & n15122 ;
  assign n15702 = ~n15700 & ~n15701 ;
  assign n15703 = \s13_data_i[22]_pad  & n15118 ;
  assign n15704 = \s0_data_i[22]_pad  & n14569 ;
  assign n15705 = ~n15703 & ~n15704 ;
  assign n15706 = n15702 & n15705 ;
  assign n15707 = n15699 & n15706 ;
  assign n15708 = n15694 & n15707 ;
  assign n15709 = ~n15679 & n15708 ;
  assign n15710 = \s15_data_i[23]_pad  & n2163 ;
  assign n15711 = ~n2258 & n15710 ;
  assign n15712 = \s8_data_i[23]_pad  & n14791 ;
  assign n15713 = \s1_data_i[23]_pad  & n14575 ;
  assign n15714 = ~n15712 & ~n15713 ;
  assign n15715 = \s4_data_i[23]_pad  & n15114 ;
  assign n15716 = \s6_data_i[23]_pad  & n14782 ;
  assign n15717 = ~n15715 & ~n15716 ;
  assign n15718 = n15714 & n15717 ;
  assign n15719 = \s5_data_i[23]_pad  & n14778 ;
  assign n15720 = \s9_data_i[23]_pad  & n15110 ;
  assign n15721 = ~n15719 & ~n15720 ;
  assign n15722 = \s10_data_i[23]_pad  & n14749 ;
  assign n15723 = \s7_data_i[23]_pad  & n14786 ;
  assign n15724 = ~n15722 & ~n15723 ;
  assign n15725 = n15721 & n15724 ;
  assign n15726 = n15718 & n15725 ;
  assign n15727 = \s11_data_i[23]_pad  & n14753 ;
  assign n15728 = \s14_data_i[23]_pad  & n14762 ;
  assign n15729 = \s3_data_i[23]_pad  & n14774 ;
  assign n15730 = ~n15728 & ~n15729 ;
  assign n15731 = ~n15727 & n15730 ;
  assign n15732 = \s2_data_i[23]_pad  & n14770 ;
  assign n15733 = \s12_data_i[23]_pad  & n15122 ;
  assign n15734 = ~n15732 & ~n15733 ;
  assign n15735 = \s13_data_i[23]_pad  & n15118 ;
  assign n15736 = \s0_data_i[23]_pad  & n14569 ;
  assign n15737 = ~n15735 & ~n15736 ;
  assign n15738 = n15734 & n15737 ;
  assign n15739 = n15731 & n15738 ;
  assign n15740 = n15726 & n15739 ;
  assign n15741 = ~n15711 & n15740 ;
  assign n15742 = \s15_data_i[24]_pad  & n2163 ;
  assign n15743 = ~n2258 & n15742 ;
  assign n15744 = \s8_data_i[24]_pad  & n14791 ;
  assign n15745 = \s1_data_i[24]_pad  & n14575 ;
  assign n15746 = ~n15744 & ~n15745 ;
  assign n15747 = \s4_data_i[24]_pad  & n15114 ;
  assign n15748 = \s6_data_i[24]_pad  & n14782 ;
  assign n15749 = ~n15747 & ~n15748 ;
  assign n15750 = n15746 & n15749 ;
  assign n15751 = \s5_data_i[24]_pad  & n14778 ;
  assign n15752 = \s9_data_i[24]_pad  & n15110 ;
  assign n15753 = ~n15751 & ~n15752 ;
  assign n15754 = \s10_data_i[24]_pad  & n14749 ;
  assign n15755 = \s7_data_i[24]_pad  & n14786 ;
  assign n15756 = ~n15754 & ~n15755 ;
  assign n15757 = n15753 & n15756 ;
  assign n15758 = n15750 & n15757 ;
  assign n15759 = \s11_data_i[24]_pad  & n14753 ;
  assign n15760 = \s14_data_i[24]_pad  & n14762 ;
  assign n15761 = \s3_data_i[24]_pad  & n14774 ;
  assign n15762 = ~n15760 & ~n15761 ;
  assign n15763 = ~n15759 & n15762 ;
  assign n15764 = \s2_data_i[24]_pad  & n14770 ;
  assign n15765 = \s12_data_i[24]_pad  & n15122 ;
  assign n15766 = ~n15764 & ~n15765 ;
  assign n15767 = \s13_data_i[24]_pad  & n15118 ;
  assign n15768 = \s0_data_i[24]_pad  & n14569 ;
  assign n15769 = ~n15767 & ~n15768 ;
  assign n15770 = n15766 & n15769 ;
  assign n15771 = n15763 & n15770 ;
  assign n15772 = n15758 & n15771 ;
  assign n15773 = ~n15743 & n15772 ;
  assign n15774 = \s15_data_i[25]_pad  & n2163 ;
  assign n15775 = ~n2258 & n15774 ;
  assign n15776 = \s8_data_i[25]_pad  & n14791 ;
  assign n15777 = \s1_data_i[25]_pad  & n14575 ;
  assign n15778 = ~n15776 & ~n15777 ;
  assign n15779 = \s4_data_i[25]_pad  & n15114 ;
  assign n15780 = \s6_data_i[25]_pad  & n14782 ;
  assign n15781 = ~n15779 & ~n15780 ;
  assign n15782 = n15778 & n15781 ;
  assign n15783 = \s5_data_i[25]_pad  & n14778 ;
  assign n15784 = \s9_data_i[25]_pad  & n15110 ;
  assign n15785 = ~n15783 & ~n15784 ;
  assign n15786 = \s10_data_i[25]_pad  & n14749 ;
  assign n15787 = \s7_data_i[25]_pad  & n14786 ;
  assign n15788 = ~n15786 & ~n15787 ;
  assign n15789 = n15785 & n15788 ;
  assign n15790 = n15782 & n15789 ;
  assign n15791 = \s11_data_i[25]_pad  & n14753 ;
  assign n15792 = \s14_data_i[25]_pad  & n14762 ;
  assign n15793 = \s3_data_i[25]_pad  & n14774 ;
  assign n15794 = ~n15792 & ~n15793 ;
  assign n15795 = ~n15791 & n15794 ;
  assign n15796 = \s2_data_i[25]_pad  & n14770 ;
  assign n15797 = \s12_data_i[25]_pad  & n15122 ;
  assign n15798 = ~n15796 & ~n15797 ;
  assign n15799 = \s13_data_i[25]_pad  & n15118 ;
  assign n15800 = \s0_data_i[25]_pad  & n14569 ;
  assign n15801 = ~n15799 & ~n15800 ;
  assign n15802 = n15798 & n15801 ;
  assign n15803 = n15795 & n15802 ;
  assign n15804 = n15790 & n15803 ;
  assign n15805 = ~n15775 & n15804 ;
  assign n15806 = \s15_data_i[26]_pad  & n2163 ;
  assign n15807 = ~n2258 & n15806 ;
  assign n15808 = \s8_data_i[26]_pad  & n14791 ;
  assign n15809 = \s1_data_i[26]_pad  & n14575 ;
  assign n15810 = ~n15808 & ~n15809 ;
  assign n15811 = \s4_data_i[26]_pad  & n15114 ;
  assign n15812 = \s6_data_i[26]_pad  & n14782 ;
  assign n15813 = ~n15811 & ~n15812 ;
  assign n15814 = n15810 & n15813 ;
  assign n15815 = \s5_data_i[26]_pad  & n14778 ;
  assign n15816 = \s9_data_i[26]_pad  & n15110 ;
  assign n15817 = ~n15815 & ~n15816 ;
  assign n15818 = \s10_data_i[26]_pad  & n14749 ;
  assign n15819 = \s7_data_i[26]_pad  & n14786 ;
  assign n15820 = ~n15818 & ~n15819 ;
  assign n15821 = n15817 & n15820 ;
  assign n15822 = n15814 & n15821 ;
  assign n15823 = \s11_data_i[26]_pad  & n14753 ;
  assign n15824 = \s14_data_i[26]_pad  & n14762 ;
  assign n15825 = \s3_data_i[26]_pad  & n14774 ;
  assign n15826 = ~n15824 & ~n15825 ;
  assign n15827 = ~n15823 & n15826 ;
  assign n15828 = \s2_data_i[26]_pad  & n14770 ;
  assign n15829 = \s12_data_i[26]_pad  & n15122 ;
  assign n15830 = ~n15828 & ~n15829 ;
  assign n15831 = \s13_data_i[26]_pad  & n15118 ;
  assign n15832 = \s0_data_i[26]_pad  & n14569 ;
  assign n15833 = ~n15831 & ~n15832 ;
  assign n15834 = n15830 & n15833 ;
  assign n15835 = n15827 & n15834 ;
  assign n15836 = n15822 & n15835 ;
  assign n15837 = ~n15807 & n15836 ;
  assign n15838 = \s15_data_i[27]_pad  & n2163 ;
  assign n15839 = ~n2258 & n15838 ;
  assign n15840 = \s8_data_i[27]_pad  & n14791 ;
  assign n15841 = \s1_data_i[27]_pad  & n14575 ;
  assign n15842 = ~n15840 & ~n15841 ;
  assign n15843 = \s4_data_i[27]_pad  & n15114 ;
  assign n15844 = \s6_data_i[27]_pad  & n14782 ;
  assign n15845 = ~n15843 & ~n15844 ;
  assign n15846 = n15842 & n15845 ;
  assign n15847 = \s5_data_i[27]_pad  & n14778 ;
  assign n15848 = \s9_data_i[27]_pad  & n15110 ;
  assign n15849 = ~n15847 & ~n15848 ;
  assign n15850 = \s10_data_i[27]_pad  & n14749 ;
  assign n15851 = \s7_data_i[27]_pad  & n14786 ;
  assign n15852 = ~n15850 & ~n15851 ;
  assign n15853 = n15849 & n15852 ;
  assign n15854 = n15846 & n15853 ;
  assign n15855 = \s11_data_i[27]_pad  & n14753 ;
  assign n15856 = \s14_data_i[27]_pad  & n14762 ;
  assign n15857 = \s3_data_i[27]_pad  & n14774 ;
  assign n15858 = ~n15856 & ~n15857 ;
  assign n15859 = ~n15855 & n15858 ;
  assign n15860 = \s2_data_i[27]_pad  & n14770 ;
  assign n15861 = \s12_data_i[27]_pad  & n15122 ;
  assign n15862 = ~n15860 & ~n15861 ;
  assign n15863 = \s13_data_i[27]_pad  & n15118 ;
  assign n15864 = \s0_data_i[27]_pad  & n14569 ;
  assign n15865 = ~n15863 & ~n15864 ;
  assign n15866 = n15862 & n15865 ;
  assign n15867 = n15859 & n15866 ;
  assign n15868 = n15854 & n15867 ;
  assign n15869 = ~n15839 & n15868 ;
  assign n15870 = \s15_data_i[28]_pad  & n2163 ;
  assign n15871 = ~n2258 & n15870 ;
  assign n15872 = \s8_data_i[28]_pad  & n14791 ;
  assign n15873 = \s1_data_i[28]_pad  & n14575 ;
  assign n15874 = ~n15872 & ~n15873 ;
  assign n15875 = \s4_data_i[28]_pad  & n15114 ;
  assign n15876 = \s6_data_i[28]_pad  & n14782 ;
  assign n15877 = ~n15875 & ~n15876 ;
  assign n15878 = n15874 & n15877 ;
  assign n15879 = \s5_data_i[28]_pad  & n14778 ;
  assign n15880 = \s9_data_i[28]_pad  & n15110 ;
  assign n15881 = ~n15879 & ~n15880 ;
  assign n15882 = \s10_data_i[28]_pad  & n14749 ;
  assign n15883 = \s7_data_i[28]_pad  & n14786 ;
  assign n15884 = ~n15882 & ~n15883 ;
  assign n15885 = n15881 & n15884 ;
  assign n15886 = n15878 & n15885 ;
  assign n15887 = \s11_data_i[28]_pad  & n14753 ;
  assign n15888 = \s14_data_i[28]_pad  & n14762 ;
  assign n15889 = \s3_data_i[28]_pad  & n14774 ;
  assign n15890 = ~n15888 & ~n15889 ;
  assign n15891 = ~n15887 & n15890 ;
  assign n15892 = \s2_data_i[28]_pad  & n14770 ;
  assign n15893 = \s12_data_i[28]_pad  & n15122 ;
  assign n15894 = ~n15892 & ~n15893 ;
  assign n15895 = \s13_data_i[28]_pad  & n15118 ;
  assign n15896 = \s0_data_i[28]_pad  & n14569 ;
  assign n15897 = ~n15895 & ~n15896 ;
  assign n15898 = n15894 & n15897 ;
  assign n15899 = n15891 & n15898 ;
  assign n15900 = n15886 & n15899 ;
  assign n15901 = ~n15871 & n15900 ;
  assign n15902 = \s15_data_i[29]_pad  & n2163 ;
  assign n15903 = ~n2258 & n15902 ;
  assign n15904 = \s8_data_i[29]_pad  & n14791 ;
  assign n15905 = \s1_data_i[29]_pad  & n14575 ;
  assign n15906 = ~n15904 & ~n15905 ;
  assign n15907 = \s4_data_i[29]_pad  & n15114 ;
  assign n15908 = \s6_data_i[29]_pad  & n14782 ;
  assign n15909 = ~n15907 & ~n15908 ;
  assign n15910 = n15906 & n15909 ;
  assign n15911 = \s5_data_i[29]_pad  & n14778 ;
  assign n15912 = \s9_data_i[29]_pad  & n15110 ;
  assign n15913 = ~n15911 & ~n15912 ;
  assign n15914 = \s10_data_i[29]_pad  & n14749 ;
  assign n15915 = \s7_data_i[29]_pad  & n14786 ;
  assign n15916 = ~n15914 & ~n15915 ;
  assign n15917 = n15913 & n15916 ;
  assign n15918 = n15910 & n15917 ;
  assign n15919 = \s11_data_i[29]_pad  & n14753 ;
  assign n15920 = \s14_data_i[29]_pad  & n14762 ;
  assign n15921 = \s3_data_i[29]_pad  & n14774 ;
  assign n15922 = ~n15920 & ~n15921 ;
  assign n15923 = ~n15919 & n15922 ;
  assign n15924 = \s2_data_i[29]_pad  & n14770 ;
  assign n15925 = \s12_data_i[29]_pad  & n15122 ;
  assign n15926 = ~n15924 & ~n15925 ;
  assign n15927 = \s13_data_i[29]_pad  & n15118 ;
  assign n15928 = \s0_data_i[29]_pad  & n14569 ;
  assign n15929 = ~n15927 & ~n15928 ;
  assign n15930 = n15926 & n15929 ;
  assign n15931 = n15923 & n15930 ;
  assign n15932 = n15918 & n15931 ;
  assign n15933 = ~n15903 & n15932 ;
  assign n15934 = \rf_rf_dout_reg[2]/P0001  & ~n2106 ;
  assign n15935 = n2153 & n15934 ;
  assign n15936 = n2257 & n15935 ;
  assign n15937 = n2163 & n15936 ;
  assign n15938 = \s15_data_i[2]_pad  & n2163 ;
  assign n15939 = ~n2258 & n15938 ;
  assign n15940 = ~n15937 & ~n15939 ;
  assign n15941 = \s8_data_i[2]_pad  & n14791 ;
  assign n15942 = \s1_data_i[2]_pad  & n14575 ;
  assign n15943 = ~n15941 & ~n15942 ;
  assign n15944 = \s4_data_i[2]_pad  & n15114 ;
  assign n15945 = \s6_data_i[2]_pad  & n14782 ;
  assign n15946 = ~n15944 & ~n15945 ;
  assign n15947 = n15943 & n15946 ;
  assign n15948 = \s5_data_i[2]_pad  & n14778 ;
  assign n15949 = \s9_data_i[2]_pad  & n15110 ;
  assign n15950 = ~n15948 & ~n15949 ;
  assign n15951 = \s10_data_i[2]_pad  & n14749 ;
  assign n15952 = \s7_data_i[2]_pad  & n14786 ;
  assign n15953 = ~n15951 & ~n15952 ;
  assign n15954 = n15950 & n15953 ;
  assign n15955 = n15947 & n15954 ;
  assign n15956 = \s11_data_i[2]_pad  & n14753 ;
  assign n15957 = \s14_data_i[2]_pad  & n14762 ;
  assign n15958 = \s3_data_i[2]_pad  & n14774 ;
  assign n15959 = ~n15957 & ~n15958 ;
  assign n15960 = ~n15956 & n15959 ;
  assign n15961 = \s2_data_i[2]_pad  & n14770 ;
  assign n15962 = \s12_data_i[2]_pad  & n15122 ;
  assign n15963 = ~n15961 & ~n15962 ;
  assign n15964 = \s13_data_i[2]_pad  & n15118 ;
  assign n15965 = \s0_data_i[2]_pad  & n14569 ;
  assign n15966 = ~n15964 & ~n15965 ;
  assign n15967 = n15963 & n15966 ;
  assign n15968 = n15960 & n15967 ;
  assign n15969 = n15955 & n15968 ;
  assign n15970 = n15940 & n15969 ;
  assign n15971 = \s15_data_i[30]_pad  & n2163 ;
  assign n15972 = ~n2258 & n15971 ;
  assign n15973 = \s8_data_i[30]_pad  & n14791 ;
  assign n15974 = \s1_data_i[30]_pad  & n14575 ;
  assign n15975 = ~n15973 & ~n15974 ;
  assign n15976 = \s4_data_i[30]_pad  & n15114 ;
  assign n15977 = \s6_data_i[30]_pad  & n14782 ;
  assign n15978 = ~n15976 & ~n15977 ;
  assign n15979 = n15975 & n15978 ;
  assign n15980 = \s5_data_i[30]_pad  & n14778 ;
  assign n15981 = \s9_data_i[30]_pad  & n15110 ;
  assign n15982 = ~n15980 & ~n15981 ;
  assign n15983 = \s10_data_i[30]_pad  & n14749 ;
  assign n15984 = \s7_data_i[30]_pad  & n14786 ;
  assign n15985 = ~n15983 & ~n15984 ;
  assign n15986 = n15982 & n15985 ;
  assign n15987 = n15979 & n15986 ;
  assign n15988 = \s11_data_i[30]_pad  & n14753 ;
  assign n15989 = \s14_data_i[30]_pad  & n14762 ;
  assign n15990 = \s3_data_i[30]_pad  & n14774 ;
  assign n15991 = ~n15989 & ~n15990 ;
  assign n15992 = ~n15988 & n15991 ;
  assign n15993 = \s2_data_i[30]_pad  & n14770 ;
  assign n15994 = \s12_data_i[30]_pad  & n15122 ;
  assign n15995 = ~n15993 & ~n15994 ;
  assign n15996 = \s13_data_i[30]_pad  & n15118 ;
  assign n15997 = \s0_data_i[30]_pad  & n14569 ;
  assign n15998 = ~n15996 & ~n15997 ;
  assign n15999 = n15995 & n15998 ;
  assign n16000 = n15992 & n15999 ;
  assign n16001 = n15987 & n16000 ;
  assign n16002 = ~n15972 & n16001 ;
  assign n16003 = \s15_data_i[31]_pad  & n2163 ;
  assign n16004 = ~n2258 & n16003 ;
  assign n16005 = \s8_data_i[31]_pad  & n14791 ;
  assign n16006 = \s1_data_i[31]_pad  & n14575 ;
  assign n16007 = ~n16005 & ~n16006 ;
  assign n16008 = \s4_data_i[31]_pad  & n15114 ;
  assign n16009 = \s6_data_i[31]_pad  & n14782 ;
  assign n16010 = ~n16008 & ~n16009 ;
  assign n16011 = n16007 & n16010 ;
  assign n16012 = \s5_data_i[31]_pad  & n14778 ;
  assign n16013 = \s9_data_i[31]_pad  & n15110 ;
  assign n16014 = ~n16012 & ~n16013 ;
  assign n16015 = \s10_data_i[31]_pad  & n14749 ;
  assign n16016 = \s7_data_i[31]_pad  & n14786 ;
  assign n16017 = ~n16015 & ~n16016 ;
  assign n16018 = n16014 & n16017 ;
  assign n16019 = n16011 & n16018 ;
  assign n16020 = \s11_data_i[31]_pad  & n14753 ;
  assign n16021 = \s14_data_i[31]_pad  & n14762 ;
  assign n16022 = \s3_data_i[31]_pad  & n14774 ;
  assign n16023 = ~n16021 & ~n16022 ;
  assign n16024 = ~n16020 & n16023 ;
  assign n16025 = \s2_data_i[31]_pad  & n14770 ;
  assign n16026 = \s12_data_i[31]_pad  & n15122 ;
  assign n16027 = ~n16025 & ~n16026 ;
  assign n16028 = \s13_data_i[31]_pad  & n15118 ;
  assign n16029 = \s0_data_i[31]_pad  & n14569 ;
  assign n16030 = ~n16028 & ~n16029 ;
  assign n16031 = n16027 & n16030 ;
  assign n16032 = n16024 & n16031 ;
  assign n16033 = n16019 & n16032 ;
  assign n16034 = ~n16004 & n16033 ;
  assign n16035 = \rf_rf_dout_reg[3]/P0001  & ~n2106 ;
  assign n16036 = n2153 & n16035 ;
  assign n16037 = n2257 & n16036 ;
  assign n16038 = n2163 & n16037 ;
  assign n16039 = \s15_data_i[3]_pad  & n2163 ;
  assign n16040 = ~n2258 & n16039 ;
  assign n16041 = ~n16038 & ~n16040 ;
  assign n16042 = \s8_data_i[3]_pad  & n14791 ;
  assign n16043 = \s1_data_i[3]_pad  & n14575 ;
  assign n16044 = ~n16042 & ~n16043 ;
  assign n16045 = \s4_data_i[3]_pad  & n15114 ;
  assign n16046 = \s6_data_i[3]_pad  & n14782 ;
  assign n16047 = ~n16045 & ~n16046 ;
  assign n16048 = n16044 & n16047 ;
  assign n16049 = \s5_data_i[3]_pad  & n14778 ;
  assign n16050 = \s9_data_i[3]_pad  & n15110 ;
  assign n16051 = ~n16049 & ~n16050 ;
  assign n16052 = \s10_data_i[3]_pad  & n14749 ;
  assign n16053 = \s7_data_i[3]_pad  & n14786 ;
  assign n16054 = ~n16052 & ~n16053 ;
  assign n16055 = n16051 & n16054 ;
  assign n16056 = n16048 & n16055 ;
  assign n16057 = \s11_data_i[3]_pad  & n14753 ;
  assign n16058 = \s14_data_i[3]_pad  & n14762 ;
  assign n16059 = \s3_data_i[3]_pad  & n14774 ;
  assign n16060 = ~n16058 & ~n16059 ;
  assign n16061 = ~n16057 & n16060 ;
  assign n16062 = \s2_data_i[3]_pad  & n14770 ;
  assign n16063 = \s12_data_i[3]_pad  & n15122 ;
  assign n16064 = ~n16062 & ~n16063 ;
  assign n16065 = \s13_data_i[3]_pad  & n15118 ;
  assign n16066 = \s0_data_i[3]_pad  & n14569 ;
  assign n16067 = ~n16065 & ~n16066 ;
  assign n16068 = n16064 & n16067 ;
  assign n16069 = n16061 & n16068 ;
  assign n16070 = n16056 & n16069 ;
  assign n16071 = n16041 & n16070 ;
  assign n16072 = \rf_rf_dout_reg[4]/P0001  & ~n2106 ;
  assign n16073 = n2153 & n16072 ;
  assign n16074 = n2257 & n16073 ;
  assign n16075 = n2163 & n16074 ;
  assign n16076 = \s15_data_i[4]_pad  & n2163 ;
  assign n16077 = ~n2258 & n16076 ;
  assign n16078 = ~n16075 & ~n16077 ;
  assign n16079 = \s8_data_i[4]_pad  & n14791 ;
  assign n16080 = \s1_data_i[4]_pad  & n14575 ;
  assign n16081 = ~n16079 & ~n16080 ;
  assign n16082 = \s4_data_i[4]_pad  & n15114 ;
  assign n16083 = \s6_data_i[4]_pad  & n14782 ;
  assign n16084 = ~n16082 & ~n16083 ;
  assign n16085 = n16081 & n16084 ;
  assign n16086 = \s5_data_i[4]_pad  & n14778 ;
  assign n16087 = \s9_data_i[4]_pad  & n15110 ;
  assign n16088 = ~n16086 & ~n16087 ;
  assign n16089 = \s10_data_i[4]_pad  & n14749 ;
  assign n16090 = \s7_data_i[4]_pad  & n14786 ;
  assign n16091 = ~n16089 & ~n16090 ;
  assign n16092 = n16088 & n16091 ;
  assign n16093 = n16085 & n16092 ;
  assign n16094 = \s11_data_i[4]_pad  & n14753 ;
  assign n16095 = \s14_data_i[4]_pad  & n14762 ;
  assign n16096 = \s3_data_i[4]_pad  & n14774 ;
  assign n16097 = ~n16095 & ~n16096 ;
  assign n16098 = ~n16094 & n16097 ;
  assign n16099 = \s2_data_i[4]_pad  & n14770 ;
  assign n16100 = \s12_data_i[4]_pad  & n15122 ;
  assign n16101 = ~n16099 & ~n16100 ;
  assign n16102 = \s13_data_i[4]_pad  & n15118 ;
  assign n16103 = \s0_data_i[4]_pad  & n14569 ;
  assign n16104 = ~n16102 & ~n16103 ;
  assign n16105 = n16101 & n16104 ;
  assign n16106 = n16098 & n16105 ;
  assign n16107 = n16093 & n16106 ;
  assign n16108 = n16078 & n16107 ;
  assign n16109 = \rf_rf_dout_reg[5]/P0001  & ~n2106 ;
  assign n16110 = n2153 & n16109 ;
  assign n16111 = n2257 & n16110 ;
  assign n16112 = n2163 & n16111 ;
  assign n16113 = \s15_data_i[5]_pad  & n2163 ;
  assign n16114 = ~n2258 & n16113 ;
  assign n16115 = ~n16112 & ~n16114 ;
  assign n16116 = \s8_data_i[5]_pad  & n14791 ;
  assign n16117 = \s1_data_i[5]_pad  & n14575 ;
  assign n16118 = ~n16116 & ~n16117 ;
  assign n16119 = \s4_data_i[5]_pad  & n15114 ;
  assign n16120 = \s6_data_i[5]_pad  & n14782 ;
  assign n16121 = ~n16119 & ~n16120 ;
  assign n16122 = n16118 & n16121 ;
  assign n16123 = \s5_data_i[5]_pad  & n14778 ;
  assign n16124 = \s9_data_i[5]_pad  & n15110 ;
  assign n16125 = ~n16123 & ~n16124 ;
  assign n16126 = \s10_data_i[5]_pad  & n14749 ;
  assign n16127 = \s7_data_i[5]_pad  & n14786 ;
  assign n16128 = ~n16126 & ~n16127 ;
  assign n16129 = n16125 & n16128 ;
  assign n16130 = n16122 & n16129 ;
  assign n16131 = \s11_data_i[5]_pad  & n14753 ;
  assign n16132 = \s14_data_i[5]_pad  & n14762 ;
  assign n16133 = \s3_data_i[5]_pad  & n14774 ;
  assign n16134 = ~n16132 & ~n16133 ;
  assign n16135 = ~n16131 & n16134 ;
  assign n16136 = \s2_data_i[5]_pad  & n14770 ;
  assign n16137 = \s12_data_i[5]_pad  & n15122 ;
  assign n16138 = ~n16136 & ~n16137 ;
  assign n16139 = \s13_data_i[5]_pad  & n15118 ;
  assign n16140 = \s0_data_i[5]_pad  & n14569 ;
  assign n16141 = ~n16139 & ~n16140 ;
  assign n16142 = n16138 & n16141 ;
  assign n16143 = n16135 & n16142 ;
  assign n16144 = n16130 & n16143 ;
  assign n16145 = n16115 & n16144 ;
  assign n16146 = \rf_rf_dout_reg[6]/P0001  & ~n2106 ;
  assign n16147 = n2153 & n16146 ;
  assign n16148 = n2257 & n16147 ;
  assign n16149 = n2163 & n16148 ;
  assign n16150 = \s15_data_i[6]_pad  & n2163 ;
  assign n16151 = ~n2258 & n16150 ;
  assign n16152 = ~n16149 & ~n16151 ;
  assign n16153 = \s8_data_i[6]_pad  & n14791 ;
  assign n16154 = \s1_data_i[6]_pad  & n14575 ;
  assign n16155 = ~n16153 & ~n16154 ;
  assign n16156 = \s4_data_i[6]_pad  & n15114 ;
  assign n16157 = \s6_data_i[6]_pad  & n14782 ;
  assign n16158 = ~n16156 & ~n16157 ;
  assign n16159 = n16155 & n16158 ;
  assign n16160 = \s5_data_i[6]_pad  & n14778 ;
  assign n16161 = \s9_data_i[6]_pad  & n15110 ;
  assign n16162 = ~n16160 & ~n16161 ;
  assign n16163 = \s10_data_i[6]_pad  & n14749 ;
  assign n16164 = \s7_data_i[6]_pad  & n14786 ;
  assign n16165 = ~n16163 & ~n16164 ;
  assign n16166 = n16162 & n16165 ;
  assign n16167 = n16159 & n16166 ;
  assign n16168 = \s11_data_i[6]_pad  & n14753 ;
  assign n16169 = \s14_data_i[6]_pad  & n14762 ;
  assign n16170 = \s3_data_i[6]_pad  & n14774 ;
  assign n16171 = ~n16169 & ~n16170 ;
  assign n16172 = ~n16168 & n16171 ;
  assign n16173 = \s2_data_i[6]_pad  & n14770 ;
  assign n16174 = \s12_data_i[6]_pad  & n15122 ;
  assign n16175 = ~n16173 & ~n16174 ;
  assign n16176 = \s13_data_i[6]_pad  & n15118 ;
  assign n16177 = \s0_data_i[6]_pad  & n14569 ;
  assign n16178 = ~n16176 & ~n16177 ;
  assign n16179 = n16175 & n16178 ;
  assign n16180 = n16172 & n16179 ;
  assign n16181 = n16167 & n16180 ;
  assign n16182 = n16152 & n16181 ;
  assign n16183 = \rf_rf_dout_reg[7]/P0001  & ~n2106 ;
  assign n16184 = n2153 & n16183 ;
  assign n16185 = n2257 & n16184 ;
  assign n16186 = n2163 & n16185 ;
  assign n16187 = \s15_data_i[7]_pad  & n2163 ;
  assign n16188 = ~n2258 & n16187 ;
  assign n16189 = ~n16186 & ~n16188 ;
  assign n16190 = \s8_data_i[7]_pad  & n14791 ;
  assign n16191 = \s1_data_i[7]_pad  & n14575 ;
  assign n16192 = ~n16190 & ~n16191 ;
  assign n16193 = \s4_data_i[7]_pad  & n15114 ;
  assign n16194 = \s6_data_i[7]_pad  & n14782 ;
  assign n16195 = ~n16193 & ~n16194 ;
  assign n16196 = n16192 & n16195 ;
  assign n16197 = \s5_data_i[7]_pad  & n14778 ;
  assign n16198 = \s9_data_i[7]_pad  & n15110 ;
  assign n16199 = ~n16197 & ~n16198 ;
  assign n16200 = \s10_data_i[7]_pad  & n14749 ;
  assign n16201 = \s7_data_i[7]_pad  & n14786 ;
  assign n16202 = ~n16200 & ~n16201 ;
  assign n16203 = n16199 & n16202 ;
  assign n16204 = n16196 & n16203 ;
  assign n16205 = \s11_data_i[7]_pad  & n14753 ;
  assign n16206 = \s14_data_i[7]_pad  & n14762 ;
  assign n16207 = \s3_data_i[7]_pad  & n14774 ;
  assign n16208 = ~n16206 & ~n16207 ;
  assign n16209 = ~n16205 & n16208 ;
  assign n16210 = \s2_data_i[7]_pad  & n14770 ;
  assign n16211 = \s12_data_i[7]_pad  & n15122 ;
  assign n16212 = ~n16210 & ~n16211 ;
  assign n16213 = \s13_data_i[7]_pad  & n15118 ;
  assign n16214 = \s0_data_i[7]_pad  & n14569 ;
  assign n16215 = ~n16213 & ~n16214 ;
  assign n16216 = n16212 & n16215 ;
  assign n16217 = n16209 & n16216 ;
  assign n16218 = n16204 & n16217 ;
  assign n16219 = n16189 & n16218 ;
  assign n16220 = \rf_rf_dout_reg[8]/P0001  & ~n2106 ;
  assign n16221 = n2153 & n16220 ;
  assign n16222 = n2257 & n16221 ;
  assign n16223 = n2163 & n16222 ;
  assign n16224 = \s15_data_i[8]_pad  & n2163 ;
  assign n16225 = ~n2258 & n16224 ;
  assign n16226 = ~n16223 & ~n16225 ;
  assign n16227 = \s8_data_i[8]_pad  & n14791 ;
  assign n16228 = \s1_data_i[8]_pad  & n14575 ;
  assign n16229 = ~n16227 & ~n16228 ;
  assign n16230 = \s4_data_i[8]_pad  & n15114 ;
  assign n16231 = \s6_data_i[8]_pad  & n14782 ;
  assign n16232 = ~n16230 & ~n16231 ;
  assign n16233 = n16229 & n16232 ;
  assign n16234 = \s5_data_i[8]_pad  & n14778 ;
  assign n16235 = \s9_data_i[8]_pad  & n15110 ;
  assign n16236 = ~n16234 & ~n16235 ;
  assign n16237 = \s10_data_i[8]_pad  & n14749 ;
  assign n16238 = \s7_data_i[8]_pad  & n14786 ;
  assign n16239 = ~n16237 & ~n16238 ;
  assign n16240 = n16236 & n16239 ;
  assign n16241 = n16233 & n16240 ;
  assign n16242 = \s11_data_i[8]_pad  & n14753 ;
  assign n16243 = \s14_data_i[8]_pad  & n14762 ;
  assign n16244 = \s3_data_i[8]_pad  & n14774 ;
  assign n16245 = ~n16243 & ~n16244 ;
  assign n16246 = ~n16242 & n16245 ;
  assign n16247 = \s2_data_i[8]_pad  & n14770 ;
  assign n16248 = \s12_data_i[8]_pad  & n15122 ;
  assign n16249 = ~n16247 & ~n16248 ;
  assign n16250 = \s13_data_i[8]_pad  & n15118 ;
  assign n16251 = \s0_data_i[8]_pad  & n14569 ;
  assign n16252 = ~n16250 & ~n16251 ;
  assign n16253 = n16249 & n16252 ;
  assign n16254 = n16246 & n16253 ;
  assign n16255 = n16241 & n16254 ;
  assign n16256 = n16226 & n16255 ;
  assign n16257 = \rf_rf_dout_reg[9]/P0001  & ~n2106 ;
  assign n16258 = n2153 & n16257 ;
  assign n16259 = n2257 & n16258 ;
  assign n16260 = n2163 & n16259 ;
  assign n16261 = \s15_data_i[9]_pad  & n2163 ;
  assign n16262 = ~n2258 & n16261 ;
  assign n16263 = ~n16260 & ~n16262 ;
  assign n16264 = \s8_data_i[9]_pad  & n14791 ;
  assign n16265 = \s1_data_i[9]_pad  & n14575 ;
  assign n16266 = ~n16264 & ~n16265 ;
  assign n16267 = \s4_data_i[9]_pad  & n15114 ;
  assign n16268 = \s6_data_i[9]_pad  & n14782 ;
  assign n16269 = ~n16267 & ~n16268 ;
  assign n16270 = n16266 & n16269 ;
  assign n16271 = \s5_data_i[9]_pad  & n14778 ;
  assign n16272 = \s9_data_i[9]_pad  & n15110 ;
  assign n16273 = ~n16271 & ~n16272 ;
  assign n16274 = \s10_data_i[9]_pad  & n14749 ;
  assign n16275 = \s7_data_i[9]_pad  & n14786 ;
  assign n16276 = ~n16274 & ~n16275 ;
  assign n16277 = n16273 & n16276 ;
  assign n16278 = n16270 & n16277 ;
  assign n16279 = \s11_data_i[9]_pad  & n14753 ;
  assign n16280 = \s14_data_i[9]_pad  & n14762 ;
  assign n16281 = \s3_data_i[9]_pad  & n14774 ;
  assign n16282 = ~n16280 & ~n16281 ;
  assign n16283 = ~n16279 & n16282 ;
  assign n16284 = \s2_data_i[9]_pad  & n14770 ;
  assign n16285 = \s12_data_i[9]_pad  & n15122 ;
  assign n16286 = ~n16284 & ~n16285 ;
  assign n16287 = \s13_data_i[9]_pad  & n15118 ;
  assign n16288 = \s0_data_i[9]_pad  & n14569 ;
  assign n16289 = ~n16287 & ~n16288 ;
  assign n16290 = n16286 & n16289 ;
  assign n16291 = n16283 & n16290 ;
  assign n16292 = n16278 & n16291 ;
  assign n16293 = n16263 & n16292 ;
  assign n16294 = \s15_err_i_pad  & n15127 ;
  assign n16295 = ~n2258 & n16294 ;
  assign n16296 = \s0_err_i_pad  & n14569 ;
  assign n16297 = n14069 & n16296 ;
  assign n16298 = n14094 & n16297 ;
  assign n16299 = \s8_err_i_pad  & n14791 ;
  assign n16300 = n13767 & n16299 ;
  assign n16301 = n13760 & n16300 ;
  assign n16302 = ~n16298 & ~n16301 ;
  assign n16303 = \s3_err_i_pad  & n14774 ;
  assign n16304 = n14451 & n16303 ;
  assign n16305 = n14476 & n16304 ;
  assign n16306 = \s14_err_i_pad  & n14762 ;
  assign n16307 = n14331 & n16306 ;
  assign n16308 = n14324 & n16307 ;
  assign n16309 = ~n16305 & ~n16308 ;
  assign n16310 = n16302 & n16309 ;
  assign n16311 = \s7_err_i_pad  & n14786 ;
  assign n16312 = n13697 & n16311 ;
  assign n16313 = n13705 & n16312 ;
  assign n16314 = \s5_err_i_pad  & n14778 ;
  assign n16315 = n13547 & n16314 ;
  assign n16316 = n13572 & n16315 ;
  assign n16317 = ~n16313 & ~n16316 ;
  assign n16318 = \s12_err_i_pad  & n15122 ;
  assign n16319 = n14140 & n16318 ;
  assign n16320 = n14165 & n16319 ;
  assign n16321 = \s13_err_i_pad  & n15118 ;
  assign n16322 = n14211 & n16321 ;
  assign n16323 = n14219 & n16322 ;
  assign n16324 = ~n16320 & ~n16323 ;
  assign n16325 = n16317 & n16324 ;
  assign n16326 = n16310 & n16325 ;
  assign n16327 = \s4_err_i_pad  & n15114 ;
  assign n16328 = n13467 & n16327 ;
  assign n16329 = n13475 & n16328 ;
  assign n16330 = \s1_err_i_pad  & n14575 ;
  assign n16331 = n14271 & n16330 ;
  assign n16332 = n14296 & n16331 ;
  assign n16333 = \s6_err_i_pad  & n14782 ;
  assign n16334 = n13627 & n16333 ;
  assign n16335 = n13620 & n16334 ;
  assign n16336 = ~n16332 & ~n16335 ;
  assign n16337 = ~n16329 & n16336 ;
  assign n16338 = \s9_err_i_pad  & n15110 ;
  assign n16339 = n13847 & n16338 ;
  assign n16340 = n13855 & n16339 ;
  assign n16341 = \s10_err_i_pad  & n14749 ;
  assign n16342 = n13928 & n16341 ;
  assign n16343 = n13945 & n16342 ;
  assign n16344 = ~n16340 & ~n16343 ;
  assign n16345 = \s11_err_i_pad  & n14753 ;
  assign n16346 = n14009 & n16345 ;
  assign n16347 = n14017 & n16346 ;
  assign n16348 = \s2_err_i_pad  & n14770 ;
  assign n16349 = n14391 & n16348 ;
  assign n16350 = n14399 & n16349 ;
  assign n16351 = ~n16347 & ~n16350 ;
  assign n16352 = n16344 & n16351 ;
  assign n16353 = n16337 & n16352 ;
  assign n16354 = n16326 & n16353 ;
  assign n16355 = ~n16295 & n16354 ;
  assign n16356 = \s15_rty_i_pad  & n15127 ;
  assign n16357 = ~n2258 & n16356 ;
  assign n16358 = \s6_rty_i_pad  & n14782 ;
  assign n16359 = n13627 & n16358 ;
  assign n16360 = n13620 & n16359 ;
  assign n16361 = \s12_rty_i_pad  & n15122 ;
  assign n16362 = n14140 & n16361 ;
  assign n16363 = n14165 & n16362 ;
  assign n16364 = ~n16360 & ~n16363 ;
  assign n16365 = \s3_rty_i_pad  & n14774 ;
  assign n16366 = n14451 & n16365 ;
  assign n16367 = n14476 & n16366 ;
  assign n16368 = \s11_rty_i_pad  & n14753 ;
  assign n16369 = n14009 & n16368 ;
  assign n16370 = n14017 & n16369 ;
  assign n16371 = ~n16367 & ~n16370 ;
  assign n16372 = n16364 & n16371 ;
  assign n16373 = \s10_rty_i_pad  & n14749 ;
  assign n16374 = n13928 & n16373 ;
  assign n16375 = n13945 & n16374 ;
  assign n16376 = \s5_rty_i_pad  & n14778 ;
  assign n16377 = n13547 & n16376 ;
  assign n16378 = n13572 & n16377 ;
  assign n16379 = ~n16375 & ~n16378 ;
  assign n16380 = \s8_rty_i_pad  & n14791 ;
  assign n16381 = n13767 & n16380 ;
  assign n16382 = n13760 & n16381 ;
  assign n16383 = \s13_rty_i_pad  & n15118 ;
  assign n16384 = n14211 & n16383 ;
  assign n16385 = n14219 & n16384 ;
  assign n16386 = ~n16382 & ~n16385 ;
  assign n16387 = n16379 & n16386 ;
  assign n16388 = n16372 & n16387 ;
  assign n16389 = \s7_rty_i_pad  & n14786 ;
  assign n16390 = n13697 & n16389 ;
  assign n16391 = n13705 & n16390 ;
  assign n16392 = \s1_rty_i_pad  & n14575 ;
  assign n16393 = n14271 & n16392 ;
  assign n16394 = n14296 & n16393 ;
  assign n16395 = \s9_rty_i_pad  & n15110 ;
  assign n16396 = n13847 & n16395 ;
  assign n16397 = n13855 & n16396 ;
  assign n16398 = ~n16394 & ~n16397 ;
  assign n16399 = ~n16391 & n16398 ;
  assign n16400 = \s0_rty_i_pad  & n14569 ;
  assign n16401 = n14069 & n16400 ;
  assign n16402 = n14094 & n16401 ;
  assign n16403 = \s4_rty_i_pad  & n15114 ;
  assign n16404 = n13467 & n16403 ;
  assign n16405 = n13475 & n16404 ;
  assign n16406 = ~n16402 & ~n16405 ;
  assign n16407 = \s14_rty_i_pad  & n14762 ;
  assign n16408 = n14331 & n16407 ;
  assign n16409 = n14324 & n16408 ;
  assign n16410 = \s2_rty_i_pad  & n14770 ;
  assign n16411 = n14391 & n16410 ;
  assign n16412 = n14399 & n16411 ;
  assign n16413 = ~n16409 & ~n16412 ;
  assign n16414 = n16406 & n16413 ;
  assign n16415 = n16399 & n16414 ;
  assign n16416 = n16388 & n16415 ;
  assign n16417 = ~n16357 & n16416 ;
  assign n16418 = n1910 & n2157 ;
  assign n16419 = n1941 & n16418 ;
  assign n16420 = ~n13416 & n16419 ;
  assign n16421 = ~n15125 & n16420 ;
  assign n16422 = \s5_ack_i_pad  & n14829 ;
  assign n16423 = ~n13547 & n16422 ;
  assign n16424 = n13572 & n16423 ;
  assign n16425 = \s1_ack_i_pad  & n14658 ;
  assign n16426 = ~n14271 & n16425 ;
  assign n16427 = n14296 & n16426 ;
  assign n16428 = ~n16424 & ~n16427 ;
  assign n16429 = \s12_ack_i_pad  & n15102 ;
  assign n16430 = ~n14140 & n16429 ;
  assign n16431 = n14165 & n16430 ;
  assign n16432 = \s10_ack_i_pad  & n14797 ;
  assign n16433 = ~n13928 & n16432 ;
  assign n16434 = n13945 & n16433 ;
  assign n16435 = ~n16431 & ~n16434 ;
  assign n16436 = n16428 & n16435 ;
  assign n16437 = \s7_ack_i_pad  & n14837 ;
  assign n16438 = ~n13697 & n16437 ;
  assign n16439 = n13705 & n16438 ;
  assign n16440 = \s14_ack_i_pad  & n14809 ;
  assign n16441 = ~n14331 & n16440 ;
  assign n16442 = n14324 & n16441 ;
  assign n16443 = ~n16439 & ~n16442 ;
  assign n16444 = \s13_ack_i_pad  & n14805 ;
  assign n16445 = ~n14211 & n16444 ;
  assign n16446 = n14219 & n16445 ;
  assign n16447 = \s9_ack_i_pad  & n14845 ;
  assign n16448 = ~n13847 & n16447 ;
  assign n16449 = n13855 & n16448 ;
  assign n16450 = ~n16446 & ~n16449 ;
  assign n16451 = n16443 & n16450 ;
  assign n16452 = n16436 & n16451 ;
  assign n16453 = \s3_ack_i_pad  & n14820 ;
  assign n16454 = ~n14451 & n16453 ;
  assign n16455 = n14476 & n16454 ;
  assign n16456 = \s11_ack_i_pad  & n15106 ;
  assign n16457 = ~n14009 & n16456 ;
  assign n16458 = n14017 & n16457 ;
  assign n16459 = \s6_ack_i_pad  & n14833 ;
  assign n16460 = ~n13627 & n16459 ;
  assign n16461 = n13620 & n16460 ;
  assign n16462 = ~n16458 & ~n16461 ;
  assign n16463 = ~n16455 & n16462 ;
  assign n16464 = \s4_ack_i_pad  & n14825 ;
  assign n16465 = ~n13467 & n16464 ;
  assign n16466 = n13475 & n16465 ;
  assign n16467 = \s0_ack_i_pad  & n14582 ;
  assign n16468 = ~n14069 & n16467 ;
  assign n16469 = n14094 & n16468 ;
  assign n16470 = ~n16466 & ~n16469 ;
  assign n16471 = \s2_ack_i_pad  & n14816 ;
  assign n16472 = ~n14391 & n16471 ;
  assign n16473 = n14399 & n16472 ;
  assign n16474 = \s8_ack_i_pad  & n14841 ;
  assign n16475 = ~n13767 & n16474 ;
  assign n16476 = n13760 & n16475 ;
  assign n16477 = ~n16473 & ~n16476 ;
  assign n16478 = n16470 & n16477 ;
  assign n16479 = n16463 & n16478 ;
  assign n16480 = n16452 & n16479 ;
  assign n16481 = ~n16421 & n16480 ;
  assign n16482 = n2157 & n15192 ;
  assign n16483 = \s15_data_i[0]_pad  & n2157 ;
  assign n16484 = ~n2258 & n16483 ;
  assign n16485 = ~n16482 & ~n16484 ;
  assign n16486 = \s12_data_i[0]_pad  & n15102 ;
  assign n16487 = \s1_data_i[0]_pad  & n14658 ;
  assign n16488 = ~n16486 & ~n16487 ;
  assign n16489 = \s0_data_i[0]_pad  & n14582 ;
  assign n16490 = \s10_data_i[0]_pad  & n14797 ;
  assign n16491 = ~n16489 & ~n16490 ;
  assign n16492 = n16488 & n16491 ;
  assign n16493 = \s3_data_i[0]_pad  & n14820 ;
  assign n16494 = \s4_data_i[0]_pad  & n14825 ;
  assign n16495 = ~n16493 & ~n16494 ;
  assign n16496 = \s9_data_i[0]_pad  & n14845 ;
  assign n16497 = \s6_data_i[0]_pad  & n14833 ;
  assign n16498 = ~n16496 & ~n16497 ;
  assign n16499 = n16495 & n16498 ;
  assign n16500 = n16492 & n16499 ;
  assign n16501 = \s14_data_i[0]_pad  & n14809 ;
  assign n16502 = \s11_data_i[0]_pad  & n15106 ;
  assign n16503 = \s7_data_i[0]_pad  & n14837 ;
  assign n16504 = ~n16502 & ~n16503 ;
  assign n16505 = ~n16501 & n16504 ;
  assign n16506 = \s5_data_i[0]_pad  & n14829 ;
  assign n16507 = \s8_data_i[0]_pad  & n14841 ;
  assign n16508 = ~n16506 & ~n16507 ;
  assign n16509 = \s2_data_i[0]_pad  & n14816 ;
  assign n16510 = \s13_data_i[0]_pad  & n14805 ;
  assign n16511 = ~n16509 & ~n16510 ;
  assign n16512 = n16508 & n16511 ;
  assign n16513 = n16505 & n16512 ;
  assign n16514 = n16500 & n16513 ;
  assign n16515 = n16485 & n16514 ;
  assign n16516 = n2157 & n15229 ;
  assign n16517 = \s15_data_i[10]_pad  & n2157 ;
  assign n16518 = ~n2258 & n16517 ;
  assign n16519 = ~n16516 & ~n16518 ;
  assign n16520 = \s12_data_i[10]_pad  & n15102 ;
  assign n16521 = \s1_data_i[10]_pad  & n14658 ;
  assign n16522 = ~n16520 & ~n16521 ;
  assign n16523 = \s0_data_i[10]_pad  & n14582 ;
  assign n16524 = \s10_data_i[10]_pad  & n14797 ;
  assign n16525 = ~n16523 & ~n16524 ;
  assign n16526 = n16522 & n16525 ;
  assign n16527 = \s3_data_i[10]_pad  & n14820 ;
  assign n16528 = \s4_data_i[10]_pad  & n14825 ;
  assign n16529 = ~n16527 & ~n16528 ;
  assign n16530 = \s9_data_i[10]_pad  & n14845 ;
  assign n16531 = \s6_data_i[10]_pad  & n14833 ;
  assign n16532 = ~n16530 & ~n16531 ;
  assign n16533 = n16529 & n16532 ;
  assign n16534 = n16526 & n16533 ;
  assign n16535 = \s14_data_i[10]_pad  & n14809 ;
  assign n16536 = \s11_data_i[10]_pad  & n15106 ;
  assign n16537 = \s7_data_i[10]_pad  & n14837 ;
  assign n16538 = ~n16536 & ~n16537 ;
  assign n16539 = ~n16535 & n16538 ;
  assign n16540 = \s5_data_i[10]_pad  & n14829 ;
  assign n16541 = \s8_data_i[10]_pad  & n14841 ;
  assign n16542 = ~n16540 & ~n16541 ;
  assign n16543 = \s2_data_i[10]_pad  & n14816 ;
  assign n16544 = \s13_data_i[10]_pad  & n14805 ;
  assign n16545 = ~n16543 & ~n16544 ;
  assign n16546 = n16542 & n16545 ;
  assign n16547 = n16539 & n16546 ;
  assign n16548 = n16534 & n16547 ;
  assign n16549 = n16519 & n16548 ;
  assign n16550 = n2157 & n15266 ;
  assign n16551 = \s15_data_i[11]_pad  & n2157 ;
  assign n16552 = ~n2258 & n16551 ;
  assign n16553 = ~n16550 & ~n16552 ;
  assign n16554 = \s14_data_i[11]_pad  & n14809 ;
  assign n16555 = \s1_data_i[11]_pad  & n14658 ;
  assign n16556 = ~n16554 & ~n16555 ;
  assign n16557 = \s10_data_i[11]_pad  & n14797 ;
  assign n16558 = \s7_data_i[11]_pad  & n14837 ;
  assign n16559 = ~n16557 & ~n16558 ;
  assign n16560 = n16556 & n16559 ;
  assign n16561 = \s5_data_i[11]_pad  & n14829 ;
  assign n16562 = \s2_data_i[11]_pad  & n14816 ;
  assign n16563 = ~n16561 & ~n16562 ;
  assign n16564 = \s6_data_i[11]_pad  & n14833 ;
  assign n16565 = \s0_data_i[11]_pad  & n14582 ;
  assign n16566 = ~n16564 & ~n16565 ;
  assign n16567 = n16563 & n16566 ;
  assign n16568 = n16560 & n16567 ;
  assign n16569 = \s11_data_i[11]_pad  & n15106 ;
  assign n16570 = \s8_data_i[11]_pad  & n14841 ;
  assign n16571 = \s4_data_i[11]_pad  & n14825 ;
  assign n16572 = ~n16570 & ~n16571 ;
  assign n16573 = ~n16569 & n16572 ;
  assign n16574 = \s3_data_i[11]_pad  & n14820 ;
  assign n16575 = \s12_data_i[11]_pad  & n15102 ;
  assign n16576 = ~n16574 & ~n16575 ;
  assign n16577 = \s13_data_i[11]_pad  & n14805 ;
  assign n16578 = \s9_data_i[11]_pad  & n14845 ;
  assign n16579 = ~n16577 & ~n16578 ;
  assign n16580 = n16576 & n16579 ;
  assign n16581 = n16573 & n16580 ;
  assign n16582 = n16568 & n16581 ;
  assign n16583 = n16553 & n16582 ;
  assign n16584 = n2157 & n15303 ;
  assign n16585 = \s15_data_i[12]_pad  & n2157 ;
  assign n16586 = ~n2258 & n16585 ;
  assign n16587 = ~n16584 & ~n16586 ;
  assign n16588 = \s12_data_i[12]_pad  & n15102 ;
  assign n16589 = \s1_data_i[12]_pad  & n14658 ;
  assign n16590 = ~n16588 & ~n16589 ;
  assign n16591 = \s0_data_i[12]_pad  & n14582 ;
  assign n16592 = \s10_data_i[12]_pad  & n14797 ;
  assign n16593 = ~n16591 & ~n16592 ;
  assign n16594 = n16590 & n16593 ;
  assign n16595 = \s3_data_i[12]_pad  & n14820 ;
  assign n16596 = \s4_data_i[12]_pad  & n14825 ;
  assign n16597 = ~n16595 & ~n16596 ;
  assign n16598 = \s9_data_i[12]_pad  & n14845 ;
  assign n16599 = \s6_data_i[12]_pad  & n14833 ;
  assign n16600 = ~n16598 & ~n16599 ;
  assign n16601 = n16597 & n16600 ;
  assign n16602 = n16594 & n16601 ;
  assign n16603 = \s14_data_i[12]_pad  & n14809 ;
  assign n16604 = \s11_data_i[12]_pad  & n15106 ;
  assign n16605 = \s7_data_i[12]_pad  & n14837 ;
  assign n16606 = ~n16604 & ~n16605 ;
  assign n16607 = ~n16603 & n16606 ;
  assign n16608 = \s5_data_i[12]_pad  & n14829 ;
  assign n16609 = \s8_data_i[12]_pad  & n14841 ;
  assign n16610 = ~n16608 & ~n16609 ;
  assign n16611 = \s2_data_i[12]_pad  & n14816 ;
  assign n16612 = \s13_data_i[12]_pad  & n14805 ;
  assign n16613 = ~n16611 & ~n16612 ;
  assign n16614 = n16610 & n16613 ;
  assign n16615 = n16607 & n16614 ;
  assign n16616 = n16602 & n16615 ;
  assign n16617 = n16587 & n16616 ;
  assign n16618 = n2157 & n15340 ;
  assign n16619 = \s15_data_i[13]_pad  & n2157 ;
  assign n16620 = ~n2258 & n16619 ;
  assign n16621 = ~n16618 & ~n16620 ;
  assign n16622 = \s12_data_i[13]_pad  & n15102 ;
  assign n16623 = \s1_data_i[13]_pad  & n14658 ;
  assign n16624 = ~n16622 & ~n16623 ;
  assign n16625 = \s0_data_i[13]_pad  & n14582 ;
  assign n16626 = \s10_data_i[13]_pad  & n14797 ;
  assign n16627 = ~n16625 & ~n16626 ;
  assign n16628 = n16624 & n16627 ;
  assign n16629 = \s3_data_i[13]_pad  & n14820 ;
  assign n16630 = \s4_data_i[13]_pad  & n14825 ;
  assign n16631 = ~n16629 & ~n16630 ;
  assign n16632 = \s9_data_i[13]_pad  & n14845 ;
  assign n16633 = \s6_data_i[13]_pad  & n14833 ;
  assign n16634 = ~n16632 & ~n16633 ;
  assign n16635 = n16631 & n16634 ;
  assign n16636 = n16628 & n16635 ;
  assign n16637 = \s14_data_i[13]_pad  & n14809 ;
  assign n16638 = \s11_data_i[13]_pad  & n15106 ;
  assign n16639 = \s7_data_i[13]_pad  & n14837 ;
  assign n16640 = ~n16638 & ~n16639 ;
  assign n16641 = ~n16637 & n16640 ;
  assign n16642 = \s5_data_i[13]_pad  & n14829 ;
  assign n16643 = \s8_data_i[13]_pad  & n14841 ;
  assign n16644 = ~n16642 & ~n16643 ;
  assign n16645 = \s2_data_i[13]_pad  & n14816 ;
  assign n16646 = \s13_data_i[13]_pad  & n14805 ;
  assign n16647 = ~n16645 & ~n16646 ;
  assign n16648 = n16644 & n16647 ;
  assign n16649 = n16641 & n16648 ;
  assign n16650 = n16636 & n16649 ;
  assign n16651 = n16621 & n16650 ;
  assign n16652 = n2157 & n15377 ;
  assign n16653 = \s15_data_i[14]_pad  & n2157 ;
  assign n16654 = ~n2258 & n16653 ;
  assign n16655 = ~n16652 & ~n16654 ;
  assign n16656 = \s12_data_i[14]_pad  & n15102 ;
  assign n16657 = \s1_data_i[14]_pad  & n14658 ;
  assign n16658 = ~n16656 & ~n16657 ;
  assign n16659 = \s0_data_i[14]_pad  & n14582 ;
  assign n16660 = \s10_data_i[14]_pad  & n14797 ;
  assign n16661 = ~n16659 & ~n16660 ;
  assign n16662 = n16658 & n16661 ;
  assign n16663 = \s3_data_i[14]_pad  & n14820 ;
  assign n16664 = \s4_data_i[14]_pad  & n14825 ;
  assign n16665 = ~n16663 & ~n16664 ;
  assign n16666 = \s9_data_i[14]_pad  & n14845 ;
  assign n16667 = \s6_data_i[14]_pad  & n14833 ;
  assign n16668 = ~n16666 & ~n16667 ;
  assign n16669 = n16665 & n16668 ;
  assign n16670 = n16662 & n16669 ;
  assign n16671 = \s14_data_i[14]_pad  & n14809 ;
  assign n16672 = \s11_data_i[14]_pad  & n15106 ;
  assign n16673 = \s7_data_i[14]_pad  & n14837 ;
  assign n16674 = ~n16672 & ~n16673 ;
  assign n16675 = ~n16671 & n16674 ;
  assign n16676 = \s5_data_i[14]_pad  & n14829 ;
  assign n16677 = \s8_data_i[14]_pad  & n14841 ;
  assign n16678 = ~n16676 & ~n16677 ;
  assign n16679 = \s2_data_i[14]_pad  & n14816 ;
  assign n16680 = \s13_data_i[14]_pad  & n14805 ;
  assign n16681 = ~n16679 & ~n16680 ;
  assign n16682 = n16678 & n16681 ;
  assign n16683 = n16675 & n16682 ;
  assign n16684 = n16670 & n16683 ;
  assign n16685 = n16655 & n16684 ;
  assign n16686 = n2157 & n15414 ;
  assign n16687 = \s15_data_i[15]_pad  & n2157 ;
  assign n16688 = ~n2258 & n16687 ;
  assign n16689 = ~n16686 & ~n16688 ;
  assign n16690 = \s12_data_i[15]_pad  & n15102 ;
  assign n16691 = \s1_data_i[15]_pad  & n14658 ;
  assign n16692 = ~n16690 & ~n16691 ;
  assign n16693 = \s0_data_i[15]_pad  & n14582 ;
  assign n16694 = \s10_data_i[15]_pad  & n14797 ;
  assign n16695 = ~n16693 & ~n16694 ;
  assign n16696 = n16692 & n16695 ;
  assign n16697 = \s3_data_i[15]_pad  & n14820 ;
  assign n16698 = \s4_data_i[15]_pad  & n14825 ;
  assign n16699 = ~n16697 & ~n16698 ;
  assign n16700 = \s9_data_i[15]_pad  & n14845 ;
  assign n16701 = \s6_data_i[15]_pad  & n14833 ;
  assign n16702 = ~n16700 & ~n16701 ;
  assign n16703 = n16699 & n16702 ;
  assign n16704 = n16696 & n16703 ;
  assign n16705 = \s14_data_i[15]_pad  & n14809 ;
  assign n16706 = \s11_data_i[15]_pad  & n15106 ;
  assign n16707 = \s7_data_i[15]_pad  & n14837 ;
  assign n16708 = ~n16706 & ~n16707 ;
  assign n16709 = ~n16705 & n16708 ;
  assign n16710 = \s5_data_i[15]_pad  & n14829 ;
  assign n16711 = \s8_data_i[15]_pad  & n14841 ;
  assign n16712 = ~n16710 & ~n16711 ;
  assign n16713 = \s2_data_i[15]_pad  & n14816 ;
  assign n16714 = \s13_data_i[15]_pad  & n14805 ;
  assign n16715 = ~n16713 & ~n16714 ;
  assign n16716 = n16712 & n16715 ;
  assign n16717 = n16709 & n16716 ;
  assign n16718 = n16704 & n16717 ;
  assign n16719 = n16689 & n16718 ;
  assign n16720 = \s15_data_i[16]_pad  & n2157 ;
  assign n16721 = ~n2258 & n16720 ;
  assign n16722 = \s8_data_i[16]_pad  & n14841 ;
  assign n16723 = \s1_data_i[16]_pad  & n14658 ;
  assign n16724 = ~n16722 & ~n16723 ;
  assign n16725 = \s7_data_i[16]_pad  & n14837 ;
  assign n16726 = \s0_data_i[16]_pad  & n14582 ;
  assign n16727 = ~n16725 & ~n16726 ;
  assign n16728 = n16724 & n16727 ;
  assign n16729 = \s3_data_i[16]_pad  & n14820 ;
  assign n16730 = \s9_data_i[16]_pad  & n14845 ;
  assign n16731 = ~n16729 & ~n16730 ;
  assign n16732 = \s10_data_i[16]_pad  & n14797 ;
  assign n16733 = \s4_data_i[16]_pad  & n14825 ;
  assign n16734 = ~n16732 & ~n16733 ;
  assign n16735 = n16731 & n16734 ;
  assign n16736 = n16728 & n16735 ;
  assign n16737 = \s11_data_i[16]_pad  & n15106 ;
  assign n16738 = \s14_data_i[16]_pad  & n14809 ;
  assign n16739 = \s2_data_i[16]_pad  & n14816 ;
  assign n16740 = ~n16738 & ~n16739 ;
  assign n16741 = ~n16737 & n16740 ;
  assign n16742 = \s5_data_i[16]_pad  & n14829 ;
  assign n16743 = \s12_data_i[16]_pad  & n15102 ;
  assign n16744 = ~n16742 & ~n16743 ;
  assign n16745 = \s13_data_i[16]_pad  & n14805 ;
  assign n16746 = \s6_data_i[16]_pad  & n14833 ;
  assign n16747 = ~n16745 & ~n16746 ;
  assign n16748 = n16744 & n16747 ;
  assign n16749 = n16741 & n16748 ;
  assign n16750 = n16736 & n16749 ;
  assign n16751 = ~n16721 & n16750 ;
  assign n16752 = \s15_data_i[17]_pad  & n2157 ;
  assign n16753 = ~n2258 & n16752 ;
  assign n16754 = \s8_data_i[17]_pad  & n14841 ;
  assign n16755 = \s1_data_i[17]_pad  & n14658 ;
  assign n16756 = ~n16754 & ~n16755 ;
  assign n16757 = \s4_data_i[17]_pad  & n14825 ;
  assign n16758 = \s6_data_i[17]_pad  & n14833 ;
  assign n16759 = ~n16757 & ~n16758 ;
  assign n16760 = n16756 & n16759 ;
  assign n16761 = \s3_data_i[17]_pad  & n14820 ;
  assign n16762 = \s9_data_i[17]_pad  & n14845 ;
  assign n16763 = ~n16761 & ~n16762 ;
  assign n16764 = \s10_data_i[17]_pad  & n14797 ;
  assign n16765 = \s7_data_i[17]_pad  & n14837 ;
  assign n16766 = ~n16764 & ~n16765 ;
  assign n16767 = n16763 & n16766 ;
  assign n16768 = n16760 & n16767 ;
  assign n16769 = \s11_data_i[17]_pad  & n15106 ;
  assign n16770 = \s14_data_i[17]_pad  & n14809 ;
  assign n16771 = \s2_data_i[17]_pad  & n14816 ;
  assign n16772 = ~n16770 & ~n16771 ;
  assign n16773 = ~n16769 & n16772 ;
  assign n16774 = \s5_data_i[17]_pad  & n14829 ;
  assign n16775 = \s12_data_i[17]_pad  & n15102 ;
  assign n16776 = ~n16774 & ~n16775 ;
  assign n16777 = \s13_data_i[17]_pad  & n14805 ;
  assign n16778 = \s0_data_i[17]_pad  & n14582 ;
  assign n16779 = ~n16777 & ~n16778 ;
  assign n16780 = n16776 & n16779 ;
  assign n16781 = n16773 & n16780 ;
  assign n16782 = n16768 & n16781 ;
  assign n16783 = ~n16753 & n16782 ;
  assign n16784 = \s15_data_i[18]_pad  & n2157 ;
  assign n16785 = ~n2258 & n16784 ;
  assign n16786 = \s8_data_i[18]_pad  & n14841 ;
  assign n16787 = \s1_data_i[18]_pad  & n14658 ;
  assign n16788 = ~n16786 & ~n16787 ;
  assign n16789 = \s7_data_i[18]_pad  & n14837 ;
  assign n16790 = \s0_data_i[18]_pad  & n14582 ;
  assign n16791 = ~n16789 & ~n16790 ;
  assign n16792 = n16788 & n16791 ;
  assign n16793 = \s3_data_i[18]_pad  & n14820 ;
  assign n16794 = \s9_data_i[18]_pad  & n14845 ;
  assign n16795 = ~n16793 & ~n16794 ;
  assign n16796 = \s10_data_i[18]_pad  & n14797 ;
  assign n16797 = \s4_data_i[18]_pad  & n14825 ;
  assign n16798 = ~n16796 & ~n16797 ;
  assign n16799 = n16795 & n16798 ;
  assign n16800 = n16792 & n16799 ;
  assign n16801 = \s11_data_i[18]_pad  & n15106 ;
  assign n16802 = \s14_data_i[18]_pad  & n14809 ;
  assign n16803 = \s2_data_i[18]_pad  & n14816 ;
  assign n16804 = ~n16802 & ~n16803 ;
  assign n16805 = ~n16801 & n16804 ;
  assign n16806 = \s5_data_i[18]_pad  & n14829 ;
  assign n16807 = \s12_data_i[18]_pad  & n15102 ;
  assign n16808 = ~n16806 & ~n16807 ;
  assign n16809 = \s13_data_i[18]_pad  & n14805 ;
  assign n16810 = \s6_data_i[18]_pad  & n14833 ;
  assign n16811 = ~n16809 & ~n16810 ;
  assign n16812 = n16808 & n16811 ;
  assign n16813 = n16805 & n16812 ;
  assign n16814 = n16800 & n16813 ;
  assign n16815 = ~n16785 & n16814 ;
  assign n16816 = \s15_data_i[19]_pad  & n2157 ;
  assign n16817 = ~n2258 & n16816 ;
  assign n16818 = \s8_data_i[19]_pad  & n14841 ;
  assign n16819 = \s1_data_i[19]_pad  & n14658 ;
  assign n16820 = ~n16818 & ~n16819 ;
  assign n16821 = \s4_data_i[19]_pad  & n14825 ;
  assign n16822 = \s6_data_i[19]_pad  & n14833 ;
  assign n16823 = ~n16821 & ~n16822 ;
  assign n16824 = n16820 & n16823 ;
  assign n16825 = \s3_data_i[19]_pad  & n14820 ;
  assign n16826 = \s9_data_i[19]_pad  & n14845 ;
  assign n16827 = ~n16825 & ~n16826 ;
  assign n16828 = \s10_data_i[19]_pad  & n14797 ;
  assign n16829 = \s7_data_i[19]_pad  & n14837 ;
  assign n16830 = ~n16828 & ~n16829 ;
  assign n16831 = n16827 & n16830 ;
  assign n16832 = n16824 & n16831 ;
  assign n16833 = \s11_data_i[19]_pad  & n15106 ;
  assign n16834 = \s14_data_i[19]_pad  & n14809 ;
  assign n16835 = \s2_data_i[19]_pad  & n14816 ;
  assign n16836 = ~n16834 & ~n16835 ;
  assign n16837 = ~n16833 & n16836 ;
  assign n16838 = \s5_data_i[19]_pad  & n14829 ;
  assign n16839 = \s12_data_i[19]_pad  & n15102 ;
  assign n16840 = ~n16838 & ~n16839 ;
  assign n16841 = \s13_data_i[19]_pad  & n14805 ;
  assign n16842 = \s0_data_i[19]_pad  & n14582 ;
  assign n16843 = ~n16841 & ~n16842 ;
  assign n16844 = n16840 & n16843 ;
  assign n16845 = n16837 & n16844 ;
  assign n16846 = n16832 & n16845 ;
  assign n16847 = ~n16817 & n16846 ;
  assign n16848 = n2157 & n15579 ;
  assign n16849 = \s15_data_i[1]_pad  & n2157 ;
  assign n16850 = ~n2258 & n16849 ;
  assign n16851 = ~n16848 & ~n16850 ;
  assign n16852 = \s12_data_i[1]_pad  & n15102 ;
  assign n16853 = \s1_data_i[1]_pad  & n14658 ;
  assign n16854 = ~n16852 & ~n16853 ;
  assign n16855 = \s0_data_i[1]_pad  & n14582 ;
  assign n16856 = \s10_data_i[1]_pad  & n14797 ;
  assign n16857 = ~n16855 & ~n16856 ;
  assign n16858 = n16854 & n16857 ;
  assign n16859 = \s3_data_i[1]_pad  & n14820 ;
  assign n16860 = \s4_data_i[1]_pad  & n14825 ;
  assign n16861 = ~n16859 & ~n16860 ;
  assign n16862 = \s9_data_i[1]_pad  & n14845 ;
  assign n16863 = \s6_data_i[1]_pad  & n14833 ;
  assign n16864 = ~n16862 & ~n16863 ;
  assign n16865 = n16861 & n16864 ;
  assign n16866 = n16858 & n16865 ;
  assign n16867 = \s14_data_i[1]_pad  & n14809 ;
  assign n16868 = \s11_data_i[1]_pad  & n15106 ;
  assign n16869 = \s7_data_i[1]_pad  & n14837 ;
  assign n16870 = ~n16868 & ~n16869 ;
  assign n16871 = ~n16867 & n16870 ;
  assign n16872 = \s5_data_i[1]_pad  & n14829 ;
  assign n16873 = \s8_data_i[1]_pad  & n14841 ;
  assign n16874 = ~n16872 & ~n16873 ;
  assign n16875 = \s2_data_i[1]_pad  & n14816 ;
  assign n16876 = \s13_data_i[1]_pad  & n14805 ;
  assign n16877 = ~n16875 & ~n16876 ;
  assign n16878 = n16874 & n16877 ;
  assign n16879 = n16871 & n16878 ;
  assign n16880 = n16866 & n16879 ;
  assign n16881 = n16851 & n16880 ;
  assign n16882 = \s15_data_i[20]_pad  & n2157 ;
  assign n16883 = ~n2258 & n16882 ;
  assign n16884 = \s8_data_i[20]_pad  & n14841 ;
  assign n16885 = \s1_data_i[20]_pad  & n14658 ;
  assign n16886 = ~n16884 & ~n16885 ;
  assign n16887 = \s4_data_i[20]_pad  & n14825 ;
  assign n16888 = \s6_data_i[20]_pad  & n14833 ;
  assign n16889 = ~n16887 & ~n16888 ;
  assign n16890 = n16886 & n16889 ;
  assign n16891 = \s3_data_i[20]_pad  & n14820 ;
  assign n16892 = \s9_data_i[20]_pad  & n14845 ;
  assign n16893 = ~n16891 & ~n16892 ;
  assign n16894 = \s10_data_i[20]_pad  & n14797 ;
  assign n16895 = \s7_data_i[20]_pad  & n14837 ;
  assign n16896 = ~n16894 & ~n16895 ;
  assign n16897 = n16893 & n16896 ;
  assign n16898 = n16890 & n16897 ;
  assign n16899 = \s11_data_i[20]_pad  & n15106 ;
  assign n16900 = \s14_data_i[20]_pad  & n14809 ;
  assign n16901 = \s2_data_i[20]_pad  & n14816 ;
  assign n16902 = ~n16900 & ~n16901 ;
  assign n16903 = ~n16899 & n16902 ;
  assign n16904 = \s5_data_i[20]_pad  & n14829 ;
  assign n16905 = \s12_data_i[20]_pad  & n15102 ;
  assign n16906 = ~n16904 & ~n16905 ;
  assign n16907 = \s13_data_i[20]_pad  & n14805 ;
  assign n16908 = \s0_data_i[20]_pad  & n14582 ;
  assign n16909 = ~n16907 & ~n16908 ;
  assign n16910 = n16906 & n16909 ;
  assign n16911 = n16903 & n16910 ;
  assign n16912 = n16898 & n16911 ;
  assign n16913 = ~n16883 & n16912 ;
  assign n16914 = \s15_data_i[21]_pad  & n2157 ;
  assign n16915 = ~n2258 & n16914 ;
  assign n16916 = \s8_data_i[21]_pad  & n14841 ;
  assign n16917 = \s1_data_i[21]_pad  & n14658 ;
  assign n16918 = ~n16916 & ~n16917 ;
  assign n16919 = \s4_data_i[21]_pad  & n14825 ;
  assign n16920 = \s6_data_i[21]_pad  & n14833 ;
  assign n16921 = ~n16919 & ~n16920 ;
  assign n16922 = n16918 & n16921 ;
  assign n16923 = \s3_data_i[21]_pad  & n14820 ;
  assign n16924 = \s9_data_i[21]_pad  & n14845 ;
  assign n16925 = ~n16923 & ~n16924 ;
  assign n16926 = \s10_data_i[21]_pad  & n14797 ;
  assign n16927 = \s7_data_i[21]_pad  & n14837 ;
  assign n16928 = ~n16926 & ~n16927 ;
  assign n16929 = n16925 & n16928 ;
  assign n16930 = n16922 & n16929 ;
  assign n16931 = \s11_data_i[21]_pad  & n15106 ;
  assign n16932 = \s14_data_i[21]_pad  & n14809 ;
  assign n16933 = \s2_data_i[21]_pad  & n14816 ;
  assign n16934 = ~n16932 & ~n16933 ;
  assign n16935 = ~n16931 & n16934 ;
  assign n16936 = \s5_data_i[21]_pad  & n14829 ;
  assign n16937 = \s12_data_i[21]_pad  & n15102 ;
  assign n16938 = ~n16936 & ~n16937 ;
  assign n16939 = \s13_data_i[21]_pad  & n14805 ;
  assign n16940 = \s0_data_i[21]_pad  & n14582 ;
  assign n16941 = ~n16939 & ~n16940 ;
  assign n16942 = n16938 & n16941 ;
  assign n16943 = n16935 & n16942 ;
  assign n16944 = n16930 & n16943 ;
  assign n16945 = ~n16915 & n16944 ;
  assign n16946 = \s15_data_i[22]_pad  & n2157 ;
  assign n16947 = ~n2258 & n16946 ;
  assign n16948 = \s8_data_i[22]_pad  & n14841 ;
  assign n16949 = \s1_data_i[22]_pad  & n14658 ;
  assign n16950 = ~n16948 & ~n16949 ;
  assign n16951 = \s4_data_i[22]_pad  & n14825 ;
  assign n16952 = \s6_data_i[22]_pad  & n14833 ;
  assign n16953 = ~n16951 & ~n16952 ;
  assign n16954 = n16950 & n16953 ;
  assign n16955 = \s3_data_i[22]_pad  & n14820 ;
  assign n16956 = \s9_data_i[22]_pad  & n14845 ;
  assign n16957 = ~n16955 & ~n16956 ;
  assign n16958 = \s10_data_i[22]_pad  & n14797 ;
  assign n16959 = \s7_data_i[22]_pad  & n14837 ;
  assign n16960 = ~n16958 & ~n16959 ;
  assign n16961 = n16957 & n16960 ;
  assign n16962 = n16954 & n16961 ;
  assign n16963 = \s11_data_i[22]_pad  & n15106 ;
  assign n16964 = \s14_data_i[22]_pad  & n14809 ;
  assign n16965 = \s2_data_i[22]_pad  & n14816 ;
  assign n16966 = ~n16964 & ~n16965 ;
  assign n16967 = ~n16963 & n16966 ;
  assign n16968 = \s5_data_i[22]_pad  & n14829 ;
  assign n16969 = \s12_data_i[22]_pad  & n15102 ;
  assign n16970 = ~n16968 & ~n16969 ;
  assign n16971 = \s13_data_i[22]_pad  & n14805 ;
  assign n16972 = \s0_data_i[22]_pad  & n14582 ;
  assign n16973 = ~n16971 & ~n16972 ;
  assign n16974 = n16970 & n16973 ;
  assign n16975 = n16967 & n16974 ;
  assign n16976 = n16962 & n16975 ;
  assign n16977 = ~n16947 & n16976 ;
  assign n16978 = \s15_data_i[23]_pad  & n2157 ;
  assign n16979 = ~n2258 & n16978 ;
  assign n16980 = \s12_data_i[23]_pad  & n15102 ;
  assign n16981 = \s1_data_i[23]_pad  & n14658 ;
  assign n16982 = ~n16980 & ~n16981 ;
  assign n16983 = \s4_data_i[23]_pad  & n14825 ;
  assign n16984 = \s6_data_i[23]_pad  & n14833 ;
  assign n16985 = ~n16983 & ~n16984 ;
  assign n16986 = n16982 & n16985 ;
  assign n16987 = \s3_data_i[23]_pad  & n14820 ;
  assign n16988 = \s9_data_i[23]_pad  & n14845 ;
  assign n16989 = ~n16987 & ~n16988 ;
  assign n16990 = \s10_data_i[23]_pad  & n14797 ;
  assign n16991 = \s7_data_i[23]_pad  & n14837 ;
  assign n16992 = ~n16990 & ~n16991 ;
  assign n16993 = n16989 & n16992 ;
  assign n16994 = n16986 & n16993 ;
  assign n16995 = \s14_data_i[23]_pad  & n14809 ;
  assign n16996 = \s11_data_i[23]_pad  & n15106 ;
  assign n16997 = \s2_data_i[23]_pad  & n14816 ;
  assign n16998 = ~n16996 & ~n16997 ;
  assign n16999 = ~n16995 & n16998 ;
  assign n17000 = \s5_data_i[23]_pad  & n14829 ;
  assign n17001 = \s8_data_i[23]_pad  & n14841 ;
  assign n17002 = ~n17000 & ~n17001 ;
  assign n17003 = \s13_data_i[23]_pad  & n14805 ;
  assign n17004 = \s0_data_i[23]_pad  & n14582 ;
  assign n17005 = ~n17003 & ~n17004 ;
  assign n17006 = n17002 & n17005 ;
  assign n17007 = n16999 & n17006 ;
  assign n17008 = n16994 & n17007 ;
  assign n17009 = ~n16979 & n17008 ;
  assign n17010 = \s15_data_i[24]_pad  & n2157 ;
  assign n17011 = ~n2258 & n17010 ;
  assign n17012 = \s8_data_i[24]_pad  & n14841 ;
  assign n17013 = \s1_data_i[24]_pad  & n14658 ;
  assign n17014 = ~n17012 & ~n17013 ;
  assign n17015 = \s4_data_i[24]_pad  & n14825 ;
  assign n17016 = \s6_data_i[24]_pad  & n14833 ;
  assign n17017 = ~n17015 & ~n17016 ;
  assign n17018 = n17014 & n17017 ;
  assign n17019 = \s3_data_i[24]_pad  & n14820 ;
  assign n17020 = \s9_data_i[24]_pad  & n14845 ;
  assign n17021 = ~n17019 & ~n17020 ;
  assign n17022 = \s10_data_i[24]_pad  & n14797 ;
  assign n17023 = \s7_data_i[24]_pad  & n14837 ;
  assign n17024 = ~n17022 & ~n17023 ;
  assign n17025 = n17021 & n17024 ;
  assign n17026 = n17018 & n17025 ;
  assign n17027 = \s11_data_i[24]_pad  & n15106 ;
  assign n17028 = \s14_data_i[24]_pad  & n14809 ;
  assign n17029 = \s2_data_i[24]_pad  & n14816 ;
  assign n17030 = ~n17028 & ~n17029 ;
  assign n17031 = ~n17027 & n17030 ;
  assign n17032 = \s5_data_i[24]_pad  & n14829 ;
  assign n17033 = \s12_data_i[24]_pad  & n15102 ;
  assign n17034 = ~n17032 & ~n17033 ;
  assign n17035 = \s13_data_i[24]_pad  & n14805 ;
  assign n17036 = \s0_data_i[24]_pad  & n14582 ;
  assign n17037 = ~n17035 & ~n17036 ;
  assign n17038 = n17034 & n17037 ;
  assign n17039 = n17031 & n17038 ;
  assign n17040 = n17026 & n17039 ;
  assign n17041 = ~n17011 & n17040 ;
  assign n17042 = \s15_data_i[25]_pad  & n2157 ;
  assign n17043 = ~n2258 & n17042 ;
  assign n17044 = \s8_data_i[25]_pad  & n14841 ;
  assign n17045 = \s1_data_i[25]_pad  & n14658 ;
  assign n17046 = ~n17044 & ~n17045 ;
  assign n17047 = \s4_data_i[25]_pad  & n14825 ;
  assign n17048 = \s6_data_i[25]_pad  & n14833 ;
  assign n17049 = ~n17047 & ~n17048 ;
  assign n17050 = n17046 & n17049 ;
  assign n17051 = \s3_data_i[25]_pad  & n14820 ;
  assign n17052 = \s9_data_i[25]_pad  & n14845 ;
  assign n17053 = ~n17051 & ~n17052 ;
  assign n17054 = \s10_data_i[25]_pad  & n14797 ;
  assign n17055 = \s7_data_i[25]_pad  & n14837 ;
  assign n17056 = ~n17054 & ~n17055 ;
  assign n17057 = n17053 & n17056 ;
  assign n17058 = n17050 & n17057 ;
  assign n17059 = \s11_data_i[25]_pad  & n15106 ;
  assign n17060 = \s14_data_i[25]_pad  & n14809 ;
  assign n17061 = \s2_data_i[25]_pad  & n14816 ;
  assign n17062 = ~n17060 & ~n17061 ;
  assign n17063 = ~n17059 & n17062 ;
  assign n17064 = \s5_data_i[25]_pad  & n14829 ;
  assign n17065 = \s12_data_i[25]_pad  & n15102 ;
  assign n17066 = ~n17064 & ~n17065 ;
  assign n17067 = \s13_data_i[25]_pad  & n14805 ;
  assign n17068 = \s0_data_i[25]_pad  & n14582 ;
  assign n17069 = ~n17067 & ~n17068 ;
  assign n17070 = n17066 & n17069 ;
  assign n17071 = n17063 & n17070 ;
  assign n17072 = n17058 & n17071 ;
  assign n17073 = ~n17043 & n17072 ;
  assign n17074 = \s15_data_i[26]_pad  & n2157 ;
  assign n17075 = ~n2258 & n17074 ;
  assign n17076 = \s8_data_i[26]_pad  & n14841 ;
  assign n17077 = \s1_data_i[26]_pad  & n14658 ;
  assign n17078 = ~n17076 & ~n17077 ;
  assign n17079 = \s4_data_i[26]_pad  & n14825 ;
  assign n17080 = \s6_data_i[26]_pad  & n14833 ;
  assign n17081 = ~n17079 & ~n17080 ;
  assign n17082 = n17078 & n17081 ;
  assign n17083 = \s3_data_i[26]_pad  & n14820 ;
  assign n17084 = \s9_data_i[26]_pad  & n14845 ;
  assign n17085 = ~n17083 & ~n17084 ;
  assign n17086 = \s10_data_i[26]_pad  & n14797 ;
  assign n17087 = \s7_data_i[26]_pad  & n14837 ;
  assign n17088 = ~n17086 & ~n17087 ;
  assign n17089 = n17085 & n17088 ;
  assign n17090 = n17082 & n17089 ;
  assign n17091 = \s11_data_i[26]_pad  & n15106 ;
  assign n17092 = \s14_data_i[26]_pad  & n14809 ;
  assign n17093 = \s2_data_i[26]_pad  & n14816 ;
  assign n17094 = ~n17092 & ~n17093 ;
  assign n17095 = ~n17091 & n17094 ;
  assign n17096 = \s5_data_i[26]_pad  & n14829 ;
  assign n17097 = \s12_data_i[26]_pad  & n15102 ;
  assign n17098 = ~n17096 & ~n17097 ;
  assign n17099 = \s13_data_i[26]_pad  & n14805 ;
  assign n17100 = \s0_data_i[26]_pad  & n14582 ;
  assign n17101 = ~n17099 & ~n17100 ;
  assign n17102 = n17098 & n17101 ;
  assign n17103 = n17095 & n17102 ;
  assign n17104 = n17090 & n17103 ;
  assign n17105 = ~n17075 & n17104 ;
  assign n17106 = \s15_data_i[27]_pad  & n2157 ;
  assign n17107 = ~n2258 & n17106 ;
  assign n17108 = \s8_data_i[27]_pad  & n14841 ;
  assign n17109 = \s1_data_i[27]_pad  & n14658 ;
  assign n17110 = ~n17108 & ~n17109 ;
  assign n17111 = \s4_data_i[27]_pad  & n14825 ;
  assign n17112 = \s6_data_i[27]_pad  & n14833 ;
  assign n17113 = ~n17111 & ~n17112 ;
  assign n17114 = n17110 & n17113 ;
  assign n17115 = \s3_data_i[27]_pad  & n14820 ;
  assign n17116 = \s9_data_i[27]_pad  & n14845 ;
  assign n17117 = ~n17115 & ~n17116 ;
  assign n17118 = \s10_data_i[27]_pad  & n14797 ;
  assign n17119 = \s7_data_i[27]_pad  & n14837 ;
  assign n17120 = ~n17118 & ~n17119 ;
  assign n17121 = n17117 & n17120 ;
  assign n17122 = n17114 & n17121 ;
  assign n17123 = \s11_data_i[27]_pad  & n15106 ;
  assign n17124 = \s14_data_i[27]_pad  & n14809 ;
  assign n17125 = \s2_data_i[27]_pad  & n14816 ;
  assign n17126 = ~n17124 & ~n17125 ;
  assign n17127 = ~n17123 & n17126 ;
  assign n17128 = \s5_data_i[27]_pad  & n14829 ;
  assign n17129 = \s12_data_i[27]_pad  & n15102 ;
  assign n17130 = ~n17128 & ~n17129 ;
  assign n17131 = \s13_data_i[27]_pad  & n14805 ;
  assign n17132 = \s0_data_i[27]_pad  & n14582 ;
  assign n17133 = ~n17131 & ~n17132 ;
  assign n17134 = n17130 & n17133 ;
  assign n17135 = n17127 & n17134 ;
  assign n17136 = n17122 & n17135 ;
  assign n17137 = ~n17107 & n17136 ;
  assign n17138 = \s15_data_i[28]_pad  & n2157 ;
  assign n17139 = ~n2258 & n17138 ;
  assign n17140 = \s8_data_i[28]_pad  & n14841 ;
  assign n17141 = \s1_data_i[28]_pad  & n14658 ;
  assign n17142 = ~n17140 & ~n17141 ;
  assign n17143 = \s4_data_i[28]_pad  & n14825 ;
  assign n17144 = \s9_data_i[28]_pad  & n14845 ;
  assign n17145 = ~n17143 & ~n17144 ;
  assign n17146 = n17142 & n17145 ;
  assign n17147 = \s3_data_i[28]_pad  & n14820 ;
  assign n17148 = \s6_data_i[28]_pad  & n14833 ;
  assign n17149 = ~n17147 & ~n17148 ;
  assign n17150 = \s7_data_i[28]_pad  & n14837 ;
  assign n17151 = \s10_data_i[28]_pad  & n14797 ;
  assign n17152 = ~n17150 & ~n17151 ;
  assign n17153 = n17149 & n17152 ;
  assign n17154 = n17146 & n17153 ;
  assign n17155 = \s11_data_i[28]_pad  & n15106 ;
  assign n17156 = \s14_data_i[28]_pad  & n14809 ;
  assign n17157 = \s2_data_i[28]_pad  & n14816 ;
  assign n17158 = ~n17156 & ~n17157 ;
  assign n17159 = ~n17155 & n17158 ;
  assign n17160 = \s5_data_i[28]_pad  & n14829 ;
  assign n17161 = \s12_data_i[28]_pad  & n15102 ;
  assign n17162 = ~n17160 & ~n17161 ;
  assign n17163 = \s13_data_i[28]_pad  & n14805 ;
  assign n17164 = \s0_data_i[28]_pad  & n14582 ;
  assign n17165 = ~n17163 & ~n17164 ;
  assign n17166 = n17162 & n17165 ;
  assign n17167 = n17159 & n17166 ;
  assign n17168 = n17154 & n17167 ;
  assign n17169 = ~n17139 & n17168 ;
  assign n17170 = \s15_data_i[29]_pad  & n2157 ;
  assign n17171 = ~n2258 & n17170 ;
  assign n17172 = \s8_data_i[29]_pad  & n14841 ;
  assign n17173 = \s1_data_i[29]_pad  & n14658 ;
  assign n17174 = ~n17172 & ~n17173 ;
  assign n17175 = \s4_data_i[29]_pad  & n14825 ;
  assign n17176 = \s6_data_i[29]_pad  & n14833 ;
  assign n17177 = ~n17175 & ~n17176 ;
  assign n17178 = n17174 & n17177 ;
  assign n17179 = \s3_data_i[29]_pad  & n14820 ;
  assign n17180 = \s9_data_i[29]_pad  & n14845 ;
  assign n17181 = ~n17179 & ~n17180 ;
  assign n17182 = \s10_data_i[29]_pad  & n14797 ;
  assign n17183 = \s7_data_i[29]_pad  & n14837 ;
  assign n17184 = ~n17182 & ~n17183 ;
  assign n17185 = n17181 & n17184 ;
  assign n17186 = n17178 & n17185 ;
  assign n17187 = \s11_data_i[29]_pad  & n15106 ;
  assign n17188 = \s14_data_i[29]_pad  & n14809 ;
  assign n17189 = \s2_data_i[29]_pad  & n14816 ;
  assign n17190 = ~n17188 & ~n17189 ;
  assign n17191 = ~n17187 & n17190 ;
  assign n17192 = \s5_data_i[29]_pad  & n14829 ;
  assign n17193 = \s12_data_i[29]_pad  & n15102 ;
  assign n17194 = ~n17192 & ~n17193 ;
  assign n17195 = \s13_data_i[29]_pad  & n14805 ;
  assign n17196 = \s0_data_i[29]_pad  & n14582 ;
  assign n17197 = ~n17195 & ~n17196 ;
  assign n17198 = n17194 & n17197 ;
  assign n17199 = n17191 & n17198 ;
  assign n17200 = n17186 & n17199 ;
  assign n17201 = ~n17171 & n17200 ;
  assign n17202 = n2157 & n15936 ;
  assign n17203 = \s15_data_i[2]_pad  & n2157 ;
  assign n17204 = ~n2258 & n17203 ;
  assign n17205 = ~n17202 & ~n17204 ;
  assign n17206 = \s12_data_i[2]_pad  & n15102 ;
  assign n17207 = \s1_data_i[2]_pad  & n14658 ;
  assign n17208 = ~n17206 & ~n17207 ;
  assign n17209 = \s0_data_i[2]_pad  & n14582 ;
  assign n17210 = \s10_data_i[2]_pad  & n14797 ;
  assign n17211 = ~n17209 & ~n17210 ;
  assign n17212 = n17208 & n17211 ;
  assign n17213 = \s3_data_i[2]_pad  & n14820 ;
  assign n17214 = \s4_data_i[2]_pad  & n14825 ;
  assign n17215 = ~n17213 & ~n17214 ;
  assign n17216 = \s9_data_i[2]_pad  & n14845 ;
  assign n17217 = \s6_data_i[2]_pad  & n14833 ;
  assign n17218 = ~n17216 & ~n17217 ;
  assign n17219 = n17215 & n17218 ;
  assign n17220 = n17212 & n17219 ;
  assign n17221 = \s14_data_i[2]_pad  & n14809 ;
  assign n17222 = \s11_data_i[2]_pad  & n15106 ;
  assign n17223 = \s7_data_i[2]_pad  & n14837 ;
  assign n17224 = ~n17222 & ~n17223 ;
  assign n17225 = ~n17221 & n17224 ;
  assign n17226 = \s5_data_i[2]_pad  & n14829 ;
  assign n17227 = \s8_data_i[2]_pad  & n14841 ;
  assign n17228 = ~n17226 & ~n17227 ;
  assign n17229 = \s2_data_i[2]_pad  & n14816 ;
  assign n17230 = \s13_data_i[2]_pad  & n14805 ;
  assign n17231 = ~n17229 & ~n17230 ;
  assign n17232 = n17228 & n17231 ;
  assign n17233 = n17225 & n17232 ;
  assign n17234 = n17220 & n17233 ;
  assign n17235 = n17205 & n17234 ;
  assign n17236 = \s15_data_i[30]_pad  & n2157 ;
  assign n17237 = ~n2258 & n17236 ;
  assign n17238 = \s8_data_i[30]_pad  & n14841 ;
  assign n17239 = \s1_data_i[30]_pad  & n14658 ;
  assign n17240 = ~n17238 & ~n17239 ;
  assign n17241 = \s4_data_i[30]_pad  & n14825 ;
  assign n17242 = \s6_data_i[30]_pad  & n14833 ;
  assign n17243 = ~n17241 & ~n17242 ;
  assign n17244 = n17240 & n17243 ;
  assign n17245 = \s3_data_i[30]_pad  & n14820 ;
  assign n17246 = \s9_data_i[30]_pad  & n14845 ;
  assign n17247 = ~n17245 & ~n17246 ;
  assign n17248 = \s10_data_i[30]_pad  & n14797 ;
  assign n17249 = \s7_data_i[30]_pad  & n14837 ;
  assign n17250 = ~n17248 & ~n17249 ;
  assign n17251 = n17247 & n17250 ;
  assign n17252 = n17244 & n17251 ;
  assign n17253 = \s11_data_i[30]_pad  & n15106 ;
  assign n17254 = \s14_data_i[30]_pad  & n14809 ;
  assign n17255 = \s2_data_i[30]_pad  & n14816 ;
  assign n17256 = ~n17254 & ~n17255 ;
  assign n17257 = ~n17253 & n17256 ;
  assign n17258 = \s5_data_i[30]_pad  & n14829 ;
  assign n17259 = \s12_data_i[30]_pad  & n15102 ;
  assign n17260 = ~n17258 & ~n17259 ;
  assign n17261 = \s13_data_i[30]_pad  & n14805 ;
  assign n17262 = \s0_data_i[30]_pad  & n14582 ;
  assign n17263 = ~n17261 & ~n17262 ;
  assign n17264 = n17260 & n17263 ;
  assign n17265 = n17257 & n17264 ;
  assign n17266 = n17252 & n17265 ;
  assign n17267 = ~n17237 & n17266 ;
  assign n17268 = \s15_data_i[31]_pad  & n2157 ;
  assign n17269 = ~n2258 & n17268 ;
  assign n17270 = \s8_data_i[31]_pad  & n14841 ;
  assign n17271 = \s1_data_i[31]_pad  & n14658 ;
  assign n17272 = ~n17270 & ~n17271 ;
  assign n17273 = \s4_data_i[31]_pad  & n14825 ;
  assign n17274 = \s6_data_i[31]_pad  & n14833 ;
  assign n17275 = ~n17273 & ~n17274 ;
  assign n17276 = n17272 & n17275 ;
  assign n17277 = \s3_data_i[31]_pad  & n14820 ;
  assign n17278 = \s9_data_i[31]_pad  & n14845 ;
  assign n17279 = ~n17277 & ~n17278 ;
  assign n17280 = \s10_data_i[31]_pad  & n14797 ;
  assign n17281 = \s7_data_i[31]_pad  & n14837 ;
  assign n17282 = ~n17280 & ~n17281 ;
  assign n17283 = n17279 & n17282 ;
  assign n17284 = n17276 & n17283 ;
  assign n17285 = \s11_data_i[31]_pad  & n15106 ;
  assign n17286 = \s14_data_i[31]_pad  & n14809 ;
  assign n17287 = \s2_data_i[31]_pad  & n14816 ;
  assign n17288 = ~n17286 & ~n17287 ;
  assign n17289 = ~n17285 & n17288 ;
  assign n17290 = \s5_data_i[31]_pad  & n14829 ;
  assign n17291 = \s12_data_i[31]_pad  & n15102 ;
  assign n17292 = ~n17290 & ~n17291 ;
  assign n17293 = \s13_data_i[31]_pad  & n14805 ;
  assign n17294 = \s0_data_i[31]_pad  & n14582 ;
  assign n17295 = ~n17293 & ~n17294 ;
  assign n17296 = n17292 & n17295 ;
  assign n17297 = n17289 & n17296 ;
  assign n17298 = n17284 & n17297 ;
  assign n17299 = ~n17269 & n17298 ;
  assign n17300 = n2157 & n16037 ;
  assign n17301 = \s15_data_i[3]_pad  & n2157 ;
  assign n17302 = ~n2258 & n17301 ;
  assign n17303 = ~n17300 & ~n17302 ;
  assign n17304 = \s12_data_i[3]_pad  & n15102 ;
  assign n17305 = \s1_data_i[3]_pad  & n14658 ;
  assign n17306 = ~n17304 & ~n17305 ;
  assign n17307 = \s7_data_i[3]_pad  & n14837 ;
  assign n17308 = \s9_data_i[3]_pad  & n14845 ;
  assign n17309 = ~n17307 & ~n17308 ;
  assign n17310 = n17306 & n17309 ;
  assign n17311 = \s3_data_i[3]_pad  & n14820 ;
  assign n17312 = \s6_data_i[3]_pad  & n14833 ;
  assign n17313 = ~n17311 & ~n17312 ;
  assign n17314 = \s10_data_i[3]_pad  & n14797 ;
  assign n17315 = \s13_data_i[3]_pad  & n14805 ;
  assign n17316 = ~n17314 & ~n17315 ;
  assign n17317 = n17313 & n17316 ;
  assign n17318 = n17310 & n17317 ;
  assign n17319 = \s14_data_i[3]_pad  & n14809 ;
  assign n17320 = \s11_data_i[3]_pad  & n15106 ;
  assign n17321 = \s2_data_i[3]_pad  & n14816 ;
  assign n17322 = ~n17320 & ~n17321 ;
  assign n17323 = ~n17319 & n17322 ;
  assign n17324 = \s5_data_i[3]_pad  & n14829 ;
  assign n17325 = \s8_data_i[3]_pad  & n14841 ;
  assign n17326 = ~n17324 & ~n17325 ;
  assign n17327 = \s4_data_i[3]_pad  & n14825 ;
  assign n17328 = \s0_data_i[3]_pad  & n14582 ;
  assign n17329 = ~n17327 & ~n17328 ;
  assign n17330 = n17326 & n17329 ;
  assign n17331 = n17323 & n17330 ;
  assign n17332 = n17318 & n17331 ;
  assign n17333 = n17303 & n17332 ;
  assign n17334 = n2157 & n16074 ;
  assign n17335 = \s15_data_i[4]_pad  & n2157 ;
  assign n17336 = ~n2258 & n17335 ;
  assign n17337 = ~n17334 & ~n17336 ;
  assign n17338 = \s12_data_i[4]_pad  & n15102 ;
  assign n17339 = \s1_data_i[4]_pad  & n14658 ;
  assign n17340 = ~n17338 & ~n17339 ;
  assign n17341 = \s0_data_i[4]_pad  & n14582 ;
  assign n17342 = \s10_data_i[4]_pad  & n14797 ;
  assign n17343 = ~n17341 & ~n17342 ;
  assign n17344 = n17340 & n17343 ;
  assign n17345 = \s3_data_i[4]_pad  & n14820 ;
  assign n17346 = \s4_data_i[4]_pad  & n14825 ;
  assign n17347 = ~n17345 & ~n17346 ;
  assign n17348 = \s9_data_i[4]_pad  & n14845 ;
  assign n17349 = \s6_data_i[4]_pad  & n14833 ;
  assign n17350 = ~n17348 & ~n17349 ;
  assign n17351 = n17347 & n17350 ;
  assign n17352 = n17344 & n17351 ;
  assign n17353 = \s14_data_i[4]_pad  & n14809 ;
  assign n17354 = \s11_data_i[4]_pad  & n15106 ;
  assign n17355 = \s7_data_i[4]_pad  & n14837 ;
  assign n17356 = ~n17354 & ~n17355 ;
  assign n17357 = ~n17353 & n17356 ;
  assign n17358 = \s5_data_i[4]_pad  & n14829 ;
  assign n17359 = \s8_data_i[4]_pad  & n14841 ;
  assign n17360 = ~n17358 & ~n17359 ;
  assign n17361 = \s2_data_i[4]_pad  & n14816 ;
  assign n17362 = \s13_data_i[4]_pad  & n14805 ;
  assign n17363 = ~n17361 & ~n17362 ;
  assign n17364 = n17360 & n17363 ;
  assign n17365 = n17357 & n17364 ;
  assign n17366 = n17352 & n17365 ;
  assign n17367 = n17337 & n17366 ;
  assign n17368 = n2157 & n16111 ;
  assign n17369 = \s15_data_i[5]_pad  & n2157 ;
  assign n17370 = ~n2258 & n17369 ;
  assign n17371 = ~n17368 & ~n17370 ;
  assign n17372 = \s14_data_i[5]_pad  & n14809 ;
  assign n17373 = \s1_data_i[5]_pad  & n14658 ;
  assign n17374 = ~n17372 & ~n17373 ;
  assign n17375 = \s10_data_i[5]_pad  & n14797 ;
  assign n17376 = \s7_data_i[5]_pad  & n14837 ;
  assign n17377 = ~n17375 & ~n17376 ;
  assign n17378 = n17374 & n17377 ;
  assign n17379 = \s5_data_i[5]_pad  & n14829 ;
  assign n17380 = \s2_data_i[5]_pad  & n14816 ;
  assign n17381 = ~n17379 & ~n17380 ;
  assign n17382 = \s6_data_i[5]_pad  & n14833 ;
  assign n17383 = \s0_data_i[5]_pad  & n14582 ;
  assign n17384 = ~n17382 & ~n17383 ;
  assign n17385 = n17381 & n17384 ;
  assign n17386 = n17378 & n17385 ;
  assign n17387 = \s11_data_i[5]_pad  & n15106 ;
  assign n17388 = \s8_data_i[5]_pad  & n14841 ;
  assign n17389 = \s4_data_i[5]_pad  & n14825 ;
  assign n17390 = ~n17388 & ~n17389 ;
  assign n17391 = ~n17387 & n17390 ;
  assign n17392 = \s3_data_i[5]_pad  & n14820 ;
  assign n17393 = \s12_data_i[5]_pad  & n15102 ;
  assign n17394 = ~n17392 & ~n17393 ;
  assign n17395 = \s13_data_i[5]_pad  & n14805 ;
  assign n17396 = \s9_data_i[5]_pad  & n14845 ;
  assign n17397 = ~n17395 & ~n17396 ;
  assign n17398 = n17394 & n17397 ;
  assign n17399 = n17391 & n17398 ;
  assign n17400 = n17386 & n17399 ;
  assign n17401 = n17371 & n17400 ;
  assign n17402 = n2157 & n16148 ;
  assign n17403 = \s15_data_i[6]_pad  & n2157 ;
  assign n17404 = ~n2258 & n17403 ;
  assign n17405 = ~n17402 & ~n17404 ;
  assign n17406 = \s12_data_i[6]_pad  & n15102 ;
  assign n17407 = \s1_data_i[6]_pad  & n14658 ;
  assign n17408 = ~n17406 & ~n17407 ;
  assign n17409 = \s0_data_i[6]_pad  & n14582 ;
  assign n17410 = \s10_data_i[6]_pad  & n14797 ;
  assign n17411 = ~n17409 & ~n17410 ;
  assign n17412 = n17408 & n17411 ;
  assign n17413 = \s3_data_i[6]_pad  & n14820 ;
  assign n17414 = \s4_data_i[6]_pad  & n14825 ;
  assign n17415 = ~n17413 & ~n17414 ;
  assign n17416 = \s9_data_i[6]_pad  & n14845 ;
  assign n17417 = \s6_data_i[6]_pad  & n14833 ;
  assign n17418 = ~n17416 & ~n17417 ;
  assign n17419 = n17415 & n17418 ;
  assign n17420 = n17412 & n17419 ;
  assign n17421 = \s14_data_i[6]_pad  & n14809 ;
  assign n17422 = \s11_data_i[6]_pad  & n15106 ;
  assign n17423 = \s7_data_i[6]_pad  & n14837 ;
  assign n17424 = ~n17422 & ~n17423 ;
  assign n17425 = ~n17421 & n17424 ;
  assign n17426 = \s5_data_i[6]_pad  & n14829 ;
  assign n17427 = \s8_data_i[6]_pad  & n14841 ;
  assign n17428 = ~n17426 & ~n17427 ;
  assign n17429 = \s2_data_i[6]_pad  & n14816 ;
  assign n17430 = \s13_data_i[6]_pad  & n14805 ;
  assign n17431 = ~n17429 & ~n17430 ;
  assign n17432 = n17428 & n17431 ;
  assign n17433 = n17425 & n17432 ;
  assign n17434 = n17420 & n17433 ;
  assign n17435 = n17405 & n17434 ;
  assign n17436 = n2157 & n16185 ;
  assign n17437 = \s15_data_i[7]_pad  & n2157 ;
  assign n17438 = ~n2258 & n17437 ;
  assign n17439 = ~n17436 & ~n17438 ;
  assign n17440 = \s12_data_i[7]_pad  & n15102 ;
  assign n17441 = \s1_data_i[7]_pad  & n14658 ;
  assign n17442 = ~n17440 & ~n17441 ;
  assign n17443 = \s0_data_i[7]_pad  & n14582 ;
  assign n17444 = \s10_data_i[7]_pad  & n14797 ;
  assign n17445 = ~n17443 & ~n17444 ;
  assign n17446 = n17442 & n17445 ;
  assign n17447 = \s3_data_i[7]_pad  & n14820 ;
  assign n17448 = \s4_data_i[7]_pad  & n14825 ;
  assign n17449 = ~n17447 & ~n17448 ;
  assign n17450 = \s9_data_i[7]_pad  & n14845 ;
  assign n17451 = \s6_data_i[7]_pad  & n14833 ;
  assign n17452 = ~n17450 & ~n17451 ;
  assign n17453 = n17449 & n17452 ;
  assign n17454 = n17446 & n17453 ;
  assign n17455 = \s14_data_i[7]_pad  & n14809 ;
  assign n17456 = \s11_data_i[7]_pad  & n15106 ;
  assign n17457 = \s7_data_i[7]_pad  & n14837 ;
  assign n17458 = ~n17456 & ~n17457 ;
  assign n17459 = ~n17455 & n17458 ;
  assign n17460 = \s5_data_i[7]_pad  & n14829 ;
  assign n17461 = \s8_data_i[7]_pad  & n14841 ;
  assign n17462 = ~n17460 & ~n17461 ;
  assign n17463 = \s2_data_i[7]_pad  & n14816 ;
  assign n17464 = \s13_data_i[7]_pad  & n14805 ;
  assign n17465 = ~n17463 & ~n17464 ;
  assign n17466 = n17462 & n17465 ;
  assign n17467 = n17459 & n17466 ;
  assign n17468 = n17454 & n17467 ;
  assign n17469 = n17439 & n17468 ;
  assign n17470 = n2157 & n16222 ;
  assign n17471 = \s15_data_i[8]_pad  & n2157 ;
  assign n17472 = ~n2258 & n17471 ;
  assign n17473 = ~n17470 & ~n17472 ;
  assign n17474 = \s12_data_i[8]_pad  & n15102 ;
  assign n17475 = \s1_data_i[8]_pad  & n14658 ;
  assign n17476 = ~n17474 & ~n17475 ;
  assign n17477 = \s0_data_i[8]_pad  & n14582 ;
  assign n17478 = \s10_data_i[8]_pad  & n14797 ;
  assign n17479 = ~n17477 & ~n17478 ;
  assign n17480 = n17476 & n17479 ;
  assign n17481 = \s3_data_i[8]_pad  & n14820 ;
  assign n17482 = \s4_data_i[8]_pad  & n14825 ;
  assign n17483 = ~n17481 & ~n17482 ;
  assign n17484 = \s9_data_i[8]_pad  & n14845 ;
  assign n17485 = \s6_data_i[8]_pad  & n14833 ;
  assign n17486 = ~n17484 & ~n17485 ;
  assign n17487 = n17483 & n17486 ;
  assign n17488 = n17480 & n17487 ;
  assign n17489 = \s14_data_i[8]_pad  & n14809 ;
  assign n17490 = \s11_data_i[8]_pad  & n15106 ;
  assign n17491 = \s7_data_i[8]_pad  & n14837 ;
  assign n17492 = ~n17490 & ~n17491 ;
  assign n17493 = ~n17489 & n17492 ;
  assign n17494 = \s5_data_i[8]_pad  & n14829 ;
  assign n17495 = \s8_data_i[8]_pad  & n14841 ;
  assign n17496 = ~n17494 & ~n17495 ;
  assign n17497 = \s2_data_i[8]_pad  & n14816 ;
  assign n17498 = \s13_data_i[8]_pad  & n14805 ;
  assign n17499 = ~n17497 & ~n17498 ;
  assign n17500 = n17496 & n17499 ;
  assign n17501 = n17493 & n17500 ;
  assign n17502 = n17488 & n17501 ;
  assign n17503 = n17473 & n17502 ;
  assign n17504 = n2157 & n16259 ;
  assign n17505 = \s15_data_i[9]_pad  & n2157 ;
  assign n17506 = ~n2258 & n17505 ;
  assign n17507 = ~n17504 & ~n17506 ;
  assign n17508 = \s8_data_i[9]_pad  & n14841 ;
  assign n17509 = \s1_data_i[9]_pad  & n14658 ;
  assign n17510 = ~n17508 & ~n17509 ;
  assign n17511 = \s0_data_i[9]_pad  & n14582 ;
  assign n17512 = \s10_data_i[9]_pad  & n14797 ;
  assign n17513 = ~n17511 & ~n17512 ;
  assign n17514 = n17510 & n17513 ;
  assign n17515 = \s3_data_i[9]_pad  & n14820 ;
  assign n17516 = \s4_data_i[9]_pad  & n14825 ;
  assign n17517 = ~n17515 & ~n17516 ;
  assign n17518 = \s9_data_i[9]_pad  & n14845 ;
  assign n17519 = \s6_data_i[9]_pad  & n14833 ;
  assign n17520 = ~n17518 & ~n17519 ;
  assign n17521 = n17517 & n17520 ;
  assign n17522 = n17514 & n17521 ;
  assign n17523 = \s11_data_i[9]_pad  & n15106 ;
  assign n17524 = \s14_data_i[9]_pad  & n14809 ;
  assign n17525 = \s7_data_i[9]_pad  & n14837 ;
  assign n17526 = ~n17524 & ~n17525 ;
  assign n17527 = ~n17523 & n17526 ;
  assign n17528 = \s5_data_i[9]_pad  & n14829 ;
  assign n17529 = \s12_data_i[9]_pad  & n15102 ;
  assign n17530 = ~n17528 & ~n17529 ;
  assign n17531 = \s2_data_i[9]_pad  & n14816 ;
  assign n17532 = \s13_data_i[9]_pad  & n14805 ;
  assign n17533 = ~n17531 & ~n17532 ;
  assign n17534 = n17530 & n17533 ;
  assign n17535 = n17527 & n17534 ;
  assign n17536 = n17522 & n17535 ;
  assign n17537 = n17507 & n17536 ;
  assign n17538 = \s15_err_i_pad  & n16419 ;
  assign n17539 = ~n2258 & n17538 ;
  assign n17540 = \s14_err_i_pad  & n14809 ;
  assign n17541 = ~n14331 & n17540 ;
  assign n17542 = n14324 & n17541 ;
  assign n17543 = \s8_err_i_pad  & n14841 ;
  assign n17544 = ~n13767 & n17543 ;
  assign n17545 = n13760 & n17544 ;
  assign n17546 = ~n17542 & ~n17545 ;
  assign n17547 = \s9_err_i_pad  & n14845 ;
  assign n17548 = ~n13847 & n17547 ;
  assign n17549 = n13855 & n17548 ;
  assign n17550 = \s0_err_i_pad  & n14582 ;
  assign n17551 = ~n14069 & n17550 ;
  assign n17552 = n14094 & n17551 ;
  assign n17553 = ~n17549 & ~n17552 ;
  assign n17554 = n17546 & n17553 ;
  assign n17555 = \s6_err_i_pad  & n14833 ;
  assign n17556 = ~n13627 & n17555 ;
  assign n17557 = n13620 & n17556 ;
  assign n17558 = \s10_err_i_pad  & n14797 ;
  assign n17559 = ~n13928 & n17558 ;
  assign n17560 = n13945 & n17559 ;
  assign n17561 = ~n17557 & ~n17560 ;
  assign n17562 = \s4_err_i_pad  & n14825 ;
  assign n17563 = ~n13467 & n17562 ;
  assign n17564 = n13475 & n17563 ;
  assign n17565 = \s13_err_i_pad  & n14805 ;
  assign n17566 = ~n14211 & n17565 ;
  assign n17567 = n14219 & n17566 ;
  assign n17568 = ~n17564 & ~n17567 ;
  assign n17569 = n17561 & n17568 ;
  assign n17570 = n17554 & n17569 ;
  assign n17571 = \s12_err_i_pad  & n15102 ;
  assign n17572 = ~n14140 & n17571 ;
  assign n17573 = n14165 & n17572 ;
  assign n17574 = \s5_err_i_pad  & n14829 ;
  assign n17575 = ~n13547 & n17574 ;
  assign n17576 = n13572 & n17575 ;
  assign n17577 = \s7_err_i_pad  & n14837 ;
  assign n17578 = ~n13697 & n17577 ;
  assign n17579 = n13705 & n17578 ;
  assign n17580 = ~n17576 & ~n17579 ;
  assign n17581 = ~n17573 & n17580 ;
  assign n17582 = \s1_err_i_pad  & n14658 ;
  assign n17583 = ~n14271 & n17582 ;
  assign n17584 = n14296 & n17583 ;
  assign n17585 = \s2_err_i_pad  & n14816 ;
  assign n17586 = ~n14391 & n17585 ;
  assign n17587 = n14399 & n17586 ;
  assign n17588 = ~n17584 & ~n17587 ;
  assign n17589 = \s11_err_i_pad  & n15106 ;
  assign n17590 = ~n14009 & n17589 ;
  assign n17591 = n14017 & n17590 ;
  assign n17592 = \s3_err_i_pad  & n14820 ;
  assign n17593 = ~n14451 & n17592 ;
  assign n17594 = n14476 & n17593 ;
  assign n17595 = ~n17591 & ~n17594 ;
  assign n17596 = n17588 & n17595 ;
  assign n17597 = n17581 & n17596 ;
  assign n17598 = n17570 & n17597 ;
  assign n17599 = ~n17539 & n17598 ;
  assign n17600 = \s15_rty_i_pad  & n16419 ;
  assign n17601 = ~n2258 & n17600 ;
  assign n17602 = \s5_rty_i_pad  & n14829 ;
  assign n17603 = ~n13547 & n17602 ;
  assign n17604 = n13572 & n17603 ;
  assign n17605 = \s12_rty_i_pad  & n15102 ;
  assign n17606 = ~n14140 & n17605 ;
  assign n17607 = n14165 & n17606 ;
  assign n17608 = ~n17604 & ~n17607 ;
  assign n17609 = \s6_rty_i_pad  & n14833 ;
  assign n17610 = ~n13627 & n17609 ;
  assign n17611 = n13620 & n17610 ;
  assign n17612 = \s9_rty_i_pad  & n14845 ;
  assign n17613 = ~n13847 & n17612 ;
  assign n17614 = n13855 & n17613 ;
  assign n17615 = ~n17611 & ~n17614 ;
  assign n17616 = n17608 & n17615 ;
  assign n17617 = \s0_rty_i_pad  & n14582 ;
  assign n17618 = ~n14069 & n17617 ;
  assign n17619 = n14094 & n17618 ;
  assign n17620 = \s7_rty_i_pad  & n14837 ;
  assign n17621 = ~n13697 & n17620 ;
  assign n17622 = n13705 & n17621 ;
  assign n17623 = ~n17619 & ~n17622 ;
  assign n17624 = \s10_rty_i_pad  & n14797 ;
  assign n17625 = ~n13928 & n17624 ;
  assign n17626 = n13945 & n17625 ;
  assign n17627 = \s13_rty_i_pad  & n14805 ;
  assign n17628 = ~n14211 & n17627 ;
  assign n17629 = n14219 & n17628 ;
  assign n17630 = ~n17626 & ~n17629 ;
  assign n17631 = n17623 & n17630 ;
  assign n17632 = n17616 & n17631 ;
  assign n17633 = \s3_rty_i_pad  & n14820 ;
  assign n17634 = ~n14451 & n17633 ;
  assign n17635 = n14476 & n17634 ;
  assign n17636 = \s2_rty_i_pad  & n14816 ;
  assign n17637 = ~n14391 & n17636 ;
  assign n17638 = n14399 & n17637 ;
  assign n17639 = \s4_rty_i_pad  & n14825 ;
  assign n17640 = ~n13467 & n17639 ;
  assign n17641 = n13475 & n17640 ;
  assign n17642 = ~n17638 & ~n17641 ;
  assign n17643 = ~n17635 & n17642 ;
  assign n17644 = \s8_rty_i_pad  & n14841 ;
  assign n17645 = ~n13767 & n17644 ;
  assign n17646 = n13760 & n17645 ;
  assign n17647 = \s11_rty_i_pad  & n15106 ;
  assign n17648 = ~n14009 & n17647 ;
  assign n17649 = n14017 & n17648 ;
  assign n17650 = ~n17646 & ~n17649 ;
  assign n17651 = \s14_rty_i_pad  & n14809 ;
  assign n17652 = ~n14331 & n17651 ;
  assign n17653 = n14324 & n17652 ;
  assign n17654 = \s1_rty_i_pad  & n14658 ;
  assign n17655 = ~n14271 & n17654 ;
  assign n17656 = n14296 & n17655 ;
  assign n17657 = ~n17653 & ~n17656 ;
  assign n17658 = n17650 & n17657 ;
  assign n17659 = n17643 & n17658 ;
  assign n17660 = n17632 & n17659 ;
  assign n17661 = ~n17601 & n17660 ;
  assign n17662 = ~n1925 & n2184 ;
  assign n17663 = n1931 & n17662 ;
  assign n17664 = ~n13416 & n17663 ;
  assign n17665 = ~n15125 & n17664 ;
  assign n17666 = \s11_ack_i_pad  & n14855 ;
  assign n17667 = n14009 & n17666 ;
  assign n17668 = n14034 & n17667 ;
  assign n17669 = \s3_ack_i_pad  & n14870 ;
  assign n17670 = n14451 & n17669 ;
  assign n17671 = n14459 & n17670 ;
  assign n17672 = ~n17668 & ~n17671 ;
  assign n17673 = \s1_ack_i_pad  & n14596 ;
  assign n17674 = n14271 & n17673 ;
  assign n17675 = n14279 & n17674 ;
  assign n17676 = \s7_ack_i_pad  & n15090 ;
  assign n17677 = n13697 & n17676 ;
  assign n17678 = n13714 & n17677 ;
  assign n17679 = ~n17675 & ~n17678 ;
  assign n17680 = n17672 & n17679 ;
  assign n17681 = \s10_ack_i_pad  & n14851 ;
  assign n17682 = n13928 & n17681 ;
  assign n17683 = n13921 & n17682 ;
  assign n17684 = \s2_ack_i_pad  & n14866 ;
  assign n17685 = n14391 & n17684 ;
  assign n17686 = n14416 & n17685 ;
  assign n17687 = ~n17683 & ~n17686 ;
  assign n17688 = \s13_ack_i_pad  & n15094 ;
  assign n17689 = n14211 & n17688 ;
  assign n17690 = n14228 & n17689 ;
  assign n17691 = \s6_ack_i_pad  & n14883 ;
  assign n17692 = n13627 & n17691 ;
  assign n17693 = n13635 & n17692 ;
  assign n17694 = ~n17690 & ~n17693 ;
  assign n17695 = n17687 & n17694 ;
  assign n17696 = n17680 & n17695 ;
  assign n17697 = \s8_ack_i_pad  & n15082 ;
  assign n17698 = n13767 & n17697 ;
  assign n17699 = n13775 & n17698 ;
  assign n17700 = \s14_ack_i_pad  & n15098 ;
  assign n17701 = n14331 & n17700 ;
  assign n17702 = n14339 & n17701 ;
  assign n17703 = \s9_ack_i_pad  & n14887 ;
  assign n17704 = n13847 & n17703 ;
  assign n17705 = n13840 & n17704 ;
  assign n17706 = ~n17702 & ~n17705 ;
  assign n17707 = ~n17699 & n17706 ;
  assign n17708 = \s4_ack_i_pad  & n14875 ;
  assign n17709 = n13467 & n17708 ;
  assign n17710 = n13484 & n17709 ;
  assign n17711 = \s0_ack_i_pad  & n14590 ;
  assign n17712 = n14069 & n17711 ;
  assign n17713 = n14086 & n17712 ;
  assign n17714 = ~n17710 & ~n17713 ;
  assign n17715 = \s5_ack_i_pad  & n14879 ;
  assign n17716 = n13547 & n17715 ;
  assign n17717 = n13540 & n17716 ;
  assign n17718 = \s12_ack_i_pad  & n14859 ;
  assign n17719 = n14140 & n17718 ;
  assign n17720 = n14133 & n17719 ;
  assign n17721 = ~n17717 & ~n17720 ;
  assign n17722 = n17714 & n17721 ;
  assign n17723 = n17707 & n17722 ;
  assign n17724 = n17696 & n17723 ;
  assign n17725 = ~n17665 & n17724 ;
  assign n17726 = n2184 & n15192 ;
  assign n17727 = \s15_data_i[0]_pad  & n2184 ;
  assign n17728 = ~n2258 & n17727 ;
  assign n17729 = ~n17726 & ~n17728 ;
  assign n17730 = \s2_data_i[0]_pad  & n14866 ;
  assign n17731 = \s13_data_i[0]_pad  & n15094 ;
  assign n17732 = ~n17730 & ~n17731 ;
  assign n17733 = \s7_data_i[0]_pad  & n15090 ;
  assign n17734 = \s3_data_i[0]_pad  & n14870 ;
  assign n17735 = ~n17733 & ~n17734 ;
  assign n17736 = n17732 & n17735 ;
  assign n17737 = \s11_data_i[0]_pad  & n14855 ;
  assign n17738 = \s5_data_i[0]_pad  & n14879 ;
  assign n17739 = ~n17737 & ~n17738 ;
  assign n17740 = \s14_data_i[0]_pad  & n15098 ;
  assign n17741 = \s8_data_i[0]_pad  & n15082 ;
  assign n17742 = ~n17740 & ~n17741 ;
  assign n17743 = n17739 & n17742 ;
  assign n17744 = n17736 & n17743 ;
  assign n17745 = \s1_data_i[0]_pad  & n14596 ;
  assign n17746 = \s4_data_i[0]_pad  & n14875 ;
  assign n17747 = \s12_data_i[0]_pad  & n14859 ;
  assign n17748 = ~n17746 & ~n17747 ;
  assign n17749 = ~n17745 & n17748 ;
  assign n17750 = \s9_data_i[0]_pad  & n14887 ;
  assign n17751 = \s10_data_i[0]_pad  & n14851 ;
  assign n17752 = ~n17750 & ~n17751 ;
  assign n17753 = \s0_data_i[0]_pad  & n14590 ;
  assign n17754 = \s6_data_i[0]_pad  & n14883 ;
  assign n17755 = ~n17753 & ~n17754 ;
  assign n17756 = n17752 & n17755 ;
  assign n17757 = n17749 & n17756 ;
  assign n17758 = n17744 & n17757 ;
  assign n17759 = n17729 & n17758 ;
  assign n17760 = n2184 & n15229 ;
  assign n17761 = \s15_data_i[10]_pad  & n2184 ;
  assign n17762 = ~n2258 & n17761 ;
  assign n17763 = ~n17760 & ~n17762 ;
  assign n17764 = \s8_data_i[10]_pad  & n15082 ;
  assign n17765 = \s13_data_i[10]_pad  & n15094 ;
  assign n17766 = ~n17764 & ~n17765 ;
  assign n17767 = \s10_data_i[10]_pad  & n14851 ;
  assign n17768 = \s1_data_i[10]_pad  & n14596 ;
  assign n17769 = ~n17767 & ~n17768 ;
  assign n17770 = n17766 & n17769 ;
  assign n17771 = \s5_data_i[10]_pad  & n14879 ;
  assign n17772 = \s6_data_i[10]_pad  & n14883 ;
  assign n17773 = ~n17771 & ~n17772 ;
  assign n17774 = \s7_data_i[10]_pad  & n15090 ;
  assign n17775 = \s2_data_i[10]_pad  & n14866 ;
  assign n17776 = ~n17774 & ~n17775 ;
  assign n17777 = n17773 & n17776 ;
  assign n17778 = n17770 & n17777 ;
  assign n17779 = \s11_data_i[10]_pad  & n14855 ;
  assign n17780 = \s4_data_i[10]_pad  & n14875 ;
  assign n17781 = \s3_data_i[10]_pad  & n14870 ;
  assign n17782 = ~n17780 & ~n17781 ;
  assign n17783 = ~n17779 & n17782 ;
  assign n17784 = \s12_data_i[10]_pad  & n14859 ;
  assign n17785 = \s14_data_i[10]_pad  & n15098 ;
  assign n17786 = ~n17784 & ~n17785 ;
  assign n17787 = \s0_data_i[10]_pad  & n14590 ;
  assign n17788 = \s9_data_i[10]_pad  & n14887 ;
  assign n17789 = ~n17787 & ~n17788 ;
  assign n17790 = n17786 & n17789 ;
  assign n17791 = n17783 & n17790 ;
  assign n17792 = n17778 & n17791 ;
  assign n17793 = n17763 & n17792 ;
  assign n17794 = n2184 & n15266 ;
  assign n17795 = \s15_data_i[11]_pad  & n2184 ;
  assign n17796 = ~n2258 & n17795 ;
  assign n17797 = ~n17794 & ~n17796 ;
  assign n17798 = \s8_data_i[11]_pad  & n15082 ;
  assign n17799 = \s13_data_i[11]_pad  & n15094 ;
  assign n17800 = ~n17798 & ~n17799 ;
  assign n17801 = \s10_data_i[11]_pad  & n14851 ;
  assign n17802 = \s1_data_i[11]_pad  & n14596 ;
  assign n17803 = ~n17801 & ~n17802 ;
  assign n17804 = n17800 & n17803 ;
  assign n17805 = \s5_data_i[11]_pad  & n14879 ;
  assign n17806 = \s6_data_i[11]_pad  & n14883 ;
  assign n17807 = ~n17805 & ~n17806 ;
  assign n17808 = \s7_data_i[11]_pad  & n15090 ;
  assign n17809 = \s2_data_i[11]_pad  & n14866 ;
  assign n17810 = ~n17808 & ~n17809 ;
  assign n17811 = n17807 & n17810 ;
  assign n17812 = n17804 & n17811 ;
  assign n17813 = \s11_data_i[11]_pad  & n14855 ;
  assign n17814 = \s4_data_i[11]_pad  & n14875 ;
  assign n17815 = \s3_data_i[11]_pad  & n14870 ;
  assign n17816 = ~n17814 & ~n17815 ;
  assign n17817 = ~n17813 & n17816 ;
  assign n17818 = \s12_data_i[11]_pad  & n14859 ;
  assign n17819 = \s14_data_i[11]_pad  & n15098 ;
  assign n17820 = ~n17818 & ~n17819 ;
  assign n17821 = \s0_data_i[11]_pad  & n14590 ;
  assign n17822 = \s9_data_i[11]_pad  & n14887 ;
  assign n17823 = ~n17821 & ~n17822 ;
  assign n17824 = n17820 & n17823 ;
  assign n17825 = n17817 & n17824 ;
  assign n17826 = n17812 & n17825 ;
  assign n17827 = n17797 & n17826 ;
  assign n17828 = n2184 & n15303 ;
  assign n17829 = \s15_data_i[12]_pad  & n2184 ;
  assign n17830 = ~n2258 & n17829 ;
  assign n17831 = ~n17828 & ~n17830 ;
  assign n17832 = \s8_data_i[12]_pad  & n15082 ;
  assign n17833 = \s13_data_i[12]_pad  & n15094 ;
  assign n17834 = ~n17832 & ~n17833 ;
  assign n17835 = \s10_data_i[12]_pad  & n14851 ;
  assign n17836 = \s1_data_i[12]_pad  & n14596 ;
  assign n17837 = ~n17835 & ~n17836 ;
  assign n17838 = n17834 & n17837 ;
  assign n17839 = \s5_data_i[12]_pad  & n14879 ;
  assign n17840 = \s6_data_i[12]_pad  & n14883 ;
  assign n17841 = ~n17839 & ~n17840 ;
  assign n17842 = \s7_data_i[12]_pad  & n15090 ;
  assign n17843 = \s2_data_i[12]_pad  & n14866 ;
  assign n17844 = ~n17842 & ~n17843 ;
  assign n17845 = n17841 & n17844 ;
  assign n17846 = n17838 & n17845 ;
  assign n17847 = \s11_data_i[12]_pad  & n14855 ;
  assign n17848 = \s4_data_i[12]_pad  & n14875 ;
  assign n17849 = \s3_data_i[12]_pad  & n14870 ;
  assign n17850 = ~n17848 & ~n17849 ;
  assign n17851 = ~n17847 & n17850 ;
  assign n17852 = \s12_data_i[12]_pad  & n14859 ;
  assign n17853 = \s14_data_i[12]_pad  & n15098 ;
  assign n17854 = ~n17852 & ~n17853 ;
  assign n17855 = \s0_data_i[12]_pad  & n14590 ;
  assign n17856 = \s9_data_i[12]_pad  & n14887 ;
  assign n17857 = ~n17855 & ~n17856 ;
  assign n17858 = n17854 & n17857 ;
  assign n17859 = n17851 & n17858 ;
  assign n17860 = n17846 & n17859 ;
  assign n17861 = n17831 & n17860 ;
  assign n17862 = n2184 & n15340 ;
  assign n17863 = \s15_data_i[13]_pad  & n2184 ;
  assign n17864 = ~n2258 & n17863 ;
  assign n17865 = ~n17862 & ~n17864 ;
  assign n17866 = \s8_data_i[13]_pad  & n15082 ;
  assign n17867 = \s1_data_i[13]_pad  & n14596 ;
  assign n17868 = ~n17866 & ~n17867 ;
  assign n17869 = \s4_data_i[13]_pad  & n14875 ;
  assign n17870 = \s6_data_i[13]_pad  & n14883 ;
  assign n17871 = ~n17869 & ~n17870 ;
  assign n17872 = n17868 & n17871 ;
  assign n17873 = \s5_data_i[13]_pad  & n14879 ;
  assign n17874 = \s9_data_i[13]_pad  & n14887 ;
  assign n17875 = ~n17873 & ~n17874 ;
  assign n17876 = \s10_data_i[13]_pad  & n14851 ;
  assign n17877 = \s7_data_i[13]_pad  & n15090 ;
  assign n17878 = ~n17876 & ~n17877 ;
  assign n17879 = n17875 & n17878 ;
  assign n17880 = n17872 & n17879 ;
  assign n17881 = \s11_data_i[13]_pad  & n14855 ;
  assign n17882 = \s13_data_i[13]_pad  & n15094 ;
  assign n17883 = \s3_data_i[13]_pad  & n14870 ;
  assign n17884 = ~n17882 & ~n17883 ;
  assign n17885 = ~n17881 & n17884 ;
  assign n17886 = \s12_data_i[13]_pad  & n14859 ;
  assign n17887 = \s14_data_i[13]_pad  & n15098 ;
  assign n17888 = ~n17886 & ~n17887 ;
  assign n17889 = \s2_data_i[13]_pad  & n14866 ;
  assign n17890 = \s0_data_i[13]_pad  & n14590 ;
  assign n17891 = ~n17889 & ~n17890 ;
  assign n17892 = n17888 & n17891 ;
  assign n17893 = n17885 & n17892 ;
  assign n17894 = n17880 & n17893 ;
  assign n17895 = n17865 & n17894 ;
  assign n17896 = n2184 & n15377 ;
  assign n17897 = \s15_data_i[14]_pad  & n2184 ;
  assign n17898 = ~n2258 & n17897 ;
  assign n17899 = ~n17896 & ~n17898 ;
  assign n17900 = \s12_data_i[14]_pad  & n14859 ;
  assign n17901 = \s13_data_i[14]_pad  & n15094 ;
  assign n17902 = ~n17900 & ~n17901 ;
  assign n17903 = \s10_data_i[14]_pad  & n14851 ;
  assign n17904 = \s1_data_i[14]_pad  & n14596 ;
  assign n17905 = ~n17903 & ~n17904 ;
  assign n17906 = n17902 & n17905 ;
  assign n17907 = \s5_data_i[14]_pad  & n14879 ;
  assign n17908 = \s0_data_i[14]_pad  & n14590 ;
  assign n17909 = ~n17907 & ~n17908 ;
  assign n17910 = \s4_data_i[14]_pad  & n14875 ;
  assign n17911 = \s2_data_i[14]_pad  & n14866 ;
  assign n17912 = ~n17910 & ~n17911 ;
  assign n17913 = n17909 & n17912 ;
  assign n17914 = n17906 & n17913 ;
  assign n17915 = \s14_data_i[14]_pad  & n15098 ;
  assign n17916 = \s7_data_i[14]_pad  & n15090 ;
  assign n17917 = \s3_data_i[14]_pad  & n14870 ;
  assign n17918 = ~n17916 & ~n17917 ;
  assign n17919 = ~n17915 & n17918 ;
  assign n17920 = \s8_data_i[14]_pad  & n15082 ;
  assign n17921 = \s11_data_i[14]_pad  & n14855 ;
  assign n17922 = ~n17920 & ~n17921 ;
  assign n17923 = \s6_data_i[14]_pad  & n14883 ;
  assign n17924 = \s9_data_i[14]_pad  & n14887 ;
  assign n17925 = ~n17923 & ~n17924 ;
  assign n17926 = n17922 & n17925 ;
  assign n17927 = n17919 & n17926 ;
  assign n17928 = n17914 & n17927 ;
  assign n17929 = n17899 & n17928 ;
  assign n17930 = n2184 & n15414 ;
  assign n17931 = \s15_data_i[15]_pad  & n2184 ;
  assign n17932 = ~n2258 & n17931 ;
  assign n17933 = ~n17930 & ~n17932 ;
  assign n17934 = \s12_data_i[15]_pad  & n14859 ;
  assign n17935 = \s13_data_i[15]_pad  & n15094 ;
  assign n17936 = ~n17934 & ~n17935 ;
  assign n17937 = \s10_data_i[15]_pad  & n14851 ;
  assign n17938 = \s3_data_i[15]_pad  & n14870 ;
  assign n17939 = ~n17937 & ~n17938 ;
  assign n17940 = n17936 & n17939 ;
  assign n17941 = \s2_data_i[15]_pad  & n14866 ;
  assign n17942 = \s0_data_i[15]_pad  & n14590 ;
  assign n17943 = ~n17941 & ~n17942 ;
  assign n17944 = \s4_data_i[15]_pad  & n14875 ;
  assign n17945 = \s5_data_i[15]_pad  & n14879 ;
  assign n17946 = ~n17944 & ~n17945 ;
  assign n17947 = n17943 & n17946 ;
  assign n17948 = n17940 & n17947 ;
  assign n17949 = \s14_data_i[15]_pad  & n15098 ;
  assign n17950 = \s7_data_i[15]_pad  & n15090 ;
  assign n17951 = \s1_data_i[15]_pad  & n14596 ;
  assign n17952 = ~n17950 & ~n17951 ;
  assign n17953 = ~n17949 & n17952 ;
  assign n17954 = \s8_data_i[15]_pad  & n15082 ;
  assign n17955 = \s11_data_i[15]_pad  & n14855 ;
  assign n17956 = ~n17954 & ~n17955 ;
  assign n17957 = \s6_data_i[15]_pad  & n14883 ;
  assign n17958 = \s9_data_i[15]_pad  & n14887 ;
  assign n17959 = ~n17957 & ~n17958 ;
  assign n17960 = n17956 & n17959 ;
  assign n17961 = n17953 & n17960 ;
  assign n17962 = n17948 & n17961 ;
  assign n17963 = n17933 & n17962 ;
  assign n17964 = \s15_data_i[16]_pad  & n2184 ;
  assign n17965 = ~n2258 & n17964 ;
  assign n17966 = \s12_data_i[16]_pad  & n14859 ;
  assign n17967 = \s13_data_i[16]_pad  & n15094 ;
  assign n17968 = ~n17966 & ~n17967 ;
  assign n17969 = \s10_data_i[16]_pad  & n14851 ;
  assign n17970 = \s3_data_i[16]_pad  & n14870 ;
  assign n17971 = ~n17969 & ~n17970 ;
  assign n17972 = n17968 & n17971 ;
  assign n17973 = \s2_data_i[16]_pad  & n14866 ;
  assign n17974 = \s6_data_i[16]_pad  & n14883 ;
  assign n17975 = ~n17973 & ~n17974 ;
  assign n17976 = \s7_data_i[16]_pad  & n15090 ;
  assign n17977 = \s5_data_i[16]_pad  & n14879 ;
  assign n17978 = ~n17976 & ~n17977 ;
  assign n17979 = n17975 & n17978 ;
  assign n17980 = n17972 & n17979 ;
  assign n17981 = \s14_data_i[16]_pad  & n15098 ;
  assign n17982 = \s4_data_i[16]_pad  & n14875 ;
  assign n17983 = \s1_data_i[16]_pad  & n14596 ;
  assign n17984 = ~n17982 & ~n17983 ;
  assign n17985 = ~n17981 & n17984 ;
  assign n17986 = \s8_data_i[16]_pad  & n15082 ;
  assign n17987 = \s11_data_i[16]_pad  & n14855 ;
  assign n17988 = ~n17986 & ~n17987 ;
  assign n17989 = \s0_data_i[16]_pad  & n14590 ;
  assign n17990 = \s9_data_i[16]_pad  & n14887 ;
  assign n17991 = ~n17989 & ~n17990 ;
  assign n17992 = n17988 & n17991 ;
  assign n17993 = n17985 & n17992 ;
  assign n17994 = n17980 & n17993 ;
  assign n17995 = ~n17965 & n17994 ;
  assign n17996 = \s15_data_i[17]_pad  & n2184 ;
  assign n17997 = ~n2258 & n17996 ;
  assign n17998 = \s12_data_i[17]_pad  & n14859 ;
  assign n17999 = \s13_data_i[17]_pad  & n15094 ;
  assign n18000 = ~n17998 & ~n17999 ;
  assign n18001 = \s10_data_i[17]_pad  & n14851 ;
  assign n18002 = \s1_data_i[17]_pad  & n14596 ;
  assign n18003 = ~n18001 & ~n18002 ;
  assign n18004 = n18000 & n18003 ;
  assign n18005 = \s5_data_i[17]_pad  & n14879 ;
  assign n18006 = \s6_data_i[17]_pad  & n14883 ;
  assign n18007 = ~n18005 & ~n18006 ;
  assign n18008 = \s7_data_i[17]_pad  & n15090 ;
  assign n18009 = \s2_data_i[17]_pad  & n14866 ;
  assign n18010 = ~n18008 & ~n18009 ;
  assign n18011 = n18007 & n18010 ;
  assign n18012 = n18004 & n18011 ;
  assign n18013 = \s14_data_i[17]_pad  & n15098 ;
  assign n18014 = \s4_data_i[17]_pad  & n14875 ;
  assign n18015 = \s3_data_i[17]_pad  & n14870 ;
  assign n18016 = ~n18014 & ~n18015 ;
  assign n18017 = ~n18013 & n18016 ;
  assign n18018 = \s8_data_i[17]_pad  & n15082 ;
  assign n18019 = \s11_data_i[17]_pad  & n14855 ;
  assign n18020 = ~n18018 & ~n18019 ;
  assign n18021 = \s0_data_i[17]_pad  & n14590 ;
  assign n18022 = \s9_data_i[17]_pad  & n14887 ;
  assign n18023 = ~n18021 & ~n18022 ;
  assign n18024 = n18020 & n18023 ;
  assign n18025 = n18017 & n18024 ;
  assign n18026 = n18012 & n18025 ;
  assign n18027 = ~n17997 & n18026 ;
  assign n18028 = \s15_data_i[18]_pad  & n2184 ;
  assign n18029 = ~n2258 & n18028 ;
  assign n18030 = \s12_data_i[18]_pad  & n14859 ;
  assign n18031 = \s13_data_i[18]_pad  & n15094 ;
  assign n18032 = ~n18030 & ~n18031 ;
  assign n18033 = \s10_data_i[18]_pad  & n14851 ;
  assign n18034 = \s1_data_i[18]_pad  & n14596 ;
  assign n18035 = ~n18033 & ~n18034 ;
  assign n18036 = n18032 & n18035 ;
  assign n18037 = \s5_data_i[18]_pad  & n14879 ;
  assign n18038 = \s6_data_i[18]_pad  & n14883 ;
  assign n18039 = ~n18037 & ~n18038 ;
  assign n18040 = \s7_data_i[18]_pad  & n15090 ;
  assign n18041 = \s2_data_i[18]_pad  & n14866 ;
  assign n18042 = ~n18040 & ~n18041 ;
  assign n18043 = n18039 & n18042 ;
  assign n18044 = n18036 & n18043 ;
  assign n18045 = \s14_data_i[18]_pad  & n15098 ;
  assign n18046 = \s4_data_i[18]_pad  & n14875 ;
  assign n18047 = \s3_data_i[18]_pad  & n14870 ;
  assign n18048 = ~n18046 & ~n18047 ;
  assign n18049 = ~n18045 & n18048 ;
  assign n18050 = \s8_data_i[18]_pad  & n15082 ;
  assign n18051 = \s11_data_i[18]_pad  & n14855 ;
  assign n18052 = ~n18050 & ~n18051 ;
  assign n18053 = \s0_data_i[18]_pad  & n14590 ;
  assign n18054 = \s9_data_i[18]_pad  & n14887 ;
  assign n18055 = ~n18053 & ~n18054 ;
  assign n18056 = n18052 & n18055 ;
  assign n18057 = n18049 & n18056 ;
  assign n18058 = n18044 & n18057 ;
  assign n18059 = ~n18029 & n18058 ;
  assign n18060 = \s15_data_i[19]_pad  & n2184 ;
  assign n18061 = ~n2258 & n18060 ;
  assign n18062 = \s12_data_i[19]_pad  & n14859 ;
  assign n18063 = \s13_data_i[19]_pad  & n15094 ;
  assign n18064 = ~n18062 & ~n18063 ;
  assign n18065 = \s10_data_i[19]_pad  & n14851 ;
  assign n18066 = \s1_data_i[19]_pad  & n14596 ;
  assign n18067 = ~n18065 & ~n18066 ;
  assign n18068 = n18064 & n18067 ;
  assign n18069 = \s5_data_i[19]_pad  & n14879 ;
  assign n18070 = \s6_data_i[19]_pad  & n14883 ;
  assign n18071 = ~n18069 & ~n18070 ;
  assign n18072 = \s7_data_i[19]_pad  & n15090 ;
  assign n18073 = \s2_data_i[19]_pad  & n14866 ;
  assign n18074 = ~n18072 & ~n18073 ;
  assign n18075 = n18071 & n18074 ;
  assign n18076 = n18068 & n18075 ;
  assign n18077 = \s14_data_i[19]_pad  & n15098 ;
  assign n18078 = \s4_data_i[19]_pad  & n14875 ;
  assign n18079 = \s3_data_i[19]_pad  & n14870 ;
  assign n18080 = ~n18078 & ~n18079 ;
  assign n18081 = ~n18077 & n18080 ;
  assign n18082 = \s8_data_i[19]_pad  & n15082 ;
  assign n18083 = \s11_data_i[19]_pad  & n14855 ;
  assign n18084 = ~n18082 & ~n18083 ;
  assign n18085 = \s0_data_i[19]_pad  & n14590 ;
  assign n18086 = \s9_data_i[19]_pad  & n14887 ;
  assign n18087 = ~n18085 & ~n18086 ;
  assign n18088 = n18084 & n18087 ;
  assign n18089 = n18081 & n18088 ;
  assign n18090 = n18076 & n18089 ;
  assign n18091 = ~n18061 & n18090 ;
  assign n18092 = n2184 & n15579 ;
  assign n18093 = \s15_data_i[1]_pad  & n2184 ;
  assign n18094 = ~n2258 & n18093 ;
  assign n18095 = ~n18092 & ~n18094 ;
  assign n18096 = \s8_data_i[1]_pad  & n15082 ;
  assign n18097 = \s10_data_i[1]_pad  & n14851 ;
  assign n18098 = ~n18096 & ~n18097 ;
  assign n18099 = \s4_data_i[1]_pad  & n14875 ;
  assign n18100 = \s1_data_i[1]_pad  & n14596 ;
  assign n18101 = ~n18099 & ~n18100 ;
  assign n18102 = n18098 & n18101 ;
  assign n18103 = \s5_data_i[1]_pad  & n14879 ;
  assign n18104 = \s0_data_i[1]_pad  & n14590 ;
  assign n18105 = ~n18103 & ~n18104 ;
  assign n18106 = \s13_data_i[1]_pad  & n15094 ;
  assign n18107 = \s2_data_i[1]_pad  & n14866 ;
  assign n18108 = ~n18106 & ~n18107 ;
  assign n18109 = n18105 & n18108 ;
  assign n18110 = n18102 & n18109 ;
  assign n18111 = \s11_data_i[1]_pad  & n14855 ;
  assign n18112 = \s7_data_i[1]_pad  & n15090 ;
  assign n18113 = \s3_data_i[1]_pad  & n14870 ;
  assign n18114 = ~n18112 & ~n18113 ;
  assign n18115 = ~n18111 & n18114 ;
  assign n18116 = \s12_data_i[1]_pad  & n14859 ;
  assign n18117 = \s14_data_i[1]_pad  & n15098 ;
  assign n18118 = ~n18116 & ~n18117 ;
  assign n18119 = \s9_data_i[1]_pad  & n14887 ;
  assign n18120 = \s6_data_i[1]_pad  & n14883 ;
  assign n18121 = ~n18119 & ~n18120 ;
  assign n18122 = n18118 & n18121 ;
  assign n18123 = n18115 & n18122 ;
  assign n18124 = n18110 & n18123 ;
  assign n18125 = n18095 & n18124 ;
  assign n18126 = \s15_data_i[20]_pad  & n2184 ;
  assign n18127 = ~n2258 & n18126 ;
  assign n18128 = \s12_data_i[20]_pad  & n14859 ;
  assign n18129 = \s13_data_i[20]_pad  & n15094 ;
  assign n18130 = ~n18128 & ~n18129 ;
  assign n18131 = \s10_data_i[20]_pad  & n14851 ;
  assign n18132 = \s1_data_i[20]_pad  & n14596 ;
  assign n18133 = ~n18131 & ~n18132 ;
  assign n18134 = n18130 & n18133 ;
  assign n18135 = \s5_data_i[20]_pad  & n14879 ;
  assign n18136 = \s6_data_i[20]_pad  & n14883 ;
  assign n18137 = ~n18135 & ~n18136 ;
  assign n18138 = \s7_data_i[20]_pad  & n15090 ;
  assign n18139 = \s2_data_i[20]_pad  & n14866 ;
  assign n18140 = ~n18138 & ~n18139 ;
  assign n18141 = n18137 & n18140 ;
  assign n18142 = n18134 & n18141 ;
  assign n18143 = \s14_data_i[20]_pad  & n15098 ;
  assign n18144 = \s4_data_i[20]_pad  & n14875 ;
  assign n18145 = \s3_data_i[20]_pad  & n14870 ;
  assign n18146 = ~n18144 & ~n18145 ;
  assign n18147 = ~n18143 & n18146 ;
  assign n18148 = \s8_data_i[20]_pad  & n15082 ;
  assign n18149 = \s11_data_i[20]_pad  & n14855 ;
  assign n18150 = ~n18148 & ~n18149 ;
  assign n18151 = \s0_data_i[20]_pad  & n14590 ;
  assign n18152 = \s9_data_i[20]_pad  & n14887 ;
  assign n18153 = ~n18151 & ~n18152 ;
  assign n18154 = n18150 & n18153 ;
  assign n18155 = n18147 & n18154 ;
  assign n18156 = n18142 & n18155 ;
  assign n18157 = ~n18127 & n18156 ;
  assign n18158 = \s15_data_i[21]_pad  & n2184 ;
  assign n18159 = ~n2258 & n18158 ;
  assign n18160 = \s12_data_i[21]_pad  & n14859 ;
  assign n18161 = \s13_data_i[21]_pad  & n15094 ;
  assign n18162 = ~n18160 & ~n18161 ;
  assign n18163 = \s10_data_i[21]_pad  & n14851 ;
  assign n18164 = \s1_data_i[21]_pad  & n14596 ;
  assign n18165 = ~n18163 & ~n18164 ;
  assign n18166 = n18162 & n18165 ;
  assign n18167 = \s5_data_i[21]_pad  & n14879 ;
  assign n18168 = \s6_data_i[21]_pad  & n14883 ;
  assign n18169 = ~n18167 & ~n18168 ;
  assign n18170 = \s7_data_i[21]_pad  & n15090 ;
  assign n18171 = \s2_data_i[21]_pad  & n14866 ;
  assign n18172 = ~n18170 & ~n18171 ;
  assign n18173 = n18169 & n18172 ;
  assign n18174 = n18166 & n18173 ;
  assign n18175 = \s14_data_i[21]_pad  & n15098 ;
  assign n18176 = \s4_data_i[21]_pad  & n14875 ;
  assign n18177 = \s3_data_i[21]_pad  & n14870 ;
  assign n18178 = ~n18176 & ~n18177 ;
  assign n18179 = ~n18175 & n18178 ;
  assign n18180 = \s8_data_i[21]_pad  & n15082 ;
  assign n18181 = \s11_data_i[21]_pad  & n14855 ;
  assign n18182 = ~n18180 & ~n18181 ;
  assign n18183 = \s0_data_i[21]_pad  & n14590 ;
  assign n18184 = \s9_data_i[21]_pad  & n14887 ;
  assign n18185 = ~n18183 & ~n18184 ;
  assign n18186 = n18182 & n18185 ;
  assign n18187 = n18179 & n18186 ;
  assign n18188 = n18174 & n18187 ;
  assign n18189 = ~n18159 & n18188 ;
  assign n18190 = \s15_data_i[22]_pad  & n2184 ;
  assign n18191 = ~n2258 & n18190 ;
  assign n18192 = \s12_data_i[22]_pad  & n14859 ;
  assign n18193 = \s13_data_i[22]_pad  & n15094 ;
  assign n18194 = ~n18192 & ~n18193 ;
  assign n18195 = \s10_data_i[22]_pad  & n14851 ;
  assign n18196 = \s1_data_i[22]_pad  & n14596 ;
  assign n18197 = ~n18195 & ~n18196 ;
  assign n18198 = n18194 & n18197 ;
  assign n18199 = \s5_data_i[22]_pad  & n14879 ;
  assign n18200 = \s6_data_i[22]_pad  & n14883 ;
  assign n18201 = ~n18199 & ~n18200 ;
  assign n18202 = \s7_data_i[22]_pad  & n15090 ;
  assign n18203 = \s2_data_i[22]_pad  & n14866 ;
  assign n18204 = ~n18202 & ~n18203 ;
  assign n18205 = n18201 & n18204 ;
  assign n18206 = n18198 & n18205 ;
  assign n18207 = \s14_data_i[22]_pad  & n15098 ;
  assign n18208 = \s4_data_i[22]_pad  & n14875 ;
  assign n18209 = \s3_data_i[22]_pad  & n14870 ;
  assign n18210 = ~n18208 & ~n18209 ;
  assign n18211 = ~n18207 & n18210 ;
  assign n18212 = \s8_data_i[22]_pad  & n15082 ;
  assign n18213 = \s11_data_i[22]_pad  & n14855 ;
  assign n18214 = ~n18212 & ~n18213 ;
  assign n18215 = \s0_data_i[22]_pad  & n14590 ;
  assign n18216 = \s9_data_i[22]_pad  & n14887 ;
  assign n18217 = ~n18215 & ~n18216 ;
  assign n18218 = n18214 & n18217 ;
  assign n18219 = n18211 & n18218 ;
  assign n18220 = n18206 & n18219 ;
  assign n18221 = ~n18191 & n18220 ;
  assign n18222 = \s15_data_i[23]_pad  & n2184 ;
  assign n18223 = ~n2258 & n18222 ;
  assign n18224 = \s12_data_i[23]_pad  & n14859 ;
  assign n18225 = \s13_data_i[23]_pad  & n15094 ;
  assign n18226 = ~n18224 & ~n18225 ;
  assign n18227 = \s10_data_i[23]_pad  & n14851 ;
  assign n18228 = \s1_data_i[23]_pad  & n14596 ;
  assign n18229 = ~n18227 & ~n18228 ;
  assign n18230 = n18226 & n18229 ;
  assign n18231 = \s5_data_i[23]_pad  & n14879 ;
  assign n18232 = \s6_data_i[23]_pad  & n14883 ;
  assign n18233 = ~n18231 & ~n18232 ;
  assign n18234 = \s7_data_i[23]_pad  & n15090 ;
  assign n18235 = \s2_data_i[23]_pad  & n14866 ;
  assign n18236 = ~n18234 & ~n18235 ;
  assign n18237 = n18233 & n18236 ;
  assign n18238 = n18230 & n18237 ;
  assign n18239 = \s14_data_i[23]_pad  & n15098 ;
  assign n18240 = \s4_data_i[23]_pad  & n14875 ;
  assign n18241 = \s3_data_i[23]_pad  & n14870 ;
  assign n18242 = ~n18240 & ~n18241 ;
  assign n18243 = ~n18239 & n18242 ;
  assign n18244 = \s8_data_i[23]_pad  & n15082 ;
  assign n18245 = \s11_data_i[23]_pad  & n14855 ;
  assign n18246 = ~n18244 & ~n18245 ;
  assign n18247 = \s0_data_i[23]_pad  & n14590 ;
  assign n18248 = \s9_data_i[23]_pad  & n14887 ;
  assign n18249 = ~n18247 & ~n18248 ;
  assign n18250 = n18246 & n18249 ;
  assign n18251 = n18243 & n18250 ;
  assign n18252 = n18238 & n18251 ;
  assign n18253 = ~n18223 & n18252 ;
  assign n18254 = \s15_data_i[24]_pad  & n2184 ;
  assign n18255 = ~n2258 & n18254 ;
  assign n18256 = \s12_data_i[24]_pad  & n14859 ;
  assign n18257 = \s13_data_i[24]_pad  & n15094 ;
  assign n18258 = ~n18256 & ~n18257 ;
  assign n18259 = \s10_data_i[24]_pad  & n14851 ;
  assign n18260 = \s1_data_i[24]_pad  & n14596 ;
  assign n18261 = ~n18259 & ~n18260 ;
  assign n18262 = n18258 & n18261 ;
  assign n18263 = \s5_data_i[24]_pad  & n14879 ;
  assign n18264 = \s6_data_i[24]_pad  & n14883 ;
  assign n18265 = ~n18263 & ~n18264 ;
  assign n18266 = \s7_data_i[24]_pad  & n15090 ;
  assign n18267 = \s2_data_i[24]_pad  & n14866 ;
  assign n18268 = ~n18266 & ~n18267 ;
  assign n18269 = n18265 & n18268 ;
  assign n18270 = n18262 & n18269 ;
  assign n18271 = \s14_data_i[24]_pad  & n15098 ;
  assign n18272 = \s4_data_i[24]_pad  & n14875 ;
  assign n18273 = \s3_data_i[24]_pad  & n14870 ;
  assign n18274 = ~n18272 & ~n18273 ;
  assign n18275 = ~n18271 & n18274 ;
  assign n18276 = \s8_data_i[24]_pad  & n15082 ;
  assign n18277 = \s11_data_i[24]_pad  & n14855 ;
  assign n18278 = ~n18276 & ~n18277 ;
  assign n18279 = \s0_data_i[24]_pad  & n14590 ;
  assign n18280 = \s9_data_i[24]_pad  & n14887 ;
  assign n18281 = ~n18279 & ~n18280 ;
  assign n18282 = n18278 & n18281 ;
  assign n18283 = n18275 & n18282 ;
  assign n18284 = n18270 & n18283 ;
  assign n18285 = ~n18255 & n18284 ;
  assign n18286 = \s15_data_i[25]_pad  & n2184 ;
  assign n18287 = ~n2258 & n18286 ;
  assign n18288 = \s12_data_i[25]_pad  & n14859 ;
  assign n18289 = \s13_data_i[25]_pad  & n15094 ;
  assign n18290 = ~n18288 & ~n18289 ;
  assign n18291 = \s10_data_i[25]_pad  & n14851 ;
  assign n18292 = \s1_data_i[25]_pad  & n14596 ;
  assign n18293 = ~n18291 & ~n18292 ;
  assign n18294 = n18290 & n18293 ;
  assign n18295 = \s5_data_i[25]_pad  & n14879 ;
  assign n18296 = \s6_data_i[25]_pad  & n14883 ;
  assign n18297 = ~n18295 & ~n18296 ;
  assign n18298 = \s7_data_i[25]_pad  & n15090 ;
  assign n18299 = \s2_data_i[25]_pad  & n14866 ;
  assign n18300 = ~n18298 & ~n18299 ;
  assign n18301 = n18297 & n18300 ;
  assign n18302 = n18294 & n18301 ;
  assign n18303 = \s14_data_i[25]_pad  & n15098 ;
  assign n18304 = \s4_data_i[25]_pad  & n14875 ;
  assign n18305 = \s3_data_i[25]_pad  & n14870 ;
  assign n18306 = ~n18304 & ~n18305 ;
  assign n18307 = ~n18303 & n18306 ;
  assign n18308 = \s8_data_i[25]_pad  & n15082 ;
  assign n18309 = \s11_data_i[25]_pad  & n14855 ;
  assign n18310 = ~n18308 & ~n18309 ;
  assign n18311 = \s0_data_i[25]_pad  & n14590 ;
  assign n18312 = \s9_data_i[25]_pad  & n14887 ;
  assign n18313 = ~n18311 & ~n18312 ;
  assign n18314 = n18310 & n18313 ;
  assign n18315 = n18307 & n18314 ;
  assign n18316 = n18302 & n18315 ;
  assign n18317 = ~n18287 & n18316 ;
  assign n18318 = \s15_data_i[26]_pad  & n2184 ;
  assign n18319 = ~n2258 & n18318 ;
  assign n18320 = \s12_data_i[26]_pad  & n14859 ;
  assign n18321 = \s13_data_i[26]_pad  & n15094 ;
  assign n18322 = ~n18320 & ~n18321 ;
  assign n18323 = \s10_data_i[26]_pad  & n14851 ;
  assign n18324 = \s1_data_i[26]_pad  & n14596 ;
  assign n18325 = ~n18323 & ~n18324 ;
  assign n18326 = n18322 & n18325 ;
  assign n18327 = \s5_data_i[26]_pad  & n14879 ;
  assign n18328 = \s6_data_i[26]_pad  & n14883 ;
  assign n18329 = ~n18327 & ~n18328 ;
  assign n18330 = \s7_data_i[26]_pad  & n15090 ;
  assign n18331 = \s2_data_i[26]_pad  & n14866 ;
  assign n18332 = ~n18330 & ~n18331 ;
  assign n18333 = n18329 & n18332 ;
  assign n18334 = n18326 & n18333 ;
  assign n18335 = \s14_data_i[26]_pad  & n15098 ;
  assign n18336 = \s4_data_i[26]_pad  & n14875 ;
  assign n18337 = \s3_data_i[26]_pad  & n14870 ;
  assign n18338 = ~n18336 & ~n18337 ;
  assign n18339 = ~n18335 & n18338 ;
  assign n18340 = \s8_data_i[26]_pad  & n15082 ;
  assign n18341 = \s11_data_i[26]_pad  & n14855 ;
  assign n18342 = ~n18340 & ~n18341 ;
  assign n18343 = \s0_data_i[26]_pad  & n14590 ;
  assign n18344 = \s9_data_i[26]_pad  & n14887 ;
  assign n18345 = ~n18343 & ~n18344 ;
  assign n18346 = n18342 & n18345 ;
  assign n18347 = n18339 & n18346 ;
  assign n18348 = n18334 & n18347 ;
  assign n18349 = ~n18319 & n18348 ;
  assign n18350 = \s15_data_i[27]_pad  & n2184 ;
  assign n18351 = ~n2258 & n18350 ;
  assign n18352 = \s12_data_i[27]_pad  & n14859 ;
  assign n18353 = \s13_data_i[27]_pad  & n15094 ;
  assign n18354 = ~n18352 & ~n18353 ;
  assign n18355 = \s10_data_i[27]_pad  & n14851 ;
  assign n18356 = \s1_data_i[27]_pad  & n14596 ;
  assign n18357 = ~n18355 & ~n18356 ;
  assign n18358 = n18354 & n18357 ;
  assign n18359 = \s5_data_i[27]_pad  & n14879 ;
  assign n18360 = \s6_data_i[27]_pad  & n14883 ;
  assign n18361 = ~n18359 & ~n18360 ;
  assign n18362 = \s7_data_i[27]_pad  & n15090 ;
  assign n18363 = \s2_data_i[27]_pad  & n14866 ;
  assign n18364 = ~n18362 & ~n18363 ;
  assign n18365 = n18361 & n18364 ;
  assign n18366 = n18358 & n18365 ;
  assign n18367 = \s14_data_i[27]_pad  & n15098 ;
  assign n18368 = \s4_data_i[27]_pad  & n14875 ;
  assign n18369 = \s3_data_i[27]_pad  & n14870 ;
  assign n18370 = ~n18368 & ~n18369 ;
  assign n18371 = ~n18367 & n18370 ;
  assign n18372 = \s8_data_i[27]_pad  & n15082 ;
  assign n18373 = \s11_data_i[27]_pad  & n14855 ;
  assign n18374 = ~n18372 & ~n18373 ;
  assign n18375 = \s0_data_i[27]_pad  & n14590 ;
  assign n18376 = \s9_data_i[27]_pad  & n14887 ;
  assign n18377 = ~n18375 & ~n18376 ;
  assign n18378 = n18374 & n18377 ;
  assign n18379 = n18371 & n18378 ;
  assign n18380 = n18366 & n18379 ;
  assign n18381 = ~n18351 & n18380 ;
  assign n18382 = \s15_data_i[28]_pad  & n2184 ;
  assign n18383 = ~n2258 & n18382 ;
  assign n18384 = \s12_data_i[28]_pad  & n14859 ;
  assign n18385 = \s13_data_i[28]_pad  & n15094 ;
  assign n18386 = ~n18384 & ~n18385 ;
  assign n18387 = \s10_data_i[28]_pad  & n14851 ;
  assign n18388 = \s1_data_i[28]_pad  & n14596 ;
  assign n18389 = ~n18387 & ~n18388 ;
  assign n18390 = n18386 & n18389 ;
  assign n18391 = \s5_data_i[28]_pad  & n14879 ;
  assign n18392 = \s6_data_i[28]_pad  & n14883 ;
  assign n18393 = ~n18391 & ~n18392 ;
  assign n18394 = \s7_data_i[28]_pad  & n15090 ;
  assign n18395 = \s2_data_i[28]_pad  & n14866 ;
  assign n18396 = ~n18394 & ~n18395 ;
  assign n18397 = n18393 & n18396 ;
  assign n18398 = n18390 & n18397 ;
  assign n18399 = \s14_data_i[28]_pad  & n15098 ;
  assign n18400 = \s4_data_i[28]_pad  & n14875 ;
  assign n18401 = \s3_data_i[28]_pad  & n14870 ;
  assign n18402 = ~n18400 & ~n18401 ;
  assign n18403 = ~n18399 & n18402 ;
  assign n18404 = \s8_data_i[28]_pad  & n15082 ;
  assign n18405 = \s11_data_i[28]_pad  & n14855 ;
  assign n18406 = ~n18404 & ~n18405 ;
  assign n18407 = \s0_data_i[28]_pad  & n14590 ;
  assign n18408 = \s9_data_i[28]_pad  & n14887 ;
  assign n18409 = ~n18407 & ~n18408 ;
  assign n18410 = n18406 & n18409 ;
  assign n18411 = n18403 & n18410 ;
  assign n18412 = n18398 & n18411 ;
  assign n18413 = ~n18383 & n18412 ;
  assign n18414 = \s15_data_i[29]_pad  & n2184 ;
  assign n18415 = ~n2258 & n18414 ;
  assign n18416 = \s12_data_i[29]_pad  & n14859 ;
  assign n18417 = \s13_data_i[29]_pad  & n15094 ;
  assign n18418 = ~n18416 & ~n18417 ;
  assign n18419 = \s10_data_i[29]_pad  & n14851 ;
  assign n18420 = \s1_data_i[29]_pad  & n14596 ;
  assign n18421 = ~n18419 & ~n18420 ;
  assign n18422 = n18418 & n18421 ;
  assign n18423 = \s5_data_i[29]_pad  & n14879 ;
  assign n18424 = \s6_data_i[29]_pad  & n14883 ;
  assign n18425 = ~n18423 & ~n18424 ;
  assign n18426 = \s7_data_i[29]_pad  & n15090 ;
  assign n18427 = \s2_data_i[29]_pad  & n14866 ;
  assign n18428 = ~n18426 & ~n18427 ;
  assign n18429 = n18425 & n18428 ;
  assign n18430 = n18422 & n18429 ;
  assign n18431 = \s14_data_i[29]_pad  & n15098 ;
  assign n18432 = \s4_data_i[29]_pad  & n14875 ;
  assign n18433 = \s3_data_i[29]_pad  & n14870 ;
  assign n18434 = ~n18432 & ~n18433 ;
  assign n18435 = ~n18431 & n18434 ;
  assign n18436 = \s8_data_i[29]_pad  & n15082 ;
  assign n18437 = \s11_data_i[29]_pad  & n14855 ;
  assign n18438 = ~n18436 & ~n18437 ;
  assign n18439 = \s0_data_i[29]_pad  & n14590 ;
  assign n18440 = \s9_data_i[29]_pad  & n14887 ;
  assign n18441 = ~n18439 & ~n18440 ;
  assign n18442 = n18438 & n18441 ;
  assign n18443 = n18435 & n18442 ;
  assign n18444 = n18430 & n18443 ;
  assign n18445 = ~n18415 & n18444 ;
  assign n18446 = n2184 & n15936 ;
  assign n18447 = \s15_data_i[2]_pad  & n2184 ;
  assign n18448 = ~n2258 & n18447 ;
  assign n18449 = ~n18446 & ~n18448 ;
  assign n18450 = \s8_data_i[2]_pad  & n15082 ;
  assign n18451 = \s1_data_i[2]_pad  & n14596 ;
  assign n18452 = ~n18450 & ~n18451 ;
  assign n18453 = \s4_data_i[2]_pad  & n14875 ;
  assign n18454 = \s6_data_i[2]_pad  & n14883 ;
  assign n18455 = ~n18453 & ~n18454 ;
  assign n18456 = n18452 & n18455 ;
  assign n18457 = \s5_data_i[2]_pad  & n14879 ;
  assign n18458 = \s9_data_i[2]_pad  & n14887 ;
  assign n18459 = ~n18457 & ~n18458 ;
  assign n18460 = \s10_data_i[2]_pad  & n14851 ;
  assign n18461 = \s7_data_i[2]_pad  & n15090 ;
  assign n18462 = ~n18460 & ~n18461 ;
  assign n18463 = n18459 & n18462 ;
  assign n18464 = n18456 & n18463 ;
  assign n18465 = \s11_data_i[2]_pad  & n14855 ;
  assign n18466 = \s13_data_i[2]_pad  & n15094 ;
  assign n18467 = \s3_data_i[2]_pad  & n14870 ;
  assign n18468 = ~n18466 & ~n18467 ;
  assign n18469 = ~n18465 & n18468 ;
  assign n18470 = \s12_data_i[2]_pad  & n14859 ;
  assign n18471 = \s14_data_i[2]_pad  & n15098 ;
  assign n18472 = ~n18470 & ~n18471 ;
  assign n18473 = \s2_data_i[2]_pad  & n14866 ;
  assign n18474 = \s0_data_i[2]_pad  & n14590 ;
  assign n18475 = ~n18473 & ~n18474 ;
  assign n18476 = n18472 & n18475 ;
  assign n18477 = n18469 & n18476 ;
  assign n18478 = n18464 & n18477 ;
  assign n18479 = n18449 & n18478 ;
  assign n18480 = \s15_data_i[30]_pad  & n2184 ;
  assign n18481 = ~n2258 & n18480 ;
  assign n18482 = \s12_data_i[30]_pad  & n14859 ;
  assign n18483 = \s13_data_i[30]_pad  & n15094 ;
  assign n18484 = ~n18482 & ~n18483 ;
  assign n18485 = \s10_data_i[30]_pad  & n14851 ;
  assign n18486 = \s1_data_i[30]_pad  & n14596 ;
  assign n18487 = ~n18485 & ~n18486 ;
  assign n18488 = n18484 & n18487 ;
  assign n18489 = \s5_data_i[30]_pad  & n14879 ;
  assign n18490 = \s6_data_i[30]_pad  & n14883 ;
  assign n18491 = ~n18489 & ~n18490 ;
  assign n18492 = \s7_data_i[30]_pad  & n15090 ;
  assign n18493 = \s2_data_i[30]_pad  & n14866 ;
  assign n18494 = ~n18492 & ~n18493 ;
  assign n18495 = n18491 & n18494 ;
  assign n18496 = n18488 & n18495 ;
  assign n18497 = \s14_data_i[30]_pad  & n15098 ;
  assign n18498 = \s4_data_i[30]_pad  & n14875 ;
  assign n18499 = \s3_data_i[30]_pad  & n14870 ;
  assign n18500 = ~n18498 & ~n18499 ;
  assign n18501 = ~n18497 & n18500 ;
  assign n18502 = \s8_data_i[30]_pad  & n15082 ;
  assign n18503 = \s11_data_i[30]_pad  & n14855 ;
  assign n18504 = ~n18502 & ~n18503 ;
  assign n18505 = \s0_data_i[30]_pad  & n14590 ;
  assign n18506 = \s9_data_i[30]_pad  & n14887 ;
  assign n18507 = ~n18505 & ~n18506 ;
  assign n18508 = n18504 & n18507 ;
  assign n18509 = n18501 & n18508 ;
  assign n18510 = n18496 & n18509 ;
  assign n18511 = ~n18481 & n18510 ;
  assign n18512 = \s15_data_i[31]_pad  & n2184 ;
  assign n18513 = ~n2258 & n18512 ;
  assign n18514 = \s12_data_i[31]_pad  & n14859 ;
  assign n18515 = \s13_data_i[31]_pad  & n15094 ;
  assign n18516 = ~n18514 & ~n18515 ;
  assign n18517 = \s10_data_i[31]_pad  & n14851 ;
  assign n18518 = \s1_data_i[31]_pad  & n14596 ;
  assign n18519 = ~n18517 & ~n18518 ;
  assign n18520 = n18516 & n18519 ;
  assign n18521 = \s5_data_i[31]_pad  & n14879 ;
  assign n18522 = \s6_data_i[31]_pad  & n14883 ;
  assign n18523 = ~n18521 & ~n18522 ;
  assign n18524 = \s7_data_i[31]_pad  & n15090 ;
  assign n18525 = \s2_data_i[31]_pad  & n14866 ;
  assign n18526 = ~n18524 & ~n18525 ;
  assign n18527 = n18523 & n18526 ;
  assign n18528 = n18520 & n18527 ;
  assign n18529 = \s14_data_i[31]_pad  & n15098 ;
  assign n18530 = \s4_data_i[31]_pad  & n14875 ;
  assign n18531 = \s3_data_i[31]_pad  & n14870 ;
  assign n18532 = ~n18530 & ~n18531 ;
  assign n18533 = ~n18529 & n18532 ;
  assign n18534 = \s8_data_i[31]_pad  & n15082 ;
  assign n18535 = \s11_data_i[31]_pad  & n14855 ;
  assign n18536 = ~n18534 & ~n18535 ;
  assign n18537 = \s0_data_i[31]_pad  & n14590 ;
  assign n18538 = \s9_data_i[31]_pad  & n14887 ;
  assign n18539 = ~n18537 & ~n18538 ;
  assign n18540 = n18536 & n18539 ;
  assign n18541 = n18533 & n18540 ;
  assign n18542 = n18528 & n18541 ;
  assign n18543 = ~n18513 & n18542 ;
  assign n18544 = n2184 & n16037 ;
  assign n18545 = \s15_data_i[3]_pad  & n2184 ;
  assign n18546 = ~n2258 & n18545 ;
  assign n18547 = ~n18544 & ~n18546 ;
  assign n18548 = \s8_data_i[3]_pad  & n15082 ;
  assign n18549 = \s13_data_i[3]_pad  & n15094 ;
  assign n18550 = ~n18548 & ~n18549 ;
  assign n18551 = \s10_data_i[3]_pad  & n14851 ;
  assign n18552 = \s1_data_i[3]_pad  & n14596 ;
  assign n18553 = ~n18551 & ~n18552 ;
  assign n18554 = n18550 & n18553 ;
  assign n18555 = \s5_data_i[3]_pad  & n14879 ;
  assign n18556 = \s6_data_i[3]_pad  & n14883 ;
  assign n18557 = ~n18555 & ~n18556 ;
  assign n18558 = \s7_data_i[3]_pad  & n15090 ;
  assign n18559 = \s2_data_i[3]_pad  & n14866 ;
  assign n18560 = ~n18558 & ~n18559 ;
  assign n18561 = n18557 & n18560 ;
  assign n18562 = n18554 & n18561 ;
  assign n18563 = \s11_data_i[3]_pad  & n14855 ;
  assign n18564 = \s4_data_i[3]_pad  & n14875 ;
  assign n18565 = \s3_data_i[3]_pad  & n14870 ;
  assign n18566 = ~n18564 & ~n18565 ;
  assign n18567 = ~n18563 & n18566 ;
  assign n18568 = \s12_data_i[3]_pad  & n14859 ;
  assign n18569 = \s14_data_i[3]_pad  & n15098 ;
  assign n18570 = ~n18568 & ~n18569 ;
  assign n18571 = \s0_data_i[3]_pad  & n14590 ;
  assign n18572 = \s9_data_i[3]_pad  & n14887 ;
  assign n18573 = ~n18571 & ~n18572 ;
  assign n18574 = n18570 & n18573 ;
  assign n18575 = n18567 & n18574 ;
  assign n18576 = n18562 & n18575 ;
  assign n18577 = n18547 & n18576 ;
  assign n18578 = n2184 & n16074 ;
  assign n18579 = \s15_data_i[4]_pad  & n2184 ;
  assign n18580 = ~n2258 & n18579 ;
  assign n18581 = ~n18578 & ~n18580 ;
  assign n18582 = \s2_data_i[4]_pad  & n14866 ;
  assign n18583 = \s13_data_i[4]_pad  & n15094 ;
  assign n18584 = ~n18582 & ~n18583 ;
  assign n18585 = \s7_data_i[4]_pad  & n15090 ;
  assign n18586 = \s3_data_i[4]_pad  & n14870 ;
  assign n18587 = ~n18585 & ~n18586 ;
  assign n18588 = n18584 & n18587 ;
  assign n18589 = \s11_data_i[4]_pad  & n14855 ;
  assign n18590 = \s5_data_i[4]_pad  & n14879 ;
  assign n18591 = ~n18589 & ~n18590 ;
  assign n18592 = \s14_data_i[4]_pad  & n15098 ;
  assign n18593 = \s8_data_i[4]_pad  & n15082 ;
  assign n18594 = ~n18592 & ~n18593 ;
  assign n18595 = n18591 & n18594 ;
  assign n18596 = n18588 & n18595 ;
  assign n18597 = \s1_data_i[4]_pad  & n14596 ;
  assign n18598 = \s4_data_i[4]_pad  & n14875 ;
  assign n18599 = \s12_data_i[4]_pad  & n14859 ;
  assign n18600 = ~n18598 & ~n18599 ;
  assign n18601 = ~n18597 & n18600 ;
  assign n18602 = \s9_data_i[4]_pad  & n14887 ;
  assign n18603 = \s10_data_i[4]_pad  & n14851 ;
  assign n18604 = ~n18602 & ~n18603 ;
  assign n18605 = \s0_data_i[4]_pad  & n14590 ;
  assign n18606 = \s6_data_i[4]_pad  & n14883 ;
  assign n18607 = ~n18605 & ~n18606 ;
  assign n18608 = n18604 & n18607 ;
  assign n18609 = n18601 & n18608 ;
  assign n18610 = n18596 & n18609 ;
  assign n18611 = n18581 & n18610 ;
  assign n18612 = n2184 & n16111 ;
  assign n18613 = \s15_data_i[5]_pad  & n2184 ;
  assign n18614 = ~n2258 & n18613 ;
  assign n18615 = ~n18612 & ~n18614 ;
  assign n18616 = \s8_data_i[5]_pad  & n15082 ;
  assign n18617 = \s13_data_i[5]_pad  & n15094 ;
  assign n18618 = ~n18616 & ~n18617 ;
  assign n18619 = \s10_data_i[5]_pad  & n14851 ;
  assign n18620 = \s1_data_i[5]_pad  & n14596 ;
  assign n18621 = ~n18619 & ~n18620 ;
  assign n18622 = n18618 & n18621 ;
  assign n18623 = \s5_data_i[5]_pad  & n14879 ;
  assign n18624 = \s6_data_i[5]_pad  & n14883 ;
  assign n18625 = ~n18623 & ~n18624 ;
  assign n18626 = \s7_data_i[5]_pad  & n15090 ;
  assign n18627 = \s2_data_i[5]_pad  & n14866 ;
  assign n18628 = ~n18626 & ~n18627 ;
  assign n18629 = n18625 & n18628 ;
  assign n18630 = n18622 & n18629 ;
  assign n18631 = \s11_data_i[5]_pad  & n14855 ;
  assign n18632 = \s4_data_i[5]_pad  & n14875 ;
  assign n18633 = \s3_data_i[5]_pad  & n14870 ;
  assign n18634 = ~n18632 & ~n18633 ;
  assign n18635 = ~n18631 & n18634 ;
  assign n18636 = \s12_data_i[5]_pad  & n14859 ;
  assign n18637 = \s14_data_i[5]_pad  & n15098 ;
  assign n18638 = ~n18636 & ~n18637 ;
  assign n18639 = \s0_data_i[5]_pad  & n14590 ;
  assign n18640 = \s9_data_i[5]_pad  & n14887 ;
  assign n18641 = ~n18639 & ~n18640 ;
  assign n18642 = n18638 & n18641 ;
  assign n18643 = n18635 & n18642 ;
  assign n18644 = n18630 & n18643 ;
  assign n18645 = n18615 & n18644 ;
  assign n18646 = n2184 & n16148 ;
  assign n18647 = \s15_data_i[6]_pad  & n2184 ;
  assign n18648 = ~n2258 & n18647 ;
  assign n18649 = ~n18646 & ~n18648 ;
  assign n18650 = \s8_data_i[6]_pad  & n15082 ;
  assign n18651 = \s13_data_i[6]_pad  & n15094 ;
  assign n18652 = ~n18650 & ~n18651 ;
  assign n18653 = \s10_data_i[6]_pad  & n14851 ;
  assign n18654 = \s1_data_i[6]_pad  & n14596 ;
  assign n18655 = ~n18653 & ~n18654 ;
  assign n18656 = n18652 & n18655 ;
  assign n18657 = \s5_data_i[6]_pad  & n14879 ;
  assign n18658 = \s6_data_i[6]_pad  & n14883 ;
  assign n18659 = ~n18657 & ~n18658 ;
  assign n18660 = \s7_data_i[6]_pad  & n15090 ;
  assign n18661 = \s2_data_i[6]_pad  & n14866 ;
  assign n18662 = ~n18660 & ~n18661 ;
  assign n18663 = n18659 & n18662 ;
  assign n18664 = n18656 & n18663 ;
  assign n18665 = \s11_data_i[6]_pad  & n14855 ;
  assign n18666 = \s4_data_i[6]_pad  & n14875 ;
  assign n18667 = \s3_data_i[6]_pad  & n14870 ;
  assign n18668 = ~n18666 & ~n18667 ;
  assign n18669 = ~n18665 & n18668 ;
  assign n18670 = \s12_data_i[6]_pad  & n14859 ;
  assign n18671 = \s14_data_i[6]_pad  & n15098 ;
  assign n18672 = ~n18670 & ~n18671 ;
  assign n18673 = \s0_data_i[6]_pad  & n14590 ;
  assign n18674 = \s9_data_i[6]_pad  & n14887 ;
  assign n18675 = ~n18673 & ~n18674 ;
  assign n18676 = n18672 & n18675 ;
  assign n18677 = n18669 & n18676 ;
  assign n18678 = n18664 & n18677 ;
  assign n18679 = n18649 & n18678 ;
  assign n18680 = n2184 & n16185 ;
  assign n18681 = \s15_data_i[7]_pad  & n2184 ;
  assign n18682 = ~n2258 & n18681 ;
  assign n18683 = ~n18680 & ~n18682 ;
  assign n18684 = \s2_data_i[7]_pad  & n14866 ;
  assign n18685 = \s13_data_i[7]_pad  & n15094 ;
  assign n18686 = ~n18684 & ~n18685 ;
  assign n18687 = \s7_data_i[7]_pad  & n15090 ;
  assign n18688 = \s3_data_i[7]_pad  & n14870 ;
  assign n18689 = ~n18687 & ~n18688 ;
  assign n18690 = n18686 & n18689 ;
  assign n18691 = \s11_data_i[7]_pad  & n14855 ;
  assign n18692 = \s5_data_i[7]_pad  & n14879 ;
  assign n18693 = ~n18691 & ~n18692 ;
  assign n18694 = \s14_data_i[7]_pad  & n15098 ;
  assign n18695 = \s8_data_i[7]_pad  & n15082 ;
  assign n18696 = ~n18694 & ~n18695 ;
  assign n18697 = n18693 & n18696 ;
  assign n18698 = n18690 & n18697 ;
  assign n18699 = \s1_data_i[7]_pad  & n14596 ;
  assign n18700 = \s4_data_i[7]_pad  & n14875 ;
  assign n18701 = \s12_data_i[7]_pad  & n14859 ;
  assign n18702 = ~n18700 & ~n18701 ;
  assign n18703 = ~n18699 & n18702 ;
  assign n18704 = \s9_data_i[7]_pad  & n14887 ;
  assign n18705 = \s10_data_i[7]_pad  & n14851 ;
  assign n18706 = ~n18704 & ~n18705 ;
  assign n18707 = \s0_data_i[7]_pad  & n14590 ;
  assign n18708 = \s6_data_i[7]_pad  & n14883 ;
  assign n18709 = ~n18707 & ~n18708 ;
  assign n18710 = n18706 & n18709 ;
  assign n18711 = n18703 & n18710 ;
  assign n18712 = n18698 & n18711 ;
  assign n18713 = n18683 & n18712 ;
  assign n18714 = n2184 & n16222 ;
  assign n18715 = \s15_data_i[8]_pad  & n2184 ;
  assign n18716 = ~n2258 & n18715 ;
  assign n18717 = ~n18714 & ~n18716 ;
  assign n18718 = \s8_data_i[8]_pad  & n15082 ;
  assign n18719 = \s13_data_i[8]_pad  & n15094 ;
  assign n18720 = ~n18718 & ~n18719 ;
  assign n18721 = \s10_data_i[8]_pad  & n14851 ;
  assign n18722 = \s1_data_i[8]_pad  & n14596 ;
  assign n18723 = ~n18721 & ~n18722 ;
  assign n18724 = n18720 & n18723 ;
  assign n18725 = \s5_data_i[8]_pad  & n14879 ;
  assign n18726 = \s6_data_i[8]_pad  & n14883 ;
  assign n18727 = ~n18725 & ~n18726 ;
  assign n18728 = \s7_data_i[8]_pad  & n15090 ;
  assign n18729 = \s2_data_i[8]_pad  & n14866 ;
  assign n18730 = ~n18728 & ~n18729 ;
  assign n18731 = n18727 & n18730 ;
  assign n18732 = n18724 & n18731 ;
  assign n18733 = \s11_data_i[8]_pad  & n14855 ;
  assign n18734 = \s4_data_i[8]_pad  & n14875 ;
  assign n18735 = \s3_data_i[8]_pad  & n14870 ;
  assign n18736 = ~n18734 & ~n18735 ;
  assign n18737 = ~n18733 & n18736 ;
  assign n18738 = \s12_data_i[8]_pad  & n14859 ;
  assign n18739 = \s14_data_i[8]_pad  & n15098 ;
  assign n18740 = ~n18738 & ~n18739 ;
  assign n18741 = \s0_data_i[8]_pad  & n14590 ;
  assign n18742 = \s9_data_i[8]_pad  & n14887 ;
  assign n18743 = ~n18741 & ~n18742 ;
  assign n18744 = n18740 & n18743 ;
  assign n18745 = n18737 & n18744 ;
  assign n18746 = n18732 & n18745 ;
  assign n18747 = n18717 & n18746 ;
  assign n18748 = n2184 & n16259 ;
  assign n18749 = \s15_data_i[9]_pad  & n2184 ;
  assign n18750 = ~n2258 & n18749 ;
  assign n18751 = ~n18748 & ~n18750 ;
  assign n18752 = \s2_data_i[9]_pad  & n14866 ;
  assign n18753 = \s13_data_i[9]_pad  & n15094 ;
  assign n18754 = ~n18752 & ~n18753 ;
  assign n18755 = \s7_data_i[9]_pad  & n15090 ;
  assign n18756 = \s3_data_i[9]_pad  & n14870 ;
  assign n18757 = ~n18755 & ~n18756 ;
  assign n18758 = n18754 & n18757 ;
  assign n18759 = \s11_data_i[9]_pad  & n14855 ;
  assign n18760 = \s5_data_i[9]_pad  & n14879 ;
  assign n18761 = ~n18759 & ~n18760 ;
  assign n18762 = \s14_data_i[9]_pad  & n15098 ;
  assign n18763 = \s8_data_i[9]_pad  & n15082 ;
  assign n18764 = ~n18762 & ~n18763 ;
  assign n18765 = n18761 & n18764 ;
  assign n18766 = n18758 & n18765 ;
  assign n18767 = \s1_data_i[9]_pad  & n14596 ;
  assign n18768 = \s4_data_i[9]_pad  & n14875 ;
  assign n18769 = \s12_data_i[9]_pad  & n14859 ;
  assign n18770 = ~n18768 & ~n18769 ;
  assign n18771 = ~n18767 & n18770 ;
  assign n18772 = \s9_data_i[9]_pad  & n14887 ;
  assign n18773 = \s10_data_i[9]_pad  & n14851 ;
  assign n18774 = ~n18772 & ~n18773 ;
  assign n18775 = \s0_data_i[9]_pad  & n14590 ;
  assign n18776 = \s6_data_i[9]_pad  & n14883 ;
  assign n18777 = ~n18775 & ~n18776 ;
  assign n18778 = n18774 & n18777 ;
  assign n18779 = n18771 & n18778 ;
  assign n18780 = n18766 & n18779 ;
  assign n18781 = n18751 & n18780 ;
  assign n18782 = \s15_err_i_pad  & n17663 ;
  assign n18783 = ~n2258 & n18782 ;
  assign n18784 = \s11_err_i_pad  & n14855 ;
  assign n18785 = n14009 & n18784 ;
  assign n18786 = n14034 & n18785 ;
  assign n18787 = \s3_err_i_pad  & n14870 ;
  assign n18788 = n14451 & n18787 ;
  assign n18789 = n14459 & n18788 ;
  assign n18790 = ~n18786 & ~n18789 ;
  assign n18791 = \s9_err_i_pad  & n14887 ;
  assign n18792 = n13847 & n18791 ;
  assign n18793 = n13840 & n18792 ;
  assign n18794 = \s0_err_i_pad  & n14590 ;
  assign n18795 = n14069 & n18794 ;
  assign n18796 = n14086 & n18795 ;
  assign n18797 = ~n18793 & ~n18796 ;
  assign n18798 = n18790 & n18797 ;
  assign n18799 = \s6_err_i_pad  & n14883 ;
  assign n18800 = n13627 & n18799 ;
  assign n18801 = n13635 & n18800 ;
  assign n18802 = \s10_err_i_pad  & n14851 ;
  assign n18803 = n13928 & n18802 ;
  assign n18804 = n13921 & n18803 ;
  assign n18805 = ~n18801 & ~n18804 ;
  assign n18806 = \s4_err_i_pad  & n14875 ;
  assign n18807 = n13467 & n18806 ;
  assign n18808 = n13484 & n18807 ;
  assign n18809 = \s13_err_i_pad  & n15094 ;
  assign n18810 = n14211 & n18809 ;
  assign n18811 = n14228 & n18810 ;
  assign n18812 = ~n18808 & ~n18811 ;
  assign n18813 = n18805 & n18812 ;
  assign n18814 = n18798 & n18813 ;
  assign n18815 = \s8_err_i_pad  & n15082 ;
  assign n18816 = n13767 & n18815 ;
  assign n18817 = n13775 & n18816 ;
  assign n18818 = \s2_err_i_pad  & n14866 ;
  assign n18819 = n14391 & n18818 ;
  assign n18820 = n14416 & n18819 ;
  assign n18821 = \s7_err_i_pad  & n15090 ;
  assign n18822 = n13697 & n18821 ;
  assign n18823 = n13714 & n18822 ;
  assign n18824 = ~n18820 & ~n18823 ;
  assign n18825 = ~n18817 & n18824 ;
  assign n18826 = \s12_err_i_pad  & n14859 ;
  assign n18827 = n14140 & n18826 ;
  assign n18828 = n14133 & n18827 ;
  assign n18829 = \s14_err_i_pad  & n15098 ;
  assign n18830 = n14331 & n18829 ;
  assign n18831 = n14339 & n18830 ;
  assign n18832 = ~n18828 & ~n18831 ;
  assign n18833 = \s5_err_i_pad  & n14879 ;
  assign n18834 = n13547 & n18833 ;
  assign n18835 = n13540 & n18834 ;
  assign n18836 = \s1_err_i_pad  & n14596 ;
  assign n18837 = n14271 & n18836 ;
  assign n18838 = n14279 & n18837 ;
  assign n18839 = ~n18835 & ~n18838 ;
  assign n18840 = n18832 & n18839 ;
  assign n18841 = n18825 & n18840 ;
  assign n18842 = n18814 & n18841 ;
  assign n18843 = ~n18783 & n18842 ;
  assign n18844 = \s15_rty_i_pad  & n17663 ;
  assign n18845 = ~n2258 & n18844 ;
  assign n18846 = \s11_rty_i_pad  & n14855 ;
  assign n18847 = n14009 & n18846 ;
  assign n18848 = n14034 & n18847 ;
  assign n18849 = \s3_rty_i_pad  & n14870 ;
  assign n18850 = n14451 & n18849 ;
  assign n18851 = n14459 & n18850 ;
  assign n18852 = ~n18848 & ~n18851 ;
  assign n18853 = \s6_rty_i_pad  & n14883 ;
  assign n18854 = n13627 & n18853 ;
  assign n18855 = n13635 & n18854 ;
  assign n18856 = \s0_rty_i_pad  & n14590 ;
  assign n18857 = n14069 & n18856 ;
  assign n18858 = n14086 & n18857 ;
  assign n18859 = ~n18855 & ~n18858 ;
  assign n18860 = n18852 & n18859 ;
  assign n18861 = \s9_rty_i_pad  & n14887 ;
  assign n18862 = n13847 & n18861 ;
  assign n18863 = n13840 & n18862 ;
  assign n18864 = \s7_rty_i_pad  & n15090 ;
  assign n18865 = n13697 & n18864 ;
  assign n18866 = n13714 & n18865 ;
  assign n18867 = ~n18863 & ~n18866 ;
  assign n18868 = \s4_rty_i_pad  & n14875 ;
  assign n18869 = n13467 & n18868 ;
  assign n18870 = n13484 & n18869 ;
  assign n18871 = \s13_rty_i_pad  & n15094 ;
  assign n18872 = n14211 & n18871 ;
  assign n18873 = n14228 & n18872 ;
  assign n18874 = ~n18870 & ~n18873 ;
  assign n18875 = n18867 & n18874 ;
  assign n18876 = n18860 & n18875 ;
  assign n18877 = \s8_rty_i_pad  & n15082 ;
  assign n18878 = n13767 & n18877 ;
  assign n18879 = n13775 & n18878 ;
  assign n18880 = \s2_rty_i_pad  & n14866 ;
  assign n18881 = n14391 & n18880 ;
  assign n18882 = n14416 & n18881 ;
  assign n18883 = \s10_rty_i_pad  & n14851 ;
  assign n18884 = n13928 & n18883 ;
  assign n18885 = n13921 & n18884 ;
  assign n18886 = ~n18882 & ~n18885 ;
  assign n18887 = ~n18879 & n18886 ;
  assign n18888 = \s12_rty_i_pad  & n14859 ;
  assign n18889 = n14140 & n18888 ;
  assign n18890 = n14133 & n18889 ;
  assign n18891 = \s14_rty_i_pad  & n15098 ;
  assign n18892 = n14331 & n18891 ;
  assign n18893 = n14339 & n18892 ;
  assign n18894 = ~n18890 & ~n18893 ;
  assign n18895 = \s5_rty_i_pad  & n14879 ;
  assign n18896 = n13547 & n18895 ;
  assign n18897 = n13540 & n18896 ;
  assign n18898 = \s1_rty_i_pad  & n14596 ;
  assign n18899 = n14271 & n18898 ;
  assign n18900 = n14279 & n18899 ;
  assign n18901 = ~n18897 & ~n18900 ;
  assign n18902 = n18894 & n18901 ;
  assign n18903 = n18887 & n18902 ;
  assign n18904 = n18876 & n18903 ;
  assign n18905 = ~n18845 & n18904 ;
  assign n18906 = n1910 & n2190 ;
  assign n18907 = n1938 & n18906 ;
  assign n18908 = ~n13416 & n18907 ;
  assign n18909 = ~n15125 & n18908 ;
  assign n18910 = \s5_ack_i_pad  & n14757 ;
  assign n18911 = ~n13547 & n18910 ;
  assign n18912 = n13540 & n18911 ;
  assign n18913 = \s1_ack_i_pad  & n14609 ;
  assign n18914 = ~n14271 & n18913 ;
  assign n18915 = n14279 & n18914 ;
  assign n18916 = ~n18912 & ~n18915 ;
  assign n18917 = \s8_ack_i_pad  & n14923 ;
  assign n18918 = ~n13767 & n18917 ;
  assign n18919 = n13775 & n18918 ;
  assign n18920 = \s10_ack_i_pad  & n14892 ;
  assign n18921 = ~n13928 & n18920 ;
  assign n18922 = n13921 & n18921 ;
  assign n18923 = ~n18919 & ~n18922 ;
  assign n18924 = n18916 & n18923 ;
  assign n18925 = \s7_ack_i_pad  & n14740 ;
  assign n18926 = ~n13697 & n18925 ;
  assign n18927 = n13714 & n18926 ;
  assign n18928 = \s11_ack_i_pad  & n14896 ;
  assign n18929 = ~n14009 & n18928 ;
  assign n18930 = n14034 & n18929 ;
  assign n18931 = ~n18927 & ~n18930 ;
  assign n18932 = \s13_ack_i_pad  & n14904 ;
  assign n18933 = ~n14211 & n18932 ;
  assign n18934 = n14228 & n18933 ;
  assign n18935 = \s9_ack_i_pad  & n14927 ;
  assign n18936 = ~n13847 & n18935 ;
  assign n18937 = n13840 & n18936 ;
  assign n18938 = ~n18934 & ~n18937 ;
  assign n18939 = n18931 & n18938 ;
  assign n18940 = n18924 & n18939 ;
  assign n18941 = \s3_ack_i_pad  & n14801 ;
  assign n18942 = ~n14451 & n18941 ;
  assign n18943 = n14459 & n18942 ;
  assign n18944 = \s14_ack_i_pad  & n14915 ;
  assign n18945 = ~n14331 & n18944 ;
  assign n18946 = n14339 & n18945 ;
  assign n18947 = \s6_ack_i_pad  & n14745 ;
  assign n18948 = ~n13627 & n18947 ;
  assign n18949 = n13635 & n18948 ;
  assign n18950 = ~n18946 & ~n18949 ;
  assign n18951 = ~n18943 & n18950 ;
  assign n18952 = \s4_ack_i_pad  & n14919 ;
  assign n18953 = ~n13467 & n18952 ;
  assign n18954 = n13484 & n18953 ;
  assign n18955 = \s0_ack_i_pad  & n14603 ;
  assign n18956 = ~n14069 & n18955 ;
  assign n18957 = n14086 & n18956 ;
  assign n18958 = ~n18954 & ~n18957 ;
  assign n18959 = \s2_ack_i_pad  & n14911 ;
  assign n18960 = ~n14391 & n18959 ;
  assign n18961 = n14416 & n18960 ;
  assign n18962 = \s12_ack_i_pad  & n14900 ;
  assign n18963 = ~n14140 & n18962 ;
  assign n18964 = n14133 & n18963 ;
  assign n18965 = ~n18961 & ~n18964 ;
  assign n18966 = n18958 & n18965 ;
  assign n18967 = n18951 & n18966 ;
  assign n18968 = n18940 & n18967 ;
  assign n18969 = ~n18909 & n18968 ;
  assign n18970 = n2190 & n15192 ;
  assign n18971 = \s15_data_i[0]_pad  & n2190 ;
  assign n18972 = ~n2258 & n18971 ;
  assign n18973 = ~n18970 & ~n18972 ;
  assign n18974 = \s8_data_i[0]_pad  & n14923 ;
  assign n18975 = \s1_data_i[0]_pad  & n14609 ;
  assign n18976 = ~n18974 & ~n18975 ;
  assign n18977 = \s4_data_i[0]_pad  & n14919 ;
  assign n18978 = \s6_data_i[0]_pad  & n14745 ;
  assign n18979 = ~n18977 & ~n18978 ;
  assign n18980 = n18976 & n18979 ;
  assign n18981 = \s5_data_i[0]_pad  & n14757 ;
  assign n18982 = \s9_data_i[0]_pad  & n14927 ;
  assign n18983 = ~n18981 & ~n18982 ;
  assign n18984 = \s10_data_i[0]_pad  & n14892 ;
  assign n18985 = \s7_data_i[0]_pad  & n14740 ;
  assign n18986 = ~n18984 & ~n18985 ;
  assign n18987 = n18983 & n18986 ;
  assign n18988 = n18980 & n18987 ;
  assign n18989 = \s11_data_i[0]_pad  & n14896 ;
  assign n18990 = \s13_data_i[0]_pad  & n14904 ;
  assign n18991 = \s3_data_i[0]_pad  & n14801 ;
  assign n18992 = ~n18990 & ~n18991 ;
  assign n18993 = ~n18989 & n18992 ;
  assign n18994 = \s12_data_i[0]_pad  & n14900 ;
  assign n18995 = \s14_data_i[0]_pad  & n14915 ;
  assign n18996 = ~n18994 & ~n18995 ;
  assign n18997 = \s2_data_i[0]_pad  & n14911 ;
  assign n18998 = \s0_data_i[0]_pad  & n14603 ;
  assign n18999 = ~n18997 & ~n18998 ;
  assign n19000 = n18996 & n18999 ;
  assign n19001 = n18993 & n19000 ;
  assign n19002 = n18988 & n19001 ;
  assign n19003 = n18973 & n19002 ;
  assign n19004 = n2190 & n15229 ;
  assign n19005 = \s15_data_i[10]_pad  & n2190 ;
  assign n19006 = ~n2258 & n19005 ;
  assign n19007 = ~n19004 & ~n19006 ;
  assign n19008 = \s8_data_i[10]_pad  & n14923 ;
  assign n19009 = \s13_data_i[10]_pad  & n14904 ;
  assign n19010 = ~n19008 & ~n19009 ;
  assign n19011 = \s10_data_i[10]_pad  & n14892 ;
  assign n19012 = \s1_data_i[10]_pad  & n14609 ;
  assign n19013 = ~n19011 & ~n19012 ;
  assign n19014 = n19010 & n19013 ;
  assign n19015 = \s5_data_i[10]_pad  & n14757 ;
  assign n19016 = \s6_data_i[10]_pad  & n14745 ;
  assign n19017 = ~n19015 & ~n19016 ;
  assign n19018 = \s7_data_i[10]_pad  & n14740 ;
  assign n19019 = \s2_data_i[10]_pad  & n14911 ;
  assign n19020 = ~n19018 & ~n19019 ;
  assign n19021 = n19017 & n19020 ;
  assign n19022 = n19014 & n19021 ;
  assign n19023 = \s11_data_i[10]_pad  & n14896 ;
  assign n19024 = \s4_data_i[10]_pad  & n14919 ;
  assign n19025 = \s3_data_i[10]_pad  & n14801 ;
  assign n19026 = ~n19024 & ~n19025 ;
  assign n19027 = ~n19023 & n19026 ;
  assign n19028 = \s12_data_i[10]_pad  & n14900 ;
  assign n19029 = \s14_data_i[10]_pad  & n14915 ;
  assign n19030 = ~n19028 & ~n19029 ;
  assign n19031 = \s0_data_i[10]_pad  & n14603 ;
  assign n19032 = \s9_data_i[10]_pad  & n14927 ;
  assign n19033 = ~n19031 & ~n19032 ;
  assign n19034 = n19030 & n19033 ;
  assign n19035 = n19027 & n19034 ;
  assign n19036 = n19022 & n19035 ;
  assign n19037 = n19007 & n19036 ;
  assign n19038 = n2190 & n15266 ;
  assign n19039 = \s15_data_i[11]_pad  & n2190 ;
  assign n19040 = ~n2258 & n19039 ;
  assign n19041 = ~n19038 & ~n19040 ;
  assign n19042 = \s8_data_i[11]_pad  & n14923 ;
  assign n19043 = \s13_data_i[11]_pad  & n14904 ;
  assign n19044 = ~n19042 & ~n19043 ;
  assign n19045 = \s10_data_i[11]_pad  & n14892 ;
  assign n19046 = \s1_data_i[11]_pad  & n14609 ;
  assign n19047 = ~n19045 & ~n19046 ;
  assign n19048 = n19044 & n19047 ;
  assign n19049 = \s5_data_i[11]_pad  & n14757 ;
  assign n19050 = \s6_data_i[11]_pad  & n14745 ;
  assign n19051 = ~n19049 & ~n19050 ;
  assign n19052 = \s7_data_i[11]_pad  & n14740 ;
  assign n19053 = \s2_data_i[11]_pad  & n14911 ;
  assign n19054 = ~n19052 & ~n19053 ;
  assign n19055 = n19051 & n19054 ;
  assign n19056 = n19048 & n19055 ;
  assign n19057 = \s11_data_i[11]_pad  & n14896 ;
  assign n19058 = \s4_data_i[11]_pad  & n14919 ;
  assign n19059 = \s3_data_i[11]_pad  & n14801 ;
  assign n19060 = ~n19058 & ~n19059 ;
  assign n19061 = ~n19057 & n19060 ;
  assign n19062 = \s12_data_i[11]_pad  & n14900 ;
  assign n19063 = \s14_data_i[11]_pad  & n14915 ;
  assign n19064 = ~n19062 & ~n19063 ;
  assign n19065 = \s0_data_i[11]_pad  & n14603 ;
  assign n19066 = \s9_data_i[11]_pad  & n14927 ;
  assign n19067 = ~n19065 & ~n19066 ;
  assign n19068 = n19064 & n19067 ;
  assign n19069 = n19061 & n19068 ;
  assign n19070 = n19056 & n19069 ;
  assign n19071 = n19041 & n19070 ;
  assign n19072 = n2190 & n15303 ;
  assign n19073 = \s15_data_i[12]_pad  & n2190 ;
  assign n19074 = ~n2258 & n19073 ;
  assign n19075 = ~n19072 & ~n19074 ;
  assign n19076 = \s8_data_i[12]_pad  & n14923 ;
  assign n19077 = \s13_data_i[12]_pad  & n14904 ;
  assign n19078 = ~n19076 & ~n19077 ;
  assign n19079 = \s10_data_i[12]_pad  & n14892 ;
  assign n19080 = \s1_data_i[12]_pad  & n14609 ;
  assign n19081 = ~n19079 & ~n19080 ;
  assign n19082 = n19078 & n19081 ;
  assign n19083 = \s5_data_i[12]_pad  & n14757 ;
  assign n19084 = \s6_data_i[12]_pad  & n14745 ;
  assign n19085 = ~n19083 & ~n19084 ;
  assign n19086 = \s7_data_i[12]_pad  & n14740 ;
  assign n19087 = \s2_data_i[12]_pad  & n14911 ;
  assign n19088 = ~n19086 & ~n19087 ;
  assign n19089 = n19085 & n19088 ;
  assign n19090 = n19082 & n19089 ;
  assign n19091 = \s11_data_i[12]_pad  & n14896 ;
  assign n19092 = \s4_data_i[12]_pad  & n14919 ;
  assign n19093 = \s3_data_i[12]_pad  & n14801 ;
  assign n19094 = ~n19092 & ~n19093 ;
  assign n19095 = ~n19091 & n19094 ;
  assign n19096 = \s12_data_i[12]_pad  & n14900 ;
  assign n19097 = \s14_data_i[12]_pad  & n14915 ;
  assign n19098 = ~n19096 & ~n19097 ;
  assign n19099 = \s0_data_i[12]_pad  & n14603 ;
  assign n19100 = \s9_data_i[12]_pad  & n14927 ;
  assign n19101 = ~n19099 & ~n19100 ;
  assign n19102 = n19098 & n19101 ;
  assign n19103 = n19095 & n19102 ;
  assign n19104 = n19090 & n19103 ;
  assign n19105 = n19075 & n19104 ;
  assign n19106 = n2190 & n15340 ;
  assign n19107 = \s15_data_i[13]_pad  & n2190 ;
  assign n19108 = ~n2258 & n19107 ;
  assign n19109 = ~n19106 & ~n19108 ;
  assign n19110 = \s8_data_i[13]_pad  & n14923 ;
  assign n19111 = \s1_data_i[13]_pad  & n14609 ;
  assign n19112 = ~n19110 & ~n19111 ;
  assign n19113 = \s4_data_i[13]_pad  & n14919 ;
  assign n19114 = \s6_data_i[13]_pad  & n14745 ;
  assign n19115 = ~n19113 & ~n19114 ;
  assign n19116 = n19112 & n19115 ;
  assign n19117 = \s5_data_i[13]_pad  & n14757 ;
  assign n19118 = \s9_data_i[13]_pad  & n14927 ;
  assign n19119 = ~n19117 & ~n19118 ;
  assign n19120 = \s10_data_i[13]_pad  & n14892 ;
  assign n19121 = \s7_data_i[13]_pad  & n14740 ;
  assign n19122 = ~n19120 & ~n19121 ;
  assign n19123 = n19119 & n19122 ;
  assign n19124 = n19116 & n19123 ;
  assign n19125 = \s11_data_i[13]_pad  & n14896 ;
  assign n19126 = \s13_data_i[13]_pad  & n14904 ;
  assign n19127 = \s3_data_i[13]_pad  & n14801 ;
  assign n19128 = ~n19126 & ~n19127 ;
  assign n19129 = ~n19125 & n19128 ;
  assign n19130 = \s12_data_i[13]_pad  & n14900 ;
  assign n19131 = \s14_data_i[13]_pad  & n14915 ;
  assign n19132 = ~n19130 & ~n19131 ;
  assign n19133 = \s2_data_i[13]_pad  & n14911 ;
  assign n19134 = \s0_data_i[13]_pad  & n14603 ;
  assign n19135 = ~n19133 & ~n19134 ;
  assign n19136 = n19132 & n19135 ;
  assign n19137 = n19129 & n19136 ;
  assign n19138 = n19124 & n19137 ;
  assign n19139 = n19109 & n19138 ;
  assign n19140 = n2190 & n15377 ;
  assign n19141 = \s15_data_i[14]_pad  & n2190 ;
  assign n19142 = ~n2258 & n19141 ;
  assign n19143 = ~n19140 & ~n19142 ;
  assign n19144 = \s8_data_i[14]_pad  & n14923 ;
  assign n19145 = \s4_data_i[14]_pad  & n14919 ;
  assign n19146 = ~n19144 & ~n19145 ;
  assign n19147 = \s7_data_i[14]_pad  & n14740 ;
  assign n19148 = \s1_data_i[14]_pad  & n14609 ;
  assign n19149 = ~n19147 & ~n19148 ;
  assign n19150 = n19146 & n19149 ;
  assign n19151 = \s5_data_i[14]_pad  & n14757 ;
  assign n19152 = \s6_data_i[14]_pad  & n14745 ;
  assign n19153 = ~n19151 & ~n19152 ;
  assign n19154 = \s13_data_i[14]_pad  & n14904 ;
  assign n19155 = \s2_data_i[14]_pad  & n14911 ;
  assign n19156 = ~n19154 & ~n19155 ;
  assign n19157 = n19153 & n19156 ;
  assign n19158 = n19150 & n19157 ;
  assign n19159 = \s11_data_i[14]_pad  & n14896 ;
  assign n19160 = \s10_data_i[14]_pad  & n14892 ;
  assign n19161 = \s3_data_i[14]_pad  & n14801 ;
  assign n19162 = ~n19160 & ~n19161 ;
  assign n19163 = ~n19159 & n19162 ;
  assign n19164 = \s12_data_i[14]_pad  & n14900 ;
  assign n19165 = \s14_data_i[14]_pad  & n14915 ;
  assign n19166 = ~n19164 & ~n19165 ;
  assign n19167 = \s0_data_i[14]_pad  & n14603 ;
  assign n19168 = \s9_data_i[14]_pad  & n14927 ;
  assign n19169 = ~n19167 & ~n19168 ;
  assign n19170 = n19166 & n19169 ;
  assign n19171 = n19163 & n19170 ;
  assign n19172 = n19158 & n19171 ;
  assign n19173 = n19143 & n19172 ;
  assign n19174 = n2190 & n15414 ;
  assign n19175 = \s15_data_i[15]_pad  & n2190 ;
  assign n19176 = ~n2258 & n19175 ;
  assign n19177 = ~n19174 & ~n19176 ;
  assign n19178 = \s8_data_i[15]_pad  & n14923 ;
  assign n19179 = \s1_data_i[15]_pad  & n14609 ;
  assign n19180 = ~n19178 & ~n19179 ;
  assign n19181 = \s4_data_i[15]_pad  & n14919 ;
  assign n19182 = \s6_data_i[15]_pad  & n14745 ;
  assign n19183 = ~n19181 & ~n19182 ;
  assign n19184 = n19180 & n19183 ;
  assign n19185 = \s5_data_i[15]_pad  & n14757 ;
  assign n19186 = \s9_data_i[15]_pad  & n14927 ;
  assign n19187 = ~n19185 & ~n19186 ;
  assign n19188 = \s10_data_i[15]_pad  & n14892 ;
  assign n19189 = \s7_data_i[15]_pad  & n14740 ;
  assign n19190 = ~n19188 & ~n19189 ;
  assign n19191 = n19187 & n19190 ;
  assign n19192 = n19184 & n19191 ;
  assign n19193 = \s11_data_i[15]_pad  & n14896 ;
  assign n19194 = \s13_data_i[15]_pad  & n14904 ;
  assign n19195 = \s3_data_i[15]_pad  & n14801 ;
  assign n19196 = ~n19194 & ~n19195 ;
  assign n19197 = ~n19193 & n19196 ;
  assign n19198 = \s12_data_i[15]_pad  & n14900 ;
  assign n19199 = \s14_data_i[15]_pad  & n14915 ;
  assign n19200 = ~n19198 & ~n19199 ;
  assign n19201 = \s2_data_i[15]_pad  & n14911 ;
  assign n19202 = \s0_data_i[15]_pad  & n14603 ;
  assign n19203 = ~n19201 & ~n19202 ;
  assign n19204 = n19200 & n19203 ;
  assign n19205 = n19197 & n19204 ;
  assign n19206 = n19192 & n19205 ;
  assign n19207 = n19177 & n19206 ;
  assign n19208 = \s15_data_i[16]_pad  & n2190 ;
  assign n19209 = ~n2258 & n19208 ;
  assign n19210 = \s12_data_i[16]_pad  & n14900 ;
  assign n19211 = \s13_data_i[16]_pad  & n14904 ;
  assign n19212 = ~n19210 & ~n19211 ;
  assign n19213 = \s10_data_i[16]_pad  & n14892 ;
  assign n19214 = \s1_data_i[16]_pad  & n14609 ;
  assign n19215 = ~n19213 & ~n19214 ;
  assign n19216 = n19212 & n19215 ;
  assign n19217 = \s5_data_i[16]_pad  & n14757 ;
  assign n19218 = \s6_data_i[16]_pad  & n14745 ;
  assign n19219 = ~n19217 & ~n19218 ;
  assign n19220 = \s7_data_i[16]_pad  & n14740 ;
  assign n19221 = \s2_data_i[16]_pad  & n14911 ;
  assign n19222 = ~n19220 & ~n19221 ;
  assign n19223 = n19219 & n19222 ;
  assign n19224 = n19216 & n19223 ;
  assign n19225 = \s14_data_i[16]_pad  & n14915 ;
  assign n19226 = \s4_data_i[16]_pad  & n14919 ;
  assign n19227 = \s3_data_i[16]_pad  & n14801 ;
  assign n19228 = ~n19226 & ~n19227 ;
  assign n19229 = ~n19225 & n19228 ;
  assign n19230 = \s8_data_i[16]_pad  & n14923 ;
  assign n19231 = \s11_data_i[16]_pad  & n14896 ;
  assign n19232 = ~n19230 & ~n19231 ;
  assign n19233 = \s0_data_i[16]_pad  & n14603 ;
  assign n19234 = \s9_data_i[16]_pad  & n14927 ;
  assign n19235 = ~n19233 & ~n19234 ;
  assign n19236 = n19232 & n19235 ;
  assign n19237 = n19229 & n19236 ;
  assign n19238 = n19224 & n19237 ;
  assign n19239 = ~n19209 & n19238 ;
  assign n19240 = \s15_data_i[17]_pad  & n2190 ;
  assign n19241 = ~n2258 & n19240 ;
  assign n19242 = \s12_data_i[17]_pad  & n14900 ;
  assign n19243 = \s13_data_i[17]_pad  & n14904 ;
  assign n19244 = ~n19242 & ~n19243 ;
  assign n19245 = \s10_data_i[17]_pad  & n14892 ;
  assign n19246 = \s1_data_i[17]_pad  & n14609 ;
  assign n19247 = ~n19245 & ~n19246 ;
  assign n19248 = n19244 & n19247 ;
  assign n19249 = \s5_data_i[17]_pad  & n14757 ;
  assign n19250 = \s6_data_i[17]_pad  & n14745 ;
  assign n19251 = ~n19249 & ~n19250 ;
  assign n19252 = \s7_data_i[17]_pad  & n14740 ;
  assign n19253 = \s2_data_i[17]_pad  & n14911 ;
  assign n19254 = ~n19252 & ~n19253 ;
  assign n19255 = n19251 & n19254 ;
  assign n19256 = n19248 & n19255 ;
  assign n19257 = \s14_data_i[17]_pad  & n14915 ;
  assign n19258 = \s4_data_i[17]_pad  & n14919 ;
  assign n19259 = \s3_data_i[17]_pad  & n14801 ;
  assign n19260 = ~n19258 & ~n19259 ;
  assign n19261 = ~n19257 & n19260 ;
  assign n19262 = \s8_data_i[17]_pad  & n14923 ;
  assign n19263 = \s11_data_i[17]_pad  & n14896 ;
  assign n19264 = ~n19262 & ~n19263 ;
  assign n19265 = \s0_data_i[17]_pad  & n14603 ;
  assign n19266 = \s9_data_i[17]_pad  & n14927 ;
  assign n19267 = ~n19265 & ~n19266 ;
  assign n19268 = n19264 & n19267 ;
  assign n19269 = n19261 & n19268 ;
  assign n19270 = n19256 & n19269 ;
  assign n19271 = ~n19241 & n19270 ;
  assign n19272 = \s15_data_i[18]_pad  & n2190 ;
  assign n19273 = ~n2258 & n19272 ;
  assign n19274 = \s12_data_i[18]_pad  & n14900 ;
  assign n19275 = \s13_data_i[18]_pad  & n14904 ;
  assign n19276 = ~n19274 & ~n19275 ;
  assign n19277 = \s10_data_i[18]_pad  & n14892 ;
  assign n19278 = \s1_data_i[18]_pad  & n14609 ;
  assign n19279 = ~n19277 & ~n19278 ;
  assign n19280 = n19276 & n19279 ;
  assign n19281 = \s5_data_i[18]_pad  & n14757 ;
  assign n19282 = \s6_data_i[18]_pad  & n14745 ;
  assign n19283 = ~n19281 & ~n19282 ;
  assign n19284 = \s7_data_i[18]_pad  & n14740 ;
  assign n19285 = \s2_data_i[18]_pad  & n14911 ;
  assign n19286 = ~n19284 & ~n19285 ;
  assign n19287 = n19283 & n19286 ;
  assign n19288 = n19280 & n19287 ;
  assign n19289 = \s14_data_i[18]_pad  & n14915 ;
  assign n19290 = \s4_data_i[18]_pad  & n14919 ;
  assign n19291 = \s3_data_i[18]_pad  & n14801 ;
  assign n19292 = ~n19290 & ~n19291 ;
  assign n19293 = ~n19289 & n19292 ;
  assign n19294 = \s8_data_i[18]_pad  & n14923 ;
  assign n19295 = \s11_data_i[18]_pad  & n14896 ;
  assign n19296 = ~n19294 & ~n19295 ;
  assign n19297 = \s0_data_i[18]_pad  & n14603 ;
  assign n19298 = \s9_data_i[18]_pad  & n14927 ;
  assign n19299 = ~n19297 & ~n19298 ;
  assign n19300 = n19296 & n19299 ;
  assign n19301 = n19293 & n19300 ;
  assign n19302 = n19288 & n19301 ;
  assign n19303 = ~n19273 & n19302 ;
  assign n19304 = \s15_data_i[19]_pad  & n2190 ;
  assign n19305 = ~n2258 & n19304 ;
  assign n19306 = \s12_data_i[19]_pad  & n14900 ;
  assign n19307 = \s13_data_i[19]_pad  & n14904 ;
  assign n19308 = ~n19306 & ~n19307 ;
  assign n19309 = \s10_data_i[19]_pad  & n14892 ;
  assign n19310 = \s1_data_i[19]_pad  & n14609 ;
  assign n19311 = ~n19309 & ~n19310 ;
  assign n19312 = n19308 & n19311 ;
  assign n19313 = \s5_data_i[19]_pad  & n14757 ;
  assign n19314 = \s6_data_i[19]_pad  & n14745 ;
  assign n19315 = ~n19313 & ~n19314 ;
  assign n19316 = \s7_data_i[19]_pad  & n14740 ;
  assign n19317 = \s2_data_i[19]_pad  & n14911 ;
  assign n19318 = ~n19316 & ~n19317 ;
  assign n19319 = n19315 & n19318 ;
  assign n19320 = n19312 & n19319 ;
  assign n19321 = \s14_data_i[19]_pad  & n14915 ;
  assign n19322 = \s4_data_i[19]_pad  & n14919 ;
  assign n19323 = \s3_data_i[19]_pad  & n14801 ;
  assign n19324 = ~n19322 & ~n19323 ;
  assign n19325 = ~n19321 & n19324 ;
  assign n19326 = \s8_data_i[19]_pad  & n14923 ;
  assign n19327 = \s11_data_i[19]_pad  & n14896 ;
  assign n19328 = ~n19326 & ~n19327 ;
  assign n19329 = \s0_data_i[19]_pad  & n14603 ;
  assign n19330 = \s9_data_i[19]_pad  & n14927 ;
  assign n19331 = ~n19329 & ~n19330 ;
  assign n19332 = n19328 & n19331 ;
  assign n19333 = n19325 & n19332 ;
  assign n19334 = n19320 & n19333 ;
  assign n19335 = ~n19305 & n19334 ;
  assign n19336 = n2190 & n15579 ;
  assign n19337 = \s15_data_i[1]_pad  & n2190 ;
  assign n19338 = ~n2258 & n19337 ;
  assign n19339 = ~n19336 & ~n19338 ;
  assign n19340 = \s8_data_i[1]_pad  & n14923 ;
  assign n19341 = \s1_data_i[1]_pad  & n14609 ;
  assign n19342 = ~n19340 & ~n19341 ;
  assign n19343 = \s4_data_i[1]_pad  & n14919 ;
  assign n19344 = \s6_data_i[1]_pad  & n14745 ;
  assign n19345 = ~n19343 & ~n19344 ;
  assign n19346 = n19342 & n19345 ;
  assign n19347 = \s5_data_i[1]_pad  & n14757 ;
  assign n19348 = \s9_data_i[1]_pad  & n14927 ;
  assign n19349 = ~n19347 & ~n19348 ;
  assign n19350 = \s10_data_i[1]_pad  & n14892 ;
  assign n19351 = \s7_data_i[1]_pad  & n14740 ;
  assign n19352 = ~n19350 & ~n19351 ;
  assign n19353 = n19349 & n19352 ;
  assign n19354 = n19346 & n19353 ;
  assign n19355 = \s11_data_i[1]_pad  & n14896 ;
  assign n19356 = \s13_data_i[1]_pad  & n14904 ;
  assign n19357 = \s3_data_i[1]_pad  & n14801 ;
  assign n19358 = ~n19356 & ~n19357 ;
  assign n19359 = ~n19355 & n19358 ;
  assign n19360 = \s12_data_i[1]_pad  & n14900 ;
  assign n19361 = \s14_data_i[1]_pad  & n14915 ;
  assign n19362 = ~n19360 & ~n19361 ;
  assign n19363 = \s2_data_i[1]_pad  & n14911 ;
  assign n19364 = \s0_data_i[1]_pad  & n14603 ;
  assign n19365 = ~n19363 & ~n19364 ;
  assign n19366 = n19362 & n19365 ;
  assign n19367 = n19359 & n19366 ;
  assign n19368 = n19354 & n19367 ;
  assign n19369 = n19339 & n19368 ;
  assign n19370 = \s15_data_i[20]_pad  & n2190 ;
  assign n19371 = ~n2258 & n19370 ;
  assign n19372 = \s12_data_i[20]_pad  & n14900 ;
  assign n19373 = \s13_data_i[20]_pad  & n14904 ;
  assign n19374 = ~n19372 & ~n19373 ;
  assign n19375 = \s10_data_i[20]_pad  & n14892 ;
  assign n19376 = \s1_data_i[20]_pad  & n14609 ;
  assign n19377 = ~n19375 & ~n19376 ;
  assign n19378 = n19374 & n19377 ;
  assign n19379 = \s5_data_i[20]_pad  & n14757 ;
  assign n19380 = \s6_data_i[20]_pad  & n14745 ;
  assign n19381 = ~n19379 & ~n19380 ;
  assign n19382 = \s7_data_i[20]_pad  & n14740 ;
  assign n19383 = \s2_data_i[20]_pad  & n14911 ;
  assign n19384 = ~n19382 & ~n19383 ;
  assign n19385 = n19381 & n19384 ;
  assign n19386 = n19378 & n19385 ;
  assign n19387 = \s14_data_i[20]_pad  & n14915 ;
  assign n19388 = \s4_data_i[20]_pad  & n14919 ;
  assign n19389 = \s3_data_i[20]_pad  & n14801 ;
  assign n19390 = ~n19388 & ~n19389 ;
  assign n19391 = ~n19387 & n19390 ;
  assign n19392 = \s8_data_i[20]_pad  & n14923 ;
  assign n19393 = \s11_data_i[20]_pad  & n14896 ;
  assign n19394 = ~n19392 & ~n19393 ;
  assign n19395 = \s0_data_i[20]_pad  & n14603 ;
  assign n19396 = \s9_data_i[20]_pad  & n14927 ;
  assign n19397 = ~n19395 & ~n19396 ;
  assign n19398 = n19394 & n19397 ;
  assign n19399 = n19391 & n19398 ;
  assign n19400 = n19386 & n19399 ;
  assign n19401 = ~n19371 & n19400 ;
  assign n19402 = \s15_data_i[21]_pad  & n2190 ;
  assign n19403 = ~n2258 & n19402 ;
  assign n19404 = \s12_data_i[21]_pad  & n14900 ;
  assign n19405 = \s13_data_i[21]_pad  & n14904 ;
  assign n19406 = ~n19404 & ~n19405 ;
  assign n19407 = \s10_data_i[21]_pad  & n14892 ;
  assign n19408 = \s1_data_i[21]_pad  & n14609 ;
  assign n19409 = ~n19407 & ~n19408 ;
  assign n19410 = n19406 & n19409 ;
  assign n19411 = \s5_data_i[21]_pad  & n14757 ;
  assign n19412 = \s6_data_i[21]_pad  & n14745 ;
  assign n19413 = ~n19411 & ~n19412 ;
  assign n19414 = \s7_data_i[21]_pad  & n14740 ;
  assign n19415 = \s2_data_i[21]_pad  & n14911 ;
  assign n19416 = ~n19414 & ~n19415 ;
  assign n19417 = n19413 & n19416 ;
  assign n19418 = n19410 & n19417 ;
  assign n19419 = \s14_data_i[21]_pad  & n14915 ;
  assign n19420 = \s4_data_i[21]_pad  & n14919 ;
  assign n19421 = \s3_data_i[21]_pad  & n14801 ;
  assign n19422 = ~n19420 & ~n19421 ;
  assign n19423 = ~n19419 & n19422 ;
  assign n19424 = \s8_data_i[21]_pad  & n14923 ;
  assign n19425 = \s11_data_i[21]_pad  & n14896 ;
  assign n19426 = ~n19424 & ~n19425 ;
  assign n19427 = \s0_data_i[21]_pad  & n14603 ;
  assign n19428 = \s9_data_i[21]_pad  & n14927 ;
  assign n19429 = ~n19427 & ~n19428 ;
  assign n19430 = n19426 & n19429 ;
  assign n19431 = n19423 & n19430 ;
  assign n19432 = n19418 & n19431 ;
  assign n19433 = ~n19403 & n19432 ;
  assign n19434 = \s15_data_i[22]_pad  & n2190 ;
  assign n19435 = ~n2258 & n19434 ;
  assign n19436 = \s12_data_i[22]_pad  & n14900 ;
  assign n19437 = \s13_data_i[22]_pad  & n14904 ;
  assign n19438 = ~n19436 & ~n19437 ;
  assign n19439 = \s10_data_i[22]_pad  & n14892 ;
  assign n19440 = \s1_data_i[22]_pad  & n14609 ;
  assign n19441 = ~n19439 & ~n19440 ;
  assign n19442 = n19438 & n19441 ;
  assign n19443 = \s5_data_i[22]_pad  & n14757 ;
  assign n19444 = \s6_data_i[22]_pad  & n14745 ;
  assign n19445 = ~n19443 & ~n19444 ;
  assign n19446 = \s7_data_i[22]_pad  & n14740 ;
  assign n19447 = \s2_data_i[22]_pad  & n14911 ;
  assign n19448 = ~n19446 & ~n19447 ;
  assign n19449 = n19445 & n19448 ;
  assign n19450 = n19442 & n19449 ;
  assign n19451 = \s14_data_i[22]_pad  & n14915 ;
  assign n19452 = \s4_data_i[22]_pad  & n14919 ;
  assign n19453 = \s3_data_i[22]_pad  & n14801 ;
  assign n19454 = ~n19452 & ~n19453 ;
  assign n19455 = ~n19451 & n19454 ;
  assign n19456 = \s8_data_i[22]_pad  & n14923 ;
  assign n19457 = \s11_data_i[22]_pad  & n14896 ;
  assign n19458 = ~n19456 & ~n19457 ;
  assign n19459 = \s0_data_i[22]_pad  & n14603 ;
  assign n19460 = \s9_data_i[22]_pad  & n14927 ;
  assign n19461 = ~n19459 & ~n19460 ;
  assign n19462 = n19458 & n19461 ;
  assign n19463 = n19455 & n19462 ;
  assign n19464 = n19450 & n19463 ;
  assign n19465 = ~n19435 & n19464 ;
  assign n19466 = \s15_data_i[23]_pad  & n2190 ;
  assign n19467 = ~n2258 & n19466 ;
  assign n19468 = \s12_data_i[23]_pad  & n14900 ;
  assign n19469 = \s13_data_i[23]_pad  & n14904 ;
  assign n19470 = ~n19468 & ~n19469 ;
  assign n19471 = \s10_data_i[23]_pad  & n14892 ;
  assign n19472 = \s1_data_i[23]_pad  & n14609 ;
  assign n19473 = ~n19471 & ~n19472 ;
  assign n19474 = n19470 & n19473 ;
  assign n19475 = \s5_data_i[23]_pad  & n14757 ;
  assign n19476 = \s6_data_i[23]_pad  & n14745 ;
  assign n19477 = ~n19475 & ~n19476 ;
  assign n19478 = \s7_data_i[23]_pad  & n14740 ;
  assign n19479 = \s2_data_i[23]_pad  & n14911 ;
  assign n19480 = ~n19478 & ~n19479 ;
  assign n19481 = n19477 & n19480 ;
  assign n19482 = n19474 & n19481 ;
  assign n19483 = \s14_data_i[23]_pad  & n14915 ;
  assign n19484 = \s4_data_i[23]_pad  & n14919 ;
  assign n19485 = \s3_data_i[23]_pad  & n14801 ;
  assign n19486 = ~n19484 & ~n19485 ;
  assign n19487 = ~n19483 & n19486 ;
  assign n19488 = \s8_data_i[23]_pad  & n14923 ;
  assign n19489 = \s11_data_i[23]_pad  & n14896 ;
  assign n19490 = ~n19488 & ~n19489 ;
  assign n19491 = \s0_data_i[23]_pad  & n14603 ;
  assign n19492 = \s9_data_i[23]_pad  & n14927 ;
  assign n19493 = ~n19491 & ~n19492 ;
  assign n19494 = n19490 & n19493 ;
  assign n19495 = n19487 & n19494 ;
  assign n19496 = n19482 & n19495 ;
  assign n19497 = ~n19467 & n19496 ;
  assign n19498 = \s15_data_i[24]_pad  & n2190 ;
  assign n19499 = ~n2258 & n19498 ;
  assign n19500 = \s12_data_i[24]_pad  & n14900 ;
  assign n19501 = \s13_data_i[24]_pad  & n14904 ;
  assign n19502 = ~n19500 & ~n19501 ;
  assign n19503 = \s10_data_i[24]_pad  & n14892 ;
  assign n19504 = \s1_data_i[24]_pad  & n14609 ;
  assign n19505 = ~n19503 & ~n19504 ;
  assign n19506 = n19502 & n19505 ;
  assign n19507 = \s5_data_i[24]_pad  & n14757 ;
  assign n19508 = \s6_data_i[24]_pad  & n14745 ;
  assign n19509 = ~n19507 & ~n19508 ;
  assign n19510 = \s7_data_i[24]_pad  & n14740 ;
  assign n19511 = \s2_data_i[24]_pad  & n14911 ;
  assign n19512 = ~n19510 & ~n19511 ;
  assign n19513 = n19509 & n19512 ;
  assign n19514 = n19506 & n19513 ;
  assign n19515 = \s14_data_i[24]_pad  & n14915 ;
  assign n19516 = \s4_data_i[24]_pad  & n14919 ;
  assign n19517 = \s3_data_i[24]_pad  & n14801 ;
  assign n19518 = ~n19516 & ~n19517 ;
  assign n19519 = ~n19515 & n19518 ;
  assign n19520 = \s8_data_i[24]_pad  & n14923 ;
  assign n19521 = \s11_data_i[24]_pad  & n14896 ;
  assign n19522 = ~n19520 & ~n19521 ;
  assign n19523 = \s0_data_i[24]_pad  & n14603 ;
  assign n19524 = \s9_data_i[24]_pad  & n14927 ;
  assign n19525 = ~n19523 & ~n19524 ;
  assign n19526 = n19522 & n19525 ;
  assign n19527 = n19519 & n19526 ;
  assign n19528 = n19514 & n19527 ;
  assign n19529 = ~n19499 & n19528 ;
  assign n19530 = \s15_data_i[25]_pad  & n2190 ;
  assign n19531 = ~n2258 & n19530 ;
  assign n19532 = \s12_data_i[25]_pad  & n14900 ;
  assign n19533 = \s13_data_i[25]_pad  & n14904 ;
  assign n19534 = ~n19532 & ~n19533 ;
  assign n19535 = \s10_data_i[25]_pad  & n14892 ;
  assign n19536 = \s1_data_i[25]_pad  & n14609 ;
  assign n19537 = ~n19535 & ~n19536 ;
  assign n19538 = n19534 & n19537 ;
  assign n19539 = \s5_data_i[25]_pad  & n14757 ;
  assign n19540 = \s6_data_i[25]_pad  & n14745 ;
  assign n19541 = ~n19539 & ~n19540 ;
  assign n19542 = \s7_data_i[25]_pad  & n14740 ;
  assign n19543 = \s2_data_i[25]_pad  & n14911 ;
  assign n19544 = ~n19542 & ~n19543 ;
  assign n19545 = n19541 & n19544 ;
  assign n19546 = n19538 & n19545 ;
  assign n19547 = \s14_data_i[25]_pad  & n14915 ;
  assign n19548 = \s4_data_i[25]_pad  & n14919 ;
  assign n19549 = \s3_data_i[25]_pad  & n14801 ;
  assign n19550 = ~n19548 & ~n19549 ;
  assign n19551 = ~n19547 & n19550 ;
  assign n19552 = \s8_data_i[25]_pad  & n14923 ;
  assign n19553 = \s11_data_i[25]_pad  & n14896 ;
  assign n19554 = ~n19552 & ~n19553 ;
  assign n19555 = \s0_data_i[25]_pad  & n14603 ;
  assign n19556 = \s9_data_i[25]_pad  & n14927 ;
  assign n19557 = ~n19555 & ~n19556 ;
  assign n19558 = n19554 & n19557 ;
  assign n19559 = n19551 & n19558 ;
  assign n19560 = n19546 & n19559 ;
  assign n19561 = ~n19531 & n19560 ;
  assign n19562 = \s15_data_i[26]_pad  & n2190 ;
  assign n19563 = ~n2258 & n19562 ;
  assign n19564 = \s12_data_i[26]_pad  & n14900 ;
  assign n19565 = \s13_data_i[26]_pad  & n14904 ;
  assign n19566 = ~n19564 & ~n19565 ;
  assign n19567 = \s10_data_i[26]_pad  & n14892 ;
  assign n19568 = \s1_data_i[26]_pad  & n14609 ;
  assign n19569 = ~n19567 & ~n19568 ;
  assign n19570 = n19566 & n19569 ;
  assign n19571 = \s5_data_i[26]_pad  & n14757 ;
  assign n19572 = \s6_data_i[26]_pad  & n14745 ;
  assign n19573 = ~n19571 & ~n19572 ;
  assign n19574 = \s7_data_i[26]_pad  & n14740 ;
  assign n19575 = \s2_data_i[26]_pad  & n14911 ;
  assign n19576 = ~n19574 & ~n19575 ;
  assign n19577 = n19573 & n19576 ;
  assign n19578 = n19570 & n19577 ;
  assign n19579 = \s14_data_i[26]_pad  & n14915 ;
  assign n19580 = \s4_data_i[26]_pad  & n14919 ;
  assign n19581 = \s3_data_i[26]_pad  & n14801 ;
  assign n19582 = ~n19580 & ~n19581 ;
  assign n19583 = ~n19579 & n19582 ;
  assign n19584 = \s8_data_i[26]_pad  & n14923 ;
  assign n19585 = \s11_data_i[26]_pad  & n14896 ;
  assign n19586 = ~n19584 & ~n19585 ;
  assign n19587 = \s0_data_i[26]_pad  & n14603 ;
  assign n19588 = \s9_data_i[26]_pad  & n14927 ;
  assign n19589 = ~n19587 & ~n19588 ;
  assign n19590 = n19586 & n19589 ;
  assign n19591 = n19583 & n19590 ;
  assign n19592 = n19578 & n19591 ;
  assign n19593 = ~n19563 & n19592 ;
  assign n19594 = \s15_data_i[27]_pad  & n2190 ;
  assign n19595 = ~n2258 & n19594 ;
  assign n19596 = \s12_data_i[27]_pad  & n14900 ;
  assign n19597 = \s13_data_i[27]_pad  & n14904 ;
  assign n19598 = ~n19596 & ~n19597 ;
  assign n19599 = \s10_data_i[27]_pad  & n14892 ;
  assign n19600 = \s1_data_i[27]_pad  & n14609 ;
  assign n19601 = ~n19599 & ~n19600 ;
  assign n19602 = n19598 & n19601 ;
  assign n19603 = \s5_data_i[27]_pad  & n14757 ;
  assign n19604 = \s6_data_i[27]_pad  & n14745 ;
  assign n19605 = ~n19603 & ~n19604 ;
  assign n19606 = \s7_data_i[27]_pad  & n14740 ;
  assign n19607 = \s2_data_i[27]_pad  & n14911 ;
  assign n19608 = ~n19606 & ~n19607 ;
  assign n19609 = n19605 & n19608 ;
  assign n19610 = n19602 & n19609 ;
  assign n19611 = \s14_data_i[27]_pad  & n14915 ;
  assign n19612 = \s4_data_i[27]_pad  & n14919 ;
  assign n19613 = \s3_data_i[27]_pad  & n14801 ;
  assign n19614 = ~n19612 & ~n19613 ;
  assign n19615 = ~n19611 & n19614 ;
  assign n19616 = \s8_data_i[27]_pad  & n14923 ;
  assign n19617 = \s11_data_i[27]_pad  & n14896 ;
  assign n19618 = ~n19616 & ~n19617 ;
  assign n19619 = \s0_data_i[27]_pad  & n14603 ;
  assign n19620 = \s9_data_i[27]_pad  & n14927 ;
  assign n19621 = ~n19619 & ~n19620 ;
  assign n19622 = n19618 & n19621 ;
  assign n19623 = n19615 & n19622 ;
  assign n19624 = n19610 & n19623 ;
  assign n19625 = ~n19595 & n19624 ;
  assign n19626 = \s15_data_i[28]_pad  & n2190 ;
  assign n19627 = ~n2258 & n19626 ;
  assign n19628 = \s12_data_i[28]_pad  & n14900 ;
  assign n19629 = \s13_data_i[28]_pad  & n14904 ;
  assign n19630 = ~n19628 & ~n19629 ;
  assign n19631 = \s10_data_i[28]_pad  & n14892 ;
  assign n19632 = \s1_data_i[28]_pad  & n14609 ;
  assign n19633 = ~n19631 & ~n19632 ;
  assign n19634 = n19630 & n19633 ;
  assign n19635 = \s5_data_i[28]_pad  & n14757 ;
  assign n19636 = \s6_data_i[28]_pad  & n14745 ;
  assign n19637 = ~n19635 & ~n19636 ;
  assign n19638 = \s7_data_i[28]_pad  & n14740 ;
  assign n19639 = \s2_data_i[28]_pad  & n14911 ;
  assign n19640 = ~n19638 & ~n19639 ;
  assign n19641 = n19637 & n19640 ;
  assign n19642 = n19634 & n19641 ;
  assign n19643 = \s14_data_i[28]_pad  & n14915 ;
  assign n19644 = \s4_data_i[28]_pad  & n14919 ;
  assign n19645 = \s3_data_i[28]_pad  & n14801 ;
  assign n19646 = ~n19644 & ~n19645 ;
  assign n19647 = ~n19643 & n19646 ;
  assign n19648 = \s8_data_i[28]_pad  & n14923 ;
  assign n19649 = \s11_data_i[28]_pad  & n14896 ;
  assign n19650 = ~n19648 & ~n19649 ;
  assign n19651 = \s0_data_i[28]_pad  & n14603 ;
  assign n19652 = \s9_data_i[28]_pad  & n14927 ;
  assign n19653 = ~n19651 & ~n19652 ;
  assign n19654 = n19650 & n19653 ;
  assign n19655 = n19647 & n19654 ;
  assign n19656 = n19642 & n19655 ;
  assign n19657 = ~n19627 & n19656 ;
  assign n19658 = \s15_data_i[29]_pad  & n2190 ;
  assign n19659 = ~n2258 & n19658 ;
  assign n19660 = \s12_data_i[29]_pad  & n14900 ;
  assign n19661 = \s13_data_i[29]_pad  & n14904 ;
  assign n19662 = ~n19660 & ~n19661 ;
  assign n19663 = \s10_data_i[29]_pad  & n14892 ;
  assign n19664 = \s1_data_i[29]_pad  & n14609 ;
  assign n19665 = ~n19663 & ~n19664 ;
  assign n19666 = n19662 & n19665 ;
  assign n19667 = \s5_data_i[29]_pad  & n14757 ;
  assign n19668 = \s6_data_i[29]_pad  & n14745 ;
  assign n19669 = ~n19667 & ~n19668 ;
  assign n19670 = \s7_data_i[29]_pad  & n14740 ;
  assign n19671 = \s2_data_i[29]_pad  & n14911 ;
  assign n19672 = ~n19670 & ~n19671 ;
  assign n19673 = n19669 & n19672 ;
  assign n19674 = n19666 & n19673 ;
  assign n19675 = \s14_data_i[29]_pad  & n14915 ;
  assign n19676 = \s4_data_i[29]_pad  & n14919 ;
  assign n19677 = \s3_data_i[29]_pad  & n14801 ;
  assign n19678 = ~n19676 & ~n19677 ;
  assign n19679 = ~n19675 & n19678 ;
  assign n19680 = \s8_data_i[29]_pad  & n14923 ;
  assign n19681 = \s11_data_i[29]_pad  & n14896 ;
  assign n19682 = ~n19680 & ~n19681 ;
  assign n19683 = \s0_data_i[29]_pad  & n14603 ;
  assign n19684 = \s9_data_i[29]_pad  & n14927 ;
  assign n19685 = ~n19683 & ~n19684 ;
  assign n19686 = n19682 & n19685 ;
  assign n19687 = n19679 & n19686 ;
  assign n19688 = n19674 & n19687 ;
  assign n19689 = ~n19659 & n19688 ;
  assign n19690 = n2190 & n15936 ;
  assign n19691 = \s15_data_i[2]_pad  & n2190 ;
  assign n19692 = ~n2258 & n19691 ;
  assign n19693 = ~n19690 & ~n19692 ;
  assign n19694 = \s8_data_i[2]_pad  & n14923 ;
  assign n19695 = \s1_data_i[2]_pad  & n14609 ;
  assign n19696 = ~n19694 & ~n19695 ;
  assign n19697 = \s4_data_i[2]_pad  & n14919 ;
  assign n19698 = \s6_data_i[2]_pad  & n14745 ;
  assign n19699 = ~n19697 & ~n19698 ;
  assign n19700 = n19696 & n19699 ;
  assign n19701 = \s5_data_i[2]_pad  & n14757 ;
  assign n19702 = \s9_data_i[2]_pad  & n14927 ;
  assign n19703 = ~n19701 & ~n19702 ;
  assign n19704 = \s10_data_i[2]_pad  & n14892 ;
  assign n19705 = \s7_data_i[2]_pad  & n14740 ;
  assign n19706 = ~n19704 & ~n19705 ;
  assign n19707 = n19703 & n19706 ;
  assign n19708 = n19700 & n19707 ;
  assign n19709 = \s11_data_i[2]_pad  & n14896 ;
  assign n19710 = \s13_data_i[2]_pad  & n14904 ;
  assign n19711 = \s3_data_i[2]_pad  & n14801 ;
  assign n19712 = ~n19710 & ~n19711 ;
  assign n19713 = ~n19709 & n19712 ;
  assign n19714 = \s12_data_i[2]_pad  & n14900 ;
  assign n19715 = \s14_data_i[2]_pad  & n14915 ;
  assign n19716 = ~n19714 & ~n19715 ;
  assign n19717 = \s2_data_i[2]_pad  & n14911 ;
  assign n19718 = \s0_data_i[2]_pad  & n14603 ;
  assign n19719 = ~n19717 & ~n19718 ;
  assign n19720 = n19716 & n19719 ;
  assign n19721 = n19713 & n19720 ;
  assign n19722 = n19708 & n19721 ;
  assign n19723 = n19693 & n19722 ;
  assign n19724 = \s15_data_i[30]_pad  & n2190 ;
  assign n19725 = ~n2258 & n19724 ;
  assign n19726 = \s12_data_i[30]_pad  & n14900 ;
  assign n19727 = \s13_data_i[30]_pad  & n14904 ;
  assign n19728 = ~n19726 & ~n19727 ;
  assign n19729 = \s10_data_i[30]_pad  & n14892 ;
  assign n19730 = \s1_data_i[30]_pad  & n14609 ;
  assign n19731 = ~n19729 & ~n19730 ;
  assign n19732 = n19728 & n19731 ;
  assign n19733 = \s5_data_i[30]_pad  & n14757 ;
  assign n19734 = \s6_data_i[30]_pad  & n14745 ;
  assign n19735 = ~n19733 & ~n19734 ;
  assign n19736 = \s7_data_i[30]_pad  & n14740 ;
  assign n19737 = \s2_data_i[30]_pad  & n14911 ;
  assign n19738 = ~n19736 & ~n19737 ;
  assign n19739 = n19735 & n19738 ;
  assign n19740 = n19732 & n19739 ;
  assign n19741 = \s14_data_i[30]_pad  & n14915 ;
  assign n19742 = \s4_data_i[30]_pad  & n14919 ;
  assign n19743 = \s3_data_i[30]_pad  & n14801 ;
  assign n19744 = ~n19742 & ~n19743 ;
  assign n19745 = ~n19741 & n19744 ;
  assign n19746 = \s8_data_i[30]_pad  & n14923 ;
  assign n19747 = \s11_data_i[30]_pad  & n14896 ;
  assign n19748 = ~n19746 & ~n19747 ;
  assign n19749 = \s0_data_i[30]_pad  & n14603 ;
  assign n19750 = \s9_data_i[30]_pad  & n14927 ;
  assign n19751 = ~n19749 & ~n19750 ;
  assign n19752 = n19748 & n19751 ;
  assign n19753 = n19745 & n19752 ;
  assign n19754 = n19740 & n19753 ;
  assign n19755 = ~n19725 & n19754 ;
  assign n19756 = \s15_data_i[31]_pad  & n2190 ;
  assign n19757 = ~n2258 & n19756 ;
  assign n19758 = \s12_data_i[31]_pad  & n14900 ;
  assign n19759 = \s13_data_i[31]_pad  & n14904 ;
  assign n19760 = ~n19758 & ~n19759 ;
  assign n19761 = \s10_data_i[31]_pad  & n14892 ;
  assign n19762 = \s1_data_i[31]_pad  & n14609 ;
  assign n19763 = ~n19761 & ~n19762 ;
  assign n19764 = n19760 & n19763 ;
  assign n19765 = \s5_data_i[31]_pad  & n14757 ;
  assign n19766 = \s6_data_i[31]_pad  & n14745 ;
  assign n19767 = ~n19765 & ~n19766 ;
  assign n19768 = \s7_data_i[31]_pad  & n14740 ;
  assign n19769 = \s2_data_i[31]_pad  & n14911 ;
  assign n19770 = ~n19768 & ~n19769 ;
  assign n19771 = n19767 & n19770 ;
  assign n19772 = n19764 & n19771 ;
  assign n19773 = \s14_data_i[31]_pad  & n14915 ;
  assign n19774 = \s4_data_i[31]_pad  & n14919 ;
  assign n19775 = \s3_data_i[31]_pad  & n14801 ;
  assign n19776 = ~n19774 & ~n19775 ;
  assign n19777 = ~n19773 & n19776 ;
  assign n19778 = \s8_data_i[31]_pad  & n14923 ;
  assign n19779 = \s11_data_i[31]_pad  & n14896 ;
  assign n19780 = ~n19778 & ~n19779 ;
  assign n19781 = \s0_data_i[31]_pad  & n14603 ;
  assign n19782 = \s9_data_i[31]_pad  & n14927 ;
  assign n19783 = ~n19781 & ~n19782 ;
  assign n19784 = n19780 & n19783 ;
  assign n19785 = n19777 & n19784 ;
  assign n19786 = n19772 & n19785 ;
  assign n19787 = ~n19757 & n19786 ;
  assign n19788 = n2190 & n16037 ;
  assign n19789 = \s15_data_i[3]_pad  & n2190 ;
  assign n19790 = ~n2258 & n19789 ;
  assign n19791 = ~n19788 & ~n19790 ;
  assign n19792 = \s8_data_i[3]_pad  & n14923 ;
  assign n19793 = \s13_data_i[3]_pad  & n14904 ;
  assign n19794 = ~n19792 & ~n19793 ;
  assign n19795 = \s10_data_i[3]_pad  & n14892 ;
  assign n19796 = \s1_data_i[3]_pad  & n14609 ;
  assign n19797 = ~n19795 & ~n19796 ;
  assign n19798 = n19794 & n19797 ;
  assign n19799 = \s5_data_i[3]_pad  & n14757 ;
  assign n19800 = \s6_data_i[3]_pad  & n14745 ;
  assign n19801 = ~n19799 & ~n19800 ;
  assign n19802 = \s7_data_i[3]_pad  & n14740 ;
  assign n19803 = \s2_data_i[3]_pad  & n14911 ;
  assign n19804 = ~n19802 & ~n19803 ;
  assign n19805 = n19801 & n19804 ;
  assign n19806 = n19798 & n19805 ;
  assign n19807 = \s11_data_i[3]_pad  & n14896 ;
  assign n19808 = \s4_data_i[3]_pad  & n14919 ;
  assign n19809 = \s3_data_i[3]_pad  & n14801 ;
  assign n19810 = ~n19808 & ~n19809 ;
  assign n19811 = ~n19807 & n19810 ;
  assign n19812 = \s12_data_i[3]_pad  & n14900 ;
  assign n19813 = \s14_data_i[3]_pad  & n14915 ;
  assign n19814 = ~n19812 & ~n19813 ;
  assign n19815 = \s0_data_i[3]_pad  & n14603 ;
  assign n19816 = \s9_data_i[3]_pad  & n14927 ;
  assign n19817 = ~n19815 & ~n19816 ;
  assign n19818 = n19814 & n19817 ;
  assign n19819 = n19811 & n19818 ;
  assign n19820 = n19806 & n19819 ;
  assign n19821 = n19791 & n19820 ;
  assign n19822 = n2190 & n16074 ;
  assign n19823 = \s15_data_i[4]_pad  & n2190 ;
  assign n19824 = ~n2258 & n19823 ;
  assign n19825 = ~n19822 & ~n19824 ;
  assign n19826 = \s8_data_i[4]_pad  & n14923 ;
  assign n19827 = \s4_data_i[4]_pad  & n14919 ;
  assign n19828 = ~n19826 & ~n19827 ;
  assign n19829 = \s7_data_i[4]_pad  & n14740 ;
  assign n19830 = \s1_data_i[4]_pad  & n14609 ;
  assign n19831 = ~n19829 & ~n19830 ;
  assign n19832 = n19828 & n19831 ;
  assign n19833 = \s5_data_i[4]_pad  & n14757 ;
  assign n19834 = \s6_data_i[4]_pad  & n14745 ;
  assign n19835 = ~n19833 & ~n19834 ;
  assign n19836 = \s13_data_i[4]_pad  & n14904 ;
  assign n19837 = \s2_data_i[4]_pad  & n14911 ;
  assign n19838 = ~n19836 & ~n19837 ;
  assign n19839 = n19835 & n19838 ;
  assign n19840 = n19832 & n19839 ;
  assign n19841 = \s11_data_i[4]_pad  & n14896 ;
  assign n19842 = \s10_data_i[4]_pad  & n14892 ;
  assign n19843 = \s3_data_i[4]_pad  & n14801 ;
  assign n19844 = ~n19842 & ~n19843 ;
  assign n19845 = ~n19841 & n19844 ;
  assign n19846 = \s12_data_i[4]_pad  & n14900 ;
  assign n19847 = \s14_data_i[4]_pad  & n14915 ;
  assign n19848 = ~n19846 & ~n19847 ;
  assign n19849 = \s0_data_i[4]_pad  & n14603 ;
  assign n19850 = \s9_data_i[4]_pad  & n14927 ;
  assign n19851 = ~n19849 & ~n19850 ;
  assign n19852 = n19848 & n19851 ;
  assign n19853 = n19845 & n19852 ;
  assign n19854 = n19840 & n19853 ;
  assign n19855 = n19825 & n19854 ;
  assign n19856 = n2190 & n16111 ;
  assign n19857 = \s15_data_i[5]_pad  & n2190 ;
  assign n19858 = ~n2258 & n19857 ;
  assign n19859 = ~n19856 & ~n19858 ;
  assign n19860 = \s8_data_i[5]_pad  & n14923 ;
  assign n19861 = \s13_data_i[5]_pad  & n14904 ;
  assign n19862 = ~n19860 & ~n19861 ;
  assign n19863 = \s10_data_i[5]_pad  & n14892 ;
  assign n19864 = \s1_data_i[5]_pad  & n14609 ;
  assign n19865 = ~n19863 & ~n19864 ;
  assign n19866 = n19862 & n19865 ;
  assign n19867 = \s5_data_i[5]_pad  & n14757 ;
  assign n19868 = \s6_data_i[5]_pad  & n14745 ;
  assign n19869 = ~n19867 & ~n19868 ;
  assign n19870 = \s7_data_i[5]_pad  & n14740 ;
  assign n19871 = \s2_data_i[5]_pad  & n14911 ;
  assign n19872 = ~n19870 & ~n19871 ;
  assign n19873 = n19869 & n19872 ;
  assign n19874 = n19866 & n19873 ;
  assign n19875 = \s11_data_i[5]_pad  & n14896 ;
  assign n19876 = \s4_data_i[5]_pad  & n14919 ;
  assign n19877 = \s3_data_i[5]_pad  & n14801 ;
  assign n19878 = ~n19876 & ~n19877 ;
  assign n19879 = ~n19875 & n19878 ;
  assign n19880 = \s12_data_i[5]_pad  & n14900 ;
  assign n19881 = \s14_data_i[5]_pad  & n14915 ;
  assign n19882 = ~n19880 & ~n19881 ;
  assign n19883 = \s0_data_i[5]_pad  & n14603 ;
  assign n19884 = \s9_data_i[5]_pad  & n14927 ;
  assign n19885 = ~n19883 & ~n19884 ;
  assign n19886 = n19882 & n19885 ;
  assign n19887 = n19879 & n19886 ;
  assign n19888 = n19874 & n19887 ;
  assign n19889 = n19859 & n19888 ;
  assign n19890 = n2190 & n16148 ;
  assign n19891 = \s15_data_i[6]_pad  & n2190 ;
  assign n19892 = ~n2258 & n19891 ;
  assign n19893 = ~n19890 & ~n19892 ;
  assign n19894 = \s8_data_i[6]_pad  & n14923 ;
  assign n19895 = \s13_data_i[6]_pad  & n14904 ;
  assign n19896 = ~n19894 & ~n19895 ;
  assign n19897 = \s10_data_i[6]_pad  & n14892 ;
  assign n19898 = \s1_data_i[6]_pad  & n14609 ;
  assign n19899 = ~n19897 & ~n19898 ;
  assign n19900 = n19896 & n19899 ;
  assign n19901 = \s5_data_i[6]_pad  & n14757 ;
  assign n19902 = \s6_data_i[6]_pad  & n14745 ;
  assign n19903 = ~n19901 & ~n19902 ;
  assign n19904 = \s7_data_i[6]_pad  & n14740 ;
  assign n19905 = \s2_data_i[6]_pad  & n14911 ;
  assign n19906 = ~n19904 & ~n19905 ;
  assign n19907 = n19903 & n19906 ;
  assign n19908 = n19900 & n19907 ;
  assign n19909 = \s11_data_i[6]_pad  & n14896 ;
  assign n19910 = \s4_data_i[6]_pad  & n14919 ;
  assign n19911 = \s3_data_i[6]_pad  & n14801 ;
  assign n19912 = ~n19910 & ~n19911 ;
  assign n19913 = ~n19909 & n19912 ;
  assign n19914 = \s12_data_i[6]_pad  & n14900 ;
  assign n19915 = \s14_data_i[6]_pad  & n14915 ;
  assign n19916 = ~n19914 & ~n19915 ;
  assign n19917 = \s0_data_i[6]_pad  & n14603 ;
  assign n19918 = \s9_data_i[6]_pad  & n14927 ;
  assign n19919 = ~n19917 & ~n19918 ;
  assign n19920 = n19916 & n19919 ;
  assign n19921 = n19913 & n19920 ;
  assign n19922 = n19908 & n19921 ;
  assign n19923 = n19893 & n19922 ;
  assign n19924 = n2190 & n16185 ;
  assign n19925 = \s15_data_i[7]_pad  & n2190 ;
  assign n19926 = ~n2258 & n19925 ;
  assign n19927 = ~n19924 & ~n19926 ;
  assign n19928 = \s2_data_i[7]_pad  & n14911 ;
  assign n19929 = \s13_data_i[7]_pad  & n14904 ;
  assign n19930 = ~n19928 & ~n19929 ;
  assign n19931 = \s11_data_i[7]_pad  & n14896 ;
  assign n19932 = \s6_data_i[7]_pad  & n14745 ;
  assign n19933 = ~n19931 & ~n19932 ;
  assign n19934 = n19930 & n19933 ;
  assign n19935 = \s4_data_i[7]_pad  & n14919 ;
  assign n19936 = \s3_data_i[7]_pad  & n14801 ;
  assign n19937 = ~n19935 & ~n19936 ;
  assign n19938 = \s12_data_i[7]_pad  & n14900 ;
  assign n19939 = \s7_data_i[7]_pad  & n14740 ;
  assign n19940 = ~n19938 & ~n19939 ;
  assign n19941 = n19937 & n19940 ;
  assign n19942 = n19934 & n19941 ;
  assign n19943 = \s1_data_i[7]_pad  & n14609 ;
  assign n19944 = \s8_data_i[7]_pad  & n14923 ;
  assign n19945 = \s0_data_i[7]_pad  & n14603 ;
  assign n19946 = ~n19944 & ~n19945 ;
  assign n19947 = ~n19943 & n19946 ;
  assign n19948 = \s9_data_i[7]_pad  & n14927 ;
  assign n19949 = \s10_data_i[7]_pad  & n14892 ;
  assign n19950 = ~n19948 & ~n19949 ;
  assign n19951 = \s5_data_i[7]_pad  & n14757 ;
  assign n19952 = \s14_data_i[7]_pad  & n14915 ;
  assign n19953 = ~n19951 & ~n19952 ;
  assign n19954 = n19950 & n19953 ;
  assign n19955 = n19947 & n19954 ;
  assign n19956 = n19942 & n19955 ;
  assign n19957 = n19927 & n19956 ;
  assign n19958 = n2190 & n16222 ;
  assign n19959 = \s15_data_i[8]_pad  & n2190 ;
  assign n19960 = ~n2258 & n19959 ;
  assign n19961 = ~n19958 & ~n19960 ;
  assign n19962 = \s8_data_i[8]_pad  & n14923 ;
  assign n19963 = \s13_data_i[8]_pad  & n14904 ;
  assign n19964 = ~n19962 & ~n19963 ;
  assign n19965 = \s10_data_i[8]_pad  & n14892 ;
  assign n19966 = \s1_data_i[8]_pad  & n14609 ;
  assign n19967 = ~n19965 & ~n19966 ;
  assign n19968 = n19964 & n19967 ;
  assign n19969 = \s5_data_i[8]_pad  & n14757 ;
  assign n19970 = \s6_data_i[8]_pad  & n14745 ;
  assign n19971 = ~n19969 & ~n19970 ;
  assign n19972 = \s7_data_i[8]_pad  & n14740 ;
  assign n19973 = \s2_data_i[8]_pad  & n14911 ;
  assign n19974 = ~n19972 & ~n19973 ;
  assign n19975 = n19971 & n19974 ;
  assign n19976 = n19968 & n19975 ;
  assign n19977 = \s11_data_i[8]_pad  & n14896 ;
  assign n19978 = \s4_data_i[8]_pad  & n14919 ;
  assign n19979 = \s3_data_i[8]_pad  & n14801 ;
  assign n19980 = ~n19978 & ~n19979 ;
  assign n19981 = ~n19977 & n19980 ;
  assign n19982 = \s12_data_i[8]_pad  & n14900 ;
  assign n19983 = \s14_data_i[8]_pad  & n14915 ;
  assign n19984 = ~n19982 & ~n19983 ;
  assign n19985 = \s0_data_i[8]_pad  & n14603 ;
  assign n19986 = \s9_data_i[8]_pad  & n14927 ;
  assign n19987 = ~n19985 & ~n19986 ;
  assign n19988 = n19984 & n19987 ;
  assign n19989 = n19981 & n19988 ;
  assign n19990 = n19976 & n19989 ;
  assign n19991 = n19961 & n19990 ;
  assign n19992 = n2190 & n16259 ;
  assign n19993 = \s15_data_i[9]_pad  & n2190 ;
  assign n19994 = ~n2258 & n19993 ;
  assign n19995 = ~n19992 & ~n19994 ;
  assign n19996 = \s2_data_i[9]_pad  & n14911 ;
  assign n19997 = \s13_data_i[9]_pad  & n14904 ;
  assign n19998 = ~n19996 & ~n19997 ;
  assign n19999 = \s11_data_i[9]_pad  & n14896 ;
  assign n20000 = \s6_data_i[9]_pad  & n14745 ;
  assign n20001 = ~n19999 & ~n20000 ;
  assign n20002 = n19998 & n20001 ;
  assign n20003 = \s4_data_i[9]_pad  & n14919 ;
  assign n20004 = \s3_data_i[9]_pad  & n14801 ;
  assign n20005 = ~n20003 & ~n20004 ;
  assign n20006 = \s12_data_i[9]_pad  & n14900 ;
  assign n20007 = \s7_data_i[9]_pad  & n14740 ;
  assign n20008 = ~n20006 & ~n20007 ;
  assign n20009 = n20005 & n20008 ;
  assign n20010 = n20002 & n20009 ;
  assign n20011 = \s1_data_i[9]_pad  & n14609 ;
  assign n20012 = \s8_data_i[9]_pad  & n14923 ;
  assign n20013 = \s0_data_i[9]_pad  & n14603 ;
  assign n20014 = ~n20012 & ~n20013 ;
  assign n20015 = ~n20011 & n20014 ;
  assign n20016 = \s9_data_i[9]_pad  & n14927 ;
  assign n20017 = \s10_data_i[9]_pad  & n14892 ;
  assign n20018 = ~n20016 & ~n20017 ;
  assign n20019 = \s5_data_i[9]_pad  & n14757 ;
  assign n20020 = \s14_data_i[9]_pad  & n14915 ;
  assign n20021 = ~n20019 & ~n20020 ;
  assign n20022 = n20018 & n20021 ;
  assign n20023 = n20015 & n20022 ;
  assign n20024 = n20010 & n20023 ;
  assign n20025 = n19995 & n20024 ;
  assign n20026 = \s15_err_i_pad  & n18907 ;
  assign n20027 = ~n2258 & n20026 ;
  assign n20028 = \s14_err_i_pad  & n14915 ;
  assign n20029 = ~n14331 & n20028 ;
  assign n20030 = n14339 & n20029 ;
  assign n20031 = \s3_err_i_pad  & n14801 ;
  assign n20032 = ~n14451 & n20031 ;
  assign n20033 = n14459 & n20032 ;
  assign n20034 = ~n20030 & ~n20033 ;
  assign n20035 = \s13_err_i_pad  & n14904 ;
  assign n20036 = ~n14211 & n20035 ;
  assign n20037 = n14228 & n20036 ;
  assign n20038 = \s6_err_i_pad  & n14745 ;
  assign n20039 = ~n13627 & n20038 ;
  assign n20040 = n13635 & n20039 ;
  assign n20041 = ~n20037 & ~n20040 ;
  assign n20042 = n20034 & n20041 ;
  assign n20043 = \s0_err_i_pad  & n14603 ;
  assign n20044 = ~n14069 & n20043 ;
  assign n20045 = n14086 & n20044 ;
  assign n20046 = \s10_err_i_pad  & n14892 ;
  assign n20047 = ~n13928 & n20046 ;
  assign n20048 = n13921 & n20047 ;
  assign n20049 = ~n20045 & ~n20048 ;
  assign n20050 = \s9_err_i_pad  & n14927 ;
  assign n20051 = ~n13847 & n20050 ;
  assign n20052 = n13840 & n20051 ;
  assign n20053 = \s7_err_i_pad  & n14740 ;
  assign n20054 = ~n13697 & n20053 ;
  assign n20055 = n13714 & n20054 ;
  assign n20056 = ~n20052 & ~n20055 ;
  assign n20057 = n20049 & n20056 ;
  assign n20058 = n20042 & n20057 ;
  assign n20059 = \s12_err_i_pad  & n14900 ;
  assign n20060 = ~n14140 & n20059 ;
  assign n20061 = n14133 & n20060 ;
  assign n20062 = \s11_err_i_pad  & n14896 ;
  assign n20063 = ~n14009 & n20062 ;
  assign n20064 = n14034 & n20063 ;
  assign n20065 = \s4_err_i_pad  & n14919 ;
  assign n20066 = ~n13467 & n20065 ;
  assign n20067 = n13484 & n20066 ;
  assign n20068 = ~n20064 & ~n20067 ;
  assign n20069 = ~n20061 & n20068 ;
  assign n20070 = \s1_err_i_pad  & n14609 ;
  assign n20071 = ~n14271 & n20070 ;
  assign n20072 = n14279 & n20071 ;
  assign n20073 = \s2_err_i_pad  & n14911 ;
  assign n20074 = ~n14391 & n20073 ;
  assign n20075 = n14416 & n20074 ;
  assign n20076 = ~n20072 & ~n20075 ;
  assign n20077 = \s5_err_i_pad  & n14757 ;
  assign n20078 = ~n13547 & n20077 ;
  assign n20079 = n13540 & n20078 ;
  assign n20080 = \s8_err_i_pad  & n14923 ;
  assign n20081 = ~n13767 & n20080 ;
  assign n20082 = n13775 & n20081 ;
  assign n20083 = ~n20079 & ~n20082 ;
  assign n20084 = n20076 & n20083 ;
  assign n20085 = n20069 & n20084 ;
  assign n20086 = n20058 & n20085 ;
  assign n20087 = ~n20027 & n20086 ;
  assign n20088 = \s15_rty_i_pad  & n18907 ;
  assign n20089 = ~n2258 & n20088 ;
  assign n20090 = \s11_rty_i_pad  & n14896 ;
  assign n20091 = ~n14009 & n20090 ;
  assign n20092 = n14034 & n20091 ;
  assign n20093 = \s3_rty_i_pad  & n14801 ;
  assign n20094 = ~n14451 & n20093 ;
  assign n20095 = n14459 & n20094 ;
  assign n20096 = ~n20092 & ~n20095 ;
  assign n20097 = \s13_rty_i_pad  & n14904 ;
  assign n20098 = ~n14211 & n20097 ;
  assign n20099 = n14228 & n20098 ;
  assign n20100 = \s0_rty_i_pad  & n14603 ;
  assign n20101 = ~n14069 & n20100 ;
  assign n20102 = n14086 & n20101 ;
  assign n20103 = ~n20099 & ~n20102 ;
  assign n20104 = n20096 & n20103 ;
  assign n20105 = \s6_rty_i_pad  & n14745 ;
  assign n20106 = ~n13627 & n20105 ;
  assign n20107 = n13635 & n20106 ;
  assign n20108 = \s10_rty_i_pad  & n14892 ;
  assign n20109 = ~n13928 & n20108 ;
  assign n20110 = n13921 & n20109 ;
  assign n20111 = ~n20107 & ~n20110 ;
  assign n20112 = \s9_rty_i_pad  & n14927 ;
  assign n20113 = ~n13847 & n20112 ;
  assign n20114 = n13840 & n20113 ;
  assign n20115 = \s4_rty_i_pad  & n14919 ;
  assign n20116 = ~n13467 & n20115 ;
  assign n20117 = n13484 & n20116 ;
  assign n20118 = ~n20114 & ~n20117 ;
  assign n20119 = n20111 & n20118 ;
  assign n20120 = n20104 & n20119 ;
  assign n20121 = \s8_rty_i_pad  & n14923 ;
  assign n20122 = ~n13767 & n20121 ;
  assign n20123 = n13775 & n20122 ;
  assign n20124 = \s14_rty_i_pad  & n14915 ;
  assign n20125 = ~n14331 & n20124 ;
  assign n20126 = n14339 & n20125 ;
  assign n20127 = \s7_rty_i_pad  & n14740 ;
  assign n20128 = ~n13697 & n20127 ;
  assign n20129 = n13714 & n20128 ;
  assign n20130 = ~n20126 & ~n20129 ;
  assign n20131 = ~n20123 & n20130 ;
  assign n20132 = \s1_rty_i_pad  & n14609 ;
  assign n20133 = ~n14271 & n20132 ;
  assign n20134 = n14279 & n20133 ;
  assign n20135 = \s2_rty_i_pad  & n14911 ;
  assign n20136 = ~n14391 & n20135 ;
  assign n20137 = n14416 & n20136 ;
  assign n20138 = ~n20134 & ~n20137 ;
  assign n20139 = \s5_rty_i_pad  & n14757 ;
  assign n20140 = ~n13547 & n20139 ;
  assign n20141 = n13540 & n20140 ;
  assign n20142 = \s12_rty_i_pad  & n14900 ;
  assign n20143 = ~n14140 & n20142 ;
  assign n20144 = n14133 & n20143 ;
  assign n20145 = ~n20141 & ~n20144 ;
  assign n20146 = n20138 & n20145 ;
  assign n20147 = n20131 & n20146 ;
  assign n20148 = n20120 & n20147 ;
  assign n20149 = ~n20089 & n20148 ;
  assign n20150 = n1925 & n2197 ;
  assign n20151 = n1918 & n20150 ;
  assign n20152 = ~n13416 & n20151 ;
  assign n20153 = ~n15125 & n20152 ;
  assign n20154 = \s14_ack_i_pad  & n14939 ;
  assign n20155 = n14331 & n20154 ;
  assign n20156 = n14356 & n20155 ;
  assign n20157 = \s3_ack_i_pad  & n14950 ;
  assign n20158 = n14451 & n20157 ;
  assign n20159 = n14444 & n20158 ;
  assign n20160 = ~n20156 & ~n20159 ;
  assign n20161 = \s8_ack_i_pad  & n14717 ;
  assign n20162 = n13767 & n20161 ;
  assign n20163 = n13792 & n20162 ;
  assign n20164 = \s7_ack_i_pad  & n14958 ;
  assign n20165 = n13697 & n20164 ;
  assign n20166 = n13722 & n20165 ;
  assign n20167 = ~n20163 & ~n20166 ;
  assign n20168 = n20160 & n20167 ;
  assign n20169 = \s10_ack_i_pad  & n14931 ;
  assign n20170 = n13928 & n20169 ;
  assign n20171 = n13953 & n20170 ;
  assign n20172 = \s11_ack_i_pad  & n14735 ;
  assign n20173 = n14009 & n20172 ;
  assign n20174 = n14002 & n20173 ;
  assign n20175 = ~n20171 & ~n20174 ;
  assign n20176 = \s13_ack_i_pad  & n14731 ;
  assign n20177 = n14211 & n20176 ;
  assign n20178 = n14236 & n20177 ;
  assign n20179 = \s6_ack_i_pad  & n14723 ;
  assign n20180 = n13627 & n20179 ;
  assign n20181 = n13652 & n20180 ;
  assign n20182 = ~n20178 & ~n20181 ;
  assign n20183 = n20175 & n20182 ;
  assign n20184 = n20168 & n20183 ;
  assign n20185 = \s12_ack_i_pad  & n14935 ;
  assign n20186 = n14140 & n20185 ;
  assign n20187 = n14157 & n20186 ;
  assign n20188 = \s2_ack_i_pad  & n14946 ;
  assign n20189 = n14391 & n20188 ;
  assign n20190 = n14384 & n20189 ;
  assign n20191 = \s9_ack_i_pad  & n14713 ;
  assign n20192 = n13847 & n20191 ;
  assign n20193 = n13872 & n20192 ;
  assign n20194 = ~n20190 & ~n20193 ;
  assign n20195 = ~n20187 & n20194 ;
  assign n20196 = \s4_ack_i_pad  & n14727 ;
  assign n20197 = n13467 & n20196 ;
  assign n20198 = n13460 & n20197 ;
  assign n20199 = \s0_ack_i_pad  & n14616 ;
  assign n20200 = n14069 & n20199 ;
  assign n20201 = n14077 & n20200 ;
  assign n20202 = ~n20198 & ~n20201 ;
  assign n20203 = \s5_ack_i_pad  & n14954 ;
  assign n20204 = n13547 & n20203 ;
  assign n20205 = n13555 & n20204 ;
  assign n20206 = \s1_ack_i_pad  & n14622 ;
  assign n20207 = n14271 & n20206 ;
  assign n20208 = n14288 & n20207 ;
  assign n20209 = ~n20205 & ~n20208 ;
  assign n20210 = n20202 & n20209 ;
  assign n20211 = n20195 & n20210 ;
  assign n20212 = n20184 & n20211 ;
  assign n20213 = ~n20153 & n20212 ;
  assign n20214 = n2197 & n15192 ;
  assign n20215 = \s15_data_i[0]_pad  & n2197 ;
  assign n20216 = ~n2258 & n20215 ;
  assign n20217 = ~n20214 & ~n20216 ;
  assign n20218 = \s8_data_i[0]_pad  & n14717 ;
  assign n20219 = \s1_data_i[0]_pad  & n14622 ;
  assign n20220 = ~n20218 & ~n20219 ;
  assign n20221 = \s4_data_i[0]_pad  & n14727 ;
  assign n20222 = \s6_data_i[0]_pad  & n14723 ;
  assign n20223 = ~n20221 & ~n20222 ;
  assign n20224 = n20220 & n20223 ;
  assign n20225 = \s3_data_i[0]_pad  & n14950 ;
  assign n20226 = \s9_data_i[0]_pad  & n14713 ;
  assign n20227 = ~n20225 & ~n20226 ;
  assign n20228 = \s10_data_i[0]_pad  & n14931 ;
  assign n20229 = \s7_data_i[0]_pad  & n14958 ;
  assign n20230 = ~n20228 & ~n20229 ;
  assign n20231 = n20227 & n20230 ;
  assign n20232 = n20224 & n20231 ;
  assign n20233 = \s11_data_i[0]_pad  & n14735 ;
  assign n20234 = \s14_data_i[0]_pad  & n14939 ;
  assign n20235 = \s2_data_i[0]_pad  & n14946 ;
  assign n20236 = ~n20234 & ~n20235 ;
  assign n20237 = ~n20233 & n20236 ;
  assign n20238 = \s5_data_i[0]_pad  & n14954 ;
  assign n20239 = \s12_data_i[0]_pad  & n14935 ;
  assign n20240 = ~n20238 & ~n20239 ;
  assign n20241 = \s13_data_i[0]_pad  & n14731 ;
  assign n20242 = \s0_data_i[0]_pad  & n14616 ;
  assign n20243 = ~n20241 & ~n20242 ;
  assign n20244 = n20240 & n20243 ;
  assign n20245 = n20237 & n20244 ;
  assign n20246 = n20232 & n20245 ;
  assign n20247 = n20217 & n20246 ;
  assign n20248 = n2197 & n15229 ;
  assign n20249 = \s15_data_i[10]_pad  & n2197 ;
  assign n20250 = ~n2258 & n20249 ;
  assign n20251 = ~n20248 & ~n20250 ;
  assign n20252 = \s8_data_i[10]_pad  & n14717 ;
  assign n20253 = \s1_data_i[10]_pad  & n14622 ;
  assign n20254 = ~n20252 & ~n20253 ;
  assign n20255 = \s4_data_i[10]_pad  & n14727 ;
  assign n20256 = \s6_data_i[10]_pad  & n14723 ;
  assign n20257 = ~n20255 & ~n20256 ;
  assign n20258 = n20254 & n20257 ;
  assign n20259 = \s3_data_i[10]_pad  & n14950 ;
  assign n20260 = \s9_data_i[10]_pad  & n14713 ;
  assign n20261 = ~n20259 & ~n20260 ;
  assign n20262 = \s10_data_i[10]_pad  & n14931 ;
  assign n20263 = \s7_data_i[10]_pad  & n14958 ;
  assign n20264 = ~n20262 & ~n20263 ;
  assign n20265 = n20261 & n20264 ;
  assign n20266 = n20258 & n20265 ;
  assign n20267 = \s11_data_i[10]_pad  & n14735 ;
  assign n20268 = \s14_data_i[10]_pad  & n14939 ;
  assign n20269 = \s2_data_i[10]_pad  & n14946 ;
  assign n20270 = ~n20268 & ~n20269 ;
  assign n20271 = ~n20267 & n20270 ;
  assign n20272 = \s5_data_i[10]_pad  & n14954 ;
  assign n20273 = \s12_data_i[10]_pad  & n14935 ;
  assign n20274 = ~n20272 & ~n20273 ;
  assign n20275 = \s13_data_i[10]_pad  & n14731 ;
  assign n20276 = \s0_data_i[10]_pad  & n14616 ;
  assign n20277 = ~n20275 & ~n20276 ;
  assign n20278 = n20274 & n20277 ;
  assign n20279 = n20271 & n20278 ;
  assign n20280 = n20266 & n20279 ;
  assign n20281 = n20251 & n20280 ;
  assign n20282 = n2197 & n15266 ;
  assign n20283 = \s15_data_i[11]_pad  & n2197 ;
  assign n20284 = ~n2258 & n20283 ;
  assign n20285 = ~n20282 & ~n20284 ;
  assign n20286 = \s8_data_i[11]_pad  & n14717 ;
  assign n20287 = \s1_data_i[11]_pad  & n14622 ;
  assign n20288 = ~n20286 & ~n20287 ;
  assign n20289 = \s4_data_i[11]_pad  & n14727 ;
  assign n20290 = \s6_data_i[11]_pad  & n14723 ;
  assign n20291 = ~n20289 & ~n20290 ;
  assign n20292 = n20288 & n20291 ;
  assign n20293 = \s3_data_i[11]_pad  & n14950 ;
  assign n20294 = \s9_data_i[11]_pad  & n14713 ;
  assign n20295 = ~n20293 & ~n20294 ;
  assign n20296 = \s10_data_i[11]_pad  & n14931 ;
  assign n20297 = \s7_data_i[11]_pad  & n14958 ;
  assign n20298 = ~n20296 & ~n20297 ;
  assign n20299 = n20295 & n20298 ;
  assign n20300 = n20292 & n20299 ;
  assign n20301 = \s11_data_i[11]_pad  & n14735 ;
  assign n20302 = \s14_data_i[11]_pad  & n14939 ;
  assign n20303 = \s2_data_i[11]_pad  & n14946 ;
  assign n20304 = ~n20302 & ~n20303 ;
  assign n20305 = ~n20301 & n20304 ;
  assign n20306 = \s5_data_i[11]_pad  & n14954 ;
  assign n20307 = \s12_data_i[11]_pad  & n14935 ;
  assign n20308 = ~n20306 & ~n20307 ;
  assign n20309 = \s13_data_i[11]_pad  & n14731 ;
  assign n20310 = \s0_data_i[11]_pad  & n14616 ;
  assign n20311 = ~n20309 & ~n20310 ;
  assign n20312 = n20308 & n20311 ;
  assign n20313 = n20305 & n20312 ;
  assign n20314 = n20300 & n20313 ;
  assign n20315 = n20285 & n20314 ;
  assign n20316 = n2197 & n15303 ;
  assign n20317 = \s15_data_i[12]_pad  & n2197 ;
  assign n20318 = ~n2258 & n20317 ;
  assign n20319 = ~n20316 & ~n20318 ;
  assign n20320 = \s8_data_i[12]_pad  & n14717 ;
  assign n20321 = \s1_data_i[12]_pad  & n14622 ;
  assign n20322 = ~n20320 & ~n20321 ;
  assign n20323 = \s4_data_i[12]_pad  & n14727 ;
  assign n20324 = \s6_data_i[12]_pad  & n14723 ;
  assign n20325 = ~n20323 & ~n20324 ;
  assign n20326 = n20322 & n20325 ;
  assign n20327 = \s3_data_i[12]_pad  & n14950 ;
  assign n20328 = \s9_data_i[12]_pad  & n14713 ;
  assign n20329 = ~n20327 & ~n20328 ;
  assign n20330 = \s10_data_i[12]_pad  & n14931 ;
  assign n20331 = \s7_data_i[12]_pad  & n14958 ;
  assign n20332 = ~n20330 & ~n20331 ;
  assign n20333 = n20329 & n20332 ;
  assign n20334 = n20326 & n20333 ;
  assign n20335 = \s11_data_i[12]_pad  & n14735 ;
  assign n20336 = \s14_data_i[12]_pad  & n14939 ;
  assign n20337 = \s2_data_i[12]_pad  & n14946 ;
  assign n20338 = ~n20336 & ~n20337 ;
  assign n20339 = ~n20335 & n20338 ;
  assign n20340 = \s5_data_i[12]_pad  & n14954 ;
  assign n20341 = \s12_data_i[12]_pad  & n14935 ;
  assign n20342 = ~n20340 & ~n20341 ;
  assign n20343 = \s13_data_i[12]_pad  & n14731 ;
  assign n20344 = \s0_data_i[12]_pad  & n14616 ;
  assign n20345 = ~n20343 & ~n20344 ;
  assign n20346 = n20342 & n20345 ;
  assign n20347 = n20339 & n20346 ;
  assign n20348 = n20334 & n20347 ;
  assign n20349 = n20319 & n20348 ;
  assign n20350 = n2197 & n15340 ;
  assign n20351 = \s15_data_i[13]_pad  & n2197 ;
  assign n20352 = ~n2258 & n20351 ;
  assign n20353 = ~n20350 & ~n20352 ;
  assign n20354 = \s8_data_i[13]_pad  & n14717 ;
  assign n20355 = \s1_data_i[13]_pad  & n14622 ;
  assign n20356 = ~n20354 & ~n20355 ;
  assign n20357 = \s4_data_i[13]_pad  & n14727 ;
  assign n20358 = \s6_data_i[13]_pad  & n14723 ;
  assign n20359 = ~n20357 & ~n20358 ;
  assign n20360 = n20356 & n20359 ;
  assign n20361 = \s3_data_i[13]_pad  & n14950 ;
  assign n20362 = \s9_data_i[13]_pad  & n14713 ;
  assign n20363 = ~n20361 & ~n20362 ;
  assign n20364 = \s10_data_i[13]_pad  & n14931 ;
  assign n20365 = \s7_data_i[13]_pad  & n14958 ;
  assign n20366 = ~n20364 & ~n20365 ;
  assign n20367 = n20363 & n20366 ;
  assign n20368 = n20360 & n20367 ;
  assign n20369 = \s11_data_i[13]_pad  & n14735 ;
  assign n20370 = \s14_data_i[13]_pad  & n14939 ;
  assign n20371 = \s2_data_i[13]_pad  & n14946 ;
  assign n20372 = ~n20370 & ~n20371 ;
  assign n20373 = ~n20369 & n20372 ;
  assign n20374 = \s5_data_i[13]_pad  & n14954 ;
  assign n20375 = \s12_data_i[13]_pad  & n14935 ;
  assign n20376 = ~n20374 & ~n20375 ;
  assign n20377 = \s13_data_i[13]_pad  & n14731 ;
  assign n20378 = \s0_data_i[13]_pad  & n14616 ;
  assign n20379 = ~n20377 & ~n20378 ;
  assign n20380 = n20376 & n20379 ;
  assign n20381 = n20373 & n20380 ;
  assign n20382 = n20368 & n20381 ;
  assign n20383 = n20353 & n20382 ;
  assign n20384 = n2197 & n15377 ;
  assign n20385 = \s15_data_i[14]_pad  & n2197 ;
  assign n20386 = ~n2258 & n20385 ;
  assign n20387 = ~n20384 & ~n20386 ;
  assign n20388 = \s8_data_i[14]_pad  & n14717 ;
  assign n20389 = \s1_data_i[14]_pad  & n14622 ;
  assign n20390 = ~n20388 & ~n20389 ;
  assign n20391 = \s10_data_i[14]_pad  & n14931 ;
  assign n20392 = \s0_data_i[14]_pad  & n14616 ;
  assign n20393 = ~n20391 & ~n20392 ;
  assign n20394 = n20390 & n20393 ;
  assign n20395 = \s3_data_i[14]_pad  & n14950 ;
  assign n20396 = \s6_data_i[14]_pad  & n14723 ;
  assign n20397 = ~n20395 & ~n20396 ;
  assign n20398 = \s7_data_i[14]_pad  & n14958 ;
  assign n20399 = \s4_data_i[14]_pad  & n14727 ;
  assign n20400 = ~n20398 & ~n20399 ;
  assign n20401 = n20397 & n20400 ;
  assign n20402 = n20394 & n20401 ;
  assign n20403 = \s11_data_i[14]_pad  & n14735 ;
  assign n20404 = \s14_data_i[14]_pad  & n14939 ;
  assign n20405 = \s2_data_i[14]_pad  & n14946 ;
  assign n20406 = ~n20404 & ~n20405 ;
  assign n20407 = ~n20403 & n20406 ;
  assign n20408 = \s5_data_i[14]_pad  & n14954 ;
  assign n20409 = \s12_data_i[14]_pad  & n14935 ;
  assign n20410 = ~n20408 & ~n20409 ;
  assign n20411 = \s13_data_i[14]_pad  & n14731 ;
  assign n20412 = \s9_data_i[14]_pad  & n14713 ;
  assign n20413 = ~n20411 & ~n20412 ;
  assign n20414 = n20410 & n20413 ;
  assign n20415 = n20407 & n20414 ;
  assign n20416 = n20402 & n20415 ;
  assign n20417 = n20387 & n20416 ;
  assign n20418 = n2197 & n15414 ;
  assign n20419 = \s15_data_i[15]_pad  & n2197 ;
  assign n20420 = ~n2258 & n20419 ;
  assign n20421 = ~n20418 & ~n20420 ;
  assign n20422 = \s8_data_i[15]_pad  & n14717 ;
  assign n20423 = \s1_data_i[15]_pad  & n14622 ;
  assign n20424 = ~n20422 & ~n20423 ;
  assign n20425 = \s4_data_i[15]_pad  & n14727 ;
  assign n20426 = \s6_data_i[15]_pad  & n14723 ;
  assign n20427 = ~n20425 & ~n20426 ;
  assign n20428 = n20424 & n20427 ;
  assign n20429 = \s3_data_i[15]_pad  & n14950 ;
  assign n20430 = \s9_data_i[15]_pad  & n14713 ;
  assign n20431 = ~n20429 & ~n20430 ;
  assign n20432 = \s10_data_i[15]_pad  & n14931 ;
  assign n20433 = \s7_data_i[15]_pad  & n14958 ;
  assign n20434 = ~n20432 & ~n20433 ;
  assign n20435 = n20431 & n20434 ;
  assign n20436 = n20428 & n20435 ;
  assign n20437 = \s11_data_i[15]_pad  & n14735 ;
  assign n20438 = \s14_data_i[15]_pad  & n14939 ;
  assign n20439 = \s2_data_i[15]_pad  & n14946 ;
  assign n20440 = ~n20438 & ~n20439 ;
  assign n20441 = ~n20437 & n20440 ;
  assign n20442 = \s5_data_i[15]_pad  & n14954 ;
  assign n20443 = \s12_data_i[15]_pad  & n14935 ;
  assign n20444 = ~n20442 & ~n20443 ;
  assign n20445 = \s13_data_i[15]_pad  & n14731 ;
  assign n20446 = \s0_data_i[15]_pad  & n14616 ;
  assign n20447 = ~n20445 & ~n20446 ;
  assign n20448 = n20444 & n20447 ;
  assign n20449 = n20441 & n20448 ;
  assign n20450 = n20436 & n20449 ;
  assign n20451 = n20421 & n20450 ;
  assign n20452 = \s15_data_i[16]_pad  & n2197 ;
  assign n20453 = ~n2258 & n20452 ;
  assign n20454 = \s8_data_i[16]_pad  & n14717 ;
  assign n20455 = \s1_data_i[16]_pad  & n14622 ;
  assign n20456 = ~n20454 & ~n20455 ;
  assign n20457 = \s4_data_i[16]_pad  & n14727 ;
  assign n20458 = \s6_data_i[16]_pad  & n14723 ;
  assign n20459 = ~n20457 & ~n20458 ;
  assign n20460 = n20456 & n20459 ;
  assign n20461 = \s3_data_i[16]_pad  & n14950 ;
  assign n20462 = \s9_data_i[16]_pad  & n14713 ;
  assign n20463 = ~n20461 & ~n20462 ;
  assign n20464 = \s10_data_i[16]_pad  & n14931 ;
  assign n20465 = \s7_data_i[16]_pad  & n14958 ;
  assign n20466 = ~n20464 & ~n20465 ;
  assign n20467 = n20463 & n20466 ;
  assign n20468 = n20460 & n20467 ;
  assign n20469 = \s11_data_i[16]_pad  & n14735 ;
  assign n20470 = \s14_data_i[16]_pad  & n14939 ;
  assign n20471 = \s2_data_i[16]_pad  & n14946 ;
  assign n20472 = ~n20470 & ~n20471 ;
  assign n20473 = ~n20469 & n20472 ;
  assign n20474 = \s5_data_i[16]_pad  & n14954 ;
  assign n20475 = \s12_data_i[16]_pad  & n14935 ;
  assign n20476 = ~n20474 & ~n20475 ;
  assign n20477 = \s13_data_i[16]_pad  & n14731 ;
  assign n20478 = \s0_data_i[16]_pad  & n14616 ;
  assign n20479 = ~n20477 & ~n20478 ;
  assign n20480 = n20476 & n20479 ;
  assign n20481 = n20473 & n20480 ;
  assign n20482 = n20468 & n20481 ;
  assign n20483 = ~n20453 & n20482 ;
  assign n20484 = \s15_data_i[17]_pad  & n2197 ;
  assign n20485 = ~n2258 & n20484 ;
  assign n20486 = \s8_data_i[17]_pad  & n14717 ;
  assign n20487 = \s1_data_i[17]_pad  & n14622 ;
  assign n20488 = ~n20486 & ~n20487 ;
  assign n20489 = \s4_data_i[17]_pad  & n14727 ;
  assign n20490 = \s6_data_i[17]_pad  & n14723 ;
  assign n20491 = ~n20489 & ~n20490 ;
  assign n20492 = n20488 & n20491 ;
  assign n20493 = \s3_data_i[17]_pad  & n14950 ;
  assign n20494 = \s9_data_i[17]_pad  & n14713 ;
  assign n20495 = ~n20493 & ~n20494 ;
  assign n20496 = \s10_data_i[17]_pad  & n14931 ;
  assign n20497 = \s7_data_i[17]_pad  & n14958 ;
  assign n20498 = ~n20496 & ~n20497 ;
  assign n20499 = n20495 & n20498 ;
  assign n20500 = n20492 & n20499 ;
  assign n20501 = \s11_data_i[17]_pad  & n14735 ;
  assign n20502 = \s14_data_i[17]_pad  & n14939 ;
  assign n20503 = \s2_data_i[17]_pad  & n14946 ;
  assign n20504 = ~n20502 & ~n20503 ;
  assign n20505 = ~n20501 & n20504 ;
  assign n20506 = \s5_data_i[17]_pad  & n14954 ;
  assign n20507 = \s12_data_i[17]_pad  & n14935 ;
  assign n20508 = ~n20506 & ~n20507 ;
  assign n20509 = \s13_data_i[17]_pad  & n14731 ;
  assign n20510 = \s0_data_i[17]_pad  & n14616 ;
  assign n20511 = ~n20509 & ~n20510 ;
  assign n20512 = n20508 & n20511 ;
  assign n20513 = n20505 & n20512 ;
  assign n20514 = n20500 & n20513 ;
  assign n20515 = ~n20485 & n20514 ;
  assign n20516 = \s15_data_i[18]_pad  & n2197 ;
  assign n20517 = ~n2258 & n20516 ;
  assign n20518 = \s12_data_i[18]_pad  & n14935 ;
  assign n20519 = \s1_data_i[18]_pad  & n14622 ;
  assign n20520 = ~n20518 & ~n20519 ;
  assign n20521 = \s4_data_i[18]_pad  & n14727 ;
  assign n20522 = \s6_data_i[18]_pad  & n14723 ;
  assign n20523 = ~n20521 & ~n20522 ;
  assign n20524 = n20520 & n20523 ;
  assign n20525 = \s3_data_i[18]_pad  & n14950 ;
  assign n20526 = \s9_data_i[18]_pad  & n14713 ;
  assign n20527 = ~n20525 & ~n20526 ;
  assign n20528 = \s10_data_i[18]_pad  & n14931 ;
  assign n20529 = \s7_data_i[18]_pad  & n14958 ;
  assign n20530 = ~n20528 & ~n20529 ;
  assign n20531 = n20527 & n20530 ;
  assign n20532 = n20524 & n20531 ;
  assign n20533 = \s14_data_i[18]_pad  & n14939 ;
  assign n20534 = \s11_data_i[18]_pad  & n14735 ;
  assign n20535 = \s2_data_i[18]_pad  & n14946 ;
  assign n20536 = ~n20534 & ~n20535 ;
  assign n20537 = ~n20533 & n20536 ;
  assign n20538 = \s5_data_i[18]_pad  & n14954 ;
  assign n20539 = \s8_data_i[18]_pad  & n14717 ;
  assign n20540 = ~n20538 & ~n20539 ;
  assign n20541 = \s13_data_i[18]_pad  & n14731 ;
  assign n20542 = \s0_data_i[18]_pad  & n14616 ;
  assign n20543 = ~n20541 & ~n20542 ;
  assign n20544 = n20540 & n20543 ;
  assign n20545 = n20537 & n20544 ;
  assign n20546 = n20532 & n20545 ;
  assign n20547 = ~n20517 & n20546 ;
  assign n20548 = \s15_data_i[19]_pad  & n2197 ;
  assign n20549 = ~n2258 & n20548 ;
  assign n20550 = \s8_data_i[19]_pad  & n14717 ;
  assign n20551 = \s1_data_i[19]_pad  & n14622 ;
  assign n20552 = ~n20550 & ~n20551 ;
  assign n20553 = \s4_data_i[19]_pad  & n14727 ;
  assign n20554 = \s6_data_i[19]_pad  & n14723 ;
  assign n20555 = ~n20553 & ~n20554 ;
  assign n20556 = n20552 & n20555 ;
  assign n20557 = \s3_data_i[19]_pad  & n14950 ;
  assign n20558 = \s9_data_i[19]_pad  & n14713 ;
  assign n20559 = ~n20557 & ~n20558 ;
  assign n20560 = \s10_data_i[19]_pad  & n14931 ;
  assign n20561 = \s7_data_i[19]_pad  & n14958 ;
  assign n20562 = ~n20560 & ~n20561 ;
  assign n20563 = n20559 & n20562 ;
  assign n20564 = n20556 & n20563 ;
  assign n20565 = \s11_data_i[19]_pad  & n14735 ;
  assign n20566 = \s14_data_i[19]_pad  & n14939 ;
  assign n20567 = \s2_data_i[19]_pad  & n14946 ;
  assign n20568 = ~n20566 & ~n20567 ;
  assign n20569 = ~n20565 & n20568 ;
  assign n20570 = \s5_data_i[19]_pad  & n14954 ;
  assign n20571 = \s12_data_i[19]_pad  & n14935 ;
  assign n20572 = ~n20570 & ~n20571 ;
  assign n20573 = \s13_data_i[19]_pad  & n14731 ;
  assign n20574 = \s0_data_i[19]_pad  & n14616 ;
  assign n20575 = ~n20573 & ~n20574 ;
  assign n20576 = n20572 & n20575 ;
  assign n20577 = n20569 & n20576 ;
  assign n20578 = n20564 & n20577 ;
  assign n20579 = ~n20549 & n20578 ;
  assign n20580 = n2197 & n15579 ;
  assign n20581 = \s15_data_i[1]_pad  & n2197 ;
  assign n20582 = ~n2258 & n20581 ;
  assign n20583 = ~n20580 & ~n20582 ;
  assign n20584 = \s8_data_i[1]_pad  & n14717 ;
  assign n20585 = \s1_data_i[1]_pad  & n14622 ;
  assign n20586 = ~n20584 & ~n20585 ;
  assign n20587 = \s4_data_i[1]_pad  & n14727 ;
  assign n20588 = \s6_data_i[1]_pad  & n14723 ;
  assign n20589 = ~n20587 & ~n20588 ;
  assign n20590 = n20586 & n20589 ;
  assign n20591 = \s3_data_i[1]_pad  & n14950 ;
  assign n20592 = \s9_data_i[1]_pad  & n14713 ;
  assign n20593 = ~n20591 & ~n20592 ;
  assign n20594 = \s10_data_i[1]_pad  & n14931 ;
  assign n20595 = \s7_data_i[1]_pad  & n14958 ;
  assign n20596 = ~n20594 & ~n20595 ;
  assign n20597 = n20593 & n20596 ;
  assign n20598 = n20590 & n20597 ;
  assign n20599 = \s11_data_i[1]_pad  & n14735 ;
  assign n20600 = \s14_data_i[1]_pad  & n14939 ;
  assign n20601 = \s2_data_i[1]_pad  & n14946 ;
  assign n20602 = ~n20600 & ~n20601 ;
  assign n20603 = ~n20599 & n20602 ;
  assign n20604 = \s5_data_i[1]_pad  & n14954 ;
  assign n20605 = \s12_data_i[1]_pad  & n14935 ;
  assign n20606 = ~n20604 & ~n20605 ;
  assign n20607 = \s13_data_i[1]_pad  & n14731 ;
  assign n20608 = \s0_data_i[1]_pad  & n14616 ;
  assign n20609 = ~n20607 & ~n20608 ;
  assign n20610 = n20606 & n20609 ;
  assign n20611 = n20603 & n20610 ;
  assign n20612 = n20598 & n20611 ;
  assign n20613 = n20583 & n20612 ;
  assign n20614 = \s15_data_i[20]_pad  & n2197 ;
  assign n20615 = ~n2258 & n20614 ;
  assign n20616 = \s8_data_i[20]_pad  & n14717 ;
  assign n20617 = \s1_data_i[20]_pad  & n14622 ;
  assign n20618 = ~n20616 & ~n20617 ;
  assign n20619 = \s4_data_i[20]_pad  & n14727 ;
  assign n20620 = \s6_data_i[20]_pad  & n14723 ;
  assign n20621 = ~n20619 & ~n20620 ;
  assign n20622 = n20618 & n20621 ;
  assign n20623 = \s3_data_i[20]_pad  & n14950 ;
  assign n20624 = \s9_data_i[20]_pad  & n14713 ;
  assign n20625 = ~n20623 & ~n20624 ;
  assign n20626 = \s10_data_i[20]_pad  & n14931 ;
  assign n20627 = \s7_data_i[20]_pad  & n14958 ;
  assign n20628 = ~n20626 & ~n20627 ;
  assign n20629 = n20625 & n20628 ;
  assign n20630 = n20622 & n20629 ;
  assign n20631 = \s11_data_i[20]_pad  & n14735 ;
  assign n20632 = \s14_data_i[20]_pad  & n14939 ;
  assign n20633 = \s2_data_i[20]_pad  & n14946 ;
  assign n20634 = ~n20632 & ~n20633 ;
  assign n20635 = ~n20631 & n20634 ;
  assign n20636 = \s5_data_i[20]_pad  & n14954 ;
  assign n20637 = \s12_data_i[20]_pad  & n14935 ;
  assign n20638 = ~n20636 & ~n20637 ;
  assign n20639 = \s13_data_i[20]_pad  & n14731 ;
  assign n20640 = \s0_data_i[20]_pad  & n14616 ;
  assign n20641 = ~n20639 & ~n20640 ;
  assign n20642 = n20638 & n20641 ;
  assign n20643 = n20635 & n20642 ;
  assign n20644 = n20630 & n20643 ;
  assign n20645 = ~n20615 & n20644 ;
  assign n20646 = \s15_data_i[21]_pad  & n2197 ;
  assign n20647 = ~n2258 & n20646 ;
  assign n20648 = \s8_data_i[21]_pad  & n14717 ;
  assign n20649 = \s1_data_i[21]_pad  & n14622 ;
  assign n20650 = ~n20648 & ~n20649 ;
  assign n20651 = \s4_data_i[21]_pad  & n14727 ;
  assign n20652 = \s6_data_i[21]_pad  & n14723 ;
  assign n20653 = ~n20651 & ~n20652 ;
  assign n20654 = n20650 & n20653 ;
  assign n20655 = \s3_data_i[21]_pad  & n14950 ;
  assign n20656 = \s9_data_i[21]_pad  & n14713 ;
  assign n20657 = ~n20655 & ~n20656 ;
  assign n20658 = \s10_data_i[21]_pad  & n14931 ;
  assign n20659 = \s7_data_i[21]_pad  & n14958 ;
  assign n20660 = ~n20658 & ~n20659 ;
  assign n20661 = n20657 & n20660 ;
  assign n20662 = n20654 & n20661 ;
  assign n20663 = \s11_data_i[21]_pad  & n14735 ;
  assign n20664 = \s14_data_i[21]_pad  & n14939 ;
  assign n20665 = \s2_data_i[21]_pad  & n14946 ;
  assign n20666 = ~n20664 & ~n20665 ;
  assign n20667 = ~n20663 & n20666 ;
  assign n20668 = \s5_data_i[21]_pad  & n14954 ;
  assign n20669 = \s12_data_i[21]_pad  & n14935 ;
  assign n20670 = ~n20668 & ~n20669 ;
  assign n20671 = \s13_data_i[21]_pad  & n14731 ;
  assign n20672 = \s0_data_i[21]_pad  & n14616 ;
  assign n20673 = ~n20671 & ~n20672 ;
  assign n20674 = n20670 & n20673 ;
  assign n20675 = n20667 & n20674 ;
  assign n20676 = n20662 & n20675 ;
  assign n20677 = ~n20647 & n20676 ;
  assign n20678 = \s15_data_i[22]_pad  & n2197 ;
  assign n20679 = ~n2258 & n20678 ;
  assign n20680 = \s8_data_i[22]_pad  & n14717 ;
  assign n20681 = \s1_data_i[22]_pad  & n14622 ;
  assign n20682 = ~n20680 & ~n20681 ;
  assign n20683 = \s4_data_i[22]_pad  & n14727 ;
  assign n20684 = \s6_data_i[22]_pad  & n14723 ;
  assign n20685 = ~n20683 & ~n20684 ;
  assign n20686 = n20682 & n20685 ;
  assign n20687 = \s3_data_i[22]_pad  & n14950 ;
  assign n20688 = \s9_data_i[22]_pad  & n14713 ;
  assign n20689 = ~n20687 & ~n20688 ;
  assign n20690 = \s10_data_i[22]_pad  & n14931 ;
  assign n20691 = \s7_data_i[22]_pad  & n14958 ;
  assign n20692 = ~n20690 & ~n20691 ;
  assign n20693 = n20689 & n20692 ;
  assign n20694 = n20686 & n20693 ;
  assign n20695 = \s11_data_i[22]_pad  & n14735 ;
  assign n20696 = \s14_data_i[22]_pad  & n14939 ;
  assign n20697 = \s2_data_i[22]_pad  & n14946 ;
  assign n20698 = ~n20696 & ~n20697 ;
  assign n20699 = ~n20695 & n20698 ;
  assign n20700 = \s5_data_i[22]_pad  & n14954 ;
  assign n20701 = \s12_data_i[22]_pad  & n14935 ;
  assign n20702 = ~n20700 & ~n20701 ;
  assign n20703 = \s13_data_i[22]_pad  & n14731 ;
  assign n20704 = \s0_data_i[22]_pad  & n14616 ;
  assign n20705 = ~n20703 & ~n20704 ;
  assign n20706 = n20702 & n20705 ;
  assign n20707 = n20699 & n20706 ;
  assign n20708 = n20694 & n20707 ;
  assign n20709 = ~n20679 & n20708 ;
  assign n20710 = \s15_data_i[23]_pad  & n2197 ;
  assign n20711 = ~n2258 & n20710 ;
  assign n20712 = \s8_data_i[23]_pad  & n14717 ;
  assign n20713 = \s1_data_i[23]_pad  & n14622 ;
  assign n20714 = ~n20712 & ~n20713 ;
  assign n20715 = \s4_data_i[23]_pad  & n14727 ;
  assign n20716 = \s6_data_i[23]_pad  & n14723 ;
  assign n20717 = ~n20715 & ~n20716 ;
  assign n20718 = n20714 & n20717 ;
  assign n20719 = \s3_data_i[23]_pad  & n14950 ;
  assign n20720 = \s9_data_i[23]_pad  & n14713 ;
  assign n20721 = ~n20719 & ~n20720 ;
  assign n20722 = \s10_data_i[23]_pad  & n14931 ;
  assign n20723 = \s7_data_i[23]_pad  & n14958 ;
  assign n20724 = ~n20722 & ~n20723 ;
  assign n20725 = n20721 & n20724 ;
  assign n20726 = n20718 & n20725 ;
  assign n20727 = \s11_data_i[23]_pad  & n14735 ;
  assign n20728 = \s14_data_i[23]_pad  & n14939 ;
  assign n20729 = \s2_data_i[23]_pad  & n14946 ;
  assign n20730 = ~n20728 & ~n20729 ;
  assign n20731 = ~n20727 & n20730 ;
  assign n20732 = \s5_data_i[23]_pad  & n14954 ;
  assign n20733 = \s12_data_i[23]_pad  & n14935 ;
  assign n20734 = ~n20732 & ~n20733 ;
  assign n20735 = \s13_data_i[23]_pad  & n14731 ;
  assign n20736 = \s0_data_i[23]_pad  & n14616 ;
  assign n20737 = ~n20735 & ~n20736 ;
  assign n20738 = n20734 & n20737 ;
  assign n20739 = n20731 & n20738 ;
  assign n20740 = n20726 & n20739 ;
  assign n20741 = ~n20711 & n20740 ;
  assign n20742 = \s15_data_i[24]_pad  & n2197 ;
  assign n20743 = ~n2258 & n20742 ;
  assign n20744 = \s8_data_i[24]_pad  & n14717 ;
  assign n20745 = \s1_data_i[24]_pad  & n14622 ;
  assign n20746 = ~n20744 & ~n20745 ;
  assign n20747 = \s4_data_i[24]_pad  & n14727 ;
  assign n20748 = \s6_data_i[24]_pad  & n14723 ;
  assign n20749 = ~n20747 & ~n20748 ;
  assign n20750 = n20746 & n20749 ;
  assign n20751 = \s3_data_i[24]_pad  & n14950 ;
  assign n20752 = \s9_data_i[24]_pad  & n14713 ;
  assign n20753 = ~n20751 & ~n20752 ;
  assign n20754 = \s10_data_i[24]_pad  & n14931 ;
  assign n20755 = \s7_data_i[24]_pad  & n14958 ;
  assign n20756 = ~n20754 & ~n20755 ;
  assign n20757 = n20753 & n20756 ;
  assign n20758 = n20750 & n20757 ;
  assign n20759 = \s11_data_i[24]_pad  & n14735 ;
  assign n20760 = \s14_data_i[24]_pad  & n14939 ;
  assign n20761 = \s2_data_i[24]_pad  & n14946 ;
  assign n20762 = ~n20760 & ~n20761 ;
  assign n20763 = ~n20759 & n20762 ;
  assign n20764 = \s5_data_i[24]_pad  & n14954 ;
  assign n20765 = \s12_data_i[24]_pad  & n14935 ;
  assign n20766 = ~n20764 & ~n20765 ;
  assign n20767 = \s13_data_i[24]_pad  & n14731 ;
  assign n20768 = \s0_data_i[24]_pad  & n14616 ;
  assign n20769 = ~n20767 & ~n20768 ;
  assign n20770 = n20766 & n20769 ;
  assign n20771 = n20763 & n20770 ;
  assign n20772 = n20758 & n20771 ;
  assign n20773 = ~n20743 & n20772 ;
  assign n20774 = \s15_data_i[25]_pad  & n2197 ;
  assign n20775 = ~n2258 & n20774 ;
  assign n20776 = \s8_data_i[25]_pad  & n14717 ;
  assign n20777 = \s1_data_i[25]_pad  & n14622 ;
  assign n20778 = ~n20776 & ~n20777 ;
  assign n20779 = \s4_data_i[25]_pad  & n14727 ;
  assign n20780 = \s6_data_i[25]_pad  & n14723 ;
  assign n20781 = ~n20779 & ~n20780 ;
  assign n20782 = n20778 & n20781 ;
  assign n20783 = \s3_data_i[25]_pad  & n14950 ;
  assign n20784 = \s9_data_i[25]_pad  & n14713 ;
  assign n20785 = ~n20783 & ~n20784 ;
  assign n20786 = \s10_data_i[25]_pad  & n14931 ;
  assign n20787 = \s7_data_i[25]_pad  & n14958 ;
  assign n20788 = ~n20786 & ~n20787 ;
  assign n20789 = n20785 & n20788 ;
  assign n20790 = n20782 & n20789 ;
  assign n20791 = \s11_data_i[25]_pad  & n14735 ;
  assign n20792 = \s14_data_i[25]_pad  & n14939 ;
  assign n20793 = \s2_data_i[25]_pad  & n14946 ;
  assign n20794 = ~n20792 & ~n20793 ;
  assign n20795 = ~n20791 & n20794 ;
  assign n20796 = \s5_data_i[25]_pad  & n14954 ;
  assign n20797 = \s12_data_i[25]_pad  & n14935 ;
  assign n20798 = ~n20796 & ~n20797 ;
  assign n20799 = \s13_data_i[25]_pad  & n14731 ;
  assign n20800 = \s0_data_i[25]_pad  & n14616 ;
  assign n20801 = ~n20799 & ~n20800 ;
  assign n20802 = n20798 & n20801 ;
  assign n20803 = n20795 & n20802 ;
  assign n20804 = n20790 & n20803 ;
  assign n20805 = ~n20775 & n20804 ;
  assign n20806 = \s15_data_i[26]_pad  & n2197 ;
  assign n20807 = ~n2258 & n20806 ;
  assign n20808 = \s8_data_i[26]_pad  & n14717 ;
  assign n20809 = \s1_data_i[26]_pad  & n14622 ;
  assign n20810 = ~n20808 & ~n20809 ;
  assign n20811 = \s4_data_i[26]_pad  & n14727 ;
  assign n20812 = \s6_data_i[26]_pad  & n14723 ;
  assign n20813 = ~n20811 & ~n20812 ;
  assign n20814 = n20810 & n20813 ;
  assign n20815 = \s3_data_i[26]_pad  & n14950 ;
  assign n20816 = \s9_data_i[26]_pad  & n14713 ;
  assign n20817 = ~n20815 & ~n20816 ;
  assign n20818 = \s10_data_i[26]_pad  & n14931 ;
  assign n20819 = \s7_data_i[26]_pad  & n14958 ;
  assign n20820 = ~n20818 & ~n20819 ;
  assign n20821 = n20817 & n20820 ;
  assign n20822 = n20814 & n20821 ;
  assign n20823 = \s11_data_i[26]_pad  & n14735 ;
  assign n20824 = \s14_data_i[26]_pad  & n14939 ;
  assign n20825 = \s2_data_i[26]_pad  & n14946 ;
  assign n20826 = ~n20824 & ~n20825 ;
  assign n20827 = ~n20823 & n20826 ;
  assign n20828 = \s5_data_i[26]_pad  & n14954 ;
  assign n20829 = \s12_data_i[26]_pad  & n14935 ;
  assign n20830 = ~n20828 & ~n20829 ;
  assign n20831 = \s13_data_i[26]_pad  & n14731 ;
  assign n20832 = \s0_data_i[26]_pad  & n14616 ;
  assign n20833 = ~n20831 & ~n20832 ;
  assign n20834 = n20830 & n20833 ;
  assign n20835 = n20827 & n20834 ;
  assign n20836 = n20822 & n20835 ;
  assign n20837 = ~n20807 & n20836 ;
  assign n20838 = \s15_data_i[27]_pad  & n2197 ;
  assign n20839 = ~n2258 & n20838 ;
  assign n20840 = \s8_data_i[27]_pad  & n14717 ;
  assign n20841 = \s1_data_i[27]_pad  & n14622 ;
  assign n20842 = ~n20840 & ~n20841 ;
  assign n20843 = \s4_data_i[27]_pad  & n14727 ;
  assign n20844 = \s6_data_i[27]_pad  & n14723 ;
  assign n20845 = ~n20843 & ~n20844 ;
  assign n20846 = n20842 & n20845 ;
  assign n20847 = \s3_data_i[27]_pad  & n14950 ;
  assign n20848 = \s9_data_i[27]_pad  & n14713 ;
  assign n20849 = ~n20847 & ~n20848 ;
  assign n20850 = \s10_data_i[27]_pad  & n14931 ;
  assign n20851 = \s7_data_i[27]_pad  & n14958 ;
  assign n20852 = ~n20850 & ~n20851 ;
  assign n20853 = n20849 & n20852 ;
  assign n20854 = n20846 & n20853 ;
  assign n20855 = \s11_data_i[27]_pad  & n14735 ;
  assign n20856 = \s14_data_i[27]_pad  & n14939 ;
  assign n20857 = \s2_data_i[27]_pad  & n14946 ;
  assign n20858 = ~n20856 & ~n20857 ;
  assign n20859 = ~n20855 & n20858 ;
  assign n20860 = \s5_data_i[27]_pad  & n14954 ;
  assign n20861 = \s12_data_i[27]_pad  & n14935 ;
  assign n20862 = ~n20860 & ~n20861 ;
  assign n20863 = \s13_data_i[27]_pad  & n14731 ;
  assign n20864 = \s0_data_i[27]_pad  & n14616 ;
  assign n20865 = ~n20863 & ~n20864 ;
  assign n20866 = n20862 & n20865 ;
  assign n20867 = n20859 & n20866 ;
  assign n20868 = n20854 & n20867 ;
  assign n20869 = ~n20839 & n20868 ;
  assign n20870 = \s15_data_i[28]_pad  & n2197 ;
  assign n20871 = ~n2258 & n20870 ;
  assign n20872 = \s8_data_i[28]_pad  & n14717 ;
  assign n20873 = \s1_data_i[28]_pad  & n14622 ;
  assign n20874 = ~n20872 & ~n20873 ;
  assign n20875 = \s4_data_i[28]_pad  & n14727 ;
  assign n20876 = \s6_data_i[28]_pad  & n14723 ;
  assign n20877 = ~n20875 & ~n20876 ;
  assign n20878 = n20874 & n20877 ;
  assign n20879 = \s3_data_i[28]_pad  & n14950 ;
  assign n20880 = \s9_data_i[28]_pad  & n14713 ;
  assign n20881 = ~n20879 & ~n20880 ;
  assign n20882 = \s10_data_i[28]_pad  & n14931 ;
  assign n20883 = \s7_data_i[28]_pad  & n14958 ;
  assign n20884 = ~n20882 & ~n20883 ;
  assign n20885 = n20881 & n20884 ;
  assign n20886 = n20878 & n20885 ;
  assign n20887 = \s11_data_i[28]_pad  & n14735 ;
  assign n20888 = \s14_data_i[28]_pad  & n14939 ;
  assign n20889 = \s2_data_i[28]_pad  & n14946 ;
  assign n20890 = ~n20888 & ~n20889 ;
  assign n20891 = ~n20887 & n20890 ;
  assign n20892 = \s5_data_i[28]_pad  & n14954 ;
  assign n20893 = \s12_data_i[28]_pad  & n14935 ;
  assign n20894 = ~n20892 & ~n20893 ;
  assign n20895 = \s13_data_i[28]_pad  & n14731 ;
  assign n20896 = \s0_data_i[28]_pad  & n14616 ;
  assign n20897 = ~n20895 & ~n20896 ;
  assign n20898 = n20894 & n20897 ;
  assign n20899 = n20891 & n20898 ;
  assign n20900 = n20886 & n20899 ;
  assign n20901 = ~n20871 & n20900 ;
  assign n20902 = \s15_data_i[29]_pad  & n2197 ;
  assign n20903 = ~n2258 & n20902 ;
  assign n20904 = \s8_data_i[29]_pad  & n14717 ;
  assign n20905 = \s1_data_i[29]_pad  & n14622 ;
  assign n20906 = ~n20904 & ~n20905 ;
  assign n20907 = \s4_data_i[29]_pad  & n14727 ;
  assign n20908 = \s6_data_i[29]_pad  & n14723 ;
  assign n20909 = ~n20907 & ~n20908 ;
  assign n20910 = n20906 & n20909 ;
  assign n20911 = \s3_data_i[29]_pad  & n14950 ;
  assign n20912 = \s9_data_i[29]_pad  & n14713 ;
  assign n20913 = ~n20911 & ~n20912 ;
  assign n20914 = \s10_data_i[29]_pad  & n14931 ;
  assign n20915 = \s7_data_i[29]_pad  & n14958 ;
  assign n20916 = ~n20914 & ~n20915 ;
  assign n20917 = n20913 & n20916 ;
  assign n20918 = n20910 & n20917 ;
  assign n20919 = \s11_data_i[29]_pad  & n14735 ;
  assign n20920 = \s14_data_i[29]_pad  & n14939 ;
  assign n20921 = \s2_data_i[29]_pad  & n14946 ;
  assign n20922 = ~n20920 & ~n20921 ;
  assign n20923 = ~n20919 & n20922 ;
  assign n20924 = \s5_data_i[29]_pad  & n14954 ;
  assign n20925 = \s12_data_i[29]_pad  & n14935 ;
  assign n20926 = ~n20924 & ~n20925 ;
  assign n20927 = \s13_data_i[29]_pad  & n14731 ;
  assign n20928 = \s0_data_i[29]_pad  & n14616 ;
  assign n20929 = ~n20927 & ~n20928 ;
  assign n20930 = n20926 & n20929 ;
  assign n20931 = n20923 & n20930 ;
  assign n20932 = n20918 & n20931 ;
  assign n20933 = ~n20903 & n20932 ;
  assign n20934 = n2197 & n15936 ;
  assign n20935 = \s15_data_i[2]_pad  & n2197 ;
  assign n20936 = ~n2258 & n20935 ;
  assign n20937 = ~n20934 & ~n20936 ;
  assign n20938 = \s8_data_i[2]_pad  & n14717 ;
  assign n20939 = \s1_data_i[2]_pad  & n14622 ;
  assign n20940 = ~n20938 & ~n20939 ;
  assign n20941 = \s4_data_i[2]_pad  & n14727 ;
  assign n20942 = \s6_data_i[2]_pad  & n14723 ;
  assign n20943 = ~n20941 & ~n20942 ;
  assign n20944 = n20940 & n20943 ;
  assign n20945 = \s3_data_i[2]_pad  & n14950 ;
  assign n20946 = \s9_data_i[2]_pad  & n14713 ;
  assign n20947 = ~n20945 & ~n20946 ;
  assign n20948 = \s10_data_i[2]_pad  & n14931 ;
  assign n20949 = \s7_data_i[2]_pad  & n14958 ;
  assign n20950 = ~n20948 & ~n20949 ;
  assign n20951 = n20947 & n20950 ;
  assign n20952 = n20944 & n20951 ;
  assign n20953 = \s11_data_i[2]_pad  & n14735 ;
  assign n20954 = \s14_data_i[2]_pad  & n14939 ;
  assign n20955 = \s2_data_i[2]_pad  & n14946 ;
  assign n20956 = ~n20954 & ~n20955 ;
  assign n20957 = ~n20953 & n20956 ;
  assign n20958 = \s5_data_i[2]_pad  & n14954 ;
  assign n20959 = \s12_data_i[2]_pad  & n14935 ;
  assign n20960 = ~n20958 & ~n20959 ;
  assign n20961 = \s13_data_i[2]_pad  & n14731 ;
  assign n20962 = \s0_data_i[2]_pad  & n14616 ;
  assign n20963 = ~n20961 & ~n20962 ;
  assign n20964 = n20960 & n20963 ;
  assign n20965 = n20957 & n20964 ;
  assign n20966 = n20952 & n20965 ;
  assign n20967 = n20937 & n20966 ;
  assign n20968 = \s15_data_i[30]_pad  & n2197 ;
  assign n20969 = ~n2258 & n20968 ;
  assign n20970 = \s8_data_i[30]_pad  & n14717 ;
  assign n20971 = \s1_data_i[30]_pad  & n14622 ;
  assign n20972 = ~n20970 & ~n20971 ;
  assign n20973 = \s4_data_i[30]_pad  & n14727 ;
  assign n20974 = \s6_data_i[30]_pad  & n14723 ;
  assign n20975 = ~n20973 & ~n20974 ;
  assign n20976 = n20972 & n20975 ;
  assign n20977 = \s3_data_i[30]_pad  & n14950 ;
  assign n20978 = \s9_data_i[30]_pad  & n14713 ;
  assign n20979 = ~n20977 & ~n20978 ;
  assign n20980 = \s10_data_i[30]_pad  & n14931 ;
  assign n20981 = \s7_data_i[30]_pad  & n14958 ;
  assign n20982 = ~n20980 & ~n20981 ;
  assign n20983 = n20979 & n20982 ;
  assign n20984 = n20976 & n20983 ;
  assign n20985 = \s11_data_i[30]_pad  & n14735 ;
  assign n20986 = \s14_data_i[30]_pad  & n14939 ;
  assign n20987 = \s2_data_i[30]_pad  & n14946 ;
  assign n20988 = ~n20986 & ~n20987 ;
  assign n20989 = ~n20985 & n20988 ;
  assign n20990 = \s5_data_i[30]_pad  & n14954 ;
  assign n20991 = \s12_data_i[30]_pad  & n14935 ;
  assign n20992 = ~n20990 & ~n20991 ;
  assign n20993 = \s13_data_i[30]_pad  & n14731 ;
  assign n20994 = \s0_data_i[30]_pad  & n14616 ;
  assign n20995 = ~n20993 & ~n20994 ;
  assign n20996 = n20992 & n20995 ;
  assign n20997 = n20989 & n20996 ;
  assign n20998 = n20984 & n20997 ;
  assign n20999 = ~n20969 & n20998 ;
  assign n21000 = \s15_data_i[31]_pad  & n2197 ;
  assign n21001 = ~n2258 & n21000 ;
  assign n21002 = \s8_data_i[31]_pad  & n14717 ;
  assign n21003 = \s1_data_i[31]_pad  & n14622 ;
  assign n21004 = ~n21002 & ~n21003 ;
  assign n21005 = \s4_data_i[31]_pad  & n14727 ;
  assign n21006 = \s6_data_i[31]_pad  & n14723 ;
  assign n21007 = ~n21005 & ~n21006 ;
  assign n21008 = n21004 & n21007 ;
  assign n21009 = \s3_data_i[31]_pad  & n14950 ;
  assign n21010 = \s9_data_i[31]_pad  & n14713 ;
  assign n21011 = ~n21009 & ~n21010 ;
  assign n21012 = \s10_data_i[31]_pad  & n14931 ;
  assign n21013 = \s7_data_i[31]_pad  & n14958 ;
  assign n21014 = ~n21012 & ~n21013 ;
  assign n21015 = n21011 & n21014 ;
  assign n21016 = n21008 & n21015 ;
  assign n21017 = \s11_data_i[31]_pad  & n14735 ;
  assign n21018 = \s14_data_i[31]_pad  & n14939 ;
  assign n21019 = \s2_data_i[31]_pad  & n14946 ;
  assign n21020 = ~n21018 & ~n21019 ;
  assign n21021 = ~n21017 & n21020 ;
  assign n21022 = \s5_data_i[31]_pad  & n14954 ;
  assign n21023 = \s12_data_i[31]_pad  & n14935 ;
  assign n21024 = ~n21022 & ~n21023 ;
  assign n21025 = \s13_data_i[31]_pad  & n14731 ;
  assign n21026 = \s0_data_i[31]_pad  & n14616 ;
  assign n21027 = ~n21025 & ~n21026 ;
  assign n21028 = n21024 & n21027 ;
  assign n21029 = n21021 & n21028 ;
  assign n21030 = n21016 & n21029 ;
  assign n21031 = ~n21001 & n21030 ;
  assign n21032 = n2197 & n16037 ;
  assign n21033 = \s15_data_i[3]_pad  & n2197 ;
  assign n21034 = ~n2258 & n21033 ;
  assign n21035 = ~n21032 & ~n21034 ;
  assign n21036 = \s8_data_i[3]_pad  & n14717 ;
  assign n21037 = \s1_data_i[3]_pad  & n14622 ;
  assign n21038 = ~n21036 & ~n21037 ;
  assign n21039 = \s4_data_i[3]_pad  & n14727 ;
  assign n21040 = \s6_data_i[3]_pad  & n14723 ;
  assign n21041 = ~n21039 & ~n21040 ;
  assign n21042 = n21038 & n21041 ;
  assign n21043 = \s3_data_i[3]_pad  & n14950 ;
  assign n21044 = \s9_data_i[3]_pad  & n14713 ;
  assign n21045 = ~n21043 & ~n21044 ;
  assign n21046 = \s10_data_i[3]_pad  & n14931 ;
  assign n21047 = \s7_data_i[3]_pad  & n14958 ;
  assign n21048 = ~n21046 & ~n21047 ;
  assign n21049 = n21045 & n21048 ;
  assign n21050 = n21042 & n21049 ;
  assign n21051 = \s11_data_i[3]_pad  & n14735 ;
  assign n21052 = \s14_data_i[3]_pad  & n14939 ;
  assign n21053 = \s2_data_i[3]_pad  & n14946 ;
  assign n21054 = ~n21052 & ~n21053 ;
  assign n21055 = ~n21051 & n21054 ;
  assign n21056 = \s5_data_i[3]_pad  & n14954 ;
  assign n21057 = \s12_data_i[3]_pad  & n14935 ;
  assign n21058 = ~n21056 & ~n21057 ;
  assign n21059 = \s13_data_i[3]_pad  & n14731 ;
  assign n21060 = \s0_data_i[3]_pad  & n14616 ;
  assign n21061 = ~n21059 & ~n21060 ;
  assign n21062 = n21058 & n21061 ;
  assign n21063 = n21055 & n21062 ;
  assign n21064 = n21050 & n21063 ;
  assign n21065 = n21035 & n21064 ;
  assign n21066 = n2197 & n16074 ;
  assign n21067 = \s15_data_i[4]_pad  & n2197 ;
  assign n21068 = ~n2258 & n21067 ;
  assign n21069 = ~n21066 & ~n21068 ;
  assign n21070 = \s8_data_i[4]_pad  & n14717 ;
  assign n21071 = \s1_data_i[4]_pad  & n14622 ;
  assign n21072 = ~n21070 & ~n21071 ;
  assign n21073 = \s4_data_i[4]_pad  & n14727 ;
  assign n21074 = \s6_data_i[4]_pad  & n14723 ;
  assign n21075 = ~n21073 & ~n21074 ;
  assign n21076 = n21072 & n21075 ;
  assign n21077 = \s3_data_i[4]_pad  & n14950 ;
  assign n21078 = \s9_data_i[4]_pad  & n14713 ;
  assign n21079 = ~n21077 & ~n21078 ;
  assign n21080 = \s10_data_i[4]_pad  & n14931 ;
  assign n21081 = \s7_data_i[4]_pad  & n14958 ;
  assign n21082 = ~n21080 & ~n21081 ;
  assign n21083 = n21079 & n21082 ;
  assign n21084 = n21076 & n21083 ;
  assign n21085 = \s11_data_i[4]_pad  & n14735 ;
  assign n21086 = \s14_data_i[4]_pad  & n14939 ;
  assign n21087 = \s2_data_i[4]_pad  & n14946 ;
  assign n21088 = ~n21086 & ~n21087 ;
  assign n21089 = ~n21085 & n21088 ;
  assign n21090 = \s5_data_i[4]_pad  & n14954 ;
  assign n21091 = \s12_data_i[4]_pad  & n14935 ;
  assign n21092 = ~n21090 & ~n21091 ;
  assign n21093 = \s13_data_i[4]_pad  & n14731 ;
  assign n21094 = \s0_data_i[4]_pad  & n14616 ;
  assign n21095 = ~n21093 & ~n21094 ;
  assign n21096 = n21092 & n21095 ;
  assign n21097 = n21089 & n21096 ;
  assign n21098 = n21084 & n21097 ;
  assign n21099 = n21069 & n21098 ;
  assign n21100 = n2197 & n16111 ;
  assign n21101 = \s15_data_i[5]_pad  & n2197 ;
  assign n21102 = ~n2258 & n21101 ;
  assign n21103 = ~n21100 & ~n21102 ;
  assign n21104 = \s8_data_i[5]_pad  & n14717 ;
  assign n21105 = \s1_data_i[5]_pad  & n14622 ;
  assign n21106 = ~n21104 & ~n21105 ;
  assign n21107 = \s4_data_i[5]_pad  & n14727 ;
  assign n21108 = \s6_data_i[5]_pad  & n14723 ;
  assign n21109 = ~n21107 & ~n21108 ;
  assign n21110 = n21106 & n21109 ;
  assign n21111 = \s3_data_i[5]_pad  & n14950 ;
  assign n21112 = \s9_data_i[5]_pad  & n14713 ;
  assign n21113 = ~n21111 & ~n21112 ;
  assign n21114 = \s10_data_i[5]_pad  & n14931 ;
  assign n21115 = \s7_data_i[5]_pad  & n14958 ;
  assign n21116 = ~n21114 & ~n21115 ;
  assign n21117 = n21113 & n21116 ;
  assign n21118 = n21110 & n21117 ;
  assign n21119 = \s11_data_i[5]_pad  & n14735 ;
  assign n21120 = \s14_data_i[5]_pad  & n14939 ;
  assign n21121 = \s2_data_i[5]_pad  & n14946 ;
  assign n21122 = ~n21120 & ~n21121 ;
  assign n21123 = ~n21119 & n21122 ;
  assign n21124 = \s5_data_i[5]_pad  & n14954 ;
  assign n21125 = \s12_data_i[5]_pad  & n14935 ;
  assign n21126 = ~n21124 & ~n21125 ;
  assign n21127 = \s13_data_i[5]_pad  & n14731 ;
  assign n21128 = \s0_data_i[5]_pad  & n14616 ;
  assign n21129 = ~n21127 & ~n21128 ;
  assign n21130 = n21126 & n21129 ;
  assign n21131 = n21123 & n21130 ;
  assign n21132 = n21118 & n21131 ;
  assign n21133 = n21103 & n21132 ;
  assign n21134 = n2197 & n16148 ;
  assign n21135 = \s15_data_i[6]_pad  & n2197 ;
  assign n21136 = ~n2258 & n21135 ;
  assign n21137 = ~n21134 & ~n21136 ;
  assign n21138 = \s11_data_i[6]_pad  & n14735 ;
  assign n21139 = \s1_data_i[6]_pad  & n14622 ;
  assign n21140 = ~n21138 & ~n21139 ;
  assign n21141 = \s4_data_i[6]_pad  & n14727 ;
  assign n21142 = \s6_data_i[6]_pad  & n14723 ;
  assign n21143 = ~n21141 & ~n21142 ;
  assign n21144 = n21140 & n21143 ;
  assign n21145 = \s5_data_i[6]_pad  & n14954 ;
  assign n21146 = \s9_data_i[6]_pad  & n14713 ;
  assign n21147 = ~n21145 & ~n21146 ;
  assign n21148 = \s10_data_i[6]_pad  & n14931 ;
  assign n21149 = \s7_data_i[6]_pad  & n14958 ;
  assign n21150 = ~n21148 & ~n21149 ;
  assign n21151 = n21147 & n21150 ;
  assign n21152 = n21144 & n21151 ;
  assign n21153 = \s12_data_i[6]_pad  & n14935 ;
  assign n21154 = \s2_data_i[6]_pad  & n14946 ;
  assign n21155 = \s3_data_i[6]_pad  & n14950 ;
  assign n21156 = ~n21154 & ~n21155 ;
  assign n21157 = ~n21153 & n21156 ;
  assign n21158 = \s8_data_i[6]_pad  & n14717 ;
  assign n21159 = \s14_data_i[6]_pad  & n14939 ;
  assign n21160 = ~n21158 & ~n21159 ;
  assign n21161 = \s13_data_i[6]_pad  & n14731 ;
  assign n21162 = \s0_data_i[6]_pad  & n14616 ;
  assign n21163 = ~n21161 & ~n21162 ;
  assign n21164 = n21160 & n21163 ;
  assign n21165 = n21157 & n21164 ;
  assign n21166 = n21152 & n21165 ;
  assign n21167 = n21137 & n21166 ;
  assign n21168 = n2197 & n16185 ;
  assign n21169 = \s15_data_i[7]_pad  & n2197 ;
  assign n21170 = ~n2258 & n21169 ;
  assign n21171 = ~n21168 & ~n21170 ;
  assign n21172 = \s8_data_i[7]_pad  & n14717 ;
  assign n21173 = \s1_data_i[7]_pad  & n14622 ;
  assign n21174 = ~n21172 & ~n21173 ;
  assign n21175 = \s4_data_i[7]_pad  & n14727 ;
  assign n21176 = \s6_data_i[7]_pad  & n14723 ;
  assign n21177 = ~n21175 & ~n21176 ;
  assign n21178 = n21174 & n21177 ;
  assign n21179 = \s3_data_i[7]_pad  & n14950 ;
  assign n21180 = \s9_data_i[7]_pad  & n14713 ;
  assign n21181 = ~n21179 & ~n21180 ;
  assign n21182 = \s10_data_i[7]_pad  & n14931 ;
  assign n21183 = \s7_data_i[7]_pad  & n14958 ;
  assign n21184 = ~n21182 & ~n21183 ;
  assign n21185 = n21181 & n21184 ;
  assign n21186 = n21178 & n21185 ;
  assign n21187 = \s11_data_i[7]_pad  & n14735 ;
  assign n21188 = \s14_data_i[7]_pad  & n14939 ;
  assign n21189 = \s2_data_i[7]_pad  & n14946 ;
  assign n21190 = ~n21188 & ~n21189 ;
  assign n21191 = ~n21187 & n21190 ;
  assign n21192 = \s5_data_i[7]_pad  & n14954 ;
  assign n21193 = \s12_data_i[7]_pad  & n14935 ;
  assign n21194 = ~n21192 & ~n21193 ;
  assign n21195 = \s13_data_i[7]_pad  & n14731 ;
  assign n21196 = \s0_data_i[7]_pad  & n14616 ;
  assign n21197 = ~n21195 & ~n21196 ;
  assign n21198 = n21194 & n21197 ;
  assign n21199 = n21191 & n21198 ;
  assign n21200 = n21186 & n21199 ;
  assign n21201 = n21171 & n21200 ;
  assign n21202 = n2197 & n16222 ;
  assign n21203 = \s15_data_i[8]_pad  & n2197 ;
  assign n21204 = ~n2258 & n21203 ;
  assign n21205 = ~n21202 & ~n21204 ;
  assign n21206 = \s8_data_i[8]_pad  & n14717 ;
  assign n21207 = \s1_data_i[8]_pad  & n14622 ;
  assign n21208 = ~n21206 & ~n21207 ;
  assign n21209 = \s4_data_i[8]_pad  & n14727 ;
  assign n21210 = \s6_data_i[8]_pad  & n14723 ;
  assign n21211 = ~n21209 & ~n21210 ;
  assign n21212 = n21208 & n21211 ;
  assign n21213 = \s3_data_i[8]_pad  & n14950 ;
  assign n21214 = \s9_data_i[8]_pad  & n14713 ;
  assign n21215 = ~n21213 & ~n21214 ;
  assign n21216 = \s10_data_i[8]_pad  & n14931 ;
  assign n21217 = \s7_data_i[8]_pad  & n14958 ;
  assign n21218 = ~n21216 & ~n21217 ;
  assign n21219 = n21215 & n21218 ;
  assign n21220 = n21212 & n21219 ;
  assign n21221 = \s11_data_i[8]_pad  & n14735 ;
  assign n21222 = \s14_data_i[8]_pad  & n14939 ;
  assign n21223 = \s2_data_i[8]_pad  & n14946 ;
  assign n21224 = ~n21222 & ~n21223 ;
  assign n21225 = ~n21221 & n21224 ;
  assign n21226 = \s5_data_i[8]_pad  & n14954 ;
  assign n21227 = \s12_data_i[8]_pad  & n14935 ;
  assign n21228 = ~n21226 & ~n21227 ;
  assign n21229 = \s13_data_i[8]_pad  & n14731 ;
  assign n21230 = \s0_data_i[8]_pad  & n14616 ;
  assign n21231 = ~n21229 & ~n21230 ;
  assign n21232 = n21228 & n21231 ;
  assign n21233 = n21225 & n21232 ;
  assign n21234 = n21220 & n21233 ;
  assign n21235 = n21205 & n21234 ;
  assign n21236 = n2197 & n16259 ;
  assign n21237 = \s15_data_i[9]_pad  & n2197 ;
  assign n21238 = ~n2258 & n21237 ;
  assign n21239 = ~n21236 & ~n21238 ;
  assign n21240 = \s8_data_i[9]_pad  & n14717 ;
  assign n21241 = \s1_data_i[9]_pad  & n14622 ;
  assign n21242 = ~n21240 & ~n21241 ;
  assign n21243 = \s4_data_i[9]_pad  & n14727 ;
  assign n21244 = \s6_data_i[9]_pad  & n14723 ;
  assign n21245 = ~n21243 & ~n21244 ;
  assign n21246 = n21242 & n21245 ;
  assign n21247 = \s3_data_i[9]_pad  & n14950 ;
  assign n21248 = \s9_data_i[9]_pad  & n14713 ;
  assign n21249 = ~n21247 & ~n21248 ;
  assign n21250 = \s10_data_i[9]_pad  & n14931 ;
  assign n21251 = \s7_data_i[9]_pad  & n14958 ;
  assign n21252 = ~n21250 & ~n21251 ;
  assign n21253 = n21249 & n21252 ;
  assign n21254 = n21246 & n21253 ;
  assign n21255 = \s11_data_i[9]_pad  & n14735 ;
  assign n21256 = \s14_data_i[9]_pad  & n14939 ;
  assign n21257 = \s2_data_i[9]_pad  & n14946 ;
  assign n21258 = ~n21256 & ~n21257 ;
  assign n21259 = ~n21255 & n21258 ;
  assign n21260 = \s5_data_i[9]_pad  & n14954 ;
  assign n21261 = \s12_data_i[9]_pad  & n14935 ;
  assign n21262 = ~n21260 & ~n21261 ;
  assign n21263 = \s13_data_i[9]_pad  & n14731 ;
  assign n21264 = \s0_data_i[9]_pad  & n14616 ;
  assign n21265 = ~n21263 & ~n21264 ;
  assign n21266 = n21262 & n21265 ;
  assign n21267 = n21259 & n21266 ;
  assign n21268 = n21254 & n21267 ;
  assign n21269 = n21239 & n21268 ;
  assign n21270 = \s15_err_i_pad  & n20151 ;
  assign n21271 = ~n2258 & n21270 ;
  assign n21272 = \s6_err_i_pad  & n14723 ;
  assign n21273 = n13627 & n21272 ;
  assign n21274 = n13652 & n21273 ;
  assign n21275 = \s1_err_i_pad  & n14622 ;
  assign n21276 = n14271 & n21275 ;
  assign n21277 = n14288 & n21276 ;
  assign n21278 = ~n21274 & ~n21277 ;
  assign n21279 = \s7_err_i_pad  & n14958 ;
  assign n21280 = n13697 & n21279 ;
  assign n21281 = n13722 & n21280 ;
  assign n21282 = \s3_err_i_pad  & n14950 ;
  assign n21283 = n14451 & n21282 ;
  assign n21284 = n14444 & n21283 ;
  assign n21285 = ~n21281 & ~n21284 ;
  assign n21286 = n21278 & n21285 ;
  assign n21287 = \s14_err_i_pad  & n14939 ;
  assign n21288 = n14331 & n21287 ;
  assign n21289 = n14356 & n21288 ;
  assign n21290 = \s13_err_i_pad  & n14731 ;
  assign n21291 = n14211 & n21290 ;
  assign n21292 = n14236 & n21291 ;
  assign n21293 = ~n21289 & ~n21292 ;
  assign n21294 = \s10_err_i_pad  & n14931 ;
  assign n21295 = n13928 & n21294 ;
  assign n21296 = n13953 & n21295 ;
  assign n21297 = \s9_err_i_pad  & n14713 ;
  assign n21298 = n13847 & n21297 ;
  assign n21299 = n13872 & n21298 ;
  assign n21300 = ~n21296 & ~n21299 ;
  assign n21301 = n21293 & n21300 ;
  assign n21302 = n21286 & n21301 ;
  assign n21303 = \s0_err_i_pad  & n14616 ;
  assign n21304 = n14069 & n21303 ;
  assign n21305 = n14077 & n21304 ;
  assign n21306 = \s11_err_i_pad  & n14735 ;
  assign n21307 = n14009 & n21306 ;
  assign n21308 = n14002 & n21307 ;
  assign n21309 = \s5_err_i_pad  & n14954 ;
  assign n21310 = n13547 & n21309 ;
  assign n21311 = n13555 & n21310 ;
  assign n21312 = ~n21308 & ~n21311 ;
  assign n21313 = ~n21305 & n21312 ;
  assign n21314 = \s12_err_i_pad  & n14935 ;
  assign n21315 = n14140 & n21314 ;
  assign n21316 = n14157 & n21315 ;
  assign n21317 = \s4_err_i_pad  & n14727 ;
  assign n21318 = n13467 & n21317 ;
  assign n21319 = n13460 & n21318 ;
  assign n21320 = ~n21316 & ~n21319 ;
  assign n21321 = \s2_err_i_pad  & n14946 ;
  assign n21322 = n14391 & n21321 ;
  assign n21323 = n14384 & n21322 ;
  assign n21324 = \s8_err_i_pad  & n14717 ;
  assign n21325 = n13767 & n21324 ;
  assign n21326 = n13792 & n21325 ;
  assign n21327 = ~n21323 & ~n21326 ;
  assign n21328 = n21320 & n21327 ;
  assign n21329 = n21313 & n21328 ;
  assign n21330 = n21302 & n21329 ;
  assign n21331 = ~n21271 & n21330 ;
  assign n21332 = \s15_rty_i_pad  & n20151 ;
  assign n21333 = ~n2258 & n21332 ;
  assign n21334 = \s14_rty_i_pad  & n14939 ;
  assign n21335 = n14331 & n21334 ;
  assign n21336 = n14356 & n21335 ;
  assign n21337 = \s1_rty_i_pad  & n14622 ;
  assign n21338 = n14271 & n21337 ;
  assign n21339 = n14288 & n21338 ;
  assign n21340 = ~n21336 & ~n21339 ;
  assign n21341 = \s10_rty_i_pad  & n14931 ;
  assign n21342 = n13928 & n21341 ;
  assign n21343 = n13953 & n21342 ;
  assign n21344 = \s7_rty_i_pad  & n14958 ;
  assign n21345 = n13697 & n21344 ;
  assign n21346 = n13722 & n21345 ;
  assign n21347 = ~n21343 & ~n21346 ;
  assign n21348 = n21340 & n21347 ;
  assign n21349 = \s8_rty_i_pad  & n14717 ;
  assign n21350 = n13767 & n21349 ;
  assign n21351 = n13792 & n21350 ;
  assign n21352 = \s9_rty_i_pad  & n14713 ;
  assign n21353 = n13847 & n21352 ;
  assign n21354 = n13872 & n21353 ;
  assign n21355 = ~n21351 & ~n21354 ;
  assign n21356 = \s6_rty_i_pad  & n14723 ;
  assign n21357 = n13627 & n21356 ;
  assign n21358 = n13652 & n21357 ;
  assign n21359 = \s13_rty_i_pad  & n14731 ;
  assign n21360 = n14211 & n21359 ;
  assign n21361 = n14236 & n21360 ;
  assign n21362 = ~n21358 & ~n21361 ;
  assign n21363 = n21355 & n21362 ;
  assign n21364 = n21348 & n21363 ;
  assign n21365 = \s12_rty_i_pad  & n14935 ;
  assign n21366 = n14140 & n21365 ;
  assign n21367 = n14157 & n21366 ;
  assign n21368 = \s5_rty_i_pad  & n14954 ;
  assign n21369 = n13547 & n21368 ;
  assign n21370 = n13555 & n21369 ;
  assign n21371 = \s4_rty_i_pad  & n14727 ;
  assign n21372 = n13467 & n21371 ;
  assign n21373 = n13460 & n21372 ;
  assign n21374 = ~n21370 & ~n21373 ;
  assign n21375 = ~n21367 & n21374 ;
  assign n21376 = \s0_rty_i_pad  & n14616 ;
  assign n21377 = n14069 & n21376 ;
  assign n21378 = n14077 & n21377 ;
  assign n21379 = \s11_rty_i_pad  & n14735 ;
  assign n21380 = n14009 & n21379 ;
  assign n21381 = n14002 & n21380 ;
  assign n21382 = ~n21378 & ~n21381 ;
  assign n21383 = \s2_rty_i_pad  & n14946 ;
  assign n21384 = n14391 & n21383 ;
  assign n21385 = n14384 & n21384 ;
  assign n21386 = \s3_rty_i_pad  & n14950 ;
  assign n21387 = n14451 & n21386 ;
  assign n21388 = n14444 & n21387 ;
  assign n21389 = ~n21385 & ~n21388 ;
  assign n21390 = n21382 & n21389 ;
  assign n21391 = n21375 & n21390 ;
  assign n21392 = n21364 & n21391 ;
  assign n21393 = ~n21333 & n21392 ;
  assign n21394 = ~n1910 & n2203 ;
  assign n21395 = n1941 & n21394 ;
  assign n21396 = ~n13416 & n21395 ;
  assign n21397 = ~n15125 & n21396 ;
  assign n21398 = \s11_ack_i_pad  & n14967 ;
  assign n21399 = ~n14009 & n21398 ;
  assign n21400 = n14002 & n21399 ;
  assign n21401 = \s3_ack_i_pad  & n14704 ;
  assign n21402 = ~n14451 & n21401 ;
  assign n21403 = n14444 & n21402 ;
  assign n21404 = ~n21400 & ~n21403 ;
  assign n21405 = \s1_ack_i_pad  & n14561 ;
  assign n21406 = ~n14271 & n21405 ;
  assign n21407 = n14288 & n21406 ;
  assign n21408 = \s7_ack_i_pad  & n14695 ;
  assign n21409 = ~n13697 & n21408 ;
  assign n21410 = n13722 & n21409 ;
  assign n21411 = ~n21407 & ~n21410 ;
  assign n21412 = n21404 & n21411 ;
  assign n21413 = \s10_ack_i_pad  & n14963 ;
  assign n21414 = ~n13928 & n21413 ;
  assign n21415 = n13953 & n21414 ;
  assign n21416 = \s2_ack_i_pad  & n14975 ;
  assign n21417 = ~n14391 & n21416 ;
  assign n21418 = n14384 & n21417 ;
  assign n21419 = ~n21415 & ~n21418 ;
  assign n21420 = \s13_ack_i_pad  & n14971 ;
  assign n21421 = ~n14211 & n21420 ;
  assign n21422 = n14236 & n21421 ;
  assign n21423 = \s6_ack_i_pad  & n14987 ;
  assign n21424 = ~n13627 & n21423 ;
  assign n21425 = n13652 & n21424 ;
  assign n21426 = ~n21422 & ~n21425 ;
  assign n21427 = n21419 & n21426 ;
  assign n21428 = n21412 & n21427 ;
  assign n21429 = \s8_ack_i_pad  & n14991 ;
  assign n21430 = ~n13767 & n21429 ;
  assign n21431 = n13792 & n21430 ;
  assign n21432 = \s14_ack_i_pad  & n14700 ;
  assign n21433 = ~n14331 & n21432 ;
  assign n21434 = n14356 & n21433 ;
  assign n21435 = \s9_ack_i_pad  & n14995 ;
  assign n21436 = ~n13847 & n21435 ;
  assign n21437 = n13872 & n21436 ;
  assign n21438 = ~n21434 & ~n21437 ;
  assign n21439 = ~n21431 & n21438 ;
  assign n21440 = \s4_ack_i_pad  & n14979 ;
  assign n21441 = ~n13467 & n21440 ;
  assign n21442 = n13460 & n21441 ;
  assign n21443 = \s0_ack_i_pad  & n14627 ;
  assign n21444 = ~n14069 & n21443 ;
  assign n21445 = n14077 & n21444 ;
  assign n21446 = ~n21442 & ~n21445 ;
  assign n21447 = \s5_ack_i_pad  & n14983 ;
  assign n21448 = ~n13547 & n21447 ;
  assign n21449 = n13555 & n21448 ;
  assign n21450 = \s12_ack_i_pad  & n14708 ;
  assign n21451 = ~n14140 & n21450 ;
  assign n21452 = n14157 & n21451 ;
  assign n21453 = ~n21449 & ~n21452 ;
  assign n21454 = n21446 & n21453 ;
  assign n21455 = n21439 & n21454 ;
  assign n21456 = n21428 & n21455 ;
  assign n21457 = ~n21397 & n21456 ;
  assign n21458 = n2203 & n15192 ;
  assign n21459 = \s15_data_i[0]_pad  & n2203 ;
  assign n21460 = ~n2258 & n21459 ;
  assign n21461 = ~n21458 & ~n21460 ;
  assign n21462 = \s12_data_i[0]_pad  & n14708 ;
  assign n21463 = \s1_data_i[0]_pad  & n14561 ;
  assign n21464 = ~n21462 & ~n21463 ;
  assign n21465 = \s0_data_i[0]_pad  & n14627 ;
  assign n21466 = \s10_data_i[0]_pad  & n14963 ;
  assign n21467 = ~n21465 & ~n21466 ;
  assign n21468 = n21464 & n21467 ;
  assign n21469 = \s3_data_i[0]_pad  & n14704 ;
  assign n21470 = \s4_data_i[0]_pad  & n14979 ;
  assign n21471 = ~n21469 & ~n21470 ;
  assign n21472 = \s9_data_i[0]_pad  & n14995 ;
  assign n21473 = \s6_data_i[0]_pad  & n14987 ;
  assign n21474 = ~n21472 & ~n21473 ;
  assign n21475 = n21471 & n21474 ;
  assign n21476 = n21468 & n21475 ;
  assign n21477 = \s14_data_i[0]_pad  & n14700 ;
  assign n21478 = \s11_data_i[0]_pad  & n14967 ;
  assign n21479 = \s7_data_i[0]_pad  & n14695 ;
  assign n21480 = ~n21478 & ~n21479 ;
  assign n21481 = ~n21477 & n21480 ;
  assign n21482 = \s5_data_i[0]_pad  & n14983 ;
  assign n21483 = \s8_data_i[0]_pad  & n14991 ;
  assign n21484 = ~n21482 & ~n21483 ;
  assign n21485 = \s2_data_i[0]_pad  & n14975 ;
  assign n21486 = \s13_data_i[0]_pad  & n14971 ;
  assign n21487 = ~n21485 & ~n21486 ;
  assign n21488 = n21484 & n21487 ;
  assign n21489 = n21481 & n21488 ;
  assign n21490 = n21476 & n21489 ;
  assign n21491 = n21461 & n21490 ;
  assign n21492 = n2203 & n15229 ;
  assign n21493 = \s15_data_i[10]_pad  & n2203 ;
  assign n21494 = ~n2258 & n21493 ;
  assign n21495 = ~n21492 & ~n21494 ;
  assign n21496 = \s12_data_i[10]_pad  & n14708 ;
  assign n21497 = \s1_data_i[10]_pad  & n14561 ;
  assign n21498 = ~n21496 & ~n21497 ;
  assign n21499 = \s0_data_i[10]_pad  & n14627 ;
  assign n21500 = \s10_data_i[10]_pad  & n14963 ;
  assign n21501 = ~n21499 & ~n21500 ;
  assign n21502 = n21498 & n21501 ;
  assign n21503 = \s3_data_i[10]_pad  & n14704 ;
  assign n21504 = \s4_data_i[10]_pad  & n14979 ;
  assign n21505 = ~n21503 & ~n21504 ;
  assign n21506 = \s9_data_i[10]_pad  & n14995 ;
  assign n21507 = \s6_data_i[10]_pad  & n14987 ;
  assign n21508 = ~n21506 & ~n21507 ;
  assign n21509 = n21505 & n21508 ;
  assign n21510 = n21502 & n21509 ;
  assign n21511 = \s14_data_i[10]_pad  & n14700 ;
  assign n21512 = \s11_data_i[10]_pad  & n14967 ;
  assign n21513 = \s7_data_i[10]_pad  & n14695 ;
  assign n21514 = ~n21512 & ~n21513 ;
  assign n21515 = ~n21511 & n21514 ;
  assign n21516 = \s5_data_i[10]_pad  & n14983 ;
  assign n21517 = \s8_data_i[10]_pad  & n14991 ;
  assign n21518 = ~n21516 & ~n21517 ;
  assign n21519 = \s2_data_i[10]_pad  & n14975 ;
  assign n21520 = \s13_data_i[10]_pad  & n14971 ;
  assign n21521 = ~n21519 & ~n21520 ;
  assign n21522 = n21518 & n21521 ;
  assign n21523 = n21515 & n21522 ;
  assign n21524 = n21510 & n21523 ;
  assign n21525 = n21495 & n21524 ;
  assign n21526 = n2203 & n15266 ;
  assign n21527 = \s15_data_i[11]_pad  & n2203 ;
  assign n21528 = ~n2258 & n21527 ;
  assign n21529 = ~n21526 & ~n21528 ;
  assign n21530 = \s7_data_i[11]_pad  & n14695 ;
  assign n21531 = \s1_data_i[11]_pad  & n14561 ;
  assign n21532 = ~n21530 & ~n21531 ;
  assign n21533 = \s2_data_i[11]_pad  & n14975 ;
  assign n21534 = \s5_data_i[11]_pad  & n14983 ;
  assign n21535 = ~n21533 & ~n21534 ;
  assign n21536 = n21532 & n21535 ;
  assign n21537 = \s12_data_i[11]_pad  & n14708 ;
  assign n21538 = \s3_data_i[11]_pad  & n14704 ;
  assign n21539 = ~n21537 & ~n21538 ;
  assign n21540 = \s8_data_i[11]_pad  & n14991 ;
  assign n21541 = \s14_data_i[11]_pad  & n14700 ;
  assign n21542 = ~n21540 & ~n21541 ;
  assign n21543 = n21539 & n21542 ;
  assign n21544 = n21536 & n21543 ;
  assign n21545 = \s0_data_i[11]_pad  & n14627 ;
  assign n21546 = \s13_data_i[11]_pad  & n14971 ;
  assign n21547 = \s11_data_i[11]_pad  & n14967 ;
  assign n21548 = ~n21546 & ~n21547 ;
  assign n21549 = ~n21545 & n21548 ;
  assign n21550 = \s6_data_i[11]_pad  & n14987 ;
  assign n21551 = \s4_data_i[11]_pad  & n14979 ;
  assign n21552 = ~n21550 & ~n21551 ;
  assign n21553 = \s9_data_i[11]_pad  & n14995 ;
  assign n21554 = \s10_data_i[11]_pad  & n14963 ;
  assign n21555 = ~n21553 & ~n21554 ;
  assign n21556 = n21552 & n21555 ;
  assign n21557 = n21549 & n21556 ;
  assign n21558 = n21544 & n21557 ;
  assign n21559 = n21529 & n21558 ;
  assign n21560 = n2203 & n15303 ;
  assign n21561 = \s15_data_i[12]_pad  & n2203 ;
  assign n21562 = ~n2258 & n21561 ;
  assign n21563 = ~n21560 & ~n21562 ;
  assign n21564 = \s12_data_i[12]_pad  & n14708 ;
  assign n21565 = \s1_data_i[12]_pad  & n14561 ;
  assign n21566 = ~n21564 & ~n21565 ;
  assign n21567 = \s0_data_i[12]_pad  & n14627 ;
  assign n21568 = \s10_data_i[12]_pad  & n14963 ;
  assign n21569 = ~n21567 & ~n21568 ;
  assign n21570 = n21566 & n21569 ;
  assign n21571 = \s3_data_i[12]_pad  & n14704 ;
  assign n21572 = \s4_data_i[12]_pad  & n14979 ;
  assign n21573 = ~n21571 & ~n21572 ;
  assign n21574 = \s9_data_i[12]_pad  & n14995 ;
  assign n21575 = \s6_data_i[12]_pad  & n14987 ;
  assign n21576 = ~n21574 & ~n21575 ;
  assign n21577 = n21573 & n21576 ;
  assign n21578 = n21570 & n21577 ;
  assign n21579 = \s14_data_i[12]_pad  & n14700 ;
  assign n21580 = \s11_data_i[12]_pad  & n14967 ;
  assign n21581 = \s7_data_i[12]_pad  & n14695 ;
  assign n21582 = ~n21580 & ~n21581 ;
  assign n21583 = ~n21579 & n21582 ;
  assign n21584 = \s5_data_i[12]_pad  & n14983 ;
  assign n21585 = \s8_data_i[12]_pad  & n14991 ;
  assign n21586 = ~n21584 & ~n21585 ;
  assign n21587 = \s2_data_i[12]_pad  & n14975 ;
  assign n21588 = \s13_data_i[12]_pad  & n14971 ;
  assign n21589 = ~n21587 & ~n21588 ;
  assign n21590 = n21586 & n21589 ;
  assign n21591 = n21583 & n21590 ;
  assign n21592 = n21578 & n21591 ;
  assign n21593 = n21563 & n21592 ;
  assign n21594 = n2203 & n15340 ;
  assign n21595 = \s15_data_i[13]_pad  & n2203 ;
  assign n21596 = ~n2258 & n21595 ;
  assign n21597 = ~n21594 & ~n21596 ;
  assign n21598 = \s12_data_i[13]_pad  & n14708 ;
  assign n21599 = \s1_data_i[13]_pad  & n14561 ;
  assign n21600 = ~n21598 & ~n21599 ;
  assign n21601 = \s0_data_i[13]_pad  & n14627 ;
  assign n21602 = \s10_data_i[13]_pad  & n14963 ;
  assign n21603 = ~n21601 & ~n21602 ;
  assign n21604 = n21600 & n21603 ;
  assign n21605 = \s3_data_i[13]_pad  & n14704 ;
  assign n21606 = \s4_data_i[13]_pad  & n14979 ;
  assign n21607 = ~n21605 & ~n21606 ;
  assign n21608 = \s9_data_i[13]_pad  & n14995 ;
  assign n21609 = \s6_data_i[13]_pad  & n14987 ;
  assign n21610 = ~n21608 & ~n21609 ;
  assign n21611 = n21607 & n21610 ;
  assign n21612 = n21604 & n21611 ;
  assign n21613 = \s14_data_i[13]_pad  & n14700 ;
  assign n21614 = \s11_data_i[13]_pad  & n14967 ;
  assign n21615 = \s7_data_i[13]_pad  & n14695 ;
  assign n21616 = ~n21614 & ~n21615 ;
  assign n21617 = ~n21613 & n21616 ;
  assign n21618 = \s5_data_i[13]_pad  & n14983 ;
  assign n21619 = \s8_data_i[13]_pad  & n14991 ;
  assign n21620 = ~n21618 & ~n21619 ;
  assign n21621 = \s2_data_i[13]_pad  & n14975 ;
  assign n21622 = \s13_data_i[13]_pad  & n14971 ;
  assign n21623 = ~n21621 & ~n21622 ;
  assign n21624 = n21620 & n21623 ;
  assign n21625 = n21617 & n21624 ;
  assign n21626 = n21612 & n21625 ;
  assign n21627 = n21597 & n21626 ;
  assign n21628 = n2203 & n15377 ;
  assign n21629 = \s15_data_i[14]_pad  & n2203 ;
  assign n21630 = ~n2258 & n21629 ;
  assign n21631 = ~n21628 & ~n21630 ;
  assign n21632 = \s12_data_i[14]_pad  & n14708 ;
  assign n21633 = \s1_data_i[14]_pad  & n14561 ;
  assign n21634 = ~n21632 & ~n21633 ;
  assign n21635 = \s0_data_i[14]_pad  & n14627 ;
  assign n21636 = \s10_data_i[14]_pad  & n14963 ;
  assign n21637 = ~n21635 & ~n21636 ;
  assign n21638 = n21634 & n21637 ;
  assign n21639 = \s3_data_i[14]_pad  & n14704 ;
  assign n21640 = \s4_data_i[14]_pad  & n14979 ;
  assign n21641 = ~n21639 & ~n21640 ;
  assign n21642 = \s9_data_i[14]_pad  & n14995 ;
  assign n21643 = \s6_data_i[14]_pad  & n14987 ;
  assign n21644 = ~n21642 & ~n21643 ;
  assign n21645 = n21641 & n21644 ;
  assign n21646 = n21638 & n21645 ;
  assign n21647 = \s14_data_i[14]_pad  & n14700 ;
  assign n21648 = \s11_data_i[14]_pad  & n14967 ;
  assign n21649 = \s7_data_i[14]_pad  & n14695 ;
  assign n21650 = ~n21648 & ~n21649 ;
  assign n21651 = ~n21647 & n21650 ;
  assign n21652 = \s5_data_i[14]_pad  & n14983 ;
  assign n21653 = \s8_data_i[14]_pad  & n14991 ;
  assign n21654 = ~n21652 & ~n21653 ;
  assign n21655 = \s2_data_i[14]_pad  & n14975 ;
  assign n21656 = \s13_data_i[14]_pad  & n14971 ;
  assign n21657 = ~n21655 & ~n21656 ;
  assign n21658 = n21654 & n21657 ;
  assign n21659 = n21651 & n21658 ;
  assign n21660 = n21646 & n21659 ;
  assign n21661 = n21631 & n21660 ;
  assign n21662 = n2203 & n15414 ;
  assign n21663 = \s15_data_i[15]_pad  & n2203 ;
  assign n21664 = ~n2258 & n21663 ;
  assign n21665 = ~n21662 & ~n21664 ;
  assign n21666 = \s12_data_i[15]_pad  & n14708 ;
  assign n21667 = \s1_data_i[15]_pad  & n14561 ;
  assign n21668 = ~n21666 & ~n21667 ;
  assign n21669 = \s0_data_i[15]_pad  & n14627 ;
  assign n21670 = \s10_data_i[15]_pad  & n14963 ;
  assign n21671 = ~n21669 & ~n21670 ;
  assign n21672 = n21668 & n21671 ;
  assign n21673 = \s3_data_i[15]_pad  & n14704 ;
  assign n21674 = \s4_data_i[15]_pad  & n14979 ;
  assign n21675 = ~n21673 & ~n21674 ;
  assign n21676 = \s9_data_i[15]_pad  & n14995 ;
  assign n21677 = \s6_data_i[15]_pad  & n14987 ;
  assign n21678 = ~n21676 & ~n21677 ;
  assign n21679 = n21675 & n21678 ;
  assign n21680 = n21672 & n21679 ;
  assign n21681 = \s14_data_i[15]_pad  & n14700 ;
  assign n21682 = \s11_data_i[15]_pad  & n14967 ;
  assign n21683 = \s7_data_i[15]_pad  & n14695 ;
  assign n21684 = ~n21682 & ~n21683 ;
  assign n21685 = ~n21681 & n21684 ;
  assign n21686 = \s5_data_i[15]_pad  & n14983 ;
  assign n21687 = \s8_data_i[15]_pad  & n14991 ;
  assign n21688 = ~n21686 & ~n21687 ;
  assign n21689 = \s2_data_i[15]_pad  & n14975 ;
  assign n21690 = \s13_data_i[15]_pad  & n14971 ;
  assign n21691 = ~n21689 & ~n21690 ;
  assign n21692 = n21688 & n21691 ;
  assign n21693 = n21685 & n21692 ;
  assign n21694 = n21680 & n21693 ;
  assign n21695 = n21665 & n21694 ;
  assign n21696 = \s15_data_i[16]_pad  & n2203 ;
  assign n21697 = ~n2258 & n21696 ;
  assign n21698 = \s8_data_i[16]_pad  & n14991 ;
  assign n21699 = \s1_data_i[16]_pad  & n14561 ;
  assign n21700 = ~n21698 & ~n21699 ;
  assign n21701 = \s4_data_i[16]_pad  & n14979 ;
  assign n21702 = \s6_data_i[16]_pad  & n14987 ;
  assign n21703 = ~n21701 & ~n21702 ;
  assign n21704 = n21700 & n21703 ;
  assign n21705 = \s3_data_i[16]_pad  & n14704 ;
  assign n21706 = \s9_data_i[16]_pad  & n14995 ;
  assign n21707 = ~n21705 & ~n21706 ;
  assign n21708 = \s10_data_i[16]_pad  & n14963 ;
  assign n21709 = \s7_data_i[16]_pad  & n14695 ;
  assign n21710 = ~n21708 & ~n21709 ;
  assign n21711 = n21707 & n21710 ;
  assign n21712 = n21704 & n21711 ;
  assign n21713 = \s11_data_i[16]_pad  & n14967 ;
  assign n21714 = \s14_data_i[16]_pad  & n14700 ;
  assign n21715 = \s2_data_i[16]_pad  & n14975 ;
  assign n21716 = ~n21714 & ~n21715 ;
  assign n21717 = ~n21713 & n21716 ;
  assign n21718 = \s5_data_i[16]_pad  & n14983 ;
  assign n21719 = \s12_data_i[16]_pad  & n14708 ;
  assign n21720 = ~n21718 & ~n21719 ;
  assign n21721 = \s13_data_i[16]_pad  & n14971 ;
  assign n21722 = \s0_data_i[16]_pad  & n14627 ;
  assign n21723 = ~n21721 & ~n21722 ;
  assign n21724 = n21720 & n21723 ;
  assign n21725 = n21717 & n21724 ;
  assign n21726 = n21712 & n21725 ;
  assign n21727 = ~n21697 & n21726 ;
  assign n21728 = \s15_data_i[17]_pad  & n2203 ;
  assign n21729 = ~n2258 & n21728 ;
  assign n21730 = \s8_data_i[17]_pad  & n14991 ;
  assign n21731 = \s1_data_i[17]_pad  & n14561 ;
  assign n21732 = ~n21730 & ~n21731 ;
  assign n21733 = \s4_data_i[17]_pad  & n14979 ;
  assign n21734 = \s6_data_i[17]_pad  & n14987 ;
  assign n21735 = ~n21733 & ~n21734 ;
  assign n21736 = n21732 & n21735 ;
  assign n21737 = \s3_data_i[17]_pad  & n14704 ;
  assign n21738 = \s9_data_i[17]_pad  & n14995 ;
  assign n21739 = ~n21737 & ~n21738 ;
  assign n21740 = \s10_data_i[17]_pad  & n14963 ;
  assign n21741 = \s7_data_i[17]_pad  & n14695 ;
  assign n21742 = ~n21740 & ~n21741 ;
  assign n21743 = n21739 & n21742 ;
  assign n21744 = n21736 & n21743 ;
  assign n21745 = \s11_data_i[17]_pad  & n14967 ;
  assign n21746 = \s14_data_i[17]_pad  & n14700 ;
  assign n21747 = \s2_data_i[17]_pad  & n14975 ;
  assign n21748 = ~n21746 & ~n21747 ;
  assign n21749 = ~n21745 & n21748 ;
  assign n21750 = \s5_data_i[17]_pad  & n14983 ;
  assign n21751 = \s12_data_i[17]_pad  & n14708 ;
  assign n21752 = ~n21750 & ~n21751 ;
  assign n21753 = \s13_data_i[17]_pad  & n14971 ;
  assign n21754 = \s0_data_i[17]_pad  & n14627 ;
  assign n21755 = ~n21753 & ~n21754 ;
  assign n21756 = n21752 & n21755 ;
  assign n21757 = n21749 & n21756 ;
  assign n21758 = n21744 & n21757 ;
  assign n21759 = ~n21729 & n21758 ;
  assign n21760 = \s15_data_i[18]_pad  & n2203 ;
  assign n21761 = ~n2258 & n21760 ;
  assign n21762 = \s8_data_i[18]_pad  & n14991 ;
  assign n21763 = \s1_data_i[18]_pad  & n14561 ;
  assign n21764 = ~n21762 & ~n21763 ;
  assign n21765 = \s4_data_i[18]_pad  & n14979 ;
  assign n21766 = \s6_data_i[18]_pad  & n14987 ;
  assign n21767 = ~n21765 & ~n21766 ;
  assign n21768 = n21764 & n21767 ;
  assign n21769 = \s3_data_i[18]_pad  & n14704 ;
  assign n21770 = \s9_data_i[18]_pad  & n14995 ;
  assign n21771 = ~n21769 & ~n21770 ;
  assign n21772 = \s10_data_i[18]_pad  & n14963 ;
  assign n21773 = \s7_data_i[18]_pad  & n14695 ;
  assign n21774 = ~n21772 & ~n21773 ;
  assign n21775 = n21771 & n21774 ;
  assign n21776 = n21768 & n21775 ;
  assign n21777 = \s11_data_i[18]_pad  & n14967 ;
  assign n21778 = \s14_data_i[18]_pad  & n14700 ;
  assign n21779 = \s2_data_i[18]_pad  & n14975 ;
  assign n21780 = ~n21778 & ~n21779 ;
  assign n21781 = ~n21777 & n21780 ;
  assign n21782 = \s5_data_i[18]_pad  & n14983 ;
  assign n21783 = \s12_data_i[18]_pad  & n14708 ;
  assign n21784 = ~n21782 & ~n21783 ;
  assign n21785 = \s13_data_i[18]_pad  & n14971 ;
  assign n21786 = \s0_data_i[18]_pad  & n14627 ;
  assign n21787 = ~n21785 & ~n21786 ;
  assign n21788 = n21784 & n21787 ;
  assign n21789 = n21781 & n21788 ;
  assign n21790 = n21776 & n21789 ;
  assign n21791 = ~n21761 & n21790 ;
  assign n21792 = \s15_data_i[19]_pad  & n2203 ;
  assign n21793 = ~n2258 & n21792 ;
  assign n21794 = \s8_data_i[19]_pad  & n14991 ;
  assign n21795 = \s1_data_i[19]_pad  & n14561 ;
  assign n21796 = ~n21794 & ~n21795 ;
  assign n21797 = \s4_data_i[19]_pad  & n14979 ;
  assign n21798 = \s6_data_i[19]_pad  & n14987 ;
  assign n21799 = ~n21797 & ~n21798 ;
  assign n21800 = n21796 & n21799 ;
  assign n21801 = \s3_data_i[19]_pad  & n14704 ;
  assign n21802 = \s9_data_i[19]_pad  & n14995 ;
  assign n21803 = ~n21801 & ~n21802 ;
  assign n21804 = \s10_data_i[19]_pad  & n14963 ;
  assign n21805 = \s7_data_i[19]_pad  & n14695 ;
  assign n21806 = ~n21804 & ~n21805 ;
  assign n21807 = n21803 & n21806 ;
  assign n21808 = n21800 & n21807 ;
  assign n21809 = \s11_data_i[19]_pad  & n14967 ;
  assign n21810 = \s14_data_i[19]_pad  & n14700 ;
  assign n21811 = \s2_data_i[19]_pad  & n14975 ;
  assign n21812 = ~n21810 & ~n21811 ;
  assign n21813 = ~n21809 & n21812 ;
  assign n21814 = \s5_data_i[19]_pad  & n14983 ;
  assign n21815 = \s12_data_i[19]_pad  & n14708 ;
  assign n21816 = ~n21814 & ~n21815 ;
  assign n21817 = \s13_data_i[19]_pad  & n14971 ;
  assign n21818 = \s0_data_i[19]_pad  & n14627 ;
  assign n21819 = ~n21817 & ~n21818 ;
  assign n21820 = n21816 & n21819 ;
  assign n21821 = n21813 & n21820 ;
  assign n21822 = n21808 & n21821 ;
  assign n21823 = ~n21793 & n21822 ;
  assign n21824 = n2203 & n15579 ;
  assign n21825 = \s15_data_i[1]_pad  & n2203 ;
  assign n21826 = ~n2258 & n21825 ;
  assign n21827 = ~n21824 & ~n21826 ;
  assign n21828 = \s12_data_i[1]_pad  & n14708 ;
  assign n21829 = \s1_data_i[1]_pad  & n14561 ;
  assign n21830 = ~n21828 & ~n21829 ;
  assign n21831 = \s0_data_i[1]_pad  & n14627 ;
  assign n21832 = \s10_data_i[1]_pad  & n14963 ;
  assign n21833 = ~n21831 & ~n21832 ;
  assign n21834 = n21830 & n21833 ;
  assign n21835 = \s3_data_i[1]_pad  & n14704 ;
  assign n21836 = \s4_data_i[1]_pad  & n14979 ;
  assign n21837 = ~n21835 & ~n21836 ;
  assign n21838 = \s9_data_i[1]_pad  & n14995 ;
  assign n21839 = \s6_data_i[1]_pad  & n14987 ;
  assign n21840 = ~n21838 & ~n21839 ;
  assign n21841 = n21837 & n21840 ;
  assign n21842 = n21834 & n21841 ;
  assign n21843 = \s14_data_i[1]_pad  & n14700 ;
  assign n21844 = \s11_data_i[1]_pad  & n14967 ;
  assign n21845 = \s7_data_i[1]_pad  & n14695 ;
  assign n21846 = ~n21844 & ~n21845 ;
  assign n21847 = ~n21843 & n21846 ;
  assign n21848 = \s5_data_i[1]_pad  & n14983 ;
  assign n21849 = \s8_data_i[1]_pad  & n14991 ;
  assign n21850 = ~n21848 & ~n21849 ;
  assign n21851 = \s2_data_i[1]_pad  & n14975 ;
  assign n21852 = \s13_data_i[1]_pad  & n14971 ;
  assign n21853 = ~n21851 & ~n21852 ;
  assign n21854 = n21850 & n21853 ;
  assign n21855 = n21847 & n21854 ;
  assign n21856 = n21842 & n21855 ;
  assign n21857 = n21827 & n21856 ;
  assign n21858 = \s15_data_i[20]_pad  & n2203 ;
  assign n21859 = ~n2258 & n21858 ;
  assign n21860 = \s8_data_i[20]_pad  & n14991 ;
  assign n21861 = \s1_data_i[20]_pad  & n14561 ;
  assign n21862 = ~n21860 & ~n21861 ;
  assign n21863 = \s4_data_i[20]_pad  & n14979 ;
  assign n21864 = \s6_data_i[20]_pad  & n14987 ;
  assign n21865 = ~n21863 & ~n21864 ;
  assign n21866 = n21862 & n21865 ;
  assign n21867 = \s3_data_i[20]_pad  & n14704 ;
  assign n21868 = \s9_data_i[20]_pad  & n14995 ;
  assign n21869 = ~n21867 & ~n21868 ;
  assign n21870 = \s10_data_i[20]_pad  & n14963 ;
  assign n21871 = \s7_data_i[20]_pad  & n14695 ;
  assign n21872 = ~n21870 & ~n21871 ;
  assign n21873 = n21869 & n21872 ;
  assign n21874 = n21866 & n21873 ;
  assign n21875 = \s11_data_i[20]_pad  & n14967 ;
  assign n21876 = \s14_data_i[20]_pad  & n14700 ;
  assign n21877 = \s2_data_i[20]_pad  & n14975 ;
  assign n21878 = ~n21876 & ~n21877 ;
  assign n21879 = ~n21875 & n21878 ;
  assign n21880 = \s5_data_i[20]_pad  & n14983 ;
  assign n21881 = \s12_data_i[20]_pad  & n14708 ;
  assign n21882 = ~n21880 & ~n21881 ;
  assign n21883 = \s13_data_i[20]_pad  & n14971 ;
  assign n21884 = \s0_data_i[20]_pad  & n14627 ;
  assign n21885 = ~n21883 & ~n21884 ;
  assign n21886 = n21882 & n21885 ;
  assign n21887 = n21879 & n21886 ;
  assign n21888 = n21874 & n21887 ;
  assign n21889 = ~n21859 & n21888 ;
  assign n21890 = \s15_data_i[21]_pad  & n2203 ;
  assign n21891 = ~n2258 & n21890 ;
  assign n21892 = \s8_data_i[21]_pad  & n14991 ;
  assign n21893 = \s1_data_i[21]_pad  & n14561 ;
  assign n21894 = ~n21892 & ~n21893 ;
  assign n21895 = \s4_data_i[21]_pad  & n14979 ;
  assign n21896 = \s6_data_i[21]_pad  & n14987 ;
  assign n21897 = ~n21895 & ~n21896 ;
  assign n21898 = n21894 & n21897 ;
  assign n21899 = \s3_data_i[21]_pad  & n14704 ;
  assign n21900 = \s9_data_i[21]_pad  & n14995 ;
  assign n21901 = ~n21899 & ~n21900 ;
  assign n21902 = \s10_data_i[21]_pad  & n14963 ;
  assign n21903 = \s7_data_i[21]_pad  & n14695 ;
  assign n21904 = ~n21902 & ~n21903 ;
  assign n21905 = n21901 & n21904 ;
  assign n21906 = n21898 & n21905 ;
  assign n21907 = \s11_data_i[21]_pad  & n14967 ;
  assign n21908 = \s14_data_i[21]_pad  & n14700 ;
  assign n21909 = \s2_data_i[21]_pad  & n14975 ;
  assign n21910 = ~n21908 & ~n21909 ;
  assign n21911 = ~n21907 & n21910 ;
  assign n21912 = \s5_data_i[21]_pad  & n14983 ;
  assign n21913 = \s12_data_i[21]_pad  & n14708 ;
  assign n21914 = ~n21912 & ~n21913 ;
  assign n21915 = \s13_data_i[21]_pad  & n14971 ;
  assign n21916 = \s0_data_i[21]_pad  & n14627 ;
  assign n21917 = ~n21915 & ~n21916 ;
  assign n21918 = n21914 & n21917 ;
  assign n21919 = n21911 & n21918 ;
  assign n21920 = n21906 & n21919 ;
  assign n21921 = ~n21891 & n21920 ;
  assign n21922 = \s15_data_i[22]_pad  & n2203 ;
  assign n21923 = ~n2258 & n21922 ;
  assign n21924 = \s8_data_i[22]_pad  & n14991 ;
  assign n21925 = \s1_data_i[22]_pad  & n14561 ;
  assign n21926 = ~n21924 & ~n21925 ;
  assign n21927 = \s4_data_i[22]_pad  & n14979 ;
  assign n21928 = \s6_data_i[22]_pad  & n14987 ;
  assign n21929 = ~n21927 & ~n21928 ;
  assign n21930 = n21926 & n21929 ;
  assign n21931 = \s3_data_i[22]_pad  & n14704 ;
  assign n21932 = \s9_data_i[22]_pad  & n14995 ;
  assign n21933 = ~n21931 & ~n21932 ;
  assign n21934 = \s10_data_i[22]_pad  & n14963 ;
  assign n21935 = \s7_data_i[22]_pad  & n14695 ;
  assign n21936 = ~n21934 & ~n21935 ;
  assign n21937 = n21933 & n21936 ;
  assign n21938 = n21930 & n21937 ;
  assign n21939 = \s11_data_i[22]_pad  & n14967 ;
  assign n21940 = \s14_data_i[22]_pad  & n14700 ;
  assign n21941 = \s2_data_i[22]_pad  & n14975 ;
  assign n21942 = ~n21940 & ~n21941 ;
  assign n21943 = ~n21939 & n21942 ;
  assign n21944 = \s5_data_i[22]_pad  & n14983 ;
  assign n21945 = \s12_data_i[22]_pad  & n14708 ;
  assign n21946 = ~n21944 & ~n21945 ;
  assign n21947 = \s13_data_i[22]_pad  & n14971 ;
  assign n21948 = \s0_data_i[22]_pad  & n14627 ;
  assign n21949 = ~n21947 & ~n21948 ;
  assign n21950 = n21946 & n21949 ;
  assign n21951 = n21943 & n21950 ;
  assign n21952 = n21938 & n21951 ;
  assign n21953 = ~n21923 & n21952 ;
  assign n21954 = \s15_data_i[23]_pad  & n2203 ;
  assign n21955 = ~n2258 & n21954 ;
  assign n21956 = \s8_data_i[23]_pad  & n14991 ;
  assign n21957 = \s1_data_i[23]_pad  & n14561 ;
  assign n21958 = ~n21956 & ~n21957 ;
  assign n21959 = \s4_data_i[23]_pad  & n14979 ;
  assign n21960 = \s6_data_i[23]_pad  & n14987 ;
  assign n21961 = ~n21959 & ~n21960 ;
  assign n21962 = n21958 & n21961 ;
  assign n21963 = \s3_data_i[23]_pad  & n14704 ;
  assign n21964 = \s9_data_i[23]_pad  & n14995 ;
  assign n21965 = ~n21963 & ~n21964 ;
  assign n21966 = \s10_data_i[23]_pad  & n14963 ;
  assign n21967 = \s7_data_i[23]_pad  & n14695 ;
  assign n21968 = ~n21966 & ~n21967 ;
  assign n21969 = n21965 & n21968 ;
  assign n21970 = n21962 & n21969 ;
  assign n21971 = \s11_data_i[23]_pad  & n14967 ;
  assign n21972 = \s14_data_i[23]_pad  & n14700 ;
  assign n21973 = \s2_data_i[23]_pad  & n14975 ;
  assign n21974 = ~n21972 & ~n21973 ;
  assign n21975 = ~n21971 & n21974 ;
  assign n21976 = \s5_data_i[23]_pad  & n14983 ;
  assign n21977 = \s12_data_i[23]_pad  & n14708 ;
  assign n21978 = ~n21976 & ~n21977 ;
  assign n21979 = \s13_data_i[23]_pad  & n14971 ;
  assign n21980 = \s0_data_i[23]_pad  & n14627 ;
  assign n21981 = ~n21979 & ~n21980 ;
  assign n21982 = n21978 & n21981 ;
  assign n21983 = n21975 & n21982 ;
  assign n21984 = n21970 & n21983 ;
  assign n21985 = ~n21955 & n21984 ;
  assign n21986 = \s15_data_i[24]_pad  & n2203 ;
  assign n21987 = ~n2258 & n21986 ;
  assign n21988 = \s8_data_i[24]_pad  & n14991 ;
  assign n21989 = \s1_data_i[24]_pad  & n14561 ;
  assign n21990 = ~n21988 & ~n21989 ;
  assign n21991 = \s4_data_i[24]_pad  & n14979 ;
  assign n21992 = \s6_data_i[24]_pad  & n14987 ;
  assign n21993 = ~n21991 & ~n21992 ;
  assign n21994 = n21990 & n21993 ;
  assign n21995 = \s3_data_i[24]_pad  & n14704 ;
  assign n21996 = \s9_data_i[24]_pad  & n14995 ;
  assign n21997 = ~n21995 & ~n21996 ;
  assign n21998 = \s10_data_i[24]_pad  & n14963 ;
  assign n21999 = \s7_data_i[24]_pad  & n14695 ;
  assign n22000 = ~n21998 & ~n21999 ;
  assign n22001 = n21997 & n22000 ;
  assign n22002 = n21994 & n22001 ;
  assign n22003 = \s11_data_i[24]_pad  & n14967 ;
  assign n22004 = \s14_data_i[24]_pad  & n14700 ;
  assign n22005 = \s2_data_i[24]_pad  & n14975 ;
  assign n22006 = ~n22004 & ~n22005 ;
  assign n22007 = ~n22003 & n22006 ;
  assign n22008 = \s5_data_i[24]_pad  & n14983 ;
  assign n22009 = \s12_data_i[24]_pad  & n14708 ;
  assign n22010 = ~n22008 & ~n22009 ;
  assign n22011 = \s13_data_i[24]_pad  & n14971 ;
  assign n22012 = \s0_data_i[24]_pad  & n14627 ;
  assign n22013 = ~n22011 & ~n22012 ;
  assign n22014 = n22010 & n22013 ;
  assign n22015 = n22007 & n22014 ;
  assign n22016 = n22002 & n22015 ;
  assign n22017 = ~n21987 & n22016 ;
  assign n22018 = \s15_data_i[25]_pad  & n2203 ;
  assign n22019 = ~n2258 & n22018 ;
  assign n22020 = \s8_data_i[25]_pad  & n14991 ;
  assign n22021 = \s1_data_i[25]_pad  & n14561 ;
  assign n22022 = ~n22020 & ~n22021 ;
  assign n22023 = \s4_data_i[25]_pad  & n14979 ;
  assign n22024 = \s6_data_i[25]_pad  & n14987 ;
  assign n22025 = ~n22023 & ~n22024 ;
  assign n22026 = n22022 & n22025 ;
  assign n22027 = \s3_data_i[25]_pad  & n14704 ;
  assign n22028 = \s9_data_i[25]_pad  & n14995 ;
  assign n22029 = ~n22027 & ~n22028 ;
  assign n22030 = \s10_data_i[25]_pad  & n14963 ;
  assign n22031 = \s7_data_i[25]_pad  & n14695 ;
  assign n22032 = ~n22030 & ~n22031 ;
  assign n22033 = n22029 & n22032 ;
  assign n22034 = n22026 & n22033 ;
  assign n22035 = \s11_data_i[25]_pad  & n14967 ;
  assign n22036 = \s14_data_i[25]_pad  & n14700 ;
  assign n22037 = \s2_data_i[25]_pad  & n14975 ;
  assign n22038 = ~n22036 & ~n22037 ;
  assign n22039 = ~n22035 & n22038 ;
  assign n22040 = \s5_data_i[25]_pad  & n14983 ;
  assign n22041 = \s12_data_i[25]_pad  & n14708 ;
  assign n22042 = ~n22040 & ~n22041 ;
  assign n22043 = \s13_data_i[25]_pad  & n14971 ;
  assign n22044 = \s0_data_i[25]_pad  & n14627 ;
  assign n22045 = ~n22043 & ~n22044 ;
  assign n22046 = n22042 & n22045 ;
  assign n22047 = n22039 & n22046 ;
  assign n22048 = n22034 & n22047 ;
  assign n22049 = ~n22019 & n22048 ;
  assign n22050 = \s15_data_i[26]_pad  & n2203 ;
  assign n22051 = ~n2258 & n22050 ;
  assign n22052 = \s8_data_i[26]_pad  & n14991 ;
  assign n22053 = \s1_data_i[26]_pad  & n14561 ;
  assign n22054 = ~n22052 & ~n22053 ;
  assign n22055 = \s4_data_i[26]_pad  & n14979 ;
  assign n22056 = \s6_data_i[26]_pad  & n14987 ;
  assign n22057 = ~n22055 & ~n22056 ;
  assign n22058 = n22054 & n22057 ;
  assign n22059 = \s3_data_i[26]_pad  & n14704 ;
  assign n22060 = \s9_data_i[26]_pad  & n14995 ;
  assign n22061 = ~n22059 & ~n22060 ;
  assign n22062 = \s10_data_i[26]_pad  & n14963 ;
  assign n22063 = \s7_data_i[26]_pad  & n14695 ;
  assign n22064 = ~n22062 & ~n22063 ;
  assign n22065 = n22061 & n22064 ;
  assign n22066 = n22058 & n22065 ;
  assign n22067 = \s11_data_i[26]_pad  & n14967 ;
  assign n22068 = \s14_data_i[26]_pad  & n14700 ;
  assign n22069 = \s2_data_i[26]_pad  & n14975 ;
  assign n22070 = ~n22068 & ~n22069 ;
  assign n22071 = ~n22067 & n22070 ;
  assign n22072 = \s5_data_i[26]_pad  & n14983 ;
  assign n22073 = \s12_data_i[26]_pad  & n14708 ;
  assign n22074 = ~n22072 & ~n22073 ;
  assign n22075 = \s13_data_i[26]_pad  & n14971 ;
  assign n22076 = \s0_data_i[26]_pad  & n14627 ;
  assign n22077 = ~n22075 & ~n22076 ;
  assign n22078 = n22074 & n22077 ;
  assign n22079 = n22071 & n22078 ;
  assign n22080 = n22066 & n22079 ;
  assign n22081 = ~n22051 & n22080 ;
  assign n22082 = \s15_data_i[27]_pad  & n2203 ;
  assign n22083 = ~n2258 & n22082 ;
  assign n22084 = \s8_data_i[27]_pad  & n14991 ;
  assign n22085 = \s1_data_i[27]_pad  & n14561 ;
  assign n22086 = ~n22084 & ~n22085 ;
  assign n22087 = \s4_data_i[27]_pad  & n14979 ;
  assign n22088 = \s6_data_i[27]_pad  & n14987 ;
  assign n22089 = ~n22087 & ~n22088 ;
  assign n22090 = n22086 & n22089 ;
  assign n22091 = \s3_data_i[27]_pad  & n14704 ;
  assign n22092 = \s9_data_i[27]_pad  & n14995 ;
  assign n22093 = ~n22091 & ~n22092 ;
  assign n22094 = \s10_data_i[27]_pad  & n14963 ;
  assign n22095 = \s7_data_i[27]_pad  & n14695 ;
  assign n22096 = ~n22094 & ~n22095 ;
  assign n22097 = n22093 & n22096 ;
  assign n22098 = n22090 & n22097 ;
  assign n22099 = \s11_data_i[27]_pad  & n14967 ;
  assign n22100 = \s14_data_i[27]_pad  & n14700 ;
  assign n22101 = \s2_data_i[27]_pad  & n14975 ;
  assign n22102 = ~n22100 & ~n22101 ;
  assign n22103 = ~n22099 & n22102 ;
  assign n22104 = \s5_data_i[27]_pad  & n14983 ;
  assign n22105 = \s12_data_i[27]_pad  & n14708 ;
  assign n22106 = ~n22104 & ~n22105 ;
  assign n22107 = \s13_data_i[27]_pad  & n14971 ;
  assign n22108 = \s0_data_i[27]_pad  & n14627 ;
  assign n22109 = ~n22107 & ~n22108 ;
  assign n22110 = n22106 & n22109 ;
  assign n22111 = n22103 & n22110 ;
  assign n22112 = n22098 & n22111 ;
  assign n22113 = ~n22083 & n22112 ;
  assign n22114 = \s15_data_i[28]_pad  & n2203 ;
  assign n22115 = ~n2258 & n22114 ;
  assign n22116 = \s8_data_i[28]_pad  & n14991 ;
  assign n22117 = \s1_data_i[28]_pad  & n14561 ;
  assign n22118 = ~n22116 & ~n22117 ;
  assign n22119 = \s4_data_i[28]_pad  & n14979 ;
  assign n22120 = \s6_data_i[28]_pad  & n14987 ;
  assign n22121 = ~n22119 & ~n22120 ;
  assign n22122 = n22118 & n22121 ;
  assign n22123 = \s3_data_i[28]_pad  & n14704 ;
  assign n22124 = \s9_data_i[28]_pad  & n14995 ;
  assign n22125 = ~n22123 & ~n22124 ;
  assign n22126 = \s10_data_i[28]_pad  & n14963 ;
  assign n22127 = \s7_data_i[28]_pad  & n14695 ;
  assign n22128 = ~n22126 & ~n22127 ;
  assign n22129 = n22125 & n22128 ;
  assign n22130 = n22122 & n22129 ;
  assign n22131 = \s11_data_i[28]_pad  & n14967 ;
  assign n22132 = \s14_data_i[28]_pad  & n14700 ;
  assign n22133 = \s2_data_i[28]_pad  & n14975 ;
  assign n22134 = ~n22132 & ~n22133 ;
  assign n22135 = ~n22131 & n22134 ;
  assign n22136 = \s5_data_i[28]_pad  & n14983 ;
  assign n22137 = \s12_data_i[28]_pad  & n14708 ;
  assign n22138 = ~n22136 & ~n22137 ;
  assign n22139 = \s13_data_i[28]_pad  & n14971 ;
  assign n22140 = \s0_data_i[28]_pad  & n14627 ;
  assign n22141 = ~n22139 & ~n22140 ;
  assign n22142 = n22138 & n22141 ;
  assign n22143 = n22135 & n22142 ;
  assign n22144 = n22130 & n22143 ;
  assign n22145 = ~n22115 & n22144 ;
  assign n22146 = \s15_data_i[29]_pad  & n2203 ;
  assign n22147 = ~n2258 & n22146 ;
  assign n22148 = \s8_data_i[29]_pad  & n14991 ;
  assign n22149 = \s1_data_i[29]_pad  & n14561 ;
  assign n22150 = ~n22148 & ~n22149 ;
  assign n22151 = \s4_data_i[29]_pad  & n14979 ;
  assign n22152 = \s6_data_i[29]_pad  & n14987 ;
  assign n22153 = ~n22151 & ~n22152 ;
  assign n22154 = n22150 & n22153 ;
  assign n22155 = \s3_data_i[29]_pad  & n14704 ;
  assign n22156 = \s9_data_i[29]_pad  & n14995 ;
  assign n22157 = ~n22155 & ~n22156 ;
  assign n22158 = \s10_data_i[29]_pad  & n14963 ;
  assign n22159 = \s7_data_i[29]_pad  & n14695 ;
  assign n22160 = ~n22158 & ~n22159 ;
  assign n22161 = n22157 & n22160 ;
  assign n22162 = n22154 & n22161 ;
  assign n22163 = \s11_data_i[29]_pad  & n14967 ;
  assign n22164 = \s14_data_i[29]_pad  & n14700 ;
  assign n22165 = \s2_data_i[29]_pad  & n14975 ;
  assign n22166 = ~n22164 & ~n22165 ;
  assign n22167 = ~n22163 & n22166 ;
  assign n22168 = \s5_data_i[29]_pad  & n14983 ;
  assign n22169 = \s12_data_i[29]_pad  & n14708 ;
  assign n22170 = ~n22168 & ~n22169 ;
  assign n22171 = \s13_data_i[29]_pad  & n14971 ;
  assign n22172 = \s0_data_i[29]_pad  & n14627 ;
  assign n22173 = ~n22171 & ~n22172 ;
  assign n22174 = n22170 & n22173 ;
  assign n22175 = n22167 & n22174 ;
  assign n22176 = n22162 & n22175 ;
  assign n22177 = ~n22147 & n22176 ;
  assign n22178 = n2203 & n15936 ;
  assign n22179 = \s15_data_i[2]_pad  & n2203 ;
  assign n22180 = ~n2258 & n22179 ;
  assign n22181 = ~n22178 & ~n22180 ;
  assign n22182 = \s12_data_i[2]_pad  & n14708 ;
  assign n22183 = \s1_data_i[2]_pad  & n14561 ;
  assign n22184 = ~n22182 & ~n22183 ;
  assign n22185 = \s0_data_i[2]_pad  & n14627 ;
  assign n22186 = \s10_data_i[2]_pad  & n14963 ;
  assign n22187 = ~n22185 & ~n22186 ;
  assign n22188 = n22184 & n22187 ;
  assign n22189 = \s3_data_i[2]_pad  & n14704 ;
  assign n22190 = \s4_data_i[2]_pad  & n14979 ;
  assign n22191 = ~n22189 & ~n22190 ;
  assign n22192 = \s9_data_i[2]_pad  & n14995 ;
  assign n22193 = \s6_data_i[2]_pad  & n14987 ;
  assign n22194 = ~n22192 & ~n22193 ;
  assign n22195 = n22191 & n22194 ;
  assign n22196 = n22188 & n22195 ;
  assign n22197 = \s14_data_i[2]_pad  & n14700 ;
  assign n22198 = \s11_data_i[2]_pad  & n14967 ;
  assign n22199 = \s7_data_i[2]_pad  & n14695 ;
  assign n22200 = ~n22198 & ~n22199 ;
  assign n22201 = ~n22197 & n22200 ;
  assign n22202 = \s5_data_i[2]_pad  & n14983 ;
  assign n22203 = \s8_data_i[2]_pad  & n14991 ;
  assign n22204 = ~n22202 & ~n22203 ;
  assign n22205 = \s2_data_i[2]_pad  & n14975 ;
  assign n22206 = \s13_data_i[2]_pad  & n14971 ;
  assign n22207 = ~n22205 & ~n22206 ;
  assign n22208 = n22204 & n22207 ;
  assign n22209 = n22201 & n22208 ;
  assign n22210 = n22196 & n22209 ;
  assign n22211 = n22181 & n22210 ;
  assign n22212 = \s15_data_i[30]_pad  & n2203 ;
  assign n22213 = ~n2258 & n22212 ;
  assign n22214 = \s8_data_i[30]_pad  & n14991 ;
  assign n22215 = \s1_data_i[30]_pad  & n14561 ;
  assign n22216 = ~n22214 & ~n22215 ;
  assign n22217 = \s4_data_i[30]_pad  & n14979 ;
  assign n22218 = \s6_data_i[30]_pad  & n14987 ;
  assign n22219 = ~n22217 & ~n22218 ;
  assign n22220 = n22216 & n22219 ;
  assign n22221 = \s3_data_i[30]_pad  & n14704 ;
  assign n22222 = \s9_data_i[30]_pad  & n14995 ;
  assign n22223 = ~n22221 & ~n22222 ;
  assign n22224 = \s10_data_i[30]_pad  & n14963 ;
  assign n22225 = \s7_data_i[30]_pad  & n14695 ;
  assign n22226 = ~n22224 & ~n22225 ;
  assign n22227 = n22223 & n22226 ;
  assign n22228 = n22220 & n22227 ;
  assign n22229 = \s11_data_i[30]_pad  & n14967 ;
  assign n22230 = \s14_data_i[30]_pad  & n14700 ;
  assign n22231 = \s2_data_i[30]_pad  & n14975 ;
  assign n22232 = ~n22230 & ~n22231 ;
  assign n22233 = ~n22229 & n22232 ;
  assign n22234 = \s5_data_i[30]_pad  & n14983 ;
  assign n22235 = \s12_data_i[30]_pad  & n14708 ;
  assign n22236 = ~n22234 & ~n22235 ;
  assign n22237 = \s13_data_i[30]_pad  & n14971 ;
  assign n22238 = \s0_data_i[30]_pad  & n14627 ;
  assign n22239 = ~n22237 & ~n22238 ;
  assign n22240 = n22236 & n22239 ;
  assign n22241 = n22233 & n22240 ;
  assign n22242 = n22228 & n22241 ;
  assign n22243 = ~n22213 & n22242 ;
  assign n22244 = \s15_data_i[31]_pad  & n2203 ;
  assign n22245 = ~n2258 & n22244 ;
  assign n22246 = \s8_data_i[31]_pad  & n14991 ;
  assign n22247 = \s1_data_i[31]_pad  & n14561 ;
  assign n22248 = ~n22246 & ~n22247 ;
  assign n22249 = \s4_data_i[31]_pad  & n14979 ;
  assign n22250 = \s6_data_i[31]_pad  & n14987 ;
  assign n22251 = ~n22249 & ~n22250 ;
  assign n22252 = n22248 & n22251 ;
  assign n22253 = \s3_data_i[31]_pad  & n14704 ;
  assign n22254 = \s9_data_i[31]_pad  & n14995 ;
  assign n22255 = ~n22253 & ~n22254 ;
  assign n22256 = \s10_data_i[31]_pad  & n14963 ;
  assign n22257 = \s7_data_i[31]_pad  & n14695 ;
  assign n22258 = ~n22256 & ~n22257 ;
  assign n22259 = n22255 & n22258 ;
  assign n22260 = n22252 & n22259 ;
  assign n22261 = \s11_data_i[31]_pad  & n14967 ;
  assign n22262 = \s14_data_i[31]_pad  & n14700 ;
  assign n22263 = \s2_data_i[31]_pad  & n14975 ;
  assign n22264 = ~n22262 & ~n22263 ;
  assign n22265 = ~n22261 & n22264 ;
  assign n22266 = \s5_data_i[31]_pad  & n14983 ;
  assign n22267 = \s12_data_i[31]_pad  & n14708 ;
  assign n22268 = ~n22266 & ~n22267 ;
  assign n22269 = \s13_data_i[31]_pad  & n14971 ;
  assign n22270 = \s0_data_i[31]_pad  & n14627 ;
  assign n22271 = ~n22269 & ~n22270 ;
  assign n22272 = n22268 & n22271 ;
  assign n22273 = n22265 & n22272 ;
  assign n22274 = n22260 & n22273 ;
  assign n22275 = ~n22245 & n22274 ;
  assign n22276 = n2203 & n16037 ;
  assign n22277 = \s15_data_i[3]_pad  & n2203 ;
  assign n22278 = ~n2258 & n22277 ;
  assign n22279 = ~n22276 & ~n22278 ;
  assign n22280 = \s12_data_i[3]_pad  & n14708 ;
  assign n22281 = \s1_data_i[3]_pad  & n14561 ;
  assign n22282 = ~n22280 & ~n22281 ;
  assign n22283 = \s4_data_i[3]_pad  & n14979 ;
  assign n22284 = \s6_data_i[3]_pad  & n14987 ;
  assign n22285 = ~n22283 & ~n22284 ;
  assign n22286 = n22282 & n22285 ;
  assign n22287 = \s3_data_i[3]_pad  & n14704 ;
  assign n22288 = \s9_data_i[3]_pad  & n14995 ;
  assign n22289 = ~n22287 & ~n22288 ;
  assign n22290 = \s10_data_i[3]_pad  & n14963 ;
  assign n22291 = \s7_data_i[3]_pad  & n14695 ;
  assign n22292 = ~n22290 & ~n22291 ;
  assign n22293 = n22289 & n22292 ;
  assign n22294 = n22286 & n22293 ;
  assign n22295 = \s14_data_i[3]_pad  & n14700 ;
  assign n22296 = \s11_data_i[3]_pad  & n14967 ;
  assign n22297 = \s2_data_i[3]_pad  & n14975 ;
  assign n22298 = ~n22296 & ~n22297 ;
  assign n22299 = ~n22295 & n22298 ;
  assign n22300 = \s5_data_i[3]_pad  & n14983 ;
  assign n22301 = \s8_data_i[3]_pad  & n14991 ;
  assign n22302 = ~n22300 & ~n22301 ;
  assign n22303 = \s13_data_i[3]_pad  & n14971 ;
  assign n22304 = \s0_data_i[3]_pad  & n14627 ;
  assign n22305 = ~n22303 & ~n22304 ;
  assign n22306 = n22302 & n22305 ;
  assign n22307 = n22299 & n22306 ;
  assign n22308 = n22294 & n22307 ;
  assign n22309 = n22279 & n22308 ;
  assign n22310 = n2203 & n16074 ;
  assign n22311 = \s15_data_i[4]_pad  & n2203 ;
  assign n22312 = ~n2258 & n22311 ;
  assign n22313 = ~n22310 & ~n22312 ;
  assign n22314 = \s12_data_i[4]_pad  & n14708 ;
  assign n22315 = \s1_data_i[4]_pad  & n14561 ;
  assign n22316 = ~n22314 & ~n22315 ;
  assign n22317 = \s0_data_i[4]_pad  & n14627 ;
  assign n22318 = \s10_data_i[4]_pad  & n14963 ;
  assign n22319 = ~n22317 & ~n22318 ;
  assign n22320 = n22316 & n22319 ;
  assign n22321 = \s3_data_i[4]_pad  & n14704 ;
  assign n22322 = \s4_data_i[4]_pad  & n14979 ;
  assign n22323 = ~n22321 & ~n22322 ;
  assign n22324 = \s9_data_i[4]_pad  & n14995 ;
  assign n22325 = \s6_data_i[4]_pad  & n14987 ;
  assign n22326 = ~n22324 & ~n22325 ;
  assign n22327 = n22323 & n22326 ;
  assign n22328 = n22320 & n22327 ;
  assign n22329 = \s14_data_i[4]_pad  & n14700 ;
  assign n22330 = \s11_data_i[4]_pad  & n14967 ;
  assign n22331 = \s7_data_i[4]_pad  & n14695 ;
  assign n22332 = ~n22330 & ~n22331 ;
  assign n22333 = ~n22329 & n22332 ;
  assign n22334 = \s5_data_i[4]_pad  & n14983 ;
  assign n22335 = \s8_data_i[4]_pad  & n14991 ;
  assign n22336 = ~n22334 & ~n22335 ;
  assign n22337 = \s2_data_i[4]_pad  & n14975 ;
  assign n22338 = \s13_data_i[4]_pad  & n14971 ;
  assign n22339 = ~n22337 & ~n22338 ;
  assign n22340 = n22336 & n22339 ;
  assign n22341 = n22333 & n22340 ;
  assign n22342 = n22328 & n22341 ;
  assign n22343 = n22313 & n22342 ;
  assign n22344 = n2203 & n16111 ;
  assign n22345 = \s15_data_i[5]_pad  & n2203 ;
  assign n22346 = ~n2258 & n22345 ;
  assign n22347 = ~n22344 & ~n22346 ;
  assign n22348 = \s12_data_i[5]_pad  & n14708 ;
  assign n22349 = \s1_data_i[5]_pad  & n14561 ;
  assign n22350 = ~n22348 & ~n22349 ;
  assign n22351 = \s7_data_i[5]_pad  & n14695 ;
  assign n22352 = \s9_data_i[5]_pad  & n14995 ;
  assign n22353 = ~n22351 & ~n22352 ;
  assign n22354 = n22350 & n22353 ;
  assign n22355 = \s3_data_i[5]_pad  & n14704 ;
  assign n22356 = \s6_data_i[5]_pad  & n14987 ;
  assign n22357 = ~n22355 & ~n22356 ;
  assign n22358 = \s10_data_i[5]_pad  & n14963 ;
  assign n22359 = \s13_data_i[5]_pad  & n14971 ;
  assign n22360 = ~n22358 & ~n22359 ;
  assign n22361 = n22357 & n22360 ;
  assign n22362 = n22354 & n22361 ;
  assign n22363 = \s14_data_i[5]_pad  & n14700 ;
  assign n22364 = \s11_data_i[5]_pad  & n14967 ;
  assign n22365 = \s2_data_i[5]_pad  & n14975 ;
  assign n22366 = ~n22364 & ~n22365 ;
  assign n22367 = ~n22363 & n22366 ;
  assign n22368 = \s5_data_i[5]_pad  & n14983 ;
  assign n22369 = \s8_data_i[5]_pad  & n14991 ;
  assign n22370 = ~n22368 & ~n22369 ;
  assign n22371 = \s4_data_i[5]_pad  & n14979 ;
  assign n22372 = \s0_data_i[5]_pad  & n14627 ;
  assign n22373 = ~n22371 & ~n22372 ;
  assign n22374 = n22370 & n22373 ;
  assign n22375 = n22367 & n22374 ;
  assign n22376 = n22362 & n22375 ;
  assign n22377 = n22347 & n22376 ;
  assign n22378 = n2203 & n16148 ;
  assign n22379 = \s15_data_i[6]_pad  & n2203 ;
  assign n22380 = ~n2258 & n22379 ;
  assign n22381 = ~n22378 & ~n22380 ;
  assign n22382 = \s12_data_i[6]_pad  & n14708 ;
  assign n22383 = \s1_data_i[6]_pad  & n14561 ;
  assign n22384 = ~n22382 & ~n22383 ;
  assign n22385 = \s0_data_i[6]_pad  & n14627 ;
  assign n22386 = \s10_data_i[6]_pad  & n14963 ;
  assign n22387 = ~n22385 & ~n22386 ;
  assign n22388 = n22384 & n22387 ;
  assign n22389 = \s3_data_i[6]_pad  & n14704 ;
  assign n22390 = \s4_data_i[6]_pad  & n14979 ;
  assign n22391 = ~n22389 & ~n22390 ;
  assign n22392 = \s9_data_i[6]_pad  & n14995 ;
  assign n22393 = \s6_data_i[6]_pad  & n14987 ;
  assign n22394 = ~n22392 & ~n22393 ;
  assign n22395 = n22391 & n22394 ;
  assign n22396 = n22388 & n22395 ;
  assign n22397 = \s14_data_i[6]_pad  & n14700 ;
  assign n22398 = \s11_data_i[6]_pad  & n14967 ;
  assign n22399 = \s7_data_i[6]_pad  & n14695 ;
  assign n22400 = ~n22398 & ~n22399 ;
  assign n22401 = ~n22397 & n22400 ;
  assign n22402 = \s5_data_i[6]_pad  & n14983 ;
  assign n22403 = \s8_data_i[6]_pad  & n14991 ;
  assign n22404 = ~n22402 & ~n22403 ;
  assign n22405 = \s2_data_i[6]_pad  & n14975 ;
  assign n22406 = \s13_data_i[6]_pad  & n14971 ;
  assign n22407 = ~n22405 & ~n22406 ;
  assign n22408 = n22404 & n22407 ;
  assign n22409 = n22401 & n22408 ;
  assign n22410 = n22396 & n22409 ;
  assign n22411 = n22381 & n22410 ;
  assign n22412 = n2203 & n16185 ;
  assign n22413 = \s15_data_i[7]_pad  & n2203 ;
  assign n22414 = ~n2258 & n22413 ;
  assign n22415 = ~n22412 & ~n22414 ;
  assign n22416 = \s12_data_i[7]_pad  & n14708 ;
  assign n22417 = \s1_data_i[7]_pad  & n14561 ;
  assign n22418 = ~n22416 & ~n22417 ;
  assign n22419 = \s0_data_i[7]_pad  & n14627 ;
  assign n22420 = \s10_data_i[7]_pad  & n14963 ;
  assign n22421 = ~n22419 & ~n22420 ;
  assign n22422 = n22418 & n22421 ;
  assign n22423 = \s3_data_i[7]_pad  & n14704 ;
  assign n22424 = \s4_data_i[7]_pad  & n14979 ;
  assign n22425 = ~n22423 & ~n22424 ;
  assign n22426 = \s9_data_i[7]_pad  & n14995 ;
  assign n22427 = \s6_data_i[7]_pad  & n14987 ;
  assign n22428 = ~n22426 & ~n22427 ;
  assign n22429 = n22425 & n22428 ;
  assign n22430 = n22422 & n22429 ;
  assign n22431 = \s14_data_i[7]_pad  & n14700 ;
  assign n22432 = \s11_data_i[7]_pad  & n14967 ;
  assign n22433 = \s7_data_i[7]_pad  & n14695 ;
  assign n22434 = ~n22432 & ~n22433 ;
  assign n22435 = ~n22431 & n22434 ;
  assign n22436 = \s5_data_i[7]_pad  & n14983 ;
  assign n22437 = \s8_data_i[7]_pad  & n14991 ;
  assign n22438 = ~n22436 & ~n22437 ;
  assign n22439 = \s2_data_i[7]_pad  & n14975 ;
  assign n22440 = \s13_data_i[7]_pad  & n14971 ;
  assign n22441 = ~n22439 & ~n22440 ;
  assign n22442 = n22438 & n22441 ;
  assign n22443 = n22435 & n22442 ;
  assign n22444 = n22430 & n22443 ;
  assign n22445 = n22415 & n22444 ;
  assign n22446 = n2203 & n16222 ;
  assign n22447 = \s15_data_i[8]_pad  & n2203 ;
  assign n22448 = ~n2258 & n22447 ;
  assign n22449 = ~n22446 & ~n22448 ;
  assign n22450 = \s12_data_i[8]_pad  & n14708 ;
  assign n22451 = \s1_data_i[8]_pad  & n14561 ;
  assign n22452 = ~n22450 & ~n22451 ;
  assign n22453 = \s0_data_i[8]_pad  & n14627 ;
  assign n22454 = \s10_data_i[8]_pad  & n14963 ;
  assign n22455 = ~n22453 & ~n22454 ;
  assign n22456 = n22452 & n22455 ;
  assign n22457 = \s3_data_i[8]_pad  & n14704 ;
  assign n22458 = \s4_data_i[8]_pad  & n14979 ;
  assign n22459 = ~n22457 & ~n22458 ;
  assign n22460 = \s9_data_i[8]_pad  & n14995 ;
  assign n22461 = \s6_data_i[8]_pad  & n14987 ;
  assign n22462 = ~n22460 & ~n22461 ;
  assign n22463 = n22459 & n22462 ;
  assign n22464 = n22456 & n22463 ;
  assign n22465 = \s14_data_i[8]_pad  & n14700 ;
  assign n22466 = \s11_data_i[8]_pad  & n14967 ;
  assign n22467 = \s7_data_i[8]_pad  & n14695 ;
  assign n22468 = ~n22466 & ~n22467 ;
  assign n22469 = ~n22465 & n22468 ;
  assign n22470 = \s5_data_i[8]_pad  & n14983 ;
  assign n22471 = \s8_data_i[8]_pad  & n14991 ;
  assign n22472 = ~n22470 & ~n22471 ;
  assign n22473 = \s2_data_i[8]_pad  & n14975 ;
  assign n22474 = \s13_data_i[8]_pad  & n14971 ;
  assign n22475 = ~n22473 & ~n22474 ;
  assign n22476 = n22472 & n22475 ;
  assign n22477 = n22469 & n22476 ;
  assign n22478 = n22464 & n22477 ;
  assign n22479 = n22449 & n22478 ;
  assign n22480 = n2203 & n16259 ;
  assign n22481 = \s15_data_i[9]_pad  & n2203 ;
  assign n22482 = ~n2258 & n22481 ;
  assign n22483 = ~n22480 & ~n22482 ;
  assign n22484 = \s12_data_i[9]_pad  & n14708 ;
  assign n22485 = \s1_data_i[9]_pad  & n14561 ;
  assign n22486 = ~n22484 & ~n22485 ;
  assign n22487 = \s0_data_i[9]_pad  & n14627 ;
  assign n22488 = \s10_data_i[9]_pad  & n14963 ;
  assign n22489 = ~n22487 & ~n22488 ;
  assign n22490 = n22486 & n22489 ;
  assign n22491 = \s3_data_i[9]_pad  & n14704 ;
  assign n22492 = \s4_data_i[9]_pad  & n14979 ;
  assign n22493 = ~n22491 & ~n22492 ;
  assign n22494 = \s9_data_i[9]_pad  & n14995 ;
  assign n22495 = \s6_data_i[9]_pad  & n14987 ;
  assign n22496 = ~n22494 & ~n22495 ;
  assign n22497 = n22493 & n22496 ;
  assign n22498 = n22490 & n22497 ;
  assign n22499 = \s14_data_i[9]_pad  & n14700 ;
  assign n22500 = \s11_data_i[9]_pad  & n14967 ;
  assign n22501 = \s7_data_i[9]_pad  & n14695 ;
  assign n22502 = ~n22500 & ~n22501 ;
  assign n22503 = ~n22499 & n22502 ;
  assign n22504 = \s5_data_i[9]_pad  & n14983 ;
  assign n22505 = \s8_data_i[9]_pad  & n14991 ;
  assign n22506 = ~n22504 & ~n22505 ;
  assign n22507 = \s2_data_i[9]_pad  & n14975 ;
  assign n22508 = \s13_data_i[9]_pad  & n14971 ;
  assign n22509 = ~n22507 & ~n22508 ;
  assign n22510 = n22506 & n22509 ;
  assign n22511 = n22503 & n22510 ;
  assign n22512 = n22498 & n22511 ;
  assign n22513 = n22483 & n22512 ;
  assign n22514 = \s15_err_i_pad  & n21395 ;
  assign n22515 = ~n2258 & n22514 ;
  assign n22516 = \s6_err_i_pad  & n14987 ;
  assign n22517 = ~n13627 & n22516 ;
  assign n22518 = n13652 & n22517 ;
  assign n22519 = \s1_err_i_pad  & n14561 ;
  assign n22520 = ~n14271 & n22519 ;
  assign n22521 = n14288 & n22520 ;
  assign n22522 = ~n22518 & ~n22521 ;
  assign n22523 = \s12_err_i_pad  & n14708 ;
  assign n22524 = ~n14140 & n22523 ;
  assign n22525 = n14157 & n22524 ;
  assign n22526 = \s13_err_i_pad  & n14971 ;
  assign n22527 = ~n14211 & n22526 ;
  assign n22528 = n14236 & n22527 ;
  assign n22529 = ~n22525 & ~n22528 ;
  assign n22530 = n22522 & n22529 ;
  assign n22531 = \s10_err_i_pad  & n14963 ;
  assign n22532 = ~n13928 & n22531 ;
  assign n22533 = n13953 & n22532 ;
  assign n22534 = \s5_err_i_pad  & n14983 ;
  assign n22535 = ~n13547 & n22534 ;
  assign n22536 = n13555 & n22535 ;
  assign n22537 = ~n22533 & ~n22536 ;
  assign n22538 = \s8_err_i_pad  & n14991 ;
  assign n22539 = ~n13767 & n22538 ;
  assign n22540 = n13792 & n22539 ;
  assign n22541 = \s0_err_i_pad  & n14627 ;
  assign n22542 = ~n14069 & n22541 ;
  assign n22543 = n14077 & n22542 ;
  assign n22544 = ~n22540 & ~n22543 ;
  assign n22545 = n22537 & n22544 ;
  assign n22546 = n22530 & n22545 ;
  assign n22547 = \s7_err_i_pad  & n14695 ;
  assign n22548 = ~n13697 & n22547 ;
  assign n22549 = n13722 & n22548 ;
  assign n22550 = \s2_err_i_pad  & n14975 ;
  assign n22551 = ~n14391 & n22550 ;
  assign n22552 = n14384 & n22551 ;
  assign n22553 = \s4_err_i_pad  & n14979 ;
  assign n22554 = ~n13467 & n22553 ;
  assign n22555 = n13460 & n22554 ;
  assign n22556 = ~n22552 & ~n22555 ;
  assign n22557 = ~n22549 & n22556 ;
  assign n22558 = \s9_err_i_pad  & n14995 ;
  assign n22559 = ~n13847 & n22558 ;
  assign n22560 = n13872 & n22559 ;
  assign n22561 = \s3_err_i_pad  & n14704 ;
  assign n22562 = ~n14451 & n22561 ;
  assign n22563 = n14444 & n22562 ;
  assign n22564 = ~n22560 & ~n22563 ;
  assign n22565 = \s11_err_i_pad  & n14967 ;
  assign n22566 = ~n14009 & n22565 ;
  assign n22567 = n14002 & n22566 ;
  assign n22568 = \s14_err_i_pad  & n14700 ;
  assign n22569 = ~n14331 & n22568 ;
  assign n22570 = n14356 & n22569 ;
  assign n22571 = ~n22567 & ~n22570 ;
  assign n22572 = n22564 & n22571 ;
  assign n22573 = n22557 & n22572 ;
  assign n22574 = n22546 & n22573 ;
  assign n22575 = ~n22515 & n22574 ;
  assign n22576 = \s15_rty_i_pad  & n21395 ;
  assign n22577 = ~n2258 & n22576 ;
  assign n22578 = \s14_rty_i_pad  & n14700 ;
  assign n22579 = ~n14331 & n22578 ;
  assign n22580 = n14356 & n22579 ;
  assign n22581 = \s1_rty_i_pad  & n14561 ;
  assign n22582 = ~n14271 & n22581 ;
  assign n22583 = n14288 & n22582 ;
  assign n22584 = ~n22580 & ~n22583 ;
  assign n22585 = \s13_rty_i_pad  & n14971 ;
  assign n22586 = ~n14211 & n22585 ;
  assign n22587 = n14236 & n22586 ;
  assign n22588 = \s9_rty_i_pad  & n14995 ;
  assign n22589 = ~n13847 & n22588 ;
  assign n22590 = n13872 & n22589 ;
  assign n22591 = ~n22587 & ~n22590 ;
  assign n22592 = n22584 & n22591 ;
  assign n22593 = \s0_rty_i_pad  & n14627 ;
  assign n22594 = ~n14069 & n22593 ;
  assign n22595 = n14077 & n22594 ;
  assign n22596 = \s6_rty_i_pad  & n14987 ;
  assign n22597 = ~n13627 & n22596 ;
  assign n22598 = n13652 & n22597 ;
  assign n22599 = ~n22595 & ~n22598 ;
  assign n22600 = \s7_rty_i_pad  & n14695 ;
  assign n22601 = ~n13697 & n22600 ;
  assign n22602 = n13722 & n22601 ;
  assign n22603 = \s10_rty_i_pad  & n14963 ;
  assign n22604 = ~n13928 & n22603 ;
  assign n22605 = n13953 & n22604 ;
  assign n22606 = ~n22602 & ~n22605 ;
  assign n22607 = n22599 & n22606 ;
  assign n22608 = n22592 & n22607 ;
  assign n22609 = \s12_rty_i_pad  & n14708 ;
  assign n22610 = ~n14140 & n22609 ;
  assign n22611 = n14157 & n22610 ;
  assign n22612 = \s11_rty_i_pad  & n14967 ;
  assign n22613 = ~n14009 & n22612 ;
  assign n22614 = n14002 & n22613 ;
  assign n22615 = \s4_rty_i_pad  & n14979 ;
  assign n22616 = ~n13467 & n22615 ;
  assign n22617 = n13460 & n22616 ;
  assign n22618 = ~n22614 & ~n22617 ;
  assign n22619 = ~n22611 & n22618 ;
  assign n22620 = \s3_rty_i_pad  & n14704 ;
  assign n22621 = ~n14451 & n22620 ;
  assign n22622 = n14444 & n22621 ;
  assign n22623 = \s5_rty_i_pad  & n14983 ;
  assign n22624 = ~n13547 & n22623 ;
  assign n22625 = n13555 & n22624 ;
  assign n22626 = ~n22622 & ~n22625 ;
  assign n22627 = \s2_rty_i_pad  & n14975 ;
  assign n22628 = ~n14391 & n22627 ;
  assign n22629 = n14384 & n22628 ;
  assign n22630 = \s8_rty_i_pad  & n14991 ;
  assign n22631 = ~n13767 & n22630 ;
  assign n22632 = n13792 & n22631 ;
  assign n22633 = ~n22629 & ~n22632 ;
  assign n22634 = n22626 & n22633 ;
  assign n22635 = n22619 & n22634 ;
  assign n22636 = n22608 & n22635 ;
  assign n22637 = ~n22577 & n22636 ;
  assign n22638 = ~n1925 & n2176 ;
  assign n22639 = n1918 & n22638 ;
  assign n22640 = ~n13416 & n22639 ;
  assign n22641 = ~n15125 & n22640 ;
  assign n22642 = \s5_ack_i_pad  & n15034 ;
  assign n22643 = n13547 & n22642 ;
  assign n22644 = n13564 & n22643 ;
  assign n22645 = \s1_ack_i_pad  & n14640 ;
  assign n22646 = n14271 & n22645 ;
  assign n22647 = n14264 & n22646 ;
  assign n22648 = ~n22644 & ~n22647 ;
  assign n22649 = \s8_ack_i_pad  & n14690 ;
  assign n22650 = n13767 & n22649 ;
  assign n22651 = n13784 & n22650 ;
  assign n22652 = \s4_ack_i_pad  & n15030 ;
  assign n22653 = n13467 & n22652 ;
  assign n22654 = n13492 & n22653 ;
  assign n22655 = ~n22651 & ~n22654 ;
  assign n22656 = n22648 & n22655 ;
  assign n22657 = \s6_ack_i_pad  & n14681 ;
  assign n22658 = n13627 & n22657 ;
  assign n22659 = n13644 & n22658 ;
  assign n22660 = \s11_ack_i_pad  & n15003 ;
  assign n22661 = n14009 & n22660 ;
  assign n22662 = n14026 & n22661 ;
  assign n22663 = ~n22659 & ~n22662 ;
  assign n22664 = \s0_ack_i_pad  & n14634 ;
  assign n22665 = n14069 & n22664 ;
  assign n22666 = n14062 & n22665 ;
  assign n22667 = \s10_ack_i_pad  & n14999 ;
  assign n22668 = n13928 & n22667 ;
  assign n22669 = n13936 & n22668 ;
  assign n22670 = ~n22666 & ~n22669 ;
  assign n22671 = n22663 & n22670 ;
  assign n22672 = n22656 & n22671 ;
  assign n22673 = \s3_ack_i_pad  & n15026 ;
  assign n22674 = n14451 & n22673 ;
  assign n22675 = n14468 & n22674 ;
  assign n22676 = \s14_ack_i_pad  & n15015 ;
  assign n22677 = n14331 & n22676 ;
  assign n22678 = n14348 & n22677 ;
  assign n22679 = \s9_ack_i_pad  & n15042 ;
  assign n22680 = n13847 & n22679 ;
  assign n22681 = n13864 & n22680 ;
  assign n22682 = ~n22678 & ~n22681 ;
  assign n22683 = ~n22675 & n22682 ;
  assign n22684 = \s7_ack_i_pad  & n15038 ;
  assign n22685 = n13697 & n22684 ;
  assign n22686 = n13690 & n22685 ;
  assign n22687 = \s13_ack_i_pad  & n15011 ;
  assign n22688 = n14211 & n22687 ;
  assign n22689 = n14204 & n22688 ;
  assign n22690 = ~n22686 & ~n22689 ;
  assign n22691 = \s2_ack_i_pad  & n15022 ;
  assign n22692 = n14391 & n22691 ;
  assign n22693 = n14408 & n22692 ;
  assign n22694 = \s12_ack_i_pad  & n15007 ;
  assign n22695 = n14140 & n22694 ;
  assign n22696 = n14148 & n22695 ;
  assign n22697 = ~n22693 & ~n22696 ;
  assign n22698 = n22690 & n22697 ;
  assign n22699 = n22683 & n22698 ;
  assign n22700 = n22672 & n22699 ;
  assign n22701 = ~n22641 & n22700 ;
  assign n22702 = n2176 & n15192 ;
  assign n22703 = \s15_data_i[0]_pad  & n2176 ;
  assign n22704 = ~n2258 & n22703 ;
  assign n22705 = ~n22702 & ~n22704 ;
  assign n22706 = \s12_data_i[0]_pad  & n15007 ;
  assign n22707 = \s1_data_i[0]_pad  & n14640 ;
  assign n22708 = ~n22706 & ~n22707 ;
  assign n22709 = \s7_data_i[0]_pad  & n15038 ;
  assign n22710 = \s9_data_i[0]_pad  & n15042 ;
  assign n22711 = ~n22709 & ~n22710 ;
  assign n22712 = n22708 & n22711 ;
  assign n22713 = \s3_data_i[0]_pad  & n15026 ;
  assign n22714 = \s6_data_i[0]_pad  & n14681 ;
  assign n22715 = ~n22713 & ~n22714 ;
  assign n22716 = \s10_data_i[0]_pad  & n14999 ;
  assign n22717 = \s13_data_i[0]_pad  & n15011 ;
  assign n22718 = ~n22716 & ~n22717 ;
  assign n22719 = n22715 & n22718 ;
  assign n22720 = n22712 & n22719 ;
  assign n22721 = \s14_data_i[0]_pad  & n15015 ;
  assign n22722 = \s11_data_i[0]_pad  & n15003 ;
  assign n22723 = \s2_data_i[0]_pad  & n15022 ;
  assign n22724 = ~n22722 & ~n22723 ;
  assign n22725 = ~n22721 & n22724 ;
  assign n22726 = \s5_data_i[0]_pad  & n15034 ;
  assign n22727 = \s8_data_i[0]_pad  & n14690 ;
  assign n22728 = ~n22726 & ~n22727 ;
  assign n22729 = \s4_data_i[0]_pad  & n15030 ;
  assign n22730 = \s0_data_i[0]_pad  & n14634 ;
  assign n22731 = ~n22729 & ~n22730 ;
  assign n22732 = n22728 & n22731 ;
  assign n22733 = n22725 & n22732 ;
  assign n22734 = n22720 & n22733 ;
  assign n22735 = n22705 & n22734 ;
  assign n22736 = n2176 & n15229 ;
  assign n22737 = \s15_data_i[10]_pad  & n2176 ;
  assign n22738 = ~n2258 & n22737 ;
  assign n22739 = ~n22736 & ~n22738 ;
  assign n22740 = \s12_data_i[10]_pad  & n15007 ;
  assign n22741 = \s1_data_i[10]_pad  & n14640 ;
  assign n22742 = ~n22740 & ~n22741 ;
  assign n22743 = \s4_data_i[10]_pad  & n15030 ;
  assign n22744 = \s6_data_i[10]_pad  & n14681 ;
  assign n22745 = ~n22743 & ~n22744 ;
  assign n22746 = n22742 & n22745 ;
  assign n22747 = \s3_data_i[10]_pad  & n15026 ;
  assign n22748 = \s9_data_i[10]_pad  & n15042 ;
  assign n22749 = ~n22747 & ~n22748 ;
  assign n22750 = \s10_data_i[10]_pad  & n14999 ;
  assign n22751 = \s7_data_i[10]_pad  & n15038 ;
  assign n22752 = ~n22750 & ~n22751 ;
  assign n22753 = n22749 & n22752 ;
  assign n22754 = n22746 & n22753 ;
  assign n22755 = \s14_data_i[10]_pad  & n15015 ;
  assign n22756 = \s11_data_i[10]_pad  & n15003 ;
  assign n22757 = \s2_data_i[10]_pad  & n15022 ;
  assign n22758 = ~n22756 & ~n22757 ;
  assign n22759 = ~n22755 & n22758 ;
  assign n22760 = \s5_data_i[10]_pad  & n15034 ;
  assign n22761 = \s8_data_i[10]_pad  & n14690 ;
  assign n22762 = ~n22760 & ~n22761 ;
  assign n22763 = \s13_data_i[10]_pad  & n15011 ;
  assign n22764 = \s0_data_i[10]_pad  & n14634 ;
  assign n22765 = ~n22763 & ~n22764 ;
  assign n22766 = n22762 & n22765 ;
  assign n22767 = n22759 & n22766 ;
  assign n22768 = n22754 & n22767 ;
  assign n22769 = n22739 & n22768 ;
  assign n22770 = n2176 & n15266 ;
  assign n22771 = \s15_data_i[11]_pad  & n2176 ;
  assign n22772 = ~n2258 & n22771 ;
  assign n22773 = ~n22770 & ~n22772 ;
  assign n22774 = \s12_data_i[11]_pad  & n15007 ;
  assign n22775 = \s1_data_i[11]_pad  & n14640 ;
  assign n22776 = ~n22774 & ~n22775 ;
  assign n22777 = \s4_data_i[11]_pad  & n15030 ;
  assign n22778 = \s6_data_i[11]_pad  & n14681 ;
  assign n22779 = ~n22777 & ~n22778 ;
  assign n22780 = n22776 & n22779 ;
  assign n22781 = \s3_data_i[11]_pad  & n15026 ;
  assign n22782 = \s9_data_i[11]_pad  & n15042 ;
  assign n22783 = ~n22781 & ~n22782 ;
  assign n22784 = \s10_data_i[11]_pad  & n14999 ;
  assign n22785 = \s7_data_i[11]_pad  & n15038 ;
  assign n22786 = ~n22784 & ~n22785 ;
  assign n22787 = n22783 & n22786 ;
  assign n22788 = n22780 & n22787 ;
  assign n22789 = \s14_data_i[11]_pad  & n15015 ;
  assign n22790 = \s11_data_i[11]_pad  & n15003 ;
  assign n22791 = \s2_data_i[11]_pad  & n15022 ;
  assign n22792 = ~n22790 & ~n22791 ;
  assign n22793 = ~n22789 & n22792 ;
  assign n22794 = \s5_data_i[11]_pad  & n15034 ;
  assign n22795 = \s8_data_i[11]_pad  & n14690 ;
  assign n22796 = ~n22794 & ~n22795 ;
  assign n22797 = \s13_data_i[11]_pad  & n15011 ;
  assign n22798 = \s0_data_i[11]_pad  & n14634 ;
  assign n22799 = ~n22797 & ~n22798 ;
  assign n22800 = n22796 & n22799 ;
  assign n22801 = n22793 & n22800 ;
  assign n22802 = n22788 & n22801 ;
  assign n22803 = n22773 & n22802 ;
  assign n22804 = n2176 & n15303 ;
  assign n22805 = \s15_data_i[12]_pad  & n2176 ;
  assign n22806 = ~n2258 & n22805 ;
  assign n22807 = ~n22804 & ~n22806 ;
  assign n22808 = \s12_data_i[12]_pad  & n15007 ;
  assign n22809 = \s1_data_i[12]_pad  & n14640 ;
  assign n22810 = ~n22808 & ~n22809 ;
  assign n22811 = \s4_data_i[12]_pad  & n15030 ;
  assign n22812 = \s6_data_i[12]_pad  & n14681 ;
  assign n22813 = ~n22811 & ~n22812 ;
  assign n22814 = n22810 & n22813 ;
  assign n22815 = \s3_data_i[12]_pad  & n15026 ;
  assign n22816 = \s9_data_i[12]_pad  & n15042 ;
  assign n22817 = ~n22815 & ~n22816 ;
  assign n22818 = \s10_data_i[12]_pad  & n14999 ;
  assign n22819 = \s7_data_i[12]_pad  & n15038 ;
  assign n22820 = ~n22818 & ~n22819 ;
  assign n22821 = n22817 & n22820 ;
  assign n22822 = n22814 & n22821 ;
  assign n22823 = \s14_data_i[12]_pad  & n15015 ;
  assign n22824 = \s11_data_i[12]_pad  & n15003 ;
  assign n22825 = \s2_data_i[12]_pad  & n15022 ;
  assign n22826 = ~n22824 & ~n22825 ;
  assign n22827 = ~n22823 & n22826 ;
  assign n22828 = \s5_data_i[12]_pad  & n15034 ;
  assign n22829 = \s8_data_i[12]_pad  & n14690 ;
  assign n22830 = ~n22828 & ~n22829 ;
  assign n22831 = \s13_data_i[12]_pad  & n15011 ;
  assign n22832 = \s0_data_i[12]_pad  & n14634 ;
  assign n22833 = ~n22831 & ~n22832 ;
  assign n22834 = n22830 & n22833 ;
  assign n22835 = n22827 & n22834 ;
  assign n22836 = n22822 & n22835 ;
  assign n22837 = n22807 & n22836 ;
  assign n22838 = n2176 & n15340 ;
  assign n22839 = \s15_data_i[13]_pad  & n2176 ;
  assign n22840 = ~n2258 & n22839 ;
  assign n22841 = ~n22838 & ~n22840 ;
  assign n22842 = \s12_data_i[13]_pad  & n15007 ;
  assign n22843 = \s1_data_i[13]_pad  & n14640 ;
  assign n22844 = ~n22842 & ~n22843 ;
  assign n22845 = \s0_data_i[13]_pad  & n14634 ;
  assign n22846 = \s10_data_i[13]_pad  & n14999 ;
  assign n22847 = ~n22845 & ~n22846 ;
  assign n22848 = n22844 & n22847 ;
  assign n22849 = \s3_data_i[13]_pad  & n15026 ;
  assign n22850 = \s4_data_i[13]_pad  & n15030 ;
  assign n22851 = ~n22849 & ~n22850 ;
  assign n22852 = \s9_data_i[13]_pad  & n15042 ;
  assign n22853 = \s6_data_i[13]_pad  & n14681 ;
  assign n22854 = ~n22852 & ~n22853 ;
  assign n22855 = n22851 & n22854 ;
  assign n22856 = n22848 & n22855 ;
  assign n22857 = \s14_data_i[13]_pad  & n15015 ;
  assign n22858 = \s11_data_i[13]_pad  & n15003 ;
  assign n22859 = \s7_data_i[13]_pad  & n15038 ;
  assign n22860 = ~n22858 & ~n22859 ;
  assign n22861 = ~n22857 & n22860 ;
  assign n22862 = \s5_data_i[13]_pad  & n15034 ;
  assign n22863 = \s8_data_i[13]_pad  & n14690 ;
  assign n22864 = ~n22862 & ~n22863 ;
  assign n22865 = \s2_data_i[13]_pad  & n15022 ;
  assign n22866 = \s13_data_i[13]_pad  & n15011 ;
  assign n22867 = ~n22865 & ~n22866 ;
  assign n22868 = n22864 & n22867 ;
  assign n22869 = n22861 & n22868 ;
  assign n22870 = n22856 & n22869 ;
  assign n22871 = n22841 & n22870 ;
  assign n22872 = n2176 & n15377 ;
  assign n22873 = \s15_data_i[14]_pad  & n2176 ;
  assign n22874 = ~n2258 & n22873 ;
  assign n22875 = ~n22872 & ~n22874 ;
  assign n22876 = \s12_data_i[14]_pad  & n15007 ;
  assign n22877 = \s1_data_i[14]_pad  & n14640 ;
  assign n22878 = ~n22876 & ~n22877 ;
  assign n22879 = \s7_data_i[14]_pad  & n15038 ;
  assign n22880 = \s0_data_i[14]_pad  & n14634 ;
  assign n22881 = ~n22879 & ~n22880 ;
  assign n22882 = n22878 & n22881 ;
  assign n22883 = \s3_data_i[14]_pad  & n15026 ;
  assign n22884 = \s9_data_i[14]_pad  & n15042 ;
  assign n22885 = ~n22883 & ~n22884 ;
  assign n22886 = \s10_data_i[14]_pad  & n14999 ;
  assign n22887 = \s4_data_i[14]_pad  & n15030 ;
  assign n22888 = ~n22886 & ~n22887 ;
  assign n22889 = n22885 & n22888 ;
  assign n22890 = n22882 & n22889 ;
  assign n22891 = \s14_data_i[14]_pad  & n15015 ;
  assign n22892 = \s11_data_i[14]_pad  & n15003 ;
  assign n22893 = \s2_data_i[14]_pad  & n15022 ;
  assign n22894 = ~n22892 & ~n22893 ;
  assign n22895 = ~n22891 & n22894 ;
  assign n22896 = \s5_data_i[14]_pad  & n15034 ;
  assign n22897 = \s8_data_i[14]_pad  & n14690 ;
  assign n22898 = ~n22896 & ~n22897 ;
  assign n22899 = \s13_data_i[14]_pad  & n15011 ;
  assign n22900 = \s6_data_i[14]_pad  & n14681 ;
  assign n22901 = ~n22899 & ~n22900 ;
  assign n22902 = n22898 & n22901 ;
  assign n22903 = n22895 & n22902 ;
  assign n22904 = n22890 & n22903 ;
  assign n22905 = n22875 & n22904 ;
  assign n22906 = n2176 & n15414 ;
  assign n22907 = \s15_data_i[15]_pad  & n2176 ;
  assign n22908 = ~n2258 & n22907 ;
  assign n22909 = ~n22906 & ~n22908 ;
  assign n22910 = \s12_data_i[15]_pad  & n15007 ;
  assign n22911 = \s1_data_i[15]_pad  & n14640 ;
  assign n22912 = ~n22910 & ~n22911 ;
  assign n22913 = \s0_data_i[15]_pad  & n14634 ;
  assign n22914 = \s10_data_i[15]_pad  & n14999 ;
  assign n22915 = ~n22913 & ~n22914 ;
  assign n22916 = n22912 & n22915 ;
  assign n22917 = \s3_data_i[15]_pad  & n15026 ;
  assign n22918 = \s4_data_i[15]_pad  & n15030 ;
  assign n22919 = ~n22917 & ~n22918 ;
  assign n22920 = \s9_data_i[15]_pad  & n15042 ;
  assign n22921 = \s6_data_i[15]_pad  & n14681 ;
  assign n22922 = ~n22920 & ~n22921 ;
  assign n22923 = n22919 & n22922 ;
  assign n22924 = n22916 & n22923 ;
  assign n22925 = \s14_data_i[15]_pad  & n15015 ;
  assign n22926 = \s11_data_i[15]_pad  & n15003 ;
  assign n22927 = \s7_data_i[15]_pad  & n15038 ;
  assign n22928 = ~n22926 & ~n22927 ;
  assign n22929 = ~n22925 & n22928 ;
  assign n22930 = \s5_data_i[15]_pad  & n15034 ;
  assign n22931 = \s8_data_i[15]_pad  & n14690 ;
  assign n22932 = ~n22930 & ~n22931 ;
  assign n22933 = \s2_data_i[15]_pad  & n15022 ;
  assign n22934 = \s13_data_i[15]_pad  & n15011 ;
  assign n22935 = ~n22933 & ~n22934 ;
  assign n22936 = n22932 & n22935 ;
  assign n22937 = n22929 & n22936 ;
  assign n22938 = n22924 & n22937 ;
  assign n22939 = n22909 & n22938 ;
  assign n22940 = \s15_data_i[16]_pad  & n2176 ;
  assign n22941 = ~n2258 & n22940 ;
  assign n22942 = \s8_data_i[16]_pad  & n14690 ;
  assign n22943 = \s1_data_i[16]_pad  & n14640 ;
  assign n22944 = ~n22942 & ~n22943 ;
  assign n22945 = \s4_data_i[16]_pad  & n15030 ;
  assign n22946 = \s6_data_i[16]_pad  & n14681 ;
  assign n22947 = ~n22945 & ~n22946 ;
  assign n22948 = n22944 & n22947 ;
  assign n22949 = \s3_data_i[16]_pad  & n15026 ;
  assign n22950 = \s9_data_i[16]_pad  & n15042 ;
  assign n22951 = ~n22949 & ~n22950 ;
  assign n22952 = \s10_data_i[16]_pad  & n14999 ;
  assign n22953 = \s7_data_i[16]_pad  & n15038 ;
  assign n22954 = ~n22952 & ~n22953 ;
  assign n22955 = n22951 & n22954 ;
  assign n22956 = n22948 & n22955 ;
  assign n22957 = \s11_data_i[16]_pad  & n15003 ;
  assign n22958 = \s14_data_i[16]_pad  & n15015 ;
  assign n22959 = \s2_data_i[16]_pad  & n15022 ;
  assign n22960 = ~n22958 & ~n22959 ;
  assign n22961 = ~n22957 & n22960 ;
  assign n22962 = \s5_data_i[16]_pad  & n15034 ;
  assign n22963 = \s12_data_i[16]_pad  & n15007 ;
  assign n22964 = ~n22962 & ~n22963 ;
  assign n22965 = \s13_data_i[16]_pad  & n15011 ;
  assign n22966 = \s0_data_i[16]_pad  & n14634 ;
  assign n22967 = ~n22965 & ~n22966 ;
  assign n22968 = n22964 & n22967 ;
  assign n22969 = n22961 & n22968 ;
  assign n22970 = n22956 & n22969 ;
  assign n22971 = ~n22941 & n22970 ;
  assign n22972 = \s15_data_i[17]_pad  & n2176 ;
  assign n22973 = ~n2258 & n22972 ;
  assign n22974 = \s8_data_i[17]_pad  & n14690 ;
  assign n22975 = \s1_data_i[17]_pad  & n14640 ;
  assign n22976 = ~n22974 & ~n22975 ;
  assign n22977 = \s4_data_i[17]_pad  & n15030 ;
  assign n22978 = \s6_data_i[17]_pad  & n14681 ;
  assign n22979 = ~n22977 & ~n22978 ;
  assign n22980 = n22976 & n22979 ;
  assign n22981 = \s3_data_i[17]_pad  & n15026 ;
  assign n22982 = \s9_data_i[17]_pad  & n15042 ;
  assign n22983 = ~n22981 & ~n22982 ;
  assign n22984 = \s10_data_i[17]_pad  & n14999 ;
  assign n22985 = \s7_data_i[17]_pad  & n15038 ;
  assign n22986 = ~n22984 & ~n22985 ;
  assign n22987 = n22983 & n22986 ;
  assign n22988 = n22980 & n22987 ;
  assign n22989 = \s11_data_i[17]_pad  & n15003 ;
  assign n22990 = \s14_data_i[17]_pad  & n15015 ;
  assign n22991 = \s2_data_i[17]_pad  & n15022 ;
  assign n22992 = ~n22990 & ~n22991 ;
  assign n22993 = ~n22989 & n22992 ;
  assign n22994 = \s5_data_i[17]_pad  & n15034 ;
  assign n22995 = \s12_data_i[17]_pad  & n15007 ;
  assign n22996 = ~n22994 & ~n22995 ;
  assign n22997 = \s13_data_i[17]_pad  & n15011 ;
  assign n22998 = \s0_data_i[17]_pad  & n14634 ;
  assign n22999 = ~n22997 & ~n22998 ;
  assign n23000 = n22996 & n22999 ;
  assign n23001 = n22993 & n23000 ;
  assign n23002 = n22988 & n23001 ;
  assign n23003 = ~n22973 & n23002 ;
  assign n23004 = \s15_data_i[18]_pad  & n2176 ;
  assign n23005 = ~n2258 & n23004 ;
  assign n23006 = \s8_data_i[18]_pad  & n14690 ;
  assign n23007 = \s1_data_i[18]_pad  & n14640 ;
  assign n23008 = ~n23006 & ~n23007 ;
  assign n23009 = \s4_data_i[18]_pad  & n15030 ;
  assign n23010 = \s6_data_i[18]_pad  & n14681 ;
  assign n23011 = ~n23009 & ~n23010 ;
  assign n23012 = n23008 & n23011 ;
  assign n23013 = \s3_data_i[18]_pad  & n15026 ;
  assign n23014 = \s9_data_i[18]_pad  & n15042 ;
  assign n23015 = ~n23013 & ~n23014 ;
  assign n23016 = \s10_data_i[18]_pad  & n14999 ;
  assign n23017 = \s7_data_i[18]_pad  & n15038 ;
  assign n23018 = ~n23016 & ~n23017 ;
  assign n23019 = n23015 & n23018 ;
  assign n23020 = n23012 & n23019 ;
  assign n23021 = \s11_data_i[18]_pad  & n15003 ;
  assign n23022 = \s14_data_i[18]_pad  & n15015 ;
  assign n23023 = \s2_data_i[18]_pad  & n15022 ;
  assign n23024 = ~n23022 & ~n23023 ;
  assign n23025 = ~n23021 & n23024 ;
  assign n23026 = \s5_data_i[18]_pad  & n15034 ;
  assign n23027 = \s12_data_i[18]_pad  & n15007 ;
  assign n23028 = ~n23026 & ~n23027 ;
  assign n23029 = \s13_data_i[18]_pad  & n15011 ;
  assign n23030 = \s0_data_i[18]_pad  & n14634 ;
  assign n23031 = ~n23029 & ~n23030 ;
  assign n23032 = n23028 & n23031 ;
  assign n23033 = n23025 & n23032 ;
  assign n23034 = n23020 & n23033 ;
  assign n23035 = ~n23005 & n23034 ;
  assign n23036 = \s15_data_i[19]_pad  & n2176 ;
  assign n23037 = ~n2258 & n23036 ;
  assign n23038 = \s8_data_i[19]_pad  & n14690 ;
  assign n23039 = \s1_data_i[19]_pad  & n14640 ;
  assign n23040 = ~n23038 & ~n23039 ;
  assign n23041 = \s4_data_i[19]_pad  & n15030 ;
  assign n23042 = \s6_data_i[19]_pad  & n14681 ;
  assign n23043 = ~n23041 & ~n23042 ;
  assign n23044 = n23040 & n23043 ;
  assign n23045 = \s3_data_i[19]_pad  & n15026 ;
  assign n23046 = \s9_data_i[19]_pad  & n15042 ;
  assign n23047 = ~n23045 & ~n23046 ;
  assign n23048 = \s10_data_i[19]_pad  & n14999 ;
  assign n23049 = \s7_data_i[19]_pad  & n15038 ;
  assign n23050 = ~n23048 & ~n23049 ;
  assign n23051 = n23047 & n23050 ;
  assign n23052 = n23044 & n23051 ;
  assign n23053 = \s11_data_i[19]_pad  & n15003 ;
  assign n23054 = \s14_data_i[19]_pad  & n15015 ;
  assign n23055 = \s2_data_i[19]_pad  & n15022 ;
  assign n23056 = ~n23054 & ~n23055 ;
  assign n23057 = ~n23053 & n23056 ;
  assign n23058 = \s5_data_i[19]_pad  & n15034 ;
  assign n23059 = \s12_data_i[19]_pad  & n15007 ;
  assign n23060 = ~n23058 & ~n23059 ;
  assign n23061 = \s13_data_i[19]_pad  & n15011 ;
  assign n23062 = \s0_data_i[19]_pad  & n14634 ;
  assign n23063 = ~n23061 & ~n23062 ;
  assign n23064 = n23060 & n23063 ;
  assign n23065 = n23057 & n23064 ;
  assign n23066 = n23052 & n23065 ;
  assign n23067 = ~n23037 & n23066 ;
  assign n23068 = n2176 & n15579 ;
  assign n23069 = \s15_data_i[1]_pad  & n2176 ;
  assign n23070 = ~n2258 & n23069 ;
  assign n23071 = ~n23068 & ~n23070 ;
  assign n23072 = \s12_data_i[1]_pad  & n15007 ;
  assign n23073 = \s1_data_i[1]_pad  & n14640 ;
  assign n23074 = ~n23072 & ~n23073 ;
  assign n23075 = \s0_data_i[1]_pad  & n14634 ;
  assign n23076 = \s10_data_i[1]_pad  & n14999 ;
  assign n23077 = ~n23075 & ~n23076 ;
  assign n23078 = n23074 & n23077 ;
  assign n23079 = \s3_data_i[1]_pad  & n15026 ;
  assign n23080 = \s4_data_i[1]_pad  & n15030 ;
  assign n23081 = ~n23079 & ~n23080 ;
  assign n23082 = \s9_data_i[1]_pad  & n15042 ;
  assign n23083 = \s6_data_i[1]_pad  & n14681 ;
  assign n23084 = ~n23082 & ~n23083 ;
  assign n23085 = n23081 & n23084 ;
  assign n23086 = n23078 & n23085 ;
  assign n23087 = \s14_data_i[1]_pad  & n15015 ;
  assign n23088 = \s11_data_i[1]_pad  & n15003 ;
  assign n23089 = \s7_data_i[1]_pad  & n15038 ;
  assign n23090 = ~n23088 & ~n23089 ;
  assign n23091 = ~n23087 & n23090 ;
  assign n23092 = \s5_data_i[1]_pad  & n15034 ;
  assign n23093 = \s8_data_i[1]_pad  & n14690 ;
  assign n23094 = ~n23092 & ~n23093 ;
  assign n23095 = \s2_data_i[1]_pad  & n15022 ;
  assign n23096 = \s13_data_i[1]_pad  & n15011 ;
  assign n23097 = ~n23095 & ~n23096 ;
  assign n23098 = n23094 & n23097 ;
  assign n23099 = n23091 & n23098 ;
  assign n23100 = n23086 & n23099 ;
  assign n23101 = n23071 & n23100 ;
  assign n23102 = \s15_data_i[20]_pad  & n2176 ;
  assign n23103 = ~n2258 & n23102 ;
  assign n23104 = \s8_data_i[20]_pad  & n14690 ;
  assign n23105 = \s1_data_i[20]_pad  & n14640 ;
  assign n23106 = ~n23104 & ~n23105 ;
  assign n23107 = \s4_data_i[20]_pad  & n15030 ;
  assign n23108 = \s6_data_i[20]_pad  & n14681 ;
  assign n23109 = ~n23107 & ~n23108 ;
  assign n23110 = n23106 & n23109 ;
  assign n23111 = \s3_data_i[20]_pad  & n15026 ;
  assign n23112 = \s9_data_i[20]_pad  & n15042 ;
  assign n23113 = ~n23111 & ~n23112 ;
  assign n23114 = \s10_data_i[20]_pad  & n14999 ;
  assign n23115 = \s7_data_i[20]_pad  & n15038 ;
  assign n23116 = ~n23114 & ~n23115 ;
  assign n23117 = n23113 & n23116 ;
  assign n23118 = n23110 & n23117 ;
  assign n23119 = \s11_data_i[20]_pad  & n15003 ;
  assign n23120 = \s14_data_i[20]_pad  & n15015 ;
  assign n23121 = \s2_data_i[20]_pad  & n15022 ;
  assign n23122 = ~n23120 & ~n23121 ;
  assign n23123 = ~n23119 & n23122 ;
  assign n23124 = \s5_data_i[20]_pad  & n15034 ;
  assign n23125 = \s12_data_i[20]_pad  & n15007 ;
  assign n23126 = ~n23124 & ~n23125 ;
  assign n23127 = \s13_data_i[20]_pad  & n15011 ;
  assign n23128 = \s0_data_i[20]_pad  & n14634 ;
  assign n23129 = ~n23127 & ~n23128 ;
  assign n23130 = n23126 & n23129 ;
  assign n23131 = n23123 & n23130 ;
  assign n23132 = n23118 & n23131 ;
  assign n23133 = ~n23103 & n23132 ;
  assign n23134 = \s15_data_i[21]_pad  & n2176 ;
  assign n23135 = ~n2258 & n23134 ;
  assign n23136 = \s8_data_i[21]_pad  & n14690 ;
  assign n23137 = \s1_data_i[21]_pad  & n14640 ;
  assign n23138 = ~n23136 & ~n23137 ;
  assign n23139 = \s4_data_i[21]_pad  & n15030 ;
  assign n23140 = \s6_data_i[21]_pad  & n14681 ;
  assign n23141 = ~n23139 & ~n23140 ;
  assign n23142 = n23138 & n23141 ;
  assign n23143 = \s3_data_i[21]_pad  & n15026 ;
  assign n23144 = \s9_data_i[21]_pad  & n15042 ;
  assign n23145 = ~n23143 & ~n23144 ;
  assign n23146 = \s10_data_i[21]_pad  & n14999 ;
  assign n23147 = \s7_data_i[21]_pad  & n15038 ;
  assign n23148 = ~n23146 & ~n23147 ;
  assign n23149 = n23145 & n23148 ;
  assign n23150 = n23142 & n23149 ;
  assign n23151 = \s11_data_i[21]_pad  & n15003 ;
  assign n23152 = \s14_data_i[21]_pad  & n15015 ;
  assign n23153 = \s2_data_i[21]_pad  & n15022 ;
  assign n23154 = ~n23152 & ~n23153 ;
  assign n23155 = ~n23151 & n23154 ;
  assign n23156 = \s5_data_i[21]_pad  & n15034 ;
  assign n23157 = \s12_data_i[21]_pad  & n15007 ;
  assign n23158 = ~n23156 & ~n23157 ;
  assign n23159 = \s13_data_i[21]_pad  & n15011 ;
  assign n23160 = \s0_data_i[21]_pad  & n14634 ;
  assign n23161 = ~n23159 & ~n23160 ;
  assign n23162 = n23158 & n23161 ;
  assign n23163 = n23155 & n23162 ;
  assign n23164 = n23150 & n23163 ;
  assign n23165 = ~n23135 & n23164 ;
  assign n23166 = \s15_data_i[22]_pad  & n2176 ;
  assign n23167 = ~n2258 & n23166 ;
  assign n23168 = \s8_data_i[22]_pad  & n14690 ;
  assign n23169 = \s1_data_i[22]_pad  & n14640 ;
  assign n23170 = ~n23168 & ~n23169 ;
  assign n23171 = \s7_data_i[22]_pad  & n15038 ;
  assign n23172 = \s0_data_i[22]_pad  & n14634 ;
  assign n23173 = ~n23171 & ~n23172 ;
  assign n23174 = n23170 & n23173 ;
  assign n23175 = \s3_data_i[22]_pad  & n15026 ;
  assign n23176 = \s9_data_i[22]_pad  & n15042 ;
  assign n23177 = ~n23175 & ~n23176 ;
  assign n23178 = \s10_data_i[22]_pad  & n14999 ;
  assign n23179 = \s4_data_i[22]_pad  & n15030 ;
  assign n23180 = ~n23178 & ~n23179 ;
  assign n23181 = n23177 & n23180 ;
  assign n23182 = n23174 & n23181 ;
  assign n23183 = \s11_data_i[22]_pad  & n15003 ;
  assign n23184 = \s14_data_i[22]_pad  & n15015 ;
  assign n23185 = \s2_data_i[22]_pad  & n15022 ;
  assign n23186 = ~n23184 & ~n23185 ;
  assign n23187 = ~n23183 & n23186 ;
  assign n23188 = \s5_data_i[22]_pad  & n15034 ;
  assign n23189 = \s12_data_i[22]_pad  & n15007 ;
  assign n23190 = ~n23188 & ~n23189 ;
  assign n23191 = \s13_data_i[22]_pad  & n15011 ;
  assign n23192 = \s6_data_i[22]_pad  & n14681 ;
  assign n23193 = ~n23191 & ~n23192 ;
  assign n23194 = n23190 & n23193 ;
  assign n23195 = n23187 & n23194 ;
  assign n23196 = n23182 & n23195 ;
  assign n23197 = ~n23167 & n23196 ;
  assign n23198 = \s15_data_i[23]_pad  & n2176 ;
  assign n23199 = ~n2258 & n23198 ;
  assign n23200 = \s8_data_i[23]_pad  & n14690 ;
  assign n23201 = \s1_data_i[23]_pad  & n14640 ;
  assign n23202 = ~n23200 & ~n23201 ;
  assign n23203 = \s4_data_i[23]_pad  & n15030 ;
  assign n23204 = \s6_data_i[23]_pad  & n14681 ;
  assign n23205 = ~n23203 & ~n23204 ;
  assign n23206 = n23202 & n23205 ;
  assign n23207 = \s5_data_i[23]_pad  & n15034 ;
  assign n23208 = \s9_data_i[23]_pad  & n15042 ;
  assign n23209 = ~n23207 & ~n23208 ;
  assign n23210 = \s10_data_i[23]_pad  & n14999 ;
  assign n23211 = \s7_data_i[23]_pad  & n15038 ;
  assign n23212 = ~n23210 & ~n23211 ;
  assign n23213 = n23209 & n23212 ;
  assign n23214 = n23206 & n23213 ;
  assign n23215 = \s11_data_i[23]_pad  & n15003 ;
  assign n23216 = \s14_data_i[23]_pad  & n15015 ;
  assign n23217 = \s3_data_i[23]_pad  & n15026 ;
  assign n23218 = ~n23216 & ~n23217 ;
  assign n23219 = ~n23215 & n23218 ;
  assign n23220 = \s2_data_i[23]_pad  & n15022 ;
  assign n23221 = \s12_data_i[23]_pad  & n15007 ;
  assign n23222 = ~n23220 & ~n23221 ;
  assign n23223 = \s13_data_i[23]_pad  & n15011 ;
  assign n23224 = \s0_data_i[23]_pad  & n14634 ;
  assign n23225 = ~n23223 & ~n23224 ;
  assign n23226 = n23222 & n23225 ;
  assign n23227 = n23219 & n23226 ;
  assign n23228 = n23214 & n23227 ;
  assign n23229 = ~n23199 & n23228 ;
  assign n23230 = \s15_data_i[24]_pad  & n2176 ;
  assign n23231 = ~n2258 & n23230 ;
  assign n23232 = \s8_data_i[24]_pad  & n14690 ;
  assign n23233 = \s1_data_i[24]_pad  & n14640 ;
  assign n23234 = ~n23232 & ~n23233 ;
  assign n23235 = \s4_data_i[24]_pad  & n15030 ;
  assign n23236 = \s6_data_i[24]_pad  & n14681 ;
  assign n23237 = ~n23235 & ~n23236 ;
  assign n23238 = n23234 & n23237 ;
  assign n23239 = \s3_data_i[24]_pad  & n15026 ;
  assign n23240 = \s9_data_i[24]_pad  & n15042 ;
  assign n23241 = ~n23239 & ~n23240 ;
  assign n23242 = \s10_data_i[24]_pad  & n14999 ;
  assign n23243 = \s7_data_i[24]_pad  & n15038 ;
  assign n23244 = ~n23242 & ~n23243 ;
  assign n23245 = n23241 & n23244 ;
  assign n23246 = n23238 & n23245 ;
  assign n23247 = \s11_data_i[24]_pad  & n15003 ;
  assign n23248 = \s14_data_i[24]_pad  & n15015 ;
  assign n23249 = \s2_data_i[24]_pad  & n15022 ;
  assign n23250 = ~n23248 & ~n23249 ;
  assign n23251 = ~n23247 & n23250 ;
  assign n23252 = \s5_data_i[24]_pad  & n15034 ;
  assign n23253 = \s12_data_i[24]_pad  & n15007 ;
  assign n23254 = ~n23252 & ~n23253 ;
  assign n23255 = \s13_data_i[24]_pad  & n15011 ;
  assign n23256 = \s0_data_i[24]_pad  & n14634 ;
  assign n23257 = ~n23255 & ~n23256 ;
  assign n23258 = n23254 & n23257 ;
  assign n23259 = n23251 & n23258 ;
  assign n23260 = n23246 & n23259 ;
  assign n23261 = ~n23231 & n23260 ;
  assign n23262 = \s15_data_i[25]_pad  & n2176 ;
  assign n23263 = ~n2258 & n23262 ;
  assign n23264 = \s8_data_i[25]_pad  & n14690 ;
  assign n23265 = \s1_data_i[25]_pad  & n14640 ;
  assign n23266 = ~n23264 & ~n23265 ;
  assign n23267 = \s4_data_i[25]_pad  & n15030 ;
  assign n23268 = \s6_data_i[25]_pad  & n14681 ;
  assign n23269 = ~n23267 & ~n23268 ;
  assign n23270 = n23266 & n23269 ;
  assign n23271 = \s3_data_i[25]_pad  & n15026 ;
  assign n23272 = \s9_data_i[25]_pad  & n15042 ;
  assign n23273 = ~n23271 & ~n23272 ;
  assign n23274 = \s10_data_i[25]_pad  & n14999 ;
  assign n23275 = \s7_data_i[25]_pad  & n15038 ;
  assign n23276 = ~n23274 & ~n23275 ;
  assign n23277 = n23273 & n23276 ;
  assign n23278 = n23270 & n23277 ;
  assign n23279 = \s11_data_i[25]_pad  & n15003 ;
  assign n23280 = \s14_data_i[25]_pad  & n15015 ;
  assign n23281 = \s2_data_i[25]_pad  & n15022 ;
  assign n23282 = ~n23280 & ~n23281 ;
  assign n23283 = ~n23279 & n23282 ;
  assign n23284 = \s5_data_i[25]_pad  & n15034 ;
  assign n23285 = \s12_data_i[25]_pad  & n15007 ;
  assign n23286 = ~n23284 & ~n23285 ;
  assign n23287 = \s13_data_i[25]_pad  & n15011 ;
  assign n23288 = \s0_data_i[25]_pad  & n14634 ;
  assign n23289 = ~n23287 & ~n23288 ;
  assign n23290 = n23286 & n23289 ;
  assign n23291 = n23283 & n23290 ;
  assign n23292 = n23278 & n23291 ;
  assign n23293 = ~n23263 & n23292 ;
  assign n23294 = \s15_data_i[26]_pad  & n2176 ;
  assign n23295 = ~n2258 & n23294 ;
  assign n23296 = \s8_data_i[26]_pad  & n14690 ;
  assign n23297 = \s1_data_i[26]_pad  & n14640 ;
  assign n23298 = ~n23296 & ~n23297 ;
  assign n23299 = \s4_data_i[26]_pad  & n15030 ;
  assign n23300 = \s6_data_i[26]_pad  & n14681 ;
  assign n23301 = ~n23299 & ~n23300 ;
  assign n23302 = n23298 & n23301 ;
  assign n23303 = \s3_data_i[26]_pad  & n15026 ;
  assign n23304 = \s9_data_i[26]_pad  & n15042 ;
  assign n23305 = ~n23303 & ~n23304 ;
  assign n23306 = \s10_data_i[26]_pad  & n14999 ;
  assign n23307 = \s7_data_i[26]_pad  & n15038 ;
  assign n23308 = ~n23306 & ~n23307 ;
  assign n23309 = n23305 & n23308 ;
  assign n23310 = n23302 & n23309 ;
  assign n23311 = \s11_data_i[26]_pad  & n15003 ;
  assign n23312 = \s14_data_i[26]_pad  & n15015 ;
  assign n23313 = \s2_data_i[26]_pad  & n15022 ;
  assign n23314 = ~n23312 & ~n23313 ;
  assign n23315 = ~n23311 & n23314 ;
  assign n23316 = \s5_data_i[26]_pad  & n15034 ;
  assign n23317 = \s12_data_i[26]_pad  & n15007 ;
  assign n23318 = ~n23316 & ~n23317 ;
  assign n23319 = \s13_data_i[26]_pad  & n15011 ;
  assign n23320 = \s0_data_i[26]_pad  & n14634 ;
  assign n23321 = ~n23319 & ~n23320 ;
  assign n23322 = n23318 & n23321 ;
  assign n23323 = n23315 & n23322 ;
  assign n23324 = n23310 & n23323 ;
  assign n23325 = ~n23295 & n23324 ;
  assign n23326 = \s15_data_i[27]_pad  & n2176 ;
  assign n23327 = ~n2258 & n23326 ;
  assign n23328 = \s8_data_i[27]_pad  & n14690 ;
  assign n23329 = \s1_data_i[27]_pad  & n14640 ;
  assign n23330 = ~n23328 & ~n23329 ;
  assign n23331 = \s4_data_i[27]_pad  & n15030 ;
  assign n23332 = \s6_data_i[27]_pad  & n14681 ;
  assign n23333 = ~n23331 & ~n23332 ;
  assign n23334 = n23330 & n23333 ;
  assign n23335 = \s3_data_i[27]_pad  & n15026 ;
  assign n23336 = \s9_data_i[27]_pad  & n15042 ;
  assign n23337 = ~n23335 & ~n23336 ;
  assign n23338 = \s10_data_i[27]_pad  & n14999 ;
  assign n23339 = \s7_data_i[27]_pad  & n15038 ;
  assign n23340 = ~n23338 & ~n23339 ;
  assign n23341 = n23337 & n23340 ;
  assign n23342 = n23334 & n23341 ;
  assign n23343 = \s11_data_i[27]_pad  & n15003 ;
  assign n23344 = \s14_data_i[27]_pad  & n15015 ;
  assign n23345 = \s2_data_i[27]_pad  & n15022 ;
  assign n23346 = ~n23344 & ~n23345 ;
  assign n23347 = ~n23343 & n23346 ;
  assign n23348 = \s5_data_i[27]_pad  & n15034 ;
  assign n23349 = \s12_data_i[27]_pad  & n15007 ;
  assign n23350 = ~n23348 & ~n23349 ;
  assign n23351 = \s13_data_i[27]_pad  & n15011 ;
  assign n23352 = \s0_data_i[27]_pad  & n14634 ;
  assign n23353 = ~n23351 & ~n23352 ;
  assign n23354 = n23350 & n23353 ;
  assign n23355 = n23347 & n23354 ;
  assign n23356 = n23342 & n23355 ;
  assign n23357 = ~n23327 & n23356 ;
  assign n23358 = \s15_data_i[28]_pad  & n2176 ;
  assign n23359 = ~n2258 & n23358 ;
  assign n23360 = \s8_data_i[28]_pad  & n14690 ;
  assign n23361 = \s1_data_i[28]_pad  & n14640 ;
  assign n23362 = ~n23360 & ~n23361 ;
  assign n23363 = \s4_data_i[28]_pad  & n15030 ;
  assign n23364 = \s6_data_i[28]_pad  & n14681 ;
  assign n23365 = ~n23363 & ~n23364 ;
  assign n23366 = n23362 & n23365 ;
  assign n23367 = \s3_data_i[28]_pad  & n15026 ;
  assign n23368 = \s9_data_i[28]_pad  & n15042 ;
  assign n23369 = ~n23367 & ~n23368 ;
  assign n23370 = \s10_data_i[28]_pad  & n14999 ;
  assign n23371 = \s7_data_i[28]_pad  & n15038 ;
  assign n23372 = ~n23370 & ~n23371 ;
  assign n23373 = n23369 & n23372 ;
  assign n23374 = n23366 & n23373 ;
  assign n23375 = \s11_data_i[28]_pad  & n15003 ;
  assign n23376 = \s14_data_i[28]_pad  & n15015 ;
  assign n23377 = \s2_data_i[28]_pad  & n15022 ;
  assign n23378 = ~n23376 & ~n23377 ;
  assign n23379 = ~n23375 & n23378 ;
  assign n23380 = \s5_data_i[28]_pad  & n15034 ;
  assign n23381 = \s12_data_i[28]_pad  & n15007 ;
  assign n23382 = ~n23380 & ~n23381 ;
  assign n23383 = \s13_data_i[28]_pad  & n15011 ;
  assign n23384 = \s0_data_i[28]_pad  & n14634 ;
  assign n23385 = ~n23383 & ~n23384 ;
  assign n23386 = n23382 & n23385 ;
  assign n23387 = n23379 & n23386 ;
  assign n23388 = n23374 & n23387 ;
  assign n23389 = ~n23359 & n23388 ;
  assign n23390 = \s15_data_i[29]_pad  & n2176 ;
  assign n23391 = ~n2258 & n23390 ;
  assign n23392 = \s8_data_i[29]_pad  & n14690 ;
  assign n23393 = \s1_data_i[29]_pad  & n14640 ;
  assign n23394 = ~n23392 & ~n23393 ;
  assign n23395 = \s4_data_i[29]_pad  & n15030 ;
  assign n23396 = \s6_data_i[29]_pad  & n14681 ;
  assign n23397 = ~n23395 & ~n23396 ;
  assign n23398 = n23394 & n23397 ;
  assign n23399 = \s3_data_i[29]_pad  & n15026 ;
  assign n23400 = \s9_data_i[29]_pad  & n15042 ;
  assign n23401 = ~n23399 & ~n23400 ;
  assign n23402 = \s10_data_i[29]_pad  & n14999 ;
  assign n23403 = \s7_data_i[29]_pad  & n15038 ;
  assign n23404 = ~n23402 & ~n23403 ;
  assign n23405 = n23401 & n23404 ;
  assign n23406 = n23398 & n23405 ;
  assign n23407 = \s11_data_i[29]_pad  & n15003 ;
  assign n23408 = \s14_data_i[29]_pad  & n15015 ;
  assign n23409 = \s2_data_i[29]_pad  & n15022 ;
  assign n23410 = ~n23408 & ~n23409 ;
  assign n23411 = ~n23407 & n23410 ;
  assign n23412 = \s5_data_i[29]_pad  & n15034 ;
  assign n23413 = \s12_data_i[29]_pad  & n15007 ;
  assign n23414 = ~n23412 & ~n23413 ;
  assign n23415 = \s13_data_i[29]_pad  & n15011 ;
  assign n23416 = \s0_data_i[29]_pad  & n14634 ;
  assign n23417 = ~n23415 & ~n23416 ;
  assign n23418 = n23414 & n23417 ;
  assign n23419 = n23411 & n23418 ;
  assign n23420 = n23406 & n23419 ;
  assign n23421 = ~n23391 & n23420 ;
  assign n23422 = n2176 & n15936 ;
  assign n23423 = \s15_data_i[2]_pad  & n2176 ;
  assign n23424 = ~n2258 & n23423 ;
  assign n23425 = ~n23422 & ~n23424 ;
  assign n23426 = \s12_data_i[2]_pad  & n15007 ;
  assign n23427 = \s1_data_i[2]_pad  & n14640 ;
  assign n23428 = ~n23426 & ~n23427 ;
  assign n23429 = \s0_data_i[2]_pad  & n14634 ;
  assign n23430 = \s10_data_i[2]_pad  & n14999 ;
  assign n23431 = ~n23429 & ~n23430 ;
  assign n23432 = n23428 & n23431 ;
  assign n23433 = \s3_data_i[2]_pad  & n15026 ;
  assign n23434 = \s4_data_i[2]_pad  & n15030 ;
  assign n23435 = ~n23433 & ~n23434 ;
  assign n23436 = \s9_data_i[2]_pad  & n15042 ;
  assign n23437 = \s6_data_i[2]_pad  & n14681 ;
  assign n23438 = ~n23436 & ~n23437 ;
  assign n23439 = n23435 & n23438 ;
  assign n23440 = n23432 & n23439 ;
  assign n23441 = \s14_data_i[2]_pad  & n15015 ;
  assign n23442 = \s11_data_i[2]_pad  & n15003 ;
  assign n23443 = \s7_data_i[2]_pad  & n15038 ;
  assign n23444 = ~n23442 & ~n23443 ;
  assign n23445 = ~n23441 & n23444 ;
  assign n23446 = \s5_data_i[2]_pad  & n15034 ;
  assign n23447 = \s8_data_i[2]_pad  & n14690 ;
  assign n23448 = ~n23446 & ~n23447 ;
  assign n23449 = \s2_data_i[2]_pad  & n15022 ;
  assign n23450 = \s13_data_i[2]_pad  & n15011 ;
  assign n23451 = ~n23449 & ~n23450 ;
  assign n23452 = n23448 & n23451 ;
  assign n23453 = n23445 & n23452 ;
  assign n23454 = n23440 & n23453 ;
  assign n23455 = n23425 & n23454 ;
  assign n23456 = \s15_data_i[30]_pad  & n2176 ;
  assign n23457 = ~n2258 & n23456 ;
  assign n23458 = \s8_data_i[30]_pad  & n14690 ;
  assign n23459 = \s1_data_i[30]_pad  & n14640 ;
  assign n23460 = ~n23458 & ~n23459 ;
  assign n23461 = \s4_data_i[30]_pad  & n15030 ;
  assign n23462 = \s6_data_i[30]_pad  & n14681 ;
  assign n23463 = ~n23461 & ~n23462 ;
  assign n23464 = n23460 & n23463 ;
  assign n23465 = \s3_data_i[30]_pad  & n15026 ;
  assign n23466 = \s9_data_i[30]_pad  & n15042 ;
  assign n23467 = ~n23465 & ~n23466 ;
  assign n23468 = \s10_data_i[30]_pad  & n14999 ;
  assign n23469 = \s7_data_i[30]_pad  & n15038 ;
  assign n23470 = ~n23468 & ~n23469 ;
  assign n23471 = n23467 & n23470 ;
  assign n23472 = n23464 & n23471 ;
  assign n23473 = \s11_data_i[30]_pad  & n15003 ;
  assign n23474 = \s14_data_i[30]_pad  & n15015 ;
  assign n23475 = \s2_data_i[30]_pad  & n15022 ;
  assign n23476 = ~n23474 & ~n23475 ;
  assign n23477 = ~n23473 & n23476 ;
  assign n23478 = \s5_data_i[30]_pad  & n15034 ;
  assign n23479 = \s12_data_i[30]_pad  & n15007 ;
  assign n23480 = ~n23478 & ~n23479 ;
  assign n23481 = \s13_data_i[30]_pad  & n15011 ;
  assign n23482 = \s0_data_i[30]_pad  & n14634 ;
  assign n23483 = ~n23481 & ~n23482 ;
  assign n23484 = n23480 & n23483 ;
  assign n23485 = n23477 & n23484 ;
  assign n23486 = n23472 & n23485 ;
  assign n23487 = ~n23457 & n23486 ;
  assign n23488 = \s15_data_i[31]_pad  & n2176 ;
  assign n23489 = ~n2258 & n23488 ;
  assign n23490 = \s8_data_i[31]_pad  & n14690 ;
  assign n23491 = \s1_data_i[31]_pad  & n14640 ;
  assign n23492 = ~n23490 & ~n23491 ;
  assign n23493 = \s4_data_i[31]_pad  & n15030 ;
  assign n23494 = \s6_data_i[31]_pad  & n14681 ;
  assign n23495 = ~n23493 & ~n23494 ;
  assign n23496 = n23492 & n23495 ;
  assign n23497 = \s3_data_i[31]_pad  & n15026 ;
  assign n23498 = \s9_data_i[31]_pad  & n15042 ;
  assign n23499 = ~n23497 & ~n23498 ;
  assign n23500 = \s10_data_i[31]_pad  & n14999 ;
  assign n23501 = \s7_data_i[31]_pad  & n15038 ;
  assign n23502 = ~n23500 & ~n23501 ;
  assign n23503 = n23499 & n23502 ;
  assign n23504 = n23496 & n23503 ;
  assign n23505 = \s11_data_i[31]_pad  & n15003 ;
  assign n23506 = \s14_data_i[31]_pad  & n15015 ;
  assign n23507 = \s2_data_i[31]_pad  & n15022 ;
  assign n23508 = ~n23506 & ~n23507 ;
  assign n23509 = ~n23505 & n23508 ;
  assign n23510 = \s5_data_i[31]_pad  & n15034 ;
  assign n23511 = \s12_data_i[31]_pad  & n15007 ;
  assign n23512 = ~n23510 & ~n23511 ;
  assign n23513 = \s13_data_i[31]_pad  & n15011 ;
  assign n23514 = \s0_data_i[31]_pad  & n14634 ;
  assign n23515 = ~n23513 & ~n23514 ;
  assign n23516 = n23512 & n23515 ;
  assign n23517 = n23509 & n23516 ;
  assign n23518 = n23504 & n23517 ;
  assign n23519 = ~n23489 & n23518 ;
  assign n23520 = n2176 & n16037 ;
  assign n23521 = \s15_data_i[3]_pad  & n2176 ;
  assign n23522 = ~n2258 & n23521 ;
  assign n23523 = ~n23520 & ~n23522 ;
  assign n23524 = \s12_data_i[3]_pad  & n15007 ;
  assign n23525 = \s1_data_i[3]_pad  & n14640 ;
  assign n23526 = ~n23524 & ~n23525 ;
  assign n23527 = \s4_data_i[3]_pad  & n15030 ;
  assign n23528 = \s6_data_i[3]_pad  & n14681 ;
  assign n23529 = ~n23527 & ~n23528 ;
  assign n23530 = n23526 & n23529 ;
  assign n23531 = \s3_data_i[3]_pad  & n15026 ;
  assign n23532 = \s9_data_i[3]_pad  & n15042 ;
  assign n23533 = ~n23531 & ~n23532 ;
  assign n23534 = \s10_data_i[3]_pad  & n14999 ;
  assign n23535 = \s7_data_i[3]_pad  & n15038 ;
  assign n23536 = ~n23534 & ~n23535 ;
  assign n23537 = n23533 & n23536 ;
  assign n23538 = n23530 & n23537 ;
  assign n23539 = \s14_data_i[3]_pad  & n15015 ;
  assign n23540 = \s11_data_i[3]_pad  & n15003 ;
  assign n23541 = \s2_data_i[3]_pad  & n15022 ;
  assign n23542 = ~n23540 & ~n23541 ;
  assign n23543 = ~n23539 & n23542 ;
  assign n23544 = \s5_data_i[3]_pad  & n15034 ;
  assign n23545 = \s8_data_i[3]_pad  & n14690 ;
  assign n23546 = ~n23544 & ~n23545 ;
  assign n23547 = \s13_data_i[3]_pad  & n15011 ;
  assign n23548 = \s0_data_i[3]_pad  & n14634 ;
  assign n23549 = ~n23547 & ~n23548 ;
  assign n23550 = n23546 & n23549 ;
  assign n23551 = n23543 & n23550 ;
  assign n23552 = n23538 & n23551 ;
  assign n23553 = n23523 & n23552 ;
  assign n23554 = n2176 & n16074 ;
  assign n23555 = \s15_data_i[4]_pad  & n2176 ;
  assign n23556 = ~n2258 & n23555 ;
  assign n23557 = ~n23554 & ~n23556 ;
  assign n23558 = \s5_data_i[4]_pad  & n15034 ;
  assign n23559 = \s1_data_i[4]_pad  & n14640 ;
  assign n23560 = ~n23558 & ~n23559 ;
  assign n23561 = \s4_data_i[4]_pad  & n15030 ;
  assign n23562 = \s14_data_i[4]_pad  & n15015 ;
  assign n23563 = ~n23561 & ~n23562 ;
  assign n23564 = n23560 & n23563 ;
  assign n23565 = \s8_data_i[4]_pad  & n14690 ;
  assign n23566 = \s6_data_i[4]_pad  & n14681 ;
  assign n23567 = ~n23565 & ~n23566 ;
  assign n23568 = \s7_data_i[4]_pad  & n15038 ;
  assign n23569 = \s12_data_i[4]_pad  & n15007 ;
  assign n23570 = ~n23568 & ~n23569 ;
  assign n23571 = n23567 & n23570 ;
  assign n23572 = n23564 & n23571 ;
  assign n23573 = \s9_data_i[4]_pad  & n15042 ;
  assign n23574 = \s2_data_i[4]_pad  & n15022 ;
  assign n23575 = \s3_data_i[4]_pad  & n15026 ;
  assign n23576 = ~n23574 & ~n23575 ;
  assign n23577 = ~n23573 & n23576 ;
  assign n23578 = \s11_data_i[4]_pad  & n15003 ;
  assign n23579 = \s10_data_i[4]_pad  & n14999 ;
  assign n23580 = ~n23578 & ~n23579 ;
  assign n23581 = \s13_data_i[4]_pad  & n15011 ;
  assign n23582 = \s0_data_i[4]_pad  & n14634 ;
  assign n23583 = ~n23581 & ~n23582 ;
  assign n23584 = n23580 & n23583 ;
  assign n23585 = n23577 & n23584 ;
  assign n23586 = n23572 & n23585 ;
  assign n23587 = n23557 & n23586 ;
  assign n23588 = n2176 & n16111 ;
  assign n23589 = \s15_data_i[5]_pad  & n2176 ;
  assign n23590 = ~n2258 & n23589 ;
  assign n23591 = ~n23588 & ~n23590 ;
  assign n23592 = \s12_data_i[5]_pad  & n15007 ;
  assign n23593 = \s1_data_i[5]_pad  & n14640 ;
  assign n23594 = ~n23592 & ~n23593 ;
  assign n23595 = \s4_data_i[5]_pad  & n15030 ;
  assign n23596 = \s6_data_i[5]_pad  & n14681 ;
  assign n23597 = ~n23595 & ~n23596 ;
  assign n23598 = n23594 & n23597 ;
  assign n23599 = \s3_data_i[5]_pad  & n15026 ;
  assign n23600 = \s9_data_i[5]_pad  & n15042 ;
  assign n23601 = ~n23599 & ~n23600 ;
  assign n23602 = \s10_data_i[5]_pad  & n14999 ;
  assign n23603 = \s7_data_i[5]_pad  & n15038 ;
  assign n23604 = ~n23602 & ~n23603 ;
  assign n23605 = n23601 & n23604 ;
  assign n23606 = n23598 & n23605 ;
  assign n23607 = \s14_data_i[5]_pad  & n15015 ;
  assign n23608 = \s11_data_i[5]_pad  & n15003 ;
  assign n23609 = \s2_data_i[5]_pad  & n15022 ;
  assign n23610 = ~n23608 & ~n23609 ;
  assign n23611 = ~n23607 & n23610 ;
  assign n23612 = \s5_data_i[5]_pad  & n15034 ;
  assign n23613 = \s8_data_i[5]_pad  & n14690 ;
  assign n23614 = ~n23612 & ~n23613 ;
  assign n23615 = \s13_data_i[5]_pad  & n15011 ;
  assign n23616 = \s0_data_i[5]_pad  & n14634 ;
  assign n23617 = ~n23615 & ~n23616 ;
  assign n23618 = n23614 & n23617 ;
  assign n23619 = n23611 & n23618 ;
  assign n23620 = n23606 & n23619 ;
  assign n23621 = n23591 & n23620 ;
  assign n23622 = n2176 & n16148 ;
  assign n23623 = \s15_data_i[6]_pad  & n2176 ;
  assign n23624 = ~n2258 & n23623 ;
  assign n23625 = ~n23622 & ~n23624 ;
  assign n23626 = \s12_data_i[6]_pad  & n15007 ;
  assign n23627 = \s1_data_i[6]_pad  & n14640 ;
  assign n23628 = ~n23626 & ~n23627 ;
  assign n23629 = \s4_data_i[6]_pad  & n15030 ;
  assign n23630 = \s6_data_i[6]_pad  & n14681 ;
  assign n23631 = ~n23629 & ~n23630 ;
  assign n23632 = n23628 & n23631 ;
  assign n23633 = \s3_data_i[6]_pad  & n15026 ;
  assign n23634 = \s9_data_i[6]_pad  & n15042 ;
  assign n23635 = ~n23633 & ~n23634 ;
  assign n23636 = \s10_data_i[6]_pad  & n14999 ;
  assign n23637 = \s7_data_i[6]_pad  & n15038 ;
  assign n23638 = ~n23636 & ~n23637 ;
  assign n23639 = n23635 & n23638 ;
  assign n23640 = n23632 & n23639 ;
  assign n23641 = \s14_data_i[6]_pad  & n15015 ;
  assign n23642 = \s11_data_i[6]_pad  & n15003 ;
  assign n23643 = \s2_data_i[6]_pad  & n15022 ;
  assign n23644 = ~n23642 & ~n23643 ;
  assign n23645 = ~n23641 & n23644 ;
  assign n23646 = \s5_data_i[6]_pad  & n15034 ;
  assign n23647 = \s8_data_i[6]_pad  & n14690 ;
  assign n23648 = ~n23646 & ~n23647 ;
  assign n23649 = \s13_data_i[6]_pad  & n15011 ;
  assign n23650 = \s0_data_i[6]_pad  & n14634 ;
  assign n23651 = ~n23649 & ~n23650 ;
  assign n23652 = n23648 & n23651 ;
  assign n23653 = n23645 & n23652 ;
  assign n23654 = n23640 & n23653 ;
  assign n23655 = n23625 & n23654 ;
  assign n23656 = n2176 & n16185 ;
  assign n23657 = \s15_data_i[7]_pad  & n2176 ;
  assign n23658 = ~n2258 & n23657 ;
  assign n23659 = ~n23656 & ~n23658 ;
  assign n23660 = \s5_data_i[7]_pad  & n15034 ;
  assign n23661 = \s1_data_i[7]_pad  & n14640 ;
  assign n23662 = ~n23660 & ~n23661 ;
  assign n23663 = \s4_data_i[7]_pad  & n15030 ;
  assign n23664 = \s14_data_i[7]_pad  & n15015 ;
  assign n23665 = ~n23663 & ~n23664 ;
  assign n23666 = n23662 & n23665 ;
  assign n23667 = \s8_data_i[7]_pad  & n14690 ;
  assign n23668 = \s6_data_i[7]_pad  & n14681 ;
  assign n23669 = ~n23667 & ~n23668 ;
  assign n23670 = \s7_data_i[7]_pad  & n15038 ;
  assign n23671 = \s12_data_i[7]_pad  & n15007 ;
  assign n23672 = ~n23670 & ~n23671 ;
  assign n23673 = n23669 & n23672 ;
  assign n23674 = n23666 & n23673 ;
  assign n23675 = \s9_data_i[7]_pad  & n15042 ;
  assign n23676 = \s2_data_i[7]_pad  & n15022 ;
  assign n23677 = \s3_data_i[7]_pad  & n15026 ;
  assign n23678 = ~n23676 & ~n23677 ;
  assign n23679 = ~n23675 & n23678 ;
  assign n23680 = \s11_data_i[7]_pad  & n15003 ;
  assign n23681 = \s10_data_i[7]_pad  & n14999 ;
  assign n23682 = ~n23680 & ~n23681 ;
  assign n23683 = \s13_data_i[7]_pad  & n15011 ;
  assign n23684 = \s0_data_i[7]_pad  & n14634 ;
  assign n23685 = ~n23683 & ~n23684 ;
  assign n23686 = n23682 & n23685 ;
  assign n23687 = n23679 & n23686 ;
  assign n23688 = n23674 & n23687 ;
  assign n23689 = n23659 & n23688 ;
  assign n23690 = n2176 & n16222 ;
  assign n23691 = \s15_data_i[8]_pad  & n2176 ;
  assign n23692 = ~n2258 & n23691 ;
  assign n23693 = ~n23690 & ~n23692 ;
  assign n23694 = \s12_data_i[8]_pad  & n15007 ;
  assign n23695 = \s1_data_i[8]_pad  & n14640 ;
  assign n23696 = ~n23694 & ~n23695 ;
  assign n23697 = \s4_data_i[8]_pad  & n15030 ;
  assign n23698 = \s6_data_i[8]_pad  & n14681 ;
  assign n23699 = ~n23697 & ~n23698 ;
  assign n23700 = n23696 & n23699 ;
  assign n23701 = \s3_data_i[8]_pad  & n15026 ;
  assign n23702 = \s9_data_i[8]_pad  & n15042 ;
  assign n23703 = ~n23701 & ~n23702 ;
  assign n23704 = \s10_data_i[8]_pad  & n14999 ;
  assign n23705 = \s7_data_i[8]_pad  & n15038 ;
  assign n23706 = ~n23704 & ~n23705 ;
  assign n23707 = n23703 & n23706 ;
  assign n23708 = n23700 & n23707 ;
  assign n23709 = \s14_data_i[8]_pad  & n15015 ;
  assign n23710 = \s11_data_i[8]_pad  & n15003 ;
  assign n23711 = \s2_data_i[8]_pad  & n15022 ;
  assign n23712 = ~n23710 & ~n23711 ;
  assign n23713 = ~n23709 & n23712 ;
  assign n23714 = \s5_data_i[8]_pad  & n15034 ;
  assign n23715 = \s8_data_i[8]_pad  & n14690 ;
  assign n23716 = ~n23714 & ~n23715 ;
  assign n23717 = \s13_data_i[8]_pad  & n15011 ;
  assign n23718 = \s0_data_i[8]_pad  & n14634 ;
  assign n23719 = ~n23717 & ~n23718 ;
  assign n23720 = n23716 & n23719 ;
  assign n23721 = n23713 & n23720 ;
  assign n23722 = n23708 & n23721 ;
  assign n23723 = n23693 & n23722 ;
  assign n23724 = n2176 & n16259 ;
  assign n23725 = \s15_data_i[9]_pad  & n2176 ;
  assign n23726 = ~n2258 & n23725 ;
  assign n23727 = ~n23724 & ~n23726 ;
  assign n23728 = \s5_data_i[9]_pad  & n15034 ;
  assign n23729 = \s1_data_i[9]_pad  & n14640 ;
  assign n23730 = ~n23728 & ~n23729 ;
  assign n23731 = \s4_data_i[9]_pad  & n15030 ;
  assign n23732 = \s14_data_i[9]_pad  & n15015 ;
  assign n23733 = ~n23731 & ~n23732 ;
  assign n23734 = n23730 & n23733 ;
  assign n23735 = \s8_data_i[9]_pad  & n14690 ;
  assign n23736 = \s6_data_i[9]_pad  & n14681 ;
  assign n23737 = ~n23735 & ~n23736 ;
  assign n23738 = \s7_data_i[9]_pad  & n15038 ;
  assign n23739 = \s12_data_i[9]_pad  & n15007 ;
  assign n23740 = ~n23738 & ~n23739 ;
  assign n23741 = n23737 & n23740 ;
  assign n23742 = n23734 & n23741 ;
  assign n23743 = \s9_data_i[9]_pad  & n15042 ;
  assign n23744 = \s2_data_i[9]_pad  & n15022 ;
  assign n23745 = \s3_data_i[9]_pad  & n15026 ;
  assign n23746 = ~n23744 & ~n23745 ;
  assign n23747 = ~n23743 & n23746 ;
  assign n23748 = \s11_data_i[9]_pad  & n15003 ;
  assign n23749 = \s10_data_i[9]_pad  & n14999 ;
  assign n23750 = ~n23748 & ~n23749 ;
  assign n23751 = \s13_data_i[9]_pad  & n15011 ;
  assign n23752 = \s0_data_i[9]_pad  & n14634 ;
  assign n23753 = ~n23751 & ~n23752 ;
  assign n23754 = n23750 & n23753 ;
  assign n23755 = n23747 & n23754 ;
  assign n23756 = n23742 & n23755 ;
  assign n23757 = n23727 & n23756 ;
  assign n23758 = \s15_err_i_pad  & n22639 ;
  assign n23759 = ~n2258 & n23758 ;
  assign n23760 = \s2_err_i_pad  & n15022 ;
  assign n23761 = n14391 & n23760 ;
  assign n23762 = n14408 & n23761 ;
  assign n23763 = \s12_err_i_pad  & n15007 ;
  assign n23764 = n14140 & n23763 ;
  assign n23765 = n14148 & n23764 ;
  assign n23766 = ~n23762 & ~n23765 ;
  assign n23767 = \s13_err_i_pad  & n15011 ;
  assign n23768 = n14211 & n23767 ;
  assign n23769 = n14204 & n23768 ;
  assign n23770 = \s9_err_i_pad  & n15042 ;
  assign n23771 = n13847 & n23770 ;
  assign n23772 = n13864 & n23771 ;
  assign n23773 = ~n23769 & ~n23772 ;
  assign n23774 = n23766 & n23773 ;
  assign n23775 = \s6_err_i_pad  & n14681 ;
  assign n23776 = n13627 & n23775 ;
  assign n23777 = n13644 & n23776 ;
  assign n23778 = \s4_err_i_pad  & n15030 ;
  assign n23779 = n13467 & n23778 ;
  assign n23780 = n13492 & n23779 ;
  assign n23781 = ~n23777 & ~n23780 ;
  assign n23782 = \s0_err_i_pad  & n14634 ;
  assign n23783 = n14069 & n23782 ;
  assign n23784 = n14062 & n23783 ;
  assign n23785 = \s10_err_i_pad  & n14999 ;
  assign n23786 = n13928 & n23785 ;
  assign n23787 = n13936 & n23786 ;
  assign n23788 = ~n23784 & ~n23787 ;
  assign n23789 = n23781 & n23788 ;
  assign n23790 = n23774 & n23789 ;
  assign n23791 = \s1_err_i_pad  & n14640 ;
  assign n23792 = n14271 & n23791 ;
  assign n23793 = n14264 & n23792 ;
  assign n23794 = \s11_err_i_pad  & n15003 ;
  assign n23795 = n14009 & n23794 ;
  assign n23796 = n14026 & n23795 ;
  assign n23797 = \s7_err_i_pad  & n15038 ;
  assign n23798 = n13697 & n23797 ;
  assign n23799 = n13690 & n23798 ;
  assign n23800 = ~n23796 & ~n23799 ;
  assign n23801 = ~n23793 & n23800 ;
  assign n23802 = \s3_err_i_pad  & n15026 ;
  assign n23803 = n14451 & n23802 ;
  assign n23804 = n14468 & n23803 ;
  assign n23805 = \s5_err_i_pad  & n15034 ;
  assign n23806 = n13547 & n23805 ;
  assign n23807 = n13564 & n23806 ;
  assign n23808 = ~n23804 & ~n23807 ;
  assign n23809 = \s14_err_i_pad  & n15015 ;
  assign n23810 = n14331 & n23809 ;
  assign n23811 = n14348 & n23810 ;
  assign n23812 = \s8_err_i_pad  & n14690 ;
  assign n23813 = n13767 & n23812 ;
  assign n23814 = n13784 & n23813 ;
  assign n23815 = ~n23811 & ~n23814 ;
  assign n23816 = n23808 & n23815 ;
  assign n23817 = n23801 & n23816 ;
  assign n23818 = n23790 & n23817 ;
  assign n23819 = ~n23759 & n23818 ;
  assign n23820 = \s15_rty_i_pad  & n22639 ;
  assign n23821 = ~n2258 & n23820 ;
  assign n23822 = \s2_rty_i_pad  & n15022 ;
  assign n23823 = n14391 & n23822 ;
  assign n23824 = n14408 & n23823 ;
  assign n23825 = \s3_rty_i_pad  & n15026 ;
  assign n23826 = n14451 & n23825 ;
  assign n23827 = n14468 & n23826 ;
  assign n23828 = ~n23824 & ~n23827 ;
  assign n23829 = \s13_rty_i_pad  & n15011 ;
  assign n23830 = n14211 & n23829 ;
  assign n23831 = n14204 & n23830 ;
  assign n23832 = \s0_rty_i_pad  & n14634 ;
  assign n23833 = n14069 & n23832 ;
  assign n23834 = n14062 & n23833 ;
  assign n23835 = ~n23831 & ~n23834 ;
  assign n23836 = n23828 & n23835 ;
  assign n23837 = \s6_rty_i_pad  & n14681 ;
  assign n23838 = n13627 & n23837 ;
  assign n23839 = n13644 & n23838 ;
  assign n23840 = \s10_rty_i_pad  & n14999 ;
  assign n23841 = n13928 & n23840 ;
  assign n23842 = n13936 & n23841 ;
  assign n23843 = ~n23839 & ~n23842 ;
  assign n23844 = \s9_rty_i_pad  & n15042 ;
  assign n23845 = n13847 & n23844 ;
  assign n23846 = n13864 & n23845 ;
  assign n23847 = \s4_rty_i_pad  & n15030 ;
  assign n23848 = n13467 & n23847 ;
  assign n23849 = n13492 & n23848 ;
  assign n23850 = ~n23846 & ~n23849 ;
  assign n23851 = n23843 & n23850 ;
  assign n23852 = n23836 & n23851 ;
  assign n23853 = \s1_rty_i_pad  & n14640 ;
  assign n23854 = n14271 & n23853 ;
  assign n23855 = n14264 & n23854 ;
  assign n23856 = \s14_rty_i_pad  & n15015 ;
  assign n23857 = n14331 & n23856 ;
  assign n23858 = n14348 & n23857 ;
  assign n23859 = \s7_rty_i_pad  & n15038 ;
  assign n23860 = n13697 & n23859 ;
  assign n23861 = n13690 & n23860 ;
  assign n23862 = ~n23858 & ~n23861 ;
  assign n23863 = ~n23855 & n23862 ;
  assign n23864 = \s8_rty_i_pad  & n14690 ;
  assign n23865 = n13767 & n23864 ;
  assign n23866 = n13784 & n23865 ;
  assign n23867 = \s11_rty_i_pad  & n15003 ;
  assign n23868 = n14009 & n23867 ;
  assign n23869 = n14026 & n23868 ;
  assign n23870 = ~n23866 & ~n23869 ;
  assign n23871 = \s5_rty_i_pad  & n15034 ;
  assign n23872 = n13547 & n23871 ;
  assign n23873 = n13564 & n23872 ;
  assign n23874 = \s12_rty_i_pad  & n15007 ;
  assign n23875 = n14140 & n23874 ;
  assign n23876 = n14148 & n23875 ;
  assign n23877 = ~n23873 & ~n23876 ;
  assign n23878 = n23870 & n23877 ;
  assign n23879 = n23863 & n23878 ;
  assign n23880 = n23852 & n23879 ;
  assign n23881 = ~n23821 & n23880 ;
  assign n23882 = ~n1910 & n2170 ;
  assign n23883 = n1938 & n23882 ;
  assign n23884 = ~n13416 & n23883 ;
  assign n23885 = ~n15125 & n23884 ;
  assign n23886 = \s5_ack_i_pad  & n14675 ;
  assign n23887 = ~n13547 & n23886 ;
  assign n23888 = n13564 & n23887 ;
  assign n23889 = \s8_ack_i_pad  & n15086 ;
  assign n23890 = ~n13767 & n23889 ;
  assign n23891 = n13784 & n23890 ;
  assign n23892 = ~n23888 & ~n23891 ;
  assign n23893 = \s12_ack_i_pad  & n14685 ;
  assign n23894 = ~n14140 & n23893 ;
  assign n23895 = n14148 & n23894 ;
  assign n23896 = \s4_ack_i_pad  & n15074 ;
  assign n23897 = ~n13467 & n23896 ;
  assign n23898 = n13492 & n23897 ;
  assign n23899 = ~n23895 & ~n23898 ;
  assign n23900 = n23892 & n23899 ;
  assign n23901 = \s6_ack_i_pad  & n15078 ;
  assign n23902 = ~n13627 & n23901 ;
  assign n23903 = n13644 & n23902 ;
  assign n23904 = \s14_ack_i_pad  & n15059 ;
  assign n23905 = ~n14331 & n23904 ;
  assign n23906 = n14348 & n23905 ;
  assign n23907 = ~n23903 & ~n23906 ;
  assign n23908 = \s0_ack_i_pad  & n14647 ;
  assign n23909 = ~n14069 & n23908 ;
  assign n23910 = n14062 & n23909 ;
  assign n23911 = \s10_ack_i_pad  & n15047 ;
  assign n23912 = ~n13928 & n23911 ;
  assign n23913 = n13936 & n23912 ;
  assign n23914 = ~n23910 & ~n23913 ;
  assign n23915 = n23907 & n23914 ;
  assign n23916 = n23900 & n23915 ;
  assign n23917 = \s3_ack_i_pad  & n15070 ;
  assign n23918 = ~n14451 & n23917 ;
  assign n23919 = n14468 & n23918 ;
  assign n23920 = \s2_ack_i_pad  & n15066 ;
  assign n23921 = ~n14391 & n23920 ;
  assign n23922 = n14408 & n23921 ;
  assign n23923 = \s9_ack_i_pad  & n14666 ;
  assign n23924 = ~n13847 & n23923 ;
  assign n23925 = n13864 & n23924 ;
  assign n23926 = ~n23922 & ~n23925 ;
  assign n23927 = ~n23919 & n23926 ;
  assign n23928 = \s7_ack_i_pad  & n14671 ;
  assign n23929 = ~n13697 & n23928 ;
  assign n23930 = n13690 & n23929 ;
  assign n23931 = \s13_ack_i_pad  & n15055 ;
  assign n23932 = ~n14211 & n23931 ;
  assign n23933 = n14204 & n23932 ;
  assign n23934 = ~n23930 & ~n23933 ;
  assign n23935 = \s11_ack_i_pad  & n15051 ;
  assign n23936 = ~n14009 & n23935 ;
  assign n23937 = n14026 & n23936 ;
  assign n23938 = \s1_ack_i_pad  & n14653 ;
  assign n23939 = ~n14271 & n23938 ;
  assign n23940 = n14264 & n23939 ;
  assign n23941 = ~n23937 & ~n23940 ;
  assign n23942 = n23934 & n23941 ;
  assign n23943 = n23927 & n23942 ;
  assign n23944 = n23916 & n23943 ;
  assign n23945 = ~n23885 & n23944 ;
  assign n23946 = n2170 & n15192 ;
  assign n23947 = \s15_data_i[0]_pad  & n2170 ;
  assign n23948 = ~n2258 & n23947 ;
  assign n23949 = ~n23946 & ~n23948 ;
  assign n23950 = \s8_data_i[0]_pad  & n15086 ;
  assign n23951 = \s1_data_i[0]_pad  & n14653 ;
  assign n23952 = ~n23950 & ~n23951 ;
  assign n23953 = \s4_data_i[0]_pad  & n15074 ;
  assign n23954 = \s6_data_i[0]_pad  & n15078 ;
  assign n23955 = ~n23953 & ~n23954 ;
  assign n23956 = n23952 & n23955 ;
  assign n23957 = \s5_data_i[0]_pad  & n14675 ;
  assign n23958 = \s9_data_i[0]_pad  & n14666 ;
  assign n23959 = ~n23957 & ~n23958 ;
  assign n23960 = \s10_data_i[0]_pad  & n15047 ;
  assign n23961 = \s7_data_i[0]_pad  & n14671 ;
  assign n23962 = ~n23960 & ~n23961 ;
  assign n23963 = n23959 & n23962 ;
  assign n23964 = n23956 & n23963 ;
  assign n23965 = \s11_data_i[0]_pad  & n15051 ;
  assign n23966 = \s13_data_i[0]_pad  & n15055 ;
  assign n23967 = \s3_data_i[0]_pad  & n15070 ;
  assign n23968 = ~n23966 & ~n23967 ;
  assign n23969 = ~n23965 & n23968 ;
  assign n23970 = \s12_data_i[0]_pad  & n14685 ;
  assign n23971 = \s14_data_i[0]_pad  & n15059 ;
  assign n23972 = ~n23970 & ~n23971 ;
  assign n23973 = \s2_data_i[0]_pad  & n15066 ;
  assign n23974 = \s0_data_i[0]_pad  & n14647 ;
  assign n23975 = ~n23973 & ~n23974 ;
  assign n23976 = n23972 & n23975 ;
  assign n23977 = n23969 & n23976 ;
  assign n23978 = n23964 & n23977 ;
  assign n23979 = n23949 & n23978 ;
  assign n23980 = n2170 & n15229 ;
  assign n23981 = \s15_data_i[10]_pad  & n2170 ;
  assign n23982 = ~n2258 & n23981 ;
  assign n23983 = ~n23980 & ~n23982 ;
  assign n23984 = \s8_data_i[10]_pad  & n15086 ;
  assign n23985 = \s1_data_i[10]_pad  & n14653 ;
  assign n23986 = ~n23984 & ~n23985 ;
  assign n23987 = \s4_data_i[10]_pad  & n15074 ;
  assign n23988 = \s6_data_i[10]_pad  & n15078 ;
  assign n23989 = ~n23987 & ~n23988 ;
  assign n23990 = n23986 & n23989 ;
  assign n23991 = \s5_data_i[10]_pad  & n14675 ;
  assign n23992 = \s9_data_i[10]_pad  & n14666 ;
  assign n23993 = ~n23991 & ~n23992 ;
  assign n23994 = \s10_data_i[10]_pad  & n15047 ;
  assign n23995 = \s7_data_i[10]_pad  & n14671 ;
  assign n23996 = ~n23994 & ~n23995 ;
  assign n23997 = n23993 & n23996 ;
  assign n23998 = n23990 & n23997 ;
  assign n23999 = \s11_data_i[10]_pad  & n15051 ;
  assign n24000 = \s13_data_i[10]_pad  & n15055 ;
  assign n24001 = \s3_data_i[10]_pad  & n15070 ;
  assign n24002 = ~n24000 & ~n24001 ;
  assign n24003 = ~n23999 & n24002 ;
  assign n24004 = \s12_data_i[10]_pad  & n14685 ;
  assign n24005 = \s14_data_i[10]_pad  & n15059 ;
  assign n24006 = ~n24004 & ~n24005 ;
  assign n24007 = \s2_data_i[10]_pad  & n15066 ;
  assign n24008 = \s0_data_i[10]_pad  & n14647 ;
  assign n24009 = ~n24007 & ~n24008 ;
  assign n24010 = n24006 & n24009 ;
  assign n24011 = n24003 & n24010 ;
  assign n24012 = n23998 & n24011 ;
  assign n24013 = n23983 & n24012 ;
  assign n24014 = n2170 & n15266 ;
  assign n24015 = \s15_data_i[11]_pad  & n2170 ;
  assign n24016 = ~n2258 & n24015 ;
  assign n24017 = ~n24014 & ~n24016 ;
  assign n24018 = \s1_data_i[11]_pad  & n14653 ;
  assign n24019 = \s6_data_i[11]_pad  & n15078 ;
  assign n24020 = ~n24018 & ~n24019 ;
  assign n24021 = \s14_data_i[11]_pad  & n15059 ;
  assign n24022 = \s8_data_i[11]_pad  & n15086 ;
  assign n24023 = ~n24021 & ~n24022 ;
  assign n24024 = n24020 & n24023 ;
  assign n24025 = \s9_data_i[11]_pad  & n14666 ;
  assign n24026 = \s11_data_i[11]_pad  & n15051 ;
  assign n24027 = ~n24025 & ~n24026 ;
  assign n24028 = \s12_data_i[11]_pad  & n14685 ;
  assign n24029 = \s5_data_i[11]_pad  & n14675 ;
  assign n24030 = ~n24028 & ~n24029 ;
  assign n24031 = n24027 & n24030 ;
  assign n24032 = n24024 & n24031 ;
  assign n24033 = \s13_data_i[11]_pad  & n15055 ;
  assign n24034 = \s0_data_i[11]_pad  & n14647 ;
  assign n24035 = \s3_data_i[11]_pad  & n15070 ;
  assign n24036 = ~n24034 & ~n24035 ;
  assign n24037 = ~n24033 & n24036 ;
  assign n24038 = \s10_data_i[11]_pad  & n15047 ;
  assign n24039 = \s2_data_i[11]_pad  & n15066 ;
  assign n24040 = ~n24038 & ~n24039 ;
  assign n24041 = \s7_data_i[11]_pad  & n14671 ;
  assign n24042 = \s4_data_i[11]_pad  & n15074 ;
  assign n24043 = ~n24041 & ~n24042 ;
  assign n24044 = n24040 & n24043 ;
  assign n24045 = n24037 & n24044 ;
  assign n24046 = n24032 & n24045 ;
  assign n24047 = n24017 & n24046 ;
  assign n24048 = n2170 & n15303 ;
  assign n24049 = \s15_data_i[12]_pad  & n2170 ;
  assign n24050 = ~n2258 & n24049 ;
  assign n24051 = ~n24048 & ~n24050 ;
  assign n24052 = \s8_data_i[12]_pad  & n15086 ;
  assign n24053 = \s1_data_i[12]_pad  & n14653 ;
  assign n24054 = ~n24052 & ~n24053 ;
  assign n24055 = \s4_data_i[12]_pad  & n15074 ;
  assign n24056 = \s6_data_i[12]_pad  & n15078 ;
  assign n24057 = ~n24055 & ~n24056 ;
  assign n24058 = n24054 & n24057 ;
  assign n24059 = \s5_data_i[12]_pad  & n14675 ;
  assign n24060 = \s9_data_i[12]_pad  & n14666 ;
  assign n24061 = ~n24059 & ~n24060 ;
  assign n24062 = \s10_data_i[12]_pad  & n15047 ;
  assign n24063 = \s7_data_i[12]_pad  & n14671 ;
  assign n24064 = ~n24062 & ~n24063 ;
  assign n24065 = n24061 & n24064 ;
  assign n24066 = n24058 & n24065 ;
  assign n24067 = \s11_data_i[12]_pad  & n15051 ;
  assign n24068 = \s13_data_i[12]_pad  & n15055 ;
  assign n24069 = \s3_data_i[12]_pad  & n15070 ;
  assign n24070 = ~n24068 & ~n24069 ;
  assign n24071 = ~n24067 & n24070 ;
  assign n24072 = \s12_data_i[12]_pad  & n14685 ;
  assign n24073 = \s14_data_i[12]_pad  & n15059 ;
  assign n24074 = ~n24072 & ~n24073 ;
  assign n24075 = \s2_data_i[12]_pad  & n15066 ;
  assign n24076 = \s0_data_i[12]_pad  & n14647 ;
  assign n24077 = ~n24075 & ~n24076 ;
  assign n24078 = n24074 & n24077 ;
  assign n24079 = n24071 & n24078 ;
  assign n24080 = n24066 & n24079 ;
  assign n24081 = n24051 & n24080 ;
  assign n24082 = n2170 & n15340 ;
  assign n24083 = \s15_data_i[13]_pad  & n2170 ;
  assign n24084 = ~n2258 & n24083 ;
  assign n24085 = ~n24082 & ~n24084 ;
  assign n24086 = \s8_data_i[13]_pad  & n15086 ;
  assign n24087 = \s1_data_i[13]_pad  & n14653 ;
  assign n24088 = ~n24086 & ~n24087 ;
  assign n24089 = \s4_data_i[13]_pad  & n15074 ;
  assign n24090 = \s6_data_i[13]_pad  & n15078 ;
  assign n24091 = ~n24089 & ~n24090 ;
  assign n24092 = n24088 & n24091 ;
  assign n24093 = \s5_data_i[13]_pad  & n14675 ;
  assign n24094 = \s9_data_i[13]_pad  & n14666 ;
  assign n24095 = ~n24093 & ~n24094 ;
  assign n24096 = \s10_data_i[13]_pad  & n15047 ;
  assign n24097 = \s7_data_i[13]_pad  & n14671 ;
  assign n24098 = ~n24096 & ~n24097 ;
  assign n24099 = n24095 & n24098 ;
  assign n24100 = n24092 & n24099 ;
  assign n24101 = \s11_data_i[13]_pad  & n15051 ;
  assign n24102 = \s13_data_i[13]_pad  & n15055 ;
  assign n24103 = \s3_data_i[13]_pad  & n15070 ;
  assign n24104 = ~n24102 & ~n24103 ;
  assign n24105 = ~n24101 & n24104 ;
  assign n24106 = \s12_data_i[13]_pad  & n14685 ;
  assign n24107 = \s14_data_i[13]_pad  & n15059 ;
  assign n24108 = ~n24106 & ~n24107 ;
  assign n24109 = \s2_data_i[13]_pad  & n15066 ;
  assign n24110 = \s0_data_i[13]_pad  & n14647 ;
  assign n24111 = ~n24109 & ~n24110 ;
  assign n24112 = n24108 & n24111 ;
  assign n24113 = n24105 & n24112 ;
  assign n24114 = n24100 & n24113 ;
  assign n24115 = n24085 & n24114 ;
  assign n24116 = n2170 & n15377 ;
  assign n24117 = \s15_data_i[14]_pad  & n2170 ;
  assign n24118 = ~n2258 & n24117 ;
  assign n24119 = ~n24116 & ~n24118 ;
  assign n24120 = \s8_data_i[14]_pad  & n15086 ;
  assign n24121 = \s1_data_i[14]_pad  & n14653 ;
  assign n24122 = ~n24120 & ~n24121 ;
  assign n24123 = \s4_data_i[14]_pad  & n15074 ;
  assign n24124 = \s6_data_i[14]_pad  & n15078 ;
  assign n24125 = ~n24123 & ~n24124 ;
  assign n24126 = n24122 & n24125 ;
  assign n24127 = \s5_data_i[14]_pad  & n14675 ;
  assign n24128 = \s9_data_i[14]_pad  & n14666 ;
  assign n24129 = ~n24127 & ~n24128 ;
  assign n24130 = \s10_data_i[14]_pad  & n15047 ;
  assign n24131 = \s7_data_i[14]_pad  & n14671 ;
  assign n24132 = ~n24130 & ~n24131 ;
  assign n24133 = n24129 & n24132 ;
  assign n24134 = n24126 & n24133 ;
  assign n24135 = \s11_data_i[14]_pad  & n15051 ;
  assign n24136 = \s13_data_i[14]_pad  & n15055 ;
  assign n24137 = \s3_data_i[14]_pad  & n15070 ;
  assign n24138 = ~n24136 & ~n24137 ;
  assign n24139 = ~n24135 & n24138 ;
  assign n24140 = \s12_data_i[14]_pad  & n14685 ;
  assign n24141 = \s14_data_i[14]_pad  & n15059 ;
  assign n24142 = ~n24140 & ~n24141 ;
  assign n24143 = \s2_data_i[14]_pad  & n15066 ;
  assign n24144 = \s0_data_i[14]_pad  & n14647 ;
  assign n24145 = ~n24143 & ~n24144 ;
  assign n24146 = n24142 & n24145 ;
  assign n24147 = n24139 & n24146 ;
  assign n24148 = n24134 & n24147 ;
  assign n24149 = n24119 & n24148 ;
  assign n24150 = n2170 & n15414 ;
  assign n24151 = \s15_data_i[15]_pad  & n2170 ;
  assign n24152 = ~n2258 & n24151 ;
  assign n24153 = ~n24150 & ~n24152 ;
  assign n24154 = \s8_data_i[15]_pad  & n15086 ;
  assign n24155 = \s1_data_i[15]_pad  & n14653 ;
  assign n24156 = ~n24154 & ~n24155 ;
  assign n24157 = \s4_data_i[15]_pad  & n15074 ;
  assign n24158 = \s6_data_i[15]_pad  & n15078 ;
  assign n24159 = ~n24157 & ~n24158 ;
  assign n24160 = n24156 & n24159 ;
  assign n24161 = \s5_data_i[15]_pad  & n14675 ;
  assign n24162 = \s9_data_i[15]_pad  & n14666 ;
  assign n24163 = ~n24161 & ~n24162 ;
  assign n24164 = \s10_data_i[15]_pad  & n15047 ;
  assign n24165 = \s7_data_i[15]_pad  & n14671 ;
  assign n24166 = ~n24164 & ~n24165 ;
  assign n24167 = n24163 & n24166 ;
  assign n24168 = n24160 & n24167 ;
  assign n24169 = \s11_data_i[15]_pad  & n15051 ;
  assign n24170 = \s13_data_i[15]_pad  & n15055 ;
  assign n24171 = \s3_data_i[15]_pad  & n15070 ;
  assign n24172 = ~n24170 & ~n24171 ;
  assign n24173 = ~n24169 & n24172 ;
  assign n24174 = \s12_data_i[15]_pad  & n14685 ;
  assign n24175 = \s14_data_i[15]_pad  & n15059 ;
  assign n24176 = ~n24174 & ~n24175 ;
  assign n24177 = \s2_data_i[15]_pad  & n15066 ;
  assign n24178 = \s0_data_i[15]_pad  & n14647 ;
  assign n24179 = ~n24177 & ~n24178 ;
  assign n24180 = n24176 & n24179 ;
  assign n24181 = n24173 & n24180 ;
  assign n24182 = n24168 & n24181 ;
  assign n24183 = n24153 & n24182 ;
  assign n24184 = \s15_data_i[16]_pad  & n2170 ;
  assign n24185 = ~n2258 & n24184 ;
  assign n24186 = \s12_data_i[16]_pad  & n14685 ;
  assign n24187 = \s13_data_i[16]_pad  & n15055 ;
  assign n24188 = ~n24186 & ~n24187 ;
  assign n24189 = \s10_data_i[16]_pad  & n15047 ;
  assign n24190 = \s1_data_i[16]_pad  & n14653 ;
  assign n24191 = ~n24189 & ~n24190 ;
  assign n24192 = n24188 & n24191 ;
  assign n24193 = \s5_data_i[16]_pad  & n14675 ;
  assign n24194 = \s6_data_i[16]_pad  & n15078 ;
  assign n24195 = ~n24193 & ~n24194 ;
  assign n24196 = \s7_data_i[16]_pad  & n14671 ;
  assign n24197 = \s2_data_i[16]_pad  & n15066 ;
  assign n24198 = ~n24196 & ~n24197 ;
  assign n24199 = n24195 & n24198 ;
  assign n24200 = n24192 & n24199 ;
  assign n24201 = \s14_data_i[16]_pad  & n15059 ;
  assign n24202 = \s4_data_i[16]_pad  & n15074 ;
  assign n24203 = \s3_data_i[16]_pad  & n15070 ;
  assign n24204 = ~n24202 & ~n24203 ;
  assign n24205 = ~n24201 & n24204 ;
  assign n24206 = \s8_data_i[16]_pad  & n15086 ;
  assign n24207 = \s11_data_i[16]_pad  & n15051 ;
  assign n24208 = ~n24206 & ~n24207 ;
  assign n24209 = \s0_data_i[16]_pad  & n14647 ;
  assign n24210 = \s9_data_i[16]_pad  & n14666 ;
  assign n24211 = ~n24209 & ~n24210 ;
  assign n24212 = n24208 & n24211 ;
  assign n24213 = n24205 & n24212 ;
  assign n24214 = n24200 & n24213 ;
  assign n24215 = ~n24185 & n24214 ;
  assign n24216 = \s15_data_i[17]_pad  & n2170 ;
  assign n24217 = ~n2258 & n24216 ;
  assign n24218 = \s12_data_i[17]_pad  & n14685 ;
  assign n24219 = \s13_data_i[17]_pad  & n15055 ;
  assign n24220 = ~n24218 & ~n24219 ;
  assign n24221 = \s10_data_i[17]_pad  & n15047 ;
  assign n24222 = \s1_data_i[17]_pad  & n14653 ;
  assign n24223 = ~n24221 & ~n24222 ;
  assign n24224 = n24220 & n24223 ;
  assign n24225 = \s5_data_i[17]_pad  & n14675 ;
  assign n24226 = \s6_data_i[17]_pad  & n15078 ;
  assign n24227 = ~n24225 & ~n24226 ;
  assign n24228 = \s7_data_i[17]_pad  & n14671 ;
  assign n24229 = \s2_data_i[17]_pad  & n15066 ;
  assign n24230 = ~n24228 & ~n24229 ;
  assign n24231 = n24227 & n24230 ;
  assign n24232 = n24224 & n24231 ;
  assign n24233 = \s14_data_i[17]_pad  & n15059 ;
  assign n24234 = \s4_data_i[17]_pad  & n15074 ;
  assign n24235 = \s3_data_i[17]_pad  & n15070 ;
  assign n24236 = ~n24234 & ~n24235 ;
  assign n24237 = ~n24233 & n24236 ;
  assign n24238 = \s8_data_i[17]_pad  & n15086 ;
  assign n24239 = \s11_data_i[17]_pad  & n15051 ;
  assign n24240 = ~n24238 & ~n24239 ;
  assign n24241 = \s0_data_i[17]_pad  & n14647 ;
  assign n24242 = \s9_data_i[17]_pad  & n14666 ;
  assign n24243 = ~n24241 & ~n24242 ;
  assign n24244 = n24240 & n24243 ;
  assign n24245 = n24237 & n24244 ;
  assign n24246 = n24232 & n24245 ;
  assign n24247 = ~n24217 & n24246 ;
  assign n24248 = \s15_data_i[18]_pad  & n2170 ;
  assign n24249 = ~n2258 & n24248 ;
  assign n24250 = \s12_data_i[18]_pad  & n14685 ;
  assign n24251 = \s13_data_i[18]_pad  & n15055 ;
  assign n24252 = ~n24250 & ~n24251 ;
  assign n24253 = \s10_data_i[18]_pad  & n15047 ;
  assign n24254 = \s1_data_i[18]_pad  & n14653 ;
  assign n24255 = ~n24253 & ~n24254 ;
  assign n24256 = n24252 & n24255 ;
  assign n24257 = \s5_data_i[18]_pad  & n14675 ;
  assign n24258 = \s6_data_i[18]_pad  & n15078 ;
  assign n24259 = ~n24257 & ~n24258 ;
  assign n24260 = \s7_data_i[18]_pad  & n14671 ;
  assign n24261 = \s2_data_i[18]_pad  & n15066 ;
  assign n24262 = ~n24260 & ~n24261 ;
  assign n24263 = n24259 & n24262 ;
  assign n24264 = n24256 & n24263 ;
  assign n24265 = \s14_data_i[18]_pad  & n15059 ;
  assign n24266 = \s4_data_i[18]_pad  & n15074 ;
  assign n24267 = \s3_data_i[18]_pad  & n15070 ;
  assign n24268 = ~n24266 & ~n24267 ;
  assign n24269 = ~n24265 & n24268 ;
  assign n24270 = \s8_data_i[18]_pad  & n15086 ;
  assign n24271 = \s11_data_i[18]_pad  & n15051 ;
  assign n24272 = ~n24270 & ~n24271 ;
  assign n24273 = \s0_data_i[18]_pad  & n14647 ;
  assign n24274 = \s9_data_i[18]_pad  & n14666 ;
  assign n24275 = ~n24273 & ~n24274 ;
  assign n24276 = n24272 & n24275 ;
  assign n24277 = n24269 & n24276 ;
  assign n24278 = n24264 & n24277 ;
  assign n24279 = ~n24249 & n24278 ;
  assign n24280 = \s15_data_i[19]_pad  & n2170 ;
  assign n24281 = ~n2258 & n24280 ;
  assign n24282 = \s12_data_i[19]_pad  & n14685 ;
  assign n24283 = \s13_data_i[19]_pad  & n15055 ;
  assign n24284 = ~n24282 & ~n24283 ;
  assign n24285 = \s10_data_i[19]_pad  & n15047 ;
  assign n24286 = \s1_data_i[19]_pad  & n14653 ;
  assign n24287 = ~n24285 & ~n24286 ;
  assign n24288 = n24284 & n24287 ;
  assign n24289 = \s5_data_i[19]_pad  & n14675 ;
  assign n24290 = \s6_data_i[19]_pad  & n15078 ;
  assign n24291 = ~n24289 & ~n24290 ;
  assign n24292 = \s7_data_i[19]_pad  & n14671 ;
  assign n24293 = \s2_data_i[19]_pad  & n15066 ;
  assign n24294 = ~n24292 & ~n24293 ;
  assign n24295 = n24291 & n24294 ;
  assign n24296 = n24288 & n24295 ;
  assign n24297 = \s14_data_i[19]_pad  & n15059 ;
  assign n24298 = \s4_data_i[19]_pad  & n15074 ;
  assign n24299 = \s3_data_i[19]_pad  & n15070 ;
  assign n24300 = ~n24298 & ~n24299 ;
  assign n24301 = ~n24297 & n24300 ;
  assign n24302 = \s8_data_i[19]_pad  & n15086 ;
  assign n24303 = \s11_data_i[19]_pad  & n15051 ;
  assign n24304 = ~n24302 & ~n24303 ;
  assign n24305 = \s0_data_i[19]_pad  & n14647 ;
  assign n24306 = \s9_data_i[19]_pad  & n14666 ;
  assign n24307 = ~n24305 & ~n24306 ;
  assign n24308 = n24304 & n24307 ;
  assign n24309 = n24301 & n24308 ;
  assign n24310 = n24296 & n24309 ;
  assign n24311 = ~n24281 & n24310 ;
  assign n24312 = n2170 & n15579 ;
  assign n24313 = \s15_data_i[1]_pad  & n2170 ;
  assign n24314 = ~n2258 & n24313 ;
  assign n24315 = ~n24312 & ~n24314 ;
  assign n24316 = \s8_data_i[1]_pad  & n15086 ;
  assign n24317 = \s1_data_i[1]_pad  & n14653 ;
  assign n24318 = ~n24316 & ~n24317 ;
  assign n24319 = \s4_data_i[1]_pad  & n15074 ;
  assign n24320 = \s6_data_i[1]_pad  & n15078 ;
  assign n24321 = ~n24319 & ~n24320 ;
  assign n24322 = n24318 & n24321 ;
  assign n24323 = \s5_data_i[1]_pad  & n14675 ;
  assign n24324 = \s9_data_i[1]_pad  & n14666 ;
  assign n24325 = ~n24323 & ~n24324 ;
  assign n24326 = \s10_data_i[1]_pad  & n15047 ;
  assign n24327 = \s7_data_i[1]_pad  & n14671 ;
  assign n24328 = ~n24326 & ~n24327 ;
  assign n24329 = n24325 & n24328 ;
  assign n24330 = n24322 & n24329 ;
  assign n24331 = \s11_data_i[1]_pad  & n15051 ;
  assign n24332 = \s13_data_i[1]_pad  & n15055 ;
  assign n24333 = \s3_data_i[1]_pad  & n15070 ;
  assign n24334 = ~n24332 & ~n24333 ;
  assign n24335 = ~n24331 & n24334 ;
  assign n24336 = \s12_data_i[1]_pad  & n14685 ;
  assign n24337 = \s14_data_i[1]_pad  & n15059 ;
  assign n24338 = ~n24336 & ~n24337 ;
  assign n24339 = \s2_data_i[1]_pad  & n15066 ;
  assign n24340 = \s0_data_i[1]_pad  & n14647 ;
  assign n24341 = ~n24339 & ~n24340 ;
  assign n24342 = n24338 & n24341 ;
  assign n24343 = n24335 & n24342 ;
  assign n24344 = n24330 & n24343 ;
  assign n24345 = n24315 & n24344 ;
  assign n24346 = \s15_data_i[20]_pad  & n2170 ;
  assign n24347 = ~n2258 & n24346 ;
  assign n24348 = \s12_data_i[20]_pad  & n14685 ;
  assign n24349 = \s13_data_i[20]_pad  & n15055 ;
  assign n24350 = ~n24348 & ~n24349 ;
  assign n24351 = \s10_data_i[20]_pad  & n15047 ;
  assign n24352 = \s1_data_i[20]_pad  & n14653 ;
  assign n24353 = ~n24351 & ~n24352 ;
  assign n24354 = n24350 & n24353 ;
  assign n24355 = \s5_data_i[20]_pad  & n14675 ;
  assign n24356 = \s6_data_i[20]_pad  & n15078 ;
  assign n24357 = ~n24355 & ~n24356 ;
  assign n24358 = \s7_data_i[20]_pad  & n14671 ;
  assign n24359 = \s2_data_i[20]_pad  & n15066 ;
  assign n24360 = ~n24358 & ~n24359 ;
  assign n24361 = n24357 & n24360 ;
  assign n24362 = n24354 & n24361 ;
  assign n24363 = \s14_data_i[20]_pad  & n15059 ;
  assign n24364 = \s4_data_i[20]_pad  & n15074 ;
  assign n24365 = \s3_data_i[20]_pad  & n15070 ;
  assign n24366 = ~n24364 & ~n24365 ;
  assign n24367 = ~n24363 & n24366 ;
  assign n24368 = \s8_data_i[20]_pad  & n15086 ;
  assign n24369 = \s11_data_i[20]_pad  & n15051 ;
  assign n24370 = ~n24368 & ~n24369 ;
  assign n24371 = \s0_data_i[20]_pad  & n14647 ;
  assign n24372 = \s9_data_i[20]_pad  & n14666 ;
  assign n24373 = ~n24371 & ~n24372 ;
  assign n24374 = n24370 & n24373 ;
  assign n24375 = n24367 & n24374 ;
  assign n24376 = n24362 & n24375 ;
  assign n24377 = ~n24347 & n24376 ;
  assign n24378 = \s15_data_i[21]_pad  & n2170 ;
  assign n24379 = ~n2258 & n24378 ;
  assign n24380 = \s12_data_i[21]_pad  & n14685 ;
  assign n24381 = \s13_data_i[21]_pad  & n15055 ;
  assign n24382 = ~n24380 & ~n24381 ;
  assign n24383 = \s10_data_i[21]_pad  & n15047 ;
  assign n24384 = \s1_data_i[21]_pad  & n14653 ;
  assign n24385 = ~n24383 & ~n24384 ;
  assign n24386 = n24382 & n24385 ;
  assign n24387 = \s5_data_i[21]_pad  & n14675 ;
  assign n24388 = \s6_data_i[21]_pad  & n15078 ;
  assign n24389 = ~n24387 & ~n24388 ;
  assign n24390 = \s7_data_i[21]_pad  & n14671 ;
  assign n24391 = \s2_data_i[21]_pad  & n15066 ;
  assign n24392 = ~n24390 & ~n24391 ;
  assign n24393 = n24389 & n24392 ;
  assign n24394 = n24386 & n24393 ;
  assign n24395 = \s14_data_i[21]_pad  & n15059 ;
  assign n24396 = \s4_data_i[21]_pad  & n15074 ;
  assign n24397 = \s3_data_i[21]_pad  & n15070 ;
  assign n24398 = ~n24396 & ~n24397 ;
  assign n24399 = ~n24395 & n24398 ;
  assign n24400 = \s8_data_i[21]_pad  & n15086 ;
  assign n24401 = \s11_data_i[21]_pad  & n15051 ;
  assign n24402 = ~n24400 & ~n24401 ;
  assign n24403 = \s0_data_i[21]_pad  & n14647 ;
  assign n24404 = \s9_data_i[21]_pad  & n14666 ;
  assign n24405 = ~n24403 & ~n24404 ;
  assign n24406 = n24402 & n24405 ;
  assign n24407 = n24399 & n24406 ;
  assign n24408 = n24394 & n24407 ;
  assign n24409 = ~n24379 & n24408 ;
  assign n24410 = \s15_data_i[22]_pad  & n2170 ;
  assign n24411 = ~n2258 & n24410 ;
  assign n24412 = \s12_data_i[22]_pad  & n14685 ;
  assign n24413 = \s13_data_i[22]_pad  & n15055 ;
  assign n24414 = ~n24412 & ~n24413 ;
  assign n24415 = \s10_data_i[22]_pad  & n15047 ;
  assign n24416 = \s1_data_i[22]_pad  & n14653 ;
  assign n24417 = ~n24415 & ~n24416 ;
  assign n24418 = n24414 & n24417 ;
  assign n24419 = \s5_data_i[22]_pad  & n14675 ;
  assign n24420 = \s6_data_i[22]_pad  & n15078 ;
  assign n24421 = ~n24419 & ~n24420 ;
  assign n24422 = \s7_data_i[22]_pad  & n14671 ;
  assign n24423 = \s2_data_i[22]_pad  & n15066 ;
  assign n24424 = ~n24422 & ~n24423 ;
  assign n24425 = n24421 & n24424 ;
  assign n24426 = n24418 & n24425 ;
  assign n24427 = \s14_data_i[22]_pad  & n15059 ;
  assign n24428 = \s4_data_i[22]_pad  & n15074 ;
  assign n24429 = \s3_data_i[22]_pad  & n15070 ;
  assign n24430 = ~n24428 & ~n24429 ;
  assign n24431 = ~n24427 & n24430 ;
  assign n24432 = \s8_data_i[22]_pad  & n15086 ;
  assign n24433 = \s11_data_i[22]_pad  & n15051 ;
  assign n24434 = ~n24432 & ~n24433 ;
  assign n24435 = \s0_data_i[22]_pad  & n14647 ;
  assign n24436 = \s9_data_i[22]_pad  & n14666 ;
  assign n24437 = ~n24435 & ~n24436 ;
  assign n24438 = n24434 & n24437 ;
  assign n24439 = n24431 & n24438 ;
  assign n24440 = n24426 & n24439 ;
  assign n24441 = ~n24411 & n24440 ;
  assign n24442 = \s15_data_i[23]_pad  & n2170 ;
  assign n24443 = ~n2258 & n24442 ;
  assign n24444 = \s12_data_i[23]_pad  & n14685 ;
  assign n24445 = \s13_data_i[23]_pad  & n15055 ;
  assign n24446 = ~n24444 & ~n24445 ;
  assign n24447 = \s10_data_i[23]_pad  & n15047 ;
  assign n24448 = \s1_data_i[23]_pad  & n14653 ;
  assign n24449 = ~n24447 & ~n24448 ;
  assign n24450 = n24446 & n24449 ;
  assign n24451 = \s5_data_i[23]_pad  & n14675 ;
  assign n24452 = \s6_data_i[23]_pad  & n15078 ;
  assign n24453 = ~n24451 & ~n24452 ;
  assign n24454 = \s7_data_i[23]_pad  & n14671 ;
  assign n24455 = \s2_data_i[23]_pad  & n15066 ;
  assign n24456 = ~n24454 & ~n24455 ;
  assign n24457 = n24453 & n24456 ;
  assign n24458 = n24450 & n24457 ;
  assign n24459 = \s14_data_i[23]_pad  & n15059 ;
  assign n24460 = \s4_data_i[23]_pad  & n15074 ;
  assign n24461 = \s3_data_i[23]_pad  & n15070 ;
  assign n24462 = ~n24460 & ~n24461 ;
  assign n24463 = ~n24459 & n24462 ;
  assign n24464 = \s8_data_i[23]_pad  & n15086 ;
  assign n24465 = \s11_data_i[23]_pad  & n15051 ;
  assign n24466 = ~n24464 & ~n24465 ;
  assign n24467 = \s0_data_i[23]_pad  & n14647 ;
  assign n24468 = \s9_data_i[23]_pad  & n14666 ;
  assign n24469 = ~n24467 & ~n24468 ;
  assign n24470 = n24466 & n24469 ;
  assign n24471 = n24463 & n24470 ;
  assign n24472 = n24458 & n24471 ;
  assign n24473 = ~n24443 & n24472 ;
  assign n24474 = \s15_data_i[24]_pad  & n2170 ;
  assign n24475 = ~n2258 & n24474 ;
  assign n24476 = \s12_data_i[24]_pad  & n14685 ;
  assign n24477 = \s13_data_i[24]_pad  & n15055 ;
  assign n24478 = ~n24476 & ~n24477 ;
  assign n24479 = \s10_data_i[24]_pad  & n15047 ;
  assign n24480 = \s1_data_i[24]_pad  & n14653 ;
  assign n24481 = ~n24479 & ~n24480 ;
  assign n24482 = n24478 & n24481 ;
  assign n24483 = \s5_data_i[24]_pad  & n14675 ;
  assign n24484 = \s6_data_i[24]_pad  & n15078 ;
  assign n24485 = ~n24483 & ~n24484 ;
  assign n24486 = \s7_data_i[24]_pad  & n14671 ;
  assign n24487 = \s2_data_i[24]_pad  & n15066 ;
  assign n24488 = ~n24486 & ~n24487 ;
  assign n24489 = n24485 & n24488 ;
  assign n24490 = n24482 & n24489 ;
  assign n24491 = \s14_data_i[24]_pad  & n15059 ;
  assign n24492 = \s4_data_i[24]_pad  & n15074 ;
  assign n24493 = \s3_data_i[24]_pad  & n15070 ;
  assign n24494 = ~n24492 & ~n24493 ;
  assign n24495 = ~n24491 & n24494 ;
  assign n24496 = \s8_data_i[24]_pad  & n15086 ;
  assign n24497 = \s11_data_i[24]_pad  & n15051 ;
  assign n24498 = ~n24496 & ~n24497 ;
  assign n24499 = \s0_data_i[24]_pad  & n14647 ;
  assign n24500 = \s9_data_i[24]_pad  & n14666 ;
  assign n24501 = ~n24499 & ~n24500 ;
  assign n24502 = n24498 & n24501 ;
  assign n24503 = n24495 & n24502 ;
  assign n24504 = n24490 & n24503 ;
  assign n24505 = ~n24475 & n24504 ;
  assign n24506 = \s15_data_i[25]_pad  & n2170 ;
  assign n24507 = ~n2258 & n24506 ;
  assign n24508 = \s12_data_i[25]_pad  & n14685 ;
  assign n24509 = \s13_data_i[25]_pad  & n15055 ;
  assign n24510 = ~n24508 & ~n24509 ;
  assign n24511 = \s10_data_i[25]_pad  & n15047 ;
  assign n24512 = \s1_data_i[25]_pad  & n14653 ;
  assign n24513 = ~n24511 & ~n24512 ;
  assign n24514 = n24510 & n24513 ;
  assign n24515 = \s5_data_i[25]_pad  & n14675 ;
  assign n24516 = \s6_data_i[25]_pad  & n15078 ;
  assign n24517 = ~n24515 & ~n24516 ;
  assign n24518 = \s7_data_i[25]_pad  & n14671 ;
  assign n24519 = \s2_data_i[25]_pad  & n15066 ;
  assign n24520 = ~n24518 & ~n24519 ;
  assign n24521 = n24517 & n24520 ;
  assign n24522 = n24514 & n24521 ;
  assign n24523 = \s14_data_i[25]_pad  & n15059 ;
  assign n24524 = \s4_data_i[25]_pad  & n15074 ;
  assign n24525 = \s3_data_i[25]_pad  & n15070 ;
  assign n24526 = ~n24524 & ~n24525 ;
  assign n24527 = ~n24523 & n24526 ;
  assign n24528 = \s8_data_i[25]_pad  & n15086 ;
  assign n24529 = \s11_data_i[25]_pad  & n15051 ;
  assign n24530 = ~n24528 & ~n24529 ;
  assign n24531 = \s0_data_i[25]_pad  & n14647 ;
  assign n24532 = \s9_data_i[25]_pad  & n14666 ;
  assign n24533 = ~n24531 & ~n24532 ;
  assign n24534 = n24530 & n24533 ;
  assign n24535 = n24527 & n24534 ;
  assign n24536 = n24522 & n24535 ;
  assign n24537 = ~n24507 & n24536 ;
  assign n24538 = \s15_data_i[26]_pad  & n2170 ;
  assign n24539 = ~n2258 & n24538 ;
  assign n24540 = \s12_data_i[26]_pad  & n14685 ;
  assign n24541 = \s13_data_i[26]_pad  & n15055 ;
  assign n24542 = ~n24540 & ~n24541 ;
  assign n24543 = \s10_data_i[26]_pad  & n15047 ;
  assign n24544 = \s1_data_i[26]_pad  & n14653 ;
  assign n24545 = ~n24543 & ~n24544 ;
  assign n24546 = n24542 & n24545 ;
  assign n24547 = \s5_data_i[26]_pad  & n14675 ;
  assign n24548 = \s6_data_i[26]_pad  & n15078 ;
  assign n24549 = ~n24547 & ~n24548 ;
  assign n24550 = \s7_data_i[26]_pad  & n14671 ;
  assign n24551 = \s2_data_i[26]_pad  & n15066 ;
  assign n24552 = ~n24550 & ~n24551 ;
  assign n24553 = n24549 & n24552 ;
  assign n24554 = n24546 & n24553 ;
  assign n24555 = \s14_data_i[26]_pad  & n15059 ;
  assign n24556 = \s4_data_i[26]_pad  & n15074 ;
  assign n24557 = \s3_data_i[26]_pad  & n15070 ;
  assign n24558 = ~n24556 & ~n24557 ;
  assign n24559 = ~n24555 & n24558 ;
  assign n24560 = \s8_data_i[26]_pad  & n15086 ;
  assign n24561 = \s11_data_i[26]_pad  & n15051 ;
  assign n24562 = ~n24560 & ~n24561 ;
  assign n24563 = \s0_data_i[26]_pad  & n14647 ;
  assign n24564 = \s9_data_i[26]_pad  & n14666 ;
  assign n24565 = ~n24563 & ~n24564 ;
  assign n24566 = n24562 & n24565 ;
  assign n24567 = n24559 & n24566 ;
  assign n24568 = n24554 & n24567 ;
  assign n24569 = ~n24539 & n24568 ;
  assign n24570 = \s15_data_i[27]_pad  & n2170 ;
  assign n24571 = ~n2258 & n24570 ;
  assign n24572 = \s12_data_i[27]_pad  & n14685 ;
  assign n24573 = \s13_data_i[27]_pad  & n15055 ;
  assign n24574 = ~n24572 & ~n24573 ;
  assign n24575 = \s10_data_i[27]_pad  & n15047 ;
  assign n24576 = \s1_data_i[27]_pad  & n14653 ;
  assign n24577 = ~n24575 & ~n24576 ;
  assign n24578 = n24574 & n24577 ;
  assign n24579 = \s5_data_i[27]_pad  & n14675 ;
  assign n24580 = \s6_data_i[27]_pad  & n15078 ;
  assign n24581 = ~n24579 & ~n24580 ;
  assign n24582 = \s7_data_i[27]_pad  & n14671 ;
  assign n24583 = \s2_data_i[27]_pad  & n15066 ;
  assign n24584 = ~n24582 & ~n24583 ;
  assign n24585 = n24581 & n24584 ;
  assign n24586 = n24578 & n24585 ;
  assign n24587 = \s14_data_i[27]_pad  & n15059 ;
  assign n24588 = \s4_data_i[27]_pad  & n15074 ;
  assign n24589 = \s3_data_i[27]_pad  & n15070 ;
  assign n24590 = ~n24588 & ~n24589 ;
  assign n24591 = ~n24587 & n24590 ;
  assign n24592 = \s8_data_i[27]_pad  & n15086 ;
  assign n24593 = \s11_data_i[27]_pad  & n15051 ;
  assign n24594 = ~n24592 & ~n24593 ;
  assign n24595 = \s0_data_i[27]_pad  & n14647 ;
  assign n24596 = \s9_data_i[27]_pad  & n14666 ;
  assign n24597 = ~n24595 & ~n24596 ;
  assign n24598 = n24594 & n24597 ;
  assign n24599 = n24591 & n24598 ;
  assign n24600 = n24586 & n24599 ;
  assign n24601 = ~n24571 & n24600 ;
  assign n24602 = \s15_data_i[28]_pad  & n2170 ;
  assign n24603 = ~n2258 & n24602 ;
  assign n24604 = \s12_data_i[28]_pad  & n14685 ;
  assign n24605 = \s13_data_i[28]_pad  & n15055 ;
  assign n24606 = ~n24604 & ~n24605 ;
  assign n24607 = \s10_data_i[28]_pad  & n15047 ;
  assign n24608 = \s1_data_i[28]_pad  & n14653 ;
  assign n24609 = ~n24607 & ~n24608 ;
  assign n24610 = n24606 & n24609 ;
  assign n24611 = \s5_data_i[28]_pad  & n14675 ;
  assign n24612 = \s6_data_i[28]_pad  & n15078 ;
  assign n24613 = ~n24611 & ~n24612 ;
  assign n24614 = \s7_data_i[28]_pad  & n14671 ;
  assign n24615 = \s2_data_i[28]_pad  & n15066 ;
  assign n24616 = ~n24614 & ~n24615 ;
  assign n24617 = n24613 & n24616 ;
  assign n24618 = n24610 & n24617 ;
  assign n24619 = \s14_data_i[28]_pad  & n15059 ;
  assign n24620 = \s4_data_i[28]_pad  & n15074 ;
  assign n24621 = \s3_data_i[28]_pad  & n15070 ;
  assign n24622 = ~n24620 & ~n24621 ;
  assign n24623 = ~n24619 & n24622 ;
  assign n24624 = \s8_data_i[28]_pad  & n15086 ;
  assign n24625 = \s11_data_i[28]_pad  & n15051 ;
  assign n24626 = ~n24624 & ~n24625 ;
  assign n24627 = \s0_data_i[28]_pad  & n14647 ;
  assign n24628 = \s9_data_i[28]_pad  & n14666 ;
  assign n24629 = ~n24627 & ~n24628 ;
  assign n24630 = n24626 & n24629 ;
  assign n24631 = n24623 & n24630 ;
  assign n24632 = n24618 & n24631 ;
  assign n24633 = ~n24603 & n24632 ;
  assign n24634 = \s15_data_i[29]_pad  & n2170 ;
  assign n24635 = ~n2258 & n24634 ;
  assign n24636 = \s12_data_i[29]_pad  & n14685 ;
  assign n24637 = \s13_data_i[29]_pad  & n15055 ;
  assign n24638 = ~n24636 & ~n24637 ;
  assign n24639 = \s10_data_i[29]_pad  & n15047 ;
  assign n24640 = \s1_data_i[29]_pad  & n14653 ;
  assign n24641 = ~n24639 & ~n24640 ;
  assign n24642 = n24638 & n24641 ;
  assign n24643 = \s5_data_i[29]_pad  & n14675 ;
  assign n24644 = \s6_data_i[29]_pad  & n15078 ;
  assign n24645 = ~n24643 & ~n24644 ;
  assign n24646 = \s7_data_i[29]_pad  & n14671 ;
  assign n24647 = \s2_data_i[29]_pad  & n15066 ;
  assign n24648 = ~n24646 & ~n24647 ;
  assign n24649 = n24645 & n24648 ;
  assign n24650 = n24642 & n24649 ;
  assign n24651 = \s14_data_i[29]_pad  & n15059 ;
  assign n24652 = \s4_data_i[29]_pad  & n15074 ;
  assign n24653 = \s3_data_i[29]_pad  & n15070 ;
  assign n24654 = ~n24652 & ~n24653 ;
  assign n24655 = ~n24651 & n24654 ;
  assign n24656 = \s8_data_i[29]_pad  & n15086 ;
  assign n24657 = \s11_data_i[29]_pad  & n15051 ;
  assign n24658 = ~n24656 & ~n24657 ;
  assign n24659 = \s0_data_i[29]_pad  & n14647 ;
  assign n24660 = \s9_data_i[29]_pad  & n14666 ;
  assign n24661 = ~n24659 & ~n24660 ;
  assign n24662 = n24658 & n24661 ;
  assign n24663 = n24655 & n24662 ;
  assign n24664 = n24650 & n24663 ;
  assign n24665 = ~n24635 & n24664 ;
  assign n24666 = n2170 & n15936 ;
  assign n24667 = \s15_data_i[2]_pad  & n2170 ;
  assign n24668 = ~n2258 & n24667 ;
  assign n24669 = ~n24666 & ~n24668 ;
  assign n24670 = \s8_data_i[2]_pad  & n15086 ;
  assign n24671 = \s1_data_i[2]_pad  & n14653 ;
  assign n24672 = ~n24670 & ~n24671 ;
  assign n24673 = \s4_data_i[2]_pad  & n15074 ;
  assign n24674 = \s6_data_i[2]_pad  & n15078 ;
  assign n24675 = ~n24673 & ~n24674 ;
  assign n24676 = n24672 & n24675 ;
  assign n24677 = \s5_data_i[2]_pad  & n14675 ;
  assign n24678 = \s9_data_i[2]_pad  & n14666 ;
  assign n24679 = ~n24677 & ~n24678 ;
  assign n24680 = \s10_data_i[2]_pad  & n15047 ;
  assign n24681 = \s7_data_i[2]_pad  & n14671 ;
  assign n24682 = ~n24680 & ~n24681 ;
  assign n24683 = n24679 & n24682 ;
  assign n24684 = n24676 & n24683 ;
  assign n24685 = \s11_data_i[2]_pad  & n15051 ;
  assign n24686 = \s13_data_i[2]_pad  & n15055 ;
  assign n24687 = \s3_data_i[2]_pad  & n15070 ;
  assign n24688 = ~n24686 & ~n24687 ;
  assign n24689 = ~n24685 & n24688 ;
  assign n24690 = \s12_data_i[2]_pad  & n14685 ;
  assign n24691 = \s14_data_i[2]_pad  & n15059 ;
  assign n24692 = ~n24690 & ~n24691 ;
  assign n24693 = \s2_data_i[2]_pad  & n15066 ;
  assign n24694 = \s0_data_i[2]_pad  & n14647 ;
  assign n24695 = ~n24693 & ~n24694 ;
  assign n24696 = n24692 & n24695 ;
  assign n24697 = n24689 & n24696 ;
  assign n24698 = n24684 & n24697 ;
  assign n24699 = n24669 & n24698 ;
  assign n24700 = \s15_data_i[30]_pad  & n2170 ;
  assign n24701 = ~n2258 & n24700 ;
  assign n24702 = \s12_data_i[30]_pad  & n14685 ;
  assign n24703 = \s13_data_i[30]_pad  & n15055 ;
  assign n24704 = ~n24702 & ~n24703 ;
  assign n24705 = \s10_data_i[30]_pad  & n15047 ;
  assign n24706 = \s1_data_i[30]_pad  & n14653 ;
  assign n24707 = ~n24705 & ~n24706 ;
  assign n24708 = n24704 & n24707 ;
  assign n24709 = \s5_data_i[30]_pad  & n14675 ;
  assign n24710 = \s6_data_i[30]_pad  & n15078 ;
  assign n24711 = ~n24709 & ~n24710 ;
  assign n24712 = \s7_data_i[30]_pad  & n14671 ;
  assign n24713 = \s2_data_i[30]_pad  & n15066 ;
  assign n24714 = ~n24712 & ~n24713 ;
  assign n24715 = n24711 & n24714 ;
  assign n24716 = n24708 & n24715 ;
  assign n24717 = \s14_data_i[30]_pad  & n15059 ;
  assign n24718 = \s4_data_i[30]_pad  & n15074 ;
  assign n24719 = \s3_data_i[30]_pad  & n15070 ;
  assign n24720 = ~n24718 & ~n24719 ;
  assign n24721 = ~n24717 & n24720 ;
  assign n24722 = \s8_data_i[30]_pad  & n15086 ;
  assign n24723 = \s11_data_i[30]_pad  & n15051 ;
  assign n24724 = ~n24722 & ~n24723 ;
  assign n24725 = \s0_data_i[30]_pad  & n14647 ;
  assign n24726 = \s9_data_i[30]_pad  & n14666 ;
  assign n24727 = ~n24725 & ~n24726 ;
  assign n24728 = n24724 & n24727 ;
  assign n24729 = n24721 & n24728 ;
  assign n24730 = n24716 & n24729 ;
  assign n24731 = ~n24701 & n24730 ;
  assign n24732 = \s15_data_i[31]_pad  & n2170 ;
  assign n24733 = ~n2258 & n24732 ;
  assign n24734 = \s12_data_i[31]_pad  & n14685 ;
  assign n24735 = \s13_data_i[31]_pad  & n15055 ;
  assign n24736 = ~n24734 & ~n24735 ;
  assign n24737 = \s10_data_i[31]_pad  & n15047 ;
  assign n24738 = \s1_data_i[31]_pad  & n14653 ;
  assign n24739 = ~n24737 & ~n24738 ;
  assign n24740 = n24736 & n24739 ;
  assign n24741 = \s5_data_i[31]_pad  & n14675 ;
  assign n24742 = \s6_data_i[31]_pad  & n15078 ;
  assign n24743 = ~n24741 & ~n24742 ;
  assign n24744 = \s7_data_i[31]_pad  & n14671 ;
  assign n24745 = \s2_data_i[31]_pad  & n15066 ;
  assign n24746 = ~n24744 & ~n24745 ;
  assign n24747 = n24743 & n24746 ;
  assign n24748 = n24740 & n24747 ;
  assign n24749 = \s14_data_i[31]_pad  & n15059 ;
  assign n24750 = \s4_data_i[31]_pad  & n15074 ;
  assign n24751 = \s3_data_i[31]_pad  & n15070 ;
  assign n24752 = ~n24750 & ~n24751 ;
  assign n24753 = ~n24749 & n24752 ;
  assign n24754 = \s8_data_i[31]_pad  & n15086 ;
  assign n24755 = \s11_data_i[31]_pad  & n15051 ;
  assign n24756 = ~n24754 & ~n24755 ;
  assign n24757 = \s0_data_i[31]_pad  & n14647 ;
  assign n24758 = \s9_data_i[31]_pad  & n14666 ;
  assign n24759 = ~n24757 & ~n24758 ;
  assign n24760 = n24756 & n24759 ;
  assign n24761 = n24753 & n24760 ;
  assign n24762 = n24748 & n24761 ;
  assign n24763 = ~n24733 & n24762 ;
  assign n24764 = n2170 & n16037 ;
  assign n24765 = \s15_data_i[3]_pad  & n2170 ;
  assign n24766 = ~n2258 & n24765 ;
  assign n24767 = ~n24764 & ~n24766 ;
  assign n24768 = \s8_data_i[3]_pad  & n15086 ;
  assign n24769 = \s7_data_i[3]_pad  & n14671 ;
  assign n24770 = ~n24768 & ~n24769 ;
  assign n24771 = \s10_data_i[3]_pad  & n15047 ;
  assign n24772 = \s1_data_i[3]_pad  & n14653 ;
  assign n24773 = ~n24771 & ~n24772 ;
  assign n24774 = n24770 & n24773 ;
  assign n24775 = \s5_data_i[3]_pad  & n14675 ;
  assign n24776 = \s9_data_i[3]_pad  & n14666 ;
  assign n24777 = ~n24775 & ~n24776 ;
  assign n24778 = \s13_data_i[3]_pad  & n15055 ;
  assign n24779 = \s2_data_i[3]_pad  & n15066 ;
  assign n24780 = ~n24778 & ~n24779 ;
  assign n24781 = n24777 & n24780 ;
  assign n24782 = n24774 & n24781 ;
  assign n24783 = \s11_data_i[3]_pad  & n15051 ;
  assign n24784 = \s4_data_i[3]_pad  & n15074 ;
  assign n24785 = \s3_data_i[3]_pad  & n15070 ;
  assign n24786 = ~n24784 & ~n24785 ;
  assign n24787 = ~n24783 & n24786 ;
  assign n24788 = \s12_data_i[3]_pad  & n14685 ;
  assign n24789 = \s14_data_i[3]_pad  & n15059 ;
  assign n24790 = ~n24788 & ~n24789 ;
  assign n24791 = \s6_data_i[3]_pad  & n15078 ;
  assign n24792 = \s0_data_i[3]_pad  & n14647 ;
  assign n24793 = ~n24791 & ~n24792 ;
  assign n24794 = n24790 & n24793 ;
  assign n24795 = n24787 & n24794 ;
  assign n24796 = n24782 & n24795 ;
  assign n24797 = n24767 & n24796 ;
  assign n24798 = n2170 & n16074 ;
  assign n24799 = \s15_data_i[4]_pad  & n2170 ;
  assign n24800 = ~n2258 & n24799 ;
  assign n24801 = ~n24798 & ~n24800 ;
  assign n24802 = \s8_data_i[4]_pad  & n15086 ;
  assign n24803 = \s1_data_i[4]_pad  & n14653 ;
  assign n24804 = ~n24802 & ~n24803 ;
  assign n24805 = \s4_data_i[4]_pad  & n15074 ;
  assign n24806 = \s6_data_i[4]_pad  & n15078 ;
  assign n24807 = ~n24805 & ~n24806 ;
  assign n24808 = n24804 & n24807 ;
  assign n24809 = \s5_data_i[4]_pad  & n14675 ;
  assign n24810 = \s9_data_i[4]_pad  & n14666 ;
  assign n24811 = ~n24809 & ~n24810 ;
  assign n24812 = \s10_data_i[4]_pad  & n15047 ;
  assign n24813 = \s7_data_i[4]_pad  & n14671 ;
  assign n24814 = ~n24812 & ~n24813 ;
  assign n24815 = n24811 & n24814 ;
  assign n24816 = n24808 & n24815 ;
  assign n24817 = \s11_data_i[4]_pad  & n15051 ;
  assign n24818 = \s13_data_i[4]_pad  & n15055 ;
  assign n24819 = \s3_data_i[4]_pad  & n15070 ;
  assign n24820 = ~n24818 & ~n24819 ;
  assign n24821 = ~n24817 & n24820 ;
  assign n24822 = \s12_data_i[4]_pad  & n14685 ;
  assign n24823 = \s14_data_i[4]_pad  & n15059 ;
  assign n24824 = ~n24822 & ~n24823 ;
  assign n24825 = \s2_data_i[4]_pad  & n15066 ;
  assign n24826 = \s0_data_i[4]_pad  & n14647 ;
  assign n24827 = ~n24825 & ~n24826 ;
  assign n24828 = n24824 & n24827 ;
  assign n24829 = n24821 & n24828 ;
  assign n24830 = n24816 & n24829 ;
  assign n24831 = n24801 & n24830 ;
  assign n24832 = n2170 & n16111 ;
  assign n24833 = \s15_data_i[5]_pad  & n2170 ;
  assign n24834 = ~n2258 & n24833 ;
  assign n24835 = ~n24832 & ~n24834 ;
  assign n24836 = \s2_data_i[5]_pad  & n15066 ;
  assign n24837 = \s13_data_i[5]_pad  & n15055 ;
  assign n24838 = ~n24836 & ~n24837 ;
  assign n24839 = \s4_data_i[5]_pad  & n15074 ;
  assign n24840 = \s12_data_i[5]_pad  & n14685 ;
  assign n24841 = ~n24839 & ~n24840 ;
  assign n24842 = n24838 & n24841 ;
  assign n24843 = \s3_data_i[5]_pad  & n15070 ;
  assign n24844 = \s14_data_i[5]_pad  & n15059 ;
  assign n24845 = ~n24843 & ~n24844 ;
  assign n24846 = \s11_data_i[5]_pad  & n15051 ;
  assign n24847 = \s8_data_i[5]_pad  & n15086 ;
  assign n24848 = ~n24846 & ~n24847 ;
  assign n24849 = n24845 & n24848 ;
  assign n24850 = n24842 & n24849 ;
  assign n24851 = \s1_data_i[5]_pad  & n14653 ;
  assign n24852 = \s7_data_i[5]_pad  & n14671 ;
  assign n24853 = \s5_data_i[5]_pad  & n14675 ;
  assign n24854 = ~n24852 & ~n24853 ;
  assign n24855 = ~n24851 & n24854 ;
  assign n24856 = \s9_data_i[5]_pad  & n14666 ;
  assign n24857 = \s10_data_i[5]_pad  & n15047 ;
  assign n24858 = ~n24856 & ~n24857 ;
  assign n24859 = \s6_data_i[5]_pad  & n15078 ;
  assign n24860 = \s0_data_i[5]_pad  & n14647 ;
  assign n24861 = ~n24859 & ~n24860 ;
  assign n24862 = n24858 & n24861 ;
  assign n24863 = n24855 & n24862 ;
  assign n24864 = n24850 & n24863 ;
  assign n24865 = n24835 & n24864 ;
  assign n24866 = n2170 & n16148 ;
  assign n24867 = \s15_data_i[6]_pad  & n2170 ;
  assign n24868 = ~n2258 & n24867 ;
  assign n24869 = ~n24866 & ~n24868 ;
  assign n24870 = \s8_data_i[6]_pad  & n15086 ;
  assign n24871 = \s1_data_i[6]_pad  & n14653 ;
  assign n24872 = ~n24870 & ~n24871 ;
  assign n24873 = \s4_data_i[6]_pad  & n15074 ;
  assign n24874 = \s6_data_i[6]_pad  & n15078 ;
  assign n24875 = ~n24873 & ~n24874 ;
  assign n24876 = n24872 & n24875 ;
  assign n24877 = \s5_data_i[6]_pad  & n14675 ;
  assign n24878 = \s9_data_i[6]_pad  & n14666 ;
  assign n24879 = ~n24877 & ~n24878 ;
  assign n24880 = \s10_data_i[6]_pad  & n15047 ;
  assign n24881 = \s7_data_i[6]_pad  & n14671 ;
  assign n24882 = ~n24880 & ~n24881 ;
  assign n24883 = n24879 & n24882 ;
  assign n24884 = n24876 & n24883 ;
  assign n24885 = \s11_data_i[6]_pad  & n15051 ;
  assign n24886 = \s13_data_i[6]_pad  & n15055 ;
  assign n24887 = \s3_data_i[6]_pad  & n15070 ;
  assign n24888 = ~n24886 & ~n24887 ;
  assign n24889 = ~n24885 & n24888 ;
  assign n24890 = \s12_data_i[6]_pad  & n14685 ;
  assign n24891 = \s14_data_i[6]_pad  & n15059 ;
  assign n24892 = ~n24890 & ~n24891 ;
  assign n24893 = \s2_data_i[6]_pad  & n15066 ;
  assign n24894 = \s0_data_i[6]_pad  & n14647 ;
  assign n24895 = ~n24893 & ~n24894 ;
  assign n24896 = n24892 & n24895 ;
  assign n24897 = n24889 & n24896 ;
  assign n24898 = n24884 & n24897 ;
  assign n24899 = n24869 & n24898 ;
  assign n24900 = n2170 & n16185 ;
  assign n24901 = \s15_data_i[7]_pad  & n2170 ;
  assign n24902 = ~n2258 & n24901 ;
  assign n24903 = ~n24900 & ~n24902 ;
  assign n24904 = \s8_data_i[7]_pad  & n15086 ;
  assign n24905 = \s1_data_i[7]_pad  & n14653 ;
  assign n24906 = ~n24904 & ~n24905 ;
  assign n24907 = \s4_data_i[7]_pad  & n15074 ;
  assign n24908 = \s6_data_i[7]_pad  & n15078 ;
  assign n24909 = ~n24907 & ~n24908 ;
  assign n24910 = n24906 & n24909 ;
  assign n24911 = \s5_data_i[7]_pad  & n14675 ;
  assign n24912 = \s9_data_i[7]_pad  & n14666 ;
  assign n24913 = ~n24911 & ~n24912 ;
  assign n24914 = \s10_data_i[7]_pad  & n15047 ;
  assign n24915 = \s7_data_i[7]_pad  & n14671 ;
  assign n24916 = ~n24914 & ~n24915 ;
  assign n24917 = n24913 & n24916 ;
  assign n24918 = n24910 & n24917 ;
  assign n24919 = \s11_data_i[7]_pad  & n15051 ;
  assign n24920 = \s13_data_i[7]_pad  & n15055 ;
  assign n24921 = \s3_data_i[7]_pad  & n15070 ;
  assign n24922 = ~n24920 & ~n24921 ;
  assign n24923 = ~n24919 & n24922 ;
  assign n24924 = \s12_data_i[7]_pad  & n14685 ;
  assign n24925 = \s14_data_i[7]_pad  & n15059 ;
  assign n24926 = ~n24924 & ~n24925 ;
  assign n24927 = \s2_data_i[7]_pad  & n15066 ;
  assign n24928 = \s0_data_i[7]_pad  & n14647 ;
  assign n24929 = ~n24927 & ~n24928 ;
  assign n24930 = n24926 & n24929 ;
  assign n24931 = n24923 & n24930 ;
  assign n24932 = n24918 & n24931 ;
  assign n24933 = n24903 & n24932 ;
  assign n24934 = n2170 & n16222 ;
  assign n24935 = \s15_data_i[8]_pad  & n2170 ;
  assign n24936 = ~n2258 & n24935 ;
  assign n24937 = ~n24934 & ~n24936 ;
  assign n24938 = \s8_data_i[8]_pad  & n15086 ;
  assign n24939 = \s1_data_i[8]_pad  & n14653 ;
  assign n24940 = ~n24938 & ~n24939 ;
  assign n24941 = \s4_data_i[8]_pad  & n15074 ;
  assign n24942 = \s6_data_i[8]_pad  & n15078 ;
  assign n24943 = ~n24941 & ~n24942 ;
  assign n24944 = n24940 & n24943 ;
  assign n24945 = \s5_data_i[8]_pad  & n14675 ;
  assign n24946 = \s9_data_i[8]_pad  & n14666 ;
  assign n24947 = ~n24945 & ~n24946 ;
  assign n24948 = \s10_data_i[8]_pad  & n15047 ;
  assign n24949 = \s7_data_i[8]_pad  & n14671 ;
  assign n24950 = ~n24948 & ~n24949 ;
  assign n24951 = n24947 & n24950 ;
  assign n24952 = n24944 & n24951 ;
  assign n24953 = \s11_data_i[8]_pad  & n15051 ;
  assign n24954 = \s13_data_i[8]_pad  & n15055 ;
  assign n24955 = \s3_data_i[8]_pad  & n15070 ;
  assign n24956 = ~n24954 & ~n24955 ;
  assign n24957 = ~n24953 & n24956 ;
  assign n24958 = \s12_data_i[8]_pad  & n14685 ;
  assign n24959 = \s14_data_i[8]_pad  & n15059 ;
  assign n24960 = ~n24958 & ~n24959 ;
  assign n24961 = \s2_data_i[8]_pad  & n15066 ;
  assign n24962 = \s0_data_i[8]_pad  & n14647 ;
  assign n24963 = ~n24961 & ~n24962 ;
  assign n24964 = n24960 & n24963 ;
  assign n24965 = n24957 & n24964 ;
  assign n24966 = n24952 & n24965 ;
  assign n24967 = n24937 & n24966 ;
  assign n24968 = n2170 & n16259 ;
  assign n24969 = \s15_data_i[9]_pad  & n2170 ;
  assign n24970 = ~n2258 & n24969 ;
  assign n24971 = ~n24968 & ~n24970 ;
  assign n24972 = \s8_data_i[9]_pad  & n15086 ;
  assign n24973 = \s1_data_i[9]_pad  & n14653 ;
  assign n24974 = ~n24972 & ~n24973 ;
  assign n24975 = \s4_data_i[9]_pad  & n15074 ;
  assign n24976 = \s6_data_i[9]_pad  & n15078 ;
  assign n24977 = ~n24975 & ~n24976 ;
  assign n24978 = n24974 & n24977 ;
  assign n24979 = \s5_data_i[9]_pad  & n14675 ;
  assign n24980 = \s9_data_i[9]_pad  & n14666 ;
  assign n24981 = ~n24979 & ~n24980 ;
  assign n24982 = \s10_data_i[9]_pad  & n15047 ;
  assign n24983 = \s7_data_i[9]_pad  & n14671 ;
  assign n24984 = ~n24982 & ~n24983 ;
  assign n24985 = n24981 & n24984 ;
  assign n24986 = n24978 & n24985 ;
  assign n24987 = \s11_data_i[9]_pad  & n15051 ;
  assign n24988 = \s13_data_i[9]_pad  & n15055 ;
  assign n24989 = \s3_data_i[9]_pad  & n15070 ;
  assign n24990 = ~n24988 & ~n24989 ;
  assign n24991 = ~n24987 & n24990 ;
  assign n24992 = \s12_data_i[9]_pad  & n14685 ;
  assign n24993 = \s14_data_i[9]_pad  & n15059 ;
  assign n24994 = ~n24992 & ~n24993 ;
  assign n24995 = \s2_data_i[9]_pad  & n15066 ;
  assign n24996 = \s0_data_i[9]_pad  & n14647 ;
  assign n24997 = ~n24995 & ~n24996 ;
  assign n24998 = n24994 & n24997 ;
  assign n24999 = n24991 & n24998 ;
  assign n25000 = n24986 & n24999 ;
  assign n25001 = n24971 & n25000 ;
  assign n25002 = \s15_err_i_pad  & n23883 ;
  assign n25003 = ~n2258 & n25002 ;
  assign n25004 = \s11_err_i_pad  & n15051 ;
  assign n25005 = ~n14009 & n25004 ;
  assign n25006 = n14026 & n25005 ;
  assign n25007 = \s3_err_i_pad  & n15070 ;
  assign n25008 = ~n14451 & n25007 ;
  assign n25009 = n14468 & n25008 ;
  assign n25010 = ~n25006 & ~n25009 ;
  assign n25011 = \s13_err_i_pad  & n15055 ;
  assign n25012 = ~n14211 & n25011 ;
  assign n25013 = n14204 & n25012 ;
  assign n25014 = \s9_err_i_pad  & n14666 ;
  assign n25015 = ~n13847 & n25014 ;
  assign n25016 = n13864 & n25015 ;
  assign n25017 = ~n25013 & ~n25016 ;
  assign n25018 = n25010 & n25017 ;
  assign n25019 = \s6_err_i_pad  & n15078 ;
  assign n25020 = ~n13627 & n25019 ;
  assign n25021 = n13644 & n25020 ;
  assign n25022 = \s0_err_i_pad  & n14647 ;
  assign n25023 = ~n14069 & n25022 ;
  assign n25024 = n14062 & n25023 ;
  assign n25025 = ~n25021 & ~n25024 ;
  assign n25026 = \s4_err_i_pad  & n15074 ;
  assign n25027 = ~n13467 & n25026 ;
  assign n25028 = n13492 & n25027 ;
  assign n25029 = \s10_err_i_pad  & n15047 ;
  assign n25030 = ~n13928 & n25029 ;
  assign n25031 = n13936 & n25030 ;
  assign n25032 = ~n25028 & ~n25031 ;
  assign n25033 = n25025 & n25032 ;
  assign n25034 = n25018 & n25033 ;
  assign n25035 = \s8_err_i_pad  & n15086 ;
  assign n25036 = ~n13767 & n25035 ;
  assign n25037 = n13784 & n25036 ;
  assign n25038 = \s2_err_i_pad  & n15066 ;
  assign n25039 = ~n14391 & n25038 ;
  assign n25040 = n14408 & n25039 ;
  assign n25041 = \s7_err_i_pad  & n14671 ;
  assign n25042 = ~n13697 & n25041 ;
  assign n25043 = n13690 & n25042 ;
  assign n25044 = ~n25040 & ~n25043 ;
  assign n25045 = ~n25037 & n25044 ;
  assign n25046 = \s12_err_i_pad  & n14685 ;
  assign n25047 = ~n14140 & n25046 ;
  assign n25048 = n14148 & n25047 ;
  assign n25049 = \s14_err_i_pad  & n15059 ;
  assign n25050 = ~n14331 & n25049 ;
  assign n25051 = n14348 & n25050 ;
  assign n25052 = ~n25048 & ~n25051 ;
  assign n25053 = \s5_err_i_pad  & n14675 ;
  assign n25054 = ~n13547 & n25053 ;
  assign n25055 = n13564 & n25054 ;
  assign n25056 = \s1_err_i_pad  & n14653 ;
  assign n25057 = ~n14271 & n25056 ;
  assign n25058 = n14264 & n25057 ;
  assign n25059 = ~n25055 & ~n25058 ;
  assign n25060 = n25052 & n25059 ;
  assign n25061 = n25045 & n25060 ;
  assign n25062 = n25034 & n25061 ;
  assign n25063 = ~n25003 & n25062 ;
  assign n25064 = \s15_rty_i_pad  & n23883 ;
  assign n25065 = ~n2258 & n25064 ;
  assign n25066 = \s2_rty_i_pad  & n15066 ;
  assign n25067 = ~n14391 & n25066 ;
  assign n25068 = n14408 & n25067 ;
  assign n25069 = \s3_rty_i_pad  & n15070 ;
  assign n25070 = ~n14451 & n25069 ;
  assign n25071 = n14468 & n25070 ;
  assign n25072 = ~n25068 & ~n25071 ;
  assign n25073 = \s13_rty_i_pad  & n15055 ;
  assign n25074 = ~n14211 & n25073 ;
  assign n25075 = n14204 & n25074 ;
  assign n25076 = \s9_rty_i_pad  & n14666 ;
  assign n25077 = ~n13847 & n25076 ;
  assign n25078 = n13864 & n25077 ;
  assign n25079 = ~n25075 & ~n25078 ;
  assign n25080 = n25072 & n25079 ;
  assign n25081 = \s0_rty_i_pad  & n14647 ;
  assign n25082 = ~n14069 & n25081 ;
  assign n25083 = n14062 & n25082 ;
  assign n25084 = \s7_rty_i_pad  & n14671 ;
  assign n25085 = ~n13697 & n25084 ;
  assign n25086 = n13690 & n25085 ;
  assign n25087 = ~n25083 & ~n25086 ;
  assign n25088 = \s6_rty_i_pad  & n15078 ;
  assign n25089 = ~n13627 & n25088 ;
  assign n25090 = n13644 & n25089 ;
  assign n25091 = \s10_rty_i_pad  & n15047 ;
  assign n25092 = ~n13928 & n25091 ;
  assign n25093 = n13936 & n25092 ;
  assign n25094 = ~n25090 & ~n25093 ;
  assign n25095 = n25087 & n25094 ;
  assign n25096 = n25080 & n25095 ;
  assign n25097 = \s1_rty_i_pad  & n14653 ;
  assign n25098 = ~n14271 & n25097 ;
  assign n25099 = n14264 & n25098 ;
  assign n25100 = \s11_rty_i_pad  & n15051 ;
  assign n25101 = ~n14009 & n25100 ;
  assign n25102 = n14026 & n25101 ;
  assign n25103 = \s4_rty_i_pad  & n15074 ;
  assign n25104 = ~n13467 & n25103 ;
  assign n25105 = n13492 & n25104 ;
  assign n25106 = ~n25102 & ~n25105 ;
  assign n25107 = ~n25099 & n25106 ;
  assign n25108 = \s12_rty_i_pad  & n14685 ;
  assign n25109 = ~n14140 & n25108 ;
  assign n25110 = n14148 & n25109 ;
  assign n25111 = \s14_rty_i_pad  & n15059 ;
  assign n25112 = ~n14331 & n25111 ;
  assign n25113 = n14348 & n25112 ;
  assign n25114 = ~n25110 & ~n25113 ;
  assign n25115 = \s5_rty_i_pad  & n14675 ;
  assign n25116 = ~n13547 & n25115 ;
  assign n25117 = n13564 & n25116 ;
  assign n25118 = \s8_rty_i_pad  & n15086 ;
  assign n25119 = ~n13767 & n25118 ;
  assign n25120 = n13784 & n25119 ;
  assign n25121 = ~n25117 & ~n25120 ;
  assign n25122 = n25114 & n25121 ;
  assign n25123 = n25107 & n25122 ;
  assign n25124 = n25096 & n25123 ;
  assign n25125 = ~n25065 & n25124 ;
  assign n25126 = \m2_addr_i[0]_pad  & n14069 ;
  assign n25127 = n14086 & n25126 ;
  assign n25128 = \m3_addr_i[0]_pad  & ~n14069 ;
  assign n25129 = n14086 & n25128 ;
  assign n25130 = ~n25127 & ~n25129 ;
  assign n25131 = \m0_addr_i[0]_pad  & n14069 ;
  assign n25132 = n14094 & n25131 ;
  assign n25133 = \m7_addr_i[0]_pad  & ~n14069 ;
  assign n25134 = n14062 & n25133 ;
  assign n25135 = ~n25132 & ~n25134 ;
  assign n25136 = n25130 & n25135 ;
  assign n25137 = \m1_addr_i[0]_pad  & ~n14069 ;
  assign n25138 = n14094 & n25137 ;
  assign n25139 = \m6_addr_i[0]_pad  & n14069 ;
  assign n25140 = n14062 & n25139 ;
  assign n25141 = ~n25138 & ~n25140 ;
  assign n25142 = \m4_addr_i[0]_pad  & n14069 ;
  assign n25143 = n14077 & n25142 ;
  assign n25144 = \m5_addr_i[0]_pad  & ~n14069 ;
  assign n25145 = n14077 & n25144 ;
  assign n25146 = ~n25143 & ~n25145 ;
  assign n25147 = n25141 & n25146 ;
  assign n25148 = n25136 & n25147 ;
  assign n25149 = \m2_addr_i[10]_pad  & n14069 ;
  assign n25150 = n14086 & n25149 ;
  assign n25151 = \m3_addr_i[10]_pad  & ~n14069 ;
  assign n25152 = n14086 & n25151 ;
  assign n25153 = ~n25150 & ~n25152 ;
  assign n25154 = \m0_addr_i[10]_pad  & n14069 ;
  assign n25155 = n14094 & n25154 ;
  assign n25156 = \m5_addr_i[10]_pad  & ~n14069 ;
  assign n25157 = n14077 & n25156 ;
  assign n25158 = ~n25155 & ~n25157 ;
  assign n25159 = n25153 & n25158 ;
  assign n25160 = \m1_addr_i[10]_pad  & ~n14069 ;
  assign n25161 = n14094 & n25160 ;
  assign n25162 = \m4_addr_i[10]_pad  & n14069 ;
  assign n25163 = n14077 & n25162 ;
  assign n25164 = ~n25161 & ~n25163 ;
  assign n25165 = \m6_addr_i[10]_pad  & n14069 ;
  assign n25166 = n14062 & n25165 ;
  assign n25167 = \m7_addr_i[10]_pad  & ~n14069 ;
  assign n25168 = n14062 & n25167 ;
  assign n25169 = ~n25166 & ~n25168 ;
  assign n25170 = n25164 & n25169 ;
  assign n25171 = n25159 & n25170 ;
  assign n25172 = \m2_addr_i[11]_pad  & n14069 ;
  assign n25173 = n14086 & n25172 ;
  assign n25174 = \m3_addr_i[11]_pad  & ~n14069 ;
  assign n25175 = n14086 & n25174 ;
  assign n25176 = ~n25173 & ~n25175 ;
  assign n25177 = \m6_addr_i[11]_pad  & n14069 ;
  assign n25178 = n14062 & n25177 ;
  assign n25179 = \m1_addr_i[11]_pad  & ~n14069 ;
  assign n25180 = n14094 & n25179 ;
  assign n25181 = ~n25178 & ~n25180 ;
  assign n25182 = n25176 & n25181 ;
  assign n25183 = \m7_addr_i[11]_pad  & ~n14069 ;
  assign n25184 = n14062 & n25183 ;
  assign n25185 = \m0_addr_i[11]_pad  & n14069 ;
  assign n25186 = n14094 & n25185 ;
  assign n25187 = ~n25184 & ~n25186 ;
  assign n25188 = \m4_addr_i[11]_pad  & n14069 ;
  assign n25189 = n14077 & n25188 ;
  assign n25190 = \m5_addr_i[11]_pad  & ~n14069 ;
  assign n25191 = n14077 & n25190 ;
  assign n25192 = ~n25189 & ~n25191 ;
  assign n25193 = n25187 & n25192 ;
  assign n25194 = n25182 & n25193 ;
  assign n25195 = \m6_addr_i[12]_pad  & n14069 ;
  assign n25196 = n14062 & n25195 ;
  assign n25197 = \m7_addr_i[12]_pad  & ~n14069 ;
  assign n25198 = n14062 & n25197 ;
  assign n25199 = ~n25196 & ~n25198 ;
  assign n25200 = \m4_addr_i[12]_pad  & n14069 ;
  assign n25201 = n14077 & n25200 ;
  assign n25202 = \m3_addr_i[12]_pad  & ~n14069 ;
  assign n25203 = n14086 & n25202 ;
  assign n25204 = ~n25201 & ~n25203 ;
  assign n25205 = n25199 & n25204 ;
  assign n25206 = \m5_addr_i[12]_pad  & ~n14069 ;
  assign n25207 = n14077 & n25206 ;
  assign n25208 = \m2_addr_i[12]_pad  & n14069 ;
  assign n25209 = n14086 & n25208 ;
  assign n25210 = ~n25207 & ~n25209 ;
  assign n25211 = \m0_addr_i[12]_pad  & n14069 ;
  assign n25212 = n14094 & n25211 ;
  assign n25213 = \m1_addr_i[12]_pad  & ~n14069 ;
  assign n25214 = n14094 & n25213 ;
  assign n25215 = ~n25212 & ~n25214 ;
  assign n25216 = n25210 & n25215 ;
  assign n25217 = n25205 & n25216 ;
  assign n25218 = \m6_addr_i[13]_pad  & n14069 ;
  assign n25219 = n14062 & n25218 ;
  assign n25220 = \m7_addr_i[13]_pad  & ~n14069 ;
  assign n25221 = n14062 & n25220 ;
  assign n25222 = ~n25219 & ~n25221 ;
  assign n25223 = \m4_addr_i[13]_pad  & n14069 ;
  assign n25224 = n14077 & n25223 ;
  assign n25225 = \m1_addr_i[13]_pad  & ~n14069 ;
  assign n25226 = n14094 & n25225 ;
  assign n25227 = ~n25224 & ~n25226 ;
  assign n25228 = n25222 & n25227 ;
  assign n25229 = \m5_addr_i[13]_pad  & ~n14069 ;
  assign n25230 = n14077 & n25229 ;
  assign n25231 = \m0_addr_i[13]_pad  & n14069 ;
  assign n25232 = n14094 & n25231 ;
  assign n25233 = ~n25230 & ~n25232 ;
  assign n25234 = \m2_addr_i[13]_pad  & n14069 ;
  assign n25235 = n14086 & n25234 ;
  assign n25236 = \m3_addr_i[13]_pad  & ~n14069 ;
  assign n25237 = n14086 & n25236 ;
  assign n25238 = ~n25235 & ~n25237 ;
  assign n25239 = n25233 & n25238 ;
  assign n25240 = n25228 & n25239 ;
  assign n25241 = \m4_addr_i[14]_pad  & n14069 ;
  assign n25242 = n14077 & n25241 ;
  assign n25243 = \m5_addr_i[14]_pad  & ~n14069 ;
  assign n25244 = n14077 & n25243 ;
  assign n25245 = ~n25242 & ~n25244 ;
  assign n25246 = \m6_addr_i[14]_pad  & n14069 ;
  assign n25247 = n14062 & n25246 ;
  assign n25248 = \m1_addr_i[14]_pad  & ~n14069 ;
  assign n25249 = n14094 & n25248 ;
  assign n25250 = ~n25247 & ~n25249 ;
  assign n25251 = n25245 & n25250 ;
  assign n25252 = \m7_addr_i[14]_pad  & ~n14069 ;
  assign n25253 = n14062 & n25252 ;
  assign n25254 = \m0_addr_i[14]_pad  & n14069 ;
  assign n25255 = n14094 & n25254 ;
  assign n25256 = ~n25253 & ~n25255 ;
  assign n25257 = \m2_addr_i[14]_pad  & n14069 ;
  assign n25258 = n14086 & n25257 ;
  assign n25259 = \m3_addr_i[14]_pad  & ~n14069 ;
  assign n25260 = n14086 & n25259 ;
  assign n25261 = ~n25258 & ~n25260 ;
  assign n25262 = n25256 & n25261 ;
  assign n25263 = n25251 & n25262 ;
  assign n25264 = \m2_addr_i[15]_pad  & n14069 ;
  assign n25265 = n14086 & n25264 ;
  assign n25266 = \m3_addr_i[15]_pad  & ~n14069 ;
  assign n25267 = n14086 & n25266 ;
  assign n25268 = ~n25265 & ~n25267 ;
  assign n25269 = \m0_addr_i[15]_pad  & n14069 ;
  assign n25270 = n14094 & n25269 ;
  assign n25271 = \m7_addr_i[15]_pad  & ~n14069 ;
  assign n25272 = n14062 & n25271 ;
  assign n25273 = ~n25270 & ~n25272 ;
  assign n25274 = n25268 & n25273 ;
  assign n25275 = \m1_addr_i[15]_pad  & ~n14069 ;
  assign n25276 = n14094 & n25275 ;
  assign n25277 = \m6_addr_i[15]_pad  & n14069 ;
  assign n25278 = n14062 & n25277 ;
  assign n25279 = ~n25276 & ~n25278 ;
  assign n25280 = \m4_addr_i[15]_pad  & n14069 ;
  assign n25281 = n14077 & n25280 ;
  assign n25282 = \m5_addr_i[15]_pad  & ~n14069 ;
  assign n25283 = n14077 & n25282 ;
  assign n25284 = ~n25281 & ~n25283 ;
  assign n25285 = n25279 & n25284 ;
  assign n25286 = n25274 & n25285 ;
  assign n25287 = \m0_addr_i[16]_pad  & n14069 ;
  assign n25288 = n14094 & n25287 ;
  assign n25289 = \m1_addr_i[16]_pad  & ~n14069 ;
  assign n25290 = n14094 & n25289 ;
  assign n25291 = ~n25288 & ~n25290 ;
  assign n25292 = \m4_addr_i[16]_pad  & n14069 ;
  assign n25293 = n14077 & n25292 ;
  assign n25294 = \m3_addr_i[16]_pad  & ~n14069 ;
  assign n25295 = n14086 & n25294 ;
  assign n25296 = ~n25293 & ~n25295 ;
  assign n25297 = n25291 & n25296 ;
  assign n25298 = \m5_addr_i[16]_pad  & ~n14069 ;
  assign n25299 = n14077 & n25298 ;
  assign n25300 = \m2_addr_i[16]_pad  & n14069 ;
  assign n25301 = n14086 & n25300 ;
  assign n25302 = ~n25299 & ~n25301 ;
  assign n25303 = \m6_addr_i[16]_pad  & n14069 ;
  assign n25304 = n14062 & n25303 ;
  assign n25305 = \m7_addr_i[16]_pad  & ~n14069 ;
  assign n25306 = n14062 & n25305 ;
  assign n25307 = ~n25304 & ~n25306 ;
  assign n25308 = n25302 & n25307 ;
  assign n25309 = n25297 & n25308 ;
  assign n25310 = \m4_addr_i[17]_pad  & n14069 ;
  assign n25311 = n14077 & n25310 ;
  assign n25312 = \m5_addr_i[17]_pad  & ~n14069 ;
  assign n25313 = n14077 & n25312 ;
  assign n25314 = ~n25311 & ~n25313 ;
  assign n25315 = \m0_addr_i[17]_pad  & n14069 ;
  assign n25316 = n14094 & n25315 ;
  assign n25317 = \m3_addr_i[17]_pad  & ~n14069 ;
  assign n25318 = n14086 & n25317 ;
  assign n25319 = ~n25316 & ~n25318 ;
  assign n25320 = n25314 & n25319 ;
  assign n25321 = \m1_addr_i[17]_pad  & ~n14069 ;
  assign n25322 = n14094 & n25321 ;
  assign n25323 = \m2_addr_i[17]_pad  & n14069 ;
  assign n25324 = n14086 & n25323 ;
  assign n25325 = ~n25322 & ~n25324 ;
  assign n25326 = \m6_addr_i[17]_pad  & n14069 ;
  assign n25327 = n14062 & n25326 ;
  assign n25328 = \m7_addr_i[17]_pad  & ~n14069 ;
  assign n25329 = n14062 & n25328 ;
  assign n25330 = ~n25327 & ~n25329 ;
  assign n25331 = n25325 & n25330 ;
  assign n25332 = n25320 & n25331 ;
  assign n25333 = \m2_addr_i[18]_pad  & n14069 ;
  assign n25334 = n14086 & n25333 ;
  assign n25335 = \m3_addr_i[18]_pad  & ~n14069 ;
  assign n25336 = n14086 & n25335 ;
  assign n25337 = ~n25334 & ~n25336 ;
  assign n25338 = \m0_addr_i[18]_pad  & n14069 ;
  assign n25339 = n14094 & n25338 ;
  assign n25340 = \m5_addr_i[18]_pad  & ~n14069 ;
  assign n25341 = n14077 & n25340 ;
  assign n25342 = ~n25339 & ~n25341 ;
  assign n25343 = n25337 & n25342 ;
  assign n25344 = \m1_addr_i[18]_pad  & ~n14069 ;
  assign n25345 = n14094 & n25344 ;
  assign n25346 = \m4_addr_i[18]_pad  & n14069 ;
  assign n25347 = n14077 & n25346 ;
  assign n25348 = ~n25345 & ~n25347 ;
  assign n25349 = \m6_addr_i[18]_pad  & n14069 ;
  assign n25350 = n14062 & n25349 ;
  assign n25351 = \m7_addr_i[18]_pad  & ~n14069 ;
  assign n25352 = n14062 & n25351 ;
  assign n25353 = ~n25350 & ~n25352 ;
  assign n25354 = n25348 & n25353 ;
  assign n25355 = n25343 & n25354 ;
  assign n25356 = \m2_addr_i[19]_pad  & n14069 ;
  assign n25357 = n14086 & n25356 ;
  assign n25358 = \m3_addr_i[19]_pad  & ~n14069 ;
  assign n25359 = n14086 & n25358 ;
  assign n25360 = ~n25357 & ~n25359 ;
  assign n25361 = \m4_addr_i[19]_pad  & n14069 ;
  assign n25362 = n14077 & n25361 ;
  assign n25363 = \m1_addr_i[19]_pad  & ~n14069 ;
  assign n25364 = n14094 & n25363 ;
  assign n25365 = ~n25362 & ~n25364 ;
  assign n25366 = n25360 & n25365 ;
  assign n25367 = \m5_addr_i[19]_pad  & ~n14069 ;
  assign n25368 = n14077 & n25367 ;
  assign n25369 = \m0_addr_i[19]_pad  & n14069 ;
  assign n25370 = n14094 & n25369 ;
  assign n25371 = ~n25368 & ~n25370 ;
  assign n25372 = \m6_addr_i[19]_pad  & n14069 ;
  assign n25373 = n14062 & n25372 ;
  assign n25374 = \m7_addr_i[19]_pad  & ~n14069 ;
  assign n25375 = n14062 & n25374 ;
  assign n25376 = ~n25373 & ~n25375 ;
  assign n25377 = n25371 & n25376 ;
  assign n25378 = n25366 & n25377 ;
  assign n25379 = \m0_addr_i[1]_pad  & n14069 ;
  assign n25380 = n14094 & n25379 ;
  assign n25381 = \m1_addr_i[1]_pad  & ~n14069 ;
  assign n25382 = n14094 & n25381 ;
  assign n25383 = ~n25380 & ~n25382 ;
  assign n25384 = \m6_addr_i[1]_pad  & n14069 ;
  assign n25385 = n14062 & n25384 ;
  assign n25386 = \m3_addr_i[1]_pad  & ~n14069 ;
  assign n25387 = n14086 & n25386 ;
  assign n25388 = ~n25385 & ~n25387 ;
  assign n25389 = n25383 & n25388 ;
  assign n25390 = \m7_addr_i[1]_pad  & ~n14069 ;
  assign n25391 = n14062 & n25390 ;
  assign n25392 = \m2_addr_i[1]_pad  & n14069 ;
  assign n25393 = n14086 & n25392 ;
  assign n25394 = ~n25391 & ~n25393 ;
  assign n25395 = \m4_addr_i[1]_pad  & n14069 ;
  assign n25396 = n14077 & n25395 ;
  assign n25397 = \m5_addr_i[1]_pad  & ~n14069 ;
  assign n25398 = n14077 & n25397 ;
  assign n25399 = ~n25396 & ~n25398 ;
  assign n25400 = n25394 & n25399 ;
  assign n25401 = n25389 & n25400 ;
  assign n25402 = \m6_addr_i[20]_pad  & n14069 ;
  assign n25403 = n14062 & n25402 ;
  assign n25404 = \m7_addr_i[20]_pad  & ~n14069 ;
  assign n25405 = n14062 & n25404 ;
  assign n25406 = ~n25403 & ~n25405 ;
  assign n25407 = \m4_addr_i[20]_pad  & n14069 ;
  assign n25408 = n14077 & n25407 ;
  assign n25409 = \m1_addr_i[20]_pad  & ~n14069 ;
  assign n25410 = n14094 & n25409 ;
  assign n25411 = ~n25408 & ~n25410 ;
  assign n25412 = n25406 & n25411 ;
  assign n25413 = \m5_addr_i[20]_pad  & ~n14069 ;
  assign n25414 = n14077 & n25413 ;
  assign n25415 = \m0_addr_i[20]_pad  & n14069 ;
  assign n25416 = n14094 & n25415 ;
  assign n25417 = ~n25414 & ~n25416 ;
  assign n25418 = \m2_addr_i[20]_pad  & n14069 ;
  assign n25419 = n14086 & n25418 ;
  assign n25420 = \m3_addr_i[20]_pad  & ~n14069 ;
  assign n25421 = n14086 & n25420 ;
  assign n25422 = ~n25419 & ~n25421 ;
  assign n25423 = n25417 & n25422 ;
  assign n25424 = n25412 & n25423 ;
  assign n25425 = \m6_addr_i[21]_pad  & n14069 ;
  assign n25426 = n14062 & n25425 ;
  assign n25427 = \m7_addr_i[21]_pad  & ~n14069 ;
  assign n25428 = n14062 & n25427 ;
  assign n25429 = ~n25426 & ~n25428 ;
  assign n25430 = \m0_addr_i[21]_pad  & n14069 ;
  assign n25431 = n14094 & n25430 ;
  assign n25432 = \m3_addr_i[21]_pad  & ~n14069 ;
  assign n25433 = n14086 & n25432 ;
  assign n25434 = ~n25431 & ~n25433 ;
  assign n25435 = n25429 & n25434 ;
  assign n25436 = \m1_addr_i[21]_pad  & ~n14069 ;
  assign n25437 = n14094 & n25436 ;
  assign n25438 = \m2_addr_i[21]_pad  & n14069 ;
  assign n25439 = n14086 & n25438 ;
  assign n25440 = ~n25437 & ~n25439 ;
  assign n25441 = \m4_addr_i[21]_pad  & n14069 ;
  assign n25442 = n14077 & n25441 ;
  assign n25443 = \m5_addr_i[21]_pad  & ~n14069 ;
  assign n25444 = n14077 & n25443 ;
  assign n25445 = ~n25442 & ~n25444 ;
  assign n25446 = n25440 & n25445 ;
  assign n25447 = n25435 & n25446 ;
  assign n25448 = \m6_addr_i[22]_pad  & n14069 ;
  assign n25449 = n14062 & n25448 ;
  assign n25450 = \m7_addr_i[22]_pad  & ~n14069 ;
  assign n25451 = n14062 & n25450 ;
  assign n25452 = ~n25449 & ~n25451 ;
  assign n25453 = \m2_addr_i[22]_pad  & n14069 ;
  assign n25454 = n14086 & n25453 ;
  assign n25455 = \m1_addr_i[22]_pad  & ~n14069 ;
  assign n25456 = n14094 & n25455 ;
  assign n25457 = ~n25454 & ~n25456 ;
  assign n25458 = n25452 & n25457 ;
  assign n25459 = \m3_addr_i[22]_pad  & ~n14069 ;
  assign n25460 = n14086 & n25459 ;
  assign n25461 = \m0_addr_i[22]_pad  & n14069 ;
  assign n25462 = n14094 & n25461 ;
  assign n25463 = ~n25460 & ~n25462 ;
  assign n25464 = \m4_addr_i[22]_pad  & n14069 ;
  assign n25465 = n14077 & n25464 ;
  assign n25466 = \m5_addr_i[22]_pad  & ~n14069 ;
  assign n25467 = n14077 & n25466 ;
  assign n25468 = ~n25465 & ~n25467 ;
  assign n25469 = n25463 & n25468 ;
  assign n25470 = n25458 & n25469 ;
  assign n25471 = \m4_addr_i[23]_pad  & n14069 ;
  assign n25472 = n14077 & n25471 ;
  assign n25473 = \m5_addr_i[23]_pad  & ~n14069 ;
  assign n25474 = n14077 & n25473 ;
  assign n25475 = ~n25472 & ~n25474 ;
  assign n25476 = \m0_addr_i[23]_pad  & n14069 ;
  assign n25477 = n14094 & n25476 ;
  assign n25478 = \m7_addr_i[23]_pad  & ~n14069 ;
  assign n25479 = n14062 & n25478 ;
  assign n25480 = ~n25477 & ~n25479 ;
  assign n25481 = n25475 & n25480 ;
  assign n25482 = \m1_addr_i[23]_pad  & ~n14069 ;
  assign n25483 = n14094 & n25482 ;
  assign n25484 = \m6_addr_i[23]_pad  & n14069 ;
  assign n25485 = n14062 & n25484 ;
  assign n25486 = ~n25483 & ~n25485 ;
  assign n25487 = \m2_addr_i[23]_pad  & n14069 ;
  assign n25488 = n14086 & n25487 ;
  assign n25489 = \m3_addr_i[23]_pad  & ~n14069 ;
  assign n25490 = n14086 & n25489 ;
  assign n25491 = ~n25488 & ~n25490 ;
  assign n25492 = n25486 & n25491 ;
  assign n25493 = n25481 & n25492 ;
  assign n25494 = \m0_addr_i[24]_pad  & n14069 ;
  assign n25495 = n14094 & n25494 ;
  assign n25496 = \m7_addr_i[24]_pad  & ~n14069 ;
  assign n25497 = n14062 & n25496 ;
  assign n25498 = ~n25495 & ~n25497 ;
  assign n25499 = \m1_addr_i[24]_pad  & ~n14069 ;
  assign n25500 = n14094 & n25499 ;
  assign n25501 = \m4_addr_i[24]_pad  & n14069 ;
  assign n25502 = n14077 & n25501 ;
  assign n25503 = ~n25500 & ~n25502 ;
  assign n25504 = n25498 & n25503 ;
  assign n25505 = \m2_addr_i[24]_pad  & n14069 ;
  assign n25506 = n14086 & n25505 ;
  assign n25507 = \m3_addr_i[24]_pad  & ~n14069 ;
  assign n25508 = n14086 & n25507 ;
  assign n25509 = ~n25506 & ~n25508 ;
  assign n25510 = \m5_addr_i[24]_pad  & ~n14069 ;
  assign n25511 = n14077 & n25510 ;
  assign n25512 = \m6_addr_i[24]_pad  & n14069 ;
  assign n25513 = n14062 & n25512 ;
  assign n25514 = ~n25511 & ~n25513 ;
  assign n25515 = n25509 & n25514 ;
  assign n25516 = n25504 & n25515 ;
  assign n25517 = \m0_addr_i[25]_pad  & n14069 ;
  assign n25518 = n14094 & n25517 ;
  assign n25519 = \m7_addr_i[25]_pad  & ~n14069 ;
  assign n25520 = n14062 & n25519 ;
  assign n25521 = ~n25518 & ~n25520 ;
  assign n25522 = \m1_addr_i[25]_pad  & ~n14069 ;
  assign n25523 = n14094 & n25522 ;
  assign n25524 = \m4_addr_i[25]_pad  & n14069 ;
  assign n25525 = n14077 & n25524 ;
  assign n25526 = ~n25523 & ~n25525 ;
  assign n25527 = n25521 & n25526 ;
  assign n25528 = \m2_addr_i[25]_pad  & n14069 ;
  assign n25529 = n14086 & n25528 ;
  assign n25530 = \m3_addr_i[25]_pad  & ~n14069 ;
  assign n25531 = n14086 & n25530 ;
  assign n25532 = ~n25529 & ~n25531 ;
  assign n25533 = \m5_addr_i[25]_pad  & ~n14069 ;
  assign n25534 = n14077 & n25533 ;
  assign n25535 = \m6_addr_i[25]_pad  & n14069 ;
  assign n25536 = n14062 & n25535 ;
  assign n25537 = ~n25534 & ~n25536 ;
  assign n25538 = n25532 & n25537 ;
  assign n25539 = n25527 & n25538 ;
  assign n25540 = \m1_addr_i[26]_pad  & ~n14069 ;
  assign n25541 = n14094 & n25540 ;
  assign n25542 = \m2_addr_i[26]_pad  & n14069 ;
  assign n25543 = n14086 & n25542 ;
  assign n25544 = ~n25541 & ~n25543 ;
  assign n25545 = \m0_addr_i[26]_pad  & n14069 ;
  assign n25546 = n14094 & n25545 ;
  assign n25547 = \m4_addr_i[26]_pad  & n14069 ;
  assign n25548 = n14077 & n25547 ;
  assign n25549 = ~n25546 & ~n25548 ;
  assign n25550 = n25544 & n25549 ;
  assign n25551 = \m7_addr_i[26]_pad  & ~n14069 ;
  assign n25552 = n14062 & n25551 ;
  assign n25553 = \m3_addr_i[26]_pad  & ~n14069 ;
  assign n25554 = n14086 & n25553 ;
  assign n25555 = ~n25552 & ~n25554 ;
  assign n25556 = \m5_addr_i[26]_pad  & ~n14069 ;
  assign n25557 = n14077 & n25556 ;
  assign n25558 = \m6_addr_i[26]_pad  & n14069 ;
  assign n25559 = n14062 & n25558 ;
  assign n25560 = ~n25557 & ~n25559 ;
  assign n25561 = n25555 & n25560 ;
  assign n25562 = n25550 & n25561 ;
  assign n25563 = \m1_addr_i[27]_pad  & ~n14069 ;
  assign n25564 = n14094 & n25563 ;
  assign n25565 = \m2_addr_i[27]_pad  & n14069 ;
  assign n25566 = n14086 & n25565 ;
  assign n25567 = ~n25564 & ~n25566 ;
  assign n25568 = \m0_addr_i[27]_pad  & n14069 ;
  assign n25569 = n14094 & n25568 ;
  assign n25570 = \m6_addr_i[27]_pad  & n14069 ;
  assign n25571 = n14062 & n25570 ;
  assign n25572 = ~n25569 & ~n25571 ;
  assign n25573 = n25567 & n25572 ;
  assign n25574 = \m7_addr_i[27]_pad  & ~n14069 ;
  assign n25575 = n14062 & n25574 ;
  assign n25576 = \m5_addr_i[27]_pad  & ~n14069 ;
  assign n25577 = n14077 & n25576 ;
  assign n25578 = ~n25575 & ~n25577 ;
  assign n25579 = \m3_addr_i[27]_pad  & ~n14069 ;
  assign n25580 = n14086 & n25579 ;
  assign n25581 = \m4_addr_i[27]_pad  & n14069 ;
  assign n25582 = n14077 & n25581 ;
  assign n25583 = ~n25580 & ~n25582 ;
  assign n25584 = n25578 & n25583 ;
  assign n25585 = n25573 & n25584 ;
  assign n25586 = \m1_addr_i[28]_pad  & ~n14069 ;
  assign n25587 = n14094 & n25586 ;
  assign n25588 = \m2_addr_i[28]_pad  & n14069 ;
  assign n25589 = n14086 & n25588 ;
  assign n25590 = ~n25587 & ~n25589 ;
  assign n25591 = \m5_addr_i[28]_pad  & ~n14069 ;
  assign n25592 = n14077 & n25591 ;
  assign n25593 = \m4_addr_i[28]_pad  & n14069 ;
  assign n25594 = n14077 & n25593 ;
  assign n25595 = ~n25592 & ~n25594 ;
  assign n25596 = n25590 & n25595 ;
  assign n25597 = \m6_addr_i[28]_pad  & n14069 ;
  assign n25598 = n14062 & n25597 ;
  assign n25599 = \m3_addr_i[28]_pad  & ~n14069 ;
  assign n25600 = n14086 & n25599 ;
  assign n25601 = ~n25598 & ~n25600 ;
  assign n25602 = \m0_addr_i[28]_pad  & n14069 ;
  assign n25603 = n14094 & n25602 ;
  assign n25604 = \m7_addr_i[28]_pad  & ~n14069 ;
  assign n25605 = n14062 & n25604 ;
  assign n25606 = ~n25603 & ~n25605 ;
  assign n25607 = n25601 & n25606 ;
  assign n25608 = n25596 & n25607 ;
  assign n25609 = \m3_addr_i[29]_pad  & ~n14069 ;
  assign n25610 = n14086 & n25609 ;
  assign n25611 = \m4_addr_i[29]_pad  & n14069 ;
  assign n25612 = n14077 & n25611 ;
  assign n25613 = ~n25610 & ~n25612 ;
  assign n25614 = \m1_addr_i[29]_pad  & ~n14069 ;
  assign n25615 = n14094 & n25614 ;
  assign n25616 = \m7_addr_i[29]_pad  & ~n14069 ;
  assign n25617 = n14062 & n25616 ;
  assign n25618 = ~n25615 & ~n25617 ;
  assign n25619 = n25613 & n25618 ;
  assign n25620 = \m2_addr_i[29]_pad  & n14069 ;
  assign n25621 = n14086 & n25620 ;
  assign n25622 = \m0_addr_i[29]_pad  & n14069 ;
  assign n25623 = n14094 & n25622 ;
  assign n25624 = ~n25621 & ~n25623 ;
  assign n25625 = \m5_addr_i[29]_pad  & ~n14069 ;
  assign n25626 = n14077 & n25625 ;
  assign n25627 = \m6_addr_i[29]_pad  & n14069 ;
  assign n25628 = n14062 & n25627 ;
  assign n25629 = ~n25626 & ~n25628 ;
  assign n25630 = n25624 & n25629 ;
  assign n25631 = n25619 & n25630 ;
  assign n25632 = \m2_addr_i[2]_pad  & n14069 ;
  assign n25633 = n14086 & n25632 ;
  assign n25634 = \m3_addr_i[2]_pad  & ~n14069 ;
  assign n25635 = n14086 & n25634 ;
  assign n25636 = ~n25633 & ~n25635 ;
  assign n25637 = \m0_addr_i[2]_pad  & n14069 ;
  assign n25638 = n14094 & n25637 ;
  assign n25639 = \m7_addr_i[2]_pad  & ~n14069 ;
  assign n25640 = n14062 & n25639 ;
  assign n25641 = ~n25638 & ~n25640 ;
  assign n25642 = n25636 & n25641 ;
  assign n25643 = \m1_addr_i[2]_pad  & ~n14069 ;
  assign n25644 = n14094 & n25643 ;
  assign n25645 = \m6_addr_i[2]_pad  & n14069 ;
  assign n25646 = n14062 & n25645 ;
  assign n25647 = ~n25644 & ~n25646 ;
  assign n25648 = \m4_addr_i[2]_pad  & n14069 ;
  assign n25649 = n14077 & n25648 ;
  assign n25650 = \m5_addr_i[2]_pad  & ~n14069 ;
  assign n25651 = n14077 & n25650 ;
  assign n25652 = ~n25649 & ~n25651 ;
  assign n25653 = n25647 & n25652 ;
  assign n25654 = n25642 & n25653 ;
  assign n25655 = \m3_addr_i[30]_pad  & ~n14069 ;
  assign n25656 = n14086 & n25655 ;
  assign n25657 = \m4_addr_i[30]_pad  & n14069 ;
  assign n25658 = n14077 & n25657 ;
  assign n25659 = ~n25656 & ~n25658 ;
  assign n25660 = \m0_addr_i[30]_pad  & n14069 ;
  assign n25661 = n14094 & n25660 ;
  assign n25662 = \m6_addr_i[30]_pad  & n14069 ;
  assign n25663 = n14062 & n25662 ;
  assign n25664 = ~n25661 & ~n25663 ;
  assign n25665 = n25659 & n25664 ;
  assign n25666 = \m7_addr_i[30]_pad  & ~n14069 ;
  assign n25667 = n14062 & n25666 ;
  assign n25668 = \m5_addr_i[30]_pad  & ~n14069 ;
  assign n25669 = n14077 & n25668 ;
  assign n25670 = ~n25667 & ~n25669 ;
  assign n25671 = \m1_addr_i[30]_pad  & ~n14069 ;
  assign n25672 = n14094 & n25671 ;
  assign n25673 = \m2_addr_i[30]_pad  & n14069 ;
  assign n25674 = n14086 & n25673 ;
  assign n25675 = ~n25672 & ~n25674 ;
  assign n25676 = n25670 & n25675 ;
  assign n25677 = n25665 & n25676 ;
  assign n25678 = \m1_addr_i[31]_pad  & ~n14069 ;
  assign n25679 = n14094 & n25678 ;
  assign n25680 = \m2_addr_i[31]_pad  & n14069 ;
  assign n25681 = n14086 & n25680 ;
  assign n25682 = ~n25679 & ~n25681 ;
  assign n25683 = \m0_addr_i[31]_pad  & n14069 ;
  assign n25684 = n14094 & n25683 ;
  assign n25685 = \m4_addr_i[31]_pad  & n14069 ;
  assign n25686 = n14077 & n25685 ;
  assign n25687 = ~n25684 & ~n25686 ;
  assign n25688 = n25682 & n25687 ;
  assign n25689 = \m7_addr_i[31]_pad  & ~n14069 ;
  assign n25690 = n14062 & n25689 ;
  assign n25691 = \m3_addr_i[31]_pad  & ~n14069 ;
  assign n25692 = n14086 & n25691 ;
  assign n25693 = ~n25690 & ~n25692 ;
  assign n25694 = \m5_addr_i[31]_pad  & ~n14069 ;
  assign n25695 = n14077 & n25694 ;
  assign n25696 = \m6_addr_i[31]_pad  & n14069 ;
  assign n25697 = n14062 & n25696 ;
  assign n25698 = ~n25695 & ~n25697 ;
  assign n25699 = n25693 & n25698 ;
  assign n25700 = n25688 & n25699 ;
  assign n25701 = \m2_addr_i[3]_pad  & n14069 ;
  assign n25702 = n14086 & n25701 ;
  assign n25703 = \m3_addr_i[3]_pad  & ~n14069 ;
  assign n25704 = n14086 & n25703 ;
  assign n25705 = ~n25702 & ~n25704 ;
  assign n25706 = \m0_addr_i[3]_pad  & n14069 ;
  assign n25707 = n14094 & n25706 ;
  assign n25708 = \m7_addr_i[3]_pad  & ~n14069 ;
  assign n25709 = n14062 & n25708 ;
  assign n25710 = ~n25707 & ~n25709 ;
  assign n25711 = n25705 & n25710 ;
  assign n25712 = \m1_addr_i[3]_pad  & ~n14069 ;
  assign n25713 = n14094 & n25712 ;
  assign n25714 = \m6_addr_i[3]_pad  & n14069 ;
  assign n25715 = n14062 & n25714 ;
  assign n25716 = ~n25713 & ~n25715 ;
  assign n25717 = \m4_addr_i[3]_pad  & n14069 ;
  assign n25718 = n14077 & n25717 ;
  assign n25719 = \m5_addr_i[3]_pad  & ~n14069 ;
  assign n25720 = n14077 & n25719 ;
  assign n25721 = ~n25718 & ~n25720 ;
  assign n25722 = n25716 & n25721 ;
  assign n25723 = n25711 & n25722 ;
  assign n25724 = \m2_addr_i[4]_pad  & n14069 ;
  assign n25725 = n14086 & n25724 ;
  assign n25726 = \m3_addr_i[4]_pad  & ~n14069 ;
  assign n25727 = n14086 & n25726 ;
  assign n25728 = ~n25725 & ~n25727 ;
  assign n25729 = \m0_addr_i[4]_pad  & n14069 ;
  assign n25730 = n14094 & n25729 ;
  assign n25731 = \m7_addr_i[4]_pad  & ~n14069 ;
  assign n25732 = n14062 & n25731 ;
  assign n25733 = ~n25730 & ~n25732 ;
  assign n25734 = n25728 & n25733 ;
  assign n25735 = \m1_addr_i[4]_pad  & ~n14069 ;
  assign n25736 = n14094 & n25735 ;
  assign n25737 = \m6_addr_i[4]_pad  & n14069 ;
  assign n25738 = n14062 & n25737 ;
  assign n25739 = ~n25736 & ~n25738 ;
  assign n25740 = \m4_addr_i[4]_pad  & n14069 ;
  assign n25741 = n14077 & n25740 ;
  assign n25742 = \m5_addr_i[4]_pad  & ~n14069 ;
  assign n25743 = n14077 & n25742 ;
  assign n25744 = ~n25741 & ~n25743 ;
  assign n25745 = n25739 & n25744 ;
  assign n25746 = n25734 & n25745 ;
  assign n25747 = \m2_addr_i[5]_pad  & n14069 ;
  assign n25748 = n14086 & n25747 ;
  assign n25749 = \m3_addr_i[5]_pad  & ~n14069 ;
  assign n25750 = n14086 & n25749 ;
  assign n25751 = ~n25748 & ~n25750 ;
  assign n25752 = \m0_addr_i[5]_pad  & n14069 ;
  assign n25753 = n14094 & n25752 ;
  assign n25754 = \m7_addr_i[5]_pad  & ~n14069 ;
  assign n25755 = n14062 & n25754 ;
  assign n25756 = ~n25753 & ~n25755 ;
  assign n25757 = n25751 & n25756 ;
  assign n25758 = \m1_addr_i[5]_pad  & ~n14069 ;
  assign n25759 = n14094 & n25758 ;
  assign n25760 = \m6_addr_i[5]_pad  & n14069 ;
  assign n25761 = n14062 & n25760 ;
  assign n25762 = ~n25759 & ~n25761 ;
  assign n25763 = \m4_addr_i[5]_pad  & n14069 ;
  assign n25764 = n14077 & n25763 ;
  assign n25765 = \m5_addr_i[5]_pad  & ~n14069 ;
  assign n25766 = n14077 & n25765 ;
  assign n25767 = ~n25764 & ~n25766 ;
  assign n25768 = n25762 & n25767 ;
  assign n25769 = n25757 & n25768 ;
  assign n25770 = \m2_addr_i[6]_pad  & n14069 ;
  assign n25771 = n14086 & n25770 ;
  assign n25772 = \m3_addr_i[6]_pad  & ~n14069 ;
  assign n25773 = n14086 & n25772 ;
  assign n25774 = ~n25771 & ~n25773 ;
  assign n25775 = \m0_addr_i[6]_pad  & n14069 ;
  assign n25776 = n14094 & n25775 ;
  assign n25777 = \m7_addr_i[6]_pad  & ~n14069 ;
  assign n25778 = n14062 & n25777 ;
  assign n25779 = ~n25776 & ~n25778 ;
  assign n25780 = n25774 & n25779 ;
  assign n25781 = \m1_addr_i[6]_pad  & ~n14069 ;
  assign n25782 = n14094 & n25781 ;
  assign n25783 = \m6_addr_i[6]_pad  & n14069 ;
  assign n25784 = n14062 & n25783 ;
  assign n25785 = ~n25782 & ~n25784 ;
  assign n25786 = \m4_addr_i[6]_pad  & n14069 ;
  assign n25787 = n14077 & n25786 ;
  assign n25788 = \m5_addr_i[6]_pad  & ~n14069 ;
  assign n25789 = n14077 & n25788 ;
  assign n25790 = ~n25787 & ~n25789 ;
  assign n25791 = n25785 & n25790 ;
  assign n25792 = n25780 & n25791 ;
  assign n25793 = \m2_addr_i[7]_pad  & n14069 ;
  assign n25794 = n14086 & n25793 ;
  assign n25795 = \m3_addr_i[7]_pad  & ~n14069 ;
  assign n25796 = n14086 & n25795 ;
  assign n25797 = ~n25794 & ~n25796 ;
  assign n25798 = \m0_addr_i[7]_pad  & n14069 ;
  assign n25799 = n14094 & n25798 ;
  assign n25800 = \m7_addr_i[7]_pad  & ~n14069 ;
  assign n25801 = n14062 & n25800 ;
  assign n25802 = ~n25799 & ~n25801 ;
  assign n25803 = n25797 & n25802 ;
  assign n25804 = \m1_addr_i[7]_pad  & ~n14069 ;
  assign n25805 = n14094 & n25804 ;
  assign n25806 = \m6_addr_i[7]_pad  & n14069 ;
  assign n25807 = n14062 & n25806 ;
  assign n25808 = ~n25805 & ~n25807 ;
  assign n25809 = \m4_addr_i[7]_pad  & n14069 ;
  assign n25810 = n14077 & n25809 ;
  assign n25811 = \m5_addr_i[7]_pad  & ~n14069 ;
  assign n25812 = n14077 & n25811 ;
  assign n25813 = ~n25810 & ~n25812 ;
  assign n25814 = n25808 & n25813 ;
  assign n25815 = n25803 & n25814 ;
  assign n25816 = \m0_addr_i[8]_pad  & n14069 ;
  assign n25817 = n14094 & n25816 ;
  assign n25818 = \m1_addr_i[8]_pad  & ~n14069 ;
  assign n25819 = n14094 & n25818 ;
  assign n25820 = ~n25817 & ~n25819 ;
  assign n25821 = \m6_addr_i[8]_pad  & n14069 ;
  assign n25822 = n14062 & n25821 ;
  assign n25823 = \m3_addr_i[8]_pad  & ~n14069 ;
  assign n25824 = n14086 & n25823 ;
  assign n25825 = ~n25822 & ~n25824 ;
  assign n25826 = n25820 & n25825 ;
  assign n25827 = \m7_addr_i[8]_pad  & ~n14069 ;
  assign n25828 = n14062 & n25827 ;
  assign n25829 = \m2_addr_i[8]_pad  & n14069 ;
  assign n25830 = n14086 & n25829 ;
  assign n25831 = ~n25828 & ~n25830 ;
  assign n25832 = \m4_addr_i[8]_pad  & n14069 ;
  assign n25833 = n14077 & n25832 ;
  assign n25834 = \m5_addr_i[8]_pad  & ~n14069 ;
  assign n25835 = n14077 & n25834 ;
  assign n25836 = ~n25833 & ~n25835 ;
  assign n25837 = n25831 & n25836 ;
  assign n25838 = n25826 & n25837 ;
  assign n25839 = \m0_addr_i[9]_pad  & n14069 ;
  assign n25840 = n14094 & n25839 ;
  assign n25841 = \m1_addr_i[9]_pad  & ~n14069 ;
  assign n25842 = n14094 & n25841 ;
  assign n25843 = ~n25840 & ~n25842 ;
  assign n25844 = \m4_addr_i[9]_pad  & n14069 ;
  assign n25845 = n14077 & n25844 ;
  assign n25846 = \m3_addr_i[9]_pad  & ~n14069 ;
  assign n25847 = n14086 & n25846 ;
  assign n25848 = ~n25845 & ~n25847 ;
  assign n25849 = n25843 & n25848 ;
  assign n25850 = \m5_addr_i[9]_pad  & ~n14069 ;
  assign n25851 = n14077 & n25850 ;
  assign n25852 = \m2_addr_i[9]_pad  & n14069 ;
  assign n25853 = n14086 & n25852 ;
  assign n25854 = ~n25851 & ~n25853 ;
  assign n25855 = \m6_addr_i[9]_pad  & n14069 ;
  assign n25856 = n14062 & n25855 ;
  assign n25857 = \m7_addr_i[9]_pad  & ~n14069 ;
  assign n25858 = n14062 & n25857 ;
  assign n25859 = ~n25856 & ~n25858 ;
  assign n25860 = n25854 & n25859 ;
  assign n25861 = n25849 & n25860 ;
  assign n25862 = \m0_data_i[0]_pad  & n14069 ;
  assign n25863 = n14094 & n25862 ;
  assign n25864 = \m1_data_i[0]_pad  & ~n14069 ;
  assign n25865 = n14094 & n25864 ;
  assign n25866 = ~n25863 & ~n25865 ;
  assign n25867 = \m4_data_i[0]_pad  & n14069 ;
  assign n25868 = n14077 & n25867 ;
  assign n25869 = \m3_data_i[0]_pad  & ~n14069 ;
  assign n25870 = n14086 & n25869 ;
  assign n25871 = ~n25868 & ~n25870 ;
  assign n25872 = n25866 & n25871 ;
  assign n25873 = \m5_data_i[0]_pad  & ~n14069 ;
  assign n25874 = n14077 & n25873 ;
  assign n25875 = \m2_data_i[0]_pad  & n14069 ;
  assign n25876 = n14086 & n25875 ;
  assign n25877 = ~n25874 & ~n25876 ;
  assign n25878 = \m6_data_i[0]_pad  & n14069 ;
  assign n25879 = n14062 & n25878 ;
  assign n25880 = \m7_data_i[0]_pad  & ~n14069 ;
  assign n25881 = n14062 & n25880 ;
  assign n25882 = ~n25879 & ~n25881 ;
  assign n25883 = n25877 & n25882 ;
  assign n25884 = n25872 & n25883 ;
  assign n25885 = \m0_data_i[10]_pad  & n14069 ;
  assign n25886 = n14094 & n25885 ;
  assign n25887 = \m1_data_i[10]_pad  & ~n14069 ;
  assign n25888 = n14094 & n25887 ;
  assign n25889 = ~n25886 & ~n25888 ;
  assign n25890 = \m6_data_i[10]_pad  & n14069 ;
  assign n25891 = n14062 & n25890 ;
  assign n25892 = \m3_data_i[10]_pad  & ~n14069 ;
  assign n25893 = n14086 & n25892 ;
  assign n25894 = ~n25891 & ~n25893 ;
  assign n25895 = n25889 & n25894 ;
  assign n25896 = \m7_data_i[10]_pad  & ~n14069 ;
  assign n25897 = n14062 & n25896 ;
  assign n25898 = \m2_data_i[10]_pad  & n14069 ;
  assign n25899 = n14086 & n25898 ;
  assign n25900 = ~n25897 & ~n25899 ;
  assign n25901 = \m4_data_i[10]_pad  & n14069 ;
  assign n25902 = n14077 & n25901 ;
  assign n25903 = \m5_data_i[10]_pad  & ~n14069 ;
  assign n25904 = n14077 & n25903 ;
  assign n25905 = ~n25902 & ~n25904 ;
  assign n25906 = n25900 & n25905 ;
  assign n25907 = n25895 & n25906 ;
  assign n25908 = \m2_data_i[11]_pad  & n14069 ;
  assign n25909 = n14086 & n25908 ;
  assign n25910 = \m3_data_i[11]_pad  & ~n14069 ;
  assign n25911 = n14086 & n25910 ;
  assign n25912 = ~n25909 & ~n25911 ;
  assign n25913 = \m6_data_i[11]_pad  & n14069 ;
  assign n25914 = n14062 & n25913 ;
  assign n25915 = \m1_data_i[11]_pad  & ~n14069 ;
  assign n25916 = n14094 & n25915 ;
  assign n25917 = ~n25914 & ~n25916 ;
  assign n25918 = n25912 & n25917 ;
  assign n25919 = \m7_data_i[11]_pad  & ~n14069 ;
  assign n25920 = n14062 & n25919 ;
  assign n25921 = \m0_data_i[11]_pad  & n14069 ;
  assign n25922 = n14094 & n25921 ;
  assign n25923 = ~n25920 & ~n25922 ;
  assign n25924 = \m4_data_i[11]_pad  & n14069 ;
  assign n25925 = n14077 & n25924 ;
  assign n25926 = \m5_data_i[11]_pad  & ~n14069 ;
  assign n25927 = n14077 & n25926 ;
  assign n25928 = ~n25925 & ~n25927 ;
  assign n25929 = n25923 & n25928 ;
  assign n25930 = n25918 & n25929 ;
  assign n25931 = \m0_data_i[12]_pad  & n14069 ;
  assign n25932 = n14094 & n25931 ;
  assign n25933 = \m1_data_i[12]_pad  & ~n14069 ;
  assign n25934 = n14094 & n25933 ;
  assign n25935 = ~n25932 & ~n25934 ;
  assign n25936 = \m4_data_i[12]_pad  & n14069 ;
  assign n25937 = n14077 & n25936 ;
  assign n25938 = \m3_data_i[12]_pad  & ~n14069 ;
  assign n25939 = n14086 & n25938 ;
  assign n25940 = ~n25937 & ~n25939 ;
  assign n25941 = n25935 & n25940 ;
  assign n25942 = \m5_data_i[12]_pad  & ~n14069 ;
  assign n25943 = n14077 & n25942 ;
  assign n25944 = \m2_data_i[12]_pad  & n14069 ;
  assign n25945 = n14086 & n25944 ;
  assign n25946 = ~n25943 & ~n25945 ;
  assign n25947 = \m6_data_i[12]_pad  & n14069 ;
  assign n25948 = n14062 & n25947 ;
  assign n25949 = \m7_data_i[12]_pad  & ~n14069 ;
  assign n25950 = n14062 & n25949 ;
  assign n25951 = ~n25948 & ~n25950 ;
  assign n25952 = n25946 & n25951 ;
  assign n25953 = n25941 & n25952 ;
  assign n25954 = \m0_data_i[13]_pad  & n14069 ;
  assign n25955 = n14094 & n25954 ;
  assign n25956 = \m1_data_i[13]_pad  & ~n14069 ;
  assign n25957 = n14094 & n25956 ;
  assign n25958 = ~n25955 & ~n25957 ;
  assign n25959 = \m2_data_i[13]_pad  & n14069 ;
  assign n25960 = n14086 & n25959 ;
  assign n25961 = \m7_data_i[13]_pad  & ~n14069 ;
  assign n25962 = n14062 & n25961 ;
  assign n25963 = ~n25960 & ~n25962 ;
  assign n25964 = n25958 & n25963 ;
  assign n25965 = \m3_data_i[13]_pad  & ~n14069 ;
  assign n25966 = n14086 & n25965 ;
  assign n25967 = \m6_data_i[13]_pad  & n14069 ;
  assign n25968 = n14062 & n25967 ;
  assign n25969 = ~n25966 & ~n25968 ;
  assign n25970 = \m4_data_i[13]_pad  & n14069 ;
  assign n25971 = n14077 & n25970 ;
  assign n25972 = \m5_data_i[13]_pad  & ~n14069 ;
  assign n25973 = n14077 & n25972 ;
  assign n25974 = ~n25971 & ~n25973 ;
  assign n25975 = n25969 & n25974 ;
  assign n25976 = n25964 & n25975 ;
  assign n25977 = \m2_data_i[14]_pad  & n14069 ;
  assign n25978 = n14086 & n25977 ;
  assign n25979 = \m3_data_i[14]_pad  & ~n14069 ;
  assign n25980 = n14086 & n25979 ;
  assign n25981 = ~n25978 & ~n25980 ;
  assign n25982 = \m6_data_i[14]_pad  & n14069 ;
  assign n25983 = n14062 & n25982 ;
  assign n25984 = \m1_data_i[14]_pad  & ~n14069 ;
  assign n25985 = n14094 & n25984 ;
  assign n25986 = ~n25983 & ~n25985 ;
  assign n25987 = n25981 & n25986 ;
  assign n25988 = \m7_data_i[14]_pad  & ~n14069 ;
  assign n25989 = n14062 & n25988 ;
  assign n25990 = \m0_data_i[14]_pad  & n14069 ;
  assign n25991 = n14094 & n25990 ;
  assign n25992 = ~n25989 & ~n25991 ;
  assign n25993 = \m4_data_i[14]_pad  & n14069 ;
  assign n25994 = n14077 & n25993 ;
  assign n25995 = \m5_data_i[14]_pad  & ~n14069 ;
  assign n25996 = n14077 & n25995 ;
  assign n25997 = ~n25994 & ~n25996 ;
  assign n25998 = n25992 & n25997 ;
  assign n25999 = n25987 & n25998 ;
  assign n26000 = \m2_data_i[15]_pad  & n14069 ;
  assign n26001 = n14086 & n26000 ;
  assign n26002 = \m3_data_i[15]_pad  & ~n14069 ;
  assign n26003 = n14086 & n26002 ;
  assign n26004 = ~n26001 & ~n26003 ;
  assign n26005 = \m0_data_i[15]_pad  & n14069 ;
  assign n26006 = n14094 & n26005 ;
  assign n26007 = \m7_data_i[15]_pad  & ~n14069 ;
  assign n26008 = n14062 & n26007 ;
  assign n26009 = ~n26006 & ~n26008 ;
  assign n26010 = n26004 & n26009 ;
  assign n26011 = \m1_data_i[15]_pad  & ~n14069 ;
  assign n26012 = n14094 & n26011 ;
  assign n26013 = \m6_data_i[15]_pad  & n14069 ;
  assign n26014 = n14062 & n26013 ;
  assign n26015 = ~n26012 & ~n26014 ;
  assign n26016 = \m4_data_i[15]_pad  & n14069 ;
  assign n26017 = n14077 & n26016 ;
  assign n26018 = \m5_data_i[15]_pad  & ~n14069 ;
  assign n26019 = n14077 & n26018 ;
  assign n26020 = ~n26017 & ~n26019 ;
  assign n26021 = n26015 & n26020 ;
  assign n26022 = n26010 & n26021 ;
  assign n26023 = \m0_data_i[16]_pad  & n14069 ;
  assign n26024 = n14094 & n26023 ;
  assign n26025 = \m1_data_i[16]_pad  & ~n14069 ;
  assign n26026 = n14094 & n26025 ;
  assign n26027 = ~n26024 & ~n26026 ;
  assign n26028 = \m4_data_i[16]_pad  & n14069 ;
  assign n26029 = n14077 & n26028 ;
  assign n26030 = \m3_data_i[16]_pad  & ~n14069 ;
  assign n26031 = n14086 & n26030 ;
  assign n26032 = ~n26029 & ~n26031 ;
  assign n26033 = n26027 & n26032 ;
  assign n26034 = \m5_data_i[16]_pad  & ~n14069 ;
  assign n26035 = n14077 & n26034 ;
  assign n26036 = \m2_data_i[16]_pad  & n14069 ;
  assign n26037 = n14086 & n26036 ;
  assign n26038 = ~n26035 & ~n26037 ;
  assign n26039 = \m6_data_i[16]_pad  & n14069 ;
  assign n26040 = n14062 & n26039 ;
  assign n26041 = \m7_data_i[16]_pad  & ~n14069 ;
  assign n26042 = n14062 & n26041 ;
  assign n26043 = ~n26040 & ~n26042 ;
  assign n26044 = n26038 & n26043 ;
  assign n26045 = n26033 & n26044 ;
  assign n26046 = \m2_data_i[17]_pad  & n14069 ;
  assign n26047 = n14086 & n26046 ;
  assign n26048 = \m3_data_i[17]_pad  & ~n14069 ;
  assign n26049 = n14086 & n26048 ;
  assign n26050 = ~n26047 & ~n26049 ;
  assign n26051 = \m0_data_i[17]_pad  & n14069 ;
  assign n26052 = n14094 & n26051 ;
  assign n26053 = \m7_data_i[17]_pad  & ~n14069 ;
  assign n26054 = n14062 & n26053 ;
  assign n26055 = ~n26052 & ~n26054 ;
  assign n26056 = n26050 & n26055 ;
  assign n26057 = \m1_data_i[17]_pad  & ~n14069 ;
  assign n26058 = n14094 & n26057 ;
  assign n26059 = \m6_data_i[17]_pad  & n14069 ;
  assign n26060 = n14062 & n26059 ;
  assign n26061 = ~n26058 & ~n26060 ;
  assign n26062 = \m4_data_i[17]_pad  & n14069 ;
  assign n26063 = n14077 & n26062 ;
  assign n26064 = \m5_data_i[17]_pad  & ~n14069 ;
  assign n26065 = n14077 & n26064 ;
  assign n26066 = ~n26063 & ~n26065 ;
  assign n26067 = n26061 & n26066 ;
  assign n26068 = n26056 & n26067 ;
  assign n26069 = \m4_data_i[18]_pad  & n14069 ;
  assign n26070 = n14077 & n26069 ;
  assign n26071 = \m5_data_i[18]_pad  & ~n14069 ;
  assign n26072 = n14077 & n26071 ;
  assign n26073 = ~n26070 & ~n26072 ;
  assign n26074 = \m0_data_i[18]_pad  & n14069 ;
  assign n26075 = n14094 & n26074 ;
  assign n26076 = \m7_data_i[18]_pad  & ~n14069 ;
  assign n26077 = n14062 & n26076 ;
  assign n26078 = ~n26075 & ~n26077 ;
  assign n26079 = n26073 & n26078 ;
  assign n26080 = \m1_data_i[18]_pad  & ~n14069 ;
  assign n26081 = n14094 & n26080 ;
  assign n26082 = \m6_data_i[18]_pad  & n14069 ;
  assign n26083 = n14062 & n26082 ;
  assign n26084 = ~n26081 & ~n26083 ;
  assign n26085 = \m2_data_i[18]_pad  & n14069 ;
  assign n26086 = n14086 & n26085 ;
  assign n26087 = \m3_data_i[18]_pad  & ~n14069 ;
  assign n26088 = n14086 & n26087 ;
  assign n26089 = ~n26086 & ~n26088 ;
  assign n26090 = n26084 & n26089 ;
  assign n26091 = n26079 & n26090 ;
  assign n26092 = \m2_data_i[19]_pad  & n14069 ;
  assign n26093 = n14086 & n26092 ;
  assign n26094 = \m3_data_i[19]_pad  & ~n14069 ;
  assign n26095 = n14086 & n26094 ;
  assign n26096 = ~n26093 & ~n26095 ;
  assign n26097 = \m0_data_i[19]_pad  & n14069 ;
  assign n26098 = n14094 & n26097 ;
  assign n26099 = \m7_data_i[19]_pad  & ~n14069 ;
  assign n26100 = n14062 & n26099 ;
  assign n26101 = ~n26098 & ~n26100 ;
  assign n26102 = n26096 & n26101 ;
  assign n26103 = \m1_data_i[19]_pad  & ~n14069 ;
  assign n26104 = n14094 & n26103 ;
  assign n26105 = \m6_data_i[19]_pad  & n14069 ;
  assign n26106 = n14062 & n26105 ;
  assign n26107 = ~n26104 & ~n26106 ;
  assign n26108 = \m4_data_i[19]_pad  & n14069 ;
  assign n26109 = n14077 & n26108 ;
  assign n26110 = \m5_data_i[19]_pad  & ~n14069 ;
  assign n26111 = n14077 & n26110 ;
  assign n26112 = ~n26109 & ~n26111 ;
  assign n26113 = n26107 & n26112 ;
  assign n26114 = n26102 & n26113 ;
  assign n26115 = \m4_data_i[1]_pad  & n14069 ;
  assign n26116 = n14077 & n26115 ;
  assign n26117 = \m5_data_i[1]_pad  & ~n14069 ;
  assign n26118 = n14077 & n26117 ;
  assign n26119 = ~n26116 & ~n26118 ;
  assign n26120 = \m6_data_i[1]_pad  & n14069 ;
  assign n26121 = n14062 & n26120 ;
  assign n26122 = \m1_data_i[1]_pad  & ~n14069 ;
  assign n26123 = n14094 & n26122 ;
  assign n26124 = ~n26121 & ~n26123 ;
  assign n26125 = n26119 & n26124 ;
  assign n26126 = \m7_data_i[1]_pad  & ~n14069 ;
  assign n26127 = n14062 & n26126 ;
  assign n26128 = \m0_data_i[1]_pad  & n14069 ;
  assign n26129 = n14094 & n26128 ;
  assign n26130 = ~n26127 & ~n26129 ;
  assign n26131 = \m2_data_i[1]_pad  & n14069 ;
  assign n26132 = n14086 & n26131 ;
  assign n26133 = \m3_data_i[1]_pad  & ~n14069 ;
  assign n26134 = n14086 & n26133 ;
  assign n26135 = ~n26132 & ~n26134 ;
  assign n26136 = n26130 & n26135 ;
  assign n26137 = n26125 & n26136 ;
  assign n26138 = \m6_data_i[20]_pad  & n14069 ;
  assign n26139 = n14062 & n26138 ;
  assign n26140 = \m7_data_i[20]_pad  & ~n14069 ;
  assign n26141 = n14062 & n26140 ;
  assign n26142 = ~n26139 & ~n26141 ;
  assign n26143 = \m2_data_i[20]_pad  & n14069 ;
  assign n26144 = n14086 & n26143 ;
  assign n26145 = \m5_data_i[20]_pad  & ~n14069 ;
  assign n26146 = n14077 & n26145 ;
  assign n26147 = ~n26144 & ~n26146 ;
  assign n26148 = n26142 & n26147 ;
  assign n26149 = \m3_data_i[20]_pad  & ~n14069 ;
  assign n26150 = n14086 & n26149 ;
  assign n26151 = \m4_data_i[20]_pad  & n14069 ;
  assign n26152 = n14077 & n26151 ;
  assign n26153 = ~n26150 & ~n26152 ;
  assign n26154 = \m0_data_i[20]_pad  & n14069 ;
  assign n26155 = n14094 & n26154 ;
  assign n26156 = \m1_data_i[20]_pad  & ~n14069 ;
  assign n26157 = n14094 & n26156 ;
  assign n26158 = ~n26155 & ~n26157 ;
  assign n26159 = n26153 & n26158 ;
  assign n26160 = n26148 & n26159 ;
  assign n26161 = \m6_data_i[21]_pad  & n14069 ;
  assign n26162 = n14062 & n26161 ;
  assign n26163 = \m7_data_i[21]_pad  & ~n14069 ;
  assign n26164 = n14062 & n26163 ;
  assign n26165 = ~n26162 & ~n26164 ;
  assign n26166 = \m2_data_i[21]_pad  & n14069 ;
  assign n26167 = n14086 & n26166 ;
  assign n26168 = \m5_data_i[21]_pad  & ~n14069 ;
  assign n26169 = n14077 & n26168 ;
  assign n26170 = ~n26167 & ~n26169 ;
  assign n26171 = n26165 & n26170 ;
  assign n26172 = \m3_data_i[21]_pad  & ~n14069 ;
  assign n26173 = n14086 & n26172 ;
  assign n26174 = \m4_data_i[21]_pad  & n14069 ;
  assign n26175 = n14077 & n26174 ;
  assign n26176 = ~n26173 & ~n26175 ;
  assign n26177 = \m0_data_i[21]_pad  & n14069 ;
  assign n26178 = n14094 & n26177 ;
  assign n26179 = \m1_data_i[21]_pad  & ~n14069 ;
  assign n26180 = n14094 & n26179 ;
  assign n26181 = ~n26178 & ~n26180 ;
  assign n26182 = n26176 & n26181 ;
  assign n26183 = n26171 & n26182 ;
  assign n26184 = \m6_data_i[22]_pad  & n14069 ;
  assign n26185 = n14062 & n26184 ;
  assign n26186 = \m7_data_i[22]_pad  & ~n14069 ;
  assign n26187 = n14062 & n26186 ;
  assign n26188 = ~n26185 & ~n26187 ;
  assign n26189 = \m4_data_i[22]_pad  & n14069 ;
  assign n26190 = n14077 & n26189 ;
  assign n26191 = \m3_data_i[22]_pad  & ~n14069 ;
  assign n26192 = n14086 & n26191 ;
  assign n26193 = ~n26190 & ~n26192 ;
  assign n26194 = n26188 & n26193 ;
  assign n26195 = \m5_data_i[22]_pad  & ~n14069 ;
  assign n26196 = n14077 & n26195 ;
  assign n26197 = \m2_data_i[22]_pad  & n14069 ;
  assign n26198 = n14086 & n26197 ;
  assign n26199 = ~n26196 & ~n26198 ;
  assign n26200 = \m0_data_i[22]_pad  & n14069 ;
  assign n26201 = n14094 & n26200 ;
  assign n26202 = \m1_data_i[22]_pad  & ~n14069 ;
  assign n26203 = n14094 & n26202 ;
  assign n26204 = ~n26201 & ~n26203 ;
  assign n26205 = n26199 & n26204 ;
  assign n26206 = n26194 & n26205 ;
  assign n26207 = \m6_data_i[23]_pad  & n14069 ;
  assign n26208 = n14062 & n26207 ;
  assign n26209 = \m7_data_i[23]_pad  & ~n14069 ;
  assign n26210 = n14062 & n26209 ;
  assign n26211 = ~n26208 & ~n26210 ;
  assign n26212 = \m4_data_i[23]_pad  & n14069 ;
  assign n26213 = n14077 & n26212 ;
  assign n26214 = \m3_data_i[23]_pad  & ~n14069 ;
  assign n26215 = n14086 & n26214 ;
  assign n26216 = ~n26213 & ~n26215 ;
  assign n26217 = n26211 & n26216 ;
  assign n26218 = \m5_data_i[23]_pad  & ~n14069 ;
  assign n26219 = n14077 & n26218 ;
  assign n26220 = \m2_data_i[23]_pad  & n14069 ;
  assign n26221 = n14086 & n26220 ;
  assign n26222 = ~n26219 & ~n26221 ;
  assign n26223 = \m0_data_i[23]_pad  & n14069 ;
  assign n26224 = n14094 & n26223 ;
  assign n26225 = \m1_data_i[23]_pad  & ~n14069 ;
  assign n26226 = n14094 & n26225 ;
  assign n26227 = ~n26224 & ~n26226 ;
  assign n26228 = n26222 & n26227 ;
  assign n26229 = n26217 & n26228 ;
  assign n26230 = \m0_data_i[24]_pad  & n14069 ;
  assign n26231 = n14094 & n26230 ;
  assign n26232 = \m1_data_i[24]_pad  & ~n14069 ;
  assign n26233 = n14094 & n26232 ;
  assign n26234 = ~n26231 & ~n26233 ;
  assign n26235 = \m4_data_i[24]_pad  & n14069 ;
  assign n26236 = n14077 & n26235 ;
  assign n26237 = \m7_data_i[24]_pad  & ~n14069 ;
  assign n26238 = n14062 & n26237 ;
  assign n26239 = ~n26236 & ~n26238 ;
  assign n26240 = n26234 & n26239 ;
  assign n26241 = \m5_data_i[24]_pad  & ~n14069 ;
  assign n26242 = n14077 & n26241 ;
  assign n26243 = \m6_data_i[24]_pad  & n14069 ;
  assign n26244 = n14062 & n26243 ;
  assign n26245 = ~n26242 & ~n26244 ;
  assign n26246 = \m2_data_i[24]_pad  & n14069 ;
  assign n26247 = n14086 & n26246 ;
  assign n26248 = \m3_data_i[24]_pad  & ~n14069 ;
  assign n26249 = n14086 & n26248 ;
  assign n26250 = ~n26247 & ~n26249 ;
  assign n26251 = n26245 & n26250 ;
  assign n26252 = n26240 & n26251 ;
  assign n26253 = \m0_data_i[25]_pad  & n14069 ;
  assign n26254 = n14094 & n26253 ;
  assign n26255 = \m1_data_i[25]_pad  & ~n14069 ;
  assign n26256 = n14094 & n26255 ;
  assign n26257 = ~n26254 & ~n26256 ;
  assign n26258 = \m6_data_i[25]_pad  & n14069 ;
  assign n26259 = n14062 & n26258 ;
  assign n26260 = \m3_data_i[25]_pad  & ~n14069 ;
  assign n26261 = n14086 & n26260 ;
  assign n26262 = ~n26259 & ~n26261 ;
  assign n26263 = n26257 & n26262 ;
  assign n26264 = \m7_data_i[25]_pad  & ~n14069 ;
  assign n26265 = n14062 & n26264 ;
  assign n26266 = \m2_data_i[25]_pad  & n14069 ;
  assign n26267 = n14086 & n26266 ;
  assign n26268 = ~n26265 & ~n26267 ;
  assign n26269 = \m4_data_i[25]_pad  & n14069 ;
  assign n26270 = n14077 & n26269 ;
  assign n26271 = \m5_data_i[25]_pad  & ~n14069 ;
  assign n26272 = n14077 & n26271 ;
  assign n26273 = ~n26270 & ~n26272 ;
  assign n26274 = n26268 & n26273 ;
  assign n26275 = n26263 & n26274 ;
  assign n26276 = \m6_data_i[26]_pad  & n14069 ;
  assign n26277 = n14062 & n26276 ;
  assign n26278 = \m7_data_i[26]_pad  & ~n14069 ;
  assign n26279 = n14062 & n26278 ;
  assign n26280 = ~n26277 & ~n26279 ;
  assign n26281 = \m4_data_i[26]_pad  & n14069 ;
  assign n26282 = n14077 & n26281 ;
  assign n26283 = \m1_data_i[26]_pad  & ~n14069 ;
  assign n26284 = n14094 & n26283 ;
  assign n26285 = ~n26282 & ~n26284 ;
  assign n26286 = n26280 & n26285 ;
  assign n26287 = \m5_data_i[26]_pad  & ~n14069 ;
  assign n26288 = n14077 & n26287 ;
  assign n26289 = \m0_data_i[26]_pad  & n14069 ;
  assign n26290 = n14094 & n26289 ;
  assign n26291 = ~n26288 & ~n26290 ;
  assign n26292 = \m2_data_i[26]_pad  & n14069 ;
  assign n26293 = n14086 & n26292 ;
  assign n26294 = \m3_data_i[26]_pad  & ~n14069 ;
  assign n26295 = n14086 & n26294 ;
  assign n26296 = ~n26293 & ~n26295 ;
  assign n26297 = n26291 & n26296 ;
  assign n26298 = n26286 & n26297 ;
  assign n26299 = \m6_data_i[27]_pad  & n14069 ;
  assign n26300 = n14062 & n26299 ;
  assign n26301 = \m7_data_i[27]_pad  & ~n14069 ;
  assign n26302 = n14062 & n26301 ;
  assign n26303 = ~n26300 & ~n26302 ;
  assign n26304 = \m4_data_i[27]_pad  & n14069 ;
  assign n26305 = n14077 & n26304 ;
  assign n26306 = \m3_data_i[27]_pad  & ~n14069 ;
  assign n26307 = n14086 & n26306 ;
  assign n26308 = ~n26305 & ~n26307 ;
  assign n26309 = n26303 & n26308 ;
  assign n26310 = \m5_data_i[27]_pad  & ~n14069 ;
  assign n26311 = n14077 & n26310 ;
  assign n26312 = \m2_data_i[27]_pad  & n14069 ;
  assign n26313 = n14086 & n26312 ;
  assign n26314 = ~n26311 & ~n26313 ;
  assign n26315 = \m0_data_i[27]_pad  & n14069 ;
  assign n26316 = n14094 & n26315 ;
  assign n26317 = \m1_data_i[27]_pad  & ~n14069 ;
  assign n26318 = n14094 & n26317 ;
  assign n26319 = ~n26316 & ~n26318 ;
  assign n26320 = n26314 & n26319 ;
  assign n26321 = n26309 & n26320 ;
  assign n26322 = \m4_data_i[28]_pad  & n14069 ;
  assign n26323 = n14077 & n26322 ;
  assign n26324 = \m5_data_i[28]_pad  & ~n14069 ;
  assign n26325 = n14077 & n26324 ;
  assign n26326 = ~n26323 & ~n26325 ;
  assign n26327 = \m6_data_i[28]_pad  & n14069 ;
  assign n26328 = n14062 & n26327 ;
  assign n26329 = \m1_data_i[28]_pad  & ~n14069 ;
  assign n26330 = n14094 & n26329 ;
  assign n26331 = ~n26328 & ~n26330 ;
  assign n26332 = n26326 & n26331 ;
  assign n26333 = \m7_data_i[28]_pad  & ~n14069 ;
  assign n26334 = n14062 & n26333 ;
  assign n26335 = \m0_data_i[28]_pad  & n14069 ;
  assign n26336 = n14094 & n26335 ;
  assign n26337 = ~n26334 & ~n26336 ;
  assign n26338 = \m2_data_i[28]_pad  & n14069 ;
  assign n26339 = n14086 & n26338 ;
  assign n26340 = \m3_data_i[28]_pad  & ~n14069 ;
  assign n26341 = n14086 & n26340 ;
  assign n26342 = ~n26339 & ~n26341 ;
  assign n26343 = n26337 & n26342 ;
  assign n26344 = n26332 & n26343 ;
  assign n26345 = \m6_data_i[29]_pad  & n14069 ;
  assign n26346 = n14062 & n26345 ;
  assign n26347 = \m7_data_i[29]_pad  & ~n14069 ;
  assign n26348 = n14062 & n26347 ;
  assign n26349 = ~n26346 & ~n26348 ;
  assign n26350 = \m4_data_i[29]_pad  & n14069 ;
  assign n26351 = n14077 & n26350 ;
  assign n26352 = \m3_data_i[29]_pad  & ~n14069 ;
  assign n26353 = n14086 & n26352 ;
  assign n26354 = ~n26351 & ~n26353 ;
  assign n26355 = n26349 & n26354 ;
  assign n26356 = \m5_data_i[29]_pad  & ~n14069 ;
  assign n26357 = n14077 & n26356 ;
  assign n26358 = \m2_data_i[29]_pad  & n14069 ;
  assign n26359 = n14086 & n26358 ;
  assign n26360 = ~n26357 & ~n26359 ;
  assign n26361 = \m0_data_i[29]_pad  & n14069 ;
  assign n26362 = n14094 & n26361 ;
  assign n26363 = \m1_data_i[29]_pad  & ~n14069 ;
  assign n26364 = n14094 & n26363 ;
  assign n26365 = ~n26362 & ~n26364 ;
  assign n26366 = n26360 & n26365 ;
  assign n26367 = n26355 & n26366 ;
  assign n26368 = \m0_data_i[2]_pad  & n14069 ;
  assign n26369 = n14094 & n26368 ;
  assign n26370 = \m1_data_i[2]_pad  & ~n14069 ;
  assign n26371 = n14094 & n26370 ;
  assign n26372 = ~n26369 & ~n26371 ;
  assign n26373 = \m2_data_i[2]_pad  & n14069 ;
  assign n26374 = n14086 & n26373 ;
  assign n26375 = \m7_data_i[2]_pad  & ~n14069 ;
  assign n26376 = n14062 & n26375 ;
  assign n26377 = ~n26374 & ~n26376 ;
  assign n26378 = n26372 & n26377 ;
  assign n26379 = \m3_data_i[2]_pad  & ~n14069 ;
  assign n26380 = n14086 & n26379 ;
  assign n26381 = \m6_data_i[2]_pad  & n14069 ;
  assign n26382 = n14062 & n26381 ;
  assign n26383 = ~n26380 & ~n26382 ;
  assign n26384 = \m4_data_i[2]_pad  & n14069 ;
  assign n26385 = n14077 & n26384 ;
  assign n26386 = \m5_data_i[2]_pad  & ~n14069 ;
  assign n26387 = n14077 & n26386 ;
  assign n26388 = ~n26385 & ~n26387 ;
  assign n26389 = n26383 & n26388 ;
  assign n26390 = n26378 & n26389 ;
  assign n26391 = \m4_data_i[30]_pad  & n14069 ;
  assign n26392 = n14077 & n26391 ;
  assign n26393 = \m5_data_i[30]_pad  & ~n14069 ;
  assign n26394 = n14077 & n26393 ;
  assign n26395 = ~n26392 & ~n26394 ;
  assign n26396 = \m0_data_i[30]_pad  & n14069 ;
  assign n26397 = n14094 & n26396 ;
  assign n26398 = \m3_data_i[30]_pad  & ~n14069 ;
  assign n26399 = n14086 & n26398 ;
  assign n26400 = ~n26397 & ~n26399 ;
  assign n26401 = n26395 & n26400 ;
  assign n26402 = \m1_data_i[30]_pad  & ~n14069 ;
  assign n26403 = n14094 & n26402 ;
  assign n26404 = \m2_data_i[30]_pad  & n14069 ;
  assign n26405 = n14086 & n26404 ;
  assign n26406 = ~n26403 & ~n26405 ;
  assign n26407 = \m6_data_i[30]_pad  & n14069 ;
  assign n26408 = n14062 & n26407 ;
  assign n26409 = \m7_data_i[30]_pad  & ~n14069 ;
  assign n26410 = n14062 & n26409 ;
  assign n26411 = ~n26408 & ~n26410 ;
  assign n26412 = n26406 & n26411 ;
  assign n26413 = n26401 & n26412 ;
  assign n26414 = \m6_data_i[31]_pad  & n14069 ;
  assign n26415 = n14062 & n26414 ;
  assign n26416 = \m7_data_i[31]_pad  & ~n14069 ;
  assign n26417 = n14062 & n26416 ;
  assign n26418 = ~n26415 & ~n26417 ;
  assign n26419 = \m4_data_i[31]_pad  & n14069 ;
  assign n26420 = n14077 & n26419 ;
  assign n26421 = \m3_data_i[31]_pad  & ~n14069 ;
  assign n26422 = n14086 & n26421 ;
  assign n26423 = ~n26420 & ~n26422 ;
  assign n26424 = n26418 & n26423 ;
  assign n26425 = \m5_data_i[31]_pad  & ~n14069 ;
  assign n26426 = n14077 & n26425 ;
  assign n26427 = \m2_data_i[31]_pad  & n14069 ;
  assign n26428 = n14086 & n26427 ;
  assign n26429 = ~n26426 & ~n26428 ;
  assign n26430 = \m0_data_i[31]_pad  & n14069 ;
  assign n26431 = n14094 & n26430 ;
  assign n26432 = \m1_data_i[31]_pad  & ~n14069 ;
  assign n26433 = n14094 & n26432 ;
  assign n26434 = ~n26431 & ~n26433 ;
  assign n26435 = n26429 & n26434 ;
  assign n26436 = n26424 & n26435 ;
  assign n26437 = \m0_data_i[3]_pad  & n14069 ;
  assign n26438 = n14094 & n26437 ;
  assign n26439 = \m1_data_i[3]_pad  & ~n14069 ;
  assign n26440 = n14094 & n26439 ;
  assign n26441 = ~n26438 & ~n26440 ;
  assign n26442 = \m4_data_i[3]_pad  & n14069 ;
  assign n26443 = n14077 & n26442 ;
  assign n26444 = \m3_data_i[3]_pad  & ~n14069 ;
  assign n26445 = n14086 & n26444 ;
  assign n26446 = ~n26443 & ~n26445 ;
  assign n26447 = n26441 & n26446 ;
  assign n26448 = \m5_data_i[3]_pad  & ~n14069 ;
  assign n26449 = n14077 & n26448 ;
  assign n26450 = \m2_data_i[3]_pad  & n14069 ;
  assign n26451 = n14086 & n26450 ;
  assign n26452 = ~n26449 & ~n26451 ;
  assign n26453 = \m6_data_i[3]_pad  & n14069 ;
  assign n26454 = n14062 & n26453 ;
  assign n26455 = \m7_data_i[3]_pad  & ~n14069 ;
  assign n26456 = n14062 & n26455 ;
  assign n26457 = ~n26454 & ~n26456 ;
  assign n26458 = n26452 & n26457 ;
  assign n26459 = n26447 & n26458 ;
  assign n26460 = \m2_data_i[4]_pad  & n14069 ;
  assign n26461 = n14086 & n26460 ;
  assign n26462 = \m3_data_i[4]_pad  & ~n14069 ;
  assign n26463 = n14086 & n26462 ;
  assign n26464 = ~n26461 & ~n26463 ;
  assign n26465 = \m4_data_i[4]_pad  & n14069 ;
  assign n26466 = n14077 & n26465 ;
  assign n26467 = \m1_data_i[4]_pad  & ~n14069 ;
  assign n26468 = n14094 & n26467 ;
  assign n26469 = ~n26466 & ~n26468 ;
  assign n26470 = n26464 & n26469 ;
  assign n26471 = \m5_data_i[4]_pad  & ~n14069 ;
  assign n26472 = n14077 & n26471 ;
  assign n26473 = \m0_data_i[4]_pad  & n14069 ;
  assign n26474 = n14094 & n26473 ;
  assign n26475 = ~n26472 & ~n26474 ;
  assign n26476 = \m6_data_i[4]_pad  & n14069 ;
  assign n26477 = n14062 & n26476 ;
  assign n26478 = \m7_data_i[4]_pad  & ~n14069 ;
  assign n26479 = n14062 & n26478 ;
  assign n26480 = ~n26477 & ~n26479 ;
  assign n26481 = n26475 & n26480 ;
  assign n26482 = n26470 & n26481 ;
  assign n26483 = \m6_data_i[5]_pad  & n14069 ;
  assign n26484 = n14062 & n26483 ;
  assign n26485 = \m7_data_i[5]_pad  & ~n14069 ;
  assign n26486 = n14062 & n26485 ;
  assign n26487 = ~n26484 & ~n26486 ;
  assign n26488 = \m4_data_i[5]_pad  & n14069 ;
  assign n26489 = n14077 & n26488 ;
  assign n26490 = \m3_data_i[5]_pad  & ~n14069 ;
  assign n26491 = n14086 & n26490 ;
  assign n26492 = ~n26489 & ~n26491 ;
  assign n26493 = n26487 & n26492 ;
  assign n26494 = \m5_data_i[5]_pad  & ~n14069 ;
  assign n26495 = n14077 & n26494 ;
  assign n26496 = \m2_data_i[5]_pad  & n14069 ;
  assign n26497 = n14086 & n26496 ;
  assign n26498 = ~n26495 & ~n26497 ;
  assign n26499 = \m0_data_i[5]_pad  & n14069 ;
  assign n26500 = n14094 & n26499 ;
  assign n26501 = \m1_data_i[5]_pad  & ~n14069 ;
  assign n26502 = n14094 & n26501 ;
  assign n26503 = ~n26500 & ~n26502 ;
  assign n26504 = n26498 & n26503 ;
  assign n26505 = n26493 & n26504 ;
  assign n26506 = \m2_data_i[6]_pad  & n14069 ;
  assign n26507 = n14086 & n26506 ;
  assign n26508 = \m3_data_i[6]_pad  & ~n14069 ;
  assign n26509 = n14086 & n26508 ;
  assign n26510 = ~n26507 & ~n26509 ;
  assign n26511 = \m6_data_i[6]_pad  & n14069 ;
  assign n26512 = n14062 & n26511 ;
  assign n26513 = \m1_data_i[6]_pad  & ~n14069 ;
  assign n26514 = n14094 & n26513 ;
  assign n26515 = ~n26512 & ~n26514 ;
  assign n26516 = n26510 & n26515 ;
  assign n26517 = \m7_data_i[6]_pad  & ~n14069 ;
  assign n26518 = n14062 & n26517 ;
  assign n26519 = \m0_data_i[6]_pad  & n14069 ;
  assign n26520 = n14094 & n26519 ;
  assign n26521 = ~n26518 & ~n26520 ;
  assign n26522 = \m4_data_i[6]_pad  & n14069 ;
  assign n26523 = n14077 & n26522 ;
  assign n26524 = \m5_data_i[6]_pad  & ~n14069 ;
  assign n26525 = n14077 & n26524 ;
  assign n26526 = ~n26523 & ~n26525 ;
  assign n26527 = n26521 & n26526 ;
  assign n26528 = n26516 & n26527 ;
  assign n26529 = \m6_data_i[7]_pad  & n14069 ;
  assign n26530 = n14062 & n26529 ;
  assign n26531 = \m7_data_i[7]_pad  & ~n14069 ;
  assign n26532 = n14062 & n26531 ;
  assign n26533 = ~n26530 & ~n26532 ;
  assign n26534 = \m4_data_i[7]_pad  & n14069 ;
  assign n26535 = n14077 & n26534 ;
  assign n26536 = \m1_data_i[7]_pad  & ~n14069 ;
  assign n26537 = n14094 & n26536 ;
  assign n26538 = ~n26535 & ~n26537 ;
  assign n26539 = n26533 & n26538 ;
  assign n26540 = \m5_data_i[7]_pad  & ~n14069 ;
  assign n26541 = n14077 & n26540 ;
  assign n26542 = \m0_data_i[7]_pad  & n14069 ;
  assign n26543 = n14094 & n26542 ;
  assign n26544 = ~n26541 & ~n26543 ;
  assign n26545 = \m2_data_i[7]_pad  & n14069 ;
  assign n26546 = n14086 & n26545 ;
  assign n26547 = \m3_data_i[7]_pad  & ~n14069 ;
  assign n26548 = n14086 & n26547 ;
  assign n26549 = ~n26546 & ~n26548 ;
  assign n26550 = n26544 & n26549 ;
  assign n26551 = n26539 & n26550 ;
  assign n26552 = \m6_data_i[8]_pad  & n14069 ;
  assign n26553 = n14062 & n26552 ;
  assign n26554 = \m7_data_i[8]_pad  & ~n14069 ;
  assign n26555 = n14062 & n26554 ;
  assign n26556 = ~n26553 & ~n26555 ;
  assign n26557 = \m4_data_i[8]_pad  & n14069 ;
  assign n26558 = n14077 & n26557 ;
  assign n26559 = \m1_data_i[8]_pad  & ~n14069 ;
  assign n26560 = n14094 & n26559 ;
  assign n26561 = ~n26558 & ~n26560 ;
  assign n26562 = n26556 & n26561 ;
  assign n26563 = \m5_data_i[8]_pad  & ~n14069 ;
  assign n26564 = n14077 & n26563 ;
  assign n26565 = \m0_data_i[8]_pad  & n14069 ;
  assign n26566 = n14094 & n26565 ;
  assign n26567 = ~n26564 & ~n26566 ;
  assign n26568 = \m2_data_i[8]_pad  & n14069 ;
  assign n26569 = n14086 & n26568 ;
  assign n26570 = \m3_data_i[8]_pad  & ~n14069 ;
  assign n26571 = n14086 & n26570 ;
  assign n26572 = ~n26569 & ~n26571 ;
  assign n26573 = n26567 & n26572 ;
  assign n26574 = n26562 & n26573 ;
  assign n26575 = \m6_data_i[9]_pad  & n14069 ;
  assign n26576 = n14062 & n26575 ;
  assign n26577 = \m7_data_i[9]_pad  & ~n14069 ;
  assign n26578 = n14062 & n26577 ;
  assign n26579 = ~n26576 & ~n26578 ;
  assign n26580 = \m4_data_i[9]_pad  & n14069 ;
  assign n26581 = n14077 & n26580 ;
  assign n26582 = \m1_data_i[9]_pad  & ~n14069 ;
  assign n26583 = n14094 & n26582 ;
  assign n26584 = ~n26581 & ~n26583 ;
  assign n26585 = n26579 & n26584 ;
  assign n26586 = \m5_data_i[9]_pad  & ~n14069 ;
  assign n26587 = n14077 & n26586 ;
  assign n26588 = \m0_data_i[9]_pad  & n14069 ;
  assign n26589 = n14094 & n26588 ;
  assign n26590 = ~n26587 & ~n26589 ;
  assign n26591 = \m2_data_i[9]_pad  & n14069 ;
  assign n26592 = n14086 & n26591 ;
  assign n26593 = \m3_data_i[9]_pad  & ~n14069 ;
  assign n26594 = n14086 & n26593 ;
  assign n26595 = ~n26592 & ~n26594 ;
  assign n26596 = n26590 & n26595 ;
  assign n26597 = n26585 & n26596 ;
  assign n26598 = \m2_sel_i[0]_pad  & n14069 ;
  assign n26599 = n14086 & n26598 ;
  assign n26600 = \m3_sel_i[0]_pad  & ~n14069 ;
  assign n26601 = n14086 & n26600 ;
  assign n26602 = ~n26599 & ~n26601 ;
  assign n26603 = \m0_sel_i[0]_pad  & n14069 ;
  assign n26604 = n14094 & n26603 ;
  assign n26605 = \m7_sel_i[0]_pad  & ~n14069 ;
  assign n26606 = n14062 & n26605 ;
  assign n26607 = ~n26604 & ~n26606 ;
  assign n26608 = n26602 & n26607 ;
  assign n26609 = \m1_sel_i[0]_pad  & ~n14069 ;
  assign n26610 = n14094 & n26609 ;
  assign n26611 = \m6_sel_i[0]_pad  & n14069 ;
  assign n26612 = n14062 & n26611 ;
  assign n26613 = ~n26610 & ~n26612 ;
  assign n26614 = \m4_sel_i[0]_pad  & n14069 ;
  assign n26615 = n14077 & n26614 ;
  assign n26616 = \m5_sel_i[0]_pad  & ~n14069 ;
  assign n26617 = n14077 & n26616 ;
  assign n26618 = ~n26615 & ~n26617 ;
  assign n26619 = n26613 & n26618 ;
  assign n26620 = n26608 & n26619 ;
  assign n26621 = \m0_sel_i[1]_pad  & n14069 ;
  assign n26622 = n14094 & n26621 ;
  assign n26623 = \m1_sel_i[1]_pad  & ~n14069 ;
  assign n26624 = n14094 & n26623 ;
  assign n26625 = ~n26622 & ~n26624 ;
  assign n26626 = \m6_sel_i[1]_pad  & n14069 ;
  assign n26627 = n14062 & n26626 ;
  assign n26628 = \m3_sel_i[1]_pad  & ~n14069 ;
  assign n26629 = n14086 & n26628 ;
  assign n26630 = ~n26627 & ~n26629 ;
  assign n26631 = n26625 & n26630 ;
  assign n26632 = \m7_sel_i[1]_pad  & ~n14069 ;
  assign n26633 = n14062 & n26632 ;
  assign n26634 = \m2_sel_i[1]_pad  & n14069 ;
  assign n26635 = n14086 & n26634 ;
  assign n26636 = ~n26633 & ~n26635 ;
  assign n26637 = \m4_sel_i[1]_pad  & n14069 ;
  assign n26638 = n14077 & n26637 ;
  assign n26639 = \m5_sel_i[1]_pad  & ~n14069 ;
  assign n26640 = n14077 & n26639 ;
  assign n26641 = ~n26638 & ~n26640 ;
  assign n26642 = n26636 & n26641 ;
  assign n26643 = n26631 & n26642 ;
  assign n26644 = \m2_sel_i[2]_pad  & n14069 ;
  assign n26645 = n14086 & n26644 ;
  assign n26646 = \m3_sel_i[2]_pad  & ~n14069 ;
  assign n26647 = n14086 & n26646 ;
  assign n26648 = ~n26645 & ~n26647 ;
  assign n26649 = \m0_sel_i[2]_pad  & n14069 ;
  assign n26650 = n14094 & n26649 ;
  assign n26651 = \m5_sel_i[2]_pad  & ~n14069 ;
  assign n26652 = n14077 & n26651 ;
  assign n26653 = ~n26650 & ~n26652 ;
  assign n26654 = n26648 & n26653 ;
  assign n26655 = \m1_sel_i[2]_pad  & ~n14069 ;
  assign n26656 = n14094 & n26655 ;
  assign n26657 = \m4_sel_i[2]_pad  & n14069 ;
  assign n26658 = n14077 & n26657 ;
  assign n26659 = ~n26656 & ~n26658 ;
  assign n26660 = \m6_sel_i[2]_pad  & n14069 ;
  assign n26661 = n14062 & n26660 ;
  assign n26662 = \m7_sel_i[2]_pad  & ~n14069 ;
  assign n26663 = n14062 & n26662 ;
  assign n26664 = ~n26661 & ~n26663 ;
  assign n26665 = n26659 & n26664 ;
  assign n26666 = n26654 & n26665 ;
  assign n26667 = \m2_sel_i[3]_pad  & n14069 ;
  assign n26668 = n14086 & n26667 ;
  assign n26669 = \m3_sel_i[3]_pad  & ~n14069 ;
  assign n26670 = n14086 & n26669 ;
  assign n26671 = ~n26668 & ~n26670 ;
  assign n26672 = \m0_sel_i[3]_pad  & n14069 ;
  assign n26673 = n14094 & n26672 ;
  assign n26674 = \m7_sel_i[3]_pad  & ~n14069 ;
  assign n26675 = n14062 & n26674 ;
  assign n26676 = ~n26673 & ~n26675 ;
  assign n26677 = n26671 & n26676 ;
  assign n26678 = \m1_sel_i[3]_pad  & ~n14069 ;
  assign n26679 = n14094 & n26678 ;
  assign n26680 = \m6_sel_i[3]_pad  & n14069 ;
  assign n26681 = n14062 & n26680 ;
  assign n26682 = ~n26679 & ~n26681 ;
  assign n26683 = \m4_sel_i[3]_pad  & n14069 ;
  assign n26684 = n14077 & n26683 ;
  assign n26685 = \m5_sel_i[3]_pad  & ~n14069 ;
  assign n26686 = n14077 & n26685 ;
  assign n26687 = ~n26684 & ~n26686 ;
  assign n26688 = n26682 & n26687 ;
  assign n26689 = n26677 & n26688 ;
  assign n26690 = \m1_stb_i_pad  & n14582 ;
  assign n26691 = ~n14069 & n26690 ;
  assign n26692 = n14094 & n26691 ;
  assign n26693 = \m7_stb_i_pad  & n14647 ;
  assign n26694 = ~n14069 & n26693 ;
  assign n26695 = n14062 & n26694 ;
  assign n26696 = ~n26692 & ~n26695 ;
  assign n26697 = \m2_stb_i_pad  & n14590 ;
  assign n26698 = n14069 & n26697 ;
  assign n26699 = n14086 & n26698 ;
  assign n26700 = \m3_stb_i_pad  & n14603 ;
  assign n26701 = ~n14069 & n26700 ;
  assign n26702 = n14086 & n26701 ;
  assign n26703 = ~n26699 & ~n26702 ;
  assign n26704 = n26696 & n26703 ;
  assign n26705 = \m0_stb_i_pad  & n14569 ;
  assign n26706 = n14069 & n26705 ;
  assign n26707 = n14094 & n26706 ;
  assign n26708 = \m5_stb_i_pad  & n14627 ;
  assign n26709 = ~n14069 & n26708 ;
  assign n26710 = n14077 & n26709 ;
  assign n26711 = ~n26707 & ~n26710 ;
  assign n26712 = \m4_stb_i_pad  & n14616 ;
  assign n26713 = n14069 & n26712 ;
  assign n26714 = n14077 & n26713 ;
  assign n26715 = \m6_stb_i_pad  & n14634 ;
  assign n26716 = n14069 & n26715 ;
  assign n26717 = n14062 & n26716 ;
  assign n26718 = ~n26714 & ~n26717 ;
  assign n26719 = n26711 & n26718 ;
  assign n26720 = n26704 & n26719 ;
  assign n26721 = \m2_we_i_pad  & n14069 ;
  assign n26722 = n14086 & n26721 ;
  assign n26723 = \m3_we_i_pad  & ~n14069 ;
  assign n26724 = n14086 & n26723 ;
  assign n26725 = ~n26722 & ~n26724 ;
  assign n26726 = \m0_we_i_pad  & n14069 ;
  assign n26727 = n14094 & n26726 ;
  assign n26728 = \m7_we_i_pad  & ~n14069 ;
  assign n26729 = n14062 & n26728 ;
  assign n26730 = ~n26727 & ~n26729 ;
  assign n26731 = n26725 & n26730 ;
  assign n26732 = \m1_we_i_pad  & ~n14069 ;
  assign n26733 = n14094 & n26732 ;
  assign n26734 = \m6_we_i_pad  & n14069 ;
  assign n26735 = n14062 & n26734 ;
  assign n26736 = ~n26733 & ~n26735 ;
  assign n26737 = \m4_we_i_pad  & n14069 ;
  assign n26738 = n14077 & n26737 ;
  assign n26739 = \m5_we_i_pad  & ~n14069 ;
  assign n26740 = n14077 & n26739 ;
  assign n26741 = ~n26738 & ~n26740 ;
  assign n26742 = n26736 & n26741 ;
  assign n26743 = n26731 & n26742 ;
  assign n26744 = \m1_addr_i[0]_pad  & ~n13928 ;
  assign n26745 = n13945 & n26744 ;
  assign n26746 = \m2_addr_i[0]_pad  & n13928 ;
  assign n26747 = n13921 & n26746 ;
  assign n26748 = ~n26745 & ~n26747 ;
  assign n26749 = \m0_addr_i[0]_pad  & n13928 ;
  assign n26750 = n13945 & n26749 ;
  assign n26751 = \m4_addr_i[0]_pad  & n13928 ;
  assign n26752 = n13953 & n26751 ;
  assign n26753 = ~n26750 & ~n26752 ;
  assign n26754 = n26748 & n26753 ;
  assign n26755 = \m7_addr_i[0]_pad  & ~n13928 ;
  assign n26756 = n13936 & n26755 ;
  assign n26757 = \m3_addr_i[0]_pad  & ~n13928 ;
  assign n26758 = n13921 & n26757 ;
  assign n26759 = ~n26756 & ~n26758 ;
  assign n26760 = \m6_addr_i[0]_pad  & n13928 ;
  assign n26761 = n13936 & n26760 ;
  assign n26762 = \m5_addr_i[0]_pad  & ~n13928 ;
  assign n26763 = n13953 & n26762 ;
  assign n26764 = ~n26761 & ~n26763 ;
  assign n26765 = n26759 & n26764 ;
  assign n26766 = n26754 & n26765 ;
  assign n26767 = \m1_addr_i[10]_pad  & ~n13928 ;
  assign n26768 = n13945 & n26767 ;
  assign n26769 = \m2_addr_i[10]_pad  & n13928 ;
  assign n26770 = n13921 & n26769 ;
  assign n26771 = ~n26768 & ~n26770 ;
  assign n26772 = \m6_addr_i[10]_pad  & n13928 ;
  assign n26773 = n13936 & n26772 ;
  assign n26774 = \m4_addr_i[10]_pad  & n13928 ;
  assign n26775 = n13953 & n26774 ;
  assign n26776 = ~n26773 & ~n26775 ;
  assign n26777 = n26771 & n26776 ;
  assign n26778 = \m5_addr_i[10]_pad  & ~n13928 ;
  assign n26779 = n13953 & n26778 ;
  assign n26780 = \m3_addr_i[10]_pad  & ~n13928 ;
  assign n26781 = n13921 & n26780 ;
  assign n26782 = ~n26779 & ~n26781 ;
  assign n26783 = \m0_addr_i[10]_pad  & n13928 ;
  assign n26784 = n13945 & n26783 ;
  assign n26785 = \m7_addr_i[10]_pad  & ~n13928 ;
  assign n26786 = n13936 & n26785 ;
  assign n26787 = ~n26784 & ~n26786 ;
  assign n26788 = n26782 & n26787 ;
  assign n26789 = n26777 & n26788 ;
  assign n26790 = \m3_addr_i[11]_pad  & ~n13928 ;
  assign n26791 = n13921 & n26790 ;
  assign n26792 = \m4_addr_i[11]_pad  & n13928 ;
  assign n26793 = n13953 & n26792 ;
  assign n26794 = ~n26791 & ~n26793 ;
  assign n26795 = \m0_addr_i[11]_pad  & n13928 ;
  assign n26796 = n13945 & n26795 ;
  assign n26797 = \m2_addr_i[11]_pad  & n13928 ;
  assign n26798 = n13921 & n26797 ;
  assign n26799 = ~n26796 & ~n26798 ;
  assign n26800 = n26794 & n26799 ;
  assign n26801 = \m7_addr_i[11]_pad  & ~n13928 ;
  assign n26802 = n13936 & n26801 ;
  assign n26803 = \m1_addr_i[11]_pad  & ~n13928 ;
  assign n26804 = n13945 & n26803 ;
  assign n26805 = ~n26802 & ~n26804 ;
  assign n26806 = \m6_addr_i[11]_pad  & n13928 ;
  assign n26807 = n13936 & n26806 ;
  assign n26808 = \m5_addr_i[11]_pad  & ~n13928 ;
  assign n26809 = n13953 & n26808 ;
  assign n26810 = ~n26807 & ~n26809 ;
  assign n26811 = n26805 & n26810 ;
  assign n26812 = n26800 & n26811 ;
  assign n26813 = \m1_addr_i[12]_pad  & ~n13928 ;
  assign n26814 = n13945 & n26813 ;
  assign n26815 = \m2_addr_i[12]_pad  & n13928 ;
  assign n26816 = n13921 & n26815 ;
  assign n26817 = ~n26814 & ~n26816 ;
  assign n26818 = \m3_addr_i[12]_pad  & ~n13928 ;
  assign n26819 = n13921 & n26818 ;
  assign n26820 = \m7_addr_i[12]_pad  & ~n13928 ;
  assign n26821 = n13936 & n26820 ;
  assign n26822 = ~n26819 & ~n26821 ;
  assign n26823 = n26817 & n26822 ;
  assign n26824 = \m4_addr_i[12]_pad  & n13928 ;
  assign n26825 = n13953 & n26824 ;
  assign n26826 = \m0_addr_i[12]_pad  & n13928 ;
  assign n26827 = n13945 & n26826 ;
  assign n26828 = ~n26825 & ~n26827 ;
  assign n26829 = \m6_addr_i[12]_pad  & n13928 ;
  assign n26830 = n13936 & n26829 ;
  assign n26831 = \m5_addr_i[12]_pad  & ~n13928 ;
  assign n26832 = n13953 & n26831 ;
  assign n26833 = ~n26830 & ~n26832 ;
  assign n26834 = n26828 & n26833 ;
  assign n26835 = n26823 & n26834 ;
  assign n26836 = \m3_addr_i[13]_pad  & ~n13928 ;
  assign n26837 = n13921 & n26836 ;
  assign n26838 = \m4_addr_i[13]_pad  & n13928 ;
  assign n26839 = n13953 & n26838 ;
  assign n26840 = ~n26837 & ~n26839 ;
  assign n26841 = \m0_addr_i[13]_pad  & n13928 ;
  assign n26842 = n13945 & n26841 ;
  assign n26843 = \m5_addr_i[13]_pad  & ~n13928 ;
  assign n26844 = n13953 & n26843 ;
  assign n26845 = ~n26842 & ~n26844 ;
  assign n26846 = n26840 & n26845 ;
  assign n26847 = \m7_addr_i[13]_pad  & ~n13928 ;
  assign n26848 = n13936 & n26847 ;
  assign n26849 = \m6_addr_i[13]_pad  & n13928 ;
  assign n26850 = n13936 & n26849 ;
  assign n26851 = ~n26848 & ~n26850 ;
  assign n26852 = \m1_addr_i[13]_pad  & ~n13928 ;
  assign n26853 = n13945 & n26852 ;
  assign n26854 = \m2_addr_i[13]_pad  & n13928 ;
  assign n26855 = n13921 & n26854 ;
  assign n26856 = ~n26853 & ~n26855 ;
  assign n26857 = n26851 & n26856 ;
  assign n26858 = n26846 & n26857 ;
  assign n26859 = \m3_addr_i[14]_pad  & ~n13928 ;
  assign n26860 = n13921 & n26859 ;
  assign n26861 = \m4_addr_i[14]_pad  & n13928 ;
  assign n26862 = n13953 & n26861 ;
  assign n26863 = ~n26860 & ~n26862 ;
  assign n26864 = \m1_addr_i[14]_pad  & ~n13928 ;
  assign n26865 = n13945 & n26864 ;
  assign n26866 = \m5_addr_i[14]_pad  & ~n13928 ;
  assign n26867 = n13953 & n26866 ;
  assign n26868 = ~n26865 & ~n26867 ;
  assign n26869 = n26863 & n26868 ;
  assign n26870 = \m2_addr_i[14]_pad  & n13928 ;
  assign n26871 = n13921 & n26870 ;
  assign n26872 = \m6_addr_i[14]_pad  & n13928 ;
  assign n26873 = n13936 & n26872 ;
  assign n26874 = ~n26871 & ~n26873 ;
  assign n26875 = \m0_addr_i[14]_pad  & n13928 ;
  assign n26876 = n13945 & n26875 ;
  assign n26877 = \m7_addr_i[14]_pad  & ~n13928 ;
  assign n26878 = n13936 & n26877 ;
  assign n26879 = ~n26876 & ~n26878 ;
  assign n26880 = n26874 & n26879 ;
  assign n26881 = n26869 & n26880 ;
  assign n26882 = \m1_addr_i[15]_pad  & ~n13928 ;
  assign n26883 = n13945 & n26882 ;
  assign n26884 = \m2_addr_i[15]_pad  & n13928 ;
  assign n26885 = n13921 & n26884 ;
  assign n26886 = ~n26883 & ~n26885 ;
  assign n26887 = \m0_addr_i[15]_pad  & n13928 ;
  assign n26888 = n13945 & n26887 ;
  assign n26889 = \m4_addr_i[15]_pad  & n13928 ;
  assign n26890 = n13953 & n26889 ;
  assign n26891 = ~n26888 & ~n26890 ;
  assign n26892 = n26886 & n26891 ;
  assign n26893 = \m7_addr_i[15]_pad  & ~n13928 ;
  assign n26894 = n13936 & n26893 ;
  assign n26895 = \m3_addr_i[15]_pad  & ~n13928 ;
  assign n26896 = n13921 & n26895 ;
  assign n26897 = ~n26894 & ~n26896 ;
  assign n26898 = \m6_addr_i[15]_pad  & n13928 ;
  assign n26899 = n13936 & n26898 ;
  assign n26900 = \m5_addr_i[15]_pad  & ~n13928 ;
  assign n26901 = n13953 & n26900 ;
  assign n26902 = ~n26899 & ~n26901 ;
  assign n26903 = n26897 & n26902 ;
  assign n26904 = n26892 & n26903 ;
  assign n26905 = \m6_addr_i[16]_pad  & n13928 ;
  assign n26906 = n13936 & n26905 ;
  assign n26907 = \m5_addr_i[16]_pad  & ~n13928 ;
  assign n26908 = n13953 & n26907 ;
  assign n26909 = ~n26906 & ~n26908 ;
  assign n26910 = \m0_addr_i[16]_pad  & n13928 ;
  assign n26911 = n13945 & n26910 ;
  assign n26912 = \m4_addr_i[16]_pad  & n13928 ;
  assign n26913 = n13953 & n26912 ;
  assign n26914 = ~n26911 & ~n26913 ;
  assign n26915 = n26909 & n26914 ;
  assign n26916 = \m7_addr_i[16]_pad  & ~n13928 ;
  assign n26917 = n13936 & n26916 ;
  assign n26918 = \m3_addr_i[16]_pad  & ~n13928 ;
  assign n26919 = n13921 & n26918 ;
  assign n26920 = ~n26917 & ~n26919 ;
  assign n26921 = \m1_addr_i[16]_pad  & ~n13928 ;
  assign n26922 = n13945 & n26921 ;
  assign n26923 = \m2_addr_i[16]_pad  & n13928 ;
  assign n26924 = n13921 & n26923 ;
  assign n26925 = ~n26922 & ~n26924 ;
  assign n26926 = n26920 & n26925 ;
  assign n26927 = n26915 & n26926 ;
  assign n26928 = \m0_addr_i[17]_pad  & n13928 ;
  assign n26929 = n13945 & n26928 ;
  assign n26930 = \m7_addr_i[17]_pad  & ~n13928 ;
  assign n26931 = n13936 & n26930 ;
  assign n26932 = ~n26929 & ~n26931 ;
  assign n26933 = \m1_addr_i[17]_pad  & ~n13928 ;
  assign n26934 = n13945 & n26933 ;
  assign n26935 = \m4_addr_i[17]_pad  & n13928 ;
  assign n26936 = n13953 & n26935 ;
  assign n26937 = ~n26934 & ~n26936 ;
  assign n26938 = n26932 & n26937 ;
  assign n26939 = \m2_addr_i[17]_pad  & n13928 ;
  assign n26940 = n13921 & n26939 ;
  assign n26941 = \m3_addr_i[17]_pad  & ~n13928 ;
  assign n26942 = n13921 & n26941 ;
  assign n26943 = ~n26940 & ~n26942 ;
  assign n26944 = \m6_addr_i[17]_pad  & n13928 ;
  assign n26945 = n13936 & n26944 ;
  assign n26946 = \m5_addr_i[17]_pad  & ~n13928 ;
  assign n26947 = n13953 & n26946 ;
  assign n26948 = ~n26945 & ~n26947 ;
  assign n26949 = n26943 & n26948 ;
  assign n26950 = n26938 & n26949 ;
  assign n26951 = \m3_addr_i[18]_pad  & ~n13928 ;
  assign n26952 = n13921 & n26951 ;
  assign n26953 = \m4_addr_i[18]_pad  & n13928 ;
  assign n26954 = n13953 & n26953 ;
  assign n26955 = ~n26952 & ~n26954 ;
  assign n26956 = \m1_addr_i[18]_pad  & ~n13928 ;
  assign n26957 = n13945 & n26956 ;
  assign n26958 = \m5_addr_i[18]_pad  & ~n13928 ;
  assign n26959 = n13953 & n26958 ;
  assign n26960 = ~n26957 & ~n26959 ;
  assign n26961 = n26955 & n26960 ;
  assign n26962 = \m2_addr_i[18]_pad  & n13928 ;
  assign n26963 = n13921 & n26962 ;
  assign n26964 = \m6_addr_i[18]_pad  & n13928 ;
  assign n26965 = n13936 & n26964 ;
  assign n26966 = ~n26963 & ~n26965 ;
  assign n26967 = \m0_addr_i[18]_pad  & n13928 ;
  assign n26968 = n13945 & n26967 ;
  assign n26969 = \m7_addr_i[18]_pad  & ~n13928 ;
  assign n26970 = n13936 & n26969 ;
  assign n26971 = ~n26968 & ~n26970 ;
  assign n26972 = n26966 & n26971 ;
  assign n26973 = n26961 & n26972 ;
  assign n26974 = \m6_addr_i[19]_pad  & n13928 ;
  assign n26975 = n13936 & n26974 ;
  assign n26976 = \m5_addr_i[19]_pad  & ~n13928 ;
  assign n26977 = n13953 & n26976 ;
  assign n26978 = ~n26975 & ~n26977 ;
  assign n26979 = \m0_addr_i[19]_pad  & n13928 ;
  assign n26980 = n13945 & n26979 ;
  assign n26981 = \m4_addr_i[19]_pad  & n13928 ;
  assign n26982 = n13953 & n26981 ;
  assign n26983 = ~n26980 & ~n26982 ;
  assign n26984 = n26978 & n26983 ;
  assign n26985 = \m7_addr_i[19]_pad  & ~n13928 ;
  assign n26986 = n13936 & n26985 ;
  assign n26987 = \m3_addr_i[19]_pad  & ~n13928 ;
  assign n26988 = n13921 & n26987 ;
  assign n26989 = ~n26986 & ~n26988 ;
  assign n26990 = \m1_addr_i[19]_pad  & ~n13928 ;
  assign n26991 = n13945 & n26990 ;
  assign n26992 = \m2_addr_i[19]_pad  & n13928 ;
  assign n26993 = n13921 & n26992 ;
  assign n26994 = ~n26991 & ~n26993 ;
  assign n26995 = n26989 & n26994 ;
  assign n26996 = n26984 & n26995 ;
  assign n26997 = \m0_addr_i[1]_pad  & n13928 ;
  assign n26998 = n13945 & n26997 ;
  assign n26999 = \m7_addr_i[1]_pad  & ~n13928 ;
  assign n27000 = n13936 & n26999 ;
  assign n27001 = ~n26998 & ~n27000 ;
  assign n27002 = \m6_addr_i[1]_pad  & n13928 ;
  assign n27003 = n13936 & n27002 ;
  assign n27004 = \m2_addr_i[1]_pad  & n13928 ;
  assign n27005 = n13921 & n27004 ;
  assign n27006 = ~n27003 & ~n27005 ;
  assign n27007 = n27001 & n27006 ;
  assign n27008 = \m5_addr_i[1]_pad  & ~n13928 ;
  assign n27009 = n13953 & n27008 ;
  assign n27010 = \m1_addr_i[1]_pad  & ~n13928 ;
  assign n27011 = n13945 & n27010 ;
  assign n27012 = ~n27009 & ~n27011 ;
  assign n27013 = \m3_addr_i[1]_pad  & ~n13928 ;
  assign n27014 = n13921 & n27013 ;
  assign n27015 = \m4_addr_i[1]_pad  & n13928 ;
  assign n27016 = n13953 & n27015 ;
  assign n27017 = ~n27014 & ~n27016 ;
  assign n27018 = n27012 & n27017 ;
  assign n27019 = n27007 & n27018 ;
  assign n27020 = \m1_addr_i[20]_pad  & ~n13928 ;
  assign n27021 = n13945 & n27020 ;
  assign n27022 = \m2_addr_i[20]_pad  & n13928 ;
  assign n27023 = n13921 & n27022 ;
  assign n27024 = ~n27021 & ~n27023 ;
  assign n27025 = \m0_addr_i[20]_pad  & n13928 ;
  assign n27026 = n13945 & n27025 ;
  assign n27027 = \m4_addr_i[20]_pad  & n13928 ;
  assign n27028 = n13953 & n27027 ;
  assign n27029 = ~n27026 & ~n27028 ;
  assign n27030 = n27024 & n27029 ;
  assign n27031 = \m7_addr_i[20]_pad  & ~n13928 ;
  assign n27032 = n13936 & n27031 ;
  assign n27033 = \m3_addr_i[20]_pad  & ~n13928 ;
  assign n27034 = n13921 & n27033 ;
  assign n27035 = ~n27032 & ~n27034 ;
  assign n27036 = \m6_addr_i[20]_pad  & n13928 ;
  assign n27037 = n13936 & n27036 ;
  assign n27038 = \m5_addr_i[20]_pad  & ~n13928 ;
  assign n27039 = n13953 & n27038 ;
  assign n27040 = ~n27037 & ~n27039 ;
  assign n27041 = n27035 & n27040 ;
  assign n27042 = n27030 & n27041 ;
  assign n27043 = \m3_addr_i[21]_pad  & ~n13928 ;
  assign n27044 = n13921 & n27043 ;
  assign n27045 = \m4_addr_i[21]_pad  & n13928 ;
  assign n27046 = n13953 & n27045 ;
  assign n27047 = ~n27044 & ~n27046 ;
  assign n27048 = \m1_addr_i[21]_pad  & ~n13928 ;
  assign n27049 = n13945 & n27048 ;
  assign n27050 = \m7_addr_i[21]_pad  & ~n13928 ;
  assign n27051 = n13936 & n27050 ;
  assign n27052 = ~n27049 & ~n27051 ;
  assign n27053 = n27047 & n27052 ;
  assign n27054 = \m2_addr_i[21]_pad  & n13928 ;
  assign n27055 = n13921 & n27054 ;
  assign n27056 = \m0_addr_i[21]_pad  & n13928 ;
  assign n27057 = n13945 & n27056 ;
  assign n27058 = ~n27055 & ~n27057 ;
  assign n27059 = \m6_addr_i[21]_pad  & n13928 ;
  assign n27060 = n13936 & n27059 ;
  assign n27061 = \m5_addr_i[21]_pad  & ~n13928 ;
  assign n27062 = n13953 & n27061 ;
  assign n27063 = ~n27060 & ~n27062 ;
  assign n27064 = n27058 & n27063 ;
  assign n27065 = n27053 & n27064 ;
  assign n27066 = \m1_addr_i[22]_pad  & ~n13928 ;
  assign n27067 = n13945 & n27066 ;
  assign n27068 = \m2_addr_i[22]_pad  & n13928 ;
  assign n27069 = n13921 & n27068 ;
  assign n27070 = ~n27067 & ~n27069 ;
  assign n27071 = \m0_addr_i[22]_pad  & n13928 ;
  assign n27072 = n13945 & n27071 ;
  assign n27073 = \m4_addr_i[22]_pad  & n13928 ;
  assign n27074 = n13953 & n27073 ;
  assign n27075 = ~n27072 & ~n27074 ;
  assign n27076 = n27070 & n27075 ;
  assign n27077 = \m7_addr_i[22]_pad  & ~n13928 ;
  assign n27078 = n13936 & n27077 ;
  assign n27079 = \m3_addr_i[22]_pad  & ~n13928 ;
  assign n27080 = n13921 & n27079 ;
  assign n27081 = ~n27078 & ~n27080 ;
  assign n27082 = \m6_addr_i[22]_pad  & n13928 ;
  assign n27083 = n13936 & n27082 ;
  assign n27084 = \m5_addr_i[22]_pad  & ~n13928 ;
  assign n27085 = n13953 & n27084 ;
  assign n27086 = ~n27083 & ~n27085 ;
  assign n27087 = n27081 & n27086 ;
  assign n27088 = n27076 & n27087 ;
  assign n27089 = \m1_addr_i[23]_pad  & ~n13928 ;
  assign n27090 = n13945 & n27089 ;
  assign n27091 = \m2_addr_i[23]_pad  & n13928 ;
  assign n27092 = n13921 & n27091 ;
  assign n27093 = ~n27090 & ~n27092 ;
  assign n27094 = \m0_addr_i[23]_pad  & n13928 ;
  assign n27095 = n13945 & n27094 ;
  assign n27096 = \m4_addr_i[23]_pad  & n13928 ;
  assign n27097 = n13953 & n27096 ;
  assign n27098 = ~n27095 & ~n27097 ;
  assign n27099 = n27093 & n27098 ;
  assign n27100 = \m7_addr_i[23]_pad  & ~n13928 ;
  assign n27101 = n13936 & n27100 ;
  assign n27102 = \m3_addr_i[23]_pad  & ~n13928 ;
  assign n27103 = n13921 & n27102 ;
  assign n27104 = ~n27101 & ~n27103 ;
  assign n27105 = \m6_addr_i[23]_pad  & n13928 ;
  assign n27106 = n13936 & n27105 ;
  assign n27107 = \m5_addr_i[23]_pad  & ~n13928 ;
  assign n27108 = n13953 & n27107 ;
  assign n27109 = ~n27106 & ~n27108 ;
  assign n27110 = n27104 & n27109 ;
  assign n27111 = n27099 & n27110 ;
  assign n27112 = \m3_addr_i[24]_pad  & ~n13928 ;
  assign n27113 = n13921 & n27112 ;
  assign n27114 = \m4_addr_i[24]_pad  & n13928 ;
  assign n27115 = n13953 & n27114 ;
  assign n27116 = ~n27113 & ~n27115 ;
  assign n27117 = \m5_addr_i[24]_pad  & ~n13928 ;
  assign n27118 = n13953 & n27117 ;
  assign n27119 = \m7_addr_i[24]_pad  & ~n13928 ;
  assign n27120 = n13936 & n27119 ;
  assign n27121 = ~n27118 & ~n27120 ;
  assign n27122 = n27116 & n27121 ;
  assign n27123 = \m6_addr_i[24]_pad  & n13928 ;
  assign n27124 = n13936 & n27123 ;
  assign n27125 = \m0_addr_i[24]_pad  & n13928 ;
  assign n27126 = n13945 & n27125 ;
  assign n27127 = ~n27124 & ~n27126 ;
  assign n27128 = \m1_addr_i[24]_pad  & ~n13928 ;
  assign n27129 = n13945 & n27128 ;
  assign n27130 = \m2_addr_i[24]_pad  & n13928 ;
  assign n27131 = n13921 & n27130 ;
  assign n27132 = ~n27129 & ~n27131 ;
  assign n27133 = n27127 & n27132 ;
  assign n27134 = n27122 & n27133 ;
  assign n27135 = \m0_addr_i[25]_pad  & n13928 ;
  assign n27136 = n13945 & n27135 ;
  assign n27137 = \m7_addr_i[25]_pad  & ~n13928 ;
  assign n27138 = n13936 & n27137 ;
  assign n27139 = ~n27136 & ~n27138 ;
  assign n27140 = \m1_addr_i[25]_pad  & ~n13928 ;
  assign n27141 = n13945 & n27140 ;
  assign n27142 = \m4_addr_i[25]_pad  & n13928 ;
  assign n27143 = n13953 & n27142 ;
  assign n27144 = ~n27141 & ~n27143 ;
  assign n27145 = n27139 & n27144 ;
  assign n27146 = \m2_addr_i[25]_pad  & n13928 ;
  assign n27147 = n13921 & n27146 ;
  assign n27148 = \m3_addr_i[25]_pad  & ~n13928 ;
  assign n27149 = n13921 & n27148 ;
  assign n27150 = ~n27147 & ~n27149 ;
  assign n27151 = \m5_addr_i[25]_pad  & ~n13928 ;
  assign n27152 = n13953 & n27151 ;
  assign n27153 = \m6_addr_i[25]_pad  & n13928 ;
  assign n27154 = n13936 & n27153 ;
  assign n27155 = ~n27152 & ~n27154 ;
  assign n27156 = n27150 & n27155 ;
  assign n27157 = n27145 & n27156 ;
  assign n27158 = \m0_addr_i[26]_pad  & n13928 ;
  assign n27159 = n13945 & n27158 ;
  assign n27160 = \m7_addr_i[26]_pad  & ~n13928 ;
  assign n27161 = n13936 & n27160 ;
  assign n27162 = ~n27159 & ~n27161 ;
  assign n27163 = \m5_addr_i[26]_pad  & ~n13928 ;
  assign n27164 = n13953 & n27163 ;
  assign n27165 = \m2_addr_i[26]_pad  & n13928 ;
  assign n27166 = n13921 & n27165 ;
  assign n27167 = ~n27164 & ~n27166 ;
  assign n27168 = n27162 & n27167 ;
  assign n27169 = \m6_addr_i[26]_pad  & n13928 ;
  assign n27170 = n13936 & n27169 ;
  assign n27171 = \m1_addr_i[26]_pad  & ~n13928 ;
  assign n27172 = n13945 & n27171 ;
  assign n27173 = ~n27170 & ~n27172 ;
  assign n27174 = \m3_addr_i[26]_pad  & ~n13928 ;
  assign n27175 = n13921 & n27174 ;
  assign n27176 = \m4_addr_i[26]_pad  & n13928 ;
  assign n27177 = n13953 & n27176 ;
  assign n27178 = ~n27175 & ~n27177 ;
  assign n27179 = n27173 & n27178 ;
  assign n27180 = n27168 & n27179 ;
  assign n27181 = \m0_addr_i[27]_pad  & n13928 ;
  assign n27182 = n13945 & n27181 ;
  assign n27183 = \m7_addr_i[27]_pad  & ~n13928 ;
  assign n27184 = n13936 & n27183 ;
  assign n27185 = ~n27182 & ~n27184 ;
  assign n27186 = \m1_addr_i[27]_pad  & ~n13928 ;
  assign n27187 = n13945 & n27186 ;
  assign n27188 = \m4_addr_i[27]_pad  & n13928 ;
  assign n27189 = n13953 & n27188 ;
  assign n27190 = ~n27187 & ~n27189 ;
  assign n27191 = n27185 & n27190 ;
  assign n27192 = \m2_addr_i[27]_pad  & n13928 ;
  assign n27193 = n13921 & n27192 ;
  assign n27194 = \m3_addr_i[27]_pad  & ~n13928 ;
  assign n27195 = n13921 & n27194 ;
  assign n27196 = ~n27193 & ~n27195 ;
  assign n27197 = \m5_addr_i[27]_pad  & ~n13928 ;
  assign n27198 = n13953 & n27197 ;
  assign n27199 = \m6_addr_i[27]_pad  & n13928 ;
  assign n27200 = n13936 & n27199 ;
  assign n27201 = ~n27198 & ~n27200 ;
  assign n27202 = n27196 & n27201 ;
  assign n27203 = n27191 & n27202 ;
  assign n27204 = \m3_addr_i[28]_pad  & ~n13928 ;
  assign n27205 = n13921 & n27204 ;
  assign n27206 = \m4_addr_i[28]_pad  & n13928 ;
  assign n27207 = n13953 & n27206 ;
  assign n27208 = ~n27205 & ~n27207 ;
  assign n27209 = \m5_addr_i[28]_pad  & ~n13928 ;
  assign n27210 = n13953 & n27209 ;
  assign n27211 = \m7_addr_i[28]_pad  & ~n13928 ;
  assign n27212 = n13936 & n27211 ;
  assign n27213 = ~n27210 & ~n27212 ;
  assign n27214 = n27208 & n27213 ;
  assign n27215 = \m6_addr_i[28]_pad  & n13928 ;
  assign n27216 = n13936 & n27215 ;
  assign n27217 = \m0_addr_i[28]_pad  & n13928 ;
  assign n27218 = n13945 & n27217 ;
  assign n27219 = ~n27216 & ~n27218 ;
  assign n27220 = \m1_addr_i[28]_pad  & ~n13928 ;
  assign n27221 = n13945 & n27220 ;
  assign n27222 = \m2_addr_i[28]_pad  & n13928 ;
  assign n27223 = n13921 & n27222 ;
  assign n27224 = ~n27221 & ~n27223 ;
  assign n27225 = n27219 & n27224 ;
  assign n27226 = n27214 & n27225 ;
  assign n27227 = \m0_addr_i[29]_pad  & n13928 ;
  assign n27228 = n13945 & n27227 ;
  assign n27229 = \m7_addr_i[29]_pad  & ~n13928 ;
  assign n27230 = n13936 & n27229 ;
  assign n27231 = ~n27228 & ~n27230 ;
  assign n27232 = \m1_addr_i[29]_pad  & ~n13928 ;
  assign n27233 = n13945 & n27232 ;
  assign n27234 = \m4_addr_i[29]_pad  & n13928 ;
  assign n27235 = n13953 & n27234 ;
  assign n27236 = ~n27233 & ~n27235 ;
  assign n27237 = n27231 & n27236 ;
  assign n27238 = \m2_addr_i[29]_pad  & n13928 ;
  assign n27239 = n13921 & n27238 ;
  assign n27240 = \m3_addr_i[29]_pad  & ~n13928 ;
  assign n27241 = n13921 & n27240 ;
  assign n27242 = ~n27239 & ~n27241 ;
  assign n27243 = \m5_addr_i[29]_pad  & ~n13928 ;
  assign n27244 = n13953 & n27243 ;
  assign n27245 = \m6_addr_i[29]_pad  & n13928 ;
  assign n27246 = n13936 & n27245 ;
  assign n27247 = ~n27244 & ~n27246 ;
  assign n27248 = n27242 & n27247 ;
  assign n27249 = n27237 & n27248 ;
  assign n27250 = \m0_addr_i[2]_pad  & n13928 ;
  assign n27251 = n13945 & n27250 ;
  assign n27252 = \m7_addr_i[2]_pad  & ~n13928 ;
  assign n27253 = n13936 & n27252 ;
  assign n27254 = ~n27251 & ~n27253 ;
  assign n27255 = \m6_addr_i[2]_pad  & n13928 ;
  assign n27256 = n13936 & n27255 ;
  assign n27257 = \m2_addr_i[2]_pad  & n13928 ;
  assign n27258 = n13921 & n27257 ;
  assign n27259 = ~n27256 & ~n27258 ;
  assign n27260 = n27254 & n27259 ;
  assign n27261 = \m5_addr_i[2]_pad  & ~n13928 ;
  assign n27262 = n13953 & n27261 ;
  assign n27263 = \m1_addr_i[2]_pad  & ~n13928 ;
  assign n27264 = n13945 & n27263 ;
  assign n27265 = ~n27262 & ~n27264 ;
  assign n27266 = \m3_addr_i[2]_pad  & ~n13928 ;
  assign n27267 = n13921 & n27266 ;
  assign n27268 = \m4_addr_i[2]_pad  & n13928 ;
  assign n27269 = n13953 & n27268 ;
  assign n27270 = ~n27267 & ~n27269 ;
  assign n27271 = n27265 & n27270 ;
  assign n27272 = n27260 & n27271 ;
  assign n27273 = \m1_addr_i[30]_pad  & ~n13928 ;
  assign n27274 = n13945 & n27273 ;
  assign n27275 = \m2_addr_i[30]_pad  & n13928 ;
  assign n27276 = n13921 & n27275 ;
  assign n27277 = ~n27274 & ~n27276 ;
  assign n27278 = \m3_addr_i[30]_pad  & ~n13928 ;
  assign n27279 = n13921 & n27278 ;
  assign n27280 = \m6_addr_i[30]_pad  & n13928 ;
  assign n27281 = n13936 & n27280 ;
  assign n27282 = ~n27279 & ~n27281 ;
  assign n27283 = n27277 & n27282 ;
  assign n27284 = \m4_addr_i[30]_pad  & n13928 ;
  assign n27285 = n13953 & n27284 ;
  assign n27286 = \m5_addr_i[30]_pad  & ~n13928 ;
  assign n27287 = n13953 & n27286 ;
  assign n27288 = ~n27285 & ~n27287 ;
  assign n27289 = \m0_addr_i[30]_pad  & n13928 ;
  assign n27290 = n13945 & n27289 ;
  assign n27291 = \m7_addr_i[30]_pad  & ~n13928 ;
  assign n27292 = n13936 & n27291 ;
  assign n27293 = ~n27290 & ~n27292 ;
  assign n27294 = n27288 & n27293 ;
  assign n27295 = n27283 & n27294 ;
  assign n27296 = \m5_addr_i[31]_pad  & ~n13928 ;
  assign n27297 = n13953 & n27296 ;
  assign n27298 = \m6_addr_i[31]_pad  & n13928 ;
  assign n27299 = n13936 & n27298 ;
  assign n27300 = ~n27297 & ~n27299 ;
  assign n27301 = \m0_addr_i[31]_pad  & n13928 ;
  assign n27302 = n13945 & n27301 ;
  assign n27303 = \m4_addr_i[31]_pad  & n13928 ;
  assign n27304 = n13953 & n27303 ;
  assign n27305 = ~n27302 & ~n27304 ;
  assign n27306 = n27300 & n27305 ;
  assign n27307 = \m7_addr_i[31]_pad  & ~n13928 ;
  assign n27308 = n13936 & n27307 ;
  assign n27309 = \m3_addr_i[31]_pad  & ~n13928 ;
  assign n27310 = n13921 & n27309 ;
  assign n27311 = ~n27308 & ~n27310 ;
  assign n27312 = \m1_addr_i[31]_pad  & ~n13928 ;
  assign n27313 = n13945 & n27312 ;
  assign n27314 = \m2_addr_i[31]_pad  & n13928 ;
  assign n27315 = n13921 & n27314 ;
  assign n27316 = ~n27313 & ~n27315 ;
  assign n27317 = n27311 & n27316 ;
  assign n27318 = n27306 & n27317 ;
  assign n27319 = \m6_addr_i[3]_pad  & n13928 ;
  assign n27320 = n13936 & n27319 ;
  assign n27321 = \m5_addr_i[3]_pad  & ~n13928 ;
  assign n27322 = n13953 & n27321 ;
  assign n27323 = ~n27320 & ~n27322 ;
  assign n27324 = \m0_addr_i[3]_pad  & n13928 ;
  assign n27325 = n13945 & n27324 ;
  assign n27326 = \m2_addr_i[3]_pad  & n13928 ;
  assign n27327 = n13921 & n27326 ;
  assign n27328 = ~n27325 & ~n27327 ;
  assign n27329 = n27323 & n27328 ;
  assign n27330 = \m7_addr_i[3]_pad  & ~n13928 ;
  assign n27331 = n13936 & n27330 ;
  assign n27332 = \m1_addr_i[3]_pad  & ~n13928 ;
  assign n27333 = n13945 & n27332 ;
  assign n27334 = ~n27331 & ~n27333 ;
  assign n27335 = \m3_addr_i[3]_pad  & ~n13928 ;
  assign n27336 = n13921 & n27335 ;
  assign n27337 = \m4_addr_i[3]_pad  & n13928 ;
  assign n27338 = n13953 & n27337 ;
  assign n27339 = ~n27336 & ~n27338 ;
  assign n27340 = n27334 & n27339 ;
  assign n27341 = n27329 & n27340 ;
  assign n27342 = \m1_addr_i[4]_pad  & ~n13928 ;
  assign n27343 = n13945 & n27342 ;
  assign n27344 = \m2_addr_i[4]_pad  & n13928 ;
  assign n27345 = n13921 & n27344 ;
  assign n27346 = ~n27343 & ~n27345 ;
  assign n27347 = \m0_addr_i[4]_pad  & n13928 ;
  assign n27348 = n13945 & n27347 ;
  assign n27349 = \m4_addr_i[4]_pad  & n13928 ;
  assign n27350 = n13953 & n27349 ;
  assign n27351 = ~n27348 & ~n27350 ;
  assign n27352 = n27346 & n27351 ;
  assign n27353 = \m7_addr_i[4]_pad  & ~n13928 ;
  assign n27354 = n13936 & n27353 ;
  assign n27355 = \m3_addr_i[4]_pad  & ~n13928 ;
  assign n27356 = n13921 & n27355 ;
  assign n27357 = ~n27354 & ~n27356 ;
  assign n27358 = \m6_addr_i[4]_pad  & n13928 ;
  assign n27359 = n13936 & n27358 ;
  assign n27360 = \m5_addr_i[4]_pad  & ~n13928 ;
  assign n27361 = n13953 & n27360 ;
  assign n27362 = ~n27359 & ~n27361 ;
  assign n27363 = n27357 & n27362 ;
  assign n27364 = n27352 & n27363 ;
  assign n27365 = \m1_addr_i[5]_pad  & ~n13928 ;
  assign n27366 = n13945 & n27365 ;
  assign n27367 = \m2_addr_i[5]_pad  & n13928 ;
  assign n27368 = n13921 & n27367 ;
  assign n27369 = ~n27366 & ~n27368 ;
  assign n27370 = \m0_addr_i[5]_pad  & n13928 ;
  assign n27371 = n13945 & n27370 ;
  assign n27372 = \m4_addr_i[5]_pad  & n13928 ;
  assign n27373 = n13953 & n27372 ;
  assign n27374 = ~n27371 & ~n27373 ;
  assign n27375 = n27369 & n27374 ;
  assign n27376 = \m7_addr_i[5]_pad  & ~n13928 ;
  assign n27377 = n13936 & n27376 ;
  assign n27378 = \m3_addr_i[5]_pad  & ~n13928 ;
  assign n27379 = n13921 & n27378 ;
  assign n27380 = ~n27377 & ~n27379 ;
  assign n27381 = \m6_addr_i[5]_pad  & n13928 ;
  assign n27382 = n13936 & n27381 ;
  assign n27383 = \m5_addr_i[5]_pad  & ~n13928 ;
  assign n27384 = n13953 & n27383 ;
  assign n27385 = ~n27382 & ~n27384 ;
  assign n27386 = n27380 & n27385 ;
  assign n27387 = n27375 & n27386 ;
  assign n27388 = \m0_addr_i[6]_pad  & n13928 ;
  assign n27389 = n13945 & n27388 ;
  assign n27390 = \m7_addr_i[6]_pad  & ~n13928 ;
  assign n27391 = n13936 & n27390 ;
  assign n27392 = ~n27389 & ~n27391 ;
  assign n27393 = \m3_addr_i[6]_pad  & ~n13928 ;
  assign n27394 = n13921 & n27393 ;
  assign n27395 = \m2_addr_i[6]_pad  & n13928 ;
  assign n27396 = n13921 & n27395 ;
  assign n27397 = ~n27394 & ~n27396 ;
  assign n27398 = n27392 & n27397 ;
  assign n27399 = \m4_addr_i[6]_pad  & n13928 ;
  assign n27400 = n13953 & n27399 ;
  assign n27401 = \m1_addr_i[6]_pad  & ~n13928 ;
  assign n27402 = n13945 & n27401 ;
  assign n27403 = ~n27400 & ~n27402 ;
  assign n27404 = \m6_addr_i[6]_pad  & n13928 ;
  assign n27405 = n13936 & n27404 ;
  assign n27406 = \m5_addr_i[6]_pad  & ~n13928 ;
  assign n27407 = n13953 & n27406 ;
  assign n27408 = ~n27405 & ~n27407 ;
  assign n27409 = n27403 & n27408 ;
  assign n27410 = n27398 & n27409 ;
  assign n27411 = \m0_addr_i[7]_pad  & n13928 ;
  assign n27412 = n13945 & n27411 ;
  assign n27413 = \m7_addr_i[7]_pad  & ~n13928 ;
  assign n27414 = n13936 & n27413 ;
  assign n27415 = ~n27412 & ~n27414 ;
  assign n27416 = \m1_addr_i[7]_pad  & ~n13928 ;
  assign n27417 = n13945 & n27416 ;
  assign n27418 = \m5_addr_i[7]_pad  & ~n13928 ;
  assign n27419 = n13953 & n27418 ;
  assign n27420 = ~n27417 & ~n27419 ;
  assign n27421 = n27415 & n27420 ;
  assign n27422 = \m2_addr_i[7]_pad  & n13928 ;
  assign n27423 = n13921 & n27422 ;
  assign n27424 = \m6_addr_i[7]_pad  & n13928 ;
  assign n27425 = n13936 & n27424 ;
  assign n27426 = ~n27423 & ~n27425 ;
  assign n27427 = \m3_addr_i[7]_pad  & ~n13928 ;
  assign n27428 = n13921 & n27427 ;
  assign n27429 = \m4_addr_i[7]_pad  & n13928 ;
  assign n27430 = n13953 & n27429 ;
  assign n27431 = ~n27428 & ~n27430 ;
  assign n27432 = n27426 & n27431 ;
  assign n27433 = n27421 & n27432 ;
  assign n27434 = \m0_addr_i[8]_pad  & n13928 ;
  assign n27435 = n13945 & n27434 ;
  assign n27436 = \m7_addr_i[8]_pad  & ~n13928 ;
  assign n27437 = n13936 & n27436 ;
  assign n27438 = ~n27435 & ~n27437 ;
  assign n27439 = \m6_addr_i[8]_pad  & n13928 ;
  assign n27440 = n13936 & n27439 ;
  assign n27441 = \m2_addr_i[8]_pad  & n13928 ;
  assign n27442 = n13921 & n27441 ;
  assign n27443 = ~n27440 & ~n27442 ;
  assign n27444 = n27438 & n27443 ;
  assign n27445 = \m5_addr_i[8]_pad  & ~n13928 ;
  assign n27446 = n13953 & n27445 ;
  assign n27447 = \m1_addr_i[8]_pad  & ~n13928 ;
  assign n27448 = n13945 & n27447 ;
  assign n27449 = ~n27446 & ~n27448 ;
  assign n27450 = \m3_addr_i[8]_pad  & ~n13928 ;
  assign n27451 = n13921 & n27450 ;
  assign n27452 = \m4_addr_i[8]_pad  & n13928 ;
  assign n27453 = n13953 & n27452 ;
  assign n27454 = ~n27451 & ~n27453 ;
  assign n27455 = n27449 & n27454 ;
  assign n27456 = n27444 & n27455 ;
  assign n27457 = \m1_addr_i[9]_pad  & ~n13928 ;
  assign n27458 = n13945 & n27457 ;
  assign n27459 = \m2_addr_i[9]_pad  & n13928 ;
  assign n27460 = n13921 & n27459 ;
  assign n27461 = ~n27458 & ~n27460 ;
  assign n27462 = \m6_addr_i[9]_pad  & n13928 ;
  assign n27463 = n13936 & n27462 ;
  assign n27464 = \m7_addr_i[9]_pad  & ~n13928 ;
  assign n27465 = n13936 & n27464 ;
  assign n27466 = ~n27463 & ~n27465 ;
  assign n27467 = n27461 & n27466 ;
  assign n27468 = \m5_addr_i[9]_pad  & ~n13928 ;
  assign n27469 = n13953 & n27468 ;
  assign n27470 = \m0_addr_i[9]_pad  & n13928 ;
  assign n27471 = n13945 & n27470 ;
  assign n27472 = ~n27469 & ~n27471 ;
  assign n27473 = \m3_addr_i[9]_pad  & ~n13928 ;
  assign n27474 = n13921 & n27473 ;
  assign n27475 = \m4_addr_i[9]_pad  & n13928 ;
  assign n27476 = n13953 & n27475 ;
  assign n27477 = ~n27474 & ~n27476 ;
  assign n27478 = n27472 & n27477 ;
  assign n27479 = n27467 & n27478 ;
  assign n27480 = \m3_data_i[0]_pad  & ~n13928 ;
  assign n27481 = n13921 & n27480 ;
  assign n27482 = \m4_data_i[0]_pad  & n13928 ;
  assign n27483 = n13953 & n27482 ;
  assign n27484 = ~n27481 & ~n27483 ;
  assign n27485 = \m1_data_i[0]_pad  & ~n13928 ;
  assign n27486 = n13945 & n27485 ;
  assign n27487 = \m5_data_i[0]_pad  & ~n13928 ;
  assign n27488 = n13953 & n27487 ;
  assign n27489 = ~n27486 & ~n27488 ;
  assign n27490 = n27484 & n27489 ;
  assign n27491 = \m2_data_i[0]_pad  & n13928 ;
  assign n27492 = n13921 & n27491 ;
  assign n27493 = \m6_data_i[0]_pad  & n13928 ;
  assign n27494 = n13936 & n27493 ;
  assign n27495 = ~n27492 & ~n27494 ;
  assign n27496 = \m0_data_i[0]_pad  & n13928 ;
  assign n27497 = n13945 & n27496 ;
  assign n27498 = \m7_data_i[0]_pad  & ~n13928 ;
  assign n27499 = n13936 & n27498 ;
  assign n27500 = ~n27497 & ~n27499 ;
  assign n27501 = n27495 & n27500 ;
  assign n27502 = n27490 & n27501 ;
  assign n27503 = \m0_data_i[10]_pad  & n13928 ;
  assign n27504 = n13945 & n27503 ;
  assign n27505 = \m7_data_i[10]_pad  & ~n13928 ;
  assign n27506 = n13936 & n27505 ;
  assign n27507 = ~n27504 & ~n27506 ;
  assign n27508 = \m1_data_i[10]_pad  & ~n13928 ;
  assign n27509 = n13945 & n27508 ;
  assign n27510 = \m4_data_i[10]_pad  & n13928 ;
  assign n27511 = n13953 & n27510 ;
  assign n27512 = ~n27509 & ~n27511 ;
  assign n27513 = n27507 & n27512 ;
  assign n27514 = \m2_data_i[10]_pad  & n13928 ;
  assign n27515 = n13921 & n27514 ;
  assign n27516 = \m3_data_i[10]_pad  & ~n13928 ;
  assign n27517 = n13921 & n27516 ;
  assign n27518 = ~n27515 & ~n27517 ;
  assign n27519 = \m6_data_i[10]_pad  & n13928 ;
  assign n27520 = n13936 & n27519 ;
  assign n27521 = \m5_data_i[10]_pad  & ~n13928 ;
  assign n27522 = n13953 & n27521 ;
  assign n27523 = ~n27520 & ~n27522 ;
  assign n27524 = n27518 & n27523 ;
  assign n27525 = n27513 & n27524 ;
  assign n27526 = \m1_data_i[11]_pad  & ~n13928 ;
  assign n27527 = n13945 & n27526 ;
  assign n27528 = \m2_data_i[11]_pad  & n13928 ;
  assign n27529 = n13921 & n27528 ;
  assign n27530 = ~n27527 & ~n27529 ;
  assign n27531 = \m0_data_i[11]_pad  & n13928 ;
  assign n27532 = n13945 & n27531 ;
  assign n27533 = \m4_data_i[11]_pad  & n13928 ;
  assign n27534 = n13953 & n27533 ;
  assign n27535 = ~n27532 & ~n27534 ;
  assign n27536 = n27530 & n27535 ;
  assign n27537 = \m7_data_i[11]_pad  & ~n13928 ;
  assign n27538 = n13936 & n27537 ;
  assign n27539 = \m3_data_i[11]_pad  & ~n13928 ;
  assign n27540 = n13921 & n27539 ;
  assign n27541 = ~n27538 & ~n27540 ;
  assign n27542 = \m6_data_i[11]_pad  & n13928 ;
  assign n27543 = n13936 & n27542 ;
  assign n27544 = \m5_data_i[11]_pad  & ~n13928 ;
  assign n27545 = n13953 & n27544 ;
  assign n27546 = ~n27543 & ~n27545 ;
  assign n27547 = n27541 & n27546 ;
  assign n27548 = n27536 & n27547 ;
  assign n27549 = \m1_data_i[12]_pad  & ~n13928 ;
  assign n27550 = n13945 & n27549 ;
  assign n27551 = \m2_data_i[12]_pad  & n13928 ;
  assign n27552 = n13921 & n27551 ;
  assign n27553 = ~n27550 & ~n27552 ;
  assign n27554 = \m0_data_i[12]_pad  & n13928 ;
  assign n27555 = n13945 & n27554 ;
  assign n27556 = \m4_data_i[12]_pad  & n13928 ;
  assign n27557 = n13953 & n27556 ;
  assign n27558 = ~n27555 & ~n27557 ;
  assign n27559 = n27553 & n27558 ;
  assign n27560 = \m7_data_i[12]_pad  & ~n13928 ;
  assign n27561 = n13936 & n27560 ;
  assign n27562 = \m3_data_i[12]_pad  & ~n13928 ;
  assign n27563 = n13921 & n27562 ;
  assign n27564 = ~n27561 & ~n27563 ;
  assign n27565 = \m6_data_i[12]_pad  & n13928 ;
  assign n27566 = n13936 & n27565 ;
  assign n27567 = \m5_data_i[12]_pad  & ~n13928 ;
  assign n27568 = n13953 & n27567 ;
  assign n27569 = ~n27566 & ~n27568 ;
  assign n27570 = n27564 & n27569 ;
  assign n27571 = n27559 & n27570 ;
  assign n27572 = \m0_data_i[13]_pad  & n13928 ;
  assign n27573 = n13945 & n27572 ;
  assign n27574 = \m7_data_i[13]_pad  & ~n13928 ;
  assign n27575 = n13936 & n27574 ;
  assign n27576 = ~n27573 & ~n27575 ;
  assign n27577 = \m6_data_i[13]_pad  & n13928 ;
  assign n27578 = n13936 & n27577 ;
  assign n27579 = \m2_data_i[13]_pad  & n13928 ;
  assign n27580 = n13921 & n27579 ;
  assign n27581 = ~n27578 & ~n27580 ;
  assign n27582 = n27576 & n27581 ;
  assign n27583 = \m5_data_i[13]_pad  & ~n13928 ;
  assign n27584 = n13953 & n27583 ;
  assign n27585 = \m1_data_i[13]_pad  & ~n13928 ;
  assign n27586 = n13945 & n27585 ;
  assign n27587 = ~n27584 & ~n27586 ;
  assign n27588 = \m3_data_i[13]_pad  & ~n13928 ;
  assign n27589 = n13921 & n27588 ;
  assign n27590 = \m4_data_i[13]_pad  & n13928 ;
  assign n27591 = n13953 & n27590 ;
  assign n27592 = ~n27589 & ~n27591 ;
  assign n27593 = n27587 & n27592 ;
  assign n27594 = n27582 & n27593 ;
  assign n27595 = \m6_data_i[14]_pad  & n13928 ;
  assign n27596 = n13936 & n27595 ;
  assign n27597 = \m5_data_i[14]_pad  & ~n13928 ;
  assign n27598 = n13953 & n27597 ;
  assign n27599 = ~n27596 & ~n27598 ;
  assign n27600 = \m3_data_i[14]_pad  & ~n13928 ;
  assign n27601 = n13921 & n27600 ;
  assign n27602 = \m2_data_i[14]_pad  & n13928 ;
  assign n27603 = n13921 & n27602 ;
  assign n27604 = ~n27601 & ~n27603 ;
  assign n27605 = n27599 & n27604 ;
  assign n27606 = \m4_data_i[14]_pad  & n13928 ;
  assign n27607 = n13953 & n27606 ;
  assign n27608 = \m1_data_i[14]_pad  & ~n13928 ;
  assign n27609 = n13945 & n27608 ;
  assign n27610 = ~n27607 & ~n27609 ;
  assign n27611 = \m0_data_i[14]_pad  & n13928 ;
  assign n27612 = n13945 & n27611 ;
  assign n27613 = \m7_data_i[14]_pad  & ~n13928 ;
  assign n27614 = n13936 & n27613 ;
  assign n27615 = ~n27612 & ~n27614 ;
  assign n27616 = n27610 & n27615 ;
  assign n27617 = n27605 & n27616 ;
  assign n27618 = \m3_data_i[15]_pad  & ~n13928 ;
  assign n27619 = n13921 & n27618 ;
  assign n27620 = \m4_data_i[15]_pad  & n13928 ;
  assign n27621 = n13953 & n27620 ;
  assign n27622 = ~n27619 & ~n27621 ;
  assign n27623 = \m1_data_i[15]_pad  & ~n13928 ;
  assign n27624 = n13945 & n27623 ;
  assign n27625 = \m5_data_i[15]_pad  & ~n13928 ;
  assign n27626 = n13953 & n27625 ;
  assign n27627 = ~n27624 & ~n27626 ;
  assign n27628 = n27622 & n27627 ;
  assign n27629 = \m2_data_i[15]_pad  & n13928 ;
  assign n27630 = n13921 & n27629 ;
  assign n27631 = \m6_data_i[15]_pad  & n13928 ;
  assign n27632 = n13936 & n27631 ;
  assign n27633 = ~n27630 & ~n27632 ;
  assign n27634 = \m0_data_i[15]_pad  & n13928 ;
  assign n27635 = n13945 & n27634 ;
  assign n27636 = \m7_data_i[15]_pad  & ~n13928 ;
  assign n27637 = n13936 & n27636 ;
  assign n27638 = ~n27635 & ~n27637 ;
  assign n27639 = n27633 & n27638 ;
  assign n27640 = n27628 & n27639 ;
  assign n27641 = \m3_data_i[16]_pad  & ~n13928 ;
  assign n27642 = n13921 & n27641 ;
  assign n27643 = \m4_data_i[16]_pad  & n13928 ;
  assign n27644 = n13953 & n27643 ;
  assign n27645 = ~n27642 & ~n27644 ;
  assign n27646 = \m1_data_i[16]_pad  & ~n13928 ;
  assign n27647 = n13945 & n27646 ;
  assign n27648 = \m5_data_i[16]_pad  & ~n13928 ;
  assign n27649 = n13953 & n27648 ;
  assign n27650 = ~n27647 & ~n27649 ;
  assign n27651 = n27645 & n27650 ;
  assign n27652 = \m2_data_i[16]_pad  & n13928 ;
  assign n27653 = n13921 & n27652 ;
  assign n27654 = \m6_data_i[16]_pad  & n13928 ;
  assign n27655 = n13936 & n27654 ;
  assign n27656 = ~n27653 & ~n27655 ;
  assign n27657 = \m0_data_i[16]_pad  & n13928 ;
  assign n27658 = n13945 & n27657 ;
  assign n27659 = \m7_data_i[16]_pad  & ~n13928 ;
  assign n27660 = n13936 & n27659 ;
  assign n27661 = ~n27658 & ~n27660 ;
  assign n27662 = n27656 & n27661 ;
  assign n27663 = n27651 & n27662 ;
  assign n27664 = \m6_data_i[17]_pad  & n13928 ;
  assign n27665 = n13936 & n27664 ;
  assign n27666 = \m5_data_i[17]_pad  & ~n13928 ;
  assign n27667 = n13953 & n27666 ;
  assign n27668 = ~n27665 & ~n27667 ;
  assign n27669 = \m1_data_i[17]_pad  & ~n13928 ;
  assign n27670 = n13945 & n27669 ;
  assign n27671 = \m4_data_i[17]_pad  & n13928 ;
  assign n27672 = n13953 & n27671 ;
  assign n27673 = ~n27670 & ~n27672 ;
  assign n27674 = n27668 & n27673 ;
  assign n27675 = \m2_data_i[17]_pad  & n13928 ;
  assign n27676 = n13921 & n27675 ;
  assign n27677 = \m3_data_i[17]_pad  & ~n13928 ;
  assign n27678 = n13921 & n27677 ;
  assign n27679 = ~n27676 & ~n27678 ;
  assign n27680 = \m0_data_i[17]_pad  & n13928 ;
  assign n27681 = n13945 & n27680 ;
  assign n27682 = \m7_data_i[17]_pad  & ~n13928 ;
  assign n27683 = n13936 & n27682 ;
  assign n27684 = ~n27681 & ~n27683 ;
  assign n27685 = n27679 & n27684 ;
  assign n27686 = n27674 & n27685 ;
  assign n27687 = \m0_data_i[18]_pad  & n13928 ;
  assign n27688 = n13945 & n27687 ;
  assign n27689 = \m7_data_i[18]_pad  & ~n13928 ;
  assign n27690 = n13936 & n27689 ;
  assign n27691 = ~n27688 & ~n27690 ;
  assign n27692 = \m1_data_i[18]_pad  & ~n13928 ;
  assign n27693 = n13945 & n27692 ;
  assign n27694 = \m4_data_i[18]_pad  & n13928 ;
  assign n27695 = n13953 & n27694 ;
  assign n27696 = ~n27693 & ~n27695 ;
  assign n27697 = n27691 & n27696 ;
  assign n27698 = \m2_data_i[18]_pad  & n13928 ;
  assign n27699 = n13921 & n27698 ;
  assign n27700 = \m3_data_i[18]_pad  & ~n13928 ;
  assign n27701 = n13921 & n27700 ;
  assign n27702 = ~n27699 & ~n27701 ;
  assign n27703 = \m6_data_i[18]_pad  & n13928 ;
  assign n27704 = n13936 & n27703 ;
  assign n27705 = \m5_data_i[18]_pad  & ~n13928 ;
  assign n27706 = n13953 & n27705 ;
  assign n27707 = ~n27704 & ~n27706 ;
  assign n27708 = n27702 & n27707 ;
  assign n27709 = n27697 & n27708 ;
  assign n27710 = \m1_data_i[19]_pad  & ~n13928 ;
  assign n27711 = n13945 & n27710 ;
  assign n27712 = \m2_data_i[19]_pad  & n13928 ;
  assign n27713 = n13921 & n27712 ;
  assign n27714 = ~n27711 & ~n27713 ;
  assign n27715 = \m6_data_i[19]_pad  & n13928 ;
  assign n27716 = n13936 & n27715 ;
  assign n27717 = \m4_data_i[19]_pad  & n13928 ;
  assign n27718 = n13953 & n27717 ;
  assign n27719 = ~n27716 & ~n27718 ;
  assign n27720 = n27714 & n27719 ;
  assign n27721 = \m5_data_i[19]_pad  & ~n13928 ;
  assign n27722 = n13953 & n27721 ;
  assign n27723 = \m3_data_i[19]_pad  & ~n13928 ;
  assign n27724 = n13921 & n27723 ;
  assign n27725 = ~n27722 & ~n27724 ;
  assign n27726 = \m0_data_i[19]_pad  & n13928 ;
  assign n27727 = n13945 & n27726 ;
  assign n27728 = \m7_data_i[19]_pad  & ~n13928 ;
  assign n27729 = n13936 & n27728 ;
  assign n27730 = ~n27727 & ~n27729 ;
  assign n27731 = n27725 & n27730 ;
  assign n27732 = n27720 & n27731 ;
  assign n27733 = \m3_data_i[1]_pad  & ~n13928 ;
  assign n27734 = n13921 & n27733 ;
  assign n27735 = \m4_data_i[1]_pad  & n13928 ;
  assign n27736 = n13953 & n27735 ;
  assign n27737 = ~n27734 & ~n27736 ;
  assign n27738 = \m1_data_i[1]_pad  & ~n13928 ;
  assign n27739 = n13945 & n27738 ;
  assign n27740 = \m5_data_i[1]_pad  & ~n13928 ;
  assign n27741 = n13953 & n27740 ;
  assign n27742 = ~n27739 & ~n27741 ;
  assign n27743 = n27737 & n27742 ;
  assign n27744 = \m2_data_i[1]_pad  & n13928 ;
  assign n27745 = n13921 & n27744 ;
  assign n27746 = \m6_data_i[1]_pad  & n13928 ;
  assign n27747 = n13936 & n27746 ;
  assign n27748 = ~n27745 & ~n27747 ;
  assign n27749 = \m0_data_i[1]_pad  & n13928 ;
  assign n27750 = n13945 & n27749 ;
  assign n27751 = \m7_data_i[1]_pad  & ~n13928 ;
  assign n27752 = n13936 & n27751 ;
  assign n27753 = ~n27750 & ~n27752 ;
  assign n27754 = n27748 & n27753 ;
  assign n27755 = n27743 & n27754 ;
  assign n27756 = \m0_data_i[20]_pad  & n13928 ;
  assign n27757 = n13945 & n27756 ;
  assign n27758 = \m7_data_i[20]_pad  & ~n13928 ;
  assign n27759 = n13936 & n27758 ;
  assign n27760 = ~n27757 & ~n27759 ;
  assign n27761 = \m1_data_i[20]_pad  & ~n13928 ;
  assign n27762 = n13945 & n27761 ;
  assign n27763 = \m4_data_i[20]_pad  & n13928 ;
  assign n27764 = n13953 & n27763 ;
  assign n27765 = ~n27762 & ~n27764 ;
  assign n27766 = n27760 & n27765 ;
  assign n27767 = \m2_data_i[20]_pad  & n13928 ;
  assign n27768 = n13921 & n27767 ;
  assign n27769 = \m3_data_i[20]_pad  & ~n13928 ;
  assign n27770 = n13921 & n27769 ;
  assign n27771 = ~n27768 & ~n27770 ;
  assign n27772 = \m6_data_i[20]_pad  & n13928 ;
  assign n27773 = n13936 & n27772 ;
  assign n27774 = \m5_data_i[20]_pad  & ~n13928 ;
  assign n27775 = n13953 & n27774 ;
  assign n27776 = ~n27773 & ~n27775 ;
  assign n27777 = n27771 & n27776 ;
  assign n27778 = n27766 & n27777 ;
  assign n27779 = \m1_data_i[21]_pad  & ~n13928 ;
  assign n27780 = n13945 & n27779 ;
  assign n27781 = \m2_data_i[21]_pad  & n13928 ;
  assign n27782 = n13921 & n27781 ;
  assign n27783 = ~n27780 & ~n27782 ;
  assign n27784 = \m0_data_i[21]_pad  & n13928 ;
  assign n27785 = n13945 & n27784 ;
  assign n27786 = \m4_data_i[21]_pad  & n13928 ;
  assign n27787 = n13953 & n27786 ;
  assign n27788 = ~n27785 & ~n27787 ;
  assign n27789 = n27783 & n27788 ;
  assign n27790 = \m7_data_i[21]_pad  & ~n13928 ;
  assign n27791 = n13936 & n27790 ;
  assign n27792 = \m3_data_i[21]_pad  & ~n13928 ;
  assign n27793 = n13921 & n27792 ;
  assign n27794 = ~n27791 & ~n27793 ;
  assign n27795 = \m6_data_i[21]_pad  & n13928 ;
  assign n27796 = n13936 & n27795 ;
  assign n27797 = \m5_data_i[21]_pad  & ~n13928 ;
  assign n27798 = n13953 & n27797 ;
  assign n27799 = ~n27796 & ~n27798 ;
  assign n27800 = n27794 & n27799 ;
  assign n27801 = n27789 & n27800 ;
  assign n27802 = \m6_data_i[22]_pad  & n13928 ;
  assign n27803 = n13936 & n27802 ;
  assign n27804 = \m5_data_i[22]_pad  & ~n13928 ;
  assign n27805 = n13953 & n27804 ;
  assign n27806 = ~n27803 & ~n27805 ;
  assign n27807 = \m3_data_i[22]_pad  & ~n13928 ;
  assign n27808 = n13921 & n27807 ;
  assign n27809 = \m7_data_i[22]_pad  & ~n13928 ;
  assign n27810 = n13936 & n27809 ;
  assign n27811 = ~n27808 & ~n27810 ;
  assign n27812 = n27806 & n27811 ;
  assign n27813 = \m4_data_i[22]_pad  & n13928 ;
  assign n27814 = n13953 & n27813 ;
  assign n27815 = \m0_data_i[22]_pad  & n13928 ;
  assign n27816 = n13945 & n27815 ;
  assign n27817 = ~n27814 & ~n27816 ;
  assign n27818 = \m1_data_i[22]_pad  & ~n13928 ;
  assign n27819 = n13945 & n27818 ;
  assign n27820 = \m2_data_i[22]_pad  & n13928 ;
  assign n27821 = n13921 & n27820 ;
  assign n27822 = ~n27819 & ~n27821 ;
  assign n27823 = n27817 & n27822 ;
  assign n27824 = n27812 & n27823 ;
  assign n27825 = \m1_data_i[23]_pad  & ~n13928 ;
  assign n27826 = n13945 & n27825 ;
  assign n27827 = \m2_data_i[23]_pad  & n13928 ;
  assign n27828 = n13921 & n27827 ;
  assign n27829 = ~n27826 & ~n27828 ;
  assign n27830 = \m0_data_i[23]_pad  & n13928 ;
  assign n27831 = n13945 & n27830 ;
  assign n27832 = \m4_data_i[23]_pad  & n13928 ;
  assign n27833 = n13953 & n27832 ;
  assign n27834 = ~n27831 & ~n27833 ;
  assign n27835 = n27829 & n27834 ;
  assign n27836 = \m7_data_i[23]_pad  & ~n13928 ;
  assign n27837 = n13936 & n27836 ;
  assign n27838 = \m3_data_i[23]_pad  & ~n13928 ;
  assign n27839 = n13921 & n27838 ;
  assign n27840 = ~n27837 & ~n27839 ;
  assign n27841 = \m6_data_i[23]_pad  & n13928 ;
  assign n27842 = n13936 & n27841 ;
  assign n27843 = \m5_data_i[23]_pad  & ~n13928 ;
  assign n27844 = n13953 & n27843 ;
  assign n27845 = ~n27842 & ~n27844 ;
  assign n27846 = n27840 & n27845 ;
  assign n27847 = n27835 & n27846 ;
  assign n27848 = \m3_data_i[24]_pad  & ~n13928 ;
  assign n27849 = n13921 & n27848 ;
  assign n27850 = \m4_data_i[24]_pad  & n13928 ;
  assign n27851 = n13953 & n27850 ;
  assign n27852 = ~n27849 & ~n27851 ;
  assign n27853 = \m1_data_i[24]_pad  & ~n13928 ;
  assign n27854 = n13945 & n27853 ;
  assign n27855 = \m5_data_i[24]_pad  & ~n13928 ;
  assign n27856 = n13953 & n27855 ;
  assign n27857 = ~n27854 & ~n27856 ;
  assign n27858 = n27852 & n27857 ;
  assign n27859 = \m2_data_i[24]_pad  & n13928 ;
  assign n27860 = n13921 & n27859 ;
  assign n27861 = \m6_data_i[24]_pad  & n13928 ;
  assign n27862 = n13936 & n27861 ;
  assign n27863 = ~n27860 & ~n27862 ;
  assign n27864 = \m0_data_i[24]_pad  & n13928 ;
  assign n27865 = n13945 & n27864 ;
  assign n27866 = \m7_data_i[24]_pad  & ~n13928 ;
  assign n27867 = n13936 & n27866 ;
  assign n27868 = ~n27865 & ~n27867 ;
  assign n27869 = n27863 & n27868 ;
  assign n27870 = n27858 & n27869 ;
  assign n27871 = \m3_data_i[25]_pad  & ~n13928 ;
  assign n27872 = n13921 & n27871 ;
  assign n27873 = \m4_data_i[25]_pad  & n13928 ;
  assign n27874 = n13953 & n27873 ;
  assign n27875 = ~n27872 & ~n27874 ;
  assign n27876 = \m0_data_i[25]_pad  & n13928 ;
  assign n27877 = n13945 & n27876 ;
  assign n27878 = \m2_data_i[25]_pad  & n13928 ;
  assign n27879 = n13921 & n27878 ;
  assign n27880 = ~n27877 & ~n27879 ;
  assign n27881 = n27875 & n27880 ;
  assign n27882 = \m7_data_i[25]_pad  & ~n13928 ;
  assign n27883 = n13936 & n27882 ;
  assign n27884 = \m1_data_i[25]_pad  & ~n13928 ;
  assign n27885 = n13945 & n27884 ;
  assign n27886 = ~n27883 & ~n27885 ;
  assign n27887 = \m6_data_i[25]_pad  & n13928 ;
  assign n27888 = n13936 & n27887 ;
  assign n27889 = \m5_data_i[25]_pad  & ~n13928 ;
  assign n27890 = n13953 & n27889 ;
  assign n27891 = ~n27888 & ~n27890 ;
  assign n27892 = n27886 & n27891 ;
  assign n27893 = n27881 & n27892 ;
  assign n27894 = \m3_data_i[26]_pad  & ~n13928 ;
  assign n27895 = n13921 & n27894 ;
  assign n27896 = \m4_data_i[26]_pad  & n13928 ;
  assign n27897 = n13953 & n27896 ;
  assign n27898 = ~n27895 & ~n27897 ;
  assign n27899 = \m0_data_i[26]_pad  & n13928 ;
  assign n27900 = n13945 & n27899 ;
  assign n27901 = \m5_data_i[26]_pad  & ~n13928 ;
  assign n27902 = n13953 & n27901 ;
  assign n27903 = ~n27900 & ~n27902 ;
  assign n27904 = n27898 & n27903 ;
  assign n27905 = \m7_data_i[26]_pad  & ~n13928 ;
  assign n27906 = n13936 & n27905 ;
  assign n27907 = \m6_data_i[26]_pad  & n13928 ;
  assign n27908 = n13936 & n27907 ;
  assign n27909 = ~n27906 & ~n27908 ;
  assign n27910 = \m1_data_i[26]_pad  & ~n13928 ;
  assign n27911 = n13945 & n27910 ;
  assign n27912 = \m2_data_i[26]_pad  & n13928 ;
  assign n27913 = n13921 & n27912 ;
  assign n27914 = ~n27911 & ~n27913 ;
  assign n27915 = n27909 & n27914 ;
  assign n27916 = n27904 & n27915 ;
  assign n27917 = \m1_data_i[27]_pad  & ~n13928 ;
  assign n27918 = n13945 & n27917 ;
  assign n27919 = \m2_data_i[27]_pad  & n13928 ;
  assign n27920 = n13921 & n27919 ;
  assign n27921 = ~n27918 & ~n27920 ;
  assign n27922 = \m0_data_i[27]_pad  & n13928 ;
  assign n27923 = n13945 & n27922 ;
  assign n27924 = \m4_data_i[27]_pad  & n13928 ;
  assign n27925 = n13953 & n27924 ;
  assign n27926 = ~n27923 & ~n27925 ;
  assign n27927 = n27921 & n27926 ;
  assign n27928 = \m7_data_i[27]_pad  & ~n13928 ;
  assign n27929 = n13936 & n27928 ;
  assign n27930 = \m3_data_i[27]_pad  & ~n13928 ;
  assign n27931 = n13921 & n27930 ;
  assign n27932 = ~n27929 & ~n27931 ;
  assign n27933 = \m6_data_i[27]_pad  & n13928 ;
  assign n27934 = n13936 & n27933 ;
  assign n27935 = \m5_data_i[27]_pad  & ~n13928 ;
  assign n27936 = n13953 & n27935 ;
  assign n27937 = ~n27934 & ~n27936 ;
  assign n27938 = n27932 & n27937 ;
  assign n27939 = n27927 & n27938 ;
  assign n27940 = \m3_data_i[28]_pad  & ~n13928 ;
  assign n27941 = n13921 & n27940 ;
  assign n27942 = \m4_data_i[28]_pad  & n13928 ;
  assign n27943 = n13953 & n27942 ;
  assign n27944 = ~n27941 & ~n27943 ;
  assign n27945 = \m6_data_i[28]_pad  & n13928 ;
  assign n27946 = n13936 & n27945 ;
  assign n27947 = \m7_data_i[28]_pad  & ~n13928 ;
  assign n27948 = n13936 & n27947 ;
  assign n27949 = ~n27946 & ~n27948 ;
  assign n27950 = n27944 & n27949 ;
  assign n27951 = \m5_data_i[28]_pad  & ~n13928 ;
  assign n27952 = n13953 & n27951 ;
  assign n27953 = \m0_data_i[28]_pad  & n13928 ;
  assign n27954 = n13945 & n27953 ;
  assign n27955 = ~n27952 & ~n27954 ;
  assign n27956 = \m1_data_i[28]_pad  & ~n13928 ;
  assign n27957 = n13945 & n27956 ;
  assign n27958 = \m2_data_i[28]_pad  & n13928 ;
  assign n27959 = n13921 & n27958 ;
  assign n27960 = ~n27957 & ~n27959 ;
  assign n27961 = n27955 & n27960 ;
  assign n27962 = n27950 & n27961 ;
  assign n27963 = \m1_data_i[29]_pad  & ~n13928 ;
  assign n27964 = n13945 & n27963 ;
  assign n27965 = \m2_data_i[29]_pad  & n13928 ;
  assign n27966 = n13921 & n27965 ;
  assign n27967 = ~n27964 & ~n27966 ;
  assign n27968 = \m0_data_i[29]_pad  & n13928 ;
  assign n27969 = n13945 & n27968 ;
  assign n27970 = \m4_data_i[29]_pad  & n13928 ;
  assign n27971 = n13953 & n27970 ;
  assign n27972 = ~n27969 & ~n27971 ;
  assign n27973 = n27967 & n27972 ;
  assign n27974 = \m7_data_i[29]_pad  & ~n13928 ;
  assign n27975 = n13936 & n27974 ;
  assign n27976 = \m3_data_i[29]_pad  & ~n13928 ;
  assign n27977 = n13921 & n27976 ;
  assign n27978 = ~n27975 & ~n27977 ;
  assign n27979 = \m6_data_i[29]_pad  & n13928 ;
  assign n27980 = n13936 & n27979 ;
  assign n27981 = \m5_data_i[29]_pad  & ~n13928 ;
  assign n27982 = n13953 & n27981 ;
  assign n27983 = ~n27980 & ~n27982 ;
  assign n27984 = n27978 & n27983 ;
  assign n27985 = n27973 & n27984 ;
  assign n27986 = \m3_data_i[2]_pad  & ~n13928 ;
  assign n27987 = n13921 & n27986 ;
  assign n27988 = \m4_data_i[2]_pad  & n13928 ;
  assign n27989 = n13953 & n27988 ;
  assign n27990 = ~n27987 & ~n27989 ;
  assign n27991 = \m0_data_i[2]_pad  & n13928 ;
  assign n27992 = n13945 & n27991 ;
  assign n27993 = \m5_data_i[2]_pad  & ~n13928 ;
  assign n27994 = n13953 & n27993 ;
  assign n27995 = ~n27992 & ~n27994 ;
  assign n27996 = n27990 & n27995 ;
  assign n27997 = \m7_data_i[2]_pad  & ~n13928 ;
  assign n27998 = n13936 & n27997 ;
  assign n27999 = \m6_data_i[2]_pad  & n13928 ;
  assign n28000 = n13936 & n27999 ;
  assign n28001 = ~n27998 & ~n28000 ;
  assign n28002 = \m1_data_i[2]_pad  & ~n13928 ;
  assign n28003 = n13945 & n28002 ;
  assign n28004 = \m2_data_i[2]_pad  & n13928 ;
  assign n28005 = n13921 & n28004 ;
  assign n28006 = ~n28003 & ~n28005 ;
  assign n28007 = n28001 & n28006 ;
  assign n28008 = n27996 & n28007 ;
  assign n28009 = \m3_data_i[30]_pad  & ~n13928 ;
  assign n28010 = n13921 & n28009 ;
  assign n28011 = \m4_data_i[30]_pad  & n13928 ;
  assign n28012 = n13953 & n28011 ;
  assign n28013 = ~n28010 & ~n28012 ;
  assign n28014 = \m6_data_i[30]_pad  & n13928 ;
  assign n28015 = n13936 & n28014 ;
  assign n28016 = \m7_data_i[30]_pad  & ~n13928 ;
  assign n28017 = n13936 & n28016 ;
  assign n28018 = ~n28015 & ~n28017 ;
  assign n28019 = n28013 & n28018 ;
  assign n28020 = \m5_data_i[30]_pad  & ~n13928 ;
  assign n28021 = n13953 & n28020 ;
  assign n28022 = \m0_data_i[30]_pad  & n13928 ;
  assign n28023 = n13945 & n28022 ;
  assign n28024 = ~n28021 & ~n28023 ;
  assign n28025 = \m1_data_i[30]_pad  & ~n13928 ;
  assign n28026 = n13945 & n28025 ;
  assign n28027 = \m2_data_i[30]_pad  & n13928 ;
  assign n28028 = n13921 & n28027 ;
  assign n28029 = ~n28026 & ~n28028 ;
  assign n28030 = n28024 & n28029 ;
  assign n28031 = n28019 & n28030 ;
  assign n28032 = \m1_data_i[31]_pad  & ~n13928 ;
  assign n28033 = n13945 & n28032 ;
  assign n28034 = \m2_data_i[31]_pad  & n13928 ;
  assign n28035 = n13921 & n28034 ;
  assign n28036 = ~n28033 & ~n28035 ;
  assign n28037 = \m3_data_i[31]_pad  & ~n13928 ;
  assign n28038 = n13921 & n28037 ;
  assign n28039 = \m7_data_i[31]_pad  & ~n13928 ;
  assign n28040 = n13936 & n28039 ;
  assign n28041 = ~n28038 & ~n28040 ;
  assign n28042 = n28036 & n28041 ;
  assign n28043 = \m4_data_i[31]_pad  & n13928 ;
  assign n28044 = n13953 & n28043 ;
  assign n28045 = \m0_data_i[31]_pad  & n13928 ;
  assign n28046 = n13945 & n28045 ;
  assign n28047 = ~n28044 & ~n28046 ;
  assign n28048 = \m6_data_i[31]_pad  & n13928 ;
  assign n28049 = n13936 & n28048 ;
  assign n28050 = \m5_data_i[31]_pad  & ~n13928 ;
  assign n28051 = n13953 & n28050 ;
  assign n28052 = ~n28049 & ~n28051 ;
  assign n28053 = n28047 & n28052 ;
  assign n28054 = n28042 & n28053 ;
  assign n28055 = \m0_data_i[3]_pad  & n13928 ;
  assign n28056 = n13945 & n28055 ;
  assign n28057 = \m7_data_i[3]_pad  & ~n13928 ;
  assign n28058 = n13936 & n28057 ;
  assign n28059 = ~n28056 & ~n28058 ;
  assign n28060 = \m1_data_i[3]_pad  & ~n13928 ;
  assign n28061 = n13945 & n28060 ;
  assign n28062 = \m5_data_i[3]_pad  & ~n13928 ;
  assign n28063 = n13953 & n28062 ;
  assign n28064 = ~n28061 & ~n28063 ;
  assign n28065 = n28059 & n28064 ;
  assign n28066 = \m2_data_i[3]_pad  & n13928 ;
  assign n28067 = n13921 & n28066 ;
  assign n28068 = \m6_data_i[3]_pad  & n13928 ;
  assign n28069 = n13936 & n28068 ;
  assign n28070 = ~n28067 & ~n28069 ;
  assign n28071 = \m3_data_i[3]_pad  & ~n13928 ;
  assign n28072 = n13921 & n28071 ;
  assign n28073 = \m4_data_i[3]_pad  & n13928 ;
  assign n28074 = n13953 & n28073 ;
  assign n28075 = ~n28072 & ~n28074 ;
  assign n28076 = n28070 & n28075 ;
  assign n28077 = n28065 & n28076 ;
  assign n28078 = \m1_data_i[4]_pad  & ~n13928 ;
  assign n28079 = n13945 & n28078 ;
  assign n28080 = \m2_data_i[4]_pad  & n13928 ;
  assign n28081 = n13921 & n28080 ;
  assign n28082 = ~n28079 & ~n28081 ;
  assign n28083 = \m0_data_i[4]_pad  & n13928 ;
  assign n28084 = n13945 & n28083 ;
  assign n28085 = \m5_data_i[4]_pad  & ~n13928 ;
  assign n28086 = n13953 & n28085 ;
  assign n28087 = ~n28084 & ~n28086 ;
  assign n28088 = n28082 & n28087 ;
  assign n28089 = \m7_data_i[4]_pad  & ~n13928 ;
  assign n28090 = n13936 & n28089 ;
  assign n28091 = \m6_data_i[4]_pad  & n13928 ;
  assign n28092 = n13936 & n28091 ;
  assign n28093 = ~n28090 & ~n28092 ;
  assign n28094 = \m3_data_i[4]_pad  & ~n13928 ;
  assign n28095 = n13921 & n28094 ;
  assign n28096 = \m4_data_i[4]_pad  & n13928 ;
  assign n28097 = n13953 & n28096 ;
  assign n28098 = ~n28095 & ~n28097 ;
  assign n28099 = n28093 & n28098 ;
  assign n28100 = n28088 & n28099 ;
  assign n28101 = \m6_data_i[5]_pad  & n13928 ;
  assign n28102 = n13936 & n28101 ;
  assign n28103 = \m5_data_i[5]_pad  & ~n13928 ;
  assign n28104 = n13953 & n28103 ;
  assign n28105 = ~n28102 & ~n28104 ;
  assign n28106 = \m1_data_i[5]_pad  & ~n13928 ;
  assign n28107 = n13945 & n28106 ;
  assign n28108 = \m7_data_i[5]_pad  & ~n13928 ;
  assign n28109 = n13936 & n28108 ;
  assign n28110 = ~n28107 & ~n28109 ;
  assign n28111 = n28105 & n28110 ;
  assign n28112 = \m2_data_i[5]_pad  & n13928 ;
  assign n28113 = n13921 & n28112 ;
  assign n28114 = \m0_data_i[5]_pad  & n13928 ;
  assign n28115 = n13945 & n28114 ;
  assign n28116 = ~n28113 & ~n28115 ;
  assign n28117 = \m3_data_i[5]_pad  & ~n13928 ;
  assign n28118 = n13921 & n28117 ;
  assign n28119 = \m4_data_i[5]_pad  & n13928 ;
  assign n28120 = n13953 & n28119 ;
  assign n28121 = ~n28118 & ~n28120 ;
  assign n28122 = n28116 & n28121 ;
  assign n28123 = n28111 & n28122 ;
  assign n28124 = \m3_data_i[6]_pad  & ~n13928 ;
  assign n28125 = n13921 & n28124 ;
  assign n28126 = \m4_data_i[6]_pad  & n13928 ;
  assign n28127 = n13953 & n28126 ;
  assign n28128 = ~n28125 & ~n28127 ;
  assign n28129 = \m1_data_i[6]_pad  & ~n13928 ;
  assign n28130 = n13945 & n28129 ;
  assign n28131 = \m5_data_i[6]_pad  & ~n13928 ;
  assign n28132 = n13953 & n28131 ;
  assign n28133 = ~n28130 & ~n28132 ;
  assign n28134 = n28128 & n28133 ;
  assign n28135 = \m2_data_i[6]_pad  & n13928 ;
  assign n28136 = n13921 & n28135 ;
  assign n28137 = \m6_data_i[6]_pad  & n13928 ;
  assign n28138 = n13936 & n28137 ;
  assign n28139 = ~n28136 & ~n28138 ;
  assign n28140 = \m0_data_i[6]_pad  & n13928 ;
  assign n28141 = n13945 & n28140 ;
  assign n28142 = \m7_data_i[6]_pad  & ~n13928 ;
  assign n28143 = n13936 & n28142 ;
  assign n28144 = ~n28141 & ~n28143 ;
  assign n28145 = n28139 & n28144 ;
  assign n28146 = n28134 & n28145 ;
  assign n28147 = \m1_data_i[7]_pad  & ~n13928 ;
  assign n28148 = n13945 & n28147 ;
  assign n28149 = \m2_data_i[7]_pad  & n13928 ;
  assign n28150 = n13921 & n28149 ;
  assign n28151 = ~n28148 & ~n28150 ;
  assign n28152 = \m0_data_i[7]_pad  & n13928 ;
  assign n28153 = n13945 & n28152 ;
  assign n28154 = \m5_data_i[7]_pad  & ~n13928 ;
  assign n28155 = n13953 & n28154 ;
  assign n28156 = ~n28153 & ~n28155 ;
  assign n28157 = n28151 & n28156 ;
  assign n28158 = \m7_data_i[7]_pad  & ~n13928 ;
  assign n28159 = n13936 & n28158 ;
  assign n28160 = \m6_data_i[7]_pad  & n13928 ;
  assign n28161 = n13936 & n28160 ;
  assign n28162 = ~n28159 & ~n28161 ;
  assign n28163 = \m3_data_i[7]_pad  & ~n13928 ;
  assign n28164 = n13921 & n28163 ;
  assign n28165 = \m4_data_i[7]_pad  & n13928 ;
  assign n28166 = n13953 & n28165 ;
  assign n28167 = ~n28164 & ~n28166 ;
  assign n28168 = n28162 & n28167 ;
  assign n28169 = n28157 & n28168 ;
  assign n28170 = \m1_data_i[8]_pad  & ~n13928 ;
  assign n28171 = n13945 & n28170 ;
  assign n28172 = \m2_data_i[8]_pad  & n13928 ;
  assign n28173 = n13921 & n28172 ;
  assign n28174 = ~n28171 & ~n28173 ;
  assign n28175 = \m0_data_i[8]_pad  & n13928 ;
  assign n28176 = n13945 & n28175 ;
  assign n28177 = \m4_data_i[8]_pad  & n13928 ;
  assign n28178 = n13953 & n28177 ;
  assign n28179 = ~n28176 & ~n28178 ;
  assign n28180 = n28174 & n28179 ;
  assign n28181 = \m7_data_i[8]_pad  & ~n13928 ;
  assign n28182 = n13936 & n28181 ;
  assign n28183 = \m3_data_i[8]_pad  & ~n13928 ;
  assign n28184 = n13921 & n28183 ;
  assign n28185 = ~n28182 & ~n28184 ;
  assign n28186 = \m6_data_i[8]_pad  & n13928 ;
  assign n28187 = n13936 & n28186 ;
  assign n28188 = \m5_data_i[8]_pad  & ~n13928 ;
  assign n28189 = n13953 & n28188 ;
  assign n28190 = ~n28187 & ~n28189 ;
  assign n28191 = n28185 & n28190 ;
  assign n28192 = n28180 & n28191 ;
  assign n28193 = \m0_data_i[9]_pad  & n13928 ;
  assign n28194 = n13945 & n28193 ;
  assign n28195 = \m7_data_i[9]_pad  & ~n13928 ;
  assign n28196 = n13936 & n28195 ;
  assign n28197 = ~n28194 & ~n28196 ;
  assign n28198 = \m1_data_i[9]_pad  & ~n13928 ;
  assign n28199 = n13945 & n28198 ;
  assign n28200 = \m5_data_i[9]_pad  & ~n13928 ;
  assign n28201 = n13953 & n28200 ;
  assign n28202 = ~n28199 & ~n28201 ;
  assign n28203 = n28197 & n28202 ;
  assign n28204 = \m2_data_i[9]_pad  & n13928 ;
  assign n28205 = n13921 & n28204 ;
  assign n28206 = \m6_data_i[9]_pad  & n13928 ;
  assign n28207 = n13936 & n28206 ;
  assign n28208 = ~n28205 & ~n28207 ;
  assign n28209 = \m3_data_i[9]_pad  & ~n13928 ;
  assign n28210 = n13921 & n28209 ;
  assign n28211 = \m4_data_i[9]_pad  & n13928 ;
  assign n28212 = n13953 & n28211 ;
  assign n28213 = ~n28210 & ~n28212 ;
  assign n28214 = n28208 & n28213 ;
  assign n28215 = n28203 & n28214 ;
  assign n28216 = \m0_sel_i[0]_pad  & n13928 ;
  assign n28217 = n13945 & n28216 ;
  assign n28218 = \m7_sel_i[0]_pad  & ~n13928 ;
  assign n28219 = n13936 & n28218 ;
  assign n28220 = ~n28217 & ~n28219 ;
  assign n28221 = \m3_sel_i[0]_pad  & ~n13928 ;
  assign n28222 = n13921 & n28221 ;
  assign n28223 = \m2_sel_i[0]_pad  & n13928 ;
  assign n28224 = n13921 & n28223 ;
  assign n28225 = ~n28222 & ~n28224 ;
  assign n28226 = n28220 & n28225 ;
  assign n28227 = \m4_sel_i[0]_pad  & n13928 ;
  assign n28228 = n13953 & n28227 ;
  assign n28229 = \m1_sel_i[0]_pad  & ~n13928 ;
  assign n28230 = n13945 & n28229 ;
  assign n28231 = ~n28228 & ~n28230 ;
  assign n28232 = \m6_sel_i[0]_pad  & n13928 ;
  assign n28233 = n13936 & n28232 ;
  assign n28234 = \m5_sel_i[0]_pad  & ~n13928 ;
  assign n28235 = n13953 & n28234 ;
  assign n28236 = ~n28233 & ~n28235 ;
  assign n28237 = n28231 & n28236 ;
  assign n28238 = n28226 & n28237 ;
  assign n28239 = \m0_sel_i[1]_pad  & n13928 ;
  assign n28240 = n13945 & n28239 ;
  assign n28241 = \m7_sel_i[1]_pad  & ~n13928 ;
  assign n28242 = n13936 & n28241 ;
  assign n28243 = ~n28240 & ~n28242 ;
  assign n28244 = \m1_sel_i[1]_pad  & ~n13928 ;
  assign n28245 = n13945 & n28244 ;
  assign n28246 = \m4_sel_i[1]_pad  & n13928 ;
  assign n28247 = n13953 & n28246 ;
  assign n28248 = ~n28245 & ~n28247 ;
  assign n28249 = n28243 & n28248 ;
  assign n28250 = \m2_sel_i[1]_pad  & n13928 ;
  assign n28251 = n13921 & n28250 ;
  assign n28252 = \m3_sel_i[1]_pad  & ~n13928 ;
  assign n28253 = n13921 & n28252 ;
  assign n28254 = ~n28251 & ~n28253 ;
  assign n28255 = \m6_sel_i[1]_pad  & n13928 ;
  assign n28256 = n13936 & n28255 ;
  assign n28257 = \m5_sel_i[1]_pad  & ~n13928 ;
  assign n28258 = n13953 & n28257 ;
  assign n28259 = ~n28256 & ~n28258 ;
  assign n28260 = n28254 & n28259 ;
  assign n28261 = n28249 & n28260 ;
  assign n28262 = \m1_sel_i[2]_pad  & ~n13928 ;
  assign n28263 = n13945 & n28262 ;
  assign n28264 = \m2_sel_i[2]_pad  & n13928 ;
  assign n28265 = n13921 & n28264 ;
  assign n28266 = ~n28263 & ~n28265 ;
  assign n28267 = \m0_sel_i[2]_pad  & n13928 ;
  assign n28268 = n13945 & n28267 ;
  assign n28269 = \m4_sel_i[2]_pad  & n13928 ;
  assign n28270 = n13953 & n28269 ;
  assign n28271 = ~n28268 & ~n28270 ;
  assign n28272 = n28266 & n28271 ;
  assign n28273 = \m7_sel_i[2]_pad  & ~n13928 ;
  assign n28274 = n13936 & n28273 ;
  assign n28275 = \m3_sel_i[2]_pad  & ~n13928 ;
  assign n28276 = n13921 & n28275 ;
  assign n28277 = ~n28274 & ~n28276 ;
  assign n28278 = \m6_sel_i[2]_pad  & n13928 ;
  assign n28279 = n13936 & n28278 ;
  assign n28280 = \m5_sel_i[2]_pad  & ~n13928 ;
  assign n28281 = n13953 & n28280 ;
  assign n28282 = ~n28279 & ~n28281 ;
  assign n28283 = n28277 & n28282 ;
  assign n28284 = n28272 & n28283 ;
  assign n28285 = \m1_sel_i[3]_pad  & ~n13928 ;
  assign n28286 = n13945 & n28285 ;
  assign n28287 = \m2_sel_i[3]_pad  & n13928 ;
  assign n28288 = n13921 & n28287 ;
  assign n28289 = ~n28286 & ~n28288 ;
  assign n28290 = \m0_sel_i[3]_pad  & n13928 ;
  assign n28291 = n13945 & n28290 ;
  assign n28292 = \m4_sel_i[3]_pad  & n13928 ;
  assign n28293 = n13953 & n28292 ;
  assign n28294 = ~n28291 & ~n28293 ;
  assign n28295 = n28289 & n28294 ;
  assign n28296 = \m7_sel_i[3]_pad  & ~n13928 ;
  assign n28297 = n13936 & n28296 ;
  assign n28298 = \m3_sel_i[3]_pad  & ~n13928 ;
  assign n28299 = n13921 & n28298 ;
  assign n28300 = ~n28297 & ~n28299 ;
  assign n28301 = \m6_sel_i[3]_pad  & n13928 ;
  assign n28302 = n13936 & n28301 ;
  assign n28303 = \m5_sel_i[3]_pad  & ~n13928 ;
  assign n28304 = n13953 & n28303 ;
  assign n28305 = ~n28302 & ~n28304 ;
  assign n28306 = n28300 & n28305 ;
  assign n28307 = n28295 & n28306 ;
  assign n28308 = \m3_stb_i_pad  & n14892 ;
  assign n28309 = ~n13928 & n28308 ;
  assign n28310 = n13921 & n28309 ;
  assign n28311 = \m2_stb_i_pad  & n14851 ;
  assign n28312 = n13928 & n28311 ;
  assign n28313 = n13921 & n28312 ;
  assign n28314 = ~n28310 & ~n28313 ;
  assign n28315 = \m6_stb_i_pad  & n14999 ;
  assign n28316 = n13928 & n28315 ;
  assign n28317 = n13936 & n28316 ;
  assign n28318 = \m1_stb_i_pad  & n14797 ;
  assign n28319 = ~n13928 & n28318 ;
  assign n28320 = n13945 & n28319 ;
  assign n28321 = ~n28317 & ~n28320 ;
  assign n28322 = n28314 & n28321 ;
  assign n28323 = \m7_stb_i_pad  & n15047 ;
  assign n28324 = ~n13928 & n28323 ;
  assign n28325 = n13936 & n28324 ;
  assign n28326 = \m5_stb_i_pad  & n14963 ;
  assign n28327 = ~n13928 & n28326 ;
  assign n28328 = n13953 & n28327 ;
  assign n28329 = ~n28325 & ~n28328 ;
  assign n28330 = \m4_stb_i_pad  & n14931 ;
  assign n28331 = n13928 & n28330 ;
  assign n28332 = n13953 & n28331 ;
  assign n28333 = \m0_stb_i_pad  & n14749 ;
  assign n28334 = n13928 & n28333 ;
  assign n28335 = n13945 & n28334 ;
  assign n28336 = ~n28332 & ~n28335 ;
  assign n28337 = n28329 & n28336 ;
  assign n28338 = n28322 & n28337 ;
  assign n28339 = \m6_we_i_pad  & n13928 ;
  assign n28340 = n13936 & n28339 ;
  assign n28341 = \m5_we_i_pad  & ~n13928 ;
  assign n28342 = n13953 & n28341 ;
  assign n28343 = ~n28340 & ~n28342 ;
  assign n28344 = \m3_we_i_pad  & ~n13928 ;
  assign n28345 = n13921 & n28344 ;
  assign n28346 = \m7_we_i_pad  & ~n13928 ;
  assign n28347 = n13936 & n28346 ;
  assign n28348 = ~n28345 & ~n28347 ;
  assign n28349 = n28343 & n28348 ;
  assign n28350 = \m4_we_i_pad  & n13928 ;
  assign n28351 = n13953 & n28350 ;
  assign n28352 = \m0_we_i_pad  & n13928 ;
  assign n28353 = n13945 & n28352 ;
  assign n28354 = ~n28351 & ~n28353 ;
  assign n28355 = \m1_we_i_pad  & ~n13928 ;
  assign n28356 = n13945 & n28355 ;
  assign n28357 = \m2_we_i_pad  & n13928 ;
  assign n28358 = n13921 & n28357 ;
  assign n28359 = ~n28356 & ~n28358 ;
  assign n28360 = n28354 & n28359 ;
  assign n28361 = n28349 & n28360 ;
  assign n28362 = \m1_addr_i[0]_pad  & ~n14009 ;
  assign n28363 = n14017 & n28362 ;
  assign n28364 = \m2_addr_i[0]_pad  & n14009 ;
  assign n28365 = n14034 & n28364 ;
  assign n28366 = ~n28363 & ~n28365 ;
  assign n28367 = \m0_addr_i[0]_pad  & n14009 ;
  assign n28368 = n14017 & n28367 ;
  assign n28369 = \m5_addr_i[0]_pad  & ~n14009 ;
  assign n28370 = n14002 & n28369 ;
  assign n28371 = ~n28368 & ~n28370 ;
  assign n28372 = n28366 & n28371 ;
  assign n28373 = \m7_addr_i[0]_pad  & ~n14009 ;
  assign n28374 = n14026 & n28373 ;
  assign n28375 = \m6_addr_i[0]_pad  & n14009 ;
  assign n28376 = n14026 & n28375 ;
  assign n28377 = ~n28374 & ~n28376 ;
  assign n28378 = \m3_addr_i[0]_pad  & ~n14009 ;
  assign n28379 = n14034 & n28378 ;
  assign n28380 = \m4_addr_i[0]_pad  & n14009 ;
  assign n28381 = n14002 & n28380 ;
  assign n28382 = ~n28379 & ~n28381 ;
  assign n28383 = n28377 & n28382 ;
  assign n28384 = n28372 & n28383 ;
  assign n28385 = \m1_addr_i[10]_pad  & ~n14009 ;
  assign n28386 = n14017 & n28385 ;
  assign n28387 = \m2_addr_i[10]_pad  & n14009 ;
  assign n28388 = n14034 & n28387 ;
  assign n28389 = ~n28386 & ~n28388 ;
  assign n28390 = \m6_addr_i[10]_pad  & n14009 ;
  assign n28391 = n14026 & n28390 ;
  assign n28392 = \m4_addr_i[10]_pad  & n14009 ;
  assign n28393 = n14002 & n28392 ;
  assign n28394 = ~n28391 & ~n28393 ;
  assign n28395 = n28389 & n28394 ;
  assign n28396 = \m5_addr_i[10]_pad  & ~n14009 ;
  assign n28397 = n14002 & n28396 ;
  assign n28398 = \m3_addr_i[10]_pad  & ~n14009 ;
  assign n28399 = n14034 & n28398 ;
  assign n28400 = ~n28397 & ~n28399 ;
  assign n28401 = \m0_addr_i[10]_pad  & n14009 ;
  assign n28402 = n14017 & n28401 ;
  assign n28403 = \m7_addr_i[10]_pad  & ~n14009 ;
  assign n28404 = n14026 & n28403 ;
  assign n28405 = ~n28402 & ~n28404 ;
  assign n28406 = n28400 & n28405 ;
  assign n28407 = n28395 & n28406 ;
  assign n28408 = \m1_addr_i[11]_pad  & ~n14009 ;
  assign n28409 = n14017 & n28408 ;
  assign n28410 = \m2_addr_i[11]_pad  & n14009 ;
  assign n28411 = n14034 & n28410 ;
  assign n28412 = ~n28409 & ~n28411 ;
  assign n28413 = \m3_addr_i[11]_pad  & ~n14009 ;
  assign n28414 = n14034 & n28413 ;
  assign n28415 = \m5_addr_i[11]_pad  & ~n14009 ;
  assign n28416 = n14002 & n28415 ;
  assign n28417 = ~n28414 & ~n28416 ;
  assign n28418 = n28412 & n28417 ;
  assign n28419 = \m4_addr_i[11]_pad  & n14009 ;
  assign n28420 = n14002 & n28419 ;
  assign n28421 = \m6_addr_i[11]_pad  & n14009 ;
  assign n28422 = n14026 & n28421 ;
  assign n28423 = ~n28420 & ~n28422 ;
  assign n28424 = \m0_addr_i[11]_pad  & n14009 ;
  assign n28425 = n14017 & n28424 ;
  assign n28426 = \m7_addr_i[11]_pad  & ~n14009 ;
  assign n28427 = n14026 & n28426 ;
  assign n28428 = ~n28425 & ~n28427 ;
  assign n28429 = n28423 & n28428 ;
  assign n28430 = n28418 & n28429 ;
  assign n28431 = \m0_addr_i[12]_pad  & n14009 ;
  assign n28432 = n14017 & n28431 ;
  assign n28433 = \m7_addr_i[12]_pad  & ~n14009 ;
  assign n28434 = n14026 & n28433 ;
  assign n28435 = ~n28432 & ~n28434 ;
  assign n28436 = \m6_addr_i[12]_pad  & n14009 ;
  assign n28437 = n14026 & n28436 ;
  assign n28438 = \m4_addr_i[12]_pad  & n14009 ;
  assign n28439 = n14002 & n28438 ;
  assign n28440 = ~n28437 & ~n28439 ;
  assign n28441 = n28435 & n28440 ;
  assign n28442 = \m5_addr_i[12]_pad  & ~n14009 ;
  assign n28443 = n14002 & n28442 ;
  assign n28444 = \m3_addr_i[12]_pad  & ~n14009 ;
  assign n28445 = n14034 & n28444 ;
  assign n28446 = ~n28443 & ~n28445 ;
  assign n28447 = \m1_addr_i[12]_pad  & ~n14009 ;
  assign n28448 = n14017 & n28447 ;
  assign n28449 = \m2_addr_i[12]_pad  & n14009 ;
  assign n28450 = n14034 & n28449 ;
  assign n28451 = ~n28448 & ~n28450 ;
  assign n28452 = n28446 & n28451 ;
  assign n28453 = n28441 & n28452 ;
  assign n28454 = \m3_addr_i[13]_pad  & ~n14009 ;
  assign n28455 = n14034 & n28454 ;
  assign n28456 = \m4_addr_i[13]_pad  & n14009 ;
  assign n28457 = n14002 & n28456 ;
  assign n28458 = ~n28455 & ~n28457 ;
  assign n28459 = \m1_addr_i[13]_pad  & ~n14009 ;
  assign n28460 = n14017 & n28459 ;
  assign n28461 = \m7_addr_i[13]_pad  & ~n14009 ;
  assign n28462 = n14026 & n28461 ;
  assign n28463 = ~n28460 & ~n28462 ;
  assign n28464 = n28458 & n28463 ;
  assign n28465 = \m2_addr_i[13]_pad  & n14009 ;
  assign n28466 = n14034 & n28465 ;
  assign n28467 = \m0_addr_i[13]_pad  & n14009 ;
  assign n28468 = n14017 & n28467 ;
  assign n28469 = ~n28466 & ~n28468 ;
  assign n28470 = \m6_addr_i[13]_pad  & n14009 ;
  assign n28471 = n14026 & n28470 ;
  assign n28472 = \m5_addr_i[13]_pad  & ~n14009 ;
  assign n28473 = n14002 & n28472 ;
  assign n28474 = ~n28471 & ~n28473 ;
  assign n28475 = n28469 & n28474 ;
  assign n28476 = n28464 & n28475 ;
  assign n28477 = \m1_addr_i[14]_pad  & ~n14009 ;
  assign n28478 = n14017 & n28477 ;
  assign n28479 = \m2_addr_i[14]_pad  & n14009 ;
  assign n28480 = n14034 & n28479 ;
  assign n28481 = ~n28478 & ~n28480 ;
  assign n28482 = \m0_addr_i[14]_pad  & n14009 ;
  assign n28483 = n14017 & n28482 ;
  assign n28484 = \m4_addr_i[14]_pad  & n14009 ;
  assign n28485 = n14002 & n28484 ;
  assign n28486 = ~n28483 & ~n28485 ;
  assign n28487 = n28481 & n28486 ;
  assign n28488 = \m7_addr_i[14]_pad  & ~n14009 ;
  assign n28489 = n14026 & n28488 ;
  assign n28490 = \m3_addr_i[14]_pad  & ~n14009 ;
  assign n28491 = n14034 & n28490 ;
  assign n28492 = ~n28489 & ~n28491 ;
  assign n28493 = \m6_addr_i[14]_pad  & n14009 ;
  assign n28494 = n14026 & n28493 ;
  assign n28495 = \m5_addr_i[14]_pad  & ~n14009 ;
  assign n28496 = n14002 & n28495 ;
  assign n28497 = ~n28494 & ~n28496 ;
  assign n28498 = n28492 & n28497 ;
  assign n28499 = n28487 & n28498 ;
  assign n28500 = \m6_addr_i[15]_pad  & n14009 ;
  assign n28501 = n14026 & n28500 ;
  assign n28502 = \m5_addr_i[15]_pad  & ~n14009 ;
  assign n28503 = n14002 & n28502 ;
  assign n28504 = ~n28501 & ~n28503 ;
  assign n28505 = \m3_addr_i[15]_pad  & ~n14009 ;
  assign n28506 = n14034 & n28505 ;
  assign n28507 = \m2_addr_i[15]_pad  & n14009 ;
  assign n28508 = n14034 & n28507 ;
  assign n28509 = ~n28506 & ~n28508 ;
  assign n28510 = n28504 & n28509 ;
  assign n28511 = \m4_addr_i[15]_pad  & n14009 ;
  assign n28512 = n14002 & n28511 ;
  assign n28513 = \m1_addr_i[15]_pad  & ~n14009 ;
  assign n28514 = n14017 & n28513 ;
  assign n28515 = ~n28512 & ~n28514 ;
  assign n28516 = \m0_addr_i[15]_pad  & n14009 ;
  assign n28517 = n14017 & n28516 ;
  assign n28518 = \m7_addr_i[15]_pad  & ~n14009 ;
  assign n28519 = n14026 & n28518 ;
  assign n28520 = ~n28517 & ~n28519 ;
  assign n28521 = n28515 & n28520 ;
  assign n28522 = n28510 & n28521 ;
  assign n28523 = \m0_addr_i[16]_pad  & n14009 ;
  assign n28524 = n14017 & n28523 ;
  assign n28525 = \m7_addr_i[16]_pad  & ~n14009 ;
  assign n28526 = n14026 & n28525 ;
  assign n28527 = ~n28524 & ~n28526 ;
  assign n28528 = \m6_addr_i[16]_pad  & n14009 ;
  assign n28529 = n14026 & n28528 ;
  assign n28530 = \m4_addr_i[16]_pad  & n14009 ;
  assign n28531 = n14002 & n28530 ;
  assign n28532 = ~n28529 & ~n28531 ;
  assign n28533 = n28527 & n28532 ;
  assign n28534 = \m5_addr_i[16]_pad  & ~n14009 ;
  assign n28535 = n14002 & n28534 ;
  assign n28536 = \m3_addr_i[16]_pad  & ~n14009 ;
  assign n28537 = n14034 & n28536 ;
  assign n28538 = ~n28535 & ~n28537 ;
  assign n28539 = \m1_addr_i[16]_pad  & ~n14009 ;
  assign n28540 = n14017 & n28539 ;
  assign n28541 = \m2_addr_i[16]_pad  & n14009 ;
  assign n28542 = n14034 & n28541 ;
  assign n28543 = ~n28540 & ~n28542 ;
  assign n28544 = n28538 & n28543 ;
  assign n28545 = n28533 & n28544 ;
  assign n28546 = \m6_addr_i[17]_pad  & n14009 ;
  assign n28547 = n14026 & n28546 ;
  assign n28548 = \m5_addr_i[17]_pad  & ~n14009 ;
  assign n28549 = n14002 & n28548 ;
  assign n28550 = ~n28547 & ~n28549 ;
  assign n28551 = \m0_addr_i[17]_pad  & n14009 ;
  assign n28552 = n14017 & n28551 ;
  assign n28553 = \m2_addr_i[17]_pad  & n14009 ;
  assign n28554 = n14034 & n28553 ;
  assign n28555 = ~n28552 & ~n28554 ;
  assign n28556 = n28550 & n28555 ;
  assign n28557 = \m7_addr_i[17]_pad  & ~n14009 ;
  assign n28558 = n14026 & n28557 ;
  assign n28559 = \m1_addr_i[17]_pad  & ~n14009 ;
  assign n28560 = n14017 & n28559 ;
  assign n28561 = ~n28558 & ~n28560 ;
  assign n28562 = \m3_addr_i[17]_pad  & ~n14009 ;
  assign n28563 = n14034 & n28562 ;
  assign n28564 = \m4_addr_i[17]_pad  & n14009 ;
  assign n28565 = n14002 & n28564 ;
  assign n28566 = ~n28563 & ~n28565 ;
  assign n28567 = n28561 & n28566 ;
  assign n28568 = n28556 & n28567 ;
  assign n28569 = \m6_addr_i[18]_pad  & n14009 ;
  assign n28570 = n14026 & n28569 ;
  assign n28571 = \m5_addr_i[18]_pad  & ~n14009 ;
  assign n28572 = n14002 & n28571 ;
  assign n28573 = ~n28570 & ~n28572 ;
  assign n28574 = \m0_addr_i[18]_pad  & n14009 ;
  assign n28575 = n14017 & n28574 ;
  assign n28576 = \m4_addr_i[18]_pad  & n14009 ;
  assign n28577 = n14002 & n28576 ;
  assign n28578 = ~n28575 & ~n28577 ;
  assign n28579 = n28573 & n28578 ;
  assign n28580 = \m7_addr_i[18]_pad  & ~n14009 ;
  assign n28581 = n14026 & n28580 ;
  assign n28582 = \m3_addr_i[18]_pad  & ~n14009 ;
  assign n28583 = n14034 & n28582 ;
  assign n28584 = ~n28581 & ~n28583 ;
  assign n28585 = \m1_addr_i[18]_pad  & ~n14009 ;
  assign n28586 = n14017 & n28585 ;
  assign n28587 = \m2_addr_i[18]_pad  & n14009 ;
  assign n28588 = n14034 & n28587 ;
  assign n28589 = ~n28586 & ~n28588 ;
  assign n28590 = n28584 & n28589 ;
  assign n28591 = n28579 & n28590 ;
  assign n28592 = \m6_addr_i[19]_pad  & n14009 ;
  assign n28593 = n14026 & n28592 ;
  assign n28594 = \m5_addr_i[19]_pad  & ~n14009 ;
  assign n28595 = n14002 & n28594 ;
  assign n28596 = ~n28593 & ~n28595 ;
  assign n28597 = \m0_addr_i[19]_pad  & n14009 ;
  assign n28598 = n14017 & n28597 ;
  assign n28599 = \m4_addr_i[19]_pad  & n14009 ;
  assign n28600 = n14002 & n28599 ;
  assign n28601 = ~n28598 & ~n28600 ;
  assign n28602 = n28596 & n28601 ;
  assign n28603 = \m7_addr_i[19]_pad  & ~n14009 ;
  assign n28604 = n14026 & n28603 ;
  assign n28605 = \m3_addr_i[19]_pad  & ~n14009 ;
  assign n28606 = n14034 & n28605 ;
  assign n28607 = ~n28604 & ~n28606 ;
  assign n28608 = \m1_addr_i[19]_pad  & ~n14009 ;
  assign n28609 = n14017 & n28608 ;
  assign n28610 = \m2_addr_i[19]_pad  & n14009 ;
  assign n28611 = n14034 & n28610 ;
  assign n28612 = ~n28609 & ~n28611 ;
  assign n28613 = n28607 & n28612 ;
  assign n28614 = n28602 & n28613 ;
  assign n28615 = \m6_addr_i[1]_pad  & n14009 ;
  assign n28616 = n14026 & n28615 ;
  assign n28617 = \m5_addr_i[1]_pad  & ~n14009 ;
  assign n28618 = n14002 & n28617 ;
  assign n28619 = ~n28616 & ~n28618 ;
  assign n28620 = \m0_addr_i[1]_pad  & n14009 ;
  assign n28621 = n14017 & n28620 ;
  assign n28622 = \m4_addr_i[1]_pad  & n14009 ;
  assign n28623 = n14002 & n28622 ;
  assign n28624 = ~n28621 & ~n28623 ;
  assign n28625 = n28619 & n28624 ;
  assign n28626 = \m7_addr_i[1]_pad  & ~n14009 ;
  assign n28627 = n14026 & n28626 ;
  assign n28628 = \m3_addr_i[1]_pad  & ~n14009 ;
  assign n28629 = n14034 & n28628 ;
  assign n28630 = ~n28627 & ~n28629 ;
  assign n28631 = \m1_addr_i[1]_pad  & ~n14009 ;
  assign n28632 = n14017 & n28631 ;
  assign n28633 = \m2_addr_i[1]_pad  & n14009 ;
  assign n28634 = n14034 & n28633 ;
  assign n28635 = ~n28632 & ~n28634 ;
  assign n28636 = n28630 & n28635 ;
  assign n28637 = n28625 & n28636 ;
  assign n28638 = \m1_addr_i[20]_pad  & ~n14009 ;
  assign n28639 = n14017 & n28638 ;
  assign n28640 = \m2_addr_i[20]_pad  & n14009 ;
  assign n28641 = n14034 & n28640 ;
  assign n28642 = ~n28639 & ~n28641 ;
  assign n28643 = \m3_addr_i[20]_pad  & ~n14009 ;
  assign n28644 = n14034 & n28643 ;
  assign n28645 = \m7_addr_i[20]_pad  & ~n14009 ;
  assign n28646 = n14026 & n28645 ;
  assign n28647 = ~n28644 & ~n28646 ;
  assign n28648 = n28642 & n28647 ;
  assign n28649 = \m4_addr_i[20]_pad  & n14009 ;
  assign n28650 = n14002 & n28649 ;
  assign n28651 = \m0_addr_i[20]_pad  & n14009 ;
  assign n28652 = n14017 & n28651 ;
  assign n28653 = ~n28650 & ~n28652 ;
  assign n28654 = \m6_addr_i[20]_pad  & n14009 ;
  assign n28655 = n14026 & n28654 ;
  assign n28656 = \m5_addr_i[20]_pad  & ~n14009 ;
  assign n28657 = n14002 & n28656 ;
  assign n28658 = ~n28655 & ~n28657 ;
  assign n28659 = n28653 & n28658 ;
  assign n28660 = n28648 & n28659 ;
  assign n28661 = \m1_addr_i[21]_pad  & ~n14009 ;
  assign n28662 = n14017 & n28661 ;
  assign n28663 = \m2_addr_i[21]_pad  & n14009 ;
  assign n28664 = n14034 & n28663 ;
  assign n28665 = ~n28662 & ~n28664 ;
  assign n28666 = \m3_addr_i[21]_pad  & ~n14009 ;
  assign n28667 = n14034 & n28666 ;
  assign n28668 = \m5_addr_i[21]_pad  & ~n14009 ;
  assign n28669 = n14002 & n28668 ;
  assign n28670 = ~n28667 & ~n28669 ;
  assign n28671 = n28665 & n28670 ;
  assign n28672 = \m4_addr_i[21]_pad  & n14009 ;
  assign n28673 = n14002 & n28672 ;
  assign n28674 = \m6_addr_i[21]_pad  & n14009 ;
  assign n28675 = n14026 & n28674 ;
  assign n28676 = ~n28673 & ~n28675 ;
  assign n28677 = \m0_addr_i[21]_pad  & n14009 ;
  assign n28678 = n14017 & n28677 ;
  assign n28679 = \m7_addr_i[21]_pad  & ~n14009 ;
  assign n28680 = n14026 & n28679 ;
  assign n28681 = ~n28678 & ~n28680 ;
  assign n28682 = n28676 & n28681 ;
  assign n28683 = n28671 & n28682 ;
  assign n28684 = \m0_addr_i[22]_pad  & n14009 ;
  assign n28685 = n14017 & n28684 ;
  assign n28686 = \m7_addr_i[22]_pad  & ~n14009 ;
  assign n28687 = n14026 & n28686 ;
  assign n28688 = ~n28685 & ~n28687 ;
  assign n28689 = \m6_addr_i[22]_pad  & n14009 ;
  assign n28690 = n14026 & n28689 ;
  assign n28691 = \m2_addr_i[22]_pad  & n14009 ;
  assign n28692 = n14034 & n28691 ;
  assign n28693 = ~n28690 & ~n28692 ;
  assign n28694 = n28688 & n28693 ;
  assign n28695 = \m5_addr_i[22]_pad  & ~n14009 ;
  assign n28696 = n14002 & n28695 ;
  assign n28697 = \m1_addr_i[22]_pad  & ~n14009 ;
  assign n28698 = n14017 & n28697 ;
  assign n28699 = ~n28696 & ~n28698 ;
  assign n28700 = \m3_addr_i[22]_pad  & ~n14009 ;
  assign n28701 = n14034 & n28700 ;
  assign n28702 = \m4_addr_i[22]_pad  & n14009 ;
  assign n28703 = n14002 & n28702 ;
  assign n28704 = ~n28701 & ~n28703 ;
  assign n28705 = n28699 & n28704 ;
  assign n28706 = n28694 & n28705 ;
  assign n28707 = \m3_addr_i[23]_pad  & ~n14009 ;
  assign n28708 = n14034 & n28707 ;
  assign n28709 = \m4_addr_i[23]_pad  & n14009 ;
  assign n28710 = n14002 & n28709 ;
  assign n28711 = ~n28708 & ~n28710 ;
  assign n28712 = \m1_addr_i[23]_pad  & ~n14009 ;
  assign n28713 = n14017 & n28712 ;
  assign n28714 = \m5_addr_i[23]_pad  & ~n14009 ;
  assign n28715 = n14002 & n28714 ;
  assign n28716 = ~n28713 & ~n28715 ;
  assign n28717 = n28711 & n28716 ;
  assign n28718 = \m2_addr_i[23]_pad  & n14009 ;
  assign n28719 = n14034 & n28718 ;
  assign n28720 = \m6_addr_i[23]_pad  & n14009 ;
  assign n28721 = n14026 & n28720 ;
  assign n28722 = ~n28719 & ~n28721 ;
  assign n28723 = \m0_addr_i[23]_pad  & n14009 ;
  assign n28724 = n14017 & n28723 ;
  assign n28725 = \m7_addr_i[23]_pad  & ~n14009 ;
  assign n28726 = n14026 & n28725 ;
  assign n28727 = ~n28724 & ~n28726 ;
  assign n28728 = n28722 & n28727 ;
  assign n28729 = n28717 & n28728 ;
  assign n28730 = \m1_addr_i[24]_pad  & ~n14009 ;
  assign n28731 = n14017 & n28730 ;
  assign n28732 = \m2_addr_i[24]_pad  & n14009 ;
  assign n28733 = n14034 & n28732 ;
  assign n28734 = ~n28731 & ~n28733 ;
  assign n28735 = \m0_addr_i[24]_pad  & n14009 ;
  assign n28736 = n14017 & n28735 ;
  assign n28737 = \m4_addr_i[24]_pad  & n14009 ;
  assign n28738 = n14002 & n28737 ;
  assign n28739 = ~n28736 & ~n28738 ;
  assign n28740 = n28734 & n28739 ;
  assign n28741 = \m7_addr_i[24]_pad  & ~n14009 ;
  assign n28742 = n14026 & n28741 ;
  assign n28743 = \m3_addr_i[24]_pad  & ~n14009 ;
  assign n28744 = n14034 & n28743 ;
  assign n28745 = ~n28742 & ~n28744 ;
  assign n28746 = \m5_addr_i[24]_pad  & ~n14009 ;
  assign n28747 = n14002 & n28746 ;
  assign n28748 = \m6_addr_i[24]_pad  & n14009 ;
  assign n28749 = n14026 & n28748 ;
  assign n28750 = ~n28747 & ~n28749 ;
  assign n28751 = n28745 & n28750 ;
  assign n28752 = n28740 & n28751 ;
  assign n28753 = \m0_addr_i[25]_pad  & n14009 ;
  assign n28754 = n14017 & n28753 ;
  assign n28755 = \m7_addr_i[25]_pad  & ~n14009 ;
  assign n28756 = n14026 & n28755 ;
  assign n28757 = ~n28754 & ~n28756 ;
  assign n28758 = \m1_addr_i[25]_pad  & ~n14009 ;
  assign n28759 = n14017 & n28758 ;
  assign n28760 = \m6_addr_i[25]_pad  & n14009 ;
  assign n28761 = n14026 & n28760 ;
  assign n28762 = ~n28759 & ~n28761 ;
  assign n28763 = n28757 & n28762 ;
  assign n28764 = \m2_addr_i[25]_pad  & n14009 ;
  assign n28765 = n14034 & n28764 ;
  assign n28766 = \m5_addr_i[25]_pad  & ~n14009 ;
  assign n28767 = n14002 & n28766 ;
  assign n28768 = ~n28765 & ~n28767 ;
  assign n28769 = \m3_addr_i[25]_pad  & ~n14009 ;
  assign n28770 = n14034 & n28769 ;
  assign n28771 = \m4_addr_i[25]_pad  & n14009 ;
  assign n28772 = n14002 & n28771 ;
  assign n28773 = ~n28770 & ~n28772 ;
  assign n28774 = n28768 & n28773 ;
  assign n28775 = n28763 & n28774 ;
  assign n28776 = \m3_addr_i[26]_pad  & ~n14009 ;
  assign n28777 = n14034 & n28776 ;
  assign n28778 = \m4_addr_i[26]_pad  & n14009 ;
  assign n28779 = n14002 & n28778 ;
  assign n28780 = ~n28777 & ~n28779 ;
  assign n28781 = \m5_addr_i[26]_pad  & ~n14009 ;
  assign n28782 = n14002 & n28781 ;
  assign n28783 = \m2_addr_i[26]_pad  & n14009 ;
  assign n28784 = n14034 & n28783 ;
  assign n28785 = ~n28782 & ~n28784 ;
  assign n28786 = n28780 & n28785 ;
  assign n28787 = \m6_addr_i[26]_pad  & n14009 ;
  assign n28788 = n14026 & n28787 ;
  assign n28789 = \m1_addr_i[26]_pad  & ~n14009 ;
  assign n28790 = n14017 & n28789 ;
  assign n28791 = ~n28788 & ~n28790 ;
  assign n28792 = \m0_addr_i[26]_pad  & n14009 ;
  assign n28793 = n14017 & n28792 ;
  assign n28794 = \m7_addr_i[26]_pad  & ~n14009 ;
  assign n28795 = n14026 & n28794 ;
  assign n28796 = ~n28793 & ~n28795 ;
  assign n28797 = n28791 & n28796 ;
  assign n28798 = n28786 & n28797 ;
  assign n28799 = \m3_addr_i[27]_pad  & ~n14009 ;
  assign n28800 = n14034 & n28799 ;
  assign n28801 = \m4_addr_i[27]_pad  & n14009 ;
  assign n28802 = n14002 & n28801 ;
  assign n28803 = ~n28800 & ~n28802 ;
  assign n28804 = \m5_addr_i[27]_pad  & ~n14009 ;
  assign n28805 = n14002 & n28804 ;
  assign n28806 = \m7_addr_i[27]_pad  & ~n14009 ;
  assign n28807 = n14026 & n28806 ;
  assign n28808 = ~n28805 & ~n28807 ;
  assign n28809 = n28803 & n28808 ;
  assign n28810 = \m6_addr_i[27]_pad  & n14009 ;
  assign n28811 = n14026 & n28810 ;
  assign n28812 = \m0_addr_i[27]_pad  & n14009 ;
  assign n28813 = n14017 & n28812 ;
  assign n28814 = ~n28811 & ~n28813 ;
  assign n28815 = \m1_addr_i[27]_pad  & ~n14009 ;
  assign n28816 = n14017 & n28815 ;
  assign n28817 = \m2_addr_i[27]_pad  & n14009 ;
  assign n28818 = n14034 & n28817 ;
  assign n28819 = ~n28816 & ~n28818 ;
  assign n28820 = n28814 & n28819 ;
  assign n28821 = n28809 & n28820 ;
  assign n28822 = \m3_addr_i[28]_pad  & ~n14009 ;
  assign n28823 = n14034 & n28822 ;
  assign n28824 = \m4_addr_i[28]_pad  & n14009 ;
  assign n28825 = n14002 & n28824 ;
  assign n28826 = ~n28823 & ~n28825 ;
  assign n28827 = \m5_addr_i[28]_pad  & ~n14009 ;
  assign n28828 = n14002 & n28827 ;
  assign n28829 = \m2_addr_i[28]_pad  & n14009 ;
  assign n28830 = n14034 & n28829 ;
  assign n28831 = ~n28828 & ~n28830 ;
  assign n28832 = n28826 & n28831 ;
  assign n28833 = \m6_addr_i[28]_pad  & n14009 ;
  assign n28834 = n14026 & n28833 ;
  assign n28835 = \m1_addr_i[28]_pad  & ~n14009 ;
  assign n28836 = n14017 & n28835 ;
  assign n28837 = ~n28834 & ~n28836 ;
  assign n28838 = \m0_addr_i[28]_pad  & n14009 ;
  assign n28839 = n14017 & n28838 ;
  assign n28840 = \m7_addr_i[28]_pad  & ~n14009 ;
  assign n28841 = n14026 & n28840 ;
  assign n28842 = ~n28839 & ~n28841 ;
  assign n28843 = n28837 & n28842 ;
  assign n28844 = n28832 & n28843 ;
  assign n28845 = \m5_addr_i[29]_pad  & ~n14009 ;
  assign n28846 = n14002 & n28845 ;
  assign n28847 = \m6_addr_i[29]_pad  & n14009 ;
  assign n28848 = n14026 & n28847 ;
  assign n28849 = ~n28846 & ~n28848 ;
  assign n28850 = \m3_addr_i[29]_pad  & ~n14009 ;
  assign n28851 = n14034 & n28850 ;
  assign n28852 = \m2_addr_i[29]_pad  & n14009 ;
  assign n28853 = n14034 & n28852 ;
  assign n28854 = ~n28851 & ~n28853 ;
  assign n28855 = n28849 & n28854 ;
  assign n28856 = \m4_addr_i[29]_pad  & n14009 ;
  assign n28857 = n14002 & n28856 ;
  assign n28858 = \m1_addr_i[29]_pad  & ~n14009 ;
  assign n28859 = n14017 & n28858 ;
  assign n28860 = ~n28857 & ~n28859 ;
  assign n28861 = \m0_addr_i[29]_pad  & n14009 ;
  assign n28862 = n14017 & n28861 ;
  assign n28863 = \m7_addr_i[29]_pad  & ~n14009 ;
  assign n28864 = n14026 & n28863 ;
  assign n28865 = ~n28862 & ~n28864 ;
  assign n28866 = n28860 & n28865 ;
  assign n28867 = n28855 & n28866 ;
  assign n28868 = \m3_addr_i[2]_pad  & ~n14009 ;
  assign n28869 = n14034 & n28868 ;
  assign n28870 = \m4_addr_i[2]_pad  & n14009 ;
  assign n28871 = n14002 & n28870 ;
  assign n28872 = ~n28869 & ~n28871 ;
  assign n28873 = \m0_addr_i[2]_pad  & n14009 ;
  assign n28874 = n14017 & n28873 ;
  assign n28875 = \m5_addr_i[2]_pad  & ~n14009 ;
  assign n28876 = n14002 & n28875 ;
  assign n28877 = ~n28874 & ~n28876 ;
  assign n28878 = n28872 & n28877 ;
  assign n28879 = \m7_addr_i[2]_pad  & ~n14009 ;
  assign n28880 = n14026 & n28879 ;
  assign n28881 = \m6_addr_i[2]_pad  & n14009 ;
  assign n28882 = n14026 & n28881 ;
  assign n28883 = ~n28880 & ~n28882 ;
  assign n28884 = \m1_addr_i[2]_pad  & ~n14009 ;
  assign n28885 = n14017 & n28884 ;
  assign n28886 = \m2_addr_i[2]_pad  & n14009 ;
  assign n28887 = n14034 & n28886 ;
  assign n28888 = ~n28885 & ~n28887 ;
  assign n28889 = n28883 & n28888 ;
  assign n28890 = n28878 & n28889 ;
  assign n28891 = \m1_addr_i[30]_pad  & ~n14009 ;
  assign n28892 = n14017 & n28891 ;
  assign n28893 = \m2_addr_i[30]_pad  & n14009 ;
  assign n28894 = n14034 & n28893 ;
  assign n28895 = ~n28892 & ~n28894 ;
  assign n28896 = \m0_addr_i[30]_pad  & n14009 ;
  assign n28897 = n14017 & n28896 ;
  assign n28898 = \m6_addr_i[30]_pad  & n14009 ;
  assign n28899 = n14026 & n28898 ;
  assign n28900 = ~n28897 & ~n28899 ;
  assign n28901 = n28895 & n28900 ;
  assign n28902 = \m7_addr_i[30]_pad  & ~n14009 ;
  assign n28903 = n14026 & n28902 ;
  assign n28904 = \m5_addr_i[30]_pad  & ~n14009 ;
  assign n28905 = n14002 & n28904 ;
  assign n28906 = ~n28903 & ~n28905 ;
  assign n28907 = \m3_addr_i[30]_pad  & ~n14009 ;
  assign n28908 = n14034 & n28907 ;
  assign n28909 = \m4_addr_i[30]_pad  & n14009 ;
  assign n28910 = n14002 & n28909 ;
  assign n28911 = ~n28908 & ~n28910 ;
  assign n28912 = n28906 & n28911 ;
  assign n28913 = n28901 & n28912 ;
  assign n28914 = \m0_addr_i[31]_pad  & n14009 ;
  assign n28915 = n14017 & n28914 ;
  assign n28916 = \m7_addr_i[31]_pad  & ~n14009 ;
  assign n28917 = n14026 & n28916 ;
  assign n28918 = ~n28915 & ~n28917 ;
  assign n28919 = \m1_addr_i[31]_pad  & ~n14009 ;
  assign n28920 = n14017 & n28919 ;
  assign n28921 = \m6_addr_i[31]_pad  & n14009 ;
  assign n28922 = n14026 & n28921 ;
  assign n28923 = ~n28920 & ~n28922 ;
  assign n28924 = n28918 & n28923 ;
  assign n28925 = \m2_addr_i[31]_pad  & n14009 ;
  assign n28926 = n14034 & n28925 ;
  assign n28927 = \m5_addr_i[31]_pad  & ~n14009 ;
  assign n28928 = n14002 & n28927 ;
  assign n28929 = ~n28926 & ~n28928 ;
  assign n28930 = \m3_addr_i[31]_pad  & ~n14009 ;
  assign n28931 = n14034 & n28930 ;
  assign n28932 = \m4_addr_i[31]_pad  & n14009 ;
  assign n28933 = n14002 & n28932 ;
  assign n28934 = ~n28931 & ~n28933 ;
  assign n28935 = n28929 & n28934 ;
  assign n28936 = n28924 & n28935 ;
  assign n28937 = \m0_addr_i[3]_pad  & n14009 ;
  assign n28938 = n14017 & n28937 ;
  assign n28939 = \m7_addr_i[3]_pad  & ~n14009 ;
  assign n28940 = n14026 & n28939 ;
  assign n28941 = ~n28938 & ~n28940 ;
  assign n28942 = \m1_addr_i[3]_pad  & ~n14009 ;
  assign n28943 = n14017 & n28942 ;
  assign n28944 = \m4_addr_i[3]_pad  & n14009 ;
  assign n28945 = n14002 & n28944 ;
  assign n28946 = ~n28943 & ~n28945 ;
  assign n28947 = n28941 & n28946 ;
  assign n28948 = \m2_addr_i[3]_pad  & n14009 ;
  assign n28949 = n14034 & n28948 ;
  assign n28950 = \m3_addr_i[3]_pad  & ~n14009 ;
  assign n28951 = n14034 & n28950 ;
  assign n28952 = ~n28949 & ~n28951 ;
  assign n28953 = \m6_addr_i[3]_pad  & n14009 ;
  assign n28954 = n14026 & n28953 ;
  assign n28955 = \m5_addr_i[3]_pad  & ~n14009 ;
  assign n28956 = n14002 & n28955 ;
  assign n28957 = ~n28954 & ~n28956 ;
  assign n28958 = n28952 & n28957 ;
  assign n28959 = n28947 & n28958 ;
  assign n28960 = \m1_addr_i[4]_pad  & ~n14009 ;
  assign n28961 = n14017 & n28960 ;
  assign n28962 = \m2_addr_i[4]_pad  & n14009 ;
  assign n28963 = n14034 & n28962 ;
  assign n28964 = ~n28961 & ~n28963 ;
  assign n28965 = \m6_addr_i[4]_pad  & n14009 ;
  assign n28966 = n14026 & n28965 ;
  assign n28967 = \m7_addr_i[4]_pad  & ~n14009 ;
  assign n28968 = n14026 & n28967 ;
  assign n28969 = ~n28966 & ~n28968 ;
  assign n28970 = n28964 & n28969 ;
  assign n28971 = \m5_addr_i[4]_pad  & ~n14009 ;
  assign n28972 = n14002 & n28971 ;
  assign n28973 = \m0_addr_i[4]_pad  & n14009 ;
  assign n28974 = n14017 & n28973 ;
  assign n28975 = ~n28972 & ~n28974 ;
  assign n28976 = \m3_addr_i[4]_pad  & ~n14009 ;
  assign n28977 = n14034 & n28976 ;
  assign n28978 = \m4_addr_i[4]_pad  & n14009 ;
  assign n28979 = n14002 & n28978 ;
  assign n28980 = ~n28977 & ~n28979 ;
  assign n28981 = n28975 & n28980 ;
  assign n28982 = n28970 & n28981 ;
  assign n28983 = \m3_addr_i[5]_pad  & ~n14009 ;
  assign n28984 = n14034 & n28983 ;
  assign n28985 = \m4_addr_i[5]_pad  & n14009 ;
  assign n28986 = n14002 & n28985 ;
  assign n28987 = ~n28984 & ~n28986 ;
  assign n28988 = \m0_addr_i[5]_pad  & n14009 ;
  assign n28989 = n14017 & n28988 ;
  assign n28990 = \m5_addr_i[5]_pad  & ~n14009 ;
  assign n28991 = n14002 & n28990 ;
  assign n28992 = ~n28989 & ~n28991 ;
  assign n28993 = n28987 & n28992 ;
  assign n28994 = \m7_addr_i[5]_pad  & ~n14009 ;
  assign n28995 = n14026 & n28994 ;
  assign n28996 = \m6_addr_i[5]_pad  & n14009 ;
  assign n28997 = n14026 & n28996 ;
  assign n28998 = ~n28995 & ~n28997 ;
  assign n28999 = \m1_addr_i[5]_pad  & ~n14009 ;
  assign n29000 = n14017 & n28999 ;
  assign n29001 = \m2_addr_i[5]_pad  & n14009 ;
  assign n29002 = n14034 & n29001 ;
  assign n29003 = ~n29000 & ~n29002 ;
  assign n29004 = n28998 & n29003 ;
  assign n29005 = n28993 & n29004 ;
  assign n29006 = \m3_addr_i[6]_pad  & ~n14009 ;
  assign n29007 = n14034 & n29006 ;
  assign n29008 = \m4_addr_i[6]_pad  & n14009 ;
  assign n29009 = n14002 & n29008 ;
  assign n29010 = ~n29007 & ~n29009 ;
  assign n29011 = \m1_addr_i[6]_pad  & ~n14009 ;
  assign n29012 = n14017 & n29011 ;
  assign n29013 = \m7_addr_i[6]_pad  & ~n14009 ;
  assign n29014 = n14026 & n29013 ;
  assign n29015 = ~n29012 & ~n29014 ;
  assign n29016 = n29010 & n29015 ;
  assign n29017 = \m2_addr_i[6]_pad  & n14009 ;
  assign n29018 = n14034 & n29017 ;
  assign n29019 = \m0_addr_i[6]_pad  & n14009 ;
  assign n29020 = n14017 & n29019 ;
  assign n29021 = ~n29018 & ~n29020 ;
  assign n29022 = \m6_addr_i[6]_pad  & n14009 ;
  assign n29023 = n14026 & n29022 ;
  assign n29024 = \m5_addr_i[6]_pad  & ~n14009 ;
  assign n29025 = n14002 & n29024 ;
  assign n29026 = ~n29023 & ~n29025 ;
  assign n29027 = n29021 & n29026 ;
  assign n29028 = n29016 & n29027 ;
  assign n29029 = \m3_addr_i[7]_pad  & ~n14009 ;
  assign n29030 = n14034 & n29029 ;
  assign n29031 = \m4_addr_i[7]_pad  & n14009 ;
  assign n29032 = n14002 & n29031 ;
  assign n29033 = ~n29030 & ~n29032 ;
  assign n29034 = \m6_addr_i[7]_pad  & n14009 ;
  assign n29035 = n14026 & n29034 ;
  assign n29036 = \m2_addr_i[7]_pad  & n14009 ;
  assign n29037 = n14034 & n29036 ;
  assign n29038 = ~n29035 & ~n29037 ;
  assign n29039 = n29033 & n29038 ;
  assign n29040 = \m5_addr_i[7]_pad  & ~n14009 ;
  assign n29041 = n14002 & n29040 ;
  assign n29042 = \m1_addr_i[7]_pad  & ~n14009 ;
  assign n29043 = n14017 & n29042 ;
  assign n29044 = ~n29041 & ~n29043 ;
  assign n29045 = \m0_addr_i[7]_pad  & n14009 ;
  assign n29046 = n14017 & n29045 ;
  assign n29047 = \m7_addr_i[7]_pad  & ~n14009 ;
  assign n29048 = n14026 & n29047 ;
  assign n29049 = ~n29046 & ~n29048 ;
  assign n29050 = n29044 & n29049 ;
  assign n29051 = n29039 & n29050 ;
  assign n29052 = \m6_addr_i[8]_pad  & n14009 ;
  assign n29053 = n14026 & n29052 ;
  assign n29054 = \m5_addr_i[8]_pad  & ~n14009 ;
  assign n29055 = n14002 & n29054 ;
  assign n29056 = ~n29053 & ~n29055 ;
  assign n29057 = \m0_addr_i[8]_pad  & n14009 ;
  assign n29058 = n14017 & n29057 ;
  assign n29059 = \m4_addr_i[8]_pad  & n14009 ;
  assign n29060 = n14002 & n29059 ;
  assign n29061 = ~n29058 & ~n29060 ;
  assign n29062 = n29056 & n29061 ;
  assign n29063 = \m7_addr_i[8]_pad  & ~n14009 ;
  assign n29064 = n14026 & n29063 ;
  assign n29065 = \m3_addr_i[8]_pad  & ~n14009 ;
  assign n29066 = n14034 & n29065 ;
  assign n29067 = ~n29064 & ~n29066 ;
  assign n29068 = \m1_addr_i[8]_pad  & ~n14009 ;
  assign n29069 = n14017 & n29068 ;
  assign n29070 = \m2_addr_i[8]_pad  & n14009 ;
  assign n29071 = n14034 & n29070 ;
  assign n29072 = ~n29069 & ~n29071 ;
  assign n29073 = n29067 & n29072 ;
  assign n29074 = n29062 & n29073 ;
  assign n29075 = \m1_addr_i[9]_pad  & ~n14009 ;
  assign n29076 = n14017 & n29075 ;
  assign n29077 = \m2_addr_i[9]_pad  & n14009 ;
  assign n29078 = n14034 & n29077 ;
  assign n29079 = ~n29076 & ~n29078 ;
  assign n29080 = \m3_addr_i[9]_pad  & ~n14009 ;
  assign n29081 = n14034 & n29080 ;
  assign n29082 = \m5_addr_i[9]_pad  & ~n14009 ;
  assign n29083 = n14002 & n29082 ;
  assign n29084 = ~n29081 & ~n29083 ;
  assign n29085 = n29079 & n29084 ;
  assign n29086 = \m4_addr_i[9]_pad  & n14009 ;
  assign n29087 = n14002 & n29086 ;
  assign n29088 = \m6_addr_i[9]_pad  & n14009 ;
  assign n29089 = n14026 & n29088 ;
  assign n29090 = ~n29087 & ~n29089 ;
  assign n29091 = \m0_addr_i[9]_pad  & n14009 ;
  assign n29092 = n14017 & n29091 ;
  assign n29093 = \m7_addr_i[9]_pad  & ~n14009 ;
  assign n29094 = n14026 & n29093 ;
  assign n29095 = ~n29092 & ~n29094 ;
  assign n29096 = n29090 & n29095 ;
  assign n29097 = n29085 & n29096 ;
  assign n29098 = \m0_data_i[0]_pad  & n14009 ;
  assign n29099 = n14017 & n29098 ;
  assign n29100 = \m7_data_i[0]_pad  & ~n14009 ;
  assign n29101 = n14026 & n29100 ;
  assign n29102 = ~n29099 & ~n29101 ;
  assign n29103 = \m6_data_i[0]_pad  & n14009 ;
  assign n29104 = n14026 & n29103 ;
  assign n29105 = \m2_data_i[0]_pad  & n14009 ;
  assign n29106 = n14034 & n29105 ;
  assign n29107 = ~n29104 & ~n29106 ;
  assign n29108 = n29102 & n29107 ;
  assign n29109 = \m5_data_i[0]_pad  & ~n14009 ;
  assign n29110 = n14002 & n29109 ;
  assign n29111 = \m1_data_i[0]_pad  & ~n14009 ;
  assign n29112 = n14017 & n29111 ;
  assign n29113 = ~n29110 & ~n29112 ;
  assign n29114 = \m3_data_i[0]_pad  & ~n14009 ;
  assign n29115 = n14034 & n29114 ;
  assign n29116 = \m4_data_i[0]_pad  & n14009 ;
  assign n29117 = n14002 & n29116 ;
  assign n29118 = ~n29115 & ~n29117 ;
  assign n29119 = n29113 & n29118 ;
  assign n29120 = n29108 & n29119 ;
  assign n29121 = \m1_data_i[10]_pad  & ~n14009 ;
  assign n29122 = n14017 & n29121 ;
  assign n29123 = \m2_data_i[10]_pad  & n14009 ;
  assign n29124 = n14034 & n29123 ;
  assign n29125 = ~n29122 & ~n29124 ;
  assign n29126 = \m0_data_i[10]_pad  & n14009 ;
  assign n29127 = n14017 & n29126 ;
  assign n29128 = \m4_data_i[10]_pad  & n14009 ;
  assign n29129 = n14002 & n29128 ;
  assign n29130 = ~n29127 & ~n29129 ;
  assign n29131 = n29125 & n29130 ;
  assign n29132 = \m7_data_i[10]_pad  & ~n14009 ;
  assign n29133 = n14026 & n29132 ;
  assign n29134 = \m3_data_i[10]_pad  & ~n14009 ;
  assign n29135 = n14034 & n29134 ;
  assign n29136 = ~n29133 & ~n29135 ;
  assign n29137 = \m6_data_i[10]_pad  & n14009 ;
  assign n29138 = n14026 & n29137 ;
  assign n29139 = \m5_data_i[10]_pad  & ~n14009 ;
  assign n29140 = n14002 & n29139 ;
  assign n29141 = ~n29138 & ~n29140 ;
  assign n29142 = n29136 & n29141 ;
  assign n29143 = n29131 & n29142 ;
  assign n29144 = \m3_data_i[11]_pad  & ~n14009 ;
  assign n29145 = n14034 & n29144 ;
  assign n29146 = \m4_data_i[11]_pad  & n14009 ;
  assign n29147 = n14002 & n29146 ;
  assign n29148 = ~n29145 & ~n29147 ;
  assign n29149 = \m0_data_i[11]_pad  & n14009 ;
  assign n29150 = n14017 & n29149 ;
  assign n29151 = \m2_data_i[11]_pad  & n14009 ;
  assign n29152 = n14034 & n29151 ;
  assign n29153 = ~n29150 & ~n29152 ;
  assign n29154 = n29148 & n29153 ;
  assign n29155 = \m7_data_i[11]_pad  & ~n14009 ;
  assign n29156 = n14026 & n29155 ;
  assign n29157 = \m1_data_i[11]_pad  & ~n14009 ;
  assign n29158 = n14017 & n29157 ;
  assign n29159 = ~n29156 & ~n29158 ;
  assign n29160 = \m6_data_i[11]_pad  & n14009 ;
  assign n29161 = n14026 & n29160 ;
  assign n29162 = \m5_data_i[11]_pad  & ~n14009 ;
  assign n29163 = n14002 & n29162 ;
  assign n29164 = ~n29161 & ~n29163 ;
  assign n29165 = n29159 & n29164 ;
  assign n29166 = n29154 & n29165 ;
  assign n29167 = \m1_data_i[12]_pad  & ~n14009 ;
  assign n29168 = n14017 & n29167 ;
  assign n29169 = \m2_data_i[12]_pad  & n14009 ;
  assign n29170 = n14034 & n29169 ;
  assign n29171 = ~n29168 & ~n29170 ;
  assign n29172 = \m0_data_i[12]_pad  & n14009 ;
  assign n29173 = n14017 & n29172 ;
  assign n29174 = \m4_data_i[12]_pad  & n14009 ;
  assign n29175 = n14002 & n29174 ;
  assign n29176 = ~n29173 & ~n29175 ;
  assign n29177 = n29171 & n29176 ;
  assign n29178 = \m7_data_i[12]_pad  & ~n14009 ;
  assign n29179 = n14026 & n29178 ;
  assign n29180 = \m3_data_i[12]_pad  & ~n14009 ;
  assign n29181 = n14034 & n29180 ;
  assign n29182 = ~n29179 & ~n29181 ;
  assign n29183 = \m6_data_i[12]_pad  & n14009 ;
  assign n29184 = n14026 & n29183 ;
  assign n29185 = \m5_data_i[12]_pad  & ~n14009 ;
  assign n29186 = n14002 & n29185 ;
  assign n29187 = ~n29184 & ~n29186 ;
  assign n29188 = n29182 & n29187 ;
  assign n29189 = n29177 & n29188 ;
  assign n29190 = \m1_data_i[13]_pad  & ~n14009 ;
  assign n29191 = n14017 & n29190 ;
  assign n29192 = \m2_data_i[13]_pad  & n14009 ;
  assign n29193 = n14034 & n29192 ;
  assign n29194 = ~n29191 & ~n29193 ;
  assign n29195 = \m0_data_i[13]_pad  & n14009 ;
  assign n29196 = n14017 & n29195 ;
  assign n29197 = \m5_data_i[13]_pad  & ~n14009 ;
  assign n29198 = n14002 & n29197 ;
  assign n29199 = ~n29196 & ~n29198 ;
  assign n29200 = n29194 & n29199 ;
  assign n29201 = \m7_data_i[13]_pad  & ~n14009 ;
  assign n29202 = n14026 & n29201 ;
  assign n29203 = \m6_data_i[13]_pad  & n14009 ;
  assign n29204 = n14026 & n29203 ;
  assign n29205 = ~n29202 & ~n29204 ;
  assign n29206 = \m3_data_i[13]_pad  & ~n14009 ;
  assign n29207 = n14034 & n29206 ;
  assign n29208 = \m4_data_i[13]_pad  & n14009 ;
  assign n29209 = n14002 & n29208 ;
  assign n29210 = ~n29207 & ~n29209 ;
  assign n29211 = n29205 & n29210 ;
  assign n29212 = n29200 & n29211 ;
  assign n29213 = \m1_data_i[14]_pad  & ~n14009 ;
  assign n29214 = n14017 & n29213 ;
  assign n29215 = \m2_data_i[14]_pad  & n14009 ;
  assign n29216 = n14034 & n29215 ;
  assign n29217 = ~n29214 & ~n29216 ;
  assign n29218 = \m0_data_i[14]_pad  & n14009 ;
  assign n29219 = n14017 & n29218 ;
  assign n29220 = \m5_data_i[14]_pad  & ~n14009 ;
  assign n29221 = n14002 & n29220 ;
  assign n29222 = ~n29219 & ~n29221 ;
  assign n29223 = n29217 & n29222 ;
  assign n29224 = \m7_data_i[14]_pad  & ~n14009 ;
  assign n29225 = n14026 & n29224 ;
  assign n29226 = \m6_data_i[14]_pad  & n14009 ;
  assign n29227 = n14026 & n29226 ;
  assign n29228 = ~n29225 & ~n29227 ;
  assign n29229 = \m3_data_i[14]_pad  & ~n14009 ;
  assign n29230 = n14034 & n29229 ;
  assign n29231 = \m4_data_i[14]_pad  & n14009 ;
  assign n29232 = n14002 & n29231 ;
  assign n29233 = ~n29230 & ~n29232 ;
  assign n29234 = n29228 & n29233 ;
  assign n29235 = n29223 & n29234 ;
  assign n29236 = \m3_data_i[15]_pad  & ~n14009 ;
  assign n29237 = n14034 & n29236 ;
  assign n29238 = \m4_data_i[15]_pad  & n14009 ;
  assign n29239 = n14002 & n29238 ;
  assign n29240 = ~n29237 & ~n29239 ;
  assign n29241 = \m1_data_i[15]_pad  & ~n14009 ;
  assign n29242 = n14017 & n29241 ;
  assign n29243 = \m5_data_i[15]_pad  & ~n14009 ;
  assign n29244 = n14002 & n29243 ;
  assign n29245 = ~n29242 & ~n29244 ;
  assign n29246 = n29240 & n29245 ;
  assign n29247 = \m2_data_i[15]_pad  & n14009 ;
  assign n29248 = n14034 & n29247 ;
  assign n29249 = \m6_data_i[15]_pad  & n14009 ;
  assign n29250 = n14026 & n29249 ;
  assign n29251 = ~n29248 & ~n29250 ;
  assign n29252 = \m0_data_i[15]_pad  & n14009 ;
  assign n29253 = n14017 & n29252 ;
  assign n29254 = \m7_data_i[15]_pad  & ~n14009 ;
  assign n29255 = n14026 & n29254 ;
  assign n29256 = ~n29253 & ~n29255 ;
  assign n29257 = n29251 & n29256 ;
  assign n29258 = n29246 & n29257 ;
  assign n29259 = \m1_data_i[16]_pad  & ~n14009 ;
  assign n29260 = n14017 & n29259 ;
  assign n29261 = \m2_data_i[16]_pad  & n14009 ;
  assign n29262 = n14034 & n29261 ;
  assign n29263 = ~n29260 & ~n29262 ;
  assign n29264 = \m0_data_i[16]_pad  & n14009 ;
  assign n29265 = n14017 & n29264 ;
  assign n29266 = \m4_data_i[16]_pad  & n14009 ;
  assign n29267 = n14002 & n29266 ;
  assign n29268 = ~n29265 & ~n29267 ;
  assign n29269 = n29263 & n29268 ;
  assign n29270 = \m7_data_i[16]_pad  & ~n14009 ;
  assign n29271 = n14026 & n29270 ;
  assign n29272 = \m3_data_i[16]_pad  & ~n14009 ;
  assign n29273 = n14034 & n29272 ;
  assign n29274 = ~n29271 & ~n29273 ;
  assign n29275 = \m6_data_i[16]_pad  & n14009 ;
  assign n29276 = n14026 & n29275 ;
  assign n29277 = \m5_data_i[16]_pad  & ~n14009 ;
  assign n29278 = n14002 & n29277 ;
  assign n29279 = ~n29276 & ~n29278 ;
  assign n29280 = n29274 & n29279 ;
  assign n29281 = n29269 & n29280 ;
  assign n29282 = \m0_data_i[17]_pad  & n14009 ;
  assign n29283 = n14017 & n29282 ;
  assign n29284 = \m7_data_i[17]_pad  & ~n14009 ;
  assign n29285 = n14026 & n29284 ;
  assign n29286 = ~n29283 & ~n29285 ;
  assign n29287 = \m6_data_i[17]_pad  & n14009 ;
  assign n29288 = n14026 & n29287 ;
  assign n29289 = \m2_data_i[17]_pad  & n14009 ;
  assign n29290 = n14034 & n29289 ;
  assign n29291 = ~n29288 & ~n29290 ;
  assign n29292 = n29286 & n29291 ;
  assign n29293 = \m5_data_i[17]_pad  & ~n14009 ;
  assign n29294 = n14002 & n29293 ;
  assign n29295 = \m1_data_i[17]_pad  & ~n14009 ;
  assign n29296 = n14017 & n29295 ;
  assign n29297 = ~n29294 & ~n29296 ;
  assign n29298 = \m3_data_i[17]_pad  & ~n14009 ;
  assign n29299 = n14034 & n29298 ;
  assign n29300 = \m4_data_i[17]_pad  & n14009 ;
  assign n29301 = n14002 & n29300 ;
  assign n29302 = ~n29299 & ~n29301 ;
  assign n29303 = n29297 & n29302 ;
  assign n29304 = n29292 & n29303 ;
  assign n29305 = \m1_data_i[18]_pad  & ~n14009 ;
  assign n29306 = n14017 & n29305 ;
  assign n29307 = \m2_data_i[18]_pad  & n14009 ;
  assign n29308 = n14034 & n29307 ;
  assign n29309 = ~n29306 & ~n29308 ;
  assign n29310 = \m3_data_i[18]_pad  & ~n14009 ;
  assign n29311 = n14034 & n29310 ;
  assign n29312 = \m7_data_i[18]_pad  & ~n14009 ;
  assign n29313 = n14026 & n29312 ;
  assign n29314 = ~n29311 & ~n29313 ;
  assign n29315 = n29309 & n29314 ;
  assign n29316 = \m4_data_i[18]_pad  & n14009 ;
  assign n29317 = n14002 & n29316 ;
  assign n29318 = \m0_data_i[18]_pad  & n14009 ;
  assign n29319 = n14017 & n29318 ;
  assign n29320 = ~n29317 & ~n29319 ;
  assign n29321 = \m6_data_i[18]_pad  & n14009 ;
  assign n29322 = n14026 & n29321 ;
  assign n29323 = \m5_data_i[18]_pad  & ~n14009 ;
  assign n29324 = n14002 & n29323 ;
  assign n29325 = ~n29322 & ~n29324 ;
  assign n29326 = n29320 & n29325 ;
  assign n29327 = n29315 & n29326 ;
  assign n29328 = \m1_data_i[19]_pad  & ~n14009 ;
  assign n29329 = n14017 & n29328 ;
  assign n29330 = \m2_data_i[19]_pad  & n14009 ;
  assign n29331 = n14034 & n29330 ;
  assign n29332 = ~n29329 & ~n29331 ;
  assign n29333 = \m0_data_i[19]_pad  & n14009 ;
  assign n29334 = n14017 & n29333 ;
  assign n29335 = \m5_data_i[19]_pad  & ~n14009 ;
  assign n29336 = n14002 & n29335 ;
  assign n29337 = ~n29334 & ~n29336 ;
  assign n29338 = n29332 & n29337 ;
  assign n29339 = \m7_data_i[19]_pad  & ~n14009 ;
  assign n29340 = n14026 & n29339 ;
  assign n29341 = \m6_data_i[19]_pad  & n14009 ;
  assign n29342 = n14026 & n29341 ;
  assign n29343 = ~n29340 & ~n29342 ;
  assign n29344 = \m3_data_i[19]_pad  & ~n14009 ;
  assign n29345 = n14034 & n29344 ;
  assign n29346 = \m4_data_i[19]_pad  & n14009 ;
  assign n29347 = n14002 & n29346 ;
  assign n29348 = ~n29345 & ~n29347 ;
  assign n29349 = n29343 & n29348 ;
  assign n29350 = n29338 & n29349 ;
  assign n29351 = \m3_data_i[1]_pad  & ~n14009 ;
  assign n29352 = n14034 & n29351 ;
  assign n29353 = \m4_data_i[1]_pad  & n14009 ;
  assign n29354 = n14002 & n29353 ;
  assign n29355 = ~n29352 & ~n29354 ;
  assign n29356 = \m0_data_i[1]_pad  & n14009 ;
  assign n29357 = n14017 & n29356 ;
  assign n29358 = \m2_data_i[1]_pad  & n14009 ;
  assign n29359 = n14034 & n29358 ;
  assign n29360 = ~n29357 & ~n29359 ;
  assign n29361 = n29355 & n29360 ;
  assign n29362 = \m7_data_i[1]_pad  & ~n14009 ;
  assign n29363 = n14026 & n29362 ;
  assign n29364 = \m1_data_i[1]_pad  & ~n14009 ;
  assign n29365 = n14017 & n29364 ;
  assign n29366 = ~n29363 & ~n29365 ;
  assign n29367 = \m6_data_i[1]_pad  & n14009 ;
  assign n29368 = n14026 & n29367 ;
  assign n29369 = \m5_data_i[1]_pad  & ~n14009 ;
  assign n29370 = n14002 & n29369 ;
  assign n29371 = ~n29368 & ~n29370 ;
  assign n29372 = n29366 & n29371 ;
  assign n29373 = n29361 & n29372 ;
  assign n29374 = \m1_data_i[20]_pad  & ~n14009 ;
  assign n29375 = n14017 & n29374 ;
  assign n29376 = \m2_data_i[20]_pad  & n14009 ;
  assign n29377 = n14034 & n29376 ;
  assign n29378 = ~n29375 & ~n29377 ;
  assign n29379 = \m0_data_i[20]_pad  & n14009 ;
  assign n29380 = n14017 & n29379 ;
  assign n29381 = \m4_data_i[20]_pad  & n14009 ;
  assign n29382 = n14002 & n29381 ;
  assign n29383 = ~n29380 & ~n29382 ;
  assign n29384 = n29378 & n29383 ;
  assign n29385 = \m7_data_i[20]_pad  & ~n14009 ;
  assign n29386 = n14026 & n29385 ;
  assign n29387 = \m3_data_i[20]_pad  & ~n14009 ;
  assign n29388 = n14034 & n29387 ;
  assign n29389 = ~n29386 & ~n29388 ;
  assign n29390 = \m6_data_i[20]_pad  & n14009 ;
  assign n29391 = n14026 & n29390 ;
  assign n29392 = \m5_data_i[20]_pad  & ~n14009 ;
  assign n29393 = n14002 & n29392 ;
  assign n29394 = ~n29391 & ~n29393 ;
  assign n29395 = n29389 & n29394 ;
  assign n29396 = n29384 & n29395 ;
  assign n29397 = \m1_data_i[21]_pad  & ~n14009 ;
  assign n29398 = n14017 & n29397 ;
  assign n29399 = \m2_data_i[21]_pad  & n14009 ;
  assign n29400 = n14034 & n29399 ;
  assign n29401 = ~n29398 & ~n29400 ;
  assign n29402 = \m0_data_i[21]_pad  & n14009 ;
  assign n29403 = n14017 & n29402 ;
  assign n29404 = \m4_data_i[21]_pad  & n14009 ;
  assign n29405 = n14002 & n29404 ;
  assign n29406 = ~n29403 & ~n29405 ;
  assign n29407 = n29401 & n29406 ;
  assign n29408 = \m7_data_i[21]_pad  & ~n14009 ;
  assign n29409 = n14026 & n29408 ;
  assign n29410 = \m3_data_i[21]_pad  & ~n14009 ;
  assign n29411 = n14034 & n29410 ;
  assign n29412 = ~n29409 & ~n29411 ;
  assign n29413 = \m6_data_i[21]_pad  & n14009 ;
  assign n29414 = n14026 & n29413 ;
  assign n29415 = \m5_data_i[21]_pad  & ~n14009 ;
  assign n29416 = n14002 & n29415 ;
  assign n29417 = ~n29414 & ~n29416 ;
  assign n29418 = n29412 & n29417 ;
  assign n29419 = n29407 & n29418 ;
  assign n29420 = \m1_data_i[22]_pad  & ~n14009 ;
  assign n29421 = n14017 & n29420 ;
  assign n29422 = \m2_data_i[22]_pad  & n14009 ;
  assign n29423 = n14034 & n29422 ;
  assign n29424 = ~n29421 & ~n29423 ;
  assign n29425 = \m0_data_i[22]_pad  & n14009 ;
  assign n29426 = n14017 & n29425 ;
  assign n29427 = \m4_data_i[22]_pad  & n14009 ;
  assign n29428 = n14002 & n29427 ;
  assign n29429 = ~n29426 & ~n29428 ;
  assign n29430 = n29424 & n29429 ;
  assign n29431 = \m7_data_i[22]_pad  & ~n14009 ;
  assign n29432 = n14026 & n29431 ;
  assign n29433 = \m3_data_i[22]_pad  & ~n14009 ;
  assign n29434 = n14034 & n29433 ;
  assign n29435 = ~n29432 & ~n29434 ;
  assign n29436 = \m6_data_i[22]_pad  & n14009 ;
  assign n29437 = n14026 & n29436 ;
  assign n29438 = \m5_data_i[22]_pad  & ~n14009 ;
  assign n29439 = n14002 & n29438 ;
  assign n29440 = ~n29437 & ~n29439 ;
  assign n29441 = n29435 & n29440 ;
  assign n29442 = n29430 & n29441 ;
  assign n29443 = \m1_data_i[23]_pad  & ~n14009 ;
  assign n29444 = n14017 & n29443 ;
  assign n29445 = \m2_data_i[23]_pad  & n14009 ;
  assign n29446 = n14034 & n29445 ;
  assign n29447 = ~n29444 & ~n29446 ;
  assign n29448 = \m0_data_i[23]_pad  & n14009 ;
  assign n29449 = n14017 & n29448 ;
  assign n29450 = \m4_data_i[23]_pad  & n14009 ;
  assign n29451 = n14002 & n29450 ;
  assign n29452 = ~n29449 & ~n29451 ;
  assign n29453 = n29447 & n29452 ;
  assign n29454 = \m7_data_i[23]_pad  & ~n14009 ;
  assign n29455 = n14026 & n29454 ;
  assign n29456 = \m3_data_i[23]_pad  & ~n14009 ;
  assign n29457 = n14034 & n29456 ;
  assign n29458 = ~n29455 & ~n29457 ;
  assign n29459 = \m6_data_i[23]_pad  & n14009 ;
  assign n29460 = n14026 & n29459 ;
  assign n29461 = \m5_data_i[23]_pad  & ~n14009 ;
  assign n29462 = n14002 & n29461 ;
  assign n29463 = ~n29460 & ~n29462 ;
  assign n29464 = n29458 & n29463 ;
  assign n29465 = n29453 & n29464 ;
  assign n29466 = \m6_data_i[24]_pad  & n14009 ;
  assign n29467 = n14026 & n29466 ;
  assign n29468 = \m5_data_i[24]_pad  & ~n14009 ;
  assign n29469 = n14002 & n29468 ;
  assign n29470 = ~n29467 & ~n29469 ;
  assign n29471 = \m1_data_i[24]_pad  & ~n14009 ;
  assign n29472 = n14017 & n29471 ;
  assign n29473 = \m4_data_i[24]_pad  & n14009 ;
  assign n29474 = n14002 & n29473 ;
  assign n29475 = ~n29472 & ~n29474 ;
  assign n29476 = n29470 & n29475 ;
  assign n29477 = \m2_data_i[24]_pad  & n14009 ;
  assign n29478 = n14034 & n29477 ;
  assign n29479 = \m3_data_i[24]_pad  & ~n14009 ;
  assign n29480 = n14034 & n29479 ;
  assign n29481 = ~n29478 & ~n29480 ;
  assign n29482 = \m0_data_i[24]_pad  & n14009 ;
  assign n29483 = n14017 & n29482 ;
  assign n29484 = \m7_data_i[24]_pad  & ~n14009 ;
  assign n29485 = n14026 & n29484 ;
  assign n29486 = ~n29483 & ~n29485 ;
  assign n29487 = n29481 & n29486 ;
  assign n29488 = n29476 & n29487 ;
  assign n29489 = \m1_data_i[25]_pad  & ~n14009 ;
  assign n29490 = n14017 & n29489 ;
  assign n29491 = \m2_data_i[25]_pad  & n14009 ;
  assign n29492 = n14034 & n29491 ;
  assign n29493 = ~n29490 & ~n29492 ;
  assign n29494 = \m0_data_i[25]_pad  & n14009 ;
  assign n29495 = n14017 & n29494 ;
  assign n29496 = \m4_data_i[25]_pad  & n14009 ;
  assign n29497 = n14002 & n29496 ;
  assign n29498 = ~n29495 & ~n29497 ;
  assign n29499 = n29493 & n29498 ;
  assign n29500 = \m7_data_i[25]_pad  & ~n14009 ;
  assign n29501 = n14026 & n29500 ;
  assign n29502 = \m3_data_i[25]_pad  & ~n14009 ;
  assign n29503 = n14034 & n29502 ;
  assign n29504 = ~n29501 & ~n29503 ;
  assign n29505 = \m6_data_i[25]_pad  & n14009 ;
  assign n29506 = n14026 & n29505 ;
  assign n29507 = \m5_data_i[25]_pad  & ~n14009 ;
  assign n29508 = n14002 & n29507 ;
  assign n29509 = ~n29506 & ~n29508 ;
  assign n29510 = n29504 & n29509 ;
  assign n29511 = n29499 & n29510 ;
  assign n29512 = \m0_data_i[26]_pad  & n14009 ;
  assign n29513 = n14017 & n29512 ;
  assign n29514 = \m7_data_i[26]_pad  & ~n14009 ;
  assign n29515 = n14026 & n29514 ;
  assign n29516 = ~n29513 & ~n29515 ;
  assign n29517 = \m1_data_i[26]_pad  & ~n14009 ;
  assign n29518 = n14017 & n29517 ;
  assign n29519 = \m4_data_i[26]_pad  & n14009 ;
  assign n29520 = n14002 & n29519 ;
  assign n29521 = ~n29518 & ~n29520 ;
  assign n29522 = n29516 & n29521 ;
  assign n29523 = \m2_data_i[26]_pad  & n14009 ;
  assign n29524 = n14034 & n29523 ;
  assign n29525 = \m3_data_i[26]_pad  & ~n14009 ;
  assign n29526 = n14034 & n29525 ;
  assign n29527 = ~n29524 & ~n29526 ;
  assign n29528 = \m6_data_i[26]_pad  & n14009 ;
  assign n29529 = n14026 & n29528 ;
  assign n29530 = \m5_data_i[26]_pad  & ~n14009 ;
  assign n29531 = n14002 & n29530 ;
  assign n29532 = ~n29529 & ~n29531 ;
  assign n29533 = n29527 & n29532 ;
  assign n29534 = n29522 & n29533 ;
  assign n29535 = \m0_data_i[27]_pad  & n14009 ;
  assign n29536 = n14017 & n29535 ;
  assign n29537 = \m7_data_i[27]_pad  & ~n14009 ;
  assign n29538 = n14026 & n29537 ;
  assign n29539 = ~n29536 & ~n29538 ;
  assign n29540 = \m1_data_i[27]_pad  & ~n14009 ;
  assign n29541 = n14017 & n29540 ;
  assign n29542 = \m4_data_i[27]_pad  & n14009 ;
  assign n29543 = n14002 & n29542 ;
  assign n29544 = ~n29541 & ~n29543 ;
  assign n29545 = n29539 & n29544 ;
  assign n29546 = \m2_data_i[27]_pad  & n14009 ;
  assign n29547 = n14034 & n29546 ;
  assign n29548 = \m3_data_i[27]_pad  & ~n14009 ;
  assign n29549 = n14034 & n29548 ;
  assign n29550 = ~n29547 & ~n29549 ;
  assign n29551 = \m6_data_i[27]_pad  & n14009 ;
  assign n29552 = n14026 & n29551 ;
  assign n29553 = \m5_data_i[27]_pad  & ~n14009 ;
  assign n29554 = n14002 & n29553 ;
  assign n29555 = ~n29552 & ~n29554 ;
  assign n29556 = n29550 & n29555 ;
  assign n29557 = n29545 & n29556 ;
  assign n29558 = \m1_data_i[28]_pad  & ~n14009 ;
  assign n29559 = n14017 & n29558 ;
  assign n29560 = \m2_data_i[28]_pad  & n14009 ;
  assign n29561 = n14034 & n29560 ;
  assign n29562 = ~n29559 & ~n29561 ;
  assign n29563 = \m0_data_i[28]_pad  & n14009 ;
  assign n29564 = n14017 & n29563 ;
  assign n29565 = \m4_data_i[28]_pad  & n14009 ;
  assign n29566 = n14002 & n29565 ;
  assign n29567 = ~n29564 & ~n29566 ;
  assign n29568 = n29562 & n29567 ;
  assign n29569 = \m7_data_i[28]_pad  & ~n14009 ;
  assign n29570 = n14026 & n29569 ;
  assign n29571 = \m3_data_i[28]_pad  & ~n14009 ;
  assign n29572 = n14034 & n29571 ;
  assign n29573 = ~n29570 & ~n29572 ;
  assign n29574 = \m6_data_i[28]_pad  & n14009 ;
  assign n29575 = n14026 & n29574 ;
  assign n29576 = \m5_data_i[28]_pad  & ~n14009 ;
  assign n29577 = n14002 & n29576 ;
  assign n29578 = ~n29575 & ~n29577 ;
  assign n29579 = n29573 & n29578 ;
  assign n29580 = n29568 & n29579 ;
  assign n29581 = \m1_data_i[29]_pad  & ~n14009 ;
  assign n29582 = n14017 & n29581 ;
  assign n29583 = \m2_data_i[29]_pad  & n14009 ;
  assign n29584 = n14034 & n29583 ;
  assign n29585 = ~n29582 & ~n29584 ;
  assign n29586 = \m0_data_i[29]_pad  & n14009 ;
  assign n29587 = n14017 & n29586 ;
  assign n29588 = \m4_data_i[29]_pad  & n14009 ;
  assign n29589 = n14002 & n29588 ;
  assign n29590 = ~n29587 & ~n29589 ;
  assign n29591 = n29585 & n29590 ;
  assign n29592 = \m7_data_i[29]_pad  & ~n14009 ;
  assign n29593 = n14026 & n29592 ;
  assign n29594 = \m3_data_i[29]_pad  & ~n14009 ;
  assign n29595 = n14034 & n29594 ;
  assign n29596 = ~n29593 & ~n29595 ;
  assign n29597 = \m6_data_i[29]_pad  & n14009 ;
  assign n29598 = n14026 & n29597 ;
  assign n29599 = \m5_data_i[29]_pad  & ~n14009 ;
  assign n29600 = n14002 & n29599 ;
  assign n29601 = ~n29598 & ~n29600 ;
  assign n29602 = n29596 & n29601 ;
  assign n29603 = n29591 & n29602 ;
  assign n29604 = \m1_data_i[2]_pad  & ~n14009 ;
  assign n29605 = n14017 & n29604 ;
  assign n29606 = \m2_data_i[2]_pad  & n14009 ;
  assign n29607 = n14034 & n29606 ;
  assign n29608 = ~n29605 & ~n29607 ;
  assign n29609 = \m0_data_i[2]_pad  & n14009 ;
  assign n29610 = n14017 & n29609 ;
  assign n29611 = \m5_data_i[2]_pad  & ~n14009 ;
  assign n29612 = n14002 & n29611 ;
  assign n29613 = ~n29610 & ~n29612 ;
  assign n29614 = n29608 & n29613 ;
  assign n29615 = \m7_data_i[2]_pad  & ~n14009 ;
  assign n29616 = n14026 & n29615 ;
  assign n29617 = \m6_data_i[2]_pad  & n14009 ;
  assign n29618 = n14026 & n29617 ;
  assign n29619 = ~n29616 & ~n29618 ;
  assign n29620 = \m3_data_i[2]_pad  & ~n14009 ;
  assign n29621 = n14034 & n29620 ;
  assign n29622 = \m4_data_i[2]_pad  & n14009 ;
  assign n29623 = n14002 & n29622 ;
  assign n29624 = ~n29621 & ~n29623 ;
  assign n29625 = n29619 & n29624 ;
  assign n29626 = n29614 & n29625 ;
  assign n29627 = \m1_data_i[30]_pad  & ~n14009 ;
  assign n29628 = n14017 & n29627 ;
  assign n29629 = \m2_data_i[30]_pad  & n14009 ;
  assign n29630 = n14034 & n29629 ;
  assign n29631 = ~n29628 & ~n29630 ;
  assign n29632 = \m0_data_i[30]_pad  & n14009 ;
  assign n29633 = n14017 & n29632 ;
  assign n29634 = \m4_data_i[30]_pad  & n14009 ;
  assign n29635 = n14002 & n29634 ;
  assign n29636 = ~n29633 & ~n29635 ;
  assign n29637 = n29631 & n29636 ;
  assign n29638 = \m7_data_i[30]_pad  & ~n14009 ;
  assign n29639 = n14026 & n29638 ;
  assign n29640 = \m3_data_i[30]_pad  & ~n14009 ;
  assign n29641 = n14034 & n29640 ;
  assign n29642 = ~n29639 & ~n29641 ;
  assign n29643 = \m6_data_i[30]_pad  & n14009 ;
  assign n29644 = n14026 & n29643 ;
  assign n29645 = \m5_data_i[30]_pad  & ~n14009 ;
  assign n29646 = n14002 & n29645 ;
  assign n29647 = ~n29644 & ~n29646 ;
  assign n29648 = n29642 & n29647 ;
  assign n29649 = n29637 & n29648 ;
  assign n29650 = \m1_data_i[31]_pad  & ~n14009 ;
  assign n29651 = n14017 & n29650 ;
  assign n29652 = \m2_data_i[31]_pad  & n14009 ;
  assign n29653 = n14034 & n29652 ;
  assign n29654 = ~n29651 & ~n29653 ;
  assign n29655 = \m0_data_i[31]_pad  & n14009 ;
  assign n29656 = n14017 & n29655 ;
  assign n29657 = \m5_data_i[31]_pad  & ~n14009 ;
  assign n29658 = n14002 & n29657 ;
  assign n29659 = ~n29656 & ~n29658 ;
  assign n29660 = n29654 & n29659 ;
  assign n29661 = \m7_data_i[31]_pad  & ~n14009 ;
  assign n29662 = n14026 & n29661 ;
  assign n29663 = \m6_data_i[31]_pad  & n14009 ;
  assign n29664 = n14026 & n29663 ;
  assign n29665 = ~n29662 & ~n29664 ;
  assign n29666 = \m3_data_i[31]_pad  & ~n14009 ;
  assign n29667 = n14034 & n29666 ;
  assign n29668 = \m4_data_i[31]_pad  & n14009 ;
  assign n29669 = n14002 & n29668 ;
  assign n29670 = ~n29667 & ~n29669 ;
  assign n29671 = n29665 & n29670 ;
  assign n29672 = n29660 & n29671 ;
  assign n29673 = \m0_data_i[3]_pad  & n14009 ;
  assign n29674 = n14017 & n29673 ;
  assign n29675 = \m7_data_i[3]_pad  & ~n14009 ;
  assign n29676 = n14026 & n29675 ;
  assign n29677 = ~n29674 & ~n29676 ;
  assign n29678 = \m1_data_i[3]_pad  & ~n14009 ;
  assign n29679 = n14017 & n29678 ;
  assign n29680 = \m5_data_i[3]_pad  & ~n14009 ;
  assign n29681 = n14002 & n29680 ;
  assign n29682 = ~n29679 & ~n29681 ;
  assign n29683 = n29677 & n29682 ;
  assign n29684 = \m2_data_i[3]_pad  & n14009 ;
  assign n29685 = n14034 & n29684 ;
  assign n29686 = \m6_data_i[3]_pad  & n14009 ;
  assign n29687 = n14026 & n29686 ;
  assign n29688 = ~n29685 & ~n29687 ;
  assign n29689 = \m3_data_i[3]_pad  & ~n14009 ;
  assign n29690 = n14034 & n29689 ;
  assign n29691 = \m4_data_i[3]_pad  & n14009 ;
  assign n29692 = n14002 & n29691 ;
  assign n29693 = ~n29690 & ~n29692 ;
  assign n29694 = n29688 & n29693 ;
  assign n29695 = n29683 & n29694 ;
  assign n29696 = \m1_data_i[4]_pad  & ~n14009 ;
  assign n29697 = n14017 & n29696 ;
  assign n29698 = \m2_data_i[4]_pad  & n14009 ;
  assign n29699 = n14034 & n29698 ;
  assign n29700 = ~n29697 & ~n29699 ;
  assign n29701 = \m0_data_i[4]_pad  & n14009 ;
  assign n29702 = n14017 & n29701 ;
  assign n29703 = \m4_data_i[4]_pad  & n14009 ;
  assign n29704 = n14002 & n29703 ;
  assign n29705 = ~n29702 & ~n29704 ;
  assign n29706 = n29700 & n29705 ;
  assign n29707 = \m7_data_i[4]_pad  & ~n14009 ;
  assign n29708 = n14026 & n29707 ;
  assign n29709 = \m3_data_i[4]_pad  & ~n14009 ;
  assign n29710 = n14034 & n29709 ;
  assign n29711 = ~n29708 & ~n29710 ;
  assign n29712 = \m6_data_i[4]_pad  & n14009 ;
  assign n29713 = n14026 & n29712 ;
  assign n29714 = \m5_data_i[4]_pad  & ~n14009 ;
  assign n29715 = n14002 & n29714 ;
  assign n29716 = ~n29713 & ~n29715 ;
  assign n29717 = n29711 & n29716 ;
  assign n29718 = n29706 & n29717 ;
  assign n29719 = \m1_data_i[5]_pad  & ~n14009 ;
  assign n29720 = n14017 & n29719 ;
  assign n29721 = \m2_data_i[5]_pad  & n14009 ;
  assign n29722 = n14034 & n29721 ;
  assign n29723 = ~n29720 & ~n29722 ;
  assign n29724 = \m0_data_i[5]_pad  & n14009 ;
  assign n29725 = n14017 & n29724 ;
  assign n29726 = \m5_data_i[5]_pad  & ~n14009 ;
  assign n29727 = n14002 & n29726 ;
  assign n29728 = ~n29725 & ~n29727 ;
  assign n29729 = n29723 & n29728 ;
  assign n29730 = \m7_data_i[5]_pad  & ~n14009 ;
  assign n29731 = n14026 & n29730 ;
  assign n29732 = \m6_data_i[5]_pad  & n14009 ;
  assign n29733 = n14026 & n29732 ;
  assign n29734 = ~n29731 & ~n29733 ;
  assign n29735 = \m3_data_i[5]_pad  & ~n14009 ;
  assign n29736 = n14034 & n29735 ;
  assign n29737 = \m4_data_i[5]_pad  & n14009 ;
  assign n29738 = n14002 & n29737 ;
  assign n29739 = ~n29736 & ~n29738 ;
  assign n29740 = n29734 & n29739 ;
  assign n29741 = n29729 & n29740 ;
  assign n29742 = \m3_data_i[6]_pad  & ~n14009 ;
  assign n29743 = n14034 & n29742 ;
  assign n29744 = \m4_data_i[6]_pad  & n14009 ;
  assign n29745 = n14002 & n29744 ;
  assign n29746 = ~n29743 & ~n29745 ;
  assign n29747 = \m1_data_i[6]_pad  & ~n14009 ;
  assign n29748 = n14017 & n29747 ;
  assign n29749 = \m5_data_i[6]_pad  & ~n14009 ;
  assign n29750 = n14002 & n29749 ;
  assign n29751 = ~n29748 & ~n29750 ;
  assign n29752 = n29746 & n29751 ;
  assign n29753 = \m2_data_i[6]_pad  & n14009 ;
  assign n29754 = n14034 & n29753 ;
  assign n29755 = \m6_data_i[6]_pad  & n14009 ;
  assign n29756 = n14026 & n29755 ;
  assign n29757 = ~n29754 & ~n29756 ;
  assign n29758 = \m0_data_i[6]_pad  & n14009 ;
  assign n29759 = n14017 & n29758 ;
  assign n29760 = \m7_data_i[6]_pad  & ~n14009 ;
  assign n29761 = n14026 & n29760 ;
  assign n29762 = ~n29759 & ~n29761 ;
  assign n29763 = n29757 & n29762 ;
  assign n29764 = n29752 & n29763 ;
  assign n29765 = \m3_data_i[7]_pad  & ~n14009 ;
  assign n29766 = n14034 & n29765 ;
  assign n29767 = \m4_data_i[7]_pad  & n14009 ;
  assign n29768 = n14002 & n29767 ;
  assign n29769 = ~n29766 & ~n29768 ;
  assign n29770 = \m0_data_i[7]_pad  & n14009 ;
  assign n29771 = n14017 & n29770 ;
  assign n29772 = \m2_data_i[7]_pad  & n14009 ;
  assign n29773 = n14034 & n29772 ;
  assign n29774 = ~n29771 & ~n29773 ;
  assign n29775 = n29769 & n29774 ;
  assign n29776 = \m7_data_i[7]_pad  & ~n14009 ;
  assign n29777 = n14026 & n29776 ;
  assign n29778 = \m1_data_i[7]_pad  & ~n14009 ;
  assign n29779 = n14017 & n29778 ;
  assign n29780 = ~n29777 & ~n29779 ;
  assign n29781 = \m6_data_i[7]_pad  & n14009 ;
  assign n29782 = n14026 & n29781 ;
  assign n29783 = \m5_data_i[7]_pad  & ~n14009 ;
  assign n29784 = n14002 & n29783 ;
  assign n29785 = ~n29782 & ~n29784 ;
  assign n29786 = n29780 & n29785 ;
  assign n29787 = n29775 & n29786 ;
  assign n29788 = \m3_data_i[8]_pad  & ~n14009 ;
  assign n29789 = n14034 & n29788 ;
  assign n29790 = \m4_data_i[8]_pad  & n14009 ;
  assign n29791 = n14002 & n29790 ;
  assign n29792 = ~n29789 & ~n29791 ;
  assign n29793 = \m1_data_i[8]_pad  & ~n14009 ;
  assign n29794 = n14017 & n29793 ;
  assign n29795 = \m7_data_i[8]_pad  & ~n14009 ;
  assign n29796 = n14026 & n29795 ;
  assign n29797 = ~n29794 & ~n29796 ;
  assign n29798 = n29792 & n29797 ;
  assign n29799 = \m2_data_i[8]_pad  & n14009 ;
  assign n29800 = n14034 & n29799 ;
  assign n29801 = \m0_data_i[8]_pad  & n14009 ;
  assign n29802 = n14017 & n29801 ;
  assign n29803 = ~n29800 & ~n29802 ;
  assign n29804 = \m6_data_i[8]_pad  & n14009 ;
  assign n29805 = n14026 & n29804 ;
  assign n29806 = \m5_data_i[8]_pad  & ~n14009 ;
  assign n29807 = n14002 & n29806 ;
  assign n29808 = ~n29805 & ~n29807 ;
  assign n29809 = n29803 & n29808 ;
  assign n29810 = n29798 & n29809 ;
  assign n29811 = \m1_data_i[9]_pad  & ~n14009 ;
  assign n29812 = n14017 & n29811 ;
  assign n29813 = \m2_data_i[9]_pad  & n14009 ;
  assign n29814 = n14034 & n29813 ;
  assign n29815 = ~n29812 & ~n29814 ;
  assign n29816 = \m0_data_i[9]_pad  & n14009 ;
  assign n29817 = n14017 & n29816 ;
  assign n29818 = \m5_data_i[9]_pad  & ~n14009 ;
  assign n29819 = n14002 & n29818 ;
  assign n29820 = ~n29817 & ~n29819 ;
  assign n29821 = n29815 & n29820 ;
  assign n29822 = \m7_data_i[9]_pad  & ~n14009 ;
  assign n29823 = n14026 & n29822 ;
  assign n29824 = \m6_data_i[9]_pad  & n14009 ;
  assign n29825 = n14026 & n29824 ;
  assign n29826 = ~n29823 & ~n29825 ;
  assign n29827 = \m3_data_i[9]_pad  & ~n14009 ;
  assign n29828 = n14034 & n29827 ;
  assign n29829 = \m4_data_i[9]_pad  & n14009 ;
  assign n29830 = n14002 & n29829 ;
  assign n29831 = ~n29828 & ~n29830 ;
  assign n29832 = n29826 & n29831 ;
  assign n29833 = n29821 & n29832 ;
  assign n29834 = \m6_sel_i[0]_pad  & n14009 ;
  assign n29835 = n14026 & n29834 ;
  assign n29836 = \m5_sel_i[0]_pad  & ~n14009 ;
  assign n29837 = n14002 & n29836 ;
  assign n29838 = ~n29835 & ~n29837 ;
  assign n29839 = \m0_sel_i[0]_pad  & n14009 ;
  assign n29840 = n14017 & n29839 ;
  assign n29841 = \m4_sel_i[0]_pad  & n14009 ;
  assign n29842 = n14002 & n29841 ;
  assign n29843 = ~n29840 & ~n29842 ;
  assign n29844 = n29838 & n29843 ;
  assign n29845 = \m7_sel_i[0]_pad  & ~n14009 ;
  assign n29846 = n14026 & n29845 ;
  assign n29847 = \m3_sel_i[0]_pad  & ~n14009 ;
  assign n29848 = n14034 & n29847 ;
  assign n29849 = ~n29846 & ~n29848 ;
  assign n29850 = \m1_sel_i[0]_pad  & ~n14009 ;
  assign n29851 = n14017 & n29850 ;
  assign n29852 = \m2_sel_i[0]_pad  & n14009 ;
  assign n29853 = n14034 & n29852 ;
  assign n29854 = ~n29851 & ~n29853 ;
  assign n29855 = n29849 & n29854 ;
  assign n29856 = n29844 & n29855 ;
  assign n29857 = \m0_sel_i[1]_pad  & n14009 ;
  assign n29858 = n14017 & n29857 ;
  assign n29859 = \m7_sel_i[1]_pad  & ~n14009 ;
  assign n29860 = n14026 & n29859 ;
  assign n29861 = ~n29858 & ~n29860 ;
  assign n29862 = \m1_sel_i[1]_pad  & ~n14009 ;
  assign n29863 = n14017 & n29862 ;
  assign n29864 = \m4_sel_i[1]_pad  & n14009 ;
  assign n29865 = n14002 & n29864 ;
  assign n29866 = ~n29863 & ~n29865 ;
  assign n29867 = n29861 & n29866 ;
  assign n29868 = \m2_sel_i[1]_pad  & n14009 ;
  assign n29869 = n14034 & n29868 ;
  assign n29870 = \m3_sel_i[1]_pad  & ~n14009 ;
  assign n29871 = n14034 & n29870 ;
  assign n29872 = ~n29869 & ~n29871 ;
  assign n29873 = \m6_sel_i[1]_pad  & n14009 ;
  assign n29874 = n14026 & n29873 ;
  assign n29875 = \m5_sel_i[1]_pad  & ~n14009 ;
  assign n29876 = n14002 & n29875 ;
  assign n29877 = ~n29874 & ~n29876 ;
  assign n29878 = n29872 & n29877 ;
  assign n29879 = n29867 & n29878 ;
  assign n29880 = \m3_sel_i[2]_pad  & ~n14009 ;
  assign n29881 = n14034 & n29880 ;
  assign n29882 = \m4_sel_i[2]_pad  & n14009 ;
  assign n29883 = n14002 & n29882 ;
  assign n29884 = ~n29881 & ~n29883 ;
  assign n29885 = \m0_sel_i[2]_pad  & n14009 ;
  assign n29886 = n14017 & n29885 ;
  assign n29887 = \m2_sel_i[2]_pad  & n14009 ;
  assign n29888 = n14034 & n29887 ;
  assign n29889 = ~n29886 & ~n29888 ;
  assign n29890 = n29884 & n29889 ;
  assign n29891 = \m7_sel_i[2]_pad  & ~n14009 ;
  assign n29892 = n14026 & n29891 ;
  assign n29893 = \m1_sel_i[2]_pad  & ~n14009 ;
  assign n29894 = n14017 & n29893 ;
  assign n29895 = ~n29892 & ~n29894 ;
  assign n29896 = \m6_sel_i[2]_pad  & n14009 ;
  assign n29897 = n14026 & n29896 ;
  assign n29898 = \m5_sel_i[2]_pad  & ~n14009 ;
  assign n29899 = n14002 & n29898 ;
  assign n29900 = ~n29897 & ~n29899 ;
  assign n29901 = n29895 & n29900 ;
  assign n29902 = n29890 & n29901 ;
  assign n29903 = \m3_sel_i[3]_pad  & ~n14009 ;
  assign n29904 = n14034 & n29903 ;
  assign n29905 = \m4_sel_i[3]_pad  & n14009 ;
  assign n29906 = n14002 & n29905 ;
  assign n29907 = ~n29904 & ~n29906 ;
  assign n29908 = \m1_sel_i[3]_pad  & ~n14009 ;
  assign n29909 = n14017 & n29908 ;
  assign n29910 = \m5_sel_i[3]_pad  & ~n14009 ;
  assign n29911 = n14002 & n29910 ;
  assign n29912 = ~n29909 & ~n29911 ;
  assign n29913 = n29907 & n29912 ;
  assign n29914 = \m2_sel_i[3]_pad  & n14009 ;
  assign n29915 = n14034 & n29914 ;
  assign n29916 = \m6_sel_i[3]_pad  & n14009 ;
  assign n29917 = n14026 & n29916 ;
  assign n29918 = ~n29915 & ~n29917 ;
  assign n29919 = \m0_sel_i[3]_pad  & n14009 ;
  assign n29920 = n14017 & n29919 ;
  assign n29921 = \m7_sel_i[3]_pad  & ~n14009 ;
  assign n29922 = n14026 & n29921 ;
  assign n29923 = ~n29920 & ~n29922 ;
  assign n29924 = n29918 & n29923 ;
  assign n29925 = n29913 & n29924 ;
  assign n29926 = \m3_stb_i_pad  & n14896 ;
  assign n29927 = ~n14009 & n29926 ;
  assign n29928 = n14034 & n29927 ;
  assign n29929 = \m1_stb_i_pad  & n15106 ;
  assign n29930 = ~n14009 & n29929 ;
  assign n29931 = n14017 & n29930 ;
  assign n29932 = ~n29928 & ~n29931 ;
  assign n29933 = \m4_stb_i_pad  & n14735 ;
  assign n29934 = n14009 & n29933 ;
  assign n29935 = n14002 & n29934 ;
  assign n29936 = \m5_stb_i_pad  & n14967 ;
  assign n29937 = ~n14009 & n29936 ;
  assign n29938 = n14002 & n29937 ;
  assign n29939 = ~n29935 & ~n29938 ;
  assign n29940 = n29932 & n29939 ;
  assign n29941 = \m2_stb_i_pad  & n14855 ;
  assign n29942 = n14009 & n29941 ;
  assign n29943 = n14034 & n29942 ;
  assign n29944 = \m7_stb_i_pad  & n15051 ;
  assign n29945 = ~n14009 & n29944 ;
  assign n29946 = n14026 & n29945 ;
  assign n29947 = ~n29943 & ~n29946 ;
  assign n29948 = \m6_stb_i_pad  & n15003 ;
  assign n29949 = n14009 & n29948 ;
  assign n29950 = n14026 & n29949 ;
  assign n29951 = \m0_stb_i_pad  & n14753 ;
  assign n29952 = n14009 & n29951 ;
  assign n29953 = n14017 & n29952 ;
  assign n29954 = ~n29950 & ~n29953 ;
  assign n29955 = n29947 & n29954 ;
  assign n29956 = n29940 & n29955 ;
  assign n29957 = \m6_we_i_pad  & n14009 ;
  assign n29958 = n14026 & n29957 ;
  assign n29959 = \m5_we_i_pad  & ~n14009 ;
  assign n29960 = n14002 & n29959 ;
  assign n29961 = ~n29958 & ~n29960 ;
  assign n29962 = \m3_we_i_pad  & ~n14009 ;
  assign n29963 = n14034 & n29962 ;
  assign n29964 = \m7_we_i_pad  & ~n14009 ;
  assign n29965 = n14026 & n29964 ;
  assign n29966 = ~n29963 & ~n29965 ;
  assign n29967 = n29961 & n29966 ;
  assign n29968 = \m4_we_i_pad  & n14009 ;
  assign n29969 = n14002 & n29968 ;
  assign n29970 = \m0_we_i_pad  & n14009 ;
  assign n29971 = n14017 & n29970 ;
  assign n29972 = ~n29969 & ~n29971 ;
  assign n29973 = \m1_we_i_pad  & ~n14009 ;
  assign n29974 = n14017 & n29973 ;
  assign n29975 = \m2_we_i_pad  & n14009 ;
  assign n29976 = n14034 & n29975 ;
  assign n29977 = ~n29974 & ~n29976 ;
  assign n29978 = n29972 & n29977 ;
  assign n29979 = n29967 & n29978 ;
  assign n29980 = \m3_addr_i[0]_pad  & ~n14140 ;
  assign n29981 = n14133 & n29980 ;
  assign n29982 = \m4_addr_i[0]_pad  & n14140 ;
  assign n29983 = n14157 & n29982 ;
  assign n29984 = ~n29981 & ~n29983 ;
  assign n29985 = \m6_addr_i[0]_pad  & n14140 ;
  assign n29986 = n14148 & n29985 ;
  assign n29987 = \m2_addr_i[0]_pad  & n14140 ;
  assign n29988 = n14133 & n29987 ;
  assign n29989 = ~n29986 & ~n29988 ;
  assign n29990 = n29984 & n29989 ;
  assign n29991 = \m5_addr_i[0]_pad  & ~n14140 ;
  assign n29992 = n14157 & n29991 ;
  assign n29993 = \m1_addr_i[0]_pad  & ~n14140 ;
  assign n29994 = n14165 & n29993 ;
  assign n29995 = ~n29992 & ~n29994 ;
  assign n29996 = \m0_addr_i[0]_pad  & n14140 ;
  assign n29997 = n14165 & n29996 ;
  assign n29998 = \m7_addr_i[0]_pad  & ~n14140 ;
  assign n29999 = n14148 & n29998 ;
  assign n30000 = ~n29997 & ~n29999 ;
  assign n30001 = n29995 & n30000 ;
  assign n30002 = n29990 & n30001 ;
  assign n30003 = \m3_addr_i[10]_pad  & ~n14140 ;
  assign n30004 = n14133 & n30003 ;
  assign n30005 = \m4_addr_i[10]_pad  & n14140 ;
  assign n30006 = n14157 & n30005 ;
  assign n30007 = ~n30004 & ~n30006 ;
  assign n30008 = \m1_addr_i[10]_pad  & ~n14140 ;
  assign n30009 = n14165 & n30008 ;
  assign n30010 = \m5_addr_i[10]_pad  & ~n14140 ;
  assign n30011 = n14157 & n30010 ;
  assign n30012 = ~n30009 & ~n30011 ;
  assign n30013 = n30007 & n30012 ;
  assign n30014 = \m2_addr_i[10]_pad  & n14140 ;
  assign n30015 = n14133 & n30014 ;
  assign n30016 = \m6_addr_i[10]_pad  & n14140 ;
  assign n30017 = n14148 & n30016 ;
  assign n30018 = ~n30015 & ~n30017 ;
  assign n30019 = \m0_addr_i[10]_pad  & n14140 ;
  assign n30020 = n14165 & n30019 ;
  assign n30021 = \m7_addr_i[10]_pad  & ~n14140 ;
  assign n30022 = n14148 & n30021 ;
  assign n30023 = ~n30020 & ~n30022 ;
  assign n30024 = n30018 & n30023 ;
  assign n30025 = n30013 & n30024 ;
  assign n30026 = \m1_addr_i[11]_pad  & ~n14140 ;
  assign n30027 = n14165 & n30026 ;
  assign n30028 = \m2_addr_i[11]_pad  & n14140 ;
  assign n30029 = n14133 & n30028 ;
  assign n30030 = ~n30027 & ~n30029 ;
  assign n30031 = \m6_addr_i[11]_pad  & n14140 ;
  assign n30032 = n14148 & n30031 ;
  assign n30033 = \m7_addr_i[11]_pad  & ~n14140 ;
  assign n30034 = n14148 & n30033 ;
  assign n30035 = ~n30032 & ~n30034 ;
  assign n30036 = n30030 & n30035 ;
  assign n30037 = \m5_addr_i[11]_pad  & ~n14140 ;
  assign n30038 = n14157 & n30037 ;
  assign n30039 = \m0_addr_i[11]_pad  & n14140 ;
  assign n30040 = n14165 & n30039 ;
  assign n30041 = ~n30038 & ~n30040 ;
  assign n30042 = \m3_addr_i[11]_pad  & ~n14140 ;
  assign n30043 = n14133 & n30042 ;
  assign n30044 = \m4_addr_i[11]_pad  & n14140 ;
  assign n30045 = n14157 & n30044 ;
  assign n30046 = ~n30043 & ~n30045 ;
  assign n30047 = n30041 & n30046 ;
  assign n30048 = n30036 & n30047 ;
  assign n30049 = \m0_addr_i[12]_pad  & n14140 ;
  assign n30050 = n14165 & n30049 ;
  assign n30051 = \m7_addr_i[12]_pad  & ~n14140 ;
  assign n30052 = n14148 & n30051 ;
  assign n30053 = ~n30050 & ~n30052 ;
  assign n30054 = \m6_addr_i[12]_pad  & n14140 ;
  assign n30055 = n14148 & n30054 ;
  assign n30056 = \m2_addr_i[12]_pad  & n14140 ;
  assign n30057 = n14133 & n30056 ;
  assign n30058 = ~n30055 & ~n30057 ;
  assign n30059 = n30053 & n30058 ;
  assign n30060 = \m5_addr_i[12]_pad  & ~n14140 ;
  assign n30061 = n14157 & n30060 ;
  assign n30062 = \m1_addr_i[12]_pad  & ~n14140 ;
  assign n30063 = n14165 & n30062 ;
  assign n30064 = ~n30061 & ~n30063 ;
  assign n30065 = \m3_addr_i[12]_pad  & ~n14140 ;
  assign n30066 = n14133 & n30065 ;
  assign n30067 = \m4_addr_i[12]_pad  & n14140 ;
  assign n30068 = n14157 & n30067 ;
  assign n30069 = ~n30066 & ~n30068 ;
  assign n30070 = n30064 & n30069 ;
  assign n30071 = n30059 & n30070 ;
  assign n30072 = \m3_addr_i[13]_pad  & ~n14140 ;
  assign n30073 = n14133 & n30072 ;
  assign n30074 = \m4_addr_i[13]_pad  & n14140 ;
  assign n30075 = n14157 & n30074 ;
  assign n30076 = ~n30073 & ~n30075 ;
  assign n30077 = \m6_addr_i[13]_pad  & n14140 ;
  assign n30078 = n14148 & n30077 ;
  assign n30079 = \m2_addr_i[13]_pad  & n14140 ;
  assign n30080 = n14133 & n30079 ;
  assign n30081 = ~n30078 & ~n30080 ;
  assign n30082 = n30076 & n30081 ;
  assign n30083 = \m5_addr_i[13]_pad  & ~n14140 ;
  assign n30084 = n14157 & n30083 ;
  assign n30085 = \m1_addr_i[13]_pad  & ~n14140 ;
  assign n30086 = n14165 & n30085 ;
  assign n30087 = ~n30084 & ~n30086 ;
  assign n30088 = \m0_addr_i[13]_pad  & n14140 ;
  assign n30089 = n14165 & n30088 ;
  assign n30090 = \m7_addr_i[13]_pad  & ~n14140 ;
  assign n30091 = n14148 & n30090 ;
  assign n30092 = ~n30089 & ~n30091 ;
  assign n30093 = n30087 & n30092 ;
  assign n30094 = n30082 & n30093 ;
  assign n30095 = \m3_addr_i[14]_pad  & ~n14140 ;
  assign n30096 = n14133 & n30095 ;
  assign n30097 = \m4_addr_i[14]_pad  & n14140 ;
  assign n30098 = n14157 & n30097 ;
  assign n30099 = ~n30096 & ~n30098 ;
  assign n30100 = \m6_addr_i[14]_pad  & n14140 ;
  assign n30101 = n14148 & n30100 ;
  assign n30102 = \m2_addr_i[14]_pad  & n14140 ;
  assign n30103 = n14133 & n30102 ;
  assign n30104 = ~n30101 & ~n30103 ;
  assign n30105 = n30099 & n30104 ;
  assign n30106 = \m5_addr_i[14]_pad  & ~n14140 ;
  assign n30107 = n14157 & n30106 ;
  assign n30108 = \m1_addr_i[14]_pad  & ~n14140 ;
  assign n30109 = n14165 & n30108 ;
  assign n30110 = ~n30107 & ~n30109 ;
  assign n30111 = \m0_addr_i[14]_pad  & n14140 ;
  assign n30112 = n14165 & n30111 ;
  assign n30113 = \m7_addr_i[14]_pad  & ~n14140 ;
  assign n30114 = n14148 & n30113 ;
  assign n30115 = ~n30112 & ~n30114 ;
  assign n30116 = n30110 & n30115 ;
  assign n30117 = n30105 & n30116 ;
  assign n30118 = \m3_addr_i[15]_pad  & ~n14140 ;
  assign n30119 = n14133 & n30118 ;
  assign n30120 = \m4_addr_i[15]_pad  & n14140 ;
  assign n30121 = n14157 & n30120 ;
  assign n30122 = ~n30119 & ~n30121 ;
  assign n30123 = \m6_addr_i[15]_pad  & n14140 ;
  assign n30124 = n14148 & n30123 ;
  assign n30125 = \m2_addr_i[15]_pad  & n14140 ;
  assign n30126 = n14133 & n30125 ;
  assign n30127 = ~n30124 & ~n30126 ;
  assign n30128 = n30122 & n30127 ;
  assign n30129 = \m5_addr_i[15]_pad  & ~n14140 ;
  assign n30130 = n14157 & n30129 ;
  assign n30131 = \m1_addr_i[15]_pad  & ~n14140 ;
  assign n30132 = n14165 & n30131 ;
  assign n30133 = ~n30130 & ~n30132 ;
  assign n30134 = \m0_addr_i[15]_pad  & n14140 ;
  assign n30135 = n14165 & n30134 ;
  assign n30136 = \m7_addr_i[15]_pad  & ~n14140 ;
  assign n30137 = n14148 & n30136 ;
  assign n30138 = ~n30135 & ~n30137 ;
  assign n30139 = n30133 & n30138 ;
  assign n30140 = n30128 & n30139 ;
  assign n30141 = \m3_addr_i[16]_pad  & ~n14140 ;
  assign n30142 = n14133 & n30141 ;
  assign n30143 = \m4_addr_i[16]_pad  & n14140 ;
  assign n30144 = n14157 & n30143 ;
  assign n30145 = ~n30142 & ~n30144 ;
  assign n30146 = \m6_addr_i[16]_pad  & n14140 ;
  assign n30147 = n14148 & n30146 ;
  assign n30148 = \m2_addr_i[16]_pad  & n14140 ;
  assign n30149 = n14133 & n30148 ;
  assign n30150 = ~n30147 & ~n30149 ;
  assign n30151 = n30145 & n30150 ;
  assign n30152 = \m5_addr_i[16]_pad  & ~n14140 ;
  assign n30153 = n14157 & n30152 ;
  assign n30154 = \m1_addr_i[16]_pad  & ~n14140 ;
  assign n30155 = n14165 & n30154 ;
  assign n30156 = ~n30153 & ~n30155 ;
  assign n30157 = \m0_addr_i[16]_pad  & n14140 ;
  assign n30158 = n14165 & n30157 ;
  assign n30159 = \m7_addr_i[16]_pad  & ~n14140 ;
  assign n30160 = n14148 & n30159 ;
  assign n30161 = ~n30158 & ~n30160 ;
  assign n30162 = n30156 & n30161 ;
  assign n30163 = n30151 & n30162 ;
  assign n30164 = \m3_addr_i[17]_pad  & ~n14140 ;
  assign n30165 = n14133 & n30164 ;
  assign n30166 = \m4_addr_i[17]_pad  & n14140 ;
  assign n30167 = n14157 & n30166 ;
  assign n30168 = ~n30165 & ~n30167 ;
  assign n30169 = \m6_addr_i[17]_pad  & n14140 ;
  assign n30170 = n14148 & n30169 ;
  assign n30171 = \m2_addr_i[17]_pad  & n14140 ;
  assign n30172 = n14133 & n30171 ;
  assign n30173 = ~n30170 & ~n30172 ;
  assign n30174 = n30168 & n30173 ;
  assign n30175 = \m5_addr_i[17]_pad  & ~n14140 ;
  assign n30176 = n14157 & n30175 ;
  assign n30177 = \m1_addr_i[17]_pad  & ~n14140 ;
  assign n30178 = n14165 & n30177 ;
  assign n30179 = ~n30176 & ~n30178 ;
  assign n30180 = \m0_addr_i[17]_pad  & n14140 ;
  assign n30181 = n14165 & n30180 ;
  assign n30182 = \m7_addr_i[17]_pad  & ~n14140 ;
  assign n30183 = n14148 & n30182 ;
  assign n30184 = ~n30181 & ~n30183 ;
  assign n30185 = n30179 & n30184 ;
  assign n30186 = n30174 & n30185 ;
  assign n30187 = \m1_addr_i[18]_pad  & ~n14140 ;
  assign n30188 = n14165 & n30187 ;
  assign n30189 = \m2_addr_i[18]_pad  & n14140 ;
  assign n30190 = n14133 & n30189 ;
  assign n30191 = ~n30188 & ~n30190 ;
  assign n30192 = \m6_addr_i[18]_pad  & n14140 ;
  assign n30193 = n14148 & n30192 ;
  assign n30194 = \m7_addr_i[18]_pad  & ~n14140 ;
  assign n30195 = n14148 & n30194 ;
  assign n30196 = ~n30193 & ~n30195 ;
  assign n30197 = n30191 & n30196 ;
  assign n30198 = \m5_addr_i[18]_pad  & ~n14140 ;
  assign n30199 = n14157 & n30198 ;
  assign n30200 = \m0_addr_i[18]_pad  & n14140 ;
  assign n30201 = n14165 & n30200 ;
  assign n30202 = ~n30199 & ~n30201 ;
  assign n30203 = \m3_addr_i[18]_pad  & ~n14140 ;
  assign n30204 = n14133 & n30203 ;
  assign n30205 = \m4_addr_i[18]_pad  & n14140 ;
  assign n30206 = n14157 & n30205 ;
  assign n30207 = ~n30204 & ~n30206 ;
  assign n30208 = n30202 & n30207 ;
  assign n30209 = n30197 & n30208 ;
  assign n30210 = \m0_addr_i[19]_pad  & n14140 ;
  assign n30211 = n14165 & n30210 ;
  assign n30212 = \m7_addr_i[19]_pad  & ~n14140 ;
  assign n30213 = n14148 & n30212 ;
  assign n30214 = ~n30211 & ~n30213 ;
  assign n30215 = \m6_addr_i[19]_pad  & n14140 ;
  assign n30216 = n14148 & n30215 ;
  assign n30217 = \m4_addr_i[19]_pad  & n14140 ;
  assign n30218 = n14157 & n30217 ;
  assign n30219 = ~n30216 & ~n30218 ;
  assign n30220 = n30214 & n30219 ;
  assign n30221 = \m5_addr_i[19]_pad  & ~n14140 ;
  assign n30222 = n14157 & n30221 ;
  assign n30223 = \m3_addr_i[19]_pad  & ~n14140 ;
  assign n30224 = n14133 & n30223 ;
  assign n30225 = ~n30222 & ~n30224 ;
  assign n30226 = \m1_addr_i[19]_pad  & ~n14140 ;
  assign n30227 = n14165 & n30226 ;
  assign n30228 = \m2_addr_i[19]_pad  & n14140 ;
  assign n30229 = n14133 & n30228 ;
  assign n30230 = ~n30227 & ~n30229 ;
  assign n30231 = n30225 & n30230 ;
  assign n30232 = n30220 & n30231 ;
  assign n30233 = \m3_addr_i[1]_pad  & ~n14140 ;
  assign n30234 = n14133 & n30233 ;
  assign n30235 = \m4_addr_i[1]_pad  & n14140 ;
  assign n30236 = n14157 & n30235 ;
  assign n30237 = ~n30234 & ~n30236 ;
  assign n30238 = \m6_addr_i[1]_pad  & n14140 ;
  assign n30239 = n14148 & n30238 ;
  assign n30240 = \m2_addr_i[1]_pad  & n14140 ;
  assign n30241 = n14133 & n30240 ;
  assign n30242 = ~n30239 & ~n30241 ;
  assign n30243 = n30237 & n30242 ;
  assign n30244 = \m5_addr_i[1]_pad  & ~n14140 ;
  assign n30245 = n14157 & n30244 ;
  assign n30246 = \m1_addr_i[1]_pad  & ~n14140 ;
  assign n30247 = n14165 & n30246 ;
  assign n30248 = ~n30245 & ~n30247 ;
  assign n30249 = \m0_addr_i[1]_pad  & n14140 ;
  assign n30250 = n14165 & n30249 ;
  assign n30251 = \m7_addr_i[1]_pad  & ~n14140 ;
  assign n30252 = n14148 & n30251 ;
  assign n30253 = ~n30250 & ~n30252 ;
  assign n30254 = n30248 & n30253 ;
  assign n30255 = n30243 & n30254 ;
  assign n30256 = \m6_addr_i[20]_pad  & n14140 ;
  assign n30257 = n14148 & n30256 ;
  assign n30258 = \m5_addr_i[20]_pad  & ~n14140 ;
  assign n30259 = n14157 & n30258 ;
  assign n30260 = ~n30257 & ~n30259 ;
  assign n30261 = \m1_addr_i[20]_pad  & ~n14140 ;
  assign n30262 = n14165 & n30261 ;
  assign n30263 = \m4_addr_i[20]_pad  & n14140 ;
  assign n30264 = n14157 & n30263 ;
  assign n30265 = ~n30262 & ~n30264 ;
  assign n30266 = n30260 & n30265 ;
  assign n30267 = \m2_addr_i[20]_pad  & n14140 ;
  assign n30268 = n14133 & n30267 ;
  assign n30269 = \m3_addr_i[20]_pad  & ~n14140 ;
  assign n30270 = n14133 & n30269 ;
  assign n30271 = ~n30268 & ~n30270 ;
  assign n30272 = \m0_addr_i[20]_pad  & n14140 ;
  assign n30273 = n14165 & n30272 ;
  assign n30274 = \m7_addr_i[20]_pad  & ~n14140 ;
  assign n30275 = n14148 & n30274 ;
  assign n30276 = ~n30273 & ~n30275 ;
  assign n30277 = n30271 & n30276 ;
  assign n30278 = n30266 & n30277 ;
  assign n30279 = \m0_addr_i[21]_pad  & n14140 ;
  assign n30280 = n14165 & n30279 ;
  assign n30281 = \m7_addr_i[21]_pad  & ~n14140 ;
  assign n30282 = n14148 & n30281 ;
  assign n30283 = ~n30280 & ~n30282 ;
  assign n30284 = \m1_addr_i[21]_pad  & ~n14140 ;
  assign n30285 = n14165 & n30284 ;
  assign n30286 = \m4_addr_i[21]_pad  & n14140 ;
  assign n30287 = n14157 & n30286 ;
  assign n30288 = ~n30285 & ~n30287 ;
  assign n30289 = n30283 & n30288 ;
  assign n30290 = \m2_addr_i[21]_pad  & n14140 ;
  assign n30291 = n14133 & n30290 ;
  assign n30292 = \m3_addr_i[21]_pad  & ~n14140 ;
  assign n30293 = n14133 & n30292 ;
  assign n30294 = ~n30291 & ~n30293 ;
  assign n30295 = \m6_addr_i[21]_pad  & n14140 ;
  assign n30296 = n14148 & n30295 ;
  assign n30297 = \m5_addr_i[21]_pad  & ~n14140 ;
  assign n30298 = n14157 & n30297 ;
  assign n30299 = ~n30296 & ~n30298 ;
  assign n30300 = n30294 & n30299 ;
  assign n30301 = n30289 & n30300 ;
  assign n30302 = \m0_addr_i[22]_pad  & n14140 ;
  assign n30303 = n14165 & n30302 ;
  assign n30304 = \m7_addr_i[22]_pad  & ~n14140 ;
  assign n30305 = n14148 & n30304 ;
  assign n30306 = ~n30303 & ~n30305 ;
  assign n30307 = \m3_addr_i[22]_pad  & ~n14140 ;
  assign n30308 = n14133 & n30307 ;
  assign n30309 = \m2_addr_i[22]_pad  & n14140 ;
  assign n30310 = n14133 & n30309 ;
  assign n30311 = ~n30308 & ~n30310 ;
  assign n30312 = n30306 & n30311 ;
  assign n30313 = \m4_addr_i[22]_pad  & n14140 ;
  assign n30314 = n14157 & n30313 ;
  assign n30315 = \m1_addr_i[22]_pad  & ~n14140 ;
  assign n30316 = n14165 & n30315 ;
  assign n30317 = ~n30314 & ~n30316 ;
  assign n30318 = \m6_addr_i[22]_pad  & n14140 ;
  assign n30319 = n14148 & n30318 ;
  assign n30320 = \m5_addr_i[22]_pad  & ~n14140 ;
  assign n30321 = n14157 & n30320 ;
  assign n30322 = ~n30319 & ~n30321 ;
  assign n30323 = n30317 & n30322 ;
  assign n30324 = n30312 & n30323 ;
  assign n30325 = \m6_addr_i[23]_pad  & n14140 ;
  assign n30326 = n14148 & n30325 ;
  assign n30327 = \m5_addr_i[23]_pad  & ~n14140 ;
  assign n30328 = n14157 & n30327 ;
  assign n30329 = ~n30326 & ~n30328 ;
  assign n30330 = \m3_addr_i[23]_pad  & ~n14140 ;
  assign n30331 = n14133 & n30330 ;
  assign n30332 = \m7_addr_i[23]_pad  & ~n14140 ;
  assign n30333 = n14148 & n30332 ;
  assign n30334 = ~n30331 & ~n30333 ;
  assign n30335 = n30329 & n30334 ;
  assign n30336 = \m4_addr_i[23]_pad  & n14140 ;
  assign n30337 = n14157 & n30336 ;
  assign n30338 = \m0_addr_i[23]_pad  & n14140 ;
  assign n30339 = n14165 & n30338 ;
  assign n30340 = ~n30337 & ~n30339 ;
  assign n30341 = \m1_addr_i[23]_pad  & ~n14140 ;
  assign n30342 = n14165 & n30341 ;
  assign n30343 = \m2_addr_i[23]_pad  & n14140 ;
  assign n30344 = n14133 & n30343 ;
  assign n30345 = ~n30342 & ~n30344 ;
  assign n30346 = n30340 & n30345 ;
  assign n30347 = n30335 & n30346 ;
  assign n30348 = \m3_addr_i[24]_pad  & ~n14140 ;
  assign n30349 = n14133 & n30348 ;
  assign n30350 = \m4_addr_i[24]_pad  & n14140 ;
  assign n30351 = n14157 & n30350 ;
  assign n30352 = ~n30349 & ~n30351 ;
  assign n30353 = \m1_addr_i[24]_pad  & ~n14140 ;
  assign n30354 = n14165 & n30353 ;
  assign n30355 = \m6_addr_i[24]_pad  & n14140 ;
  assign n30356 = n14148 & n30355 ;
  assign n30357 = ~n30354 & ~n30356 ;
  assign n30358 = n30352 & n30357 ;
  assign n30359 = \m2_addr_i[24]_pad  & n14140 ;
  assign n30360 = n14133 & n30359 ;
  assign n30361 = \m5_addr_i[24]_pad  & ~n14140 ;
  assign n30362 = n14157 & n30361 ;
  assign n30363 = ~n30360 & ~n30362 ;
  assign n30364 = \m0_addr_i[24]_pad  & n14140 ;
  assign n30365 = n14165 & n30364 ;
  assign n30366 = \m7_addr_i[24]_pad  & ~n14140 ;
  assign n30367 = n14148 & n30366 ;
  assign n30368 = ~n30365 & ~n30367 ;
  assign n30369 = n30363 & n30368 ;
  assign n30370 = n30358 & n30369 ;
  assign n30371 = \m0_addr_i[25]_pad  & n14140 ;
  assign n30372 = n14165 & n30371 ;
  assign n30373 = \m7_addr_i[25]_pad  & ~n14140 ;
  assign n30374 = n14148 & n30373 ;
  assign n30375 = ~n30372 & ~n30374 ;
  assign n30376 = \m3_addr_i[25]_pad  & ~n14140 ;
  assign n30377 = n14133 & n30376 ;
  assign n30378 = \m6_addr_i[25]_pad  & n14140 ;
  assign n30379 = n14148 & n30378 ;
  assign n30380 = ~n30377 & ~n30379 ;
  assign n30381 = n30375 & n30380 ;
  assign n30382 = \m4_addr_i[25]_pad  & n14140 ;
  assign n30383 = n14157 & n30382 ;
  assign n30384 = \m5_addr_i[25]_pad  & ~n14140 ;
  assign n30385 = n14157 & n30384 ;
  assign n30386 = ~n30383 & ~n30385 ;
  assign n30387 = \m1_addr_i[25]_pad  & ~n14140 ;
  assign n30388 = n14165 & n30387 ;
  assign n30389 = \m2_addr_i[25]_pad  & n14140 ;
  assign n30390 = n14133 & n30389 ;
  assign n30391 = ~n30388 & ~n30390 ;
  assign n30392 = n30386 & n30391 ;
  assign n30393 = n30381 & n30392 ;
  assign n30394 = \m1_addr_i[26]_pad  & ~n14140 ;
  assign n30395 = n14165 & n30394 ;
  assign n30396 = \m2_addr_i[26]_pad  & n14140 ;
  assign n30397 = n14133 & n30396 ;
  assign n30398 = ~n30395 & ~n30397 ;
  assign n30399 = \m3_addr_i[26]_pad  & ~n14140 ;
  assign n30400 = n14133 & n30399 ;
  assign n30401 = \m6_addr_i[26]_pad  & n14140 ;
  assign n30402 = n14148 & n30401 ;
  assign n30403 = ~n30400 & ~n30402 ;
  assign n30404 = n30398 & n30403 ;
  assign n30405 = \m4_addr_i[26]_pad  & n14140 ;
  assign n30406 = n14157 & n30405 ;
  assign n30407 = \m5_addr_i[26]_pad  & ~n14140 ;
  assign n30408 = n14157 & n30407 ;
  assign n30409 = ~n30406 & ~n30408 ;
  assign n30410 = \m0_addr_i[26]_pad  & n14140 ;
  assign n30411 = n14165 & n30410 ;
  assign n30412 = \m7_addr_i[26]_pad  & ~n14140 ;
  assign n30413 = n14148 & n30412 ;
  assign n30414 = ~n30411 & ~n30413 ;
  assign n30415 = n30409 & n30414 ;
  assign n30416 = n30404 & n30415 ;
  assign n30417 = \m3_addr_i[27]_pad  & ~n14140 ;
  assign n30418 = n14133 & n30417 ;
  assign n30419 = \m4_addr_i[27]_pad  & n14140 ;
  assign n30420 = n14157 & n30419 ;
  assign n30421 = ~n30418 & ~n30420 ;
  assign n30422 = \m5_addr_i[27]_pad  & ~n14140 ;
  assign n30423 = n14157 & n30422 ;
  assign n30424 = \m7_addr_i[27]_pad  & ~n14140 ;
  assign n30425 = n14148 & n30424 ;
  assign n30426 = ~n30423 & ~n30425 ;
  assign n30427 = n30421 & n30426 ;
  assign n30428 = \m6_addr_i[27]_pad  & n14140 ;
  assign n30429 = n14148 & n30428 ;
  assign n30430 = \m0_addr_i[27]_pad  & n14140 ;
  assign n30431 = n14165 & n30430 ;
  assign n30432 = ~n30429 & ~n30431 ;
  assign n30433 = \m1_addr_i[27]_pad  & ~n14140 ;
  assign n30434 = n14165 & n30433 ;
  assign n30435 = \m2_addr_i[27]_pad  & n14140 ;
  assign n30436 = n14133 & n30435 ;
  assign n30437 = ~n30434 & ~n30436 ;
  assign n30438 = n30432 & n30437 ;
  assign n30439 = n30427 & n30438 ;
  assign n30440 = \m1_addr_i[28]_pad  & ~n14140 ;
  assign n30441 = n14165 & n30440 ;
  assign n30442 = \m2_addr_i[28]_pad  & n14140 ;
  assign n30443 = n14133 & n30442 ;
  assign n30444 = ~n30441 & ~n30443 ;
  assign n30445 = \m3_addr_i[28]_pad  & ~n14140 ;
  assign n30446 = n14133 & n30445 ;
  assign n30447 = \m7_addr_i[28]_pad  & ~n14140 ;
  assign n30448 = n14148 & n30447 ;
  assign n30449 = ~n30446 & ~n30448 ;
  assign n30450 = n30444 & n30449 ;
  assign n30451 = \m4_addr_i[28]_pad  & n14140 ;
  assign n30452 = n14157 & n30451 ;
  assign n30453 = \m0_addr_i[28]_pad  & n14140 ;
  assign n30454 = n14165 & n30453 ;
  assign n30455 = ~n30452 & ~n30454 ;
  assign n30456 = \m5_addr_i[28]_pad  & ~n14140 ;
  assign n30457 = n14157 & n30456 ;
  assign n30458 = \m6_addr_i[28]_pad  & n14140 ;
  assign n30459 = n14148 & n30458 ;
  assign n30460 = ~n30457 & ~n30459 ;
  assign n30461 = n30455 & n30460 ;
  assign n30462 = n30450 & n30461 ;
  assign n30463 = \m3_addr_i[29]_pad  & ~n14140 ;
  assign n30464 = n14133 & n30463 ;
  assign n30465 = \m4_addr_i[29]_pad  & n14140 ;
  assign n30466 = n14157 & n30465 ;
  assign n30467 = ~n30464 & ~n30466 ;
  assign n30468 = \m5_addr_i[29]_pad  & ~n14140 ;
  assign n30469 = n14157 & n30468 ;
  assign n30470 = \m2_addr_i[29]_pad  & n14140 ;
  assign n30471 = n14133 & n30470 ;
  assign n30472 = ~n30469 & ~n30471 ;
  assign n30473 = n30467 & n30472 ;
  assign n30474 = \m6_addr_i[29]_pad  & n14140 ;
  assign n30475 = n14148 & n30474 ;
  assign n30476 = \m1_addr_i[29]_pad  & ~n14140 ;
  assign n30477 = n14165 & n30476 ;
  assign n30478 = ~n30475 & ~n30477 ;
  assign n30479 = \m0_addr_i[29]_pad  & n14140 ;
  assign n30480 = n14165 & n30479 ;
  assign n30481 = \m7_addr_i[29]_pad  & ~n14140 ;
  assign n30482 = n14148 & n30481 ;
  assign n30483 = ~n30480 & ~n30482 ;
  assign n30484 = n30478 & n30483 ;
  assign n30485 = n30473 & n30484 ;
  assign n30486 = \m3_addr_i[2]_pad  & ~n14140 ;
  assign n30487 = n14133 & n30486 ;
  assign n30488 = \m4_addr_i[2]_pad  & n14140 ;
  assign n30489 = n14157 & n30488 ;
  assign n30490 = ~n30487 & ~n30489 ;
  assign n30491 = \m6_addr_i[2]_pad  & n14140 ;
  assign n30492 = n14148 & n30491 ;
  assign n30493 = \m2_addr_i[2]_pad  & n14140 ;
  assign n30494 = n14133 & n30493 ;
  assign n30495 = ~n30492 & ~n30494 ;
  assign n30496 = n30490 & n30495 ;
  assign n30497 = \m5_addr_i[2]_pad  & ~n14140 ;
  assign n30498 = n14157 & n30497 ;
  assign n30499 = \m1_addr_i[2]_pad  & ~n14140 ;
  assign n30500 = n14165 & n30499 ;
  assign n30501 = ~n30498 & ~n30500 ;
  assign n30502 = \m0_addr_i[2]_pad  & n14140 ;
  assign n30503 = n14165 & n30502 ;
  assign n30504 = \m7_addr_i[2]_pad  & ~n14140 ;
  assign n30505 = n14148 & n30504 ;
  assign n30506 = ~n30503 & ~n30505 ;
  assign n30507 = n30501 & n30506 ;
  assign n30508 = n30496 & n30507 ;
  assign n30509 = \m1_addr_i[30]_pad  & ~n14140 ;
  assign n30510 = n14165 & n30509 ;
  assign n30511 = \m2_addr_i[30]_pad  & n14140 ;
  assign n30512 = n14133 & n30511 ;
  assign n30513 = ~n30510 & ~n30512 ;
  assign n30514 = \m5_addr_i[30]_pad  & ~n14140 ;
  assign n30515 = n14157 & n30514 ;
  assign n30516 = \m4_addr_i[30]_pad  & n14140 ;
  assign n30517 = n14157 & n30516 ;
  assign n30518 = ~n30515 & ~n30517 ;
  assign n30519 = n30513 & n30518 ;
  assign n30520 = \m6_addr_i[30]_pad  & n14140 ;
  assign n30521 = n14148 & n30520 ;
  assign n30522 = \m3_addr_i[30]_pad  & ~n14140 ;
  assign n30523 = n14133 & n30522 ;
  assign n30524 = ~n30521 & ~n30523 ;
  assign n30525 = \m0_addr_i[30]_pad  & n14140 ;
  assign n30526 = n14165 & n30525 ;
  assign n30527 = \m7_addr_i[30]_pad  & ~n14140 ;
  assign n30528 = n14148 & n30527 ;
  assign n30529 = ~n30526 & ~n30528 ;
  assign n30530 = n30524 & n30529 ;
  assign n30531 = n30519 & n30530 ;
  assign n30532 = \m0_addr_i[31]_pad  & n14140 ;
  assign n30533 = n14165 & n30532 ;
  assign n30534 = \m7_addr_i[31]_pad  & ~n14140 ;
  assign n30535 = n14148 & n30534 ;
  assign n30536 = ~n30533 & ~n30535 ;
  assign n30537 = \m1_addr_i[31]_pad  & ~n14140 ;
  assign n30538 = n14165 & n30537 ;
  assign n30539 = \m6_addr_i[31]_pad  & n14140 ;
  assign n30540 = n14148 & n30539 ;
  assign n30541 = ~n30538 & ~n30540 ;
  assign n30542 = n30536 & n30541 ;
  assign n30543 = \m2_addr_i[31]_pad  & n14140 ;
  assign n30544 = n14133 & n30543 ;
  assign n30545 = \m5_addr_i[31]_pad  & ~n14140 ;
  assign n30546 = n14157 & n30545 ;
  assign n30547 = ~n30544 & ~n30546 ;
  assign n30548 = \m3_addr_i[31]_pad  & ~n14140 ;
  assign n30549 = n14133 & n30548 ;
  assign n30550 = \m4_addr_i[31]_pad  & n14140 ;
  assign n30551 = n14157 & n30550 ;
  assign n30552 = ~n30549 & ~n30551 ;
  assign n30553 = n30547 & n30552 ;
  assign n30554 = n30542 & n30553 ;
  assign n30555 = \m3_addr_i[3]_pad  & ~n14140 ;
  assign n30556 = n14133 & n30555 ;
  assign n30557 = \m4_addr_i[3]_pad  & n14140 ;
  assign n30558 = n14157 & n30557 ;
  assign n30559 = ~n30556 & ~n30558 ;
  assign n30560 = \m6_addr_i[3]_pad  & n14140 ;
  assign n30561 = n14148 & n30560 ;
  assign n30562 = \m2_addr_i[3]_pad  & n14140 ;
  assign n30563 = n14133 & n30562 ;
  assign n30564 = ~n30561 & ~n30563 ;
  assign n30565 = n30559 & n30564 ;
  assign n30566 = \m5_addr_i[3]_pad  & ~n14140 ;
  assign n30567 = n14157 & n30566 ;
  assign n30568 = \m1_addr_i[3]_pad  & ~n14140 ;
  assign n30569 = n14165 & n30568 ;
  assign n30570 = ~n30567 & ~n30569 ;
  assign n30571 = \m0_addr_i[3]_pad  & n14140 ;
  assign n30572 = n14165 & n30571 ;
  assign n30573 = \m7_addr_i[3]_pad  & ~n14140 ;
  assign n30574 = n14148 & n30573 ;
  assign n30575 = ~n30572 & ~n30574 ;
  assign n30576 = n30570 & n30575 ;
  assign n30577 = n30565 & n30576 ;
  assign n30578 = \m3_addr_i[4]_pad  & ~n14140 ;
  assign n30579 = n14133 & n30578 ;
  assign n30580 = \m4_addr_i[4]_pad  & n14140 ;
  assign n30581 = n14157 & n30580 ;
  assign n30582 = ~n30579 & ~n30581 ;
  assign n30583 = \m6_addr_i[4]_pad  & n14140 ;
  assign n30584 = n14148 & n30583 ;
  assign n30585 = \m2_addr_i[4]_pad  & n14140 ;
  assign n30586 = n14133 & n30585 ;
  assign n30587 = ~n30584 & ~n30586 ;
  assign n30588 = n30582 & n30587 ;
  assign n30589 = \m5_addr_i[4]_pad  & ~n14140 ;
  assign n30590 = n14157 & n30589 ;
  assign n30591 = \m1_addr_i[4]_pad  & ~n14140 ;
  assign n30592 = n14165 & n30591 ;
  assign n30593 = ~n30590 & ~n30592 ;
  assign n30594 = \m0_addr_i[4]_pad  & n14140 ;
  assign n30595 = n14165 & n30594 ;
  assign n30596 = \m7_addr_i[4]_pad  & ~n14140 ;
  assign n30597 = n14148 & n30596 ;
  assign n30598 = ~n30595 & ~n30597 ;
  assign n30599 = n30593 & n30598 ;
  assign n30600 = n30588 & n30599 ;
  assign n30601 = \m3_addr_i[5]_pad  & ~n14140 ;
  assign n30602 = n14133 & n30601 ;
  assign n30603 = \m4_addr_i[5]_pad  & n14140 ;
  assign n30604 = n14157 & n30603 ;
  assign n30605 = ~n30602 & ~n30604 ;
  assign n30606 = \m6_addr_i[5]_pad  & n14140 ;
  assign n30607 = n14148 & n30606 ;
  assign n30608 = \m2_addr_i[5]_pad  & n14140 ;
  assign n30609 = n14133 & n30608 ;
  assign n30610 = ~n30607 & ~n30609 ;
  assign n30611 = n30605 & n30610 ;
  assign n30612 = \m5_addr_i[5]_pad  & ~n14140 ;
  assign n30613 = n14157 & n30612 ;
  assign n30614 = \m1_addr_i[5]_pad  & ~n14140 ;
  assign n30615 = n14165 & n30614 ;
  assign n30616 = ~n30613 & ~n30615 ;
  assign n30617 = \m0_addr_i[5]_pad  & n14140 ;
  assign n30618 = n14165 & n30617 ;
  assign n30619 = \m7_addr_i[5]_pad  & ~n14140 ;
  assign n30620 = n14148 & n30619 ;
  assign n30621 = ~n30618 & ~n30620 ;
  assign n30622 = n30616 & n30621 ;
  assign n30623 = n30611 & n30622 ;
  assign n30624 = \m3_addr_i[6]_pad  & ~n14140 ;
  assign n30625 = n14133 & n30624 ;
  assign n30626 = \m4_addr_i[6]_pad  & n14140 ;
  assign n30627 = n14157 & n30626 ;
  assign n30628 = ~n30625 & ~n30627 ;
  assign n30629 = \m6_addr_i[6]_pad  & n14140 ;
  assign n30630 = n14148 & n30629 ;
  assign n30631 = \m2_addr_i[6]_pad  & n14140 ;
  assign n30632 = n14133 & n30631 ;
  assign n30633 = ~n30630 & ~n30632 ;
  assign n30634 = n30628 & n30633 ;
  assign n30635 = \m5_addr_i[6]_pad  & ~n14140 ;
  assign n30636 = n14157 & n30635 ;
  assign n30637 = \m1_addr_i[6]_pad  & ~n14140 ;
  assign n30638 = n14165 & n30637 ;
  assign n30639 = ~n30636 & ~n30638 ;
  assign n30640 = \m0_addr_i[6]_pad  & n14140 ;
  assign n30641 = n14165 & n30640 ;
  assign n30642 = \m7_addr_i[6]_pad  & ~n14140 ;
  assign n30643 = n14148 & n30642 ;
  assign n30644 = ~n30641 & ~n30643 ;
  assign n30645 = n30639 & n30644 ;
  assign n30646 = n30634 & n30645 ;
  assign n30647 = \m1_addr_i[7]_pad  & ~n14140 ;
  assign n30648 = n14165 & n30647 ;
  assign n30649 = \m2_addr_i[7]_pad  & n14140 ;
  assign n30650 = n14133 & n30649 ;
  assign n30651 = ~n30648 & ~n30650 ;
  assign n30652 = \m6_addr_i[7]_pad  & n14140 ;
  assign n30653 = n14148 & n30652 ;
  assign n30654 = \m4_addr_i[7]_pad  & n14140 ;
  assign n30655 = n14157 & n30654 ;
  assign n30656 = ~n30653 & ~n30655 ;
  assign n30657 = n30651 & n30656 ;
  assign n30658 = \m5_addr_i[7]_pad  & ~n14140 ;
  assign n30659 = n14157 & n30658 ;
  assign n30660 = \m3_addr_i[7]_pad  & ~n14140 ;
  assign n30661 = n14133 & n30660 ;
  assign n30662 = ~n30659 & ~n30661 ;
  assign n30663 = \m0_addr_i[7]_pad  & n14140 ;
  assign n30664 = n14165 & n30663 ;
  assign n30665 = \m7_addr_i[7]_pad  & ~n14140 ;
  assign n30666 = n14148 & n30665 ;
  assign n30667 = ~n30664 & ~n30666 ;
  assign n30668 = n30662 & n30667 ;
  assign n30669 = n30657 & n30668 ;
  assign n30670 = \m0_addr_i[8]_pad  & n14140 ;
  assign n30671 = n14165 & n30670 ;
  assign n30672 = \m7_addr_i[8]_pad  & ~n14140 ;
  assign n30673 = n14148 & n30672 ;
  assign n30674 = ~n30671 & ~n30673 ;
  assign n30675 = \m6_addr_i[8]_pad  & n14140 ;
  assign n30676 = n14148 & n30675 ;
  assign n30677 = \m2_addr_i[8]_pad  & n14140 ;
  assign n30678 = n14133 & n30677 ;
  assign n30679 = ~n30676 & ~n30678 ;
  assign n30680 = n30674 & n30679 ;
  assign n30681 = \m5_addr_i[8]_pad  & ~n14140 ;
  assign n30682 = n14157 & n30681 ;
  assign n30683 = \m1_addr_i[8]_pad  & ~n14140 ;
  assign n30684 = n14165 & n30683 ;
  assign n30685 = ~n30682 & ~n30684 ;
  assign n30686 = \m3_addr_i[8]_pad  & ~n14140 ;
  assign n30687 = n14133 & n30686 ;
  assign n30688 = \m4_addr_i[8]_pad  & n14140 ;
  assign n30689 = n14157 & n30688 ;
  assign n30690 = ~n30687 & ~n30689 ;
  assign n30691 = n30685 & n30690 ;
  assign n30692 = n30680 & n30691 ;
  assign n30693 = \m6_addr_i[9]_pad  & n14140 ;
  assign n30694 = n14148 & n30693 ;
  assign n30695 = \m5_addr_i[9]_pad  & ~n14140 ;
  assign n30696 = n14157 & n30695 ;
  assign n30697 = ~n30694 & ~n30696 ;
  assign n30698 = \m0_addr_i[9]_pad  & n14140 ;
  assign n30699 = n14165 & n30698 ;
  assign n30700 = \m4_addr_i[9]_pad  & n14140 ;
  assign n30701 = n14157 & n30700 ;
  assign n30702 = ~n30699 & ~n30701 ;
  assign n30703 = n30697 & n30702 ;
  assign n30704 = \m7_addr_i[9]_pad  & ~n14140 ;
  assign n30705 = n14148 & n30704 ;
  assign n30706 = \m3_addr_i[9]_pad  & ~n14140 ;
  assign n30707 = n14133 & n30706 ;
  assign n30708 = ~n30705 & ~n30707 ;
  assign n30709 = \m1_addr_i[9]_pad  & ~n14140 ;
  assign n30710 = n14165 & n30709 ;
  assign n30711 = \m2_addr_i[9]_pad  & n14140 ;
  assign n30712 = n14133 & n30711 ;
  assign n30713 = ~n30710 & ~n30712 ;
  assign n30714 = n30708 & n30713 ;
  assign n30715 = n30703 & n30714 ;
  assign n30716 = \m1_data_i[0]_pad  & ~n14140 ;
  assign n30717 = n14165 & n30716 ;
  assign n30718 = \m2_data_i[0]_pad  & n14140 ;
  assign n30719 = n14133 & n30718 ;
  assign n30720 = ~n30717 & ~n30719 ;
  assign n30721 = \m0_data_i[0]_pad  & n14140 ;
  assign n30722 = n14165 & n30721 ;
  assign n30723 = \m5_data_i[0]_pad  & ~n14140 ;
  assign n30724 = n14157 & n30723 ;
  assign n30725 = ~n30722 & ~n30724 ;
  assign n30726 = n30720 & n30725 ;
  assign n30727 = \m7_data_i[0]_pad  & ~n14140 ;
  assign n30728 = n14148 & n30727 ;
  assign n30729 = \m6_data_i[0]_pad  & n14140 ;
  assign n30730 = n14148 & n30729 ;
  assign n30731 = ~n30728 & ~n30730 ;
  assign n30732 = \m3_data_i[0]_pad  & ~n14140 ;
  assign n30733 = n14133 & n30732 ;
  assign n30734 = \m4_data_i[0]_pad  & n14140 ;
  assign n30735 = n14157 & n30734 ;
  assign n30736 = ~n30733 & ~n30735 ;
  assign n30737 = n30731 & n30736 ;
  assign n30738 = n30726 & n30737 ;
  assign n30739 = \m0_data_i[10]_pad  & n14140 ;
  assign n30740 = n14165 & n30739 ;
  assign n30741 = \m7_data_i[10]_pad  & ~n14140 ;
  assign n30742 = n14148 & n30741 ;
  assign n30743 = ~n30740 & ~n30742 ;
  assign n30744 = \m1_data_i[10]_pad  & ~n14140 ;
  assign n30745 = n14165 & n30744 ;
  assign n30746 = \m4_data_i[10]_pad  & n14140 ;
  assign n30747 = n14157 & n30746 ;
  assign n30748 = ~n30745 & ~n30747 ;
  assign n30749 = n30743 & n30748 ;
  assign n30750 = \m2_data_i[10]_pad  & n14140 ;
  assign n30751 = n14133 & n30750 ;
  assign n30752 = \m3_data_i[10]_pad  & ~n14140 ;
  assign n30753 = n14133 & n30752 ;
  assign n30754 = ~n30751 & ~n30753 ;
  assign n30755 = \m6_data_i[10]_pad  & n14140 ;
  assign n30756 = n14148 & n30755 ;
  assign n30757 = \m5_data_i[10]_pad  & ~n14140 ;
  assign n30758 = n14157 & n30757 ;
  assign n30759 = ~n30756 & ~n30758 ;
  assign n30760 = n30754 & n30759 ;
  assign n30761 = n30749 & n30760 ;
  assign n30762 = \m1_data_i[11]_pad  & ~n14140 ;
  assign n30763 = n14165 & n30762 ;
  assign n30764 = \m2_data_i[11]_pad  & n14140 ;
  assign n30765 = n14133 & n30764 ;
  assign n30766 = ~n30763 & ~n30765 ;
  assign n30767 = \m0_data_i[11]_pad  & n14140 ;
  assign n30768 = n14165 & n30767 ;
  assign n30769 = \m5_data_i[11]_pad  & ~n14140 ;
  assign n30770 = n14157 & n30769 ;
  assign n30771 = ~n30768 & ~n30770 ;
  assign n30772 = n30766 & n30771 ;
  assign n30773 = \m7_data_i[11]_pad  & ~n14140 ;
  assign n30774 = n14148 & n30773 ;
  assign n30775 = \m6_data_i[11]_pad  & n14140 ;
  assign n30776 = n14148 & n30775 ;
  assign n30777 = ~n30774 & ~n30776 ;
  assign n30778 = \m3_data_i[11]_pad  & ~n14140 ;
  assign n30779 = n14133 & n30778 ;
  assign n30780 = \m4_data_i[11]_pad  & n14140 ;
  assign n30781 = n14157 & n30780 ;
  assign n30782 = ~n30779 & ~n30781 ;
  assign n30783 = n30777 & n30782 ;
  assign n30784 = n30772 & n30783 ;
  assign n30785 = \m0_data_i[12]_pad  & n14140 ;
  assign n30786 = n14165 & n30785 ;
  assign n30787 = \m7_data_i[12]_pad  & ~n14140 ;
  assign n30788 = n14148 & n30787 ;
  assign n30789 = ~n30786 & ~n30788 ;
  assign n30790 = \m1_data_i[12]_pad  & ~n14140 ;
  assign n30791 = n14165 & n30790 ;
  assign n30792 = \m4_data_i[12]_pad  & n14140 ;
  assign n30793 = n14157 & n30792 ;
  assign n30794 = ~n30791 & ~n30793 ;
  assign n30795 = n30789 & n30794 ;
  assign n30796 = \m2_data_i[12]_pad  & n14140 ;
  assign n30797 = n14133 & n30796 ;
  assign n30798 = \m3_data_i[12]_pad  & ~n14140 ;
  assign n30799 = n14133 & n30798 ;
  assign n30800 = ~n30797 & ~n30799 ;
  assign n30801 = \m6_data_i[12]_pad  & n14140 ;
  assign n30802 = n14148 & n30801 ;
  assign n30803 = \m5_data_i[12]_pad  & ~n14140 ;
  assign n30804 = n14157 & n30803 ;
  assign n30805 = ~n30802 & ~n30804 ;
  assign n30806 = n30800 & n30805 ;
  assign n30807 = n30795 & n30806 ;
  assign n30808 = \m1_data_i[13]_pad  & ~n14140 ;
  assign n30809 = n14165 & n30808 ;
  assign n30810 = \m2_data_i[13]_pad  & n14140 ;
  assign n30811 = n14133 & n30810 ;
  assign n30812 = ~n30809 & ~n30811 ;
  assign n30813 = \m0_data_i[13]_pad  & n14140 ;
  assign n30814 = n14165 & n30813 ;
  assign n30815 = \m4_data_i[13]_pad  & n14140 ;
  assign n30816 = n14157 & n30815 ;
  assign n30817 = ~n30814 & ~n30816 ;
  assign n30818 = n30812 & n30817 ;
  assign n30819 = \m7_data_i[13]_pad  & ~n14140 ;
  assign n30820 = n14148 & n30819 ;
  assign n30821 = \m3_data_i[13]_pad  & ~n14140 ;
  assign n30822 = n14133 & n30821 ;
  assign n30823 = ~n30820 & ~n30822 ;
  assign n30824 = \m6_data_i[13]_pad  & n14140 ;
  assign n30825 = n14148 & n30824 ;
  assign n30826 = \m5_data_i[13]_pad  & ~n14140 ;
  assign n30827 = n14157 & n30826 ;
  assign n30828 = ~n30825 & ~n30827 ;
  assign n30829 = n30823 & n30828 ;
  assign n30830 = n30818 & n30829 ;
  assign n30831 = \m3_data_i[14]_pad  & ~n14140 ;
  assign n30832 = n14133 & n30831 ;
  assign n30833 = \m4_data_i[14]_pad  & n14140 ;
  assign n30834 = n14157 & n30833 ;
  assign n30835 = ~n30832 & ~n30834 ;
  assign n30836 = \m6_data_i[14]_pad  & n14140 ;
  assign n30837 = n14148 & n30836 ;
  assign n30838 = \m2_data_i[14]_pad  & n14140 ;
  assign n30839 = n14133 & n30838 ;
  assign n30840 = ~n30837 & ~n30839 ;
  assign n30841 = n30835 & n30840 ;
  assign n30842 = \m5_data_i[14]_pad  & ~n14140 ;
  assign n30843 = n14157 & n30842 ;
  assign n30844 = \m1_data_i[14]_pad  & ~n14140 ;
  assign n30845 = n14165 & n30844 ;
  assign n30846 = ~n30843 & ~n30845 ;
  assign n30847 = \m0_data_i[14]_pad  & n14140 ;
  assign n30848 = n14165 & n30847 ;
  assign n30849 = \m7_data_i[14]_pad  & ~n14140 ;
  assign n30850 = n14148 & n30849 ;
  assign n30851 = ~n30848 & ~n30850 ;
  assign n30852 = n30846 & n30851 ;
  assign n30853 = n30841 & n30852 ;
  assign n30854 = \m0_data_i[15]_pad  & n14140 ;
  assign n30855 = n14165 & n30854 ;
  assign n30856 = \m7_data_i[15]_pad  & ~n14140 ;
  assign n30857 = n14148 & n30856 ;
  assign n30858 = ~n30855 & ~n30857 ;
  assign n30859 = \m6_data_i[15]_pad  & n14140 ;
  assign n30860 = n14148 & n30859 ;
  assign n30861 = \m4_data_i[15]_pad  & n14140 ;
  assign n30862 = n14157 & n30861 ;
  assign n30863 = ~n30860 & ~n30862 ;
  assign n30864 = n30858 & n30863 ;
  assign n30865 = \m5_data_i[15]_pad  & ~n14140 ;
  assign n30866 = n14157 & n30865 ;
  assign n30867 = \m3_data_i[15]_pad  & ~n14140 ;
  assign n30868 = n14133 & n30867 ;
  assign n30869 = ~n30866 & ~n30868 ;
  assign n30870 = \m1_data_i[15]_pad  & ~n14140 ;
  assign n30871 = n14165 & n30870 ;
  assign n30872 = \m2_data_i[15]_pad  & n14140 ;
  assign n30873 = n14133 & n30872 ;
  assign n30874 = ~n30871 & ~n30873 ;
  assign n30875 = n30869 & n30874 ;
  assign n30876 = n30864 & n30875 ;
  assign n30877 = \m6_data_i[16]_pad  & n14140 ;
  assign n30878 = n14148 & n30877 ;
  assign n30879 = \m5_data_i[16]_pad  & ~n14140 ;
  assign n30880 = n14157 & n30879 ;
  assign n30881 = ~n30878 & ~n30880 ;
  assign n30882 = \m3_data_i[16]_pad  & ~n14140 ;
  assign n30883 = n14133 & n30882 ;
  assign n30884 = \m7_data_i[16]_pad  & ~n14140 ;
  assign n30885 = n14148 & n30884 ;
  assign n30886 = ~n30883 & ~n30885 ;
  assign n30887 = n30881 & n30886 ;
  assign n30888 = \m4_data_i[16]_pad  & n14140 ;
  assign n30889 = n14157 & n30888 ;
  assign n30890 = \m0_data_i[16]_pad  & n14140 ;
  assign n30891 = n14165 & n30890 ;
  assign n30892 = ~n30889 & ~n30891 ;
  assign n30893 = \m1_data_i[16]_pad  & ~n14140 ;
  assign n30894 = n14165 & n30893 ;
  assign n30895 = \m2_data_i[16]_pad  & n14140 ;
  assign n30896 = n14133 & n30895 ;
  assign n30897 = ~n30894 & ~n30896 ;
  assign n30898 = n30892 & n30897 ;
  assign n30899 = n30887 & n30898 ;
  assign n30900 = \m1_data_i[17]_pad  & ~n14140 ;
  assign n30901 = n14165 & n30900 ;
  assign n30902 = \m2_data_i[17]_pad  & n14140 ;
  assign n30903 = n14133 & n30902 ;
  assign n30904 = ~n30901 & ~n30903 ;
  assign n30905 = \m0_data_i[17]_pad  & n14140 ;
  assign n30906 = n14165 & n30905 ;
  assign n30907 = \m5_data_i[17]_pad  & ~n14140 ;
  assign n30908 = n14157 & n30907 ;
  assign n30909 = ~n30906 & ~n30908 ;
  assign n30910 = n30904 & n30909 ;
  assign n30911 = \m7_data_i[17]_pad  & ~n14140 ;
  assign n30912 = n14148 & n30911 ;
  assign n30913 = \m6_data_i[17]_pad  & n14140 ;
  assign n30914 = n14148 & n30913 ;
  assign n30915 = ~n30912 & ~n30914 ;
  assign n30916 = \m3_data_i[17]_pad  & ~n14140 ;
  assign n30917 = n14133 & n30916 ;
  assign n30918 = \m4_data_i[17]_pad  & n14140 ;
  assign n30919 = n14157 & n30918 ;
  assign n30920 = ~n30917 & ~n30919 ;
  assign n30921 = n30915 & n30920 ;
  assign n30922 = n30910 & n30921 ;
  assign n30923 = \m1_data_i[18]_pad  & ~n14140 ;
  assign n30924 = n14165 & n30923 ;
  assign n30925 = \m2_data_i[18]_pad  & n14140 ;
  assign n30926 = n14133 & n30925 ;
  assign n30927 = ~n30924 & ~n30926 ;
  assign n30928 = \m0_data_i[18]_pad  & n14140 ;
  assign n30929 = n14165 & n30928 ;
  assign n30930 = \m5_data_i[18]_pad  & ~n14140 ;
  assign n30931 = n14157 & n30930 ;
  assign n30932 = ~n30929 & ~n30931 ;
  assign n30933 = n30927 & n30932 ;
  assign n30934 = \m7_data_i[18]_pad  & ~n14140 ;
  assign n30935 = n14148 & n30934 ;
  assign n30936 = \m6_data_i[18]_pad  & n14140 ;
  assign n30937 = n14148 & n30936 ;
  assign n30938 = ~n30935 & ~n30937 ;
  assign n30939 = \m3_data_i[18]_pad  & ~n14140 ;
  assign n30940 = n14133 & n30939 ;
  assign n30941 = \m4_data_i[18]_pad  & n14140 ;
  assign n30942 = n14157 & n30941 ;
  assign n30943 = ~n30940 & ~n30942 ;
  assign n30944 = n30938 & n30943 ;
  assign n30945 = n30933 & n30944 ;
  assign n30946 = \m1_data_i[19]_pad  & ~n14140 ;
  assign n30947 = n14165 & n30946 ;
  assign n30948 = \m2_data_i[19]_pad  & n14140 ;
  assign n30949 = n14133 & n30948 ;
  assign n30950 = ~n30947 & ~n30949 ;
  assign n30951 = \m0_data_i[19]_pad  & n14140 ;
  assign n30952 = n14165 & n30951 ;
  assign n30953 = \m4_data_i[19]_pad  & n14140 ;
  assign n30954 = n14157 & n30953 ;
  assign n30955 = ~n30952 & ~n30954 ;
  assign n30956 = n30950 & n30955 ;
  assign n30957 = \m7_data_i[19]_pad  & ~n14140 ;
  assign n30958 = n14148 & n30957 ;
  assign n30959 = \m3_data_i[19]_pad  & ~n14140 ;
  assign n30960 = n14133 & n30959 ;
  assign n30961 = ~n30958 & ~n30960 ;
  assign n30962 = \m6_data_i[19]_pad  & n14140 ;
  assign n30963 = n14148 & n30962 ;
  assign n30964 = \m5_data_i[19]_pad  & ~n14140 ;
  assign n30965 = n14157 & n30964 ;
  assign n30966 = ~n30963 & ~n30965 ;
  assign n30967 = n30961 & n30966 ;
  assign n30968 = n30956 & n30967 ;
  assign n30969 = \m3_data_i[1]_pad  & ~n14140 ;
  assign n30970 = n14133 & n30969 ;
  assign n30971 = \m4_data_i[1]_pad  & n14140 ;
  assign n30972 = n14157 & n30971 ;
  assign n30973 = ~n30970 & ~n30972 ;
  assign n30974 = \m1_data_i[1]_pad  & ~n14140 ;
  assign n30975 = n14165 & n30974 ;
  assign n30976 = \m7_data_i[1]_pad  & ~n14140 ;
  assign n30977 = n14148 & n30976 ;
  assign n30978 = ~n30975 & ~n30977 ;
  assign n30979 = n30973 & n30978 ;
  assign n30980 = \m2_data_i[1]_pad  & n14140 ;
  assign n30981 = n14133 & n30980 ;
  assign n30982 = \m0_data_i[1]_pad  & n14140 ;
  assign n30983 = n14165 & n30982 ;
  assign n30984 = ~n30981 & ~n30983 ;
  assign n30985 = \m6_data_i[1]_pad  & n14140 ;
  assign n30986 = n14148 & n30985 ;
  assign n30987 = \m5_data_i[1]_pad  & ~n14140 ;
  assign n30988 = n14157 & n30987 ;
  assign n30989 = ~n30986 & ~n30988 ;
  assign n30990 = n30984 & n30989 ;
  assign n30991 = n30979 & n30990 ;
  assign n30992 = \m6_data_i[20]_pad  & n14140 ;
  assign n30993 = n14148 & n30992 ;
  assign n30994 = \m5_data_i[20]_pad  & ~n14140 ;
  assign n30995 = n14157 & n30994 ;
  assign n30996 = ~n30993 & ~n30995 ;
  assign n30997 = \m0_data_i[20]_pad  & n14140 ;
  assign n30998 = n14165 & n30997 ;
  assign n30999 = \m4_data_i[20]_pad  & n14140 ;
  assign n31000 = n14157 & n30999 ;
  assign n31001 = ~n30998 & ~n31000 ;
  assign n31002 = n30996 & n31001 ;
  assign n31003 = \m7_data_i[20]_pad  & ~n14140 ;
  assign n31004 = n14148 & n31003 ;
  assign n31005 = \m3_data_i[20]_pad  & ~n14140 ;
  assign n31006 = n14133 & n31005 ;
  assign n31007 = ~n31004 & ~n31006 ;
  assign n31008 = \m1_data_i[20]_pad  & ~n14140 ;
  assign n31009 = n14165 & n31008 ;
  assign n31010 = \m2_data_i[20]_pad  & n14140 ;
  assign n31011 = n14133 & n31010 ;
  assign n31012 = ~n31009 & ~n31011 ;
  assign n31013 = n31007 & n31012 ;
  assign n31014 = n31002 & n31013 ;
  assign n31015 = \m3_data_i[21]_pad  & ~n14140 ;
  assign n31016 = n14133 & n31015 ;
  assign n31017 = \m4_data_i[21]_pad  & n14140 ;
  assign n31018 = n14157 & n31017 ;
  assign n31019 = ~n31016 & ~n31018 ;
  assign n31020 = \m1_data_i[21]_pad  & ~n14140 ;
  assign n31021 = n14165 & n31020 ;
  assign n31022 = \m5_data_i[21]_pad  & ~n14140 ;
  assign n31023 = n14157 & n31022 ;
  assign n31024 = ~n31021 & ~n31023 ;
  assign n31025 = n31019 & n31024 ;
  assign n31026 = \m2_data_i[21]_pad  & n14140 ;
  assign n31027 = n14133 & n31026 ;
  assign n31028 = \m6_data_i[21]_pad  & n14140 ;
  assign n31029 = n14148 & n31028 ;
  assign n31030 = ~n31027 & ~n31029 ;
  assign n31031 = \m0_data_i[21]_pad  & n14140 ;
  assign n31032 = n14165 & n31031 ;
  assign n31033 = \m7_data_i[21]_pad  & ~n14140 ;
  assign n31034 = n14148 & n31033 ;
  assign n31035 = ~n31032 & ~n31034 ;
  assign n31036 = n31030 & n31035 ;
  assign n31037 = n31025 & n31036 ;
  assign n31038 = \m6_data_i[22]_pad  & n14140 ;
  assign n31039 = n14148 & n31038 ;
  assign n31040 = \m5_data_i[22]_pad  & ~n14140 ;
  assign n31041 = n14157 & n31040 ;
  assign n31042 = ~n31039 & ~n31041 ;
  assign n31043 = \m3_data_i[22]_pad  & ~n14140 ;
  assign n31044 = n14133 & n31043 ;
  assign n31045 = \m2_data_i[22]_pad  & n14140 ;
  assign n31046 = n14133 & n31045 ;
  assign n31047 = ~n31044 & ~n31046 ;
  assign n31048 = n31042 & n31047 ;
  assign n31049 = \m4_data_i[22]_pad  & n14140 ;
  assign n31050 = n14157 & n31049 ;
  assign n31051 = \m1_data_i[22]_pad  & ~n14140 ;
  assign n31052 = n14165 & n31051 ;
  assign n31053 = ~n31050 & ~n31052 ;
  assign n31054 = \m0_data_i[22]_pad  & n14140 ;
  assign n31055 = n14165 & n31054 ;
  assign n31056 = \m7_data_i[22]_pad  & ~n14140 ;
  assign n31057 = n14148 & n31056 ;
  assign n31058 = ~n31055 & ~n31057 ;
  assign n31059 = n31053 & n31058 ;
  assign n31060 = n31048 & n31059 ;
  assign n31061 = \m6_data_i[23]_pad  & n14140 ;
  assign n31062 = n14148 & n31061 ;
  assign n31063 = \m5_data_i[23]_pad  & ~n14140 ;
  assign n31064 = n14157 & n31063 ;
  assign n31065 = ~n31062 & ~n31064 ;
  assign n31066 = \m0_data_i[23]_pad  & n14140 ;
  assign n31067 = n14165 & n31066 ;
  assign n31068 = \m2_data_i[23]_pad  & n14140 ;
  assign n31069 = n14133 & n31068 ;
  assign n31070 = ~n31067 & ~n31069 ;
  assign n31071 = n31065 & n31070 ;
  assign n31072 = \m7_data_i[23]_pad  & ~n14140 ;
  assign n31073 = n14148 & n31072 ;
  assign n31074 = \m1_data_i[23]_pad  & ~n14140 ;
  assign n31075 = n14165 & n31074 ;
  assign n31076 = ~n31073 & ~n31075 ;
  assign n31077 = \m3_data_i[23]_pad  & ~n14140 ;
  assign n31078 = n14133 & n31077 ;
  assign n31079 = \m4_data_i[23]_pad  & n14140 ;
  assign n31080 = n14157 & n31079 ;
  assign n31081 = ~n31078 & ~n31080 ;
  assign n31082 = n31076 & n31081 ;
  assign n31083 = n31071 & n31082 ;
  assign n31084 = \m6_data_i[24]_pad  & n14140 ;
  assign n31085 = n14148 & n31084 ;
  assign n31086 = \m5_data_i[24]_pad  & ~n14140 ;
  assign n31087 = n14157 & n31086 ;
  assign n31088 = ~n31085 & ~n31087 ;
  assign n31089 = \m1_data_i[24]_pad  & ~n14140 ;
  assign n31090 = n14165 & n31089 ;
  assign n31091 = \m7_data_i[24]_pad  & ~n14140 ;
  assign n31092 = n14148 & n31091 ;
  assign n31093 = ~n31090 & ~n31092 ;
  assign n31094 = n31088 & n31093 ;
  assign n31095 = \m2_data_i[24]_pad  & n14140 ;
  assign n31096 = n14133 & n31095 ;
  assign n31097 = \m0_data_i[24]_pad  & n14140 ;
  assign n31098 = n14165 & n31097 ;
  assign n31099 = ~n31096 & ~n31098 ;
  assign n31100 = \m3_data_i[24]_pad  & ~n14140 ;
  assign n31101 = n14133 & n31100 ;
  assign n31102 = \m4_data_i[24]_pad  & n14140 ;
  assign n31103 = n14157 & n31102 ;
  assign n31104 = ~n31101 & ~n31103 ;
  assign n31105 = n31099 & n31104 ;
  assign n31106 = n31094 & n31105 ;
  assign n31107 = \m3_data_i[25]_pad  & ~n14140 ;
  assign n31108 = n14133 & n31107 ;
  assign n31109 = \m4_data_i[25]_pad  & n14140 ;
  assign n31110 = n14157 & n31109 ;
  assign n31111 = ~n31108 & ~n31110 ;
  assign n31112 = \m0_data_i[25]_pad  & n14140 ;
  assign n31113 = n14165 & n31112 ;
  assign n31114 = \m2_data_i[25]_pad  & n14140 ;
  assign n31115 = n14133 & n31114 ;
  assign n31116 = ~n31113 & ~n31115 ;
  assign n31117 = n31111 & n31116 ;
  assign n31118 = \m7_data_i[25]_pad  & ~n14140 ;
  assign n31119 = n14148 & n31118 ;
  assign n31120 = \m1_data_i[25]_pad  & ~n14140 ;
  assign n31121 = n14165 & n31120 ;
  assign n31122 = ~n31119 & ~n31121 ;
  assign n31123 = \m6_data_i[25]_pad  & n14140 ;
  assign n31124 = n14148 & n31123 ;
  assign n31125 = \m5_data_i[25]_pad  & ~n14140 ;
  assign n31126 = n14157 & n31125 ;
  assign n31127 = ~n31124 & ~n31126 ;
  assign n31128 = n31122 & n31127 ;
  assign n31129 = n31117 & n31128 ;
  assign n31130 = \m1_data_i[26]_pad  & ~n14140 ;
  assign n31131 = n14165 & n31130 ;
  assign n31132 = \m2_data_i[26]_pad  & n14140 ;
  assign n31133 = n14133 & n31132 ;
  assign n31134 = ~n31131 & ~n31133 ;
  assign n31135 = \m0_data_i[26]_pad  & n14140 ;
  assign n31136 = n14165 & n31135 ;
  assign n31137 = \m5_data_i[26]_pad  & ~n14140 ;
  assign n31138 = n14157 & n31137 ;
  assign n31139 = ~n31136 & ~n31138 ;
  assign n31140 = n31134 & n31139 ;
  assign n31141 = \m7_data_i[26]_pad  & ~n14140 ;
  assign n31142 = n14148 & n31141 ;
  assign n31143 = \m6_data_i[26]_pad  & n14140 ;
  assign n31144 = n14148 & n31143 ;
  assign n31145 = ~n31142 & ~n31144 ;
  assign n31146 = \m3_data_i[26]_pad  & ~n14140 ;
  assign n31147 = n14133 & n31146 ;
  assign n31148 = \m4_data_i[26]_pad  & n14140 ;
  assign n31149 = n14157 & n31148 ;
  assign n31150 = ~n31147 & ~n31149 ;
  assign n31151 = n31145 & n31150 ;
  assign n31152 = n31140 & n31151 ;
  assign n31153 = \m1_data_i[27]_pad  & ~n14140 ;
  assign n31154 = n14165 & n31153 ;
  assign n31155 = \m2_data_i[27]_pad  & n14140 ;
  assign n31156 = n14133 & n31155 ;
  assign n31157 = ~n31154 & ~n31156 ;
  assign n31158 = \m3_data_i[27]_pad  & ~n14140 ;
  assign n31159 = n14133 & n31158 ;
  assign n31160 = \m7_data_i[27]_pad  & ~n14140 ;
  assign n31161 = n14148 & n31160 ;
  assign n31162 = ~n31159 & ~n31161 ;
  assign n31163 = n31157 & n31162 ;
  assign n31164 = \m4_data_i[27]_pad  & n14140 ;
  assign n31165 = n14157 & n31164 ;
  assign n31166 = \m0_data_i[27]_pad  & n14140 ;
  assign n31167 = n14165 & n31166 ;
  assign n31168 = ~n31165 & ~n31167 ;
  assign n31169 = \m6_data_i[27]_pad  & n14140 ;
  assign n31170 = n14148 & n31169 ;
  assign n31171 = \m5_data_i[27]_pad  & ~n14140 ;
  assign n31172 = n14157 & n31171 ;
  assign n31173 = ~n31170 & ~n31172 ;
  assign n31174 = n31168 & n31173 ;
  assign n31175 = n31163 & n31174 ;
  assign n31176 = \m3_data_i[28]_pad  & ~n14140 ;
  assign n31177 = n14133 & n31176 ;
  assign n31178 = \m4_data_i[28]_pad  & n14140 ;
  assign n31179 = n14157 & n31178 ;
  assign n31180 = ~n31177 & ~n31179 ;
  assign n31181 = \m6_data_i[28]_pad  & n14140 ;
  assign n31182 = n14148 & n31181 ;
  assign n31183 = \m2_data_i[28]_pad  & n14140 ;
  assign n31184 = n14133 & n31183 ;
  assign n31185 = ~n31182 & ~n31184 ;
  assign n31186 = n31180 & n31185 ;
  assign n31187 = \m5_data_i[28]_pad  & ~n14140 ;
  assign n31188 = n14157 & n31187 ;
  assign n31189 = \m1_data_i[28]_pad  & ~n14140 ;
  assign n31190 = n14165 & n31189 ;
  assign n31191 = ~n31188 & ~n31190 ;
  assign n31192 = \m0_data_i[28]_pad  & n14140 ;
  assign n31193 = n14165 & n31192 ;
  assign n31194 = \m7_data_i[28]_pad  & ~n14140 ;
  assign n31195 = n14148 & n31194 ;
  assign n31196 = ~n31193 & ~n31195 ;
  assign n31197 = n31191 & n31196 ;
  assign n31198 = n31186 & n31197 ;
  assign n31199 = \m6_data_i[29]_pad  & n14140 ;
  assign n31200 = n14148 & n31199 ;
  assign n31201 = \m5_data_i[29]_pad  & ~n14140 ;
  assign n31202 = n14157 & n31201 ;
  assign n31203 = ~n31200 & ~n31202 ;
  assign n31204 = \m0_data_i[29]_pad  & n14140 ;
  assign n31205 = n14165 & n31204 ;
  assign n31206 = \m2_data_i[29]_pad  & n14140 ;
  assign n31207 = n14133 & n31206 ;
  assign n31208 = ~n31205 & ~n31207 ;
  assign n31209 = n31203 & n31208 ;
  assign n31210 = \m7_data_i[29]_pad  & ~n14140 ;
  assign n31211 = n14148 & n31210 ;
  assign n31212 = \m1_data_i[29]_pad  & ~n14140 ;
  assign n31213 = n14165 & n31212 ;
  assign n31214 = ~n31211 & ~n31213 ;
  assign n31215 = \m3_data_i[29]_pad  & ~n14140 ;
  assign n31216 = n14133 & n31215 ;
  assign n31217 = \m4_data_i[29]_pad  & n14140 ;
  assign n31218 = n14157 & n31217 ;
  assign n31219 = ~n31216 & ~n31218 ;
  assign n31220 = n31214 & n31219 ;
  assign n31221 = n31209 & n31220 ;
  assign n31222 = \m1_data_i[2]_pad  & ~n14140 ;
  assign n31223 = n14165 & n31222 ;
  assign n31224 = \m2_data_i[2]_pad  & n14140 ;
  assign n31225 = n14133 & n31224 ;
  assign n31226 = ~n31223 & ~n31225 ;
  assign n31227 = \m0_data_i[2]_pad  & n14140 ;
  assign n31228 = n14165 & n31227 ;
  assign n31229 = \m5_data_i[2]_pad  & ~n14140 ;
  assign n31230 = n14157 & n31229 ;
  assign n31231 = ~n31228 & ~n31230 ;
  assign n31232 = n31226 & n31231 ;
  assign n31233 = \m7_data_i[2]_pad  & ~n14140 ;
  assign n31234 = n14148 & n31233 ;
  assign n31235 = \m6_data_i[2]_pad  & n14140 ;
  assign n31236 = n14148 & n31235 ;
  assign n31237 = ~n31234 & ~n31236 ;
  assign n31238 = \m3_data_i[2]_pad  & ~n14140 ;
  assign n31239 = n14133 & n31238 ;
  assign n31240 = \m4_data_i[2]_pad  & n14140 ;
  assign n31241 = n14157 & n31240 ;
  assign n31242 = ~n31239 & ~n31241 ;
  assign n31243 = n31237 & n31242 ;
  assign n31244 = n31232 & n31243 ;
  assign n31245 = \m3_data_i[30]_pad  & ~n14140 ;
  assign n31246 = n14133 & n31245 ;
  assign n31247 = \m4_data_i[30]_pad  & n14140 ;
  assign n31248 = n14157 & n31247 ;
  assign n31249 = ~n31246 & ~n31248 ;
  assign n31250 = \m0_data_i[30]_pad  & n14140 ;
  assign n31251 = n14165 & n31250 ;
  assign n31252 = \m5_data_i[30]_pad  & ~n14140 ;
  assign n31253 = n14157 & n31252 ;
  assign n31254 = ~n31251 & ~n31253 ;
  assign n31255 = n31249 & n31254 ;
  assign n31256 = \m7_data_i[30]_pad  & ~n14140 ;
  assign n31257 = n14148 & n31256 ;
  assign n31258 = \m6_data_i[30]_pad  & n14140 ;
  assign n31259 = n14148 & n31258 ;
  assign n31260 = ~n31257 & ~n31259 ;
  assign n31261 = \m1_data_i[30]_pad  & ~n14140 ;
  assign n31262 = n14165 & n31261 ;
  assign n31263 = \m2_data_i[30]_pad  & n14140 ;
  assign n31264 = n14133 & n31263 ;
  assign n31265 = ~n31262 & ~n31264 ;
  assign n31266 = n31260 & n31265 ;
  assign n31267 = n31255 & n31266 ;
  assign n31268 = \m1_data_i[31]_pad  & ~n14140 ;
  assign n31269 = n14165 & n31268 ;
  assign n31270 = \m2_data_i[31]_pad  & n14140 ;
  assign n31271 = n14133 & n31270 ;
  assign n31272 = ~n31269 & ~n31271 ;
  assign n31273 = \m0_data_i[31]_pad  & n14140 ;
  assign n31274 = n14165 & n31273 ;
  assign n31275 = \m4_data_i[31]_pad  & n14140 ;
  assign n31276 = n14157 & n31275 ;
  assign n31277 = ~n31274 & ~n31276 ;
  assign n31278 = n31272 & n31277 ;
  assign n31279 = \m7_data_i[31]_pad  & ~n14140 ;
  assign n31280 = n14148 & n31279 ;
  assign n31281 = \m3_data_i[31]_pad  & ~n14140 ;
  assign n31282 = n14133 & n31281 ;
  assign n31283 = ~n31280 & ~n31282 ;
  assign n31284 = \m6_data_i[31]_pad  & n14140 ;
  assign n31285 = n14148 & n31284 ;
  assign n31286 = \m5_data_i[31]_pad  & ~n14140 ;
  assign n31287 = n14157 & n31286 ;
  assign n31288 = ~n31285 & ~n31287 ;
  assign n31289 = n31283 & n31288 ;
  assign n31290 = n31278 & n31289 ;
  assign n31291 = \m6_data_i[3]_pad  & n14140 ;
  assign n31292 = n14148 & n31291 ;
  assign n31293 = \m5_data_i[3]_pad  & ~n14140 ;
  assign n31294 = n14157 & n31293 ;
  assign n31295 = ~n31292 & ~n31294 ;
  assign n31296 = \m1_data_i[3]_pad  & ~n14140 ;
  assign n31297 = n14165 & n31296 ;
  assign n31298 = \m4_data_i[3]_pad  & n14140 ;
  assign n31299 = n14157 & n31298 ;
  assign n31300 = ~n31297 & ~n31299 ;
  assign n31301 = n31295 & n31300 ;
  assign n31302 = \m2_data_i[3]_pad  & n14140 ;
  assign n31303 = n14133 & n31302 ;
  assign n31304 = \m3_data_i[3]_pad  & ~n14140 ;
  assign n31305 = n14133 & n31304 ;
  assign n31306 = ~n31303 & ~n31305 ;
  assign n31307 = \m0_data_i[3]_pad  & n14140 ;
  assign n31308 = n14165 & n31307 ;
  assign n31309 = \m7_data_i[3]_pad  & ~n14140 ;
  assign n31310 = n14148 & n31309 ;
  assign n31311 = ~n31308 & ~n31310 ;
  assign n31312 = n31306 & n31311 ;
  assign n31313 = n31301 & n31312 ;
  assign n31314 = \m1_data_i[4]_pad  & ~n14140 ;
  assign n31315 = n14165 & n31314 ;
  assign n31316 = \m2_data_i[4]_pad  & n14140 ;
  assign n31317 = n14133 & n31316 ;
  assign n31318 = ~n31315 & ~n31317 ;
  assign n31319 = \m0_data_i[4]_pad  & n14140 ;
  assign n31320 = n14165 & n31319 ;
  assign n31321 = \m4_data_i[4]_pad  & n14140 ;
  assign n31322 = n14157 & n31321 ;
  assign n31323 = ~n31320 & ~n31322 ;
  assign n31324 = n31318 & n31323 ;
  assign n31325 = \m7_data_i[4]_pad  & ~n14140 ;
  assign n31326 = n14148 & n31325 ;
  assign n31327 = \m3_data_i[4]_pad  & ~n14140 ;
  assign n31328 = n14133 & n31327 ;
  assign n31329 = ~n31326 & ~n31328 ;
  assign n31330 = \m6_data_i[4]_pad  & n14140 ;
  assign n31331 = n14148 & n31330 ;
  assign n31332 = \m5_data_i[4]_pad  & ~n14140 ;
  assign n31333 = n14157 & n31332 ;
  assign n31334 = ~n31331 & ~n31333 ;
  assign n31335 = n31329 & n31334 ;
  assign n31336 = n31324 & n31335 ;
  assign n31337 = \m3_data_i[5]_pad  & ~n14140 ;
  assign n31338 = n14133 & n31337 ;
  assign n31339 = \m4_data_i[5]_pad  & n14140 ;
  assign n31340 = n14157 & n31339 ;
  assign n31341 = ~n31338 & ~n31340 ;
  assign n31342 = \m0_data_i[5]_pad  & n14140 ;
  assign n31343 = n14165 & n31342 ;
  assign n31344 = \m2_data_i[5]_pad  & n14140 ;
  assign n31345 = n14133 & n31344 ;
  assign n31346 = ~n31343 & ~n31345 ;
  assign n31347 = n31341 & n31346 ;
  assign n31348 = \m7_data_i[5]_pad  & ~n14140 ;
  assign n31349 = n14148 & n31348 ;
  assign n31350 = \m1_data_i[5]_pad  & ~n14140 ;
  assign n31351 = n14165 & n31350 ;
  assign n31352 = ~n31349 & ~n31351 ;
  assign n31353 = \m6_data_i[5]_pad  & n14140 ;
  assign n31354 = n14148 & n31353 ;
  assign n31355 = \m5_data_i[5]_pad  & ~n14140 ;
  assign n31356 = n14157 & n31355 ;
  assign n31357 = ~n31354 & ~n31356 ;
  assign n31358 = n31352 & n31357 ;
  assign n31359 = n31347 & n31358 ;
  assign n31360 = \m3_data_i[6]_pad  & ~n14140 ;
  assign n31361 = n14133 & n31360 ;
  assign n31362 = \m4_data_i[6]_pad  & n14140 ;
  assign n31363 = n14157 & n31362 ;
  assign n31364 = ~n31361 & ~n31363 ;
  assign n31365 = \m6_data_i[6]_pad  & n14140 ;
  assign n31366 = n14148 & n31365 ;
  assign n31367 = \m7_data_i[6]_pad  & ~n14140 ;
  assign n31368 = n14148 & n31367 ;
  assign n31369 = ~n31366 & ~n31368 ;
  assign n31370 = n31364 & n31369 ;
  assign n31371 = \m5_data_i[6]_pad  & ~n14140 ;
  assign n31372 = n14157 & n31371 ;
  assign n31373 = \m0_data_i[6]_pad  & n14140 ;
  assign n31374 = n14165 & n31373 ;
  assign n31375 = ~n31372 & ~n31374 ;
  assign n31376 = \m1_data_i[6]_pad  & ~n14140 ;
  assign n31377 = n14165 & n31376 ;
  assign n31378 = \m2_data_i[6]_pad  & n14140 ;
  assign n31379 = n14133 & n31378 ;
  assign n31380 = ~n31377 & ~n31379 ;
  assign n31381 = n31375 & n31380 ;
  assign n31382 = n31370 & n31381 ;
  assign n31383 = \m3_data_i[7]_pad  & ~n14140 ;
  assign n31384 = n14133 & n31383 ;
  assign n31385 = \m4_data_i[7]_pad  & n14140 ;
  assign n31386 = n14157 & n31385 ;
  assign n31387 = ~n31384 & ~n31386 ;
  assign n31388 = \m0_data_i[7]_pad  & n14140 ;
  assign n31389 = n14165 & n31388 ;
  assign n31390 = \m2_data_i[7]_pad  & n14140 ;
  assign n31391 = n14133 & n31390 ;
  assign n31392 = ~n31389 & ~n31391 ;
  assign n31393 = n31387 & n31392 ;
  assign n31394 = \m7_data_i[7]_pad  & ~n14140 ;
  assign n31395 = n14148 & n31394 ;
  assign n31396 = \m1_data_i[7]_pad  & ~n14140 ;
  assign n31397 = n14165 & n31396 ;
  assign n31398 = ~n31395 & ~n31397 ;
  assign n31399 = \m6_data_i[7]_pad  & n14140 ;
  assign n31400 = n14148 & n31399 ;
  assign n31401 = \m5_data_i[7]_pad  & ~n14140 ;
  assign n31402 = n14157 & n31401 ;
  assign n31403 = ~n31400 & ~n31402 ;
  assign n31404 = n31398 & n31403 ;
  assign n31405 = n31393 & n31404 ;
  assign n31406 = \m1_data_i[8]_pad  & ~n14140 ;
  assign n31407 = n14165 & n31406 ;
  assign n31408 = \m2_data_i[8]_pad  & n14140 ;
  assign n31409 = n14133 & n31408 ;
  assign n31410 = ~n31407 & ~n31409 ;
  assign n31411 = \m0_data_i[8]_pad  & n14140 ;
  assign n31412 = n14165 & n31411 ;
  assign n31413 = \m4_data_i[8]_pad  & n14140 ;
  assign n31414 = n14157 & n31413 ;
  assign n31415 = ~n31412 & ~n31414 ;
  assign n31416 = n31410 & n31415 ;
  assign n31417 = \m7_data_i[8]_pad  & ~n14140 ;
  assign n31418 = n14148 & n31417 ;
  assign n31419 = \m3_data_i[8]_pad  & ~n14140 ;
  assign n31420 = n14133 & n31419 ;
  assign n31421 = ~n31418 & ~n31420 ;
  assign n31422 = \m6_data_i[8]_pad  & n14140 ;
  assign n31423 = n14148 & n31422 ;
  assign n31424 = \m5_data_i[8]_pad  & ~n14140 ;
  assign n31425 = n14157 & n31424 ;
  assign n31426 = ~n31423 & ~n31425 ;
  assign n31427 = n31421 & n31426 ;
  assign n31428 = n31416 & n31427 ;
  assign n31429 = \m1_data_i[9]_pad  & ~n14140 ;
  assign n31430 = n14165 & n31429 ;
  assign n31431 = \m2_data_i[9]_pad  & n14140 ;
  assign n31432 = n14133 & n31431 ;
  assign n31433 = ~n31430 & ~n31432 ;
  assign n31434 = \m0_data_i[9]_pad  & n14140 ;
  assign n31435 = n14165 & n31434 ;
  assign n31436 = \m4_data_i[9]_pad  & n14140 ;
  assign n31437 = n14157 & n31436 ;
  assign n31438 = ~n31435 & ~n31437 ;
  assign n31439 = n31433 & n31438 ;
  assign n31440 = \m7_data_i[9]_pad  & ~n14140 ;
  assign n31441 = n14148 & n31440 ;
  assign n31442 = \m3_data_i[9]_pad  & ~n14140 ;
  assign n31443 = n14133 & n31442 ;
  assign n31444 = ~n31441 & ~n31443 ;
  assign n31445 = \m6_data_i[9]_pad  & n14140 ;
  assign n31446 = n14148 & n31445 ;
  assign n31447 = \m5_data_i[9]_pad  & ~n14140 ;
  assign n31448 = n14157 & n31447 ;
  assign n31449 = ~n31446 & ~n31448 ;
  assign n31450 = n31444 & n31449 ;
  assign n31451 = n31439 & n31450 ;
  assign n31452 = \m3_sel_i[0]_pad  & ~n14140 ;
  assign n31453 = n14133 & n31452 ;
  assign n31454 = \m4_sel_i[0]_pad  & n14140 ;
  assign n31455 = n14157 & n31454 ;
  assign n31456 = ~n31453 & ~n31455 ;
  assign n31457 = \m6_sel_i[0]_pad  & n14140 ;
  assign n31458 = n14148 & n31457 ;
  assign n31459 = \m2_sel_i[0]_pad  & n14140 ;
  assign n31460 = n14133 & n31459 ;
  assign n31461 = ~n31458 & ~n31460 ;
  assign n31462 = n31456 & n31461 ;
  assign n31463 = \m5_sel_i[0]_pad  & ~n14140 ;
  assign n31464 = n14157 & n31463 ;
  assign n31465 = \m1_sel_i[0]_pad  & ~n14140 ;
  assign n31466 = n14165 & n31465 ;
  assign n31467 = ~n31464 & ~n31466 ;
  assign n31468 = \m0_sel_i[0]_pad  & n14140 ;
  assign n31469 = n14165 & n31468 ;
  assign n31470 = \m7_sel_i[0]_pad  & ~n14140 ;
  assign n31471 = n14148 & n31470 ;
  assign n31472 = ~n31469 & ~n31471 ;
  assign n31473 = n31467 & n31472 ;
  assign n31474 = n31462 & n31473 ;
  assign n31475 = \m3_sel_i[1]_pad  & ~n14140 ;
  assign n31476 = n14133 & n31475 ;
  assign n31477 = \m4_sel_i[1]_pad  & n14140 ;
  assign n31478 = n14157 & n31477 ;
  assign n31479 = ~n31476 & ~n31478 ;
  assign n31480 = \m6_sel_i[1]_pad  & n14140 ;
  assign n31481 = n14148 & n31480 ;
  assign n31482 = \m2_sel_i[1]_pad  & n14140 ;
  assign n31483 = n14133 & n31482 ;
  assign n31484 = ~n31481 & ~n31483 ;
  assign n31485 = n31479 & n31484 ;
  assign n31486 = \m5_sel_i[1]_pad  & ~n14140 ;
  assign n31487 = n14157 & n31486 ;
  assign n31488 = \m1_sel_i[1]_pad  & ~n14140 ;
  assign n31489 = n14165 & n31488 ;
  assign n31490 = ~n31487 & ~n31489 ;
  assign n31491 = \m0_sel_i[1]_pad  & n14140 ;
  assign n31492 = n14165 & n31491 ;
  assign n31493 = \m7_sel_i[1]_pad  & ~n14140 ;
  assign n31494 = n14148 & n31493 ;
  assign n31495 = ~n31492 & ~n31494 ;
  assign n31496 = n31490 & n31495 ;
  assign n31497 = n31485 & n31496 ;
  assign n31498 = \m3_sel_i[2]_pad  & ~n14140 ;
  assign n31499 = n14133 & n31498 ;
  assign n31500 = \m4_sel_i[2]_pad  & n14140 ;
  assign n31501 = n14157 & n31500 ;
  assign n31502 = ~n31499 & ~n31501 ;
  assign n31503 = \m6_sel_i[2]_pad  & n14140 ;
  assign n31504 = n14148 & n31503 ;
  assign n31505 = \m2_sel_i[2]_pad  & n14140 ;
  assign n31506 = n14133 & n31505 ;
  assign n31507 = ~n31504 & ~n31506 ;
  assign n31508 = n31502 & n31507 ;
  assign n31509 = \m5_sel_i[2]_pad  & ~n14140 ;
  assign n31510 = n14157 & n31509 ;
  assign n31511 = \m1_sel_i[2]_pad  & ~n14140 ;
  assign n31512 = n14165 & n31511 ;
  assign n31513 = ~n31510 & ~n31512 ;
  assign n31514 = \m0_sel_i[2]_pad  & n14140 ;
  assign n31515 = n14165 & n31514 ;
  assign n31516 = \m7_sel_i[2]_pad  & ~n14140 ;
  assign n31517 = n14148 & n31516 ;
  assign n31518 = ~n31515 & ~n31517 ;
  assign n31519 = n31513 & n31518 ;
  assign n31520 = n31508 & n31519 ;
  assign n31521 = \m3_sel_i[3]_pad  & ~n14140 ;
  assign n31522 = n14133 & n31521 ;
  assign n31523 = \m4_sel_i[3]_pad  & n14140 ;
  assign n31524 = n14157 & n31523 ;
  assign n31525 = ~n31522 & ~n31524 ;
  assign n31526 = \m6_sel_i[3]_pad  & n14140 ;
  assign n31527 = n14148 & n31526 ;
  assign n31528 = \m2_sel_i[3]_pad  & n14140 ;
  assign n31529 = n14133 & n31528 ;
  assign n31530 = ~n31527 & ~n31529 ;
  assign n31531 = n31525 & n31530 ;
  assign n31532 = \m5_sel_i[3]_pad  & ~n14140 ;
  assign n31533 = n14157 & n31532 ;
  assign n31534 = \m1_sel_i[3]_pad  & ~n14140 ;
  assign n31535 = n14165 & n31534 ;
  assign n31536 = ~n31533 & ~n31535 ;
  assign n31537 = \m0_sel_i[3]_pad  & n14140 ;
  assign n31538 = n14165 & n31537 ;
  assign n31539 = \m7_sel_i[3]_pad  & ~n14140 ;
  assign n31540 = n14148 & n31539 ;
  assign n31541 = ~n31538 & ~n31540 ;
  assign n31542 = n31536 & n31541 ;
  assign n31543 = n31531 & n31542 ;
  assign n31544 = \m7_stb_i_pad  & n14685 ;
  assign n31545 = ~n14140 & n31544 ;
  assign n31546 = n14148 & n31545 ;
  assign n31547 = \m6_stb_i_pad  & n15007 ;
  assign n31548 = n14140 & n31547 ;
  assign n31549 = n14148 & n31548 ;
  assign n31550 = ~n31546 & ~n31549 ;
  assign n31551 = \m4_stb_i_pad  & n14935 ;
  assign n31552 = n14140 & n31551 ;
  assign n31553 = n14157 & n31552 ;
  assign n31554 = \m1_stb_i_pad  & n15102 ;
  assign n31555 = ~n14140 & n31554 ;
  assign n31556 = n14165 & n31555 ;
  assign n31557 = ~n31553 & ~n31556 ;
  assign n31558 = n31550 & n31557 ;
  assign n31559 = \m5_stb_i_pad  & n14708 ;
  assign n31560 = ~n14140 & n31559 ;
  assign n31561 = n14157 & n31560 ;
  assign n31562 = \m3_stb_i_pad  & n14900 ;
  assign n31563 = ~n14140 & n31562 ;
  assign n31564 = n14133 & n31563 ;
  assign n31565 = ~n31561 & ~n31564 ;
  assign n31566 = \m2_stb_i_pad  & n14859 ;
  assign n31567 = n14140 & n31566 ;
  assign n31568 = n14133 & n31567 ;
  assign n31569 = \m0_stb_i_pad  & n15122 ;
  assign n31570 = n14140 & n31569 ;
  assign n31571 = n14165 & n31570 ;
  assign n31572 = ~n31568 & ~n31571 ;
  assign n31573 = n31565 & n31572 ;
  assign n31574 = n31558 & n31573 ;
  assign n31575 = \m3_we_i_pad  & ~n14140 ;
  assign n31576 = n14133 & n31575 ;
  assign n31577 = \m4_we_i_pad  & n14140 ;
  assign n31578 = n14157 & n31577 ;
  assign n31579 = ~n31576 & ~n31578 ;
  assign n31580 = \m6_we_i_pad  & n14140 ;
  assign n31581 = n14148 & n31580 ;
  assign n31582 = \m2_we_i_pad  & n14140 ;
  assign n31583 = n14133 & n31582 ;
  assign n31584 = ~n31581 & ~n31583 ;
  assign n31585 = n31579 & n31584 ;
  assign n31586 = \m5_we_i_pad  & ~n14140 ;
  assign n31587 = n14157 & n31586 ;
  assign n31588 = \m1_we_i_pad  & ~n14140 ;
  assign n31589 = n14165 & n31588 ;
  assign n31590 = ~n31587 & ~n31589 ;
  assign n31591 = \m0_we_i_pad  & n14140 ;
  assign n31592 = n14165 & n31591 ;
  assign n31593 = \m7_we_i_pad  & ~n14140 ;
  assign n31594 = n14148 & n31593 ;
  assign n31595 = ~n31592 & ~n31594 ;
  assign n31596 = n31590 & n31595 ;
  assign n31597 = n31585 & n31596 ;
  assign n31598 = \m6_addr_i[0]_pad  & n14211 ;
  assign n31599 = n14204 & n31598 ;
  assign n31600 = \m5_addr_i[0]_pad  & ~n14211 ;
  assign n31601 = n14236 & n31600 ;
  assign n31602 = ~n31599 & ~n31601 ;
  assign n31603 = \m0_addr_i[0]_pad  & n14211 ;
  assign n31604 = n14219 & n31603 ;
  assign n31605 = \m4_addr_i[0]_pad  & n14211 ;
  assign n31606 = n14236 & n31605 ;
  assign n31607 = ~n31604 & ~n31606 ;
  assign n31608 = n31602 & n31607 ;
  assign n31609 = \m7_addr_i[0]_pad  & ~n14211 ;
  assign n31610 = n14204 & n31609 ;
  assign n31611 = \m3_addr_i[0]_pad  & ~n14211 ;
  assign n31612 = n14228 & n31611 ;
  assign n31613 = ~n31610 & ~n31612 ;
  assign n31614 = \m1_addr_i[0]_pad  & ~n14211 ;
  assign n31615 = n14219 & n31614 ;
  assign n31616 = \m2_addr_i[0]_pad  & n14211 ;
  assign n31617 = n14228 & n31616 ;
  assign n31618 = ~n31615 & ~n31617 ;
  assign n31619 = n31613 & n31618 ;
  assign n31620 = n31608 & n31619 ;
  assign n31621 = \m3_addr_i[10]_pad  & ~n14211 ;
  assign n31622 = n14228 & n31621 ;
  assign n31623 = \m4_addr_i[10]_pad  & n14211 ;
  assign n31624 = n14236 & n31623 ;
  assign n31625 = ~n31622 & ~n31624 ;
  assign n31626 = \m6_addr_i[10]_pad  & n14211 ;
  assign n31627 = n14204 & n31626 ;
  assign n31628 = \m2_addr_i[10]_pad  & n14211 ;
  assign n31629 = n14228 & n31628 ;
  assign n31630 = ~n31627 & ~n31629 ;
  assign n31631 = n31625 & n31630 ;
  assign n31632 = \m5_addr_i[10]_pad  & ~n14211 ;
  assign n31633 = n14236 & n31632 ;
  assign n31634 = \m1_addr_i[10]_pad  & ~n14211 ;
  assign n31635 = n14219 & n31634 ;
  assign n31636 = ~n31633 & ~n31635 ;
  assign n31637 = \m0_addr_i[10]_pad  & n14211 ;
  assign n31638 = n14219 & n31637 ;
  assign n31639 = \m7_addr_i[10]_pad  & ~n14211 ;
  assign n31640 = n14204 & n31639 ;
  assign n31641 = ~n31638 & ~n31640 ;
  assign n31642 = n31636 & n31641 ;
  assign n31643 = n31631 & n31642 ;
  assign n31644 = \m3_addr_i[11]_pad  & ~n14211 ;
  assign n31645 = n14228 & n31644 ;
  assign n31646 = \m4_addr_i[11]_pad  & n14211 ;
  assign n31647 = n14236 & n31646 ;
  assign n31648 = ~n31645 & ~n31647 ;
  assign n31649 = \m6_addr_i[11]_pad  & n14211 ;
  assign n31650 = n14204 & n31649 ;
  assign n31651 = \m2_addr_i[11]_pad  & n14211 ;
  assign n31652 = n14228 & n31651 ;
  assign n31653 = ~n31650 & ~n31652 ;
  assign n31654 = n31648 & n31653 ;
  assign n31655 = \m5_addr_i[11]_pad  & ~n14211 ;
  assign n31656 = n14236 & n31655 ;
  assign n31657 = \m1_addr_i[11]_pad  & ~n14211 ;
  assign n31658 = n14219 & n31657 ;
  assign n31659 = ~n31656 & ~n31658 ;
  assign n31660 = \m0_addr_i[11]_pad  & n14211 ;
  assign n31661 = n14219 & n31660 ;
  assign n31662 = \m7_addr_i[11]_pad  & ~n14211 ;
  assign n31663 = n14204 & n31662 ;
  assign n31664 = ~n31661 & ~n31663 ;
  assign n31665 = n31659 & n31664 ;
  assign n31666 = n31654 & n31665 ;
  assign n31667 = \m3_addr_i[12]_pad  & ~n14211 ;
  assign n31668 = n14228 & n31667 ;
  assign n31669 = \m4_addr_i[12]_pad  & n14211 ;
  assign n31670 = n14236 & n31669 ;
  assign n31671 = ~n31668 & ~n31670 ;
  assign n31672 = \m6_addr_i[12]_pad  & n14211 ;
  assign n31673 = n14204 & n31672 ;
  assign n31674 = \m2_addr_i[12]_pad  & n14211 ;
  assign n31675 = n14228 & n31674 ;
  assign n31676 = ~n31673 & ~n31675 ;
  assign n31677 = n31671 & n31676 ;
  assign n31678 = \m5_addr_i[12]_pad  & ~n14211 ;
  assign n31679 = n14236 & n31678 ;
  assign n31680 = \m1_addr_i[12]_pad  & ~n14211 ;
  assign n31681 = n14219 & n31680 ;
  assign n31682 = ~n31679 & ~n31681 ;
  assign n31683 = \m0_addr_i[12]_pad  & n14211 ;
  assign n31684 = n14219 & n31683 ;
  assign n31685 = \m7_addr_i[12]_pad  & ~n14211 ;
  assign n31686 = n14204 & n31685 ;
  assign n31687 = ~n31684 & ~n31686 ;
  assign n31688 = n31682 & n31687 ;
  assign n31689 = n31677 & n31688 ;
  assign n31690 = \m3_addr_i[13]_pad  & ~n14211 ;
  assign n31691 = n14228 & n31690 ;
  assign n31692 = \m4_addr_i[13]_pad  & n14211 ;
  assign n31693 = n14236 & n31692 ;
  assign n31694 = ~n31691 & ~n31693 ;
  assign n31695 = \m6_addr_i[13]_pad  & n14211 ;
  assign n31696 = n14204 & n31695 ;
  assign n31697 = \m2_addr_i[13]_pad  & n14211 ;
  assign n31698 = n14228 & n31697 ;
  assign n31699 = ~n31696 & ~n31698 ;
  assign n31700 = n31694 & n31699 ;
  assign n31701 = \m5_addr_i[13]_pad  & ~n14211 ;
  assign n31702 = n14236 & n31701 ;
  assign n31703 = \m1_addr_i[13]_pad  & ~n14211 ;
  assign n31704 = n14219 & n31703 ;
  assign n31705 = ~n31702 & ~n31704 ;
  assign n31706 = \m0_addr_i[13]_pad  & n14211 ;
  assign n31707 = n14219 & n31706 ;
  assign n31708 = \m7_addr_i[13]_pad  & ~n14211 ;
  assign n31709 = n14204 & n31708 ;
  assign n31710 = ~n31707 & ~n31709 ;
  assign n31711 = n31705 & n31710 ;
  assign n31712 = n31700 & n31711 ;
  assign n31713 = \m3_addr_i[14]_pad  & ~n14211 ;
  assign n31714 = n14228 & n31713 ;
  assign n31715 = \m4_addr_i[14]_pad  & n14211 ;
  assign n31716 = n14236 & n31715 ;
  assign n31717 = ~n31714 & ~n31716 ;
  assign n31718 = \m6_addr_i[14]_pad  & n14211 ;
  assign n31719 = n14204 & n31718 ;
  assign n31720 = \m2_addr_i[14]_pad  & n14211 ;
  assign n31721 = n14228 & n31720 ;
  assign n31722 = ~n31719 & ~n31721 ;
  assign n31723 = n31717 & n31722 ;
  assign n31724 = \m5_addr_i[14]_pad  & ~n14211 ;
  assign n31725 = n14236 & n31724 ;
  assign n31726 = \m1_addr_i[14]_pad  & ~n14211 ;
  assign n31727 = n14219 & n31726 ;
  assign n31728 = ~n31725 & ~n31727 ;
  assign n31729 = \m0_addr_i[14]_pad  & n14211 ;
  assign n31730 = n14219 & n31729 ;
  assign n31731 = \m7_addr_i[14]_pad  & ~n14211 ;
  assign n31732 = n14204 & n31731 ;
  assign n31733 = ~n31730 & ~n31732 ;
  assign n31734 = n31728 & n31733 ;
  assign n31735 = n31723 & n31734 ;
  assign n31736 = \m3_addr_i[15]_pad  & ~n14211 ;
  assign n31737 = n14228 & n31736 ;
  assign n31738 = \m4_addr_i[15]_pad  & n14211 ;
  assign n31739 = n14236 & n31738 ;
  assign n31740 = ~n31737 & ~n31739 ;
  assign n31741 = \m6_addr_i[15]_pad  & n14211 ;
  assign n31742 = n14204 & n31741 ;
  assign n31743 = \m2_addr_i[15]_pad  & n14211 ;
  assign n31744 = n14228 & n31743 ;
  assign n31745 = ~n31742 & ~n31744 ;
  assign n31746 = n31740 & n31745 ;
  assign n31747 = \m5_addr_i[15]_pad  & ~n14211 ;
  assign n31748 = n14236 & n31747 ;
  assign n31749 = \m1_addr_i[15]_pad  & ~n14211 ;
  assign n31750 = n14219 & n31749 ;
  assign n31751 = ~n31748 & ~n31750 ;
  assign n31752 = \m0_addr_i[15]_pad  & n14211 ;
  assign n31753 = n14219 & n31752 ;
  assign n31754 = \m7_addr_i[15]_pad  & ~n14211 ;
  assign n31755 = n14204 & n31754 ;
  assign n31756 = ~n31753 & ~n31755 ;
  assign n31757 = n31751 & n31756 ;
  assign n31758 = n31746 & n31757 ;
  assign n31759 = \m3_addr_i[16]_pad  & ~n14211 ;
  assign n31760 = n14228 & n31759 ;
  assign n31761 = \m4_addr_i[16]_pad  & n14211 ;
  assign n31762 = n14236 & n31761 ;
  assign n31763 = ~n31760 & ~n31762 ;
  assign n31764 = \m6_addr_i[16]_pad  & n14211 ;
  assign n31765 = n14204 & n31764 ;
  assign n31766 = \m2_addr_i[16]_pad  & n14211 ;
  assign n31767 = n14228 & n31766 ;
  assign n31768 = ~n31765 & ~n31767 ;
  assign n31769 = n31763 & n31768 ;
  assign n31770 = \m5_addr_i[16]_pad  & ~n14211 ;
  assign n31771 = n14236 & n31770 ;
  assign n31772 = \m1_addr_i[16]_pad  & ~n14211 ;
  assign n31773 = n14219 & n31772 ;
  assign n31774 = ~n31771 & ~n31773 ;
  assign n31775 = \m0_addr_i[16]_pad  & n14211 ;
  assign n31776 = n14219 & n31775 ;
  assign n31777 = \m7_addr_i[16]_pad  & ~n14211 ;
  assign n31778 = n14204 & n31777 ;
  assign n31779 = ~n31776 & ~n31778 ;
  assign n31780 = n31774 & n31779 ;
  assign n31781 = n31769 & n31780 ;
  assign n31782 = \m3_addr_i[17]_pad  & ~n14211 ;
  assign n31783 = n14228 & n31782 ;
  assign n31784 = \m4_addr_i[17]_pad  & n14211 ;
  assign n31785 = n14236 & n31784 ;
  assign n31786 = ~n31783 & ~n31785 ;
  assign n31787 = \m6_addr_i[17]_pad  & n14211 ;
  assign n31788 = n14204 & n31787 ;
  assign n31789 = \m2_addr_i[17]_pad  & n14211 ;
  assign n31790 = n14228 & n31789 ;
  assign n31791 = ~n31788 & ~n31790 ;
  assign n31792 = n31786 & n31791 ;
  assign n31793 = \m5_addr_i[17]_pad  & ~n14211 ;
  assign n31794 = n14236 & n31793 ;
  assign n31795 = \m1_addr_i[17]_pad  & ~n14211 ;
  assign n31796 = n14219 & n31795 ;
  assign n31797 = ~n31794 & ~n31796 ;
  assign n31798 = \m0_addr_i[17]_pad  & n14211 ;
  assign n31799 = n14219 & n31798 ;
  assign n31800 = \m7_addr_i[17]_pad  & ~n14211 ;
  assign n31801 = n14204 & n31800 ;
  assign n31802 = ~n31799 & ~n31801 ;
  assign n31803 = n31797 & n31802 ;
  assign n31804 = n31792 & n31803 ;
  assign n31805 = \m3_addr_i[18]_pad  & ~n14211 ;
  assign n31806 = n14228 & n31805 ;
  assign n31807 = \m4_addr_i[18]_pad  & n14211 ;
  assign n31808 = n14236 & n31807 ;
  assign n31809 = ~n31806 & ~n31808 ;
  assign n31810 = \m6_addr_i[18]_pad  & n14211 ;
  assign n31811 = n14204 & n31810 ;
  assign n31812 = \m2_addr_i[18]_pad  & n14211 ;
  assign n31813 = n14228 & n31812 ;
  assign n31814 = ~n31811 & ~n31813 ;
  assign n31815 = n31809 & n31814 ;
  assign n31816 = \m5_addr_i[18]_pad  & ~n14211 ;
  assign n31817 = n14236 & n31816 ;
  assign n31818 = \m1_addr_i[18]_pad  & ~n14211 ;
  assign n31819 = n14219 & n31818 ;
  assign n31820 = ~n31817 & ~n31819 ;
  assign n31821 = \m0_addr_i[18]_pad  & n14211 ;
  assign n31822 = n14219 & n31821 ;
  assign n31823 = \m7_addr_i[18]_pad  & ~n14211 ;
  assign n31824 = n14204 & n31823 ;
  assign n31825 = ~n31822 & ~n31824 ;
  assign n31826 = n31820 & n31825 ;
  assign n31827 = n31815 & n31826 ;
  assign n31828 = \m3_addr_i[19]_pad  & ~n14211 ;
  assign n31829 = n14228 & n31828 ;
  assign n31830 = \m4_addr_i[19]_pad  & n14211 ;
  assign n31831 = n14236 & n31830 ;
  assign n31832 = ~n31829 & ~n31831 ;
  assign n31833 = \m6_addr_i[19]_pad  & n14211 ;
  assign n31834 = n14204 & n31833 ;
  assign n31835 = \m2_addr_i[19]_pad  & n14211 ;
  assign n31836 = n14228 & n31835 ;
  assign n31837 = ~n31834 & ~n31836 ;
  assign n31838 = n31832 & n31837 ;
  assign n31839 = \m5_addr_i[19]_pad  & ~n14211 ;
  assign n31840 = n14236 & n31839 ;
  assign n31841 = \m1_addr_i[19]_pad  & ~n14211 ;
  assign n31842 = n14219 & n31841 ;
  assign n31843 = ~n31840 & ~n31842 ;
  assign n31844 = \m0_addr_i[19]_pad  & n14211 ;
  assign n31845 = n14219 & n31844 ;
  assign n31846 = \m7_addr_i[19]_pad  & ~n14211 ;
  assign n31847 = n14204 & n31846 ;
  assign n31848 = ~n31845 & ~n31847 ;
  assign n31849 = n31843 & n31848 ;
  assign n31850 = n31838 & n31849 ;
  assign n31851 = \m3_addr_i[1]_pad  & ~n14211 ;
  assign n31852 = n14228 & n31851 ;
  assign n31853 = \m4_addr_i[1]_pad  & n14211 ;
  assign n31854 = n14236 & n31853 ;
  assign n31855 = ~n31852 & ~n31854 ;
  assign n31856 = \m6_addr_i[1]_pad  & n14211 ;
  assign n31857 = n14204 & n31856 ;
  assign n31858 = \m2_addr_i[1]_pad  & n14211 ;
  assign n31859 = n14228 & n31858 ;
  assign n31860 = ~n31857 & ~n31859 ;
  assign n31861 = n31855 & n31860 ;
  assign n31862 = \m5_addr_i[1]_pad  & ~n14211 ;
  assign n31863 = n14236 & n31862 ;
  assign n31864 = \m1_addr_i[1]_pad  & ~n14211 ;
  assign n31865 = n14219 & n31864 ;
  assign n31866 = ~n31863 & ~n31865 ;
  assign n31867 = \m0_addr_i[1]_pad  & n14211 ;
  assign n31868 = n14219 & n31867 ;
  assign n31869 = \m7_addr_i[1]_pad  & ~n14211 ;
  assign n31870 = n14204 & n31869 ;
  assign n31871 = ~n31868 & ~n31870 ;
  assign n31872 = n31866 & n31871 ;
  assign n31873 = n31861 & n31872 ;
  assign n31874 = \m3_addr_i[20]_pad  & ~n14211 ;
  assign n31875 = n14228 & n31874 ;
  assign n31876 = \m4_addr_i[20]_pad  & n14211 ;
  assign n31877 = n14236 & n31876 ;
  assign n31878 = ~n31875 & ~n31877 ;
  assign n31879 = \m6_addr_i[20]_pad  & n14211 ;
  assign n31880 = n14204 & n31879 ;
  assign n31881 = \m2_addr_i[20]_pad  & n14211 ;
  assign n31882 = n14228 & n31881 ;
  assign n31883 = ~n31880 & ~n31882 ;
  assign n31884 = n31878 & n31883 ;
  assign n31885 = \m5_addr_i[20]_pad  & ~n14211 ;
  assign n31886 = n14236 & n31885 ;
  assign n31887 = \m1_addr_i[20]_pad  & ~n14211 ;
  assign n31888 = n14219 & n31887 ;
  assign n31889 = ~n31886 & ~n31888 ;
  assign n31890 = \m0_addr_i[20]_pad  & n14211 ;
  assign n31891 = n14219 & n31890 ;
  assign n31892 = \m7_addr_i[20]_pad  & ~n14211 ;
  assign n31893 = n14204 & n31892 ;
  assign n31894 = ~n31891 & ~n31893 ;
  assign n31895 = n31889 & n31894 ;
  assign n31896 = n31884 & n31895 ;
  assign n31897 = \m3_addr_i[21]_pad  & ~n14211 ;
  assign n31898 = n14228 & n31897 ;
  assign n31899 = \m4_addr_i[21]_pad  & n14211 ;
  assign n31900 = n14236 & n31899 ;
  assign n31901 = ~n31898 & ~n31900 ;
  assign n31902 = \m6_addr_i[21]_pad  & n14211 ;
  assign n31903 = n14204 & n31902 ;
  assign n31904 = \m2_addr_i[21]_pad  & n14211 ;
  assign n31905 = n14228 & n31904 ;
  assign n31906 = ~n31903 & ~n31905 ;
  assign n31907 = n31901 & n31906 ;
  assign n31908 = \m5_addr_i[21]_pad  & ~n14211 ;
  assign n31909 = n14236 & n31908 ;
  assign n31910 = \m1_addr_i[21]_pad  & ~n14211 ;
  assign n31911 = n14219 & n31910 ;
  assign n31912 = ~n31909 & ~n31911 ;
  assign n31913 = \m0_addr_i[21]_pad  & n14211 ;
  assign n31914 = n14219 & n31913 ;
  assign n31915 = \m7_addr_i[21]_pad  & ~n14211 ;
  assign n31916 = n14204 & n31915 ;
  assign n31917 = ~n31914 & ~n31916 ;
  assign n31918 = n31912 & n31917 ;
  assign n31919 = n31907 & n31918 ;
  assign n31920 = \m3_addr_i[22]_pad  & ~n14211 ;
  assign n31921 = n14228 & n31920 ;
  assign n31922 = \m4_addr_i[22]_pad  & n14211 ;
  assign n31923 = n14236 & n31922 ;
  assign n31924 = ~n31921 & ~n31923 ;
  assign n31925 = \m6_addr_i[22]_pad  & n14211 ;
  assign n31926 = n14204 & n31925 ;
  assign n31927 = \m2_addr_i[22]_pad  & n14211 ;
  assign n31928 = n14228 & n31927 ;
  assign n31929 = ~n31926 & ~n31928 ;
  assign n31930 = n31924 & n31929 ;
  assign n31931 = \m5_addr_i[22]_pad  & ~n14211 ;
  assign n31932 = n14236 & n31931 ;
  assign n31933 = \m1_addr_i[22]_pad  & ~n14211 ;
  assign n31934 = n14219 & n31933 ;
  assign n31935 = ~n31932 & ~n31934 ;
  assign n31936 = \m0_addr_i[22]_pad  & n14211 ;
  assign n31937 = n14219 & n31936 ;
  assign n31938 = \m7_addr_i[22]_pad  & ~n14211 ;
  assign n31939 = n14204 & n31938 ;
  assign n31940 = ~n31937 & ~n31939 ;
  assign n31941 = n31935 & n31940 ;
  assign n31942 = n31930 & n31941 ;
  assign n31943 = \m3_addr_i[23]_pad  & ~n14211 ;
  assign n31944 = n14228 & n31943 ;
  assign n31945 = \m4_addr_i[23]_pad  & n14211 ;
  assign n31946 = n14236 & n31945 ;
  assign n31947 = ~n31944 & ~n31946 ;
  assign n31948 = \m6_addr_i[23]_pad  & n14211 ;
  assign n31949 = n14204 & n31948 ;
  assign n31950 = \m2_addr_i[23]_pad  & n14211 ;
  assign n31951 = n14228 & n31950 ;
  assign n31952 = ~n31949 & ~n31951 ;
  assign n31953 = n31947 & n31952 ;
  assign n31954 = \m5_addr_i[23]_pad  & ~n14211 ;
  assign n31955 = n14236 & n31954 ;
  assign n31956 = \m1_addr_i[23]_pad  & ~n14211 ;
  assign n31957 = n14219 & n31956 ;
  assign n31958 = ~n31955 & ~n31957 ;
  assign n31959 = \m0_addr_i[23]_pad  & n14211 ;
  assign n31960 = n14219 & n31959 ;
  assign n31961 = \m7_addr_i[23]_pad  & ~n14211 ;
  assign n31962 = n14204 & n31961 ;
  assign n31963 = ~n31960 & ~n31962 ;
  assign n31964 = n31958 & n31963 ;
  assign n31965 = n31953 & n31964 ;
  assign n31966 = \m3_addr_i[24]_pad  & ~n14211 ;
  assign n31967 = n14228 & n31966 ;
  assign n31968 = \m4_addr_i[24]_pad  & n14211 ;
  assign n31969 = n14236 & n31968 ;
  assign n31970 = ~n31967 & ~n31969 ;
  assign n31971 = \m5_addr_i[24]_pad  & ~n14211 ;
  assign n31972 = n14236 & n31971 ;
  assign n31973 = \m2_addr_i[24]_pad  & n14211 ;
  assign n31974 = n14228 & n31973 ;
  assign n31975 = ~n31972 & ~n31974 ;
  assign n31976 = n31970 & n31975 ;
  assign n31977 = \m6_addr_i[24]_pad  & n14211 ;
  assign n31978 = n14204 & n31977 ;
  assign n31979 = \m1_addr_i[24]_pad  & ~n14211 ;
  assign n31980 = n14219 & n31979 ;
  assign n31981 = ~n31978 & ~n31980 ;
  assign n31982 = \m0_addr_i[24]_pad  & n14211 ;
  assign n31983 = n14219 & n31982 ;
  assign n31984 = \m7_addr_i[24]_pad  & ~n14211 ;
  assign n31985 = n14204 & n31984 ;
  assign n31986 = ~n31983 & ~n31985 ;
  assign n31987 = n31981 & n31986 ;
  assign n31988 = n31976 & n31987 ;
  assign n31989 = \m3_addr_i[25]_pad  & ~n14211 ;
  assign n31990 = n14228 & n31989 ;
  assign n31991 = \m4_addr_i[25]_pad  & n14211 ;
  assign n31992 = n14236 & n31991 ;
  assign n31993 = ~n31990 & ~n31992 ;
  assign n31994 = \m5_addr_i[25]_pad  & ~n14211 ;
  assign n31995 = n14236 & n31994 ;
  assign n31996 = \m2_addr_i[25]_pad  & n14211 ;
  assign n31997 = n14228 & n31996 ;
  assign n31998 = ~n31995 & ~n31997 ;
  assign n31999 = n31993 & n31998 ;
  assign n32000 = \m6_addr_i[25]_pad  & n14211 ;
  assign n32001 = n14204 & n32000 ;
  assign n32002 = \m1_addr_i[25]_pad  & ~n14211 ;
  assign n32003 = n14219 & n32002 ;
  assign n32004 = ~n32001 & ~n32003 ;
  assign n32005 = \m0_addr_i[25]_pad  & n14211 ;
  assign n32006 = n14219 & n32005 ;
  assign n32007 = \m7_addr_i[25]_pad  & ~n14211 ;
  assign n32008 = n14204 & n32007 ;
  assign n32009 = ~n32006 & ~n32008 ;
  assign n32010 = n32004 & n32009 ;
  assign n32011 = n31999 & n32010 ;
  assign n32012 = \m3_addr_i[26]_pad  & ~n14211 ;
  assign n32013 = n14228 & n32012 ;
  assign n32014 = \m4_addr_i[26]_pad  & n14211 ;
  assign n32015 = n14236 & n32014 ;
  assign n32016 = ~n32013 & ~n32015 ;
  assign n32017 = \m5_addr_i[26]_pad  & ~n14211 ;
  assign n32018 = n14236 & n32017 ;
  assign n32019 = \m2_addr_i[26]_pad  & n14211 ;
  assign n32020 = n14228 & n32019 ;
  assign n32021 = ~n32018 & ~n32020 ;
  assign n32022 = n32016 & n32021 ;
  assign n32023 = \m6_addr_i[26]_pad  & n14211 ;
  assign n32024 = n14204 & n32023 ;
  assign n32025 = \m1_addr_i[26]_pad  & ~n14211 ;
  assign n32026 = n14219 & n32025 ;
  assign n32027 = ~n32024 & ~n32026 ;
  assign n32028 = \m0_addr_i[26]_pad  & n14211 ;
  assign n32029 = n14219 & n32028 ;
  assign n32030 = \m7_addr_i[26]_pad  & ~n14211 ;
  assign n32031 = n14204 & n32030 ;
  assign n32032 = ~n32029 & ~n32031 ;
  assign n32033 = n32027 & n32032 ;
  assign n32034 = n32022 & n32033 ;
  assign n32035 = \m3_addr_i[27]_pad  & ~n14211 ;
  assign n32036 = n14228 & n32035 ;
  assign n32037 = \m4_addr_i[27]_pad  & n14211 ;
  assign n32038 = n14236 & n32037 ;
  assign n32039 = ~n32036 & ~n32038 ;
  assign n32040 = \m5_addr_i[27]_pad  & ~n14211 ;
  assign n32041 = n14236 & n32040 ;
  assign n32042 = \m2_addr_i[27]_pad  & n14211 ;
  assign n32043 = n14228 & n32042 ;
  assign n32044 = ~n32041 & ~n32043 ;
  assign n32045 = n32039 & n32044 ;
  assign n32046 = \m6_addr_i[27]_pad  & n14211 ;
  assign n32047 = n14204 & n32046 ;
  assign n32048 = \m1_addr_i[27]_pad  & ~n14211 ;
  assign n32049 = n14219 & n32048 ;
  assign n32050 = ~n32047 & ~n32049 ;
  assign n32051 = \m0_addr_i[27]_pad  & n14211 ;
  assign n32052 = n14219 & n32051 ;
  assign n32053 = \m7_addr_i[27]_pad  & ~n14211 ;
  assign n32054 = n14204 & n32053 ;
  assign n32055 = ~n32052 & ~n32054 ;
  assign n32056 = n32050 & n32055 ;
  assign n32057 = n32045 & n32056 ;
  assign n32058 = \m3_addr_i[28]_pad  & ~n14211 ;
  assign n32059 = n14228 & n32058 ;
  assign n32060 = \m4_addr_i[28]_pad  & n14211 ;
  assign n32061 = n14236 & n32060 ;
  assign n32062 = ~n32059 & ~n32061 ;
  assign n32063 = \m5_addr_i[28]_pad  & ~n14211 ;
  assign n32064 = n14236 & n32063 ;
  assign n32065 = \m2_addr_i[28]_pad  & n14211 ;
  assign n32066 = n14228 & n32065 ;
  assign n32067 = ~n32064 & ~n32066 ;
  assign n32068 = n32062 & n32067 ;
  assign n32069 = \m6_addr_i[28]_pad  & n14211 ;
  assign n32070 = n14204 & n32069 ;
  assign n32071 = \m1_addr_i[28]_pad  & ~n14211 ;
  assign n32072 = n14219 & n32071 ;
  assign n32073 = ~n32070 & ~n32072 ;
  assign n32074 = \m0_addr_i[28]_pad  & n14211 ;
  assign n32075 = n14219 & n32074 ;
  assign n32076 = \m7_addr_i[28]_pad  & ~n14211 ;
  assign n32077 = n14204 & n32076 ;
  assign n32078 = ~n32075 & ~n32077 ;
  assign n32079 = n32073 & n32078 ;
  assign n32080 = n32068 & n32079 ;
  assign n32081 = \m0_addr_i[29]_pad  & n14211 ;
  assign n32082 = n14219 & n32081 ;
  assign n32083 = \m7_addr_i[29]_pad  & ~n14211 ;
  assign n32084 = n14204 & n32083 ;
  assign n32085 = ~n32082 & ~n32084 ;
  assign n32086 = \m1_addr_i[29]_pad  & ~n14211 ;
  assign n32087 = n14219 & n32086 ;
  assign n32088 = \m4_addr_i[29]_pad  & n14211 ;
  assign n32089 = n14236 & n32088 ;
  assign n32090 = ~n32087 & ~n32089 ;
  assign n32091 = n32085 & n32090 ;
  assign n32092 = \m2_addr_i[29]_pad  & n14211 ;
  assign n32093 = n14228 & n32092 ;
  assign n32094 = \m3_addr_i[29]_pad  & ~n14211 ;
  assign n32095 = n14228 & n32094 ;
  assign n32096 = ~n32093 & ~n32095 ;
  assign n32097 = \m5_addr_i[29]_pad  & ~n14211 ;
  assign n32098 = n14236 & n32097 ;
  assign n32099 = \m6_addr_i[29]_pad  & n14211 ;
  assign n32100 = n14204 & n32099 ;
  assign n32101 = ~n32098 & ~n32100 ;
  assign n32102 = n32096 & n32101 ;
  assign n32103 = n32091 & n32102 ;
  assign n32104 = \m3_addr_i[2]_pad  & ~n14211 ;
  assign n32105 = n14228 & n32104 ;
  assign n32106 = \m4_addr_i[2]_pad  & n14211 ;
  assign n32107 = n14236 & n32106 ;
  assign n32108 = ~n32105 & ~n32107 ;
  assign n32109 = \m6_addr_i[2]_pad  & n14211 ;
  assign n32110 = n14204 & n32109 ;
  assign n32111 = \m2_addr_i[2]_pad  & n14211 ;
  assign n32112 = n14228 & n32111 ;
  assign n32113 = ~n32110 & ~n32112 ;
  assign n32114 = n32108 & n32113 ;
  assign n32115 = \m5_addr_i[2]_pad  & ~n14211 ;
  assign n32116 = n14236 & n32115 ;
  assign n32117 = \m1_addr_i[2]_pad  & ~n14211 ;
  assign n32118 = n14219 & n32117 ;
  assign n32119 = ~n32116 & ~n32118 ;
  assign n32120 = \m0_addr_i[2]_pad  & n14211 ;
  assign n32121 = n14219 & n32120 ;
  assign n32122 = \m7_addr_i[2]_pad  & ~n14211 ;
  assign n32123 = n14204 & n32122 ;
  assign n32124 = ~n32121 & ~n32123 ;
  assign n32125 = n32119 & n32124 ;
  assign n32126 = n32114 & n32125 ;
  assign n32127 = \m5_addr_i[30]_pad  & ~n14211 ;
  assign n32128 = n14236 & n32127 ;
  assign n32129 = \m6_addr_i[30]_pad  & n14211 ;
  assign n32130 = n14204 & n32129 ;
  assign n32131 = ~n32128 & ~n32130 ;
  assign n32132 = \m0_addr_i[30]_pad  & n14211 ;
  assign n32133 = n14219 & n32132 ;
  assign n32134 = \m4_addr_i[30]_pad  & n14211 ;
  assign n32135 = n14236 & n32134 ;
  assign n32136 = ~n32133 & ~n32135 ;
  assign n32137 = n32131 & n32136 ;
  assign n32138 = \m7_addr_i[30]_pad  & ~n14211 ;
  assign n32139 = n14204 & n32138 ;
  assign n32140 = \m3_addr_i[30]_pad  & ~n14211 ;
  assign n32141 = n14228 & n32140 ;
  assign n32142 = ~n32139 & ~n32141 ;
  assign n32143 = \m1_addr_i[30]_pad  & ~n14211 ;
  assign n32144 = n14219 & n32143 ;
  assign n32145 = \m2_addr_i[30]_pad  & n14211 ;
  assign n32146 = n14228 & n32145 ;
  assign n32147 = ~n32144 & ~n32146 ;
  assign n32148 = n32142 & n32147 ;
  assign n32149 = n32137 & n32148 ;
  assign n32150 = \m5_addr_i[31]_pad  & ~n14211 ;
  assign n32151 = n14236 & n32150 ;
  assign n32152 = \m6_addr_i[31]_pad  & n14211 ;
  assign n32153 = n14204 & n32152 ;
  assign n32154 = ~n32151 & ~n32153 ;
  assign n32155 = \m3_addr_i[31]_pad  & ~n14211 ;
  assign n32156 = n14228 & n32155 ;
  assign n32157 = \m7_addr_i[31]_pad  & ~n14211 ;
  assign n32158 = n14204 & n32157 ;
  assign n32159 = ~n32156 & ~n32158 ;
  assign n32160 = n32154 & n32159 ;
  assign n32161 = \m4_addr_i[31]_pad  & n14211 ;
  assign n32162 = n14236 & n32161 ;
  assign n32163 = \m0_addr_i[31]_pad  & n14211 ;
  assign n32164 = n14219 & n32163 ;
  assign n32165 = ~n32162 & ~n32164 ;
  assign n32166 = \m1_addr_i[31]_pad  & ~n14211 ;
  assign n32167 = n14219 & n32166 ;
  assign n32168 = \m2_addr_i[31]_pad  & n14211 ;
  assign n32169 = n14228 & n32168 ;
  assign n32170 = ~n32167 & ~n32169 ;
  assign n32171 = n32165 & n32170 ;
  assign n32172 = n32160 & n32171 ;
  assign n32173 = \m3_addr_i[3]_pad  & ~n14211 ;
  assign n32174 = n14228 & n32173 ;
  assign n32175 = \m4_addr_i[3]_pad  & n14211 ;
  assign n32176 = n14236 & n32175 ;
  assign n32177 = ~n32174 & ~n32176 ;
  assign n32178 = \m6_addr_i[3]_pad  & n14211 ;
  assign n32179 = n14204 & n32178 ;
  assign n32180 = \m2_addr_i[3]_pad  & n14211 ;
  assign n32181 = n14228 & n32180 ;
  assign n32182 = ~n32179 & ~n32181 ;
  assign n32183 = n32177 & n32182 ;
  assign n32184 = \m5_addr_i[3]_pad  & ~n14211 ;
  assign n32185 = n14236 & n32184 ;
  assign n32186 = \m1_addr_i[3]_pad  & ~n14211 ;
  assign n32187 = n14219 & n32186 ;
  assign n32188 = ~n32185 & ~n32187 ;
  assign n32189 = \m0_addr_i[3]_pad  & n14211 ;
  assign n32190 = n14219 & n32189 ;
  assign n32191 = \m7_addr_i[3]_pad  & ~n14211 ;
  assign n32192 = n14204 & n32191 ;
  assign n32193 = ~n32190 & ~n32192 ;
  assign n32194 = n32188 & n32193 ;
  assign n32195 = n32183 & n32194 ;
  assign n32196 = \m3_addr_i[4]_pad  & ~n14211 ;
  assign n32197 = n14228 & n32196 ;
  assign n32198 = \m4_addr_i[4]_pad  & n14211 ;
  assign n32199 = n14236 & n32198 ;
  assign n32200 = ~n32197 & ~n32199 ;
  assign n32201 = \m6_addr_i[4]_pad  & n14211 ;
  assign n32202 = n14204 & n32201 ;
  assign n32203 = \m2_addr_i[4]_pad  & n14211 ;
  assign n32204 = n14228 & n32203 ;
  assign n32205 = ~n32202 & ~n32204 ;
  assign n32206 = n32200 & n32205 ;
  assign n32207 = \m5_addr_i[4]_pad  & ~n14211 ;
  assign n32208 = n14236 & n32207 ;
  assign n32209 = \m1_addr_i[4]_pad  & ~n14211 ;
  assign n32210 = n14219 & n32209 ;
  assign n32211 = ~n32208 & ~n32210 ;
  assign n32212 = \m0_addr_i[4]_pad  & n14211 ;
  assign n32213 = n14219 & n32212 ;
  assign n32214 = \m7_addr_i[4]_pad  & ~n14211 ;
  assign n32215 = n14204 & n32214 ;
  assign n32216 = ~n32213 & ~n32215 ;
  assign n32217 = n32211 & n32216 ;
  assign n32218 = n32206 & n32217 ;
  assign n32219 = \m3_addr_i[5]_pad  & ~n14211 ;
  assign n32220 = n14228 & n32219 ;
  assign n32221 = \m4_addr_i[5]_pad  & n14211 ;
  assign n32222 = n14236 & n32221 ;
  assign n32223 = ~n32220 & ~n32222 ;
  assign n32224 = \m6_addr_i[5]_pad  & n14211 ;
  assign n32225 = n14204 & n32224 ;
  assign n32226 = \m2_addr_i[5]_pad  & n14211 ;
  assign n32227 = n14228 & n32226 ;
  assign n32228 = ~n32225 & ~n32227 ;
  assign n32229 = n32223 & n32228 ;
  assign n32230 = \m5_addr_i[5]_pad  & ~n14211 ;
  assign n32231 = n14236 & n32230 ;
  assign n32232 = \m1_addr_i[5]_pad  & ~n14211 ;
  assign n32233 = n14219 & n32232 ;
  assign n32234 = ~n32231 & ~n32233 ;
  assign n32235 = \m0_addr_i[5]_pad  & n14211 ;
  assign n32236 = n14219 & n32235 ;
  assign n32237 = \m7_addr_i[5]_pad  & ~n14211 ;
  assign n32238 = n14204 & n32237 ;
  assign n32239 = ~n32236 & ~n32238 ;
  assign n32240 = n32234 & n32239 ;
  assign n32241 = n32229 & n32240 ;
  assign n32242 = \m1_addr_i[6]_pad  & ~n14211 ;
  assign n32243 = n14219 & n32242 ;
  assign n32244 = \m2_addr_i[6]_pad  & n14211 ;
  assign n32245 = n14228 & n32244 ;
  assign n32246 = ~n32243 & ~n32245 ;
  assign n32247 = \m6_addr_i[6]_pad  & n14211 ;
  assign n32248 = n14204 & n32247 ;
  assign n32249 = \m4_addr_i[6]_pad  & n14211 ;
  assign n32250 = n14236 & n32249 ;
  assign n32251 = ~n32248 & ~n32250 ;
  assign n32252 = n32246 & n32251 ;
  assign n32253 = \m5_addr_i[6]_pad  & ~n14211 ;
  assign n32254 = n14236 & n32253 ;
  assign n32255 = \m3_addr_i[6]_pad  & ~n14211 ;
  assign n32256 = n14228 & n32255 ;
  assign n32257 = ~n32254 & ~n32256 ;
  assign n32258 = \m0_addr_i[6]_pad  & n14211 ;
  assign n32259 = n14219 & n32258 ;
  assign n32260 = \m7_addr_i[6]_pad  & ~n14211 ;
  assign n32261 = n14204 & n32260 ;
  assign n32262 = ~n32259 & ~n32261 ;
  assign n32263 = n32257 & n32262 ;
  assign n32264 = n32252 & n32263 ;
  assign n32265 = \m6_addr_i[7]_pad  & n14211 ;
  assign n32266 = n14204 & n32265 ;
  assign n32267 = \m5_addr_i[7]_pad  & ~n14211 ;
  assign n32268 = n14236 & n32267 ;
  assign n32269 = ~n32266 & ~n32268 ;
  assign n32270 = \m3_addr_i[7]_pad  & ~n14211 ;
  assign n32271 = n14228 & n32270 ;
  assign n32272 = \m2_addr_i[7]_pad  & n14211 ;
  assign n32273 = n14228 & n32272 ;
  assign n32274 = ~n32271 & ~n32273 ;
  assign n32275 = n32269 & n32274 ;
  assign n32276 = \m4_addr_i[7]_pad  & n14211 ;
  assign n32277 = n14236 & n32276 ;
  assign n32278 = \m1_addr_i[7]_pad  & ~n14211 ;
  assign n32279 = n14219 & n32278 ;
  assign n32280 = ~n32277 & ~n32279 ;
  assign n32281 = \m0_addr_i[7]_pad  & n14211 ;
  assign n32282 = n14219 & n32281 ;
  assign n32283 = \m7_addr_i[7]_pad  & ~n14211 ;
  assign n32284 = n14204 & n32283 ;
  assign n32285 = ~n32282 & ~n32284 ;
  assign n32286 = n32280 & n32285 ;
  assign n32287 = n32275 & n32286 ;
  assign n32288 = \m6_addr_i[8]_pad  & n14211 ;
  assign n32289 = n14204 & n32288 ;
  assign n32290 = \m5_addr_i[8]_pad  & ~n14211 ;
  assign n32291 = n14236 & n32290 ;
  assign n32292 = ~n32289 & ~n32291 ;
  assign n32293 = \m0_addr_i[8]_pad  & n14211 ;
  assign n32294 = n14219 & n32293 ;
  assign n32295 = \m4_addr_i[8]_pad  & n14211 ;
  assign n32296 = n14236 & n32295 ;
  assign n32297 = ~n32294 & ~n32296 ;
  assign n32298 = n32292 & n32297 ;
  assign n32299 = \m7_addr_i[8]_pad  & ~n14211 ;
  assign n32300 = n14204 & n32299 ;
  assign n32301 = \m3_addr_i[8]_pad  & ~n14211 ;
  assign n32302 = n14228 & n32301 ;
  assign n32303 = ~n32300 & ~n32302 ;
  assign n32304 = \m1_addr_i[8]_pad  & ~n14211 ;
  assign n32305 = n14219 & n32304 ;
  assign n32306 = \m2_addr_i[8]_pad  & n14211 ;
  assign n32307 = n14228 & n32306 ;
  assign n32308 = ~n32305 & ~n32307 ;
  assign n32309 = n32303 & n32308 ;
  assign n32310 = n32298 & n32309 ;
  assign n32311 = \m3_addr_i[9]_pad  & ~n14211 ;
  assign n32312 = n14228 & n32311 ;
  assign n32313 = \m4_addr_i[9]_pad  & n14211 ;
  assign n32314 = n14236 & n32313 ;
  assign n32315 = ~n32312 & ~n32314 ;
  assign n32316 = \m6_addr_i[9]_pad  & n14211 ;
  assign n32317 = n14204 & n32316 ;
  assign n32318 = \m2_addr_i[9]_pad  & n14211 ;
  assign n32319 = n14228 & n32318 ;
  assign n32320 = ~n32317 & ~n32319 ;
  assign n32321 = n32315 & n32320 ;
  assign n32322 = \m5_addr_i[9]_pad  & ~n14211 ;
  assign n32323 = n14236 & n32322 ;
  assign n32324 = \m1_addr_i[9]_pad  & ~n14211 ;
  assign n32325 = n14219 & n32324 ;
  assign n32326 = ~n32323 & ~n32325 ;
  assign n32327 = \m0_addr_i[9]_pad  & n14211 ;
  assign n32328 = n14219 & n32327 ;
  assign n32329 = \m7_addr_i[9]_pad  & ~n14211 ;
  assign n32330 = n14204 & n32329 ;
  assign n32331 = ~n32328 & ~n32330 ;
  assign n32332 = n32326 & n32331 ;
  assign n32333 = n32321 & n32332 ;
  assign n32334 = \m6_data_i[0]_pad  & n14211 ;
  assign n32335 = n14204 & n32334 ;
  assign n32336 = \m5_data_i[0]_pad  & ~n14211 ;
  assign n32337 = n14236 & n32336 ;
  assign n32338 = ~n32335 & ~n32337 ;
  assign n32339 = \m3_data_i[0]_pad  & ~n14211 ;
  assign n32340 = n14228 & n32339 ;
  assign n32341 = \m2_data_i[0]_pad  & n14211 ;
  assign n32342 = n14228 & n32341 ;
  assign n32343 = ~n32340 & ~n32342 ;
  assign n32344 = n32338 & n32343 ;
  assign n32345 = \m4_data_i[0]_pad  & n14211 ;
  assign n32346 = n14236 & n32345 ;
  assign n32347 = \m1_data_i[0]_pad  & ~n14211 ;
  assign n32348 = n14219 & n32347 ;
  assign n32349 = ~n32346 & ~n32348 ;
  assign n32350 = \m0_data_i[0]_pad  & n14211 ;
  assign n32351 = n14219 & n32350 ;
  assign n32352 = \m7_data_i[0]_pad  & ~n14211 ;
  assign n32353 = n14204 & n32352 ;
  assign n32354 = ~n32351 & ~n32353 ;
  assign n32355 = n32349 & n32354 ;
  assign n32356 = n32344 & n32355 ;
  assign n32357 = \m0_data_i[10]_pad  & n14211 ;
  assign n32358 = n14219 & n32357 ;
  assign n32359 = \m7_data_i[10]_pad  & ~n14211 ;
  assign n32360 = n14204 & n32359 ;
  assign n32361 = ~n32358 & ~n32360 ;
  assign n32362 = \m6_data_i[10]_pad  & n14211 ;
  assign n32363 = n14204 & n32362 ;
  assign n32364 = \m2_data_i[10]_pad  & n14211 ;
  assign n32365 = n14228 & n32364 ;
  assign n32366 = ~n32363 & ~n32365 ;
  assign n32367 = n32361 & n32366 ;
  assign n32368 = \m5_data_i[10]_pad  & ~n14211 ;
  assign n32369 = n14236 & n32368 ;
  assign n32370 = \m1_data_i[10]_pad  & ~n14211 ;
  assign n32371 = n14219 & n32370 ;
  assign n32372 = ~n32369 & ~n32371 ;
  assign n32373 = \m3_data_i[10]_pad  & ~n14211 ;
  assign n32374 = n14228 & n32373 ;
  assign n32375 = \m4_data_i[10]_pad  & n14211 ;
  assign n32376 = n14236 & n32375 ;
  assign n32377 = ~n32374 & ~n32376 ;
  assign n32378 = n32372 & n32377 ;
  assign n32379 = n32367 & n32378 ;
  assign n32380 = \m0_data_i[11]_pad  & n14211 ;
  assign n32381 = n14219 & n32380 ;
  assign n32382 = \m7_data_i[11]_pad  & ~n14211 ;
  assign n32383 = n14204 & n32382 ;
  assign n32384 = ~n32381 & ~n32383 ;
  assign n32385 = \m1_data_i[11]_pad  & ~n14211 ;
  assign n32386 = n14219 & n32385 ;
  assign n32387 = \m4_data_i[11]_pad  & n14211 ;
  assign n32388 = n14236 & n32387 ;
  assign n32389 = ~n32386 & ~n32388 ;
  assign n32390 = n32384 & n32389 ;
  assign n32391 = \m2_data_i[11]_pad  & n14211 ;
  assign n32392 = n14228 & n32391 ;
  assign n32393 = \m3_data_i[11]_pad  & ~n14211 ;
  assign n32394 = n14228 & n32393 ;
  assign n32395 = ~n32392 & ~n32394 ;
  assign n32396 = \m6_data_i[11]_pad  & n14211 ;
  assign n32397 = n14204 & n32396 ;
  assign n32398 = \m5_data_i[11]_pad  & ~n14211 ;
  assign n32399 = n14236 & n32398 ;
  assign n32400 = ~n32397 & ~n32399 ;
  assign n32401 = n32395 & n32400 ;
  assign n32402 = n32390 & n32401 ;
  assign n32403 = \m3_data_i[12]_pad  & ~n14211 ;
  assign n32404 = n14228 & n32403 ;
  assign n32405 = \m4_data_i[12]_pad  & n14211 ;
  assign n32406 = n14236 & n32405 ;
  assign n32407 = ~n32404 & ~n32406 ;
  assign n32408 = \m0_data_i[12]_pad  & n14211 ;
  assign n32409 = n14219 & n32408 ;
  assign n32410 = \m5_data_i[12]_pad  & ~n14211 ;
  assign n32411 = n14236 & n32410 ;
  assign n32412 = ~n32409 & ~n32411 ;
  assign n32413 = n32407 & n32412 ;
  assign n32414 = \m7_data_i[12]_pad  & ~n14211 ;
  assign n32415 = n14204 & n32414 ;
  assign n32416 = \m6_data_i[12]_pad  & n14211 ;
  assign n32417 = n14204 & n32416 ;
  assign n32418 = ~n32415 & ~n32417 ;
  assign n32419 = \m1_data_i[12]_pad  & ~n14211 ;
  assign n32420 = n14219 & n32419 ;
  assign n32421 = \m2_data_i[12]_pad  & n14211 ;
  assign n32422 = n14228 & n32421 ;
  assign n32423 = ~n32420 & ~n32422 ;
  assign n32424 = n32418 & n32423 ;
  assign n32425 = n32413 & n32424 ;
  assign n32426 = \m3_data_i[13]_pad  & ~n14211 ;
  assign n32427 = n14228 & n32426 ;
  assign n32428 = \m4_data_i[13]_pad  & n14211 ;
  assign n32429 = n14236 & n32428 ;
  assign n32430 = ~n32427 & ~n32429 ;
  assign n32431 = \m0_data_i[13]_pad  & n14211 ;
  assign n32432 = n14219 & n32431 ;
  assign n32433 = \m2_data_i[13]_pad  & n14211 ;
  assign n32434 = n14228 & n32433 ;
  assign n32435 = ~n32432 & ~n32434 ;
  assign n32436 = n32430 & n32435 ;
  assign n32437 = \m7_data_i[13]_pad  & ~n14211 ;
  assign n32438 = n14204 & n32437 ;
  assign n32439 = \m1_data_i[13]_pad  & ~n14211 ;
  assign n32440 = n14219 & n32439 ;
  assign n32441 = ~n32438 & ~n32440 ;
  assign n32442 = \m6_data_i[13]_pad  & n14211 ;
  assign n32443 = n14204 & n32442 ;
  assign n32444 = \m5_data_i[13]_pad  & ~n14211 ;
  assign n32445 = n14236 & n32444 ;
  assign n32446 = ~n32443 & ~n32445 ;
  assign n32447 = n32441 & n32446 ;
  assign n32448 = n32436 & n32447 ;
  assign n32449 = \m3_data_i[14]_pad  & ~n14211 ;
  assign n32450 = n14228 & n32449 ;
  assign n32451 = \m4_data_i[14]_pad  & n14211 ;
  assign n32452 = n14236 & n32451 ;
  assign n32453 = ~n32450 & ~n32452 ;
  assign n32454 = \m6_data_i[14]_pad  & n14211 ;
  assign n32455 = n14204 & n32454 ;
  assign n32456 = \m2_data_i[14]_pad  & n14211 ;
  assign n32457 = n14228 & n32456 ;
  assign n32458 = ~n32455 & ~n32457 ;
  assign n32459 = n32453 & n32458 ;
  assign n32460 = \m5_data_i[14]_pad  & ~n14211 ;
  assign n32461 = n14236 & n32460 ;
  assign n32462 = \m1_data_i[14]_pad  & ~n14211 ;
  assign n32463 = n14219 & n32462 ;
  assign n32464 = ~n32461 & ~n32463 ;
  assign n32465 = \m0_data_i[14]_pad  & n14211 ;
  assign n32466 = n14219 & n32465 ;
  assign n32467 = \m7_data_i[14]_pad  & ~n14211 ;
  assign n32468 = n14204 & n32467 ;
  assign n32469 = ~n32466 & ~n32468 ;
  assign n32470 = n32464 & n32469 ;
  assign n32471 = n32459 & n32470 ;
  assign n32472 = \m3_data_i[15]_pad  & ~n14211 ;
  assign n32473 = n14228 & n32472 ;
  assign n32474 = \m4_data_i[15]_pad  & n14211 ;
  assign n32475 = n14236 & n32474 ;
  assign n32476 = ~n32473 & ~n32475 ;
  assign n32477 = \m6_data_i[15]_pad  & n14211 ;
  assign n32478 = n14204 & n32477 ;
  assign n32479 = \m2_data_i[15]_pad  & n14211 ;
  assign n32480 = n14228 & n32479 ;
  assign n32481 = ~n32478 & ~n32480 ;
  assign n32482 = n32476 & n32481 ;
  assign n32483 = \m5_data_i[15]_pad  & ~n14211 ;
  assign n32484 = n14236 & n32483 ;
  assign n32485 = \m1_data_i[15]_pad  & ~n14211 ;
  assign n32486 = n14219 & n32485 ;
  assign n32487 = ~n32484 & ~n32486 ;
  assign n32488 = \m0_data_i[15]_pad  & n14211 ;
  assign n32489 = n14219 & n32488 ;
  assign n32490 = \m7_data_i[15]_pad  & ~n14211 ;
  assign n32491 = n14204 & n32490 ;
  assign n32492 = ~n32489 & ~n32491 ;
  assign n32493 = n32487 & n32492 ;
  assign n32494 = n32482 & n32493 ;
  assign n32495 = \m3_data_i[16]_pad  & ~n14211 ;
  assign n32496 = n14228 & n32495 ;
  assign n32497 = \m4_data_i[16]_pad  & n14211 ;
  assign n32498 = n14236 & n32497 ;
  assign n32499 = ~n32496 & ~n32498 ;
  assign n32500 = \m6_data_i[16]_pad  & n14211 ;
  assign n32501 = n14204 & n32500 ;
  assign n32502 = \m2_data_i[16]_pad  & n14211 ;
  assign n32503 = n14228 & n32502 ;
  assign n32504 = ~n32501 & ~n32503 ;
  assign n32505 = n32499 & n32504 ;
  assign n32506 = \m5_data_i[16]_pad  & ~n14211 ;
  assign n32507 = n14236 & n32506 ;
  assign n32508 = \m1_data_i[16]_pad  & ~n14211 ;
  assign n32509 = n14219 & n32508 ;
  assign n32510 = ~n32507 & ~n32509 ;
  assign n32511 = \m0_data_i[16]_pad  & n14211 ;
  assign n32512 = n14219 & n32511 ;
  assign n32513 = \m7_data_i[16]_pad  & ~n14211 ;
  assign n32514 = n14204 & n32513 ;
  assign n32515 = ~n32512 & ~n32514 ;
  assign n32516 = n32510 & n32515 ;
  assign n32517 = n32505 & n32516 ;
  assign n32518 = \m3_data_i[17]_pad  & ~n14211 ;
  assign n32519 = n14228 & n32518 ;
  assign n32520 = \m4_data_i[17]_pad  & n14211 ;
  assign n32521 = n14236 & n32520 ;
  assign n32522 = ~n32519 & ~n32521 ;
  assign n32523 = \m6_data_i[17]_pad  & n14211 ;
  assign n32524 = n14204 & n32523 ;
  assign n32525 = \m2_data_i[17]_pad  & n14211 ;
  assign n32526 = n14228 & n32525 ;
  assign n32527 = ~n32524 & ~n32526 ;
  assign n32528 = n32522 & n32527 ;
  assign n32529 = \m5_data_i[17]_pad  & ~n14211 ;
  assign n32530 = n14236 & n32529 ;
  assign n32531 = \m1_data_i[17]_pad  & ~n14211 ;
  assign n32532 = n14219 & n32531 ;
  assign n32533 = ~n32530 & ~n32532 ;
  assign n32534 = \m0_data_i[17]_pad  & n14211 ;
  assign n32535 = n14219 & n32534 ;
  assign n32536 = \m7_data_i[17]_pad  & ~n14211 ;
  assign n32537 = n14204 & n32536 ;
  assign n32538 = ~n32535 & ~n32537 ;
  assign n32539 = n32533 & n32538 ;
  assign n32540 = n32528 & n32539 ;
  assign n32541 = \m3_data_i[18]_pad  & ~n14211 ;
  assign n32542 = n14228 & n32541 ;
  assign n32543 = \m4_data_i[18]_pad  & n14211 ;
  assign n32544 = n14236 & n32543 ;
  assign n32545 = ~n32542 & ~n32544 ;
  assign n32546 = \m6_data_i[18]_pad  & n14211 ;
  assign n32547 = n14204 & n32546 ;
  assign n32548 = \m2_data_i[18]_pad  & n14211 ;
  assign n32549 = n14228 & n32548 ;
  assign n32550 = ~n32547 & ~n32549 ;
  assign n32551 = n32545 & n32550 ;
  assign n32552 = \m5_data_i[18]_pad  & ~n14211 ;
  assign n32553 = n14236 & n32552 ;
  assign n32554 = \m1_data_i[18]_pad  & ~n14211 ;
  assign n32555 = n14219 & n32554 ;
  assign n32556 = ~n32553 & ~n32555 ;
  assign n32557 = \m0_data_i[18]_pad  & n14211 ;
  assign n32558 = n14219 & n32557 ;
  assign n32559 = \m7_data_i[18]_pad  & ~n14211 ;
  assign n32560 = n14204 & n32559 ;
  assign n32561 = ~n32558 & ~n32560 ;
  assign n32562 = n32556 & n32561 ;
  assign n32563 = n32551 & n32562 ;
  assign n32564 = \m3_data_i[19]_pad  & ~n14211 ;
  assign n32565 = n14228 & n32564 ;
  assign n32566 = \m4_data_i[19]_pad  & n14211 ;
  assign n32567 = n14236 & n32566 ;
  assign n32568 = ~n32565 & ~n32567 ;
  assign n32569 = \m6_data_i[19]_pad  & n14211 ;
  assign n32570 = n14204 & n32569 ;
  assign n32571 = \m2_data_i[19]_pad  & n14211 ;
  assign n32572 = n14228 & n32571 ;
  assign n32573 = ~n32570 & ~n32572 ;
  assign n32574 = n32568 & n32573 ;
  assign n32575 = \m5_data_i[19]_pad  & ~n14211 ;
  assign n32576 = n14236 & n32575 ;
  assign n32577 = \m1_data_i[19]_pad  & ~n14211 ;
  assign n32578 = n14219 & n32577 ;
  assign n32579 = ~n32576 & ~n32578 ;
  assign n32580 = \m0_data_i[19]_pad  & n14211 ;
  assign n32581 = n14219 & n32580 ;
  assign n32582 = \m7_data_i[19]_pad  & ~n14211 ;
  assign n32583 = n14204 & n32582 ;
  assign n32584 = ~n32581 & ~n32583 ;
  assign n32585 = n32579 & n32584 ;
  assign n32586 = n32574 & n32585 ;
  assign n32587 = \m1_data_i[1]_pad  & ~n14211 ;
  assign n32588 = n14219 & n32587 ;
  assign n32589 = \m2_data_i[1]_pad  & n14211 ;
  assign n32590 = n14228 & n32589 ;
  assign n32591 = ~n32588 & ~n32590 ;
  assign n32592 = \m0_data_i[1]_pad  & n14211 ;
  assign n32593 = n14219 & n32592 ;
  assign n32594 = \m5_data_i[1]_pad  & ~n14211 ;
  assign n32595 = n14236 & n32594 ;
  assign n32596 = ~n32593 & ~n32595 ;
  assign n32597 = n32591 & n32596 ;
  assign n32598 = \m7_data_i[1]_pad  & ~n14211 ;
  assign n32599 = n14204 & n32598 ;
  assign n32600 = \m6_data_i[1]_pad  & n14211 ;
  assign n32601 = n14204 & n32600 ;
  assign n32602 = ~n32599 & ~n32601 ;
  assign n32603 = \m3_data_i[1]_pad  & ~n14211 ;
  assign n32604 = n14228 & n32603 ;
  assign n32605 = \m4_data_i[1]_pad  & n14211 ;
  assign n32606 = n14236 & n32605 ;
  assign n32607 = ~n32604 & ~n32606 ;
  assign n32608 = n32602 & n32607 ;
  assign n32609 = n32597 & n32608 ;
  assign n32610 = \m1_data_i[20]_pad  & ~n14211 ;
  assign n32611 = n14219 & n32610 ;
  assign n32612 = \m2_data_i[20]_pad  & n14211 ;
  assign n32613 = n14228 & n32612 ;
  assign n32614 = ~n32611 & ~n32613 ;
  assign n32615 = \m0_data_i[20]_pad  & n14211 ;
  assign n32616 = n14219 & n32615 ;
  assign n32617 = \m4_data_i[20]_pad  & n14211 ;
  assign n32618 = n14236 & n32617 ;
  assign n32619 = ~n32616 & ~n32618 ;
  assign n32620 = n32614 & n32619 ;
  assign n32621 = \m7_data_i[20]_pad  & ~n14211 ;
  assign n32622 = n14204 & n32621 ;
  assign n32623 = \m3_data_i[20]_pad  & ~n14211 ;
  assign n32624 = n14228 & n32623 ;
  assign n32625 = ~n32622 & ~n32624 ;
  assign n32626 = \m6_data_i[20]_pad  & n14211 ;
  assign n32627 = n14204 & n32626 ;
  assign n32628 = \m5_data_i[20]_pad  & ~n14211 ;
  assign n32629 = n14236 & n32628 ;
  assign n32630 = ~n32627 & ~n32629 ;
  assign n32631 = n32625 & n32630 ;
  assign n32632 = n32620 & n32631 ;
  assign n32633 = \m1_data_i[21]_pad  & ~n14211 ;
  assign n32634 = n14219 & n32633 ;
  assign n32635 = \m2_data_i[21]_pad  & n14211 ;
  assign n32636 = n14228 & n32635 ;
  assign n32637 = ~n32634 & ~n32636 ;
  assign n32638 = \m0_data_i[21]_pad  & n14211 ;
  assign n32639 = n14219 & n32638 ;
  assign n32640 = \m4_data_i[21]_pad  & n14211 ;
  assign n32641 = n14236 & n32640 ;
  assign n32642 = ~n32639 & ~n32641 ;
  assign n32643 = n32637 & n32642 ;
  assign n32644 = \m7_data_i[21]_pad  & ~n14211 ;
  assign n32645 = n14204 & n32644 ;
  assign n32646 = \m3_data_i[21]_pad  & ~n14211 ;
  assign n32647 = n14228 & n32646 ;
  assign n32648 = ~n32645 & ~n32647 ;
  assign n32649 = \m6_data_i[21]_pad  & n14211 ;
  assign n32650 = n14204 & n32649 ;
  assign n32651 = \m5_data_i[21]_pad  & ~n14211 ;
  assign n32652 = n14236 & n32651 ;
  assign n32653 = ~n32650 & ~n32652 ;
  assign n32654 = n32648 & n32653 ;
  assign n32655 = n32643 & n32654 ;
  assign n32656 = \m1_data_i[22]_pad  & ~n14211 ;
  assign n32657 = n14219 & n32656 ;
  assign n32658 = \m2_data_i[22]_pad  & n14211 ;
  assign n32659 = n14228 & n32658 ;
  assign n32660 = ~n32657 & ~n32659 ;
  assign n32661 = \m0_data_i[22]_pad  & n14211 ;
  assign n32662 = n14219 & n32661 ;
  assign n32663 = \m5_data_i[22]_pad  & ~n14211 ;
  assign n32664 = n14236 & n32663 ;
  assign n32665 = ~n32662 & ~n32664 ;
  assign n32666 = n32660 & n32665 ;
  assign n32667 = \m7_data_i[22]_pad  & ~n14211 ;
  assign n32668 = n14204 & n32667 ;
  assign n32669 = \m6_data_i[22]_pad  & n14211 ;
  assign n32670 = n14204 & n32669 ;
  assign n32671 = ~n32668 & ~n32670 ;
  assign n32672 = \m3_data_i[22]_pad  & ~n14211 ;
  assign n32673 = n14228 & n32672 ;
  assign n32674 = \m4_data_i[22]_pad  & n14211 ;
  assign n32675 = n14236 & n32674 ;
  assign n32676 = ~n32673 & ~n32675 ;
  assign n32677 = n32671 & n32676 ;
  assign n32678 = n32666 & n32677 ;
  assign n32679 = \m1_data_i[23]_pad  & ~n14211 ;
  assign n32680 = n14219 & n32679 ;
  assign n32681 = \m2_data_i[23]_pad  & n14211 ;
  assign n32682 = n14228 & n32681 ;
  assign n32683 = ~n32680 & ~n32682 ;
  assign n32684 = \m0_data_i[23]_pad  & n14211 ;
  assign n32685 = n14219 & n32684 ;
  assign n32686 = \m4_data_i[23]_pad  & n14211 ;
  assign n32687 = n14236 & n32686 ;
  assign n32688 = ~n32685 & ~n32687 ;
  assign n32689 = n32683 & n32688 ;
  assign n32690 = \m7_data_i[23]_pad  & ~n14211 ;
  assign n32691 = n14204 & n32690 ;
  assign n32692 = \m3_data_i[23]_pad  & ~n14211 ;
  assign n32693 = n14228 & n32692 ;
  assign n32694 = ~n32691 & ~n32693 ;
  assign n32695 = \m6_data_i[23]_pad  & n14211 ;
  assign n32696 = n14204 & n32695 ;
  assign n32697 = \m5_data_i[23]_pad  & ~n14211 ;
  assign n32698 = n14236 & n32697 ;
  assign n32699 = ~n32696 & ~n32698 ;
  assign n32700 = n32694 & n32699 ;
  assign n32701 = n32689 & n32700 ;
  assign n32702 = \m3_data_i[24]_pad  & ~n14211 ;
  assign n32703 = n14228 & n32702 ;
  assign n32704 = \m4_data_i[24]_pad  & n14211 ;
  assign n32705 = n14236 & n32704 ;
  assign n32706 = ~n32703 & ~n32705 ;
  assign n32707 = \m6_data_i[24]_pad  & n14211 ;
  assign n32708 = n14204 & n32707 ;
  assign n32709 = \m2_data_i[24]_pad  & n14211 ;
  assign n32710 = n14228 & n32709 ;
  assign n32711 = ~n32708 & ~n32710 ;
  assign n32712 = n32706 & n32711 ;
  assign n32713 = \m5_data_i[24]_pad  & ~n14211 ;
  assign n32714 = n14236 & n32713 ;
  assign n32715 = \m1_data_i[24]_pad  & ~n14211 ;
  assign n32716 = n14219 & n32715 ;
  assign n32717 = ~n32714 & ~n32716 ;
  assign n32718 = \m0_data_i[24]_pad  & n14211 ;
  assign n32719 = n14219 & n32718 ;
  assign n32720 = \m7_data_i[24]_pad  & ~n14211 ;
  assign n32721 = n14204 & n32720 ;
  assign n32722 = ~n32719 & ~n32721 ;
  assign n32723 = n32717 & n32722 ;
  assign n32724 = n32712 & n32723 ;
  assign n32725 = \m3_data_i[25]_pad  & ~n14211 ;
  assign n32726 = n14228 & n32725 ;
  assign n32727 = \m4_data_i[25]_pad  & n14211 ;
  assign n32728 = n14236 & n32727 ;
  assign n32729 = ~n32726 & ~n32728 ;
  assign n32730 = \m6_data_i[25]_pad  & n14211 ;
  assign n32731 = n14204 & n32730 ;
  assign n32732 = \m2_data_i[25]_pad  & n14211 ;
  assign n32733 = n14228 & n32732 ;
  assign n32734 = ~n32731 & ~n32733 ;
  assign n32735 = n32729 & n32734 ;
  assign n32736 = \m5_data_i[25]_pad  & ~n14211 ;
  assign n32737 = n14236 & n32736 ;
  assign n32738 = \m1_data_i[25]_pad  & ~n14211 ;
  assign n32739 = n14219 & n32738 ;
  assign n32740 = ~n32737 & ~n32739 ;
  assign n32741 = \m0_data_i[25]_pad  & n14211 ;
  assign n32742 = n14219 & n32741 ;
  assign n32743 = \m7_data_i[25]_pad  & ~n14211 ;
  assign n32744 = n14204 & n32743 ;
  assign n32745 = ~n32742 & ~n32744 ;
  assign n32746 = n32740 & n32745 ;
  assign n32747 = n32735 & n32746 ;
  assign n32748 = \m3_data_i[26]_pad  & ~n14211 ;
  assign n32749 = n14228 & n32748 ;
  assign n32750 = \m4_data_i[26]_pad  & n14211 ;
  assign n32751 = n14236 & n32750 ;
  assign n32752 = ~n32749 & ~n32751 ;
  assign n32753 = \m6_data_i[26]_pad  & n14211 ;
  assign n32754 = n14204 & n32753 ;
  assign n32755 = \m2_data_i[26]_pad  & n14211 ;
  assign n32756 = n14228 & n32755 ;
  assign n32757 = ~n32754 & ~n32756 ;
  assign n32758 = n32752 & n32757 ;
  assign n32759 = \m5_data_i[26]_pad  & ~n14211 ;
  assign n32760 = n14236 & n32759 ;
  assign n32761 = \m1_data_i[26]_pad  & ~n14211 ;
  assign n32762 = n14219 & n32761 ;
  assign n32763 = ~n32760 & ~n32762 ;
  assign n32764 = \m0_data_i[26]_pad  & n14211 ;
  assign n32765 = n14219 & n32764 ;
  assign n32766 = \m7_data_i[26]_pad  & ~n14211 ;
  assign n32767 = n14204 & n32766 ;
  assign n32768 = ~n32765 & ~n32767 ;
  assign n32769 = n32763 & n32768 ;
  assign n32770 = n32758 & n32769 ;
  assign n32771 = \m3_data_i[27]_pad  & ~n14211 ;
  assign n32772 = n14228 & n32771 ;
  assign n32773 = \m4_data_i[27]_pad  & n14211 ;
  assign n32774 = n14236 & n32773 ;
  assign n32775 = ~n32772 & ~n32774 ;
  assign n32776 = \m6_data_i[27]_pad  & n14211 ;
  assign n32777 = n14204 & n32776 ;
  assign n32778 = \m2_data_i[27]_pad  & n14211 ;
  assign n32779 = n14228 & n32778 ;
  assign n32780 = ~n32777 & ~n32779 ;
  assign n32781 = n32775 & n32780 ;
  assign n32782 = \m5_data_i[27]_pad  & ~n14211 ;
  assign n32783 = n14236 & n32782 ;
  assign n32784 = \m1_data_i[27]_pad  & ~n14211 ;
  assign n32785 = n14219 & n32784 ;
  assign n32786 = ~n32783 & ~n32785 ;
  assign n32787 = \m0_data_i[27]_pad  & n14211 ;
  assign n32788 = n14219 & n32787 ;
  assign n32789 = \m7_data_i[27]_pad  & ~n14211 ;
  assign n32790 = n14204 & n32789 ;
  assign n32791 = ~n32788 & ~n32790 ;
  assign n32792 = n32786 & n32791 ;
  assign n32793 = n32781 & n32792 ;
  assign n32794 = \m3_data_i[28]_pad  & ~n14211 ;
  assign n32795 = n14228 & n32794 ;
  assign n32796 = \m4_data_i[28]_pad  & n14211 ;
  assign n32797 = n14236 & n32796 ;
  assign n32798 = ~n32795 & ~n32797 ;
  assign n32799 = \m6_data_i[28]_pad  & n14211 ;
  assign n32800 = n14204 & n32799 ;
  assign n32801 = \m2_data_i[28]_pad  & n14211 ;
  assign n32802 = n14228 & n32801 ;
  assign n32803 = ~n32800 & ~n32802 ;
  assign n32804 = n32798 & n32803 ;
  assign n32805 = \m5_data_i[28]_pad  & ~n14211 ;
  assign n32806 = n14236 & n32805 ;
  assign n32807 = \m1_data_i[28]_pad  & ~n14211 ;
  assign n32808 = n14219 & n32807 ;
  assign n32809 = ~n32806 & ~n32808 ;
  assign n32810 = \m0_data_i[28]_pad  & n14211 ;
  assign n32811 = n14219 & n32810 ;
  assign n32812 = \m7_data_i[28]_pad  & ~n14211 ;
  assign n32813 = n14204 & n32812 ;
  assign n32814 = ~n32811 & ~n32813 ;
  assign n32815 = n32809 & n32814 ;
  assign n32816 = n32804 & n32815 ;
  assign n32817 = \m3_data_i[29]_pad  & ~n14211 ;
  assign n32818 = n14228 & n32817 ;
  assign n32819 = \m4_data_i[29]_pad  & n14211 ;
  assign n32820 = n14236 & n32819 ;
  assign n32821 = ~n32818 & ~n32820 ;
  assign n32822 = \m6_data_i[29]_pad  & n14211 ;
  assign n32823 = n14204 & n32822 ;
  assign n32824 = \m2_data_i[29]_pad  & n14211 ;
  assign n32825 = n14228 & n32824 ;
  assign n32826 = ~n32823 & ~n32825 ;
  assign n32827 = n32821 & n32826 ;
  assign n32828 = \m5_data_i[29]_pad  & ~n14211 ;
  assign n32829 = n14236 & n32828 ;
  assign n32830 = \m1_data_i[29]_pad  & ~n14211 ;
  assign n32831 = n14219 & n32830 ;
  assign n32832 = ~n32829 & ~n32831 ;
  assign n32833 = \m0_data_i[29]_pad  & n14211 ;
  assign n32834 = n14219 & n32833 ;
  assign n32835 = \m7_data_i[29]_pad  & ~n14211 ;
  assign n32836 = n14204 & n32835 ;
  assign n32837 = ~n32834 & ~n32836 ;
  assign n32838 = n32832 & n32837 ;
  assign n32839 = n32827 & n32838 ;
  assign n32840 = \m0_data_i[2]_pad  & n14211 ;
  assign n32841 = n14219 & n32840 ;
  assign n32842 = \m7_data_i[2]_pad  & ~n14211 ;
  assign n32843 = n14204 & n32842 ;
  assign n32844 = ~n32841 & ~n32843 ;
  assign n32845 = \m1_data_i[2]_pad  & ~n14211 ;
  assign n32846 = n14219 & n32845 ;
  assign n32847 = \m5_data_i[2]_pad  & ~n14211 ;
  assign n32848 = n14236 & n32847 ;
  assign n32849 = ~n32846 & ~n32848 ;
  assign n32850 = n32844 & n32849 ;
  assign n32851 = \m2_data_i[2]_pad  & n14211 ;
  assign n32852 = n14228 & n32851 ;
  assign n32853 = \m6_data_i[2]_pad  & n14211 ;
  assign n32854 = n14204 & n32853 ;
  assign n32855 = ~n32852 & ~n32854 ;
  assign n32856 = \m3_data_i[2]_pad  & ~n14211 ;
  assign n32857 = n14228 & n32856 ;
  assign n32858 = \m4_data_i[2]_pad  & n14211 ;
  assign n32859 = n14236 & n32858 ;
  assign n32860 = ~n32857 & ~n32859 ;
  assign n32861 = n32855 & n32860 ;
  assign n32862 = n32850 & n32861 ;
  assign n32863 = \m3_data_i[30]_pad  & ~n14211 ;
  assign n32864 = n14228 & n32863 ;
  assign n32865 = \m4_data_i[30]_pad  & n14211 ;
  assign n32866 = n14236 & n32865 ;
  assign n32867 = ~n32864 & ~n32866 ;
  assign n32868 = \m6_data_i[30]_pad  & n14211 ;
  assign n32869 = n14204 & n32868 ;
  assign n32870 = \m2_data_i[30]_pad  & n14211 ;
  assign n32871 = n14228 & n32870 ;
  assign n32872 = ~n32869 & ~n32871 ;
  assign n32873 = n32867 & n32872 ;
  assign n32874 = \m5_data_i[30]_pad  & ~n14211 ;
  assign n32875 = n14236 & n32874 ;
  assign n32876 = \m1_data_i[30]_pad  & ~n14211 ;
  assign n32877 = n14219 & n32876 ;
  assign n32878 = ~n32875 & ~n32877 ;
  assign n32879 = \m0_data_i[30]_pad  & n14211 ;
  assign n32880 = n14219 & n32879 ;
  assign n32881 = \m7_data_i[30]_pad  & ~n14211 ;
  assign n32882 = n14204 & n32881 ;
  assign n32883 = ~n32880 & ~n32882 ;
  assign n32884 = n32878 & n32883 ;
  assign n32885 = n32873 & n32884 ;
  assign n32886 = \m3_data_i[31]_pad  & ~n14211 ;
  assign n32887 = n14228 & n32886 ;
  assign n32888 = \m4_data_i[31]_pad  & n14211 ;
  assign n32889 = n14236 & n32888 ;
  assign n32890 = ~n32887 & ~n32889 ;
  assign n32891 = \m6_data_i[31]_pad  & n14211 ;
  assign n32892 = n14204 & n32891 ;
  assign n32893 = \m2_data_i[31]_pad  & n14211 ;
  assign n32894 = n14228 & n32893 ;
  assign n32895 = ~n32892 & ~n32894 ;
  assign n32896 = n32890 & n32895 ;
  assign n32897 = \m5_data_i[31]_pad  & ~n14211 ;
  assign n32898 = n14236 & n32897 ;
  assign n32899 = \m1_data_i[31]_pad  & ~n14211 ;
  assign n32900 = n14219 & n32899 ;
  assign n32901 = ~n32898 & ~n32900 ;
  assign n32902 = \m0_data_i[31]_pad  & n14211 ;
  assign n32903 = n14219 & n32902 ;
  assign n32904 = \m7_data_i[31]_pad  & ~n14211 ;
  assign n32905 = n14204 & n32904 ;
  assign n32906 = ~n32903 & ~n32905 ;
  assign n32907 = n32901 & n32906 ;
  assign n32908 = n32896 & n32907 ;
  assign n32909 = \m3_data_i[3]_pad  & ~n14211 ;
  assign n32910 = n14228 & n32909 ;
  assign n32911 = \m4_data_i[3]_pad  & n14211 ;
  assign n32912 = n14236 & n32911 ;
  assign n32913 = ~n32910 & ~n32912 ;
  assign n32914 = \m6_data_i[3]_pad  & n14211 ;
  assign n32915 = n14204 & n32914 ;
  assign n32916 = \m7_data_i[3]_pad  & ~n14211 ;
  assign n32917 = n14204 & n32916 ;
  assign n32918 = ~n32915 & ~n32917 ;
  assign n32919 = n32913 & n32918 ;
  assign n32920 = \m5_data_i[3]_pad  & ~n14211 ;
  assign n32921 = n14236 & n32920 ;
  assign n32922 = \m0_data_i[3]_pad  & n14211 ;
  assign n32923 = n14219 & n32922 ;
  assign n32924 = ~n32921 & ~n32923 ;
  assign n32925 = \m1_data_i[3]_pad  & ~n14211 ;
  assign n32926 = n14219 & n32925 ;
  assign n32927 = \m2_data_i[3]_pad  & n14211 ;
  assign n32928 = n14228 & n32927 ;
  assign n32929 = ~n32926 & ~n32928 ;
  assign n32930 = n32924 & n32929 ;
  assign n32931 = n32919 & n32930 ;
  assign n32932 = \m6_data_i[4]_pad  & n14211 ;
  assign n32933 = n14204 & n32932 ;
  assign n32934 = \m5_data_i[4]_pad  & ~n14211 ;
  assign n32935 = n14236 & n32934 ;
  assign n32936 = ~n32933 & ~n32935 ;
  assign n32937 = \m1_data_i[4]_pad  & ~n14211 ;
  assign n32938 = n14219 & n32937 ;
  assign n32939 = \m4_data_i[4]_pad  & n14211 ;
  assign n32940 = n14236 & n32939 ;
  assign n32941 = ~n32938 & ~n32940 ;
  assign n32942 = n32936 & n32941 ;
  assign n32943 = \m2_data_i[4]_pad  & n14211 ;
  assign n32944 = n14228 & n32943 ;
  assign n32945 = \m3_data_i[4]_pad  & ~n14211 ;
  assign n32946 = n14228 & n32945 ;
  assign n32947 = ~n32944 & ~n32946 ;
  assign n32948 = \m0_data_i[4]_pad  & n14211 ;
  assign n32949 = n14219 & n32948 ;
  assign n32950 = \m7_data_i[4]_pad  & ~n14211 ;
  assign n32951 = n14204 & n32950 ;
  assign n32952 = ~n32949 & ~n32951 ;
  assign n32953 = n32947 & n32952 ;
  assign n32954 = n32942 & n32953 ;
  assign n32955 = \m1_data_i[5]_pad  & ~n14211 ;
  assign n32956 = n14219 & n32955 ;
  assign n32957 = \m2_data_i[5]_pad  & n14211 ;
  assign n32958 = n14228 & n32957 ;
  assign n32959 = ~n32956 & ~n32958 ;
  assign n32960 = \m3_data_i[5]_pad  & ~n14211 ;
  assign n32961 = n14228 & n32960 ;
  assign n32962 = \m7_data_i[5]_pad  & ~n14211 ;
  assign n32963 = n14204 & n32962 ;
  assign n32964 = ~n32961 & ~n32963 ;
  assign n32965 = n32959 & n32964 ;
  assign n32966 = \m4_data_i[5]_pad  & n14211 ;
  assign n32967 = n14236 & n32966 ;
  assign n32968 = \m0_data_i[5]_pad  & n14211 ;
  assign n32969 = n14219 & n32968 ;
  assign n32970 = ~n32967 & ~n32969 ;
  assign n32971 = \m6_data_i[5]_pad  & n14211 ;
  assign n32972 = n14204 & n32971 ;
  assign n32973 = \m5_data_i[5]_pad  & ~n14211 ;
  assign n32974 = n14236 & n32973 ;
  assign n32975 = ~n32972 & ~n32974 ;
  assign n32976 = n32970 & n32975 ;
  assign n32977 = n32965 & n32976 ;
  assign n32978 = \m3_data_i[6]_pad  & ~n14211 ;
  assign n32979 = n14228 & n32978 ;
  assign n32980 = \m4_data_i[6]_pad  & n14211 ;
  assign n32981 = n14236 & n32980 ;
  assign n32982 = ~n32979 & ~n32981 ;
  assign n32983 = \m0_data_i[6]_pad  & n14211 ;
  assign n32984 = n14219 & n32983 ;
  assign n32985 = \m5_data_i[6]_pad  & ~n14211 ;
  assign n32986 = n14236 & n32985 ;
  assign n32987 = ~n32984 & ~n32986 ;
  assign n32988 = n32982 & n32987 ;
  assign n32989 = \m7_data_i[6]_pad  & ~n14211 ;
  assign n32990 = n14204 & n32989 ;
  assign n32991 = \m6_data_i[6]_pad  & n14211 ;
  assign n32992 = n14204 & n32991 ;
  assign n32993 = ~n32990 & ~n32992 ;
  assign n32994 = \m1_data_i[6]_pad  & ~n14211 ;
  assign n32995 = n14219 & n32994 ;
  assign n32996 = \m2_data_i[6]_pad  & n14211 ;
  assign n32997 = n14228 & n32996 ;
  assign n32998 = ~n32995 & ~n32997 ;
  assign n32999 = n32993 & n32998 ;
  assign n33000 = n32988 & n32999 ;
  assign n33001 = \m3_data_i[7]_pad  & ~n14211 ;
  assign n33002 = n14228 & n33001 ;
  assign n33003 = \m4_data_i[7]_pad  & n14211 ;
  assign n33004 = n14236 & n33003 ;
  assign n33005 = ~n33002 & ~n33004 ;
  assign n33006 = \m6_data_i[7]_pad  & n14211 ;
  assign n33007 = n14204 & n33006 ;
  assign n33008 = \m2_data_i[7]_pad  & n14211 ;
  assign n33009 = n14228 & n33008 ;
  assign n33010 = ~n33007 & ~n33009 ;
  assign n33011 = n33005 & n33010 ;
  assign n33012 = \m5_data_i[7]_pad  & ~n14211 ;
  assign n33013 = n14236 & n33012 ;
  assign n33014 = \m1_data_i[7]_pad  & ~n14211 ;
  assign n33015 = n14219 & n33014 ;
  assign n33016 = ~n33013 & ~n33015 ;
  assign n33017 = \m0_data_i[7]_pad  & n14211 ;
  assign n33018 = n14219 & n33017 ;
  assign n33019 = \m7_data_i[7]_pad  & ~n14211 ;
  assign n33020 = n14204 & n33019 ;
  assign n33021 = ~n33018 & ~n33020 ;
  assign n33022 = n33016 & n33021 ;
  assign n33023 = n33011 & n33022 ;
  assign n33024 = \m0_data_i[8]_pad  & n14211 ;
  assign n33025 = n14219 & n33024 ;
  assign n33026 = \m7_data_i[8]_pad  & ~n14211 ;
  assign n33027 = n14204 & n33026 ;
  assign n33028 = ~n33025 & ~n33027 ;
  assign n33029 = \m1_data_i[8]_pad  & ~n14211 ;
  assign n33030 = n14219 & n33029 ;
  assign n33031 = \m4_data_i[8]_pad  & n14211 ;
  assign n33032 = n14236 & n33031 ;
  assign n33033 = ~n33030 & ~n33032 ;
  assign n33034 = n33028 & n33033 ;
  assign n33035 = \m2_data_i[8]_pad  & n14211 ;
  assign n33036 = n14228 & n33035 ;
  assign n33037 = \m3_data_i[8]_pad  & ~n14211 ;
  assign n33038 = n14228 & n33037 ;
  assign n33039 = ~n33036 & ~n33038 ;
  assign n33040 = \m6_data_i[8]_pad  & n14211 ;
  assign n33041 = n14204 & n33040 ;
  assign n33042 = \m5_data_i[8]_pad  & ~n14211 ;
  assign n33043 = n14236 & n33042 ;
  assign n33044 = ~n33041 & ~n33043 ;
  assign n33045 = n33039 & n33044 ;
  assign n33046 = n33034 & n33045 ;
  assign n33047 = \m6_data_i[9]_pad  & n14211 ;
  assign n33048 = n14204 & n33047 ;
  assign n33049 = \m5_data_i[9]_pad  & ~n14211 ;
  assign n33050 = n14236 & n33049 ;
  assign n33051 = ~n33048 & ~n33050 ;
  assign n33052 = \m3_data_i[9]_pad  & ~n14211 ;
  assign n33053 = n14228 & n33052 ;
  assign n33054 = \m7_data_i[9]_pad  & ~n14211 ;
  assign n33055 = n14204 & n33054 ;
  assign n33056 = ~n33053 & ~n33055 ;
  assign n33057 = n33051 & n33056 ;
  assign n33058 = \m4_data_i[9]_pad  & n14211 ;
  assign n33059 = n14236 & n33058 ;
  assign n33060 = \m0_data_i[9]_pad  & n14211 ;
  assign n33061 = n14219 & n33060 ;
  assign n33062 = ~n33059 & ~n33061 ;
  assign n33063 = \m1_data_i[9]_pad  & ~n14211 ;
  assign n33064 = n14219 & n33063 ;
  assign n33065 = \m2_data_i[9]_pad  & n14211 ;
  assign n33066 = n14228 & n33065 ;
  assign n33067 = ~n33064 & ~n33066 ;
  assign n33068 = n33062 & n33067 ;
  assign n33069 = n33057 & n33068 ;
  assign n33070 = \m3_sel_i[0]_pad  & ~n14211 ;
  assign n33071 = n14228 & n33070 ;
  assign n33072 = \m4_sel_i[0]_pad  & n14211 ;
  assign n33073 = n14236 & n33072 ;
  assign n33074 = ~n33071 & ~n33073 ;
  assign n33075 = \m6_sel_i[0]_pad  & n14211 ;
  assign n33076 = n14204 & n33075 ;
  assign n33077 = \m2_sel_i[0]_pad  & n14211 ;
  assign n33078 = n14228 & n33077 ;
  assign n33079 = ~n33076 & ~n33078 ;
  assign n33080 = n33074 & n33079 ;
  assign n33081 = \m5_sel_i[0]_pad  & ~n14211 ;
  assign n33082 = n14236 & n33081 ;
  assign n33083 = \m1_sel_i[0]_pad  & ~n14211 ;
  assign n33084 = n14219 & n33083 ;
  assign n33085 = ~n33082 & ~n33084 ;
  assign n33086 = \m0_sel_i[0]_pad  & n14211 ;
  assign n33087 = n14219 & n33086 ;
  assign n33088 = \m7_sel_i[0]_pad  & ~n14211 ;
  assign n33089 = n14204 & n33088 ;
  assign n33090 = ~n33087 & ~n33089 ;
  assign n33091 = n33085 & n33090 ;
  assign n33092 = n33080 & n33091 ;
  assign n33093 = \m3_sel_i[1]_pad  & ~n14211 ;
  assign n33094 = n14228 & n33093 ;
  assign n33095 = \m4_sel_i[1]_pad  & n14211 ;
  assign n33096 = n14236 & n33095 ;
  assign n33097 = ~n33094 & ~n33096 ;
  assign n33098 = \m6_sel_i[1]_pad  & n14211 ;
  assign n33099 = n14204 & n33098 ;
  assign n33100 = \m2_sel_i[1]_pad  & n14211 ;
  assign n33101 = n14228 & n33100 ;
  assign n33102 = ~n33099 & ~n33101 ;
  assign n33103 = n33097 & n33102 ;
  assign n33104 = \m5_sel_i[1]_pad  & ~n14211 ;
  assign n33105 = n14236 & n33104 ;
  assign n33106 = \m1_sel_i[1]_pad  & ~n14211 ;
  assign n33107 = n14219 & n33106 ;
  assign n33108 = ~n33105 & ~n33107 ;
  assign n33109 = \m0_sel_i[1]_pad  & n14211 ;
  assign n33110 = n14219 & n33109 ;
  assign n33111 = \m7_sel_i[1]_pad  & ~n14211 ;
  assign n33112 = n14204 & n33111 ;
  assign n33113 = ~n33110 & ~n33112 ;
  assign n33114 = n33108 & n33113 ;
  assign n33115 = n33103 & n33114 ;
  assign n33116 = \m6_sel_i[2]_pad  & n14211 ;
  assign n33117 = n14204 & n33116 ;
  assign n33118 = \m5_sel_i[2]_pad  & ~n14211 ;
  assign n33119 = n14236 & n33118 ;
  assign n33120 = ~n33117 & ~n33119 ;
  assign n33121 = \m0_sel_i[2]_pad  & n14211 ;
  assign n33122 = n14219 & n33121 ;
  assign n33123 = \m4_sel_i[2]_pad  & n14211 ;
  assign n33124 = n14236 & n33123 ;
  assign n33125 = ~n33122 & ~n33124 ;
  assign n33126 = n33120 & n33125 ;
  assign n33127 = \m7_sel_i[2]_pad  & ~n14211 ;
  assign n33128 = n14204 & n33127 ;
  assign n33129 = \m3_sel_i[2]_pad  & ~n14211 ;
  assign n33130 = n14228 & n33129 ;
  assign n33131 = ~n33128 & ~n33130 ;
  assign n33132 = \m1_sel_i[2]_pad  & ~n14211 ;
  assign n33133 = n14219 & n33132 ;
  assign n33134 = \m2_sel_i[2]_pad  & n14211 ;
  assign n33135 = n14228 & n33134 ;
  assign n33136 = ~n33133 & ~n33135 ;
  assign n33137 = n33131 & n33136 ;
  assign n33138 = n33126 & n33137 ;
  assign n33139 = \m6_sel_i[3]_pad  & n14211 ;
  assign n33140 = n14204 & n33139 ;
  assign n33141 = \m5_sel_i[3]_pad  & ~n14211 ;
  assign n33142 = n14236 & n33141 ;
  assign n33143 = ~n33140 & ~n33142 ;
  assign n33144 = \m0_sel_i[3]_pad  & n14211 ;
  assign n33145 = n14219 & n33144 ;
  assign n33146 = \m4_sel_i[3]_pad  & n14211 ;
  assign n33147 = n14236 & n33146 ;
  assign n33148 = ~n33145 & ~n33147 ;
  assign n33149 = n33143 & n33148 ;
  assign n33150 = \m7_sel_i[3]_pad  & ~n14211 ;
  assign n33151 = n14204 & n33150 ;
  assign n33152 = \m3_sel_i[3]_pad  & ~n14211 ;
  assign n33153 = n14228 & n33152 ;
  assign n33154 = ~n33151 & ~n33153 ;
  assign n33155 = \m1_sel_i[3]_pad  & ~n14211 ;
  assign n33156 = n14219 & n33155 ;
  assign n33157 = \m2_sel_i[3]_pad  & n14211 ;
  assign n33158 = n14228 & n33157 ;
  assign n33159 = ~n33156 & ~n33158 ;
  assign n33160 = n33154 & n33159 ;
  assign n33161 = n33149 & n33160 ;
  assign n33162 = \m3_stb_i_pad  & n14904 ;
  assign n33163 = ~n14211 & n33162 ;
  assign n33164 = n14228 & n33163 ;
  assign n33165 = \m2_stb_i_pad  & n15094 ;
  assign n33166 = n14211 & n33165 ;
  assign n33167 = n14228 & n33166 ;
  assign n33168 = ~n33164 & ~n33167 ;
  assign n33169 = \m6_stb_i_pad  & n15011 ;
  assign n33170 = n14211 & n33169 ;
  assign n33171 = n14204 & n33170 ;
  assign n33172 = \m7_stb_i_pad  & n15055 ;
  assign n33173 = ~n14211 & n33172 ;
  assign n33174 = n14204 & n33173 ;
  assign n33175 = ~n33171 & ~n33174 ;
  assign n33176 = n33168 & n33175 ;
  assign n33177 = \m1_stb_i_pad  & n14805 ;
  assign n33178 = ~n14211 & n33177 ;
  assign n33179 = n14219 & n33178 ;
  assign n33180 = \m5_stb_i_pad  & n14971 ;
  assign n33181 = ~n14211 & n33180 ;
  assign n33182 = n14236 & n33181 ;
  assign n33183 = ~n33179 & ~n33182 ;
  assign n33184 = \m4_stb_i_pad  & n14731 ;
  assign n33185 = n14211 & n33184 ;
  assign n33186 = n14236 & n33185 ;
  assign n33187 = \m0_stb_i_pad  & n15118 ;
  assign n33188 = n14211 & n33187 ;
  assign n33189 = n14219 & n33188 ;
  assign n33190 = ~n33186 & ~n33189 ;
  assign n33191 = n33183 & n33190 ;
  assign n33192 = n33176 & n33191 ;
  assign n33193 = \m3_we_i_pad  & ~n14211 ;
  assign n33194 = n14228 & n33193 ;
  assign n33195 = \m4_we_i_pad  & n14211 ;
  assign n33196 = n14236 & n33195 ;
  assign n33197 = ~n33194 & ~n33196 ;
  assign n33198 = \m6_we_i_pad  & n14211 ;
  assign n33199 = n14204 & n33198 ;
  assign n33200 = \m2_we_i_pad  & n14211 ;
  assign n33201 = n14228 & n33200 ;
  assign n33202 = ~n33199 & ~n33201 ;
  assign n33203 = n33197 & n33202 ;
  assign n33204 = \m5_we_i_pad  & ~n14211 ;
  assign n33205 = n14236 & n33204 ;
  assign n33206 = \m1_we_i_pad  & ~n14211 ;
  assign n33207 = n14219 & n33206 ;
  assign n33208 = ~n33205 & ~n33207 ;
  assign n33209 = \m0_we_i_pad  & n14211 ;
  assign n33210 = n14219 & n33209 ;
  assign n33211 = \m7_we_i_pad  & ~n14211 ;
  assign n33212 = n14204 & n33211 ;
  assign n33213 = ~n33210 & ~n33212 ;
  assign n33214 = n33208 & n33213 ;
  assign n33215 = n33203 & n33214 ;
  assign n33216 = \m3_addr_i[0]_pad  & ~n14331 ;
  assign n33217 = n14339 & n33216 ;
  assign n33218 = \m4_addr_i[0]_pad  & n14331 ;
  assign n33219 = n14356 & n33218 ;
  assign n33220 = ~n33217 & ~n33219 ;
  assign n33221 = \m6_addr_i[0]_pad  & n14331 ;
  assign n33222 = n14348 & n33221 ;
  assign n33223 = \m2_addr_i[0]_pad  & n14331 ;
  assign n33224 = n14339 & n33223 ;
  assign n33225 = ~n33222 & ~n33224 ;
  assign n33226 = n33220 & n33225 ;
  assign n33227 = \m5_addr_i[0]_pad  & ~n14331 ;
  assign n33228 = n14356 & n33227 ;
  assign n33229 = \m1_addr_i[0]_pad  & ~n14331 ;
  assign n33230 = n14324 & n33229 ;
  assign n33231 = ~n33228 & ~n33230 ;
  assign n33232 = \m0_addr_i[0]_pad  & n14331 ;
  assign n33233 = n14324 & n33232 ;
  assign n33234 = \m7_addr_i[0]_pad  & ~n14331 ;
  assign n33235 = n14348 & n33234 ;
  assign n33236 = ~n33233 & ~n33235 ;
  assign n33237 = n33231 & n33236 ;
  assign n33238 = n33226 & n33237 ;
  assign n33239 = \m1_addr_i[10]_pad  & ~n14331 ;
  assign n33240 = n14324 & n33239 ;
  assign n33241 = \m2_addr_i[10]_pad  & n14331 ;
  assign n33242 = n14339 & n33241 ;
  assign n33243 = ~n33240 & ~n33242 ;
  assign n33244 = \m6_addr_i[10]_pad  & n14331 ;
  assign n33245 = n14348 & n33244 ;
  assign n33246 = \m7_addr_i[10]_pad  & ~n14331 ;
  assign n33247 = n14348 & n33246 ;
  assign n33248 = ~n33245 & ~n33247 ;
  assign n33249 = n33243 & n33248 ;
  assign n33250 = \m5_addr_i[10]_pad  & ~n14331 ;
  assign n33251 = n14356 & n33250 ;
  assign n33252 = \m0_addr_i[10]_pad  & n14331 ;
  assign n33253 = n14324 & n33252 ;
  assign n33254 = ~n33251 & ~n33253 ;
  assign n33255 = \m3_addr_i[10]_pad  & ~n14331 ;
  assign n33256 = n14339 & n33255 ;
  assign n33257 = \m4_addr_i[10]_pad  & n14331 ;
  assign n33258 = n14356 & n33257 ;
  assign n33259 = ~n33256 & ~n33258 ;
  assign n33260 = n33254 & n33259 ;
  assign n33261 = n33249 & n33260 ;
  assign n33262 = \m3_addr_i[11]_pad  & ~n14331 ;
  assign n33263 = n14339 & n33262 ;
  assign n33264 = \m4_addr_i[11]_pad  & n14331 ;
  assign n33265 = n14356 & n33264 ;
  assign n33266 = ~n33263 & ~n33265 ;
  assign n33267 = \m6_addr_i[11]_pad  & n14331 ;
  assign n33268 = n14348 & n33267 ;
  assign n33269 = \m2_addr_i[11]_pad  & n14331 ;
  assign n33270 = n14339 & n33269 ;
  assign n33271 = ~n33268 & ~n33270 ;
  assign n33272 = n33266 & n33271 ;
  assign n33273 = \m5_addr_i[11]_pad  & ~n14331 ;
  assign n33274 = n14356 & n33273 ;
  assign n33275 = \m1_addr_i[11]_pad  & ~n14331 ;
  assign n33276 = n14324 & n33275 ;
  assign n33277 = ~n33274 & ~n33276 ;
  assign n33278 = \m0_addr_i[11]_pad  & n14331 ;
  assign n33279 = n14324 & n33278 ;
  assign n33280 = \m7_addr_i[11]_pad  & ~n14331 ;
  assign n33281 = n14348 & n33280 ;
  assign n33282 = ~n33279 & ~n33281 ;
  assign n33283 = n33277 & n33282 ;
  assign n33284 = n33272 & n33283 ;
  assign n33285 = \m3_addr_i[12]_pad  & ~n14331 ;
  assign n33286 = n14339 & n33285 ;
  assign n33287 = \m4_addr_i[12]_pad  & n14331 ;
  assign n33288 = n14356 & n33287 ;
  assign n33289 = ~n33286 & ~n33288 ;
  assign n33290 = \m6_addr_i[12]_pad  & n14331 ;
  assign n33291 = n14348 & n33290 ;
  assign n33292 = \m2_addr_i[12]_pad  & n14331 ;
  assign n33293 = n14339 & n33292 ;
  assign n33294 = ~n33291 & ~n33293 ;
  assign n33295 = n33289 & n33294 ;
  assign n33296 = \m5_addr_i[12]_pad  & ~n14331 ;
  assign n33297 = n14356 & n33296 ;
  assign n33298 = \m1_addr_i[12]_pad  & ~n14331 ;
  assign n33299 = n14324 & n33298 ;
  assign n33300 = ~n33297 & ~n33299 ;
  assign n33301 = \m0_addr_i[12]_pad  & n14331 ;
  assign n33302 = n14324 & n33301 ;
  assign n33303 = \m7_addr_i[12]_pad  & ~n14331 ;
  assign n33304 = n14348 & n33303 ;
  assign n33305 = ~n33302 & ~n33304 ;
  assign n33306 = n33300 & n33305 ;
  assign n33307 = n33295 & n33306 ;
  assign n33308 = \m3_addr_i[13]_pad  & ~n14331 ;
  assign n33309 = n14339 & n33308 ;
  assign n33310 = \m4_addr_i[13]_pad  & n14331 ;
  assign n33311 = n14356 & n33310 ;
  assign n33312 = ~n33309 & ~n33311 ;
  assign n33313 = \m6_addr_i[13]_pad  & n14331 ;
  assign n33314 = n14348 & n33313 ;
  assign n33315 = \m2_addr_i[13]_pad  & n14331 ;
  assign n33316 = n14339 & n33315 ;
  assign n33317 = ~n33314 & ~n33316 ;
  assign n33318 = n33312 & n33317 ;
  assign n33319 = \m5_addr_i[13]_pad  & ~n14331 ;
  assign n33320 = n14356 & n33319 ;
  assign n33321 = \m1_addr_i[13]_pad  & ~n14331 ;
  assign n33322 = n14324 & n33321 ;
  assign n33323 = ~n33320 & ~n33322 ;
  assign n33324 = \m0_addr_i[13]_pad  & n14331 ;
  assign n33325 = n14324 & n33324 ;
  assign n33326 = \m7_addr_i[13]_pad  & ~n14331 ;
  assign n33327 = n14348 & n33326 ;
  assign n33328 = ~n33325 & ~n33327 ;
  assign n33329 = n33323 & n33328 ;
  assign n33330 = n33318 & n33329 ;
  assign n33331 = \m1_addr_i[14]_pad  & ~n14331 ;
  assign n33332 = n14324 & n33331 ;
  assign n33333 = \m2_addr_i[14]_pad  & n14331 ;
  assign n33334 = n14339 & n33333 ;
  assign n33335 = ~n33332 & ~n33334 ;
  assign n33336 = \m6_addr_i[14]_pad  & n14331 ;
  assign n33337 = n14348 & n33336 ;
  assign n33338 = \m7_addr_i[14]_pad  & ~n14331 ;
  assign n33339 = n14348 & n33338 ;
  assign n33340 = ~n33337 & ~n33339 ;
  assign n33341 = n33335 & n33340 ;
  assign n33342 = \m5_addr_i[14]_pad  & ~n14331 ;
  assign n33343 = n14356 & n33342 ;
  assign n33344 = \m0_addr_i[14]_pad  & n14331 ;
  assign n33345 = n14324 & n33344 ;
  assign n33346 = ~n33343 & ~n33345 ;
  assign n33347 = \m3_addr_i[14]_pad  & ~n14331 ;
  assign n33348 = n14339 & n33347 ;
  assign n33349 = \m4_addr_i[14]_pad  & n14331 ;
  assign n33350 = n14356 & n33349 ;
  assign n33351 = ~n33348 & ~n33350 ;
  assign n33352 = n33346 & n33351 ;
  assign n33353 = n33341 & n33352 ;
  assign n33354 = \m6_addr_i[15]_pad  & n14331 ;
  assign n33355 = n14348 & n33354 ;
  assign n33356 = \m5_addr_i[15]_pad  & ~n14331 ;
  assign n33357 = n14356 & n33356 ;
  assign n33358 = ~n33355 & ~n33357 ;
  assign n33359 = \m0_addr_i[15]_pad  & n14331 ;
  assign n33360 = n14324 & n33359 ;
  assign n33361 = \m4_addr_i[15]_pad  & n14331 ;
  assign n33362 = n14356 & n33361 ;
  assign n33363 = ~n33360 & ~n33362 ;
  assign n33364 = n33358 & n33363 ;
  assign n33365 = \m7_addr_i[15]_pad  & ~n14331 ;
  assign n33366 = n14348 & n33365 ;
  assign n33367 = \m3_addr_i[15]_pad  & ~n14331 ;
  assign n33368 = n14339 & n33367 ;
  assign n33369 = ~n33366 & ~n33368 ;
  assign n33370 = \m1_addr_i[15]_pad  & ~n14331 ;
  assign n33371 = n14324 & n33370 ;
  assign n33372 = \m2_addr_i[15]_pad  & n14331 ;
  assign n33373 = n14339 & n33372 ;
  assign n33374 = ~n33371 & ~n33373 ;
  assign n33375 = n33369 & n33374 ;
  assign n33376 = n33364 & n33375 ;
  assign n33377 = \m3_addr_i[16]_pad  & ~n14331 ;
  assign n33378 = n14339 & n33377 ;
  assign n33379 = \m4_addr_i[16]_pad  & n14331 ;
  assign n33380 = n14356 & n33379 ;
  assign n33381 = ~n33378 & ~n33380 ;
  assign n33382 = \m6_addr_i[16]_pad  & n14331 ;
  assign n33383 = n14348 & n33382 ;
  assign n33384 = \m7_addr_i[16]_pad  & ~n14331 ;
  assign n33385 = n14348 & n33384 ;
  assign n33386 = ~n33383 & ~n33385 ;
  assign n33387 = n33381 & n33386 ;
  assign n33388 = \m5_addr_i[16]_pad  & ~n14331 ;
  assign n33389 = n14356 & n33388 ;
  assign n33390 = \m0_addr_i[16]_pad  & n14331 ;
  assign n33391 = n14324 & n33390 ;
  assign n33392 = ~n33389 & ~n33391 ;
  assign n33393 = \m1_addr_i[16]_pad  & ~n14331 ;
  assign n33394 = n14324 & n33393 ;
  assign n33395 = \m2_addr_i[16]_pad  & n14331 ;
  assign n33396 = n14339 & n33395 ;
  assign n33397 = ~n33394 & ~n33396 ;
  assign n33398 = n33392 & n33397 ;
  assign n33399 = n33387 & n33398 ;
  assign n33400 = \m3_addr_i[17]_pad  & ~n14331 ;
  assign n33401 = n14339 & n33400 ;
  assign n33402 = \m4_addr_i[17]_pad  & n14331 ;
  assign n33403 = n14356 & n33402 ;
  assign n33404 = ~n33401 & ~n33403 ;
  assign n33405 = \m6_addr_i[17]_pad  & n14331 ;
  assign n33406 = n14348 & n33405 ;
  assign n33407 = \m2_addr_i[17]_pad  & n14331 ;
  assign n33408 = n14339 & n33407 ;
  assign n33409 = ~n33406 & ~n33408 ;
  assign n33410 = n33404 & n33409 ;
  assign n33411 = \m5_addr_i[17]_pad  & ~n14331 ;
  assign n33412 = n14356 & n33411 ;
  assign n33413 = \m1_addr_i[17]_pad  & ~n14331 ;
  assign n33414 = n14324 & n33413 ;
  assign n33415 = ~n33412 & ~n33414 ;
  assign n33416 = \m0_addr_i[17]_pad  & n14331 ;
  assign n33417 = n14324 & n33416 ;
  assign n33418 = \m7_addr_i[17]_pad  & ~n14331 ;
  assign n33419 = n14348 & n33418 ;
  assign n33420 = ~n33417 & ~n33419 ;
  assign n33421 = n33415 & n33420 ;
  assign n33422 = n33410 & n33421 ;
  assign n33423 = \m3_addr_i[18]_pad  & ~n14331 ;
  assign n33424 = n14339 & n33423 ;
  assign n33425 = \m4_addr_i[18]_pad  & n14331 ;
  assign n33426 = n14356 & n33425 ;
  assign n33427 = ~n33424 & ~n33426 ;
  assign n33428 = \m6_addr_i[18]_pad  & n14331 ;
  assign n33429 = n14348 & n33428 ;
  assign n33430 = \m7_addr_i[18]_pad  & ~n14331 ;
  assign n33431 = n14348 & n33430 ;
  assign n33432 = ~n33429 & ~n33431 ;
  assign n33433 = n33427 & n33432 ;
  assign n33434 = \m5_addr_i[18]_pad  & ~n14331 ;
  assign n33435 = n14356 & n33434 ;
  assign n33436 = \m0_addr_i[18]_pad  & n14331 ;
  assign n33437 = n14324 & n33436 ;
  assign n33438 = ~n33435 & ~n33437 ;
  assign n33439 = \m1_addr_i[18]_pad  & ~n14331 ;
  assign n33440 = n14324 & n33439 ;
  assign n33441 = \m2_addr_i[18]_pad  & n14331 ;
  assign n33442 = n14339 & n33441 ;
  assign n33443 = ~n33440 & ~n33442 ;
  assign n33444 = n33438 & n33443 ;
  assign n33445 = n33433 & n33444 ;
  assign n33446 = \m3_addr_i[19]_pad  & ~n14331 ;
  assign n33447 = n14339 & n33446 ;
  assign n33448 = \m4_addr_i[19]_pad  & n14331 ;
  assign n33449 = n14356 & n33448 ;
  assign n33450 = ~n33447 & ~n33449 ;
  assign n33451 = \m6_addr_i[19]_pad  & n14331 ;
  assign n33452 = n14348 & n33451 ;
  assign n33453 = \m2_addr_i[19]_pad  & n14331 ;
  assign n33454 = n14339 & n33453 ;
  assign n33455 = ~n33452 & ~n33454 ;
  assign n33456 = n33450 & n33455 ;
  assign n33457 = \m5_addr_i[19]_pad  & ~n14331 ;
  assign n33458 = n14356 & n33457 ;
  assign n33459 = \m1_addr_i[19]_pad  & ~n14331 ;
  assign n33460 = n14324 & n33459 ;
  assign n33461 = ~n33458 & ~n33460 ;
  assign n33462 = \m0_addr_i[19]_pad  & n14331 ;
  assign n33463 = n14324 & n33462 ;
  assign n33464 = \m7_addr_i[19]_pad  & ~n14331 ;
  assign n33465 = n14348 & n33464 ;
  assign n33466 = ~n33463 & ~n33465 ;
  assign n33467 = n33461 & n33466 ;
  assign n33468 = n33456 & n33467 ;
  assign n33469 = \m3_addr_i[1]_pad  & ~n14331 ;
  assign n33470 = n14339 & n33469 ;
  assign n33471 = \m4_addr_i[1]_pad  & n14331 ;
  assign n33472 = n14356 & n33471 ;
  assign n33473 = ~n33470 & ~n33472 ;
  assign n33474 = \m6_addr_i[1]_pad  & n14331 ;
  assign n33475 = n14348 & n33474 ;
  assign n33476 = \m2_addr_i[1]_pad  & n14331 ;
  assign n33477 = n14339 & n33476 ;
  assign n33478 = ~n33475 & ~n33477 ;
  assign n33479 = n33473 & n33478 ;
  assign n33480 = \m5_addr_i[1]_pad  & ~n14331 ;
  assign n33481 = n14356 & n33480 ;
  assign n33482 = \m1_addr_i[1]_pad  & ~n14331 ;
  assign n33483 = n14324 & n33482 ;
  assign n33484 = ~n33481 & ~n33483 ;
  assign n33485 = \m0_addr_i[1]_pad  & n14331 ;
  assign n33486 = n14324 & n33485 ;
  assign n33487 = \m7_addr_i[1]_pad  & ~n14331 ;
  assign n33488 = n14348 & n33487 ;
  assign n33489 = ~n33486 & ~n33488 ;
  assign n33490 = n33484 & n33489 ;
  assign n33491 = n33479 & n33490 ;
  assign n33492 = \m3_addr_i[20]_pad  & ~n14331 ;
  assign n33493 = n14339 & n33492 ;
  assign n33494 = \m4_addr_i[20]_pad  & n14331 ;
  assign n33495 = n14356 & n33494 ;
  assign n33496 = ~n33493 & ~n33495 ;
  assign n33497 = \m6_addr_i[20]_pad  & n14331 ;
  assign n33498 = n14348 & n33497 ;
  assign n33499 = \m2_addr_i[20]_pad  & n14331 ;
  assign n33500 = n14339 & n33499 ;
  assign n33501 = ~n33498 & ~n33500 ;
  assign n33502 = n33496 & n33501 ;
  assign n33503 = \m5_addr_i[20]_pad  & ~n14331 ;
  assign n33504 = n14356 & n33503 ;
  assign n33505 = \m1_addr_i[20]_pad  & ~n14331 ;
  assign n33506 = n14324 & n33505 ;
  assign n33507 = ~n33504 & ~n33506 ;
  assign n33508 = \m0_addr_i[20]_pad  & n14331 ;
  assign n33509 = n14324 & n33508 ;
  assign n33510 = \m7_addr_i[20]_pad  & ~n14331 ;
  assign n33511 = n14348 & n33510 ;
  assign n33512 = ~n33509 & ~n33511 ;
  assign n33513 = n33507 & n33512 ;
  assign n33514 = n33502 & n33513 ;
  assign n33515 = \m3_addr_i[21]_pad  & ~n14331 ;
  assign n33516 = n14339 & n33515 ;
  assign n33517 = \m4_addr_i[21]_pad  & n14331 ;
  assign n33518 = n14356 & n33517 ;
  assign n33519 = ~n33516 & ~n33518 ;
  assign n33520 = \m6_addr_i[21]_pad  & n14331 ;
  assign n33521 = n14348 & n33520 ;
  assign n33522 = \m2_addr_i[21]_pad  & n14331 ;
  assign n33523 = n14339 & n33522 ;
  assign n33524 = ~n33521 & ~n33523 ;
  assign n33525 = n33519 & n33524 ;
  assign n33526 = \m5_addr_i[21]_pad  & ~n14331 ;
  assign n33527 = n14356 & n33526 ;
  assign n33528 = \m1_addr_i[21]_pad  & ~n14331 ;
  assign n33529 = n14324 & n33528 ;
  assign n33530 = ~n33527 & ~n33529 ;
  assign n33531 = \m0_addr_i[21]_pad  & n14331 ;
  assign n33532 = n14324 & n33531 ;
  assign n33533 = \m7_addr_i[21]_pad  & ~n14331 ;
  assign n33534 = n14348 & n33533 ;
  assign n33535 = ~n33532 & ~n33534 ;
  assign n33536 = n33530 & n33535 ;
  assign n33537 = n33525 & n33536 ;
  assign n33538 = \m3_addr_i[22]_pad  & ~n14331 ;
  assign n33539 = n14339 & n33538 ;
  assign n33540 = \m4_addr_i[22]_pad  & n14331 ;
  assign n33541 = n14356 & n33540 ;
  assign n33542 = ~n33539 & ~n33541 ;
  assign n33543 = \m6_addr_i[22]_pad  & n14331 ;
  assign n33544 = n14348 & n33543 ;
  assign n33545 = \m2_addr_i[22]_pad  & n14331 ;
  assign n33546 = n14339 & n33545 ;
  assign n33547 = ~n33544 & ~n33546 ;
  assign n33548 = n33542 & n33547 ;
  assign n33549 = \m5_addr_i[22]_pad  & ~n14331 ;
  assign n33550 = n14356 & n33549 ;
  assign n33551 = \m1_addr_i[22]_pad  & ~n14331 ;
  assign n33552 = n14324 & n33551 ;
  assign n33553 = ~n33550 & ~n33552 ;
  assign n33554 = \m0_addr_i[22]_pad  & n14331 ;
  assign n33555 = n14324 & n33554 ;
  assign n33556 = \m7_addr_i[22]_pad  & ~n14331 ;
  assign n33557 = n14348 & n33556 ;
  assign n33558 = ~n33555 & ~n33557 ;
  assign n33559 = n33553 & n33558 ;
  assign n33560 = n33548 & n33559 ;
  assign n33561 = \m3_addr_i[23]_pad  & ~n14331 ;
  assign n33562 = n14339 & n33561 ;
  assign n33563 = \m4_addr_i[23]_pad  & n14331 ;
  assign n33564 = n14356 & n33563 ;
  assign n33565 = ~n33562 & ~n33564 ;
  assign n33566 = \m6_addr_i[23]_pad  & n14331 ;
  assign n33567 = n14348 & n33566 ;
  assign n33568 = \m2_addr_i[23]_pad  & n14331 ;
  assign n33569 = n14339 & n33568 ;
  assign n33570 = ~n33567 & ~n33569 ;
  assign n33571 = n33565 & n33570 ;
  assign n33572 = \m5_addr_i[23]_pad  & ~n14331 ;
  assign n33573 = n14356 & n33572 ;
  assign n33574 = \m1_addr_i[23]_pad  & ~n14331 ;
  assign n33575 = n14324 & n33574 ;
  assign n33576 = ~n33573 & ~n33575 ;
  assign n33577 = \m0_addr_i[23]_pad  & n14331 ;
  assign n33578 = n14324 & n33577 ;
  assign n33579 = \m7_addr_i[23]_pad  & ~n14331 ;
  assign n33580 = n14348 & n33579 ;
  assign n33581 = ~n33578 & ~n33580 ;
  assign n33582 = n33576 & n33581 ;
  assign n33583 = n33571 & n33582 ;
  assign n33584 = \m3_addr_i[24]_pad  & ~n14331 ;
  assign n33585 = n14339 & n33584 ;
  assign n33586 = \m4_addr_i[24]_pad  & n14331 ;
  assign n33587 = n14356 & n33586 ;
  assign n33588 = ~n33585 & ~n33587 ;
  assign n33589 = \m5_addr_i[24]_pad  & ~n14331 ;
  assign n33590 = n14356 & n33589 ;
  assign n33591 = \m2_addr_i[24]_pad  & n14331 ;
  assign n33592 = n14339 & n33591 ;
  assign n33593 = ~n33590 & ~n33592 ;
  assign n33594 = n33588 & n33593 ;
  assign n33595 = \m6_addr_i[24]_pad  & n14331 ;
  assign n33596 = n14348 & n33595 ;
  assign n33597 = \m1_addr_i[24]_pad  & ~n14331 ;
  assign n33598 = n14324 & n33597 ;
  assign n33599 = ~n33596 & ~n33598 ;
  assign n33600 = \m0_addr_i[24]_pad  & n14331 ;
  assign n33601 = n14324 & n33600 ;
  assign n33602 = \m7_addr_i[24]_pad  & ~n14331 ;
  assign n33603 = n14348 & n33602 ;
  assign n33604 = ~n33601 & ~n33603 ;
  assign n33605 = n33599 & n33604 ;
  assign n33606 = n33594 & n33605 ;
  assign n33607 = \m3_addr_i[25]_pad  & ~n14331 ;
  assign n33608 = n14339 & n33607 ;
  assign n33609 = \m4_addr_i[25]_pad  & n14331 ;
  assign n33610 = n14356 & n33609 ;
  assign n33611 = ~n33608 & ~n33610 ;
  assign n33612 = \m5_addr_i[25]_pad  & ~n14331 ;
  assign n33613 = n14356 & n33612 ;
  assign n33614 = \m2_addr_i[25]_pad  & n14331 ;
  assign n33615 = n14339 & n33614 ;
  assign n33616 = ~n33613 & ~n33615 ;
  assign n33617 = n33611 & n33616 ;
  assign n33618 = \m6_addr_i[25]_pad  & n14331 ;
  assign n33619 = n14348 & n33618 ;
  assign n33620 = \m1_addr_i[25]_pad  & ~n14331 ;
  assign n33621 = n14324 & n33620 ;
  assign n33622 = ~n33619 & ~n33621 ;
  assign n33623 = \m0_addr_i[25]_pad  & n14331 ;
  assign n33624 = n14324 & n33623 ;
  assign n33625 = \m7_addr_i[25]_pad  & ~n14331 ;
  assign n33626 = n14348 & n33625 ;
  assign n33627 = ~n33624 & ~n33626 ;
  assign n33628 = n33622 & n33627 ;
  assign n33629 = n33617 & n33628 ;
  assign n33630 = \m3_addr_i[26]_pad  & ~n14331 ;
  assign n33631 = n14339 & n33630 ;
  assign n33632 = \m4_addr_i[26]_pad  & n14331 ;
  assign n33633 = n14356 & n33632 ;
  assign n33634 = ~n33631 & ~n33633 ;
  assign n33635 = \m5_addr_i[26]_pad  & ~n14331 ;
  assign n33636 = n14356 & n33635 ;
  assign n33637 = \m2_addr_i[26]_pad  & n14331 ;
  assign n33638 = n14339 & n33637 ;
  assign n33639 = ~n33636 & ~n33638 ;
  assign n33640 = n33634 & n33639 ;
  assign n33641 = \m6_addr_i[26]_pad  & n14331 ;
  assign n33642 = n14348 & n33641 ;
  assign n33643 = \m1_addr_i[26]_pad  & ~n14331 ;
  assign n33644 = n14324 & n33643 ;
  assign n33645 = ~n33642 & ~n33644 ;
  assign n33646 = \m0_addr_i[26]_pad  & n14331 ;
  assign n33647 = n14324 & n33646 ;
  assign n33648 = \m7_addr_i[26]_pad  & ~n14331 ;
  assign n33649 = n14348 & n33648 ;
  assign n33650 = ~n33647 & ~n33649 ;
  assign n33651 = n33645 & n33650 ;
  assign n33652 = n33640 & n33651 ;
  assign n33653 = \m3_addr_i[27]_pad  & ~n14331 ;
  assign n33654 = n14339 & n33653 ;
  assign n33655 = \m4_addr_i[27]_pad  & n14331 ;
  assign n33656 = n14356 & n33655 ;
  assign n33657 = ~n33654 & ~n33656 ;
  assign n33658 = \m5_addr_i[27]_pad  & ~n14331 ;
  assign n33659 = n14356 & n33658 ;
  assign n33660 = \m2_addr_i[27]_pad  & n14331 ;
  assign n33661 = n14339 & n33660 ;
  assign n33662 = ~n33659 & ~n33661 ;
  assign n33663 = n33657 & n33662 ;
  assign n33664 = \m6_addr_i[27]_pad  & n14331 ;
  assign n33665 = n14348 & n33664 ;
  assign n33666 = \m1_addr_i[27]_pad  & ~n14331 ;
  assign n33667 = n14324 & n33666 ;
  assign n33668 = ~n33665 & ~n33667 ;
  assign n33669 = \m0_addr_i[27]_pad  & n14331 ;
  assign n33670 = n14324 & n33669 ;
  assign n33671 = \m7_addr_i[27]_pad  & ~n14331 ;
  assign n33672 = n14348 & n33671 ;
  assign n33673 = ~n33670 & ~n33672 ;
  assign n33674 = n33668 & n33673 ;
  assign n33675 = n33663 & n33674 ;
  assign n33676 = \m3_addr_i[28]_pad  & ~n14331 ;
  assign n33677 = n14339 & n33676 ;
  assign n33678 = \m4_addr_i[28]_pad  & n14331 ;
  assign n33679 = n14356 & n33678 ;
  assign n33680 = ~n33677 & ~n33679 ;
  assign n33681 = \m5_addr_i[28]_pad  & ~n14331 ;
  assign n33682 = n14356 & n33681 ;
  assign n33683 = \m2_addr_i[28]_pad  & n14331 ;
  assign n33684 = n14339 & n33683 ;
  assign n33685 = ~n33682 & ~n33684 ;
  assign n33686 = n33680 & n33685 ;
  assign n33687 = \m6_addr_i[28]_pad  & n14331 ;
  assign n33688 = n14348 & n33687 ;
  assign n33689 = \m1_addr_i[28]_pad  & ~n14331 ;
  assign n33690 = n14324 & n33689 ;
  assign n33691 = ~n33688 & ~n33690 ;
  assign n33692 = \m0_addr_i[28]_pad  & n14331 ;
  assign n33693 = n14324 & n33692 ;
  assign n33694 = \m7_addr_i[28]_pad  & ~n14331 ;
  assign n33695 = n14348 & n33694 ;
  assign n33696 = ~n33693 & ~n33695 ;
  assign n33697 = n33691 & n33696 ;
  assign n33698 = n33686 & n33697 ;
  assign n33699 = \m3_addr_i[29]_pad  & ~n14331 ;
  assign n33700 = n14339 & n33699 ;
  assign n33701 = \m4_addr_i[29]_pad  & n14331 ;
  assign n33702 = n14356 & n33701 ;
  assign n33703 = ~n33700 & ~n33702 ;
  assign n33704 = \m5_addr_i[29]_pad  & ~n14331 ;
  assign n33705 = n14356 & n33704 ;
  assign n33706 = \m2_addr_i[29]_pad  & n14331 ;
  assign n33707 = n14339 & n33706 ;
  assign n33708 = ~n33705 & ~n33707 ;
  assign n33709 = n33703 & n33708 ;
  assign n33710 = \m6_addr_i[29]_pad  & n14331 ;
  assign n33711 = n14348 & n33710 ;
  assign n33712 = \m1_addr_i[29]_pad  & ~n14331 ;
  assign n33713 = n14324 & n33712 ;
  assign n33714 = ~n33711 & ~n33713 ;
  assign n33715 = \m0_addr_i[29]_pad  & n14331 ;
  assign n33716 = n14324 & n33715 ;
  assign n33717 = \m7_addr_i[29]_pad  & ~n14331 ;
  assign n33718 = n14348 & n33717 ;
  assign n33719 = ~n33716 & ~n33718 ;
  assign n33720 = n33714 & n33719 ;
  assign n33721 = n33709 & n33720 ;
  assign n33722 = \m6_addr_i[2]_pad  & n14331 ;
  assign n33723 = n14348 & n33722 ;
  assign n33724 = \m5_addr_i[2]_pad  & ~n14331 ;
  assign n33725 = n14356 & n33724 ;
  assign n33726 = ~n33723 & ~n33725 ;
  assign n33727 = \m0_addr_i[2]_pad  & n14331 ;
  assign n33728 = n14324 & n33727 ;
  assign n33729 = \m4_addr_i[2]_pad  & n14331 ;
  assign n33730 = n14356 & n33729 ;
  assign n33731 = ~n33728 & ~n33730 ;
  assign n33732 = n33726 & n33731 ;
  assign n33733 = \m7_addr_i[2]_pad  & ~n14331 ;
  assign n33734 = n14348 & n33733 ;
  assign n33735 = \m3_addr_i[2]_pad  & ~n14331 ;
  assign n33736 = n14339 & n33735 ;
  assign n33737 = ~n33734 & ~n33736 ;
  assign n33738 = \m1_addr_i[2]_pad  & ~n14331 ;
  assign n33739 = n14324 & n33738 ;
  assign n33740 = \m2_addr_i[2]_pad  & n14331 ;
  assign n33741 = n14339 & n33740 ;
  assign n33742 = ~n33739 & ~n33741 ;
  assign n33743 = n33737 & n33742 ;
  assign n33744 = n33732 & n33743 ;
  assign n33745 = \m3_addr_i[30]_pad  & ~n14331 ;
  assign n33746 = n14339 & n33745 ;
  assign n33747 = \m4_addr_i[30]_pad  & n14331 ;
  assign n33748 = n14356 & n33747 ;
  assign n33749 = ~n33746 & ~n33748 ;
  assign n33750 = \m5_addr_i[30]_pad  & ~n14331 ;
  assign n33751 = n14356 & n33750 ;
  assign n33752 = \m2_addr_i[30]_pad  & n14331 ;
  assign n33753 = n14339 & n33752 ;
  assign n33754 = ~n33751 & ~n33753 ;
  assign n33755 = n33749 & n33754 ;
  assign n33756 = \m6_addr_i[30]_pad  & n14331 ;
  assign n33757 = n14348 & n33756 ;
  assign n33758 = \m1_addr_i[30]_pad  & ~n14331 ;
  assign n33759 = n14324 & n33758 ;
  assign n33760 = ~n33757 & ~n33759 ;
  assign n33761 = \m0_addr_i[30]_pad  & n14331 ;
  assign n33762 = n14324 & n33761 ;
  assign n33763 = \m7_addr_i[30]_pad  & ~n14331 ;
  assign n33764 = n14348 & n33763 ;
  assign n33765 = ~n33762 & ~n33764 ;
  assign n33766 = n33760 & n33765 ;
  assign n33767 = n33755 & n33766 ;
  assign n33768 = \m3_addr_i[31]_pad  & ~n14331 ;
  assign n33769 = n14339 & n33768 ;
  assign n33770 = \m4_addr_i[31]_pad  & n14331 ;
  assign n33771 = n14356 & n33770 ;
  assign n33772 = ~n33769 & ~n33771 ;
  assign n33773 = \m5_addr_i[31]_pad  & ~n14331 ;
  assign n33774 = n14356 & n33773 ;
  assign n33775 = \m2_addr_i[31]_pad  & n14331 ;
  assign n33776 = n14339 & n33775 ;
  assign n33777 = ~n33774 & ~n33776 ;
  assign n33778 = n33772 & n33777 ;
  assign n33779 = \m6_addr_i[31]_pad  & n14331 ;
  assign n33780 = n14348 & n33779 ;
  assign n33781 = \m1_addr_i[31]_pad  & ~n14331 ;
  assign n33782 = n14324 & n33781 ;
  assign n33783 = ~n33780 & ~n33782 ;
  assign n33784 = \m0_addr_i[31]_pad  & n14331 ;
  assign n33785 = n14324 & n33784 ;
  assign n33786 = \m7_addr_i[31]_pad  & ~n14331 ;
  assign n33787 = n14348 & n33786 ;
  assign n33788 = ~n33785 & ~n33787 ;
  assign n33789 = n33783 & n33788 ;
  assign n33790 = n33778 & n33789 ;
  assign n33791 = \m3_addr_i[3]_pad  & ~n14331 ;
  assign n33792 = n14339 & n33791 ;
  assign n33793 = \m4_addr_i[3]_pad  & n14331 ;
  assign n33794 = n14356 & n33793 ;
  assign n33795 = ~n33792 & ~n33794 ;
  assign n33796 = \m6_addr_i[3]_pad  & n14331 ;
  assign n33797 = n14348 & n33796 ;
  assign n33798 = \m2_addr_i[3]_pad  & n14331 ;
  assign n33799 = n14339 & n33798 ;
  assign n33800 = ~n33797 & ~n33799 ;
  assign n33801 = n33795 & n33800 ;
  assign n33802 = \m5_addr_i[3]_pad  & ~n14331 ;
  assign n33803 = n14356 & n33802 ;
  assign n33804 = \m1_addr_i[3]_pad  & ~n14331 ;
  assign n33805 = n14324 & n33804 ;
  assign n33806 = ~n33803 & ~n33805 ;
  assign n33807 = \m0_addr_i[3]_pad  & n14331 ;
  assign n33808 = n14324 & n33807 ;
  assign n33809 = \m7_addr_i[3]_pad  & ~n14331 ;
  assign n33810 = n14348 & n33809 ;
  assign n33811 = ~n33808 & ~n33810 ;
  assign n33812 = n33806 & n33811 ;
  assign n33813 = n33801 & n33812 ;
  assign n33814 = \m6_addr_i[4]_pad  & n14331 ;
  assign n33815 = n14348 & n33814 ;
  assign n33816 = \m5_addr_i[4]_pad  & ~n14331 ;
  assign n33817 = n14356 & n33816 ;
  assign n33818 = ~n33815 & ~n33817 ;
  assign n33819 = \m0_addr_i[4]_pad  & n14331 ;
  assign n33820 = n14324 & n33819 ;
  assign n33821 = \m4_addr_i[4]_pad  & n14331 ;
  assign n33822 = n14356 & n33821 ;
  assign n33823 = ~n33820 & ~n33822 ;
  assign n33824 = n33818 & n33823 ;
  assign n33825 = \m7_addr_i[4]_pad  & ~n14331 ;
  assign n33826 = n14348 & n33825 ;
  assign n33827 = \m3_addr_i[4]_pad  & ~n14331 ;
  assign n33828 = n14339 & n33827 ;
  assign n33829 = ~n33826 & ~n33828 ;
  assign n33830 = \m1_addr_i[4]_pad  & ~n14331 ;
  assign n33831 = n14324 & n33830 ;
  assign n33832 = \m2_addr_i[4]_pad  & n14331 ;
  assign n33833 = n14339 & n33832 ;
  assign n33834 = ~n33831 & ~n33833 ;
  assign n33835 = n33829 & n33834 ;
  assign n33836 = n33824 & n33835 ;
  assign n33837 = \m3_addr_i[5]_pad  & ~n14331 ;
  assign n33838 = n14339 & n33837 ;
  assign n33839 = \m4_addr_i[5]_pad  & n14331 ;
  assign n33840 = n14356 & n33839 ;
  assign n33841 = ~n33838 & ~n33840 ;
  assign n33842 = \m6_addr_i[5]_pad  & n14331 ;
  assign n33843 = n14348 & n33842 ;
  assign n33844 = \m2_addr_i[5]_pad  & n14331 ;
  assign n33845 = n14339 & n33844 ;
  assign n33846 = ~n33843 & ~n33845 ;
  assign n33847 = n33841 & n33846 ;
  assign n33848 = \m5_addr_i[5]_pad  & ~n14331 ;
  assign n33849 = n14356 & n33848 ;
  assign n33850 = \m1_addr_i[5]_pad  & ~n14331 ;
  assign n33851 = n14324 & n33850 ;
  assign n33852 = ~n33849 & ~n33851 ;
  assign n33853 = \m0_addr_i[5]_pad  & n14331 ;
  assign n33854 = n14324 & n33853 ;
  assign n33855 = \m7_addr_i[5]_pad  & ~n14331 ;
  assign n33856 = n14348 & n33855 ;
  assign n33857 = ~n33854 & ~n33856 ;
  assign n33858 = n33852 & n33857 ;
  assign n33859 = n33847 & n33858 ;
  assign n33860 = \m3_addr_i[6]_pad  & ~n14331 ;
  assign n33861 = n14339 & n33860 ;
  assign n33862 = \m4_addr_i[6]_pad  & n14331 ;
  assign n33863 = n14356 & n33862 ;
  assign n33864 = ~n33861 & ~n33863 ;
  assign n33865 = \m6_addr_i[6]_pad  & n14331 ;
  assign n33866 = n14348 & n33865 ;
  assign n33867 = \m2_addr_i[6]_pad  & n14331 ;
  assign n33868 = n14339 & n33867 ;
  assign n33869 = ~n33866 & ~n33868 ;
  assign n33870 = n33864 & n33869 ;
  assign n33871 = \m5_addr_i[6]_pad  & ~n14331 ;
  assign n33872 = n14356 & n33871 ;
  assign n33873 = \m1_addr_i[6]_pad  & ~n14331 ;
  assign n33874 = n14324 & n33873 ;
  assign n33875 = ~n33872 & ~n33874 ;
  assign n33876 = \m0_addr_i[6]_pad  & n14331 ;
  assign n33877 = n14324 & n33876 ;
  assign n33878 = \m7_addr_i[6]_pad  & ~n14331 ;
  assign n33879 = n14348 & n33878 ;
  assign n33880 = ~n33877 & ~n33879 ;
  assign n33881 = n33875 & n33880 ;
  assign n33882 = n33870 & n33881 ;
  assign n33883 = \m3_addr_i[7]_pad  & ~n14331 ;
  assign n33884 = n14339 & n33883 ;
  assign n33885 = \m4_addr_i[7]_pad  & n14331 ;
  assign n33886 = n14356 & n33885 ;
  assign n33887 = ~n33884 & ~n33886 ;
  assign n33888 = \m6_addr_i[7]_pad  & n14331 ;
  assign n33889 = n14348 & n33888 ;
  assign n33890 = \m2_addr_i[7]_pad  & n14331 ;
  assign n33891 = n14339 & n33890 ;
  assign n33892 = ~n33889 & ~n33891 ;
  assign n33893 = n33887 & n33892 ;
  assign n33894 = \m5_addr_i[7]_pad  & ~n14331 ;
  assign n33895 = n14356 & n33894 ;
  assign n33896 = \m1_addr_i[7]_pad  & ~n14331 ;
  assign n33897 = n14324 & n33896 ;
  assign n33898 = ~n33895 & ~n33897 ;
  assign n33899 = \m0_addr_i[7]_pad  & n14331 ;
  assign n33900 = n14324 & n33899 ;
  assign n33901 = \m7_addr_i[7]_pad  & ~n14331 ;
  assign n33902 = n14348 & n33901 ;
  assign n33903 = ~n33900 & ~n33902 ;
  assign n33904 = n33898 & n33903 ;
  assign n33905 = n33893 & n33904 ;
  assign n33906 = \m3_addr_i[8]_pad  & ~n14331 ;
  assign n33907 = n14339 & n33906 ;
  assign n33908 = \m4_addr_i[8]_pad  & n14331 ;
  assign n33909 = n14356 & n33908 ;
  assign n33910 = ~n33907 & ~n33909 ;
  assign n33911 = \m6_addr_i[8]_pad  & n14331 ;
  assign n33912 = n14348 & n33911 ;
  assign n33913 = \m2_addr_i[8]_pad  & n14331 ;
  assign n33914 = n14339 & n33913 ;
  assign n33915 = ~n33912 & ~n33914 ;
  assign n33916 = n33910 & n33915 ;
  assign n33917 = \m5_addr_i[8]_pad  & ~n14331 ;
  assign n33918 = n14356 & n33917 ;
  assign n33919 = \m1_addr_i[8]_pad  & ~n14331 ;
  assign n33920 = n14324 & n33919 ;
  assign n33921 = ~n33918 & ~n33920 ;
  assign n33922 = \m0_addr_i[8]_pad  & n14331 ;
  assign n33923 = n14324 & n33922 ;
  assign n33924 = \m7_addr_i[8]_pad  & ~n14331 ;
  assign n33925 = n14348 & n33924 ;
  assign n33926 = ~n33923 & ~n33925 ;
  assign n33927 = n33921 & n33926 ;
  assign n33928 = n33916 & n33927 ;
  assign n33929 = \m3_addr_i[9]_pad  & ~n14331 ;
  assign n33930 = n14339 & n33929 ;
  assign n33931 = \m4_addr_i[9]_pad  & n14331 ;
  assign n33932 = n14356 & n33931 ;
  assign n33933 = ~n33930 & ~n33932 ;
  assign n33934 = \m6_addr_i[9]_pad  & n14331 ;
  assign n33935 = n14348 & n33934 ;
  assign n33936 = \m2_addr_i[9]_pad  & n14331 ;
  assign n33937 = n14339 & n33936 ;
  assign n33938 = ~n33935 & ~n33937 ;
  assign n33939 = n33933 & n33938 ;
  assign n33940 = \m5_addr_i[9]_pad  & ~n14331 ;
  assign n33941 = n14356 & n33940 ;
  assign n33942 = \m1_addr_i[9]_pad  & ~n14331 ;
  assign n33943 = n14324 & n33942 ;
  assign n33944 = ~n33941 & ~n33943 ;
  assign n33945 = \m0_addr_i[9]_pad  & n14331 ;
  assign n33946 = n14324 & n33945 ;
  assign n33947 = \m7_addr_i[9]_pad  & ~n14331 ;
  assign n33948 = n14348 & n33947 ;
  assign n33949 = ~n33946 & ~n33948 ;
  assign n33950 = n33944 & n33949 ;
  assign n33951 = n33939 & n33950 ;
  assign n33952 = \m3_data_i[0]_pad  & ~n14331 ;
  assign n33953 = n14339 & n33952 ;
  assign n33954 = \m4_data_i[0]_pad  & n14331 ;
  assign n33955 = n14356 & n33954 ;
  assign n33956 = ~n33953 & ~n33955 ;
  assign n33957 = \m6_data_i[0]_pad  & n14331 ;
  assign n33958 = n14348 & n33957 ;
  assign n33959 = \m2_data_i[0]_pad  & n14331 ;
  assign n33960 = n14339 & n33959 ;
  assign n33961 = ~n33958 & ~n33960 ;
  assign n33962 = n33956 & n33961 ;
  assign n33963 = \m5_data_i[0]_pad  & ~n14331 ;
  assign n33964 = n14356 & n33963 ;
  assign n33965 = \m1_data_i[0]_pad  & ~n14331 ;
  assign n33966 = n14324 & n33965 ;
  assign n33967 = ~n33964 & ~n33966 ;
  assign n33968 = \m0_data_i[0]_pad  & n14331 ;
  assign n33969 = n14324 & n33968 ;
  assign n33970 = \m7_data_i[0]_pad  & ~n14331 ;
  assign n33971 = n14348 & n33970 ;
  assign n33972 = ~n33969 & ~n33971 ;
  assign n33973 = n33967 & n33972 ;
  assign n33974 = n33962 & n33973 ;
  assign n33975 = \m3_data_i[10]_pad  & ~n14331 ;
  assign n33976 = n14339 & n33975 ;
  assign n33977 = \m4_data_i[10]_pad  & n14331 ;
  assign n33978 = n14356 & n33977 ;
  assign n33979 = ~n33976 & ~n33978 ;
  assign n33980 = \m6_data_i[10]_pad  & n14331 ;
  assign n33981 = n14348 & n33980 ;
  assign n33982 = \m7_data_i[10]_pad  & ~n14331 ;
  assign n33983 = n14348 & n33982 ;
  assign n33984 = ~n33981 & ~n33983 ;
  assign n33985 = n33979 & n33984 ;
  assign n33986 = \m5_data_i[10]_pad  & ~n14331 ;
  assign n33987 = n14356 & n33986 ;
  assign n33988 = \m0_data_i[10]_pad  & n14331 ;
  assign n33989 = n14324 & n33988 ;
  assign n33990 = ~n33987 & ~n33989 ;
  assign n33991 = \m1_data_i[10]_pad  & ~n14331 ;
  assign n33992 = n14324 & n33991 ;
  assign n33993 = \m2_data_i[10]_pad  & n14331 ;
  assign n33994 = n14339 & n33993 ;
  assign n33995 = ~n33992 & ~n33994 ;
  assign n33996 = n33990 & n33995 ;
  assign n33997 = n33985 & n33996 ;
  assign n33998 = \m3_data_i[11]_pad  & ~n14331 ;
  assign n33999 = n14339 & n33998 ;
  assign n34000 = \m4_data_i[11]_pad  & n14331 ;
  assign n34001 = n14356 & n34000 ;
  assign n34002 = ~n33999 & ~n34001 ;
  assign n34003 = \m6_data_i[11]_pad  & n14331 ;
  assign n34004 = n14348 & n34003 ;
  assign n34005 = \m2_data_i[11]_pad  & n14331 ;
  assign n34006 = n14339 & n34005 ;
  assign n34007 = ~n34004 & ~n34006 ;
  assign n34008 = n34002 & n34007 ;
  assign n34009 = \m5_data_i[11]_pad  & ~n14331 ;
  assign n34010 = n14356 & n34009 ;
  assign n34011 = \m1_data_i[11]_pad  & ~n14331 ;
  assign n34012 = n14324 & n34011 ;
  assign n34013 = ~n34010 & ~n34012 ;
  assign n34014 = \m0_data_i[11]_pad  & n14331 ;
  assign n34015 = n14324 & n34014 ;
  assign n34016 = \m7_data_i[11]_pad  & ~n14331 ;
  assign n34017 = n14348 & n34016 ;
  assign n34018 = ~n34015 & ~n34017 ;
  assign n34019 = n34013 & n34018 ;
  assign n34020 = n34008 & n34019 ;
  assign n34021 = \m3_data_i[12]_pad  & ~n14331 ;
  assign n34022 = n14339 & n34021 ;
  assign n34023 = \m4_data_i[12]_pad  & n14331 ;
  assign n34024 = n14356 & n34023 ;
  assign n34025 = ~n34022 & ~n34024 ;
  assign n34026 = \m6_data_i[12]_pad  & n14331 ;
  assign n34027 = n14348 & n34026 ;
  assign n34028 = \m2_data_i[12]_pad  & n14331 ;
  assign n34029 = n14339 & n34028 ;
  assign n34030 = ~n34027 & ~n34029 ;
  assign n34031 = n34025 & n34030 ;
  assign n34032 = \m5_data_i[12]_pad  & ~n14331 ;
  assign n34033 = n14356 & n34032 ;
  assign n34034 = \m1_data_i[12]_pad  & ~n14331 ;
  assign n34035 = n14324 & n34034 ;
  assign n34036 = ~n34033 & ~n34035 ;
  assign n34037 = \m0_data_i[12]_pad  & n14331 ;
  assign n34038 = n14324 & n34037 ;
  assign n34039 = \m7_data_i[12]_pad  & ~n14331 ;
  assign n34040 = n14348 & n34039 ;
  assign n34041 = ~n34038 & ~n34040 ;
  assign n34042 = n34036 & n34041 ;
  assign n34043 = n34031 & n34042 ;
  assign n34044 = \m3_data_i[13]_pad  & ~n14331 ;
  assign n34045 = n14339 & n34044 ;
  assign n34046 = \m4_data_i[13]_pad  & n14331 ;
  assign n34047 = n14356 & n34046 ;
  assign n34048 = ~n34045 & ~n34047 ;
  assign n34049 = \m6_data_i[13]_pad  & n14331 ;
  assign n34050 = n14348 & n34049 ;
  assign n34051 = \m2_data_i[13]_pad  & n14331 ;
  assign n34052 = n14339 & n34051 ;
  assign n34053 = ~n34050 & ~n34052 ;
  assign n34054 = n34048 & n34053 ;
  assign n34055 = \m5_data_i[13]_pad  & ~n14331 ;
  assign n34056 = n14356 & n34055 ;
  assign n34057 = \m1_data_i[13]_pad  & ~n14331 ;
  assign n34058 = n14324 & n34057 ;
  assign n34059 = ~n34056 & ~n34058 ;
  assign n34060 = \m0_data_i[13]_pad  & n14331 ;
  assign n34061 = n14324 & n34060 ;
  assign n34062 = \m7_data_i[13]_pad  & ~n14331 ;
  assign n34063 = n14348 & n34062 ;
  assign n34064 = ~n34061 & ~n34063 ;
  assign n34065 = n34059 & n34064 ;
  assign n34066 = n34054 & n34065 ;
  assign n34067 = \m3_data_i[14]_pad  & ~n14331 ;
  assign n34068 = n14339 & n34067 ;
  assign n34069 = \m4_data_i[14]_pad  & n14331 ;
  assign n34070 = n14356 & n34069 ;
  assign n34071 = ~n34068 & ~n34070 ;
  assign n34072 = \m6_data_i[14]_pad  & n14331 ;
  assign n34073 = n14348 & n34072 ;
  assign n34074 = \m2_data_i[14]_pad  & n14331 ;
  assign n34075 = n14339 & n34074 ;
  assign n34076 = ~n34073 & ~n34075 ;
  assign n34077 = n34071 & n34076 ;
  assign n34078 = \m5_data_i[14]_pad  & ~n14331 ;
  assign n34079 = n14356 & n34078 ;
  assign n34080 = \m1_data_i[14]_pad  & ~n14331 ;
  assign n34081 = n14324 & n34080 ;
  assign n34082 = ~n34079 & ~n34081 ;
  assign n34083 = \m0_data_i[14]_pad  & n14331 ;
  assign n34084 = n14324 & n34083 ;
  assign n34085 = \m7_data_i[14]_pad  & ~n14331 ;
  assign n34086 = n14348 & n34085 ;
  assign n34087 = ~n34084 & ~n34086 ;
  assign n34088 = n34082 & n34087 ;
  assign n34089 = n34077 & n34088 ;
  assign n34090 = \m3_data_i[15]_pad  & ~n14331 ;
  assign n34091 = n14339 & n34090 ;
  assign n34092 = \m4_data_i[15]_pad  & n14331 ;
  assign n34093 = n14356 & n34092 ;
  assign n34094 = ~n34091 & ~n34093 ;
  assign n34095 = \m6_data_i[15]_pad  & n14331 ;
  assign n34096 = n14348 & n34095 ;
  assign n34097 = \m2_data_i[15]_pad  & n14331 ;
  assign n34098 = n14339 & n34097 ;
  assign n34099 = ~n34096 & ~n34098 ;
  assign n34100 = n34094 & n34099 ;
  assign n34101 = \m5_data_i[15]_pad  & ~n14331 ;
  assign n34102 = n14356 & n34101 ;
  assign n34103 = \m1_data_i[15]_pad  & ~n14331 ;
  assign n34104 = n14324 & n34103 ;
  assign n34105 = ~n34102 & ~n34104 ;
  assign n34106 = \m0_data_i[15]_pad  & n14331 ;
  assign n34107 = n14324 & n34106 ;
  assign n34108 = \m7_data_i[15]_pad  & ~n14331 ;
  assign n34109 = n14348 & n34108 ;
  assign n34110 = ~n34107 & ~n34109 ;
  assign n34111 = n34105 & n34110 ;
  assign n34112 = n34100 & n34111 ;
  assign n34113 = \m3_data_i[16]_pad  & ~n14331 ;
  assign n34114 = n14339 & n34113 ;
  assign n34115 = \m4_data_i[16]_pad  & n14331 ;
  assign n34116 = n14356 & n34115 ;
  assign n34117 = ~n34114 & ~n34116 ;
  assign n34118 = \m6_data_i[16]_pad  & n14331 ;
  assign n34119 = n14348 & n34118 ;
  assign n34120 = \m2_data_i[16]_pad  & n14331 ;
  assign n34121 = n14339 & n34120 ;
  assign n34122 = ~n34119 & ~n34121 ;
  assign n34123 = n34117 & n34122 ;
  assign n34124 = \m5_data_i[16]_pad  & ~n14331 ;
  assign n34125 = n14356 & n34124 ;
  assign n34126 = \m1_data_i[16]_pad  & ~n14331 ;
  assign n34127 = n14324 & n34126 ;
  assign n34128 = ~n34125 & ~n34127 ;
  assign n34129 = \m0_data_i[16]_pad  & n14331 ;
  assign n34130 = n14324 & n34129 ;
  assign n34131 = \m7_data_i[16]_pad  & ~n14331 ;
  assign n34132 = n14348 & n34131 ;
  assign n34133 = ~n34130 & ~n34132 ;
  assign n34134 = n34128 & n34133 ;
  assign n34135 = n34123 & n34134 ;
  assign n34136 = \m3_data_i[17]_pad  & ~n14331 ;
  assign n34137 = n14339 & n34136 ;
  assign n34138 = \m4_data_i[17]_pad  & n14331 ;
  assign n34139 = n14356 & n34138 ;
  assign n34140 = ~n34137 & ~n34139 ;
  assign n34141 = \m6_data_i[17]_pad  & n14331 ;
  assign n34142 = n14348 & n34141 ;
  assign n34143 = \m2_data_i[17]_pad  & n14331 ;
  assign n34144 = n14339 & n34143 ;
  assign n34145 = ~n34142 & ~n34144 ;
  assign n34146 = n34140 & n34145 ;
  assign n34147 = \m5_data_i[17]_pad  & ~n14331 ;
  assign n34148 = n14356 & n34147 ;
  assign n34149 = \m1_data_i[17]_pad  & ~n14331 ;
  assign n34150 = n14324 & n34149 ;
  assign n34151 = ~n34148 & ~n34150 ;
  assign n34152 = \m0_data_i[17]_pad  & n14331 ;
  assign n34153 = n14324 & n34152 ;
  assign n34154 = \m7_data_i[17]_pad  & ~n14331 ;
  assign n34155 = n14348 & n34154 ;
  assign n34156 = ~n34153 & ~n34155 ;
  assign n34157 = n34151 & n34156 ;
  assign n34158 = n34146 & n34157 ;
  assign n34159 = \m3_data_i[18]_pad  & ~n14331 ;
  assign n34160 = n14339 & n34159 ;
  assign n34161 = \m4_data_i[18]_pad  & n14331 ;
  assign n34162 = n14356 & n34161 ;
  assign n34163 = ~n34160 & ~n34162 ;
  assign n34164 = \m6_data_i[18]_pad  & n14331 ;
  assign n34165 = n14348 & n34164 ;
  assign n34166 = \m2_data_i[18]_pad  & n14331 ;
  assign n34167 = n14339 & n34166 ;
  assign n34168 = ~n34165 & ~n34167 ;
  assign n34169 = n34163 & n34168 ;
  assign n34170 = \m5_data_i[18]_pad  & ~n14331 ;
  assign n34171 = n14356 & n34170 ;
  assign n34172 = \m1_data_i[18]_pad  & ~n14331 ;
  assign n34173 = n14324 & n34172 ;
  assign n34174 = ~n34171 & ~n34173 ;
  assign n34175 = \m0_data_i[18]_pad  & n14331 ;
  assign n34176 = n14324 & n34175 ;
  assign n34177 = \m7_data_i[18]_pad  & ~n14331 ;
  assign n34178 = n14348 & n34177 ;
  assign n34179 = ~n34176 & ~n34178 ;
  assign n34180 = n34174 & n34179 ;
  assign n34181 = n34169 & n34180 ;
  assign n34182 = \m6_data_i[19]_pad  & n14331 ;
  assign n34183 = n14348 & n34182 ;
  assign n34184 = \m5_data_i[19]_pad  & ~n14331 ;
  assign n34185 = n14356 & n34184 ;
  assign n34186 = ~n34183 & ~n34185 ;
  assign n34187 = \m0_data_i[19]_pad  & n14331 ;
  assign n34188 = n14324 & n34187 ;
  assign n34189 = \m4_data_i[19]_pad  & n14331 ;
  assign n34190 = n14356 & n34189 ;
  assign n34191 = ~n34188 & ~n34190 ;
  assign n34192 = n34186 & n34191 ;
  assign n34193 = \m7_data_i[19]_pad  & ~n14331 ;
  assign n34194 = n14348 & n34193 ;
  assign n34195 = \m3_data_i[19]_pad  & ~n14331 ;
  assign n34196 = n14339 & n34195 ;
  assign n34197 = ~n34194 & ~n34196 ;
  assign n34198 = \m1_data_i[19]_pad  & ~n14331 ;
  assign n34199 = n14324 & n34198 ;
  assign n34200 = \m2_data_i[19]_pad  & n14331 ;
  assign n34201 = n14339 & n34200 ;
  assign n34202 = ~n34199 & ~n34201 ;
  assign n34203 = n34197 & n34202 ;
  assign n34204 = n34192 & n34203 ;
  assign n34205 = \m3_data_i[1]_pad  & ~n14331 ;
  assign n34206 = n14339 & n34205 ;
  assign n34207 = \m4_data_i[1]_pad  & n14331 ;
  assign n34208 = n14356 & n34207 ;
  assign n34209 = ~n34206 & ~n34208 ;
  assign n34210 = \m6_data_i[1]_pad  & n14331 ;
  assign n34211 = n14348 & n34210 ;
  assign n34212 = \m2_data_i[1]_pad  & n14331 ;
  assign n34213 = n14339 & n34212 ;
  assign n34214 = ~n34211 & ~n34213 ;
  assign n34215 = n34209 & n34214 ;
  assign n34216 = \m5_data_i[1]_pad  & ~n14331 ;
  assign n34217 = n14356 & n34216 ;
  assign n34218 = \m1_data_i[1]_pad  & ~n14331 ;
  assign n34219 = n14324 & n34218 ;
  assign n34220 = ~n34217 & ~n34219 ;
  assign n34221 = \m0_data_i[1]_pad  & n14331 ;
  assign n34222 = n14324 & n34221 ;
  assign n34223 = \m7_data_i[1]_pad  & ~n14331 ;
  assign n34224 = n14348 & n34223 ;
  assign n34225 = ~n34222 & ~n34224 ;
  assign n34226 = n34220 & n34225 ;
  assign n34227 = n34215 & n34226 ;
  assign n34228 = \m3_data_i[20]_pad  & ~n14331 ;
  assign n34229 = n14339 & n34228 ;
  assign n34230 = \m4_data_i[20]_pad  & n14331 ;
  assign n34231 = n14356 & n34230 ;
  assign n34232 = ~n34229 & ~n34231 ;
  assign n34233 = \m6_data_i[20]_pad  & n14331 ;
  assign n34234 = n14348 & n34233 ;
  assign n34235 = \m2_data_i[20]_pad  & n14331 ;
  assign n34236 = n14339 & n34235 ;
  assign n34237 = ~n34234 & ~n34236 ;
  assign n34238 = n34232 & n34237 ;
  assign n34239 = \m5_data_i[20]_pad  & ~n14331 ;
  assign n34240 = n14356 & n34239 ;
  assign n34241 = \m1_data_i[20]_pad  & ~n14331 ;
  assign n34242 = n14324 & n34241 ;
  assign n34243 = ~n34240 & ~n34242 ;
  assign n34244 = \m0_data_i[20]_pad  & n14331 ;
  assign n34245 = n14324 & n34244 ;
  assign n34246 = \m7_data_i[20]_pad  & ~n14331 ;
  assign n34247 = n14348 & n34246 ;
  assign n34248 = ~n34245 & ~n34247 ;
  assign n34249 = n34243 & n34248 ;
  assign n34250 = n34238 & n34249 ;
  assign n34251 = \m1_data_i[21]_pad  & ~n14331 ;
  assign n34252 = n14324 & n34251 ;
  assign n34253 = \m2_data_i[21]_pad  & n14331 ;
  assign n34254 = n14339 & n34253 ;
  assign n34255 = ~n34252 & ~n34254 ;
  assign n34256 = \m6_data_i[21]_pad  & n14331 ;
  assign n34257 = n14348 & n34256 ;
  assign n34258 = \m7_data_i[21]_pad  & ~n14331 ;
  assign n34259 = n14348 & n34258 ;
  assign n34260 = ~n34257 & ~n34259 ;
  assign n34261 = n34255 & n34260 ;
  assign n34262 = \m5_data_i[21]_pad  & ~n14331 ;
  assign n34263 = n14356 & n34262 ;
  assign n34264 = \m0_data_i[21]_pad  & n14331 ;
  assign n34265 = n14324 & n34264 ;
  assign n34266 = ~n34263 & ~n34265 ;
  assign n34267 = \m3_data_i[21]_pad  & ~n14331 ;
  assign n34268 = n14339 & n34267 ;
  assign n34269 = \m4_data_i[21]_pad  & n14331 ;
  assign n34270 = n14356 & n34269 ;
  assign n34271 = ~n34268 & ~n34270 ;
  assign n34272 = n34266 & n34271 ;
  assign n34273 = n34261 & n34272 ;
  assign n34274 = \m3_data_i[22]_pad  & ~n14331 ;
  assign n34275 = n14339 & n34274 ;
  assign n34276 = \m4_data_i[22]_pad  & n14331 ;
  assign n34277 = n14356 & n34276 ;
  assign n34278 = ~n34275 & ~n34277 ;
  assign n34279 = \m6_data_i[22]_pad  & n14331 ;
  assign n34280 = n14348 & n34279 ;
  assign n34281 = \m2_data_i[22]_pad  & n14331 ;
  assign n34282 = n14339 & n34281 ;
  assign n34283 = ~n34280 & ~n34282 ;
  assign n34284 = n34278 & n34283 ;
  assign n34285 = \m5_data_i[22]_pad  & ~n14331 ;
  assign n34286 = n14356 & n34285 ;
  assign n34287 = \m1_data_i[22]_pad  & ~n14331 ;
  assign n34288 = n14324 & n34287 ;
  assign n34289 = ~n34286 & ~n34288 ;
  assign n34290 = \m0_data_i[22]_pad  & n14331 ;
  assign n34291 = n14324 & n34290 ;
  assign n34292 = \m7_data_i[22]_pad  & ~n14331 ;
  assign n34293 = n14348 & n34292 ;
  assign n34294 = ~n34291 & ~n34293 ;
  assign n34295 = n34289 & n34294 ;
  assign n34296 = n34284 & n34295 ;
  assign n34297 = \m3_data_i[23]_pad  & ~n14331 ;
  assign n34298 = n14339 & n34297 ;
  assign n34299 = \m4_data_i[23]_pad  & n14331 ;
  assign n34300 = n14356 & n34299 ;
  assign n34301 = ~n34298 & ~n34300 ;
  assign n34302 = \m6_data_i[23]_pad  & n14331 ;
  assign n34303 = n14348 & n34302 ;
  assign n34304 = \m2_data_i[23]_pad  & n14331 ;
  assign n34305 = n14339 & n34304 ;
  assign n34306 = ~n34303 & ~n34305 ;
  assign n34307 = n34301 & n34306 ;
  assign n34308 = \m5_data_i[23]_pad  & ~n14331 ;
  assign n34309 = n14356 & n34308 ;
  assign n34310 = \m1_data_i[23]_pad  & ~n14331 ;
  assign n34311 = n14324 & n34310 ;
  assign n34312 = ~n34309 & ~n34311 ;
  assign n34313 = \m0_data_i[23]_pad  & n14331 ;
  assign n34314 = n14324 & n34313 ;
  assign n34315 = \m7_data_i[23]_pad  & ~n14331 ;
  assign n34316 = n14348 & n34315 ;
  assign n34317 = ~n34314 & ~n34316 ;
  assign n34318 = n34312 & n34317 ;
  assign n34319 = n34307 & n34318 ;
  assign n34320 = \m3_data_i[24]_pad  & ~n14331 ;
  assign n34321 = n14339 & n34320 ;
  assign n34322 = \m4_data_i[24]_pad  & n14331 ;
  assign n34323 = n14356 & n34322 ;
  assign n34324 = ~n34321 & ~n34323 ;
  assign n34325 = \m6_data_i[24]_pad  & n14331 ;
  assign n34326 = n14348 & n34325 ;
  assign n34327 = \m2_data_i[24]_pad  & n14331 ;
  assign n34328 = n14339 & n34327 ;
  assign n34329 = ~n34326 & ~n34328 ;
  assign n34330 = n34324 & n34329 ;
  assign n34331 = \m5_data_i[24]_pad  & ~n14331 ;
  assign n34332 = n14356 & n34331 ;
  assign n34333 = \m1_data_i[24]_pad  & ~n14331 ;
  assign n34334 = n14324 & n34333 ;
  assign n34335 = ~n34332 & ~n34334 ;
  assign n34336 = \m0_data_i[24]_pad  & n14331 ;
  assign n34337 = n14324 & n34336 ;
  assign n34338 = \m7_data_i[24]_pad  & ~n14331 ;
  assign n34339 = n14348 & n34338 ;
  assign n34340 = ~n34337 & ~n34339 ;
  assign n34341 = n34335 & n34340 ;
  assign n34342 = n34330 & n34341 ;
  assign n34343 = \m3_data_i[25]_pad  & ~n14331 ;
  assign n34344 = n14339 & n34343 ;
  assign n34345 = \m4_data_i[25]_pad  & n14331 ;
  assign n34346 = n14356 & n34345 ;
  assign n34347 = ~n34344 & ~n34346 ;
  assign n34348 = \m6_data_i[25]_pad  & n14331 ;
  assign n34349 = n14348 & n34348 ;
  assign n34350 = \m2_data_i[25]_pad  & n14331 ;
  assign n34351 = n14339 & n34350 ;
  assign n34352 = ~n34349 & ~n34351 ;
  assign n34353 = n34347 & n34352 ;
  assign n34354 = \m5_data_i[25]_pad  & ~n14331 ;
  assign n34355 = n14356 & n34354 ;
  assign n34356 = \m1_data_i[25]_pad  & ~n14331 ;
  assign n34357 = n14324 & n34356 ;
  assign n34358 = ~n34355 & ~n34357 ;
  assign n34359 = \m0_data_i[25]_pad  & n14331 ;
  assign n34360 = n14324 & n34359 ;
  assign n34361 = \m7_data_i[25]_pad  & ~n14331 ;
  assign n34362 = n14348 & n34361 ;
  assign n34363 = ~n34360 & ~n34362 ;
  assign n34364 = n34358 & n34363 ;
  assign n34365 = n34353 & n34364 ;
  assign n34366 = \m3_data_i[26]_pad  & ~n14331 ;
  assign n34367 = n14339 & n34366 ;
  assign n34368 = \m4_data_i[26]_pad  & n14331 ;
  assign n34369 = n14356 & n34368 ;
  assign n34370 = ~n34367 & ~n34369 ;
  assign n34371 = \m6_data_i[26]_pad  & n14331 ;
  assign n34372 = n14348 & n34371 ;
  assign n34373 = \m2_data_i[26]_pad  & n14331 ;
  assign n34374 = n14339 & n34373 ;
  assign n34375 = ~n34372 & ~n34374 ;
  assign n34376 = n34370 & n34375 ;
  assign n34377 = \m5_data_i[26]_pad  & ~n14331 ;
  assign n34378 = n14356 & n34377 ;
  assign n34379 = \m1_data_i[26]_pad  & ~n14331 ;
  assign n34380 = n14324 & n34379 ;
  assign n34381 = ~n34378 & ~n34380 ;
  assign n34382 = \m0_data_i[26]_pad  & n14331 ;
  assign n34383 = n14324 & n34382 ;
  assign n34384 = \m7_data_i[26]_pad  & ~n14331 ;
  assign n34385 = n14348 & n34384 ;
  assign n34386 = ~n34383 & ~n34385 ;
  assign n34387 = n34381 & n34386 ;
  assign n34388 = n34376 & n34387 ;
  assign n34389 = \m3_data_i[27]_pad  & ~n14331 ;
  assign n34390 = n14339 & n34389 ;
  assign n34391 = \m4_data_i[27]_pad  & n14331 ;
  assign n34392 = n14356 & n34391 ;
  assign n34393 = ~n34390 & ~n34392 ;
  assign n34394 = \m6_data_i[27]_pad  & n14331 ;
  assign n34395 = n14348 & n34394 ;
  assign n34396 = \m2_data_i[27]_pad  & n14331 ;
  assign n34397 = n14339 & n34396 ;
  assign n34398 = ~n34395 & ~n34397 ;
  assign n34399 = n34393 & n34398 ;
  assign n34400 = \m5_data_i[27]_pad  & ~n14331 ;
  assign n34401 = n14356 & n34400 ;
  assign n34402 = \m1_data_i[27]_pad  & ~n14331 ;
  assign n34403 = n14324 & n34402 ;
  assign n34404 = ~n34401 & ~n34403 ;
  assign n34405 = \m0_data_i[27]_pad  & n14331 ;
  assign n34406 = n14324 & n34405 ;
  assign n34407 = \m7_data_i[27]_pad  & ~n14331 ;
  assign n34408 = n14348 & n34407 ;
  assign n34409 = ~n34406 & ~n34408 ;
  assign n34410 = n34404 & n34409 ;
  assign n34411 = n34399 & n34410 ;
  assign n34412 = \m3_data_i[28]_pad  & ~n14331 ;
  assign n34413 = n14339 & n34412 ;
  assign n34414 = \m4_data_i[28]_pad  & n14331 ;
  assign n34415 = n14356 & n34414 ;
  assign n34416 = ~n34413 & ~n34415 ;
  assign n34417 = \m6_data_i[28]_pad  & n14331 ;
  assign n34418 = n14348 & n34417 ;
  assign n34419 = \m2_data_i[28]_pad  & n14331 ;
  assign n34420 = n14339 & n34419 ;
  assign n34421 = ~n34418 & ~n34420 ;
  assign n34422 = n34416 & n34421 ;
  assign n34423 = \m5_data_i[28]_pad  & ~n14331 ;
  assign n34424 = n14356 & n34423 ;
  assign n34425 = \m1_data_i[28]_pad  & ~n14331 ;
  assign n34426 = n14324 & n34425 ;
  assign n34427 = ~n34424 & ~n34426 ;
  assign n34428 = \m0_data_i[28]_pad  & n14331 ;
  assign n34429 = n14324 & n34428 ;
  assign n34430 = \m7_data_i[28]_pad  & ~n14331 ;
  assign n34431 = n14348 & n34430 ;
  assign n34432 = ~n34429 & ~n34431 ;
  assign n34433 = n34427 & n34432 ;
  assign n34434 = n34422 & n34433 ;
  assign n34435 = \m3_data_i[29]_pad  & ~n14331 ;
  assign n34436 = n14339 & n34435 ;
  assign n34437 = \m4_data_i[29]_pad  & n14331 ;
  assign n34438 = n14356 & n34437 ;
  assign n34439 = ~n34436 & ~n34438 ;
  assign n34440 = \m0_data_i[29]_pad  & n14331 ;
  assign n34441 = n14324 & n34440 ;
  assign n34442 = \m5_data_i[29]_pad  & ~n14331 ;
  assign n34443 = n14356 & n34442 ;
  assign n34444 = ~n34441 & ~n34443 ;
  assign n34445 = n34439 & n34444 ;
  assign n34446 = \m7_data_i[29]_pad  & ~n14331 ;
  assign n34447 = n14348 & n34446 ;
  assign n34448 = \m6_data_i[29]_pad  & n14331 ;
  assign n34449 = n14348 & n34448 ;
  assign n34450 = ~n34447 & ~n34449 ;
  assign n34451 = \m1_data_i[29]_pad  & ~n14331 ;
  assign n34452 = n14324 & n34451 ;
  assign n34453 = \m2_data_i[29]_pad  & n14331 ;
  assign n34454 = n14339 & n34453 ;
  assign n34455 = ~n34452 & ~n34454 ;
  assign n34456 = n34450 & n34455 ;
  assign n34457 = n34445 & n34456 ;
  assign n34458 = \m3_data_i[2]_pad  & ~n14331 ;
  assign n34459 = n14339 & n34458 ;
  assign n34460 = \m4_data_i[2]_pad  & n14331 ;
  assign n34461 = n14356 & n34460 ;
  assign n34462 = ~n34459 & ~n34461 ;
  assign n34463 = \m6_data_i[2]_pad  & n14331 ;
  assign n34464 = n14348 & n34463 ;
  assign n34465 = \m2_data_i[2]_pad  & n14331 ;
  assign n34466 = n14339 & n34465 ;
  assign n34467 = ~n34464 & ~n34466 ;
  assign n34468 = n34462 & n34467 ;
  assign n34469 = \m5_data_i[2]_pad  & ~n14331 ;
  assign n34470 = n14356 & n34469 ;
  assign n34471 = \m1_data_i[2]_pad  & ~n14331 ;
  assign n34472 = n14324 & n34471 ;
  assign n34473 = ~n34470 & ~n34472 ;
  assign n34474 = \m0_data_i[2]_pad  & n14331 ;
  assign n34475 = n14324 & n34474 ;
  assign n34476 = \m7_data_i[2]_pad  & ~n14331 ;
  assign n34477 = n14348 & n34476 ;
  assign n34478 = ~n34475 & ~n34477 ;
  assign n34479 = n34473 & n34478 ;
  assign n34480 = n34468 & n34479 ;
  assign n34481 = \m3_data_i[30]_pad  & ~n14331 ;
  assign n34482 = n14339 & n34481 ;
  assign n34483 = \m4_data_i[30]_pad  & n14331 ;
  assign n34484 = n14356 & n34483 ;
  assign n34485 = ~n34482 & ~n34484 ;
  assign n34486 = \m0_data_i[30]_pad  & n14331 ;
  assign n34487 = n14324 & n34486 ;
  assign n34488 = \m5_data_i[30]_pad  & ~n14331 ;
  assign n34489 = n14356 & n34488 ;
  assign n34490 = ~n34487 & ~n34489 ;
  assign n34491 = n34485 & n34490 ;
  assign n34492 = \m7_data_i[30]_pad  & ~n14331 ;
  assign n34493 = n14348 & n34492 ;
  assign n34494 = \m6_data_i[30]_pad  & n14331 ;
  assign n34495 = n14348 & n34494 ;
  assign n34496 = ~n34493 & ~n34495 ;
  assign n34497 = \m1_data_i[30]_pad  & ~n14331 ;
  assign n34498 = n14324 & n34497 ;
  assign n34499 = \m2_data_i[30]_pad  & n14331 ;
  assign n34500 = n14339 & n34499 ;
  assign n34501 = ~n34498 & ~n34500 ;
  assign n34502 = n34496 & n34501 ;
  assign n34503 = n34491 & n34502 ;
  assign n34504 = \m1_data_i[31]_pad  & ~n14331 ;
  assign n34505 = n14324 & n34504 ;
  assign n34506 = \m2_data_i[31]_pad  & n14331 ;
  assign n34507 = n14339 & n34506 ;
  assign n34508 = ~n34505 & ~n34507 ;
  assign n34509 = \m6_data_i[31]_pad  & n14331 ;
  assign n34510 = n14348 & n34509 ;
  assign n34511 = \m7_data_i[31]_pad  & ~n14331 ;
  assign n34512 = n14348 & n34511 ;
  assign n34513 = ~n34510 & ~n34512 ;
  assign n34514 = n34508 & n34513 ;
  assign n34515 = \m5_data_i[31]_pad  & ~n14331 ;
  assign n34516 = n14356 & n34515 ;
  assign n34517 = \m0_data_i[31]_pad  & n14331 ;
  assign n34518 = n14324 & n34517 ;
  assign n34519 = ~n34516 & ~n34518 ;
  assign n34520 = \m3_data_i[31]_pad  & ~n14331 ;
  assign n34521 = n14339 & n34520 ;
  assign n34522 = \m4_data_i[31]_pad  & n14331 ;
  assign n34523 = n14356 & n34522 ;
  assign n34524 = ~n34521 & ~n34523 ;
  assign n34525 = n34519 & n34524 ;
  assign n34526 = n34514 & n34525 ;
  assign n34527 = \m3_data_i[3]_pad  & ~n14331 ;
  assign n34528 = n14339 & n34527 ;
  assign n34529 = \m4_data_i[3]_pad  & n14331 ;
  assign n34530 = n14356 & n34529 ;
  assign n34531 = ~n34528 & ~n34530 ;
  assign n34532 = \m6_data_i[3]_pad  & n14331 ;
  assign n34533 = n14348 & n34532 ;
  assign n34534 = \m2_data_i[3]_pad  & n14331 ;
  assign n34535 = n14339 & n34534 ;
  assign n34536 = ~n34533 & ~n34535 ;
  assign n34537 = n34531 & n34536 ;
  assign n34538 = \m5_data_i[3]_pad  & ~n14331 ;
  assign n34539 = n14356 & n34538 ;
  assign n34540 = \m1_data_i[3]_pad  & ~n14331 ;
  assign n34541 = n14324 & n34540 ;
  assign n34542 = ~n34539 & ~n34541 ;
  assign n34543 = \m0_data_i[3]_pad  & n14331 ;
  assign n34544 = n14324 & n34543 ;
  assign n34545 = \m7_data_i[3]_pad  & ~n14331 ;
  assign n34546 = n14348 & n34545 ;
  assign n34547 = ~n34544 & ~n34546 ;
  assign n34548 = n34542 & n34547 ;
  assign n34549 = n34537 & n34548 ;
  assign n34550 = \m6_data_i[4]_pad  & n14331 ;
  assign n34551 = n14348 & n34550 ;
  assign n34552 = \m5_data_i[4]_pad  & ~n14331 ;
  assign n34553 = n14356 & n34552 ;
  assign n34554 = ~n34551 & ~n34553 ;
  assign n34555 = \m3_data_i[4]_pad  & ~n14331 ;
  assign n34556 = n14339 & n34555 ;
  assign n34557 = \m2_data_i[4]_pad  & n14331 ;
  assign n34558 = n14339 & n34557 ;
  assign n34559 = ~n34556 & ~n34558 ;
  assign n34560 = n34554 & n34559 ;
  assign n34561 = \m4_data_i[4]_pad  & n14331 ;
  assign n34562 = n14356 & n34561 ;
  assign n34563 = \m1_data_i[4]_pad  & ~n14331 ;
  assign n34564 = n14324 & n34563 ;
  assign n34565 = ~n34562 & ~n34564 ;
  assign n34566 = \m0_data_i[4]_pad  & n14331 ;
  assign n34567 = n14324 & n34566 ;
  assign n34568 = \m7_data_i[4]_pad  & ~n14331 ;
  assign n34569 = n14348 & n34568 ;
  assign n34570 = ~n34567 & ~n34569 ;
  assign n34571 = n34565 & n34570 ;
  assign n34572 = n34560 & n34571 ;
  assign n34573 = \m3_data_i[5]_pad  & ~n14331 ;
  assign n34574 = n14339 & n34573 ;
  assign n34575 = \m4_data_i[5]_pad  & n14331 ;
  assign n34576 = n14356 & n34575 ;
  assign n34577 = ~n34574 & ~n34576 ;
  assign n34578 = \m6_data_i[5]_pad  & n14331 ;
  assign n34579 = n14348 & n34578 ;
  assign n34580 = \m2_data_i[5]_pad  & n14331 ;
  assign n34581 = n14339 & n34580 ;
  assign n34582 = ~n34579 & ~n34581 ;
  assign n34583 = n34577 & n34582 ;
  assign n34584 = \m5_data_i[5]_pad  & ~n14331 ;
  assign n34585 = n14356 & n34584 ;
  assign n34586 = \m1_data_i[5]_pad  & ~n14331 ;
  assign n34587 = n14324 & n34586 ;
  assign n34588 = ~n34585 & ~n34587 ;
  assign n34589 = \m0_data_i[5]_pad  & n14331 ;
  assign n34590 = n14324 & n34589 ;
  assign n34591 = \m7_data_i[5]_pad  & ~n14331 ;
  assign n34592 = n14348 & n34591 ;
  assign n34593 = ~n34590 & ~n34592 ;
  assign n34594 = n34588 & n34593 ;
  assign n34595 = n34583 & n34594 ;
  assign n34596 = \m3_data_i[6]_pad  & ~n14331 ;
  assign n34597 = n14339 & n34596 ;
  assign n34598 = \m4_data_i[6]_pad  & n14331 ;
  assign n34599 = n14356 & n34598 ;
  assign n34600 = ~n34597 & ~n34599 ;
  assign n34601 = \m6_data_i[6]_pad  & n14331 ;
  assign n34602 = n14348 & n34601 ;
  assign n34603 = \m2_data_i[6]_pad  & n14331 ;
  assign n34604 = n14339 & n34603 ;
  assign n34605 = ~n34602 & ~n34604 ;
  assign n34606 = n34600 & n34605 ;
  assign n34607 = \m5_data_i[6]_pad  & ~n14331 ;
  assign n34608 = n14356 & n34607 ;
  assign n34609 = \m1_data_i[6]_pad  & ~n14331 ;
  assign n34610 = n14324 & n34609 ;
  assign n34611 = ~n34608 & ~n34610 ;
  assign n34612 = \m0_data_i[6]_pad  & n14331 ;
  assign n34613 = n14324 & n34612 ;
  assign n34614 = \m7_data_i[6]_pad  & ~n14331 ;
  assign n34615 = n14348 & n34614 ;
  assign n34616 = ~n34613 & ~n34615 ;
  assign n34617 = n34611 & n34616 ;
  assign n34618 = n34606 & n34617 ;
  assign n34619 = \m6_data_i[7]_pad  & n14331 ;
  assign n34620 = n14348 & n34619 ;
  assign n34621 = \m5_data_i[7]_pad  & ~n14331 ;
  assign n34622 = n14356 & n34621 ;
  assign n34623 = ~n34620 & ~n34622 ;
  assign n34624 = \m0_data_i[7]_pad  & n14331 ;
  assign n34625 = n14324 & n34624 ;
  assign n34626 = \m4_data_i[7]_pad  & n14331 ;
  assign n34627 = n14356 & n34626 ;
  assign n34628 = ~n34625 & ~n34627 ;
  assign n34629 = n34623 & n34628 ;
  assign n34630 = \m7_data_i[7]_pad  & ~n14331 ;
  assign n34631 = n14348 & n34630 ;
  assign n34632 = \m3_data_i[7]_pad  & ~n14331 ;
  assign n34633 = n14339 & n34632 ;
  assign n34634 = ~n34631 & ~n34633 ;
  assign n34635 = \m1_data_i[7]_pad  & ~n14331 ;
  assign n34636 = n14324 & n34635 ;
  assign n34637 = \m2_data_i[7]_pad  & n14331 ;
  assign n34638 = n14339 & n34637 ;
  assign n34639 = ~n34636 & ~n34638 ;
  assign n34640 = n34634 & n34639 ;
  assign n34641 = n34629 & n34640 ;
  assign n34642 = \m3_data_i[8]_pad  & ~n14331 ;
  assign n34643 = n14339 & n34642 ;
  assign n34644 = \m4_data_i[8]_pad  & n14331 ;
  assign n34645 = n14356 & n34644 ;
  assign n34646 = ~n34643 & ~n34645 ;
  assign n34647 = \m6_data_i[8]_pad  & n14331 ;
  assign n34648 = n14348 & n34647 ;
  assign n34649 = \m2_data_i[8]_pad  & n14331 ;
  assign n34650 = n14339 & n34649 ;
  assign n34651 = ~n34648 & ~n34650 ;
  assign n34652 = n34646 & n34651 ;
  assign n34653 = \m5_data_i[8]_pad  & ~n14331 ;
  assign n34654 = n14356 & n34653 ;
  assign n34655 = \m1_data_i[8]_pad  & ~n14331 ;
  assign n34656 = n14324 & n34655 ;
  assign n34657 = ~n34654 & ~n34656 ;
  assign n34658 = \m0_data_i[8]_pad  & n14331 ;
  assign n34659 = n14324 & n34658 ;
  assign n34660 = \m7_data_i[8]_pad  & ~n14331 ;
  assign n34661 = n14348 & n34660 ;
  assign n34662 = ~n34659 & ~n34661 ;
  assign n34663 = n34657 & n34662 ;
  assign n34664 = n34652 & n34663 ;
  assign n34665 = \m3_data_i[9]_pad  & ~n14331 ;
  assign n34666 = n14339 & n34665 ;
  assign n34667 = \m4_data_i[9]_pad  & n14331 ;
  assign n34668 = n14356 & n34667 ;
  assign n34669 = ~n34666 & ~n34668 ;
  assign n34670 = \m6_data_i[9]_pad  & n14331 ;
  assign n34671 = n14348 & n34670 ;
  assign n34672 = \m2_data_i[9]_pad  & n14331 ;
  assign n34673 = n14339 & n34672 ;
  assign n34674 = ~n34671 & ~n34673 ;
  assign n34675 = n34669 & n34674 ;
  assign n34676 = \m5_data_i[9]_pad  & ~n14331 ;
  assign n34677 = n14356 & n34676 ;
  assign n34678 = \m1_data_i[9]_pad  & ~n14331 ;
  assign n34679 = n14324 & n34678 ;
  assign n34680 = ~n34677 & ~n34679 ;
  assign n34681 = \m0_data_i[9]_pad  & n14331 ;
  assign n34682 = n14324 & n34681 ;
  assign n34683 = \m7_data_i[9]_pad  & ~n14331 ;
  assign n34684 = n14348 & n34683 ;
  assign n34685 = ~n34682 & ~n34684 ;
  assign n34686 = n34680 & n34685 ;
  assign n34687 = n34675 & n34686 ;
  assign n34688 = \m3_sel_i[0]_pad  & ~n14331 ;
  assign n34689 = n14339 & n34688 ;
  assign n34690 = \m4_sel_i[0]_pad  & n14331 ;
  assign n34691 = n14356 & n34690 ;
  assign n34692 = ~n34689 & ~n34691 ;
  assign n34693 = \m6_sel_i[0]_pad  & n14331 ;
  assign n34694 = n14348 & n34693 ;
  assign n34695 = \m2_sel_i[0]_pad  & n14331 ;
  assign n34696 = n14339 & n34695 ;
  assign n34697 = ~n34694 & ~n34696 ;
  assign n34698 = n34692 & n34697 ;
  assign n34699 = \m5_sel_i[0]_pad  & ~n14331 ;
  assign n34700 = n14356 & n34699 ;
  assign n34701 = \m1_sel_i[0]_pad  & ~n14331 ;
  assign n34702 = n14324 & n34701 ;
  assign n34703 = ~n34700 & ~n34702 ;
  assign n34704 = \m0_sel_i[0]_pad  & n14331 ;
  assign n34705 = n14324 & n34704 ;
  assign n34706 = \m7_sel_i[0]_pad  & ~n14331 ;
  assign n34707 = n14348 & n34706 ;
  assign n34708 = ~n34705 & ~n34707 ;
  assign n34709 = n34703 & n34708 ;
  assign n34710 = n34698 & n34709 ;
  assign n34711 = \m3_sel_i[1]_pad  & ~n14331 ;
  assign n34712 = n14339 & n34711 ;
  assign n34713 = \m4_sel_i[1]_pad  & n14331 ;
  assign n34714 = n14356 & n34713 ;
  assign n34715 = ~n34712 & ~n34714 ;
  assign n34716 = \m6_sel_i[1]_pad  & n14331 ;
  assign n34717 = n14348 & n34716 ;
  assign n34718 = \m2_sel_i[1]_pad  & n14331 ;
  assign n34719 = n14339 & n34718 ;
  assign n34720 = ~n34717 & ~n34719 ;
  assign n34721 = n34715 & n34720 ;
  assign n34722 = \m5_sel_i[1]_pad  & ~n14331 ;
  assign n34723 = n14356 & n34722 ;
  assign n34724 = \m1_sel_i[1]_pad  & ~n14331 ;
  assign n34725 = n14324 & n34724 ;
  assign n34726 = ~n34723 & ~n34725 ;
  assign n34727 = \m0_sel_i[1]_pad  & n14331 ;
  assign n34728 = n14324 & n34727 ;
  assign n34729 = \m7_sel_i[1]_pad  & ~n14331 ;
  assign n34730 = n14348 & n34729 ;
  assign n34731 = ~n34728 & ~n34730 ;
  assign n34732 = n34726 & n34731 ;
  assign n34733 = n34721 & n34732 ;
  assign n34734 = \m6_sel_i[2]_pad  & n14331 ;
  assign n34735 = n14348 & n34734 ;
  assign n34736 = \m5_sel_i[2]_pad  & ~n14331 ;
  assign n34737 = n14356 & n34736 ;
  assign n34738 = ~n34735 & ~n34737 ;
  assign n34739 = \m3_sel_i[2]_pad  & ~n14331 ;
  assign n34740 = n14339 & n34739 ;
  assign n34741 = \m2_sel_i[2]_pad  & n14331 ;
  assign n34742 = n14339 & n34741 ;
  assign n34743 = ~n34740 & ~n34742 ;
  assign n34744 = n34738 & n34743 ;
  assign n34745 = \m4_sel_i[2]_pad  & n14331 ;
  assign n34746 = n14356 & n34745 ;
  assign n34747 = \m1_sel_i[2]_pad  & ~n14331 ;
  assign n34748 = n14324 & n34747 ;
  assign n34749 = ~n34746 & ~n34748 ;
  assign n34750 = \m0_sel_i[2]_pad  & n14331 ;
  assign n34751 = n14324 & n34750 ;
  assign n34752 = \m7_sel_i[2]_pad  & ~n14331 ;
  assign n34753 = n14348 & n34752 ;
  assign n34754 = ~n34751 & ~n34753 ;
  assign n34755 = n34749 & n34754 ;
  assign n34756 = n34744 & n34755 ;
  assign n34757 = \m1_sel_i[3]_pad  & ~n14331 ;
  assign n34758 = n14324 & n34757 ;
  assign n34759 = \m2_sel_i[3]_pad  & n14331 ;
  assign n34760 = n14339 & n34759 ;
  assign n34761 = ~n34758 & ~n34760 ;
  assign n34762 = \m6_sel_i[3]_pad  & n14331 ;
  assign n34763 = n14348 & n34762 ;
  assign n34764 = \m4_sel_i[3]_pad  & n14331 ;
  assign n34765 = n14356 & n34764 ;
  assign n34766 = ~n34763 & ~n34765 ;
  assign n34767 = n34761 & n34766 ;
  assign n34768 = \m5_sel_i[3]_pad  & ~n14331 ;
  assign n34769 = n14356 & n34768 ;
  assign n34770 = \m3_sel_i[3]_pad  & ~n14331 ;
  assign n34771 = n14339 & n34770 ;
  assign n34772 = ~n34769 & ~n34771 ;
  assign n34773 = \m0_sel_i[3]_pad  & n14331 ;
  assign n34774 = n14324 & n34773 ;
  assign n34775 = \m7_sel_i[3]_pad  & ~n14331 ;
  assign n34776 = n14348 & n34775 ;
  assign n34777 = ~n34774 & ~n34776 ;
  assign n34778 = n34772 & n34777 ;
  assign n34779 = n34767 & n34778 ;
  assign n34780 = \m3_stb_i_pad  & n14915 ;
  assign n34781 = ~n14331 & n34780 ;
  assign n34782 = n14339 & n34781 ;
  assign n34783 = \m2_stb_i_pad  & n15098 ;
  assign n34784 = n14331 & n34783 ;
  assign n34785 = n14339 & n34784 ;
  assign n34786 = ~n34782 & ~n34785 ;
  assign n34787 = \m4_stb_i_pad  & n14939 ;
  assign n34788 = n14331 & n34787 ;
  assign n34789 = n14356 & n34788 ;
  assign n34790 = \m6_stb_i_pad  & n15015 ;
  assign n34791 = n14331 & n34790 ;
  assign n34792 = n14348 & n34791 ;
  assign n34793 = ~n34789 & ~n34792 ;
  assign n34794 = n34786 & n34793 ;
  assign n34795 = \m5_stb_i_pad  & n14700 ;
  assign n34796 = ~n14331 & n34795 ;
  assign n34797 = n14356 & n34796 ;
  assign n34798 = \m7_stb_i_pad  & n15059 ;
  assign n34799 = ~n14331 & n34798 ;
  assign n34800 = n14348 & n34799 ;
  assign n34801 = ~n34797 & ~n34800 ;
  assign n34802 = \m1_stb_i_pad  & n14809 ;
  assign n34803 = ~n14331 & n34802 ;
  assign n34804 = n14324 & n34803 ;
  assign n34805 = \m0_stb_i_pad  & n14762 ;
  assign n34806 = n14331 & n34805 ;
  assign n34807 = n14324 & n34806 ;
  assign n34808 = ~n34804 & ~n34807 ;
  assign n34809 = n34801 & n34808 ;
  assign n34810 = n34794 & n34809 ;
  assign n34811 = \m3_we_i_pad  & ~n14331 ;
  assign n34812 = n14339 & n34811 ;
  assign n34813 = \m4_we_i_pad  & n14331 ;
  assign n34814 = n14356 & n34813 ;
  assign n34815 = ~n34812 & ~n34814 ;
  assign n34816 = \m6_we_i_pad  & n14331 ;
  assign n34817 = n14348 & n34816 ;
  assign n34818 = \m2_we_i_pad  & n14331 ;
  assign n34819 = n14339 & n34818 ;
  assign n34820 = ~n34817 & ~n34819 ;
  assign n34821 = n34815 & n34820 ;
  assign n34822 = \m5_we_i_pad  & ~n14331 ;
  assign n34823 = n14356 & n34822 ;
  assign n34824 = \m1_we_i_pad  & ~n14331 ;
  assign n34825 = n14324 & n34824 ;
  assign n34826 = ~n34823 & ~n34825 ;
  assign n34827 = \m0_we_i_pad  & n14331 ;
  assign n34828 = n14324 & n34827 ;
  assign n34829 = \m7_we_i_pad  & ~n14331 ;
  assign n34830 = n14348 & n34829 ;
  assign n34831 = ~n34828 & ~n34830 ;
  assign n34832 = n34826 & n34831 ;
  assign n34833 = n34821 & n34832 ;
  assign n34834 = \m7_addr_i[0]_pad  & ~n1910 ;
  assign n34835 = n1938 & n34834 ;
  assign n34836 = \m6_addr_i[0]_pad  & ~n1925 ;
  assign n34837 = n1918 & n34836 ;
  assign n34838 = ~n34835 & ~n34837 ;
  assign n34839 = \m5_addr_i[0]_pad  & ~n1910 ;
  assign n34840 = n1941 & n34839 ;
  assign n34841 = \m2_addr_i[0]_pad  & ~n1925 ;
  assign n34842 = n1931 & n34841 ;
  assign n34843 = ~n34840 & ~n34842 ;
  assign n34844 = n34838 & n34843 ;
  assign n34845 = \m4_addr_i[0]_pad  & n1925 ;
  assign n34846 = n1918 & n34845 ;
  assign n34847 = \m3_addr_i[0]_pad  & n1910 ;
  assign n34848 = n1938 & n34847 ;
  assign n34849 = ~n34846 & ~n34848 ;
  assign n34850 = \m1_addr_i[0]_pad  & n1910 ;
  assign n34851 = n1941 & n34850 ;
  assign n34852 = \m0_addr_i[0]_pad  & n1925 ;
  assign n34853 = n1931 & n34852 ;
  assign n34854 = ~n34851 & ~n34853 ;
  assign n34855 = n34849 & n34854 ;
  assign n34856 = n34844 & n34855 ;
  assign n34857 = \m7_addr_i[10]_pad  & ~n1910 ;
  assign n34858 = n1938 & n34857 ;
  assign n34859 = \m6_addr_i[10]_pad  & ~n1925 ;
  assign n34860 = n1918 & n34859 ;
  assign n34861 = ~n34858 & ~n34860 ;
  assign n34862 = \m5_addr_i[10]_pad  & ~n1910 ;
  assign n34863 = n1941 & n34862 ;
  assign n34864 = \m2_addr_i[10]_pad  & ~n1925 ;
  assign n34865 = n1931 & n34864 ;
  assign n34866 = ~n34863 & ~n34865 ;
  assign n34867 = n34861 & n34866 ;
  assign n34868 = \m4_addr_i[10]_pad  & n1925 ;
  assign n34869 = n1918 & n34868 ;
  assign n34870 = \m3_addr_i[10]_pad  & n1910 ;
  assign n34871 = n1938 & n34870 ;
  assign n34872 = ~n34869 & ~n34871 ;
  assign n34873 = \m1_addr_i[10]_pad  & n1910 ;
  assign n34874 = n1941 & n34873 ;
  assign n34875 = \m0_addr_i[10]_pad  & n1925 ;
  assign n34876 = n1931 & n34875 ;
  assign n34877 = ~n34874 & ~n34876 ;
  assign n34878 = n34872 & n34877 ;
  assign n34879 = n34867 & n34878 ;
  assign n34880 = \m7_addr_i[11]_pad  & ~n1910 ;
  assign n34881 = n1938 & n34880 ;
  assign n34882 = \m6_addr_i[11]_pad  & ~n1925 ;
  assign n34883 = n1918 & n34882 ;
  assign n34884 = ~n34881 & ~n34883 ;
  assign n34885 = \m5_addr_i[11]_pad  & ~n1910 ;
  assign n34886 = n1941 & n34885 ;
  assign n34887 = \m2_addr_i[11]_pad  & ~n1925 ;
  assign n34888 = n1931 & n34887 ;
  assign n34889 = ~n34886 & ~n34888 ;
  assign n34890 = n34884 & n34889 ;
  assign n34891 = \m4_addr_i[11]_pad  & n1925 ;
  assign n34892 = n1918 & n34891 ;
  assign n34893 = \m3_addr_i[11]_pad  & n1910 ;
  assign n34894 = n1938 & n34893 ;
  assign n34895 = ~n34892 & ~n34894 ;
  assign n34896 = \m1_addr_i[11]_pad  & n1910 ;
  assign n34897 = n1941 & n34896 ;
  assign n34898 = \m0_addr_i[11]_pad  & n1925 ;
  assign n34899 = n1931 & n34898 ;
  assign n34900 = ~n34897 & ~n34899 ;
  assign n34901 = n34895 & n34900 ;
  assign n34902 = n34890 & n34901 ;
  assign n34903 = \m7_addr_i[12]_pad  & ~n1910 ;
  assign n34904 = n1938 & n34903 ;
  assign n34905 = \m6_addr_i[12]_pad  & ~n1925 ;
  assign n34906 = n1918 & n34905 ;
  assign n34907 = ~n34904 & ~n34906 ;
  assign n34908 = \m5_addr_i[12]_pad  & ~n1910 ;
  assign n34909 = n1941 & n34908 ;
  assign n34910 = \m2_addr_i[12]_pad  & ~n1925 ;
  assign n34911 = n1931 & n34910 ;
  assign n34912 = ~n34909 & ~n34911 ;
  assign n34913 = n34907 & n34912 ;
  assign n34914 = \m4_addr_i[12]_pad  & n1925 ;
  assign n34915 = n1918 & n34914 ;
  assign n34916 = \m3_addr_i[12]_pad  & n1910 ;
  assign n34917 = n1938 & n34916 ;
  assign n34918 = ~n34915 & ~n34917 ;
  assign n34919 = \m1_addr_i[12]_pad  & n1910 ;
  assign n34920 = n1941 & n34919 ;
  assign n34921 = \m0_addr_i[12]_pad  & n1925 ;
  assign n34922 = n1931 & n34921 ;
  assign n34923 = ~n34920 & ~n34922 ;
  assign n34924 = n34918 & n34923 ;
  assign n34925 = n34913 & n34924 ;
  assign n34926 = \m7_addr_i[13]_pad  & ~n1910 ;
  assign n34927 = n1938 & n34926 ;
  assign n34928 = \m6_addr_i[13]_pad  & ~n1925 ;
  assign n34929 = n1918 & n34928 ;
  assign n34930 = ~n34927 & ~n34929 ;
  assign n34931 = \m5_addr_i[13]_pad  & ~n1910 ;
  assign n34932 = n1941 & n34931 ;
  assign n34933 = \m2_addr_i[13]_pad  & ~n1925 ;
  assign n34934 = n1931 & n34933 ;
  assign n34935 = ~n34932 & ~n34934 ;
  assign n34936 = n34930 & n34935 ;
  assign n34937 = \m4_addr_i[13]_pad  & n1925 ;
  assign n34938 = n1918 & n34937 ;
  assign n34939 = \m3_addr_i[13]_pad  & n1910 ;
  assign n34940 = n1938 & n34939 ;
  assign n34941 = ~n34938 & ~n34940 ;
  assign n34942 = \m1_addr_i[13]_pad  & n1910 ;
  assign n34943 = n1941 & n34942 ;
  assign n34944 = \m0_addr_i[13]_pad  & n1925 ;
  assign n34945 = n1931 & n34944 ;
  assign n34946 = ~n34943 & ~n34945 ;
  assign n34947 = n34941 & n34946 ;
  assign n34948 = n34936 & n34947 ;
  assign n34949 = \m7_addr_i[14]_pad  & ~n1910 ;
  assign n34950 = n1938 & n34949 ;
  assign n34951 = \m6_addr_i[14]_pad  & ~n1925 ;
  assign n34952 = n1918 & n34951 ;
  assign n34953 = ~n34950 & ~n34952 ;
  assign n34954 = \m5_addr_i[14]_pad  & ~n1910 ;
  assign n34955 = n1941 & n34954 ;
  assign n34956 = \m2_addr_i[14]_pad  & ~n1925 ;
  assign n34957 = n1931 & n34956 ;
  assign n34958 = ~n34955 & ~n34957 ;
  assign n34959 = n34953 & n34958 ;
  assign n34960 = \m4_addr_i[14]_pad  & n1925 ;
  assign n34961 = n1918 & n34960 ;
  assign n34962 = \m3_addr_i[14]_pad  & n1910 ;
  assign n34963 = n1938 & n34962 ;
  assign n34964 = ~n34961 & ~n34963 ;
  assign n34965 = \m1_addr_i[14]_pad  & n1910 ;
  assign n34966 = n1941 & n34965 ;
  assign n34967 = \m0_addr_i[14]_pad  & n1925 ;
  assign n34968 = n1931 & n34967 ;
  assign n34969 = ~n34966 & ~n34968 ;
  assign n34970 = n34964 & n34969 ;
  assign n34971 = n34959 & n34970 ;
  assign n34972 = \m3_addr_i[15]_pad  & n1910 ;
  assign n34973 = n1938 & n34972 ;
  assign n34974 = \m2_addr_i[15]_pad  & ~n1925 ;
  assign n34975 = n1931 & n34974 ;
  assign n34976 = ~n34973 & ~n34975 ;
  assign n34977 = \m5_addr_i[15]_pad  & ~n1910 ;
  assign n34978 = n1941 & n34977 ;
  assign n34979 = \m0_addr_i[15]_pad  & n1925 ;
  assign n34980 = n1931 & n34979 ;
  assign n34981 = ~n34978 & ~n34980 ;
  assign n34982 = n34976 & n34981 ;
  assign n34983 = \m4_addr_i[15]_pad  & n1925 ;
  assign n34984 = n1918 & n34983 ;
  assign n34985 = \m1_addr_i[15]_pad  & n1910 ;
  assign n34986 = n1941 & n34985 ;
  assign n34987 = ~n34984 & ~n34986 ;
  assign n34988 = \m7_addr_i[15]_pad  & ~n1910 ;
  assign n34989 = n1938 & n34988 ;
  assign n34990 = \m6_addr_i[15]_pad  & ~n1925 ;
  assign n34991 = n1918 & n34990 ;
  assign n34992 = ~n34989 & ~n34991 ;
  assign n34993 = n34987 & n34992 ;
  assign n34994 = n34982 & n34993 ;
  assign n34995 = \m7_addr_i[16]_pad  & ~n1910 ;
  assign n34996 = n1938 & n34995 ;
  assign n34997 = \m6_addr_i[16]_pad  & ~n1925 ;
  assign n34998 = n1918 & n34997 ;
  assign n34999 = ~n34996 & ~n34998 ;
  assign n35000 = \m5_addr_i[16]_pad  & ~n1910 ;
  assign n35001 = n1941 & n35000 ;
  assign n35002 = \m2_addr_i[16]_pad  & ~n1925 ;
  assign n35003 = n1931 & n35002 ;
  assign n35004 = ~n35001 & ~n35003 ;
  assign n35005 = n34999 & n35004 ;
  assign n35006 = \m4_addr_i[16]_pad  & n1925 ;
  assign n35007 = n1918 & n35006 ;
  assign n35008 = \m3_addr_i[16]_pad  & n1910 ;
  assign n35009 = n1938 & n35008 ;
  assign n35010 = ~n35007 & ~n35009 ;
  assign n35011 = \m1_addr_i[16]_pad  & n1910 ;
  assign n35012 = n1941 & n35011 ;
  assign n35013 = \m0_addr_i[16]_pad  & n1925 ;
  assign n35014 = n1931 & n35013 ;
  assign n35015 = ~n35012 & ~n35014 ;
  assign n35016 = n35010 & n35015 ;
  assign n35017 = n35005 & n35016 ;
  assign n35018 = \m5_addr_i[17]_pad  & ~n1910 ;
  assign n35019 = n1941 & n35018 ;
  assign n35020 = \m4_addr_i[17]_pad  & n1925 ;
  assign n35021 = n1918 & n35020 ;
  assign n35022 = ~n35019 & ~n35021 ;
  assign n35023 = \m7_addr_i[17]_pad  & ~n1910 ;
  assign n35024 = n1938 & n35023 ;
  assign n35025 = \m2_addr_i[17]_pad  & ~n1925 ;
  assign n35026 = n1931 & n35025 ;
  assign n35027 = ~n35024 & ~n35026 ;
  assign n35028 = n35022 & n35027 ;
  assign n35029 = \m6_addr_i[17]_pad  & ~n1925 ;
  assign n35030 = n1918 & n35029 ;
  assign n35031 = \m3_addr_i[17]_pad  & n1910 ;
  assign n35032 = n1938 & n35031 ;
  assign n35033 = ~n35030 & ~n35032 ;
  assign n35034 = \m1_addr_i[17]_pad  & n1910 ;
  assign n35035 = n1941 & n35034 ;
  assign n35036 = \m0_addr_i[17]_pad  & n1925 ;
  assign n35037 = n1931 & n35036 ;
  assign n35038 = ~n35035 & ~n35037 ;
  assign n35039 = n35033 & n35038 ;
  assign n35040 = n35028 & n35039 ;
  assign n35041 = \m7_addr_i[18]_pad  & ~n1910 ;
  assign n35042 = n1938 & n35041 ;
  assign n35043 = \m6_addr_i[18]_pad  & ~n1925 ;
  assign n35044 = n1918 & n35043 ;
  assign n35045 = ~n35042 & ~n35044 ;
  assign n35046 = \m5_addr_i[18]_pad  & ~n1910 ;
  assign n35047 = n1941 & n35046 ;
  assign n35048 = \m2_addr_i[18]_pad  & ~n1925 ;
  assign n35049 = n1931 & n35048 ;
  assign n35050 = ~n35047 & ~n35049 ;
  assign n35051 = n35045 & n35050 ;
  assign n35052 = \m4_addr_i[18]_pad  & n1925 ;
  assign n35053 = n1918 & n35052 ;
  assign n35054 = \m3_addr_i[18]_pad  & n1910 ;
  assign n35055 = n1938 & n35054 ;
  assign n35056 = ~n35053 & ~n35055 ;
  assign n35057 = \m1_addr_i[18]_pad  & n1910 ;
  assign n35058 = n1941 & n35057 ;
  assign n35059 = \m0_addr_i[18]_pad  & n1925 ;
  assign n35060 = n1931 & n35059 ;
  assign n35061 = ~n35058 & ~n35060 ;
  assign n35062 = n35056 & n35061 ;
  assign n35063 = n35051 & n35062 ;
  assign n35064 = \m7_addr_i[19]_pad  & ~n1910 ;
  assign n35065 = n1938 & n35064 ;
  assign n35066 = \m6_addr_i[19]_pad  & ~n1925 ;
  assign n35067 = n1918 & n35066 ;
  assign n35068 = ~n35065 & ~n35067 ;
  assign n35069 = \m5_addr_i[19]_pad  & ~n1910 ;
  assign n35070 = n1941 & n35069 ;
  assign n35071 = \m2_addr_i[19]_pad  & ~n1925 ;
  assign n35072 = n1931 & n35071 ;
  assign n35073 = ~n35070 & ~n35072 ;
  assign n35074 = n35068 & n35073 ;
  assign n35075 = \m4_addr_i[19]_pad  & n1925 ;
  assign n35076 = n1918 & n35075 ;
  assign n35077 = \m3_addr_i[19]_pad  & n1910 ;
  assign n35078 = n1938 & n35077 ;
  assign n35079 = ~n35076 & ~n35078 ;
  assign n35080 = \m1_addr_i[19]_pad  & n1910 ;
  assign n35081 = n1941 & n35080 ;
  assign n35082 = \m0_addr_i[19]_pad  & n1925 ;
  assign n35083 = n1931 & n35082 ;
  assign n35084 = ~n35081 & ~n35083 ;
  assign n35085 = n35079 & n35084 ;
  assign n35086 = n35074 & n35085 ;
  assign n35087 = \m7_addr_i[1]_pad  & ~n1910 ;
  assign n35088 = n1938 & n35087 ;
  assign n35089 = \m6_addr_i[1]_pad  & ~n1925 ;
  assign n35090 = n1918 & n35089 ;
  assign n35091 = ~n35088 & ~n35090 ;
  assign n35092 = \m5_addr_i[1]_pad  & ~n1910 ;
  assign n35093 = n1941 & n35092 ;
  assign n35094 = \m2_addr_i[1]_pad  & ~n1925 ;
  assign n35095 = n1931 & n35094 ;
  assign n35096 = ~n35093 & ~n35095 ;
  assign n35097 = n35091 & n35096 ;
  assign n35098 = \m4_addr_i[1]_pad  & n1925 ;
  assign n35099 = n1918 & n35098 ;
  assign n35100 = \m3_addr_i[1]_pad  & n1910 ;
  assign n35101 = n1938 & n35100 ;
  assign n35102 = ~n35099 & ~n35101 ;
  assign n35103 = \m1_addr_i[1]_pad  & n1910 ;
  assign n35104 = n1941 & n35103 ;
  assign n35105 = \m0_addr_i[1]_pad  & n1925 ;
  assign n35106 = n1931 & n35105 ;
  assign n35107 = ~n35104 & ~n35106 ;
  assign n35108 = n35102 & n35107 ;
  assign n35109 = n35097 & n35108 ;
  assign n35110 = \m7_addr_i[20]_pad  & ~n1910 ;
  assign n35111 = n1938 & n35110 ;
  assign n35112 = \m6_addr_i[20]_pad  & ~n1925 ;
  assign n35113 = n1918 & n35112 ;
  assign n35114 = ~n35111 & ~n35113 ;
  assign n35115 = \m5_addr_i[20]_pad  & ~n1910 ;
  assign n35116 = n1941 & n35115 ;
  assign n35117 = \m2_addr_i[20]_pad  & ~n1925 ;
  assign n35118 = n1931 & n35117 ;
  assign n35119 = ~n35116 & ~n35118 ;
  assign n35120 = n35114 & n35119 ;
  assign n35121 = \m4_addr_i[20]_pad  & n1925 ;
  assign n35122 = n1918 & n35121 ;
  assign n35123 = \m3_addr_i[20]_pad  & n1910 ;
  assign n35124 = n1938 & n35123 ;
  assign n35125 = ~n35122 & ~n35124 ;
  assign n35126 = \m1_addr_i[20]_pad  & n1910 ;
  assign n35127 = n1941 & n35126 ;
  assign n35128 = \m0_addr_i[20]_pad  & n1925 ;
  assign n35129 = n1931 & n35128 ;
  assign n35130 = ~n35127 & ~n35129 ;
  assign n35131 = n35125 & n35130 ;
  assign n35132 = n35120 & n35131 ;
  assign n35133 = \m3_addr_i[21]_pad  & n1910 ;
  assign n35134 = n1938 & n35133 ;
  assign n35135 = \m2_addr_i[21]_pad  & ~n1925 ;
  assign n35136 = n1931 & n35135 ;
  assign n35137 = ~n35134 & ~n35136 ;
  assign n35138 = \m5_addr_i[21]_pad  & ~n1910 ;
  assign n35139 = n1941 & n35138 ;
  assign n35140 = \m0_addr_i[21]_pad  & n1925 ;
  assign n35141 = n1931 & n35140 ;
  assign n35142 = ~n35139 & ~n35141 ;
  assign n35143 = n35137 & n35142 ;
  assign n35144 = \m4_addr_i[21]_pad  & n1925 ;
  assign n35145 = n1918 & n35144 ;
  assign n35146 = \m1_addr_i[21]_pad  & n1910 ;
  assign n35147 = n1941 & n35146 ;
  assign n35148 = ~n35145 & ~n35147 ;
  assign n35149 = \m7_addr_i[21]_pad  & ~n1910 ;
  assign n35150 = n1938 & n35149 ;
  assign n35151 = \m6_addr_i[21]_pad  & ~n1925 ;
  assign n35152 = n1918 & n35151 ;
  assign n35153 = ~n35150 & ~n35152 ;
  assign n35154 = n35148 & n35153 ;
  assign n35155 = n35143 & n35154 ;
  assign n35156 = \m7_addr_i[22]_pad  & ~n1910 ;
  assign n35157 = n1938 & n35156 ;
  assign n35158 = \m6_addr_i[22]_pad  & ~n1925 ;
  assign n35159 = n1918 & n35158 ;
  assign n35160 = ~n35157 & ~n35159 ;
  assign n35161 = \m5_addr_i[22]_pad  & ~n1910 ;
  assign n35162 = n1941 & n35161 ;
  assign n35163 = \m2_addr_i[22]_pad  & ~n1925 ;
  assign n35164 = n1931 & n35163 ;
  assign n35165 = ~n35162 & ~n35164 ;
  assign n35166 = n35160 & n35165 ;
  assign n35167 = \m4_addr_i[22]_pad  & n1925 ;
  assign n35168 = n1918 & n35167 ;
  assign n35169 = \m3_addr_i[22]_pad  & n1910 ;
  assign n35170 = n1938 & n35169 ;
  assign n35171 = ~n35168 & ~n35170 ;
  assign n35172 = \m1_addr_i[22]_pad  & n1910 ;
  assign n35173 = n1941 & n35172 ;
  assign n35174 = \m0_addr_i[22]_pad  & n1925 ;
  assign n35175 = n1931 & n35174 ;
  assign n35176 = ~n35173 & ~n35175 ;
  assign n35177 = n35171 & n35176 ;
  assign n35178 = n35166 & n35177 ;
  assign n35179 = \m7_addr_i[23]_pad  & ~n1910 ;
  assign n35180 = n1938 & n35179 ;
  assign n35181 = \m6_addr_i[23]_pad  & ~n1925 ;
  assign n35182 = n1918 & n35181 ;
  assign n35183 = ~n35180 & ~n35182 ;
  assign n35184 = \m5_addr_i[23]_pad  & ~n1910 ;
  assign n35185 = n1941 & n35184 ;
  assign n35186 = \m2_addr_i[23]_pad  & ~n1925 ;
  assign n35187 = n1931 & n35186 ;
  assign n35188 = ~n35185 & ~n35187 ;
  assign n35189 = n35183 & n35188 ;
  assign n35190 = \m4_addr_i[23]_pad  & n1925 ;
  assign n35191 = n1918 & n35190 ;
  assign n35192 = \m3_addr_i[23]_pad  & n1910 ;
  assign n35193 = n1938 & n35192 ;
  assign n35194 = ~n35191 & ~n35193 ;
  assign n35195 = \m1_addr_i[23]_pad  & n1910 ;
  assign n35196 = n1941 & n35195 ;
  assign n35197 = \m0_addr_i[23]_pad  & n1925 ;
  assign n35198 = n1931 & n35197 ;
  assign n35199 = ~n35196 & ~n35198 ;
  assign n35200 = n35194 & n35199 ;
  assign n35201 = n35189 & n35200 ;
  assign n35202 = \m4_addr_i[28]_pad  & n1925 ;
  assign n35203 = n1918 & n35202 ;
  assign n35204 = \m3_addr_i[28]_pad  & n1910 ;
  assign n35205 = n1938 & n35204 ;
  assign n35206 = ~n35203 & ~n35205 ;
  assign n35207 = \m1_addr_i[28]_pad  & n1910 ;
  assign n35208 = n1941 & n35207 ;
  assign n35209 = \m6_addr_i[28]_pad  & ~n1925 ;
  assign n35210 = n1918 & n35209 ;
  assign n35211 = ~n35208 & ~n35210 ;
  assign n35212 = n35206 & n35211 ;
  assign n35213 = \m2_addr_i[28]_pad  & ~n1925 ;
  assign n35214 = n1931 & n35213 ;
  assign n35215 = \m5_addr_i[28]_pad  & ~n1910 ;
  assign n35216 = n1941 & n35215 ;
  assign n35217 = ~n35214 & ~n35216 ;
  assign n35218 = \m0_addr_i[28]_pad  & n1925 ;
  assign n35219 = n1931 & n35218 ;
  assign n35220 = \m7_addr_i[28]_pad  & ~n1910 ;
  assign n35221 = n1938 & n35220 ;
  assign n35222 = ~n35219 & ~n35221 ;
  assign n35223 = n35217 & n35222 ;
  assign n35224 = n35212 & n35223 ;
  assign n35225 = \m1_addr_i[29]_pad  & n1910 ;
  assign n35226 = n1941 & n35225 ;
  assign n35227 = \m2_addr_i[29]_pad  & ~n1925 ;
  assign n35228 = n1931 & n35227 ;
  assign n35229 = ~n35226 & ~n35228 ;
  assign n35230 = \m0_addr_i[29]_pad  & n1925 ;
  assign n35231 = n1931 & n35230 ;
  assign n35232 = \m3_addr_i[29]_pad  & n1910 ;
  assign n35233 = n1938 & n35232 ;
  assign n35234 = ~n35231 & ~n35233 ;
  assign n35235 = n35229 & n35234 ;
  assign n35236 = \m7_addr_i[29]_pad  & ~n1910 ;
  assign n35237 = n1938 & n35236 ;
  assign n35238 = \m4_addr_i[29]_pad  & n1925 ;
  assign n35239 = n1918 & n35238 ;
  assign n35240 = ~n35237 & ~n35239 ;
  assign n35241 = \m5_addr_i[29]_pad  & ~n1910 ;
  assign n35242 = n1941 & n35241 ;
  assign n35243 = \m6_addr_i[29]_pad  & ~n1925 ;
  assign n35244 = n1918 & n35243 ;
  assign n35245 = ~n35242 & ~n35244 ;
  assign n35246 = n35240 & n35245 ;
  assign n35247 = n35235 & n35246 ;
  assign n35248 = \m4_addr_i[30]_pad  & n1925 ;
  assign n35249 = n1918 & n35248 ;
  assign n35250 = \m3_addr_i[30]_pad  & n1910 ;
  assign n35251 = n1938 & n35250 ;
  assign n35252 = ~n35249 & ~n35251 ;
  assign n35253 = \m1_addr_i[30]_pad  & n1910 ;
  assign n35254 = n1941 & n35253 ;
  assign n35255 = \m6_addr_i[30]_pad  & ~n1925 ;
  assign n35256 = n1918 & n35255 ;
  assign n35257 = ~n35254 & ~n35256 ;
  assign n35258 = n35252 & n35257 ;
  assign n35259 = \m2_addr_i[30]_pad  & ~n1925 ;
  assign n35260 = n1931 & n35259 ;
  assign n35261 = \m5_addr_i[30]_pad  & ~n1910 ;
  assign n35262 = n1941 & n35261 ;
  assign n35263 = ~n35260 & ~n35262 ;
  assign n35264 = \m0_addr_i[30]_pad  & n1925 ;
  assign n35265 = n1931 & n35264 ;
  assign n35266 = \m7_addr_i[30]_pad  & ~n1910 ;
  assign n35267 = n1938 & n35266 ;
  assign n35268 = ~n35265 & ~n35267 ;
  assign n35269 = n35263 & n35268 ;
  assign n35270 = n35258 & n35269 ;
  assign n35271 = \m4_addr_i[31]_pad  & n1925 ;
  assign n35272 = n1918 & n35271 ;
  assign n35273 = \m3_addr_i[31]_pad  & n1910 ;
  assign n35274 = n1938 & n35273 ;
  assign n35275 = ~n35272 & ~n35274 ;
  assign n35276 = \m1_addr_i[31]_pad  & n1910 ;
  assign n35277 = n1941 & n35276 ;
  assign n35278 = \m6_addr_i[31]_pad  & ~n1925 ;
  assign n35279 = n1918 & n35278 ;
  assign n35280 = ~n35277 & ~n35279 ;
  assign n35281 = n35275 & n35280 ;
  assign n35282 = \m2_addr_i[31]_pad  & ~n1925 ;
  assign n35283 = n1931 & n35282 ;
  assign n35284 = \m5_addr_i[31]_pad  & ~n1910 ;
  assign n35285 = n1941 & n35284 ;
  assign n35286 = ~n35283 & ~n35285 ;
  assign n35287 = \m0_addr_i[31]_pad  & n1925 ;
  assign n35288 = n1931 & n35287 ;
  assign n35289 = \m7_addr_i[31]_pad  & ~n1910 ;
  assign n35290 = n1938 & n35289 ;
  assign n35291 = ~n35288 & ~n35290 ;
  assign n35292 = n35286 & n35291 ;
  assign n35293 = n35281 & n35292 ;
  assign n35294 = \m7_addr_i[6]_pad  & ~n1910 ;
  assign n35295 = n1938 & n35294 ;
  assign n35296 = \m6_addr_i[6]_pad  & ~n1925 ;
  assign n35297 = n1918 & n35296 ;
  assign n35298 = ~n35295 & ~n35297 ;
  assign n35299 = \m5_addr_i[6]_pad  & ~n1910 ;
  assign n35300 = n1941 & n35299 ;
  assign n35301 = \m2_addr_i[6]_pad  & ~n1925 ;
  assign n35302 = n1931 & n35301 ;
  assign n35303 = ~n35300 & ~n35302 ;
  assign n35304 = n35298 & n35303 ;
  assign n35305 = \m4_addr_i[6]_pad  & n1925 ;
  assign n35306 = n1918 & n35305 ;
  assign n35307 = \m3_addr_i[6]_pad  & n1910 ;
  assign n35308 = n1938 & n35307 ;
  assign n35309 = ~n35306 & ~n35308 ;
  assign n35310 = \m1_addr_i[6]_pad  & n1910 ;
  assign n35311 = n1941 & n35310 ;
  assign n35312 = \m0_addr_i[6]_pad  & n1925 ;
  assign n35313 = n1931 & n35312 ;
  assign n35314 = ~n35311 & ~n35313 ;
  assign n35315 = n35309 & n35314 ;
  assign n35316 = n35304 & n35315 ;
  assign n35317 = \m7_addr_i[7]_pad  & ~n1910 ;
  assign n35318 = n1938 & n35317 ;
  assign n35319 = \m6_addr_i[7]_pad  & ~n1925 ;
  assign n35320 = n1918 & n35319 ;
  assign n35321 = ~n35318 & ~n35320 ;
  assign n35322 = \m5_addr_i[7]_pad  & ~n1910 ;
  assign n35323 = n1941 & n35322 ;
  assign n35324 = \m2_addr_i[7]_pad  & ~n1925 ;
  assign n35325 = n1931 & n35324 ;
  assign n35326 = ~n35323 & ~n35325 ;
  assign n35327 = n35321 & n35326 ;
  assign n35328 = \m4_addr_i[7]_pad  & n1925 ;
  assign n35329 = n1918 & n35328 ;
  assign n35330 = \m3_addr_i[7]_pad  & n1910 ;
  assign n35331 = n1938 & n35330 ;
  assign n35332 = ~n35329 & ~n35331 ;
  assign n35333 = \m1_addr_i[7]_pad  & n1910 ;
  assign n35334 = n1941 & n35333 ;
  assign n35335 = \m0_addr_i[7]_pad  & n1925 ;
  assign n35336 = n1931 & n35335 ;
  assign n35337 = ~n35334 & ~n35336 ;
  assign n35338 = n35332 & n35337 ;
  assign n35339 = n35327 & n35338 ;
  assign n35340 = \m7_addr_i[8]_pad  & ~n1910 ;
  assign n35341 = n1938 & n35340 ;
  assign n35342 = \m6_addr_i[8]_pad  & ~n1925 ;
  assign n35343 = n1918 & n35342 ;
  assign n35344 = ~n35341 & ~n35343 ;
  assign n35345 = \m5_addr_i[8]_pad  & ~n1910 ;
  assign n35346 = n1941 & n35345 ;
  assign n35347 = \m2_addr_i[8]_pad  & ~n1925 ;
  assign n35348 = n1931 & n35347 ;
  assign n35349 = ~n35346 & ~n35348 ;
  assign n35350 = n35344 & n35349 ;
  assign n35351 = \m4_addr_i[8]_pad  & n1925 ;
  assign n35352 = n1918 & n35351 ;
  assign n35353 = \m3_addr_i[8]_pad  & n1910 ;
  assign n35354 = n1938 & n35353 ;
  assign n35355 = ~n35352 & ~n35354 ;
  assign n35356 = \m1_addr_i[8]_pad  & n1910 ;
  assign n35357 = n1941 & n35356 ;
  assign n35358 = \m0_addr_i[8]_pad  & n1925 ;
  assign n35359 = n1931 & n35358 ;
  assign n35360 = ~n35357 & ~n35359 ;
  assign n35361 = n35355 & n35360 ;
  assign n35362 = n35350 & n35361 ;
  assign n35363 = \m3_addr_i[9]_pad  & n1910 ;
  assign n35364 = n1938 & n35363 ;
  assign n35365 = \m2_addr_i[9]_pad  & ~n1925 ;
  assign n35366 = n1931 & n35365 ;
  assign n35367 = ~n35364 & ~n35366 ;
  assign n35368 = \m5_addr_i[9]_pad  & ~n1910 ;
  assign n35369 = n1941 & n35368 ;
  assign n35370 = \m0_addr_i[9]_pad  & n1925 ;
  assign n35371 = n1931 & n35370 ;
  assign n35372 = ~n35369 & ~n35371 ;
  assign n35373 = n35367 & n35372 ;
  assign n35374 = \m4_addr_i[9]_pad  & n1925 ;
  assign n35375 = n1918 & n35374 ;
  assign n35376 = \m1_addr_i[9]_pad  & n1910 ;
  assign n35377 = n1941 & n35376 ;
  assign n35378 = ~n35375 & ~n35377 ;
  assign n35379 = \m7_addr_i[9]_pad  & ~n1910 ;
  assign n35380 = n1938 & n35379 ;
  assign n35381 = \m6_addr_i[9]_pad  & ~n1925 ;
  assign n35382 = n1918 & n35381 ;
  assign n35383 = ~n35380 & ~n35382 ;
  assign n35384 = n35378 & n35383 ;
  assign n35385 = n35373 & n35384 ;
  assign n35386 = ~n2106 & ~n2258 ;
  assign n35387 = \m7_data_i[16]_pad  & ~n1910 ;
  assign n35388 = n1938 & n35387 ;
  assign n35389 = \m6_data_i[16]_pad  & ~n1925 ;
  assign n35390 = n1918 & n35389 ;
  assign n35391 = ~n35388 & ~n35390 ;
  assign n35392 = \m5_data_i[16]_pad  & ~n1910 ;
  assign n35393 = n1941 & n35392 ;
  assign n35394 = \m2_data_i[16]_pad  & ~n1925 ;
  assign n35395 = n1931 & n35394 ;
  assign n35396 = ~n35393 & ~n35395 ;
  assign n35397 = n35391 & n35396 ;
  assign n35398 = \m4_data_i[16]_pad  & n1925 ;
  assign n35399 = n1918 & n35398 ;
  assign n35400 = \m3_data_i[16]_pad  & n1910 ;
  assign n35401 = n1938 & n35400 ;
  assign n35402 = ~n35399 & ~n35401 ;
  assign n35403 = \m1_data_i[16]_pad  & n1910 ;
  assign n35404 = n1941 & n35403 ;
  assign n35405 = \m0_data_i[16]_pad  & n1925 ;
  assign n35406 = n1931 & n35405 ;
  assign n35407 = ~n35404 & ~n35406 ;
  assign n35408 = n35402 & n35407 ;
  assign n35409 = n35397 & n35408 ;
  assign n35410 = \m7_data_i[17]_pad  & ~n1910 ;
  assign n35411 = n1938 & n35410 ;
  assign n35412 = \m6_data_i[17]_pad  & ~n1925 ;
  assign n35413 = n1918 & n35412 ;
  assign n35414 = ~n35411 & ~n35413 ;
  assign n35415 = \m5_data_i[17]_pad  & ~n1910 ;
  assign n35416 = n1941 & n35415 ;
  assign n35417 = \m0_data_i[17]_pad  & n1925 ;
  assign n35418 = n1931 & n35417 ;
  assign n35419 = ~n35416 & ~n35418 ;
  assign n35420 = n35414 & n35419 ;
  assign n35421 = \m4_data_i[17]_pad  & n1925 ;
  assign n35422 = n1918 & n35421 ;
  assign n35423 = \m1_data_i[17]_pad  & n1910 ;
  assign n35424 = n1941 & n35423 ;
  assign n35425 = ~n35422 & ~n35424 ;
  assign n35426 = \m3_data_i[17]_pad  & n1910 ;
  assign n35427 = n1938 & n35426 ;
  assign n35428 = \m2_data_i[17]_pad  & ~n1925 ;
  assign n35429 = n1931 & n35428 ;
  assign n35430 = ~n35427 & ~n35429 ;
  assign n35431 = n35425 & n35430 ;
  assign n35432 = n35420 & n35431 ;
  assign n35433 = \m7_data_i[18]_pad  & ~n1910 ;
  assign n35434 = n1938 & n35433 ;
  assign n35435 = \m6_data_i[18]_pad  & ~n1925 ;
  assign n35436 = n1918 & n35435 ;
  assign n35437 = ~n35434 & ~n35436 ;
  assign n35438 = \m5_data_i[18]_pad  & ~n1910 ;
  assign n35439 = n1941 & n35438 ;
  assign n35440 = \m2_data_i[18]_pad  & ~n1925 ;
  assign n35441 = n1931 & n35440 ;
  assign n35442 = ~n35439 & ~n35441 ;
  assign n35443 = n35437 & n35442 ;
  assign n35444 = \m4_data_i[18]_pad  & n1925 ;
  assign n35445 = n1918 & n35444 ;
  assign n35446 = \m3_data_i[18]_pad  & n1910 ;
  assign n35447 = n1938 & n35446 ;
  assign n35448 = ~n35445 & ~n35447 ;
  assign n35449 = \m1_data_i[18]_pad  & n1910 ;
  assign n35450 = n1941 & n35449 ;
  assign n35451 = \m0_data_i[18]_pad  & n1925 ;
  assign n35452 = n1931 & n35451 ;
  assign n35453 = ~n35450 & ~n35452 ;
  assign n35454 = n35448 & n35453 ;
  assign n35455 = n35443 & n35454 ;
  assign n35456 = \m5_data_i[19]_pad  & ~n1910 ;
  assign n35457 = n1941 & n35456 ;
  assign n35458 = \m4_data_i[19]_pad  & n1925 ;
  assign n35459 = n1918 & n35458 ;
  assign n35460 = ~n35457 & ~n35459 ;
  assign n35461 = \m7_data_i[19]_pad  & ~n1910 ;
  assign n35462 = n1938 & n35461 ;
  assign n35463 = \m2_data_i[19]_pad  & ~n1925 ;
  assign n35464 = n1931 & n35463 ;
  assign n35465 = ~n35462 & ~n35464 ;
  assign n35466 = n35460 & n35465 ;
  assign n35467 = \m6_data_i[19]_pad  & ~n1925 ;
  assign n35468 = n1918 & n35467 ;
  assign n35469 = \m3_data_i[19]_pad  & n1910 ;
  assign n35470 = n1938 & n35469 ;
  assign n35471 = ~n35468 & ~n35470 ;
  assign n35472 = \m1_data_i[19]_pad  & n1910 ;
  assign n35473 = n1941 & n35472 ;
  assign n35474 = \m0_data_i[19]_pad  & n1925 ;
  assign n35475 = n1931 & n35474 ;
  assign n35476 = ~n35473 & ~n35475 ;
  assign n35477 = n35471 & n35476 ;
  assign n35478 = n35466 & n35477 ;
  assign n35479 = \m7_data_i[20]_pad  & ~n1910 ;
  assign n35480 = n1938 & n35479 ;
  assign n35481 = \m6_data_i[20]_pad  & ~n1925 ;
  assign n35482 = n1918 & n35481 ;
  assign n35483 = ~n35480 & ~n35482 ;
  assign n35484 = \m5_data_i[20]_pad  & ~n1910 ;
  assign n35485 = n1941 & n35484 ;
  assign n35486 = \m2_data_i[20]_pad  & ~n1925 ;
  assign n35487 = n1931 & n35486 ;
  assign n35488 = ~n35485 & ~n35487 ;
  assign n35489 = n35483 & n35488 ;
  assign n35490 = \m4_data_i[20]_pad  & n1925 ;
  assign n35491 = n1918 & n35490 ;
  assign n35492 = \m3_data_i[20]_pad  & n1910 ;
  assign n35493 = n1938 & n35492 ;
  assign n35494 = ~n35491 & ~n35493 ;
  assign n35495 = \m1_data_i[20]_pad  & n1910 ;
  assign n35496 = n1941 & n35495 ;
  assign n35497 = \m0_data_i[20]_pad  & n1925 ;
  assign n35498 = n1931 & n35497 ;
  assign n35499 = ~n35496 & ~n35498 ;
  assign n35500 = n35494 & n35499 ;
  assign n35501 = n35489 & n35500 ;
  assign n35502 = \m5_data_i[21]_pad  & ~n1910 ;
  assign n35503 = n1941 & n35502 ;
  assign n35504 = \m4_data_i[21]_pad  & n1925 ;
  assign n35505 = n1918 & n35504 ;
  assign n35506 = ~n35503 & ~n35505 ;
  assign n35507 = \m7_data_i[21]_pad  & ~n1910 ;
  assign n35508 = n1938 & n35507 ;
  assign n35509 = \m2_data_i[21]_pad  & ~n1925 ;
  assign n35510 = n1931 & n35509 ;
  assign n35511 = ~n35508 & ~n35510 ;
  assign n35512 = n35506 & n35511 ;
  assign n35513 = \m6_data_i[21]_pad  & ~n1925 ;
  assign n35514 = n1918 & n35513 ;
  assign n35515 = \m3_data_i[21]_pad  & n1910 ;
  assign n35516 = n1938 & n35515 ;
  assign n35517 = ~n35514 & ~n35516 ;
  assign n35518 = \m1_data_i[21]_pad  & n1910 ;
  assign n35519 = n1941 & n35518 ;
  assign n35520 = \m0_data_i[21]_pad  & n1925 ;
  assign n35521 = n1931 & n35520 ;
  assign n35522 = ~n35519 & ~n35521 ;
  assign n35523 = n35517 & n35522 ;
  assign n35524 = n35512 & n35523 ;
  assign n35525 = \m7_data_i[22]_pad  & ~n1910 ;
  assign n35526 = n1938 & n35525 ;
  assign n35527 = \m6_data_i[22]_pad  & ~n1925 ;
  assign n35528 = n1918 & n35527 ;
  assign n35529 = ~n35526 & ~n35528 ;
  assign n35530 = \m5_data_i[22]_pad  & ~n1910 ;
  assign n35531 = n1941 & n35530 ;
  assign n35532 = \m2_data_i[22]_pad  & ~n1925 ;
  assign n35533 = n1931 & n35532 ;
  assign n35534 = ~n35531 & ~n35533 ;
  assign n35535 = n35529 & n35534 ;
  assign n35536 = \m4_data_i[22]_pad  & n1925 ;
  assign n35537 = n1918 & n35536 ;
  assign n35538 = \m3_data_i[22]_pad  & n1910 ;
  assign n35539 = n1938 & n35538 ;
  assign n35540 = ~n35537 & ~n35539 ;
  assign n35541 = \m1_data_i[22]_pad  & n1910 ;
  assign n35542 = n1941 & n35541 ;
  assign n35543 = \m0_data_i[22]_pad  & n1925 ;
  assign n35544 = n1931 & n35543 ;
  assign n35545 = ~n35542 & ~n35544 ;
  assign n35546 = n35540 & n35545 ;
  assign n35547 = n35535 & n35546 ;
  assign n35548 = \m7_data_i[23]_pad  & ~n1910 ;
  assign n35549 = n1938 & n35548 ;
  assign n35550 = \m6_data_i[23]_pad  & ~n1925 ;
  assign n35551 = n1918 & n35550 ;
  assign n35552 = ~n35549 & ~n35551 ;
  assign n35553 = \m5_data_i[23]_pad  & ~n1910 ;
  assign n35554 = n1941 & n35553 ;
  assign n35555 = \m2_data_i[23]_pad  & ~n1925 ;
  assign n35556 = n1931 & n35555 ;
  assign n35557 = ~n35554 & ~n35556 ;
  assign n35558 = n35552 & n35557 ;
  assign n35559 = \m4_data_i[23]_pad  & n1925 ;
  assign n35560 = n1918 & n35559 ;
  assign n35561 = \m3_data_i[23]_pad  & n1910 ;
  assign n35562 = n1938 & n35561 ;
  assign n35563 = ~n35560 & ~n35562 ;
  assign n35564 = \m1_data_i[23]_pad  & n1910 ;
  assign n35565 = n1941 & n35564 ;
  assign n35566 = \m0_data_i[23]_pad  & n1925 ;
  assign n35567 = n1931 & n35566 ;
  assign n35568 = ~n35565 & ~n35567 ;
  assign n35569 = n35563 & n35568 ;
  assign n35570 = n35558 & n35569 ;
  assign n35571 = \m7_data_i[24]_pad  & ~n1910 ;
  assign n35572 = n1938 & n35571 ;
  assign n35573 = \m6_data_i[24]_pad  & ~n1925 ;
  assign n35574 = n1918 & n35573 ;
  assign n35575 = ~n35572 & ~n35574 ;
  assign n35576 = \m5_data_i[24]_pad  & ~n1910 ;
  assign n35577 = n1941 & n35576 ;
  assign n35578 = \m2_data_i[24]_pad  & ~n1925 ;
  assign n35579 = n1931 & n35578 ;
  assign n35580 = ~n35577 & ~n35579 ;
  assign n35581 = n35575 & n35580 ;
  assign n35582 = \m4_data_i[24]_pad  & n1925 ;
  assign n35583 = n1918 & n35582 ;
  assign n35584 = \m3_data_i[24]_pad  & n1910 ;
  assign n35585 = n1938 & n35584 ;
  assign n35586 = ~n35583 & ~n35585 ;
  assign n35587 = \m1_data_i[24]_pad  & n1910 ;
  assign n35588 = n1941 & n35587 ;
  assign n35589 = \m0_data_i[24]_pad  & n1925 ;
  assign n35590 = n1931 & n35589 ;
  assign n35591 = ~n35588 & ~n35590 ;
  assign n35592 = n35586 & n35591 ;
  assign n35593 = n35581 & n35592 ;
  assign n35594 = \m7_data_i[25]_pad  & ~n1910 ;
  assign n35595 = n1938 & n35594 ;
  assign n35596 = \m6_data_i[25]_pad  & ~n1925 ;
  assign n35597 = n1918 & n35596 ;
  assign n35598 = ~n35595 & ~n35597 ;
  assign n35599 = \m5_data_i[25]_pad  & ~n1910 ;
  assign n35600 = n1941 & n35599 ;
  assign n35601 = \m2_data_i[25]_pad  & ~n1925 ;
  assign n35602 = n1931 & n35601 ;
  assign n35603 = ~n35600 & ~n35602 ;
  assign n35604 = n35598 & n35603 ;
  assign n35605 = \m4_data_i[25]_pad  & n1925 ;
  assign n35606 = n1918 & n35605 ;
  assign n35607 = \m3_data_i[25]_pad  & n1910 ;
  assign n35608 = n1938 & n35607 ;
  assign n35609 = ~n35606 & ~n35608 ;
  assign n35610 = \m1_data_i[25]_pad  & n1910 ;
  assign n35611 = n1941 & n35610 ;
  assign n35612 = \m0_data_i[25]_pad  & n1925 ;
  assign n35613 = n1931 & n35612 ;
  assign n35614 = ~n35611 & ~n35613 ;
  assign n35615 = n35609 & n35614 ;
  assign n35616 = n35604 & n35615 ;
  assign n35617 = \m7_data_i[26]_pad  & ~n1910 ;
  assign n35618 = n1938 & n35617 ;
  assign n35619 = \m6_data_i[26]_pad  & ~n1925 ;
  assign n35620 = n1918 & n35619 ;
  assign n35621 = ~n35618 & ~n35620 ;
  assign n35622 = \m5_data_i[26]_pad  & ~n1910 ;
  assign n35623 = n1941 & n35622 ;
  assign n35624 = \m2_data_i[26]_pad  & ~n1925 ;
  assign n35625 = n1931 & n35624 ;
  assign n35626 = ~n35623 & ~n35625 ;
  assign n35627 = n35621 & n35626 ;
  assign n35628 = \m4_data_i[26]_pad  & n1925 ;
  assign n35629 = n1918 & n35628 ;
  assign n35630 = \m3_data_i[26]_pad  & n1910 ;
  assign n35631 = n1938 & n35630 ;
  assign n35632 = ~n35629 & ~n35631 ;
  assign n35633 = \m1_data_i[26]_pad  & n1910 ;
  assign n35634 = n1941 & n35633 ;
  assign n35635 = \m0_data_i[26]_pad  & n1925 ;
  assign n35636 = n1931 & n35635 ;
  assign n35637 = ~n35634 & ~n35636 ;
  assign n35638 = n35632 & n35637 ;
  assign n35639 = n35627 & n35638 ;
  assign n35640 = \m7_data_i[27]_pad  & ~n1910 ;
  assign n35641 = n1938 & n35640 ;
  assign n35642 = \m6_data_i[27]_pad  & ~n1925 ;
  assign n35643 = n1918 & n35642 ;
  assign n35644 = ~n35641 & ~n35643 ;
  assign n35645 = \m5_data_i[27]_pad  & ~n1910 ;
  assign n35646 = n1941 & n35645 ;
  assign n35647 = \m2_data_i[27]_pad  & ~n1925 ;
  assign n35648 = n1931 & n35647 ;
  assign n35649 = ~n35646 & ~n35648 ;
  assign n35650 = n35644 & n35649 ;
  assign n35651 = \m4_data_i[27]_pad  & n1925 ;
  assign n35652 = n1918 & n35651 ;
  assign n35653 = \m3_data_i[27]_pad  & n1910 ;
  assign n35654 = n1938 & n35653 ;
  assign n35655 = ~n35652 & ~n35654 ;
  assign n35656 = \m1_data_i[27]_pad  & n1910 ;
  assign n35657 = n1941 & n35656 ;
  assign n35658 = \m0_data_i[27]_pad  & n1925 ;
  assign n35659 = n1931 & n35658 ;
  assign n35660 = ~n35657 & ~n35659 ;
  assign n35661 = n35655 & n35660 ;
  assign n35662 = n35650 & n35661 ;
  assign n35663 = \m7_data_i[28]_pad  & ~n1910 ;
  assign n35664 = n1938 & n35663 ;
  assign n35665 = \m6_data_i[28]_pad  & ~n1925 ;
  assign n35666 = n1918 & n35665 ;
  assign n35667 = ~n35664 & ~n35666 ;
  assign n35668 = \m5_data_i[28]_pad  & ~n1910 ;
  assign n35669 = n1941 & n35668 ;
  assign n35670 = \m2_data_i[28]_pad  & ~n1925 ;
  assign n35671 = n1931 & n35670 ;
  assign n35672 = ~n35669 & ~n35671 ;
  assign n35673 = n35667 & n35672 ;
  assign n35674 = \m4_data_i[28]_pad  & n1925 ;
  assign n35675 = n1918 & n35674 ;
  assign n35676 = \m3_data_i[28]_pad  & n1910 ;
  assign n35677 = n1938 & n35676 ;
  assign n35678 = ~n35675 & ~n35677 ;
  assign n35679 = \m1_data_i[28]_pad  & n1910 ;
  assign n35680 = n1941 & n35679 ;
  assign n35681 = \m0_data_i[28]_pad  & n1925 ;
  assign n35682 = n1931 & n35681 ;
  assign n35683 = ~n35680 & ~n35682 ;
  assign n35684 = n35678 & n35683 ;
  assign n35685 = n35673 & n35684 ;
  assign n35686 = \m5_data_i[29]_pad  & ~n1910 ;
  assign n35687 = n1941 & n35686 ;
  assign n35688 = \m4_data_i[29]_pad  & n1925 ;
  assign n35689 = n1918 & n35688 ;
  assign n35690 = ~n35687 & ~n35689 ;
  assign n35691 = \m3_data_i[29]_pad  & n1910 ;
  assign n35692 = n1938 & n35691 ;
  assign n35693 = \m0_data_i[29]_pad  & n1925 ;
  assign n35694 = n1931 & n35693 ;
  assign n35695 = ~n35692 & ~n35694 ;
  assign n35696 = n35690 & n35695 ;
  assign n35697 = \m2_data_i[29]_pad  & ~n1925 ;
  assign n35698 = n1931 & n35697 ;
  assign n35699 = \m1_data_i[29]_pad  & n1910 ;
  assign n35700 = n1941 & n35699 ;
  assign n35701 = ~n35698 & ~n35700 ;
  assign n35702 = \m7_data_i[29]_pad  & ~n1910 ;
  assign n35703 = n1938 & n35702 ;
  assign n35704 = \m6_data_i[29]_pad  & ~n1925 ;
  assign n35705 = n1918 & n35704 ;
  assign n35706 = ~n35703 & ~n35705 ;
  assign n35707 = n35701 & n35706 ;
  assign n35708 = n35696 & n35707 ;
  assign n35709 = \m3_data_i[30]_pad  & n1910 ;
  assign n35710 = n1938 & n35709 ;
  assign n35711 = \m2_data_i[30]_pad  & ~n1925 ;
  assign n35712 = n1931 & n35711 ;
  assign n35713 = ~n35710 & ~n35712 ;
  assign n35714 = \m5_data_i[30]_pad  & ~n1910 ;
  assign n35715 = n1941 & n35714 ;
  assign n35716 = \m6_data_i[30]_pad  & ~n1925 ;
  assign n35717 = n1918 & n35716 ;
  assign n35718 = ~n35715 & ~n35717 ;
  assign n35719 = n35713 & n35718 ;
  assign n35720 = \m4_data_i[30]_pad  & n1925 ;
  assign n35721 = n1918 & n35720 ;
  assign n35722 = \m7_data_i[30]_pad  & ~n1910 ;
  assign n35723 = n1938 & n35722 ;
  assign n35724 = ~n35721 & ~n35723 ;
  assign n35725 = \m1_data_i[30]_pad  & n1910 ;
  assign n35726 = n1941 & n35725 ;
  assign n35727 = \m0_data_i[30]_pad  & n1925 ;
  assign n35728 = n1931 & n35727 ;
  assign n35729 = ~n35726 & ~n35728 ;
  assign n35730 = n35724 & n35729 ;
  assign n35731 = n35719 & n35730 ;
  assign n35732 = \m7_data_i[31]_pad  & ~n1910 ;
  assign n35733 = n1938 & n35732 ;
  assign n35734 = \m6_data_i[31]_pad  & ~n1925 ;
  assign n35735 = n1918 & n35734 ;
  assign n35736 = ~n35733 & ~n35735 ;
  assign n35737 = \m5_data_i[31]_pad  & ~n1910 ;
  assign n35738 = n1941 & n35737 ;
  assign n35739 = \m2_data_i[31]_pad  & ~n1925 ;
  assign n35740 = n1931 & n35739 ;
  assign n35741 = ~n35738 & ~n35740 ;
  assign n35742 = n35736 & n35741 ;
  assign n35743 = \m4_data_i[31]_pad  & n1925 ;
  assign n35744 = n1918 & n35743 ;
  assign n35745 = \m3_data_i[31]_pad  & n1910 ;
  assign n35746 = n1938 & n35745 ;
  assign n35747 = ~n35744 & ~n35746 ;
  assign n35748 = \m1_data_i[31]_pad  & n1910 ;
  assign n35749 = n1941 & n35748 ;
  assign n35750 = \m0_data_i[31]_pad  & n1925 ;
  assign n35751 = n1931 & n35750 ;
  assign n35752 = ~n35749 & ~n35751 ;
  assign n35753 = n35747 & n35752 ;
  assign n35754 = n35742 & n35753 ;
  assign n35755 = \m7_sel_i[0]_pad  & ~n1910 ;
  assign n35756 = n1938 & n35755 ;
  assign n35757 = \m6_sel_i[0]_pad  & ~n1925 ;
  assign n35758 = n1918 & n35757 ;
  assign n35759 = ~n35756 & ~n35758 ;
  assign n35760 = \m5_sel_i[0]_pad  & ~n1910 ;
  assign n35761 = n1941 & n35760 ;
  assign n35762 = \m2_sel_i[0]_pad  & ~n1925 ;
  assign n35763 = n1931 & n35762 ;
  assign n35764 = ~n35761 & ~n35763 ;
  assign n35765 = n35759 & n35764 ;
  assign n35766 = \m4_sel_i[0]_pad  & n1925 ;
  assign n35767 = n1918 & n35766 ;
  assign n35768 = \m3_sel_i[0]_pad  & n1910 ;
  assign n35769 = n1938 & n35768 ;
  assign n35770 = ~n35767 & ~n35769 ;
  assign n35771 = \m1_sel_i[0]_pad  & n1910 ;
  assign n35772 = n1941 & n35771 ;
  assign n35773 = \m0_sel_i[0]_pad  & n1925 ;
  assign n35774 = n1931 & n35773 ;
  assign n35775 = ~n35772 & ~n35774 ;
  assign n35776 = n35770 & n35775 ;
  assign n35777 = n35765 & n35776 ;
  assign n35778 = \m7_sel_i[1]_pad  & ~n1910 ;
  assign n35779 = n1938 & n35778 ;
  assign n35780 = \m6_sel_i[1]_pad  & ~n1925 ;
  assign n35781 = n1918 & n35780 ;
  assign n35782 = ~n35779 & ~n35781 ;
  assign n35783 = \m5_sel_i[1]_pad  & ~n1910 ;
  assign n35784 = n1941 & n35783 ;
  assign n35785 = \m2_sel_i[1]_pad  & ~n1925 ;
  assign n35786 = n1931 & n35785 ;
  assign n35787 = ~n35784 & ~n35786 ;
  assign n35788 = n35782 & n35787 ;
  assign n35789 = \m4_sel_i[1]_pad  & n1925 ;
  assign n35790 = n1918 & n35789 ;
  assign n35791 = \m3_sel_i[1]_pad  & n1910 ;
  assign n35792 = n1938 & n35791 ;
  assign n35793 = ~n35790 & ~n35792 ;
  assign n35794 = \m1_sel_i[1]_pad  & n1910 ;
  assign n35795 = n1941 & n35794 ;
  assign n35796 = \m0_sel_i[1]_pad  & n1925 ;
  assign n35797 = n1931 & n35796 ;
  assign n35798 = ~n35795 & ~n35797 ;
  assign n35799 = n35793 & n35798 ;
  assign n35800 = n35788 & n35799 ;
  assign n35801 = \m7_sel_i[2]_pad  & ~n1910 ;
  assign n35802 = n1938 & n35801 ;
  assign n35803 = \m6_sel_i[2]_pad  & ~n1925 ;
  assign n35804 = n1918 & n35803 ;
  assign n35805 = ~n35802 & ~n35804 ;
  assign n35806 = \m5_sel_i[2]_pad  & ~n1910 ;
  assign n35807 = n1941 & n35806 ;
  assign n35808 = \m2_sel_i[2]_pad  & ~n1925 ;
  assign n35809 = n1931 & n35808 ;
  assign n35810 = ~n35807 & ~n35809 ;
  assign n35811 = n35805 & n35810 ;
  assign n35812 = \m4_sel_i[2]_pad  & n1925 ;
  assign n35813 = n1918 & n35812 ;
  assign n35814 = \m3_sel_i[2]_pad  & n1910 ;
  assign n35815 = n1938 & n35814 ;
  assign n35816 = ~n35813 & ~n35815 ;
  assign n35817 = \m1_sel_i[2]_pad  & n1910 ;
  assign n35818 = n1941 & n35817 ;
  assign n35819 = \m0_sel_i[2]_pad  & n1925 ;
  assign n35820 = n1931 & n35819 ;
  assign n35821 = ~n35818 & ~n35820 ;
  assign n35822 = n35816 & n35821 ;
  assign n35823 = n35811 & n35822 ;
  assign n35824 = \m3_sel_i[3]_pad  & n1910 ;
  assign n35825 = n1938 & n35824 ;
  assign n35826 = \m2_sel_i[3]_pad  & ~n1925 ;
  assign n35827 = n1931 & n35826 ;
  assign n35828 = ~n35825 & ~n35827 ;
  assign n35829 = \m5_sel_i[3]_pad  & ~n1910 ;
  assign n35830 = n1941 & n35829 ;
  assign n35831 = \m0_sel_i[3]_pad  & n1925 ;
  assign n35832 = n1931 & n35831 ;
  assign n35833 = ~n35830 & ~n35832 ;
  assign n35834 = n35828 & n35833 ;
  assign n35835 = \m4_sel_i[3]_pad  & n1925 ;
  assign n35836 = n1918 & n35835 ;
  assign n35837 = \m1_sel_i[3]_pad  & n1910 ;
  assign n35838 = n1941 & n35837 ;
  assign n35839 = ~n35836 & ~n35838 ;
  assign n35840 = \m7_sel_i[3]_pad  & ~n1910 ;
  assign n35841 = n1938 & n35840 ;
  assign n35842 = \m6_sel_i[3]_pad  & ~n1925 ;
  assign n35843 = n1918 & n35842 ;
  assign n35844 = ~n35841 & ~n35843 ;
  assign n35845 = n35839 & n35844 ;
  assign n35846 = n35834 & n35845 ;
  assign n35847 = \m3_addr_i[0]_pad  & ~n14271 ;
  assign n35848 = n14279 & n35847 ;
  assign n35849 = \m4_addr_i[0]_pad  & n14271 ;
  assign n35850 = n14288 & n35849 ;
  assign n35851 = ~n35848 & ~n35850 ;
  assign n35852 = \m6_addr_i[0]_pad  & n14271 ;
  assign n35853 = n14264 & n35852 ;
  assign n35854 = \m2_addr_i[0]_pad  & n14271 ;
  assign n35855 = n14279 & n35854 ;
  assign n35856 = ~n35853 & ~n35855 ;
  assign n35857 = n35851 & n35856 ;
  assign n35858 = \m5_addr_i[0]_pad  & ~n14271 ;
  assign n35859 = n14288 & n35858 ;
  assign n35860 = \m1_addr_i[0]_pad  & ~n14271 ;
  assign n35861 = n14296 & n35860 ;
  assign n35862 = ~n35859 & ~n35861 ;
  assign n35863 = \m0_addr_i[0]_pad  & n14271 ;
  assign n35864 = n14296 & n35863 ;
  assign n35865 = \m7_addr_i[0]_pad  & ~n14271 ;
  assign n35866 = n14264 & n35865 ;
  assign n35867 = ~n35864 & ~n35866 ;
  assign n35868 = n35862 & n35867 ;
  assign n35869 = n35857 & n35868 ;
  assign n35870 = \m3_addr_i[10]_pad  & ~n14271 ;
  assign n35871 = n14279 & n35870 ;
  assign n35872 = \m4_addr_i[10]_pad  & n14271 ;
  assign n35873 = n14288 & n35872 ;
  assign n35874 = ~n35871 & ~n35873 ;
  assign n35875 = \m6_addr_i[10]_pad  & n14271 ;
  assign n35876 = n14264 & n35875 ;
  assign n35877 = \m2_addr_i[10]_pad  & n14271 ;
  assign n35878 = n14279 & n35877 ;
  assign n35879 = ~n35876 & ~n35878 ;
  assign n35880 = n35874 & n35879 ;
  assign n35881 = \m5_addr_i[10]_pad  & ~n14271 ;
  assign n35882 = n14288 & n35881 ;
  assign n35883 = \m1_addr_i[10]_pad  & ~n14271 ;
  assign n35884 = n14296 & n35883 ;
  assign n35885 = ~n35882 & ~n35884 ;
  assign n35886 = \m0_addr_i[10]_pad  & n14271 ;
  assign n35887 = n14296 & n35886 ;
  assign n35888 = \m7_addr_i[10]_pad  & ~n14271 ;
  assign n35889 = n14264 & n35888 ;
  assign n35890 = ~n35887 & ~n35889 ;
  assign n35891 = n35885 & n35890 ;
  assign n35892 = n35880 & n35891 ;
  assign n35893 = \m0_addr_i[11]_pad  & n14271 ;
  assign n35894 = n14296 & n35893 ;
  assign n35895 = \m7_addr_i[11]_pad  & ~n14271 ;
  assign n35896 = n14264 & n35895 ;
  assign n35897 = ~n35894 & ~n35896 ;
  assign n35898 = \m6_addr_i[11]_pad  & n14271 ;
  assign n35899 = n14264 & n35898 ;
  assign n35900 = \m2_addr_i[11]_pad  & n14271 ;
  assign n35901 = n14279 & n35900 ;
  assign n35902 = ~n35899 & ~n35901 ;
  assign n35903 = n35897 & n35902 ;
  assign n35904 = \m5_addr_i[11]_pad  & ~n14271 ;
  assign n35905 = n14288 & n35904 ;
  assign n35906 = \m1_addr_i[11]_pad  & ~n14271 ;
  assign n35907 = n14296 & n35906 ;
  assign n35908 = ~n35905 & ~n35907 ;
  assign n35909 = \m3_addr_i[11]_pad  & ~n14271 ;
  assign n35910 = n14279 & n35909 ;
  assign n35911 = \m4_addr_i[11]_pad  & n14271 ;
  assign n35912 = n14288 & n35911 ;
  assign n35913 = ~n35910 & ~n35912 ;
  assign n35914 = n35908 & n35913 ;
  assign n35915 = n35903 & n35914 ;
  assign n35916 = \m1_addr_i[12]_pad  & ~n14271 ;
  assign n35917 = n14296 & n35916 ;
  assign n35918 = \m2_addr_i[12]_pad  & n14271 ;
  assign n35919 = n14279 & n35918 ;
  assign n35920 = ~n35917 & ~n35919 ;
  assign n35921 = \m0_addr_i[12]_pad  & n14271 ;
  assign n35922 = n14296 & n35921 ;
  assign n35923 = \m4_addr_i[12]_pad  & n14271 ;
  assign n35924 = n14288 & n35923 ;
  assign n35925 = ~n35922 & ~n35924 ;
  assign n35926 = n35920 & n35925 ;
  assign n35927 = \m7_addr_i[12]_pad  & ~n14271 ;
  assign n35928 = n14264 & n35927 ;
  assign n35929 = \m3_addr_i[12]_pad  & ~n14271 ;
  assign n35930 = n14279 & n35929 ;
  assign n35931 = ~n35928 & ~n35930 ;
  assign n35932 = \m6_addr_i[12]_pad  & n14271 ;
  assign n35933 = n14264 & n35932 ;
  assign n35934 = \m5_addr_i[12]_pad  & ~n14271 ;
  assign n35935 = n14288 & n35934 ;
  assign n35936 = ~n35933 & ~n35935 ;
  assign n35937 = n35931 & n35936 ;
  assign n35938 = n35926 & n35937 ;
  assign n35939 = \m3_addr_i[13]_pad  & ~n14271 ;
  assign n35940 = n14279 & n35939 ;
  assign n35941 = \m4_addr_i[13]_pad  & n14271 ;
  assign n35942 = n14288 & n35941 ;
  assign n35943 = ~n35940 & ~n35942 ;
  assign n35944 = \m6_addr_i[13]_pad  & n14271 ;
  assign n35945 = n14264 & n35944 ;
  assign n35946 = \m7_addr_i[13]_pad  & ~n14271 ;
  assign n35947 = n14264 & n35946 ;
  assign n35948 = ~n35945 & ~n35947 ;
  assign n35949 = n35943 & n35948 ;
  assign n35950 = \m5_addr_i[13]_pad  & ~n14271 ;
  assign n35951 = n14288 & n35950 ;
  assign n35952 = \m0_addr_i[13]_pad  & n14271 ;
  assign n35953 = n14296 & n35952 ;
  assign n35954 = ~n35951 & ~n35953 ;
  assign n35955 = \m1_addr_i[13]_pad  & ~n14271 ;
  assign n35956 = n14296 & n35955 ;
  assign n35957 = \m2_addr_i[13]_pad  & n14271 ;
  assign n35958 = n14279 & n35957 ;
  assign n35959 = ~n35956 & ~n35958 ;
  assign n35960 = n35954 & n35959 ;
  assign n35961 = n35949 & n35960 ;
  assign n35962 = \m3_addr_i[14]_pad  & ~n14271 ;
  assign n35963 = n14279 & n35962 ;
  assign n35964 = \m4_addr_i[14]_pad  & n14271 ;
  assign n35965 = n14288 & n35964 ;
  assign n35966 = ~n35963 & ~n35965 ;
  assign n35967 = \m6_addr_i[14]_pad  & n14271 ;
  assign n35968 = n14264 & n35967 ;
  assign n35969 = \m2_addr_i[14]_pad  & n14271 ;
  assign n35970 = n14279 & n35969 ;
  assign n35971 = ~n35968 & ~n35970 ;
  assign n35972 = n35966 & n35971 ;
  assign n35973 = \m5_addr_i[14]_pad  & ~n14271 ;
  assign n35974 = n14288 & n35973 ;
  assign n35975 = \m1_addr_i[14]_pad  & ~n14271 ;
  assign n35976 = n14296 & n35975 ;
  assign n35977 = ~n35974 & ~n35976 ;
  assign n35978 = \m0_addr_i[14]_pad  & n14271 ;
  assign n35979 = n14296 & n35978 ;
  assign n35980 = \m7_addr_i[14]_pad  & ~n14271 ;
  assign n35981 = n14264 & n35980 ;
  assign n35982 = ~n35979 & ~n35981 ;
  assign n35983 = n35977 & n35982 ;
  assign n35984 = n35972 & n35983 ;
  assign n35985 = \m3_addr_i[15]_pad  & ~n14271 ;
  assign n35986 = n14279 & n35985 ;
  assign n35987 = \m4_addr_i[15]_pad  & n14271 ;
  assign n35988 = n14288 & n35987 ;
  assign n35989 = ~n35986 & ~n35988 ;
  assign n35990 = \m6_addr_i[15]_pad  & n14271 ;
  assign n35991 = n14264 & n35990 ;
  assign n35992 = \m2_addr_i[15]_pad  & n14271 ;
  assign n35993 = n14279 & n35992 ;
  assign n35994 = ~n35991 & ~n35993 ;
  assign n35995 = n35989 & n35994 ;
  assign n35996 = \m5_addr_i[15]_pad  & ~n14271 ;
  assign n35997 = n14288 & n35996 ;
  assign n35998 = \m1_addr_i[15]_pad  & ~n14271 ;
  assign n35999 = n14296 & n35998 ;
  assign n36000 = ~n35997 & ~n35999 ;
  assign n36001 = \m0_addr_i[15]_pad  & n14271 ;
  assign n36002 = n14296 & n36001 ;
  assign n36003 = \m7_addr_i[15]_pad  & ~n14271 ;
  assign n36004 = n14264 & n36003 ;
  assign n36005 = ~n36002 & ~n36004 ;
  assign n36006 = n36000 & n36005 ;
  assign n36007 = n35995 & n36006 ;
  assign n36008 = \m1_addr_i[16]_pad  & ~n14271 ;
  assign n36009 = n14296 & n36008 ;
  assign n36010 = \m2_addr_i[16]_pad  & n14271 ;
  assign n36011 = n14279 & n36010 ;
  assign n36012 = ~n36009 & ~n36011 ;
  assign n36013 = \m6_addr_i[16]_pad  & n14271 ;
  assign n36014 = n14264 & n36013 ;
  assign n36015 = \m7_addr_i[16]_pad  & ~n14271 ;
  assign n36016 = n14264 & n36015 ;
  assign n36017 = ~n36014 & ~n36016 ;
  assign n36018 = n36012 & n36017 ;
  assign n36019 = \m5_addr_i[16]_pad  & ~n14271 ;
  assign n36020 = n14288 & n36019 ;
  assign n36021 = \m0_addr_i[16]_pad  & n14271 ;
  assign n36022 = n14296 & n36021 ;
  assign n36023 = ~n36020 & ~n36022 ;
  assign n36024 = \m3_addr_i[16]_pad  & ~n14271 ;
  assign n36025 = n14279 & n36024 ;
  assign n36026 = \m4_addr_i[16]_pad  & n14271 ;
  assign n36027 = n14288 & n36026 ;
  assign n36028 = ~n36025 & ~n36027 ;
  assign n36029 = n36023 & n36028 ;
  assign n36030 = n36018 & n36029 ;
  assign n36031 = \m6_addr_i[17]_pad  & n14271 ;
  assign n36032 = n14264 & n36031 ;
  assign n36033 = \m5_addr_i[17]_pad  & ~n14271 ;
  assign n36034 = n14288 & n36033 ;
  assign n36035 = ~n36032 & ~n36034 ;
  assign n36036 = \m0_addr_i[17]_pad  & n14271 ;
  assign n36037 = n14296 & n36036 ;
  assign n36038 = \m4_addr_i[17]_pad  & n14271 ;
  assign n36039 = n14288 & n36038 ;
  assign n36040 = ~n36037 & ~n36039 ;
  assign n36041 = n36035 & n36040 ;
  assign n36042 = \m7_addr_i[17]_pad  & ~n14271 ;
  assign n36043 = n14264 & n36042 ;
  assign n36044 = \m3_addr_i[17]_pad  & ~n14271 ;
  assign n36045 = n14279 & n36044 ;
  assign n36046 = ~n36043 & ~n36045 ;
  assign n36047 = \m1_addr_i[17]_pad  & ~n14271 ;
  assign n36048 = n14296 & n36047 ;
  assign n36049 = \m2_addr_i[17]_pad  & n14271 ;
  assign n36050 = n14279 & n36049 ;
  assign n36051 = ~n36048 & ~n36050 ;
  assign n36052 = n36046 & n36051 ;
  assign n36053 = n36041 & n36052 ;
  assign n36054 = \m3_addr_i[18]_pad  & ~n14271 ;
  assign n36055 = n14279 & n36054 ;
  assign n36056 = \m4_addr_i[18]_pad  & n14271 ;
  assign n36057 = n14288 & n36056 ;
  assign n36058 = ~n36055 & ~n36057 ;
  assign n36059 = \m6_addr_i[18]_pad  & n14271 ;
  assign n36060 = n14264 & n36059 ;
  assign n36061 = \m2_addr_i[18]_pad  & n14271 ;
  assign n36062 = n14279 & n36061 ;
  assign n36063 = ~n36060 & ~n36062 ;
  assign n36064 = n36058 & n36063 ;
  assign n36065 = \m5_addr_i[18]_pad  & ~n14271 ;
  assign n36066 = n14288 & n36065 ;
  assign n36067 = \m1_addr_i[18]_pad  & ~n14271 ;
  assign n36068 = n14296 & n36067 ;
  assign n36069 = ~n36066 & ~n36068 ;
  assign n36070 = \m0_addr_i[18]_pad  & n14271 ;
  assign n36071 = n14296 & n36070 ;
  assign n36072 = \m7_addr_i[18]_pad  & ~n14271 ;
  assign n36073 = n14264 & n36072 ;
  assign n36074 = ~n36071 & ~n36073 ;
  assign n36075 = n36069 & n36074 ;
  assign n36076 = n36064 & n36075 ;
  assign n36077 = \m3_addr_i[19]_pad  & ~n14271 ;
  assign n36078 = n14279 & n36077 ;
  assign n36079 = \m4_addr_i[19]_pad  & n14271 ;
  assign n36080 = n14288 & n36079 ;
  assign n36081 = ~n36078 & ~n36080 ;
  assign n36082 = \m6_addr_i[19]_pad  & n14271 ;
  assign n36083 = n14264 & n36082 ;
  assign n36084 = \m2_addr_i[19]_pad  & n14271 ;
  assign n36085 = n14279 & n36084 ;
  assign n36086 = ~n36083 & ~n36085 ;
  assign n36087 = n36081 & n36086 ;
  assign n36088 = \m5_addr_i[19]_pad  & ~n14271 ;
  assign n36089 = n14288 & n36088 ;
  assign n36090 = \m1_addr_i[19]_pad  & ~n14271 ;
  assign n36091 = n14296 & n36090 ;
  assign n36092 = ~n36089 & ~n36091 ;
  assign n36093 = \m0_addr_i[19]_pad  & n14271 ;
  assign n36094 = n14296 & n36093 ;
  assign n36095 = \m7_addr_i[19]_pad  & ~n14271 ;
  assign n36096 = n14264 & n36095 ;
  assign n36097 = ~n36094 & ~n36096 ;
  assign n36098 = n36092 & n36097 ;
  assign n36099 = n36087 & n36098 ;
  assign n36100 = \m3_addr_i[1]_pad  & ~n14271 ;
  assign n36101 = n14279 & n36100 ;
  assign n36102 = \m4_addr_i[1]_pad  & n14271 ;
  assign n36103 = n14288 & n36102 ;
  assign n36104 = ~n36101 & ~n36103 ;
  assign n36105 = \m6_addr_i[1]_pad  & n14271 ;
  assign n36106 = n14264 & n36105 ;
  assign n36107 = \m2_addr_i[1]_pad  & n14271 ;
  assign n36108 = n14279 & n36107 ;
  assign n36109 = ~n36106 & ~n36108 ;
  assign n36110 = n36104 & n36109 ;
  assign n36111 = \m5_addr_i[1]_pad  & ~n14271 ;
  assign n36112 = n14288 & n36111 ;
  assign n36113 = \m1_addr_i[1]_pad  & ~n14271 ;
  assign n36114 = n14296 & n36113 ;
  assign n36115 = ~n36112 & ~n36114 ;
  assign n36116 = \m0_addr_i[1]_pad  & n14271 ;
  assign n36117 = n14296 & n36116 ;
  assign n36118 = \m7_addr_i[1]_pad  & ~n14271 ;
  assign n36119 = n14264 & n36118 ;
  assign n36120 = ~n36117 & ~n36119 ;
  assign n36121 = n36115 & n36120 ;
  assign n36122 = n36110 & n36121 ;
  assign n36123 = \m1_addr_i[20]_pad  & ~n14271 ;
  assign n36124 = n14296 & n36123 ;
  assign n36125 = \m2_addr_i[20]_pad  & n14271 ;
  assign n36126 = n14279 & n36125 ;
  assign n36127 = ~n36124 & ~n36126 ;
  assign n36128 = \m3_addr_i[20]_pad  & ~n14271 ;
  assign n36129 = n14279 & n36128 ;
  assign n36130 = \m7_addr_i[20]_pad  & ~n14271 ;
  assign n36131 = n14264 & n36130 ;
  assign n36132 = ~n36129 & ~n36131 ;
  assign n36133 = n36127 & n36132 ;
  assign n36134 = \m4_addr_i[20]_pad  & n14271 ;
  assign n36135 = n14288 & n36134 ;
  assign n36136 = \m0_addr_i[20]_pad  & n14271 ;
  assign n36137 = n14296 & n36136 ;
  assign n36138 = ~n36135 & ~n36137 ;
  assign n36139 = \m6_addr_i[20]_pad  & n14271 ;
  assign n36140 = n14264 & n36139 ;
  assign n36141 = \m5_addr_i[20]_pad  & ~n14271 ;
  assign n36142 = n14288 & n36141 ;
  assign n36143 = ~n36140 & ~n36142 ;
  assign n36144 = n36138 & n36143 ;
  assign n36145 = n36133 & n36144 ;
  assign n36146 = \m0_addr_i[21]_pad  & n14271 ;
  assign n36147 = n14296 & n36146 ;
  assign n36148 = \m7_addr_i[21]_pad  & ~n14271 ;
  assign n36149 = n14264 & n36148 ;
  assign n36150 = ~n36147 & ~n36149 ;
  assign n36151 = \m1_addr_i[21]_pad  & ~n14271 ;
  assign n36152 = n14296 & n36151 ;
  assign n36153 = \m5_addr_i[21]_pad  & ~n14271 ;
  assign n36154 = n14288 & n36153 ;
  assign n36155 = ~n36152 & ~n36154 ;
  assign n36156 = n36150 & n36155 ;
  assign n36157 = \m2_addr_i[21]_pad  & n14271 ;
  assign n36158 = n14279 & n36157 ;
  assign n36159 = \m6_addr_i[21]_pad  & n14271 ;
  assign n36160 = n14264 & n36159 ;
  assign n36161 = ~n36158 & ~n36160 ;
  assign n36162 = \m3_addr_i[21]_pad  & ~n14271 ;
  assign n36163 = n14279 & n36162 ;
  assign n36164 = \m4_addr_i[21]_pad  & n14271 ;
  assign n36165 = n14288 & n36164 ;
  assign n36166 = ~n36163 & ~n36165 ;
  assign n36167 = n36161 & n36166 ;
  assign n36168 = n36156 & n36167 ;
  assign n36169 = \m1_addr_i[22]_pad  & ~n14271 ;
  assign n36170 = n14296 & n36169 ;
  assign n36171 = \m2_addr_i[22]_pad  & n14271 ;
  assign n36172 = n14279 & n36171 ;
  assign n36173 = ~n36170 & ~n36172 ;
  assign n36174 = \m3_addr_i[22]_pad  & ~n14271 ;
  assign n36175 = n14279 & n36174 ;
  assign n36176 = \m7_addr_i[22]_pad  & ~n14271 ;
  assign n36177 = n14264 & n36176 ;
  assign n36178 = ~n36175 & ~n36177 ;
  assign n36179 = n36173 & n36178 ;
  assign n36180 = \m4_addr_i[22]_pad  & n14271 ;
  assign n36181 = n14288 & n36180 ;
  assign n36182 = \m0_addr_i[22]_pad  & n14271 ;
  assign n36183 = n14296 & n36182 ;
  assign n36184 = ~n36181 & ~n36183 ;
  assign n36185 = \m6_addr_i[22]_pad  & n14271 ;
  assign n36186 = n14264 & n36185 ;
  assign n36187 = \m5_addr_i[22]_pad  & ~n14271 ;
  assign n36188 = n14288 & n36187 ;
  assign n36189 = ~n36186 & ~n36188 ;
  assign n36190 = n36184 & n36189 ;
  assign n36191 = n36179 & n36190 ;
  assign n36192 = \m1_addr_i[23]_pad  & ~n14271 ;
  assign n36193 = n14296 & n36192 ;
  assign n36194 = \m2_addr_i[23]_pad  & n14271 ;
  assign n36195 = n14279 & n36194 ;
  assign n36196 = ~n36193 & ~n36195 ;
  assign n36197 = \m0_addr_i[23]_pad  & n14271 ;
  assign n36198 = n14296 & n36197 ;
  assign n36199 = \m5_addr_i[23]_pad  & ~n14271 ;
  assign n36200 = n14288 & n36199 ;
  assign n36201 = ~n36198 & ~n36200 ;
  assign n36202 = n36196 & n36201 ;
  assign n36203 = \m7_addr_i[23]_pad  & ~n14271 ;
  assign n36204 = n14264 & n36203 ;
  assign n36205 = \m6_addr_i[23]_pad  & n14271 ;
  assign n36206 = n14264 & n36205 ;
  assign n36207 = ~n36204 & ~n36206 ;
  assign n36208 = \m3_addr_i[23]_pad  & ~n14271 ;
  assign n36209 = n14279 & n36208 ;
  assign n36210 = \m4_addr_i[23]_pad  & n14271 ;
  assign n36211 = n14288 & n36210 ;
  assign n36212 = ~n36209 & ~n36211 ;
  assign n36213 = n36207 & n36212 ;
  assign n36214 = n36202 & n36213 ;
  assign n36215 = \m5_addr_i[24]_pad  & ~n14271 ;
  assign n36216 = n14288 & n36215 ;
  assign n36217 = \m6_addr_i[24]_pad  & n14271 ;
  assign n36218 = n14264 & n36217 ;
  assign n36219 = ~n36216 & ~n36218 ;
  assign n36220 = \m1_addr_i[24]_pad  & ~n14271 ;
  assign n36221 = n14296 & n36220 ;
  assign n36222 = \m7_addr_i[24]_pad  & ~n14271 ;
  assign n36223 = n14264 & n36222 ;
  assign n36224 = ~n36221 & ~n36223 ;
  assign n36225 = n36219 & n36224 ;
  assign n36226 = \m2_addr_i[24]_pad  & n14271 ;
  assign n36227 = n14279 & n36226 ;
  assign n36228 = \m0_addr_i[24]_pad  & n14271 ;
  assign n36229 = n14296 & n36228 ;
  assign n36230 = ~n36227 & ~n36229 ;
  assign n36231 = \m3_addr_i[24]_pad  & ~n14271 ;
  assign n36232 = n14279 & n36231 ;
  assign n36233 = \m4_addr_i[24]_pad  & n14271 ;
  assign n36234 = n14288 & n36233 ;
  assign n36235 = ~n36232 & ~n36234 ;
  assign n36236 = n36230 & n36235 ;
  assign n36237 = n36225 & n36236 ;
  assign n36238 = \m1_addr_i[25]_pad  & ~n14271 ;
  assign n36239 = n14296 & n36238 ;
  assign n36240 = \m2_addr_i[25]_pad  & n14271 ;
  assign n36241 = n14279 & n36240 ;
  assign n36242 = ~n36239 & ~n36241 ;
  assign n36243 = \m0_addr_i[25]_pad  & n14271 ;
  assign n36244 = n14296 & n36243 ;
  assign n36245 = \m4_addr_i[25]_pad  & n14271 ;
  assign n36246 = n14288 & n36245 ;
  assign n36247 = ~n36244 & ~n36246 ;
  assign n36248 = n36242 & n36247 ;
  assign n36249 = \m7_addr_i[25]_pad  & ~n14271 ;
  assign n36250 = n14264 & n36249 ;
  assign n36251 = \m3_addr_i[25]_pad  & ~n14271 ;
  assign n36252 = n14279 & n36251 ;
  assign n36253 = ~n36250 & ~n36252 ;
  assign n36254 = \m5_addr_i[25]_pad  & ~n14271 ;
  assign n36255 = n14288 & n36254 ;
  assign n36256 = \m6_addr_i[25]_pad  & n14271 ;
  assign n36257 = n14264 & n36256 ;
  assign n36258 = ~n36255 & ~n36257 ;
  assign n36259 = n36253 & n36258 ;
  assign n36260 = n36248 & n36259 ;
  assign n36261 = \m3_addr_i[26]_pad  & ~n14271 ;
  assign n36262 = n14279 & n36261 ;
  assign n36263 = \m4_addr_i[26]_pad  & n14271 ;
  assign n36264 = n14288 & n36263 ;
  assign n36265 = ~n36262 & ~n36264 ;
  assign n36266 = \m1_addr_i[26]_pad  & ~n14271 ;
  assign n36267 = n14296 & n36266 ;
  assign n36268 = \m7_addr_i[26]_pad  & ~n14271 ;
  assign n36269 = n14264 & n36268 ;
  assign n36270 = ~n36267 & ~n36269 ;
  assign n36271 = n36265 & n36270 ;
  assign n36272 = \m2_addr_i[26]_pad  & n14271 ;
  assign n36273 = n14279 & n36272 ;
  assign n36274 = \m0_addr_i[26]_pad  & n14271 ;
  assign n36275 = n14296 & n36274 ;
  assign n36276 = ~n36273 & ~n36275 ;
  assign n36277 = \m5_addr_i[26]_pad  & ~n14271 ;
  assign n36278 = n14288 & n36277 ;
  assign n36279 = \m6_addr_i[26]_pad  & n14271 ;
  assign n36280 = n14264 & n36279 ;
  assign n36281 = ~n36278 & ~n36280 ;
  assign n36282 = n36276 & n36281 ;
  assign n36283 = n36271 & n36282 ;
  assign n36284 = \m1_addr_i[27]_pad  & ~n14271 ;
  assign n36285 = n14296 & n36284 ;
  assign n36286 = \m2_addr_i[27]_pad  & n14271 ;
  assign n36287 = n14279 & n36286 ;
  assign n36288 = ~n36285 & ~n36287 ;
  assign n36289 = \m0_addr_i[27]_pad  & n14271 ;
  assign n36290 = n14296 & n36289 ;
  assign n36291 = \m6_addr_i[27]_pad  & n14271 ;
  assign n36292 = n14264 & n36291 ;
  assign n36293 = ~n36290 & ~n36292 ;
  assign n36294 = n36288 & n36293 ;
  assign n36295 = \m7_addr_i[27]_pad  & ~n14271 ;
  assign n36296 = n14264 & n36295 ;
  assign n36297 = \m5_addr_i[27]_pad  & ~n14271 ;
  assign n36298 = n14288 & n36297 ;
  assign n36299 = ~n36296 & ~n36298 ;
  assign n36300 = \m3_addr_i[27]_pad  & ~n14271 ;
  assign n36301 = n14279 & n36300 ;
  assign n36302 = \m4_addr_i[27]_pad  & n14271 ;
  assign n36303 = n14288 & n36302 ;
  assign n36304 = ~n36301 & ~n36303 ;
  assign n36305 = n36299 & n36304 ;
  assign n36306 = n36294 & n36305 ;
  assign n36307 = \m1_addr_i[28]_pad  & ~n14271 ;
  assign n36308 = n14296 & n36307 ;
  assign n36309 = \m2_addr_i[28]_pad  & n14271 ;
  assign n36310 = n14279 & n36309 ;
  assign n36311 = ~n36308 & ~n36310 ;
  assign n36312 = \m0_addr_i[28]_pad  & n14271 ;
  assign n36313 = n14296 & n36312 ;
  assign n36314 = \m4_addr_i[28]_pad  & n14271 ;
  assign n36315 = n14288 & n36314 ;
  assign n36316 = ~n36313 & ~n36315 ;
  assign n36317 = n36311 & n36316 ;
  assign n36318 = \m7_addr_i[28]_pad  & ~n14271 ;
  assign n36319 = n14264 & n36318 ;
  assign n36320 = \m3_addr_i[28]_pad  & ~n14271 ;
  assign n36321 = n14279 & n36320 ;
  assign n36322 = ~n36319 & ~n36321 ;
  assign n36323 = \m5_addr_i[28]_pad  & ~n14271 ;
  assign n36324 = n14288 & n36323 ;
  assign n36325 = \m6_addr_i[28]_pad  & n14271 ;
  assign n36326 = n14264 & n36325 ;
  assign n36327 = ~n36324 & ~n36326 ;
  assign n36328 = n36322 & n36327 ;
  assign n36329 = n36317 & n36328 ;
  assign n36330 = \m0_addr_i[29]_pad  & n14271 ;
  assign n36331 = n14296 & n36330 ;
  assign n36332 = \m7_addr_i[29]_pad  & ~n14271 ;
  assign n36333 = n14264 & n36332 ;
  assign n36334 = ~n36331 & ~n36333 ;
  assign n36335 = \m5_addr_i[29]_pad  & ~n14271 ;
  assign n36336 = n14288 & n36335 ;
  assign n36337 = \m4_addr_i[29]_pad  & n14271 ;
  assign n36338 = n14288 & n36337 ;
  assign n36339 = ~n36336 & ~n36338 ;
  assign n36340 = n36334 & n36339 ;
  assign n36341 = \m6_addr_i[29]_pad  & n14271 ;
  assign n36342 = n14264 & n36341 ;
  assign n36343 = \m3_addr_i[29]_pad  & ~n14271 ;
  assign n36344 = n14279 & n36343 ;
  assign n36345 = ~n36342 & ~n36344 ;
  assign n36346 = \m1_addr_i[29]_pad  & ~n14271 ;
  assign n36347 = n14296 & n36346 ;
  assign n36348 = \m2_addr_i[29]_pad  & n14271 ;
  assign n36349 = n14279 & n36348 ;
  assign n36350 = ~n36347 & ~n36349 ;
  assign n36351 = n36345 & n36350 ;
  assign n36352 = n36340 & n36351 ;
  assign n36353 = \m3_addr_i[2]_pad  & ~n14271 ;
  assign n36354 = n14279 & n36353 ;
  assign n36355 = \m4_addr_i[2]_pad  & n14271 ;
  assign n36356 = n14288 & n36355 ;
  assign n36357 = ~n36354 & ~n36356 ;
  assign n36358 = \m6_addr_i[2]_pad  & n14271 ;
  assign n36359 = n14264 & n36358 ;
  assign n36360 = \m2_addr_i[2]_pad  & n14271 ;
  assign n36361 = n14279 & n36360 ;
  assign n36362 = ~n36359 & ~n36361 ;
  assign n36363 = n36357 & n36362 ;
  assign n36364 = \m5_addr_i[2]_pad  & ~n14271 ;
  assign n36365 = n14288 & n36364 ;
  assign n36366 = \m1_addr_i[2]_pad  & ~n14271 ;
  assign n36367 = n14296 & n36366 ;
  assign n36368 = ~n36365 & ~n36367 ;
  assign n36369 = \m0_addr_i[2]_pad  & n14271 ;
  assign n36370 = n14296 & n36369 ;
  assign n36371 = \m7_addr_i[2]_pad  & ~n14271 ;
  assign n36372 = n14264 & n36371 ;
  assign n36373 = ~n36370 & ~n36372 ;
  assign n36374 = n36368 & n36373 ;
  assign n36375 = n36363 & n36374 ;
  assign n36376 = \m3_addr_i[30]_pad  & ~n14271 ;
  assign n36377 = n14279 & n36376 ;
  assign n36378 = \m4_addr_i[30]_pad  & n14271 ;
  assign n36379 = n14288 & n36378 ;
  assign n36380 = ~n36377 & ~n36379 ;
  assign n36381 = \m0_addr_i[30]_pad  & n14271 ;
  assign n36382 = n14296 & n36381 ;
  assign n36383 = \m6_addr_i[30]_pad  & n14271 ;
  assign n36384 = n14264 & n36383 ;
  assign n36385 = ~n36382 & ~n36384 ;
  assign n36386 = n36380 & n36385 ;
  assign n36387 = \m7_addr_i[30]_pad  & ~n14271 ;
  assign n36388 = n14264 & n36387 ;
  assign n36389 = \m5_addr_i[30]_pad  & ~n14271 ;
  assign n36390 = n14288 & n36389 ;
  assign n36391 = ~n36388 & ~n36390 ;
  assign n36392 = \m1_addr_i[30]_pad  & ~n14271 ;
  assign n36393 = n14296 & n36392 ;
  assign n36394 = \m2_addr_i[30]_pad  & n14271 ;
  assign n36395 = n14279 & n36394 ;
  assign n36396 = ~n36393 & ~n36395 ;
  assign n36397 = n36391 & n36396 ;
  assign n36398 = n36386 & n36397 ;
  assign n36399 = \m5_addr_i[31]_pad  & ~n14271 ;
  assign n36400 = n14288 & n36399 ;
  assign n36401 = \m6_addr_i[31]_pad  & n14271 ;
  assign n36402 = n14264 & n36401 ;
  assign n36403 = ~n36400 & ~n36402 ;
  assign n36404 = \m1_addr_i[31]_pad  & ~n14271 ;
  assign n36405 = n14296 & n36404 ;
  assign n36406 = \m4_addr_i[31]_pad  & n14271 ;
  assign n36407 = n14288 & n36406 ;
  assign n36408 = ~n36405 & ~n36407 ;
  assign n36409 = n36403 & n36408 ;
  assign n36410 = \m2_addr_i[31]_pad  & n14271 ;
  assign n36411 = n14279 & n36410 ;
  assign n36412 = \m3_addr_i[31]_pad  & ~n14271 ;
  assign n36413 = n14279 & n36412 ;
  assign n36414 = ~n36411 & ~n36413 ;
  assign n36415 = \m0_addr_i[31]_pad  & n14271 ;
  assign n36416 = n14296 & n36415 ;
  assign n36417 = \m7_addr_i[31]_pad  & ~n14271 ;
  assign n36418 = n14264 & n36417 ;
  assign n36419 = ~n36416 & ~n36418 ;
  assign n36420 = n36414 & n36419 ;
  assign n36421 = n36409 & n36420 ;
  assign n36422 = \m3_addr_i[3]_pad  & ~n14271 ;
  assign n36423 = n14279 & n36422 ;
  assign n36424 = \m4_addr_i[3]_pad  & n14271 ;
  assign n36425 = n14288 & n36424 ;
  assign n36426 = ~n36423 & ~n36425 ;
  assign n36427 = \m6_addr_i[3]_pad  & n14271 ;
  assign n36428 = n14264 & n36427 ;
  assign n36429 = \m2_addr_i[3]_pad  & n14271 ;
  assign n36430 = n14279 & n36429 ;
  assign n36431 = ~n36428 & ~n36430 ;
  assign n36432 = n36426 & n36431 ;
  assign n36433 = \m5_addr_i[3]_pad  & ~n14271 ;
  assign n36434 = n14288 & n36433 ;
  assign n36435 = \m1_addr_i[3]_pad  & ~n14271 ;
  assign n36436 = n14296 & n36435 ;
  assign n36437 = ~n36434 & ~n36436 ;
  assign n36438 = \m0_addr_i[3]_pad  & n14271 ;
  assign n36439 = n14296 & n36438 ;
  assign n36440 = \m7_addr_i[3]_pad  & ~n14271 ;
  assign n36441 = n14264 & n36440 ;
  assign n36442 = ~n36439 & ~n36441 ;
  assign n36443 = n36437 & n36442 ;
  assign n36444 = n36432 & n36443 ;
  assign n36445 = \m3_addr_i[4]_pad  & ~n14271 ;
  assign n36446 = n14279 & n36445 ;
  assign n36447 = \m4_addr_i[4]_pad  & n14271 ;
  assign n36448 = n14288 & n36447 ;
  assign n36449 = ~n36446 & ~n36448 ;
  assign n36450 = \m6_addr_i[4]_pad  & n14271 ;
  assign n36451 = n14264 & n36450 ;
  assign n36452 = \m2_addr_i[4]_pad  & n14271 ;
  assign n36453 = n14279 & n36452 ;
  assign n36454 = ~n36451 & ~n36453 ;
  assign n36455 = n36449 & n36454 ;
  assign n36456 = \m5_addr_i[4]_pad  & ~n14271 ;
  assign n36457 = n14288 & n36456 ;
  assign n36458 = \m1_addr_i[4]_pad  & ~n14271 ;
  assign n36459 = n14296 & n36458 ;
  assign n36460 = ~n36457 & ~n36459 ;
  assign n36461 = \m0_addr_i[4]_pad  & n14271 ;
  assign n36462 = n14296 & n36461 ;
  assign n36463 = \m7_addr_i[4]_pad  & ~n14271 ;
  assign n36464 = n14264 & n36463 ;
  assign n36465 = ~n36462 & ~n36464 ;
  assign n36466 = n36460 & n36465 ;
  assign n36467 = n36455 & n36466 ;
  assign n36468 = \m3_addr_i[5]_pad  & ~n14271 ;
  assign n36469 = n14279 & n36468 ;
  assign n36470 = \m4_addr_i[5]_pad  & n14271 ;
  assign n36471 = n14288 & n36470 ;
  assign n36472 = ~n36469 & ~n36471 ;
  assign n36473 = \m6_addr_i[5]_pad  & n14271 ;
  assign n36474 = n14264 & n36473 ;
  assign n36475 = \m2_addr_i[5]_pad  & n14271 ;
  assign n36476 = n14279 & n36475 ;
  assign n36477 = ~n36474 & ~n36476 ;
  assign n36478 = n36472 & n36477 ;
  assign n36479 = \m5_addr_i[5]_pad  & ~n14271 ;
  assign n36480 = n14288 & n36479 ;
  assign n36481 = \m1_addr_i[5]_pad  & ~n14271 ;
  assign n36482 = n14296 & n36481 ;
  assign n36483 = ~n36480 & ~n36482 ;
  assign n36484 = \m0_addr_i[5]_pad  & n14271 ;
  assign n36485 = n14296 & n36484 ;
  assign n36486 = \m7_addr_i[5]_pad  & ~n14271 ;
  assign n36487 = n14264 & n36486 ;
  assign n36488 = ~n36485 & ~n36487 ;
  assign n36489 = n36483 & n36488 ;
  assign n36490 = n36478 & n36489 ;
  assign n36491 = \m3_addr_i[6]_pad  & ~n14271 ;
  assign n36492 = n14279 & n36491 ;
  assign n36493 = \m4_addr_i[6]_pad  & n14271 ;
  assign n36494 = n14288 & n36493 ;
  assign n36495 = ~n36492 & ~n36494 ;
  assign n36496 = \m6_addr_i[6]_pad  & n14271 ;
  assign n36497 = n14264 & n36496 ;
  assign n36498 = \m2_addr_i[6]_pad  & n14271 ;
  assign n36499 = n14279 & n36498 ;
  assign n36500 = ~n36497 & ~n36499 ;
  assign n36501 = n36495 & n36500 ;
  assign n36502 = \m5_addr_i[6]_pad  & ~n14271 ;
  assign n36503 = n14288 & n36502 ;
  assign n36504 = \m1_addr_i[6]_pad  & ~n14271 ;
  assign n36505 = n14296 & n36504 ;
  assign n36506 = ~n36503 & ~n36505 ;
  assign n36507 = \m0_addr_i[6]_pad  & n14271 ;
  assign n36508 = n14296 & n36507 ;
  assign n36509 = \m7_addr_i[6]_pad  & ~n14271 ;
  assign n36510 = n14264 & n36509 ;
  assign n36511 = ~n36508 & ~n36510 ;
  assign n36512 = n36506 & n36511 ;
  assign n36513 = n36501 & n36512 ;
  assign n36514 = \m3_addr_i[7]_pad  & ~n14271 ;
  assign n36515 = n14279 & n36514 ;
  assign n36516 = \m4_addr_i[7]_pad  & n14271 ;
  assign n36517 = n14288 & n36516 ;
  assign n36518 = ~n36515 & ~n36517 ;
  assign n36519 = \m6_addr_i[7]_pad  & n14271 ;
  assign n36520 = n14264 & n36519 ;
  assign n36521 = \m2_addr_i[7]_pad  & n14271 ;
  assign n36522 = n14279 & n36521 ;
  assign n36523 = ~n36520 & ~n36522 ;
  assign n36524 = n36518 & n36523 ;
  assign n36525 = \m5_addr_i[7]_pad  & ~n14271 ;
  assign n36526 = n14288 & n36525 ;
  assign n36527 = \m1_addr_i[7]_pad  & ~n14271 ;
  assign n36528 = n14296 & n36527 ;
  assign n36529 = ~n36526 & ~n36528 ;
  assign n36530 = \m0_addr_i[7]_pad  & n14271 ;
  assign n36531 = n14296 & n36530 ;
  assign n36532 = \m7_addr_i[7]_pad  & ~n14271 ;
  assign n36533 = n14264 & n36532 ;
  assign n36534 = ~n36531 & ~n36533 ;
  assign n36535 = n36529 & n36534 ;
  assign n36536 = n36524 & n36535 ;
  assign n36537 = \m3_addr_i[8]_pad  & ~n14271 ;
  assign n36538 = n14279 & n36537 ;
  assign n36539 = \m4_addr_i[8]_pad  & n14271 ;
  assign n36540 = n14288 & n36539 ;
  assign n36541 = ~n36538 & ~n36540 ;
  assign n36542 = \m6_addr_i[8]_pad  & n14271 ;
  assign n36543 = n14264 & n36542 ;
  assign n36544 = \m2_addr_i[8]_pad  & n14271 ;
  assign n36545 = n14279 & n36544 ;
  assign n36546 = ~n36543 & ~n36545 ;
  assign n36547 = n36541 & n36546 ;
  assign n36548 = \m5_addr_i[8]_pad  & ~n14271 ;
  assign n36549 = n14288 & n36548 ;
  assign n36550 = \m1_addr_i[8]_pad  & ~n14271 ;
  assign n36551 = n14296 & n36550 ;
  assign n36552 = ~n36549 & ~n36551 ;
  assign n36553 = \m0_addr_i[8]_pad  & n14271 ;
  assign n36554 = n14296 & n36553 ;
  assign n36555 = \m7_addr_i[8]_pad  & ~n14271 ;
  assign n36556 = n14264 & n36555 ;
  assign n36557 = ~n36554 & ~n36556 ;
  assign n36558 = n36552 & n36557 ;
  assign n36559 = n36547 & n36558 ;
  assign n36560 = \m3_addr_i[9]_pad  & ~n14271 ;
  assign n36561 = n14279 & n36560 ;
  assign n36562 = \m4_addr_i[9]_pad  & n14271 ;
  assign n36563 = n14288 & n36562 ;
  assign n36564 = ~n36561 & ~n36563 ;
  assign n36565 = \m6_addr_i[9]_pad  & n14271 ;
  assign n36566 = n14264 & n36565 ;
  assign n36567 = \m2_addr_i[9]_pad  & n14271 ;
  assign n36568 = n14279 & n36567 ;
  assign n36569 = ~n36566 & ~n36568 ;
  assign n36570 = n36564 & n36569 ;
  assign n36571 = \m5_addr_i[9]_pad  & ~n14271 ;
  assign n36572 = n14288 & n36571 ;
  assign n36573 = \m1_addr_i[9]_pad  & ~n14271 ;
  assign n36574 = n14296 & n36573 ;
  assign n36575 = ~n36572 & ~n36574 ;
  assign n36576 = \m0_addr_i[9]_pad  & n14271 ;
  assign n36577 = n14296 & n36576 ;
  assign n36578 = \m7_addr_i[9]_pad  & ~n14271 ;
  assign n36579 = n14264 & n36578 ;
  assign n36580 = ~n36577 & ~n36579 ;
  assign n36581 = n36575 & n36580 ;
  assign n36582 = n36570 & n36581 ;
  assign n36583 = \m1_data_i[0]_pad  & ~n14271 ;
  assign n36584 = n14296 & n36583 ;
  assign n36585 = \m2_data_i[0]_pad  & n14271 ;
  assign n36586 = n14279 & n36585 ;
  assign n36587 = ~n36584 & ~n36586 ;
  assign n36588 = \m0_data_i[0]_pad  & n14271 ;
  assign n36589 = n14296 & n36588 ;
  assign n36590 = \m4_data_i[0]_pad  & n14271 ;
  assign n36591 = n14288 & n36590 ;
  assign n36592 = ~n36589 & ~n36591 ;
  assign n36593 = n36587 & n36592 ;
  assign n36594 = \m7_data_i[0]_pad  & ~n14271 ;
  assign n36595 = n14264 & n36594 ;
  assign n36596 = \m3_data_i[0]_pad  & ~n14271 ;
  assign n36597 = n14279 & n36596 ;
  assign n36598 = ~n36595 & ~n36597 ;
  assign n36599 = \m6_data_i[0]_pad  & n14271 ;
  assign n36600 = n14264 & n36599 ;
  assign n36601 = \m5_data_i[0]_pad  & ~n14271 ;
  assign n36602 = n14288 & n36601 ;
  assign n36603 = ~n36600 & ~n36602 ;
  assign n36604 = n36598 & n36603 ;
  assign n36605 = n36593 & n36604 ;
  assign n36606 = \m6_data_i[10]_pad  & n14271 ;
  assign n36607 = n14264 & n36606 ;
  assign n36608 = \m5_data_i[10]_pad  & ~n14271 ;
  assign n36609 = n14288 & n36608 ;
  assign n36610 = ~n36607 & ~n36609 ;
  assign n36611 = \m1_data_i[10]_pad  & ~n14271 ;
  assign n36612 = n14296 & n36611 ;
  assign n36613 = \m4_data_i[10]_pad  & n14271 ;
  assign n36614 = n14288 & n36613 ;
  assign n36615 = ~n36612 & ~n36614 ;
  assign n36616 = n36610 & n36615 ;
  assign n36617 = \m2_data_i[10]_pad  & n14271 ;
  assign n36618 = n14279 & n36617 ;
  assign n36619 = \m3_data_i[10]_pad  & ~n14271 ;
  assign n36620 = n14279 & n36619 ;
  assign n36621 = ~n36618 & ~n36620 ;
  assign n36622 = \m0_data_i[10]_pad  & n14271 ;
  assign n36623 = n14296 & n36622 ;
  assign n36624 = \m7_data_i[10]_pad  & ~n14271 ;
  assign n36625 = n14264 & n36624 ;
  assign n36626 = ~n36623 & ~n36625 ;
  assign n36627 = n36621 & n36626 ;
  assign n36628 = n36616 & n36627 ;
  assign n36629 = \m6_data_i[11]_pad  & n14271 ;
  assign n36630 = n14264 & n36629 ;
  assign n36631 = \m5_data_i[11]_pad  & ~n14271 ;
  assign n36632 = n14288 & n36631 ;
  assign n36633 = ~n36630 & ~n36632 ;
  assign n36634 = \m3_data_i[11]_pad  & ~n14271 ;
  assign n36635 = n14279 & n36634 ;
  assign n36636 = \m2_data_i[11]_pad  & n14271 ;
  assign n36637 = n14279 & n36636 ;
  assign n36638 = ~n36635 & ~n36637 ;
  assign n36639 = n36633 & n36638 ;
  assign n36640 = \m4_data_i[11]_pad  & n14271 ;
  assign n36641 = n14288 & n36640 ;
  assign n36642 = \m1_data_i[11]_pad  & ~n14271 ;
  assign n36643 = n14296 & n36642 ;
  assign n36644 = ~n36641 & ~n36643 ;
  assign n36645 = \m0_data_i[11]_pad  & n14271 ;
  assign n36646 = n14296 & n36645 ;
  assign n36647 = \m7_data_i[11]_pad  & ~n14271 ;
  assign n36648 = n14264 & n36647 ;
  assign n36649 = ~n36646 & ~n36648 ;
  assign n36650 = n36644 & n36649 ;
  assign n36651 = n36639 & n36650 ;
  assign n36652 = \m0_data_i[12]_pad  & n14271 ;
  assign n36653 = n14296 & n36652 ;
  assign n36654 = \m7_data_i[12]_pad  & ~n14271 ;
  assign n36655 = n14264 & n36654 ;
  assign n36656 = ~n36653 & ~n36655 ;
  assign n36657 = \m6_data_i[12]_pad  & n14271 ;
  assign n36658 = n14264 & n36657 ;
  assign n36659 = \m4_data_i[12]_pad  & n14271 ;
  assign n36660 = n14288 & n36659 ;
  assign n36661 = ~n36658 & ~n36660 ;
  assign n36662 = n36656 & n36661 ;
  assign n36663 = \m5_data_i[12]_pad  & ~n14271 ;
  assign n36664 = n14288 & n36663 ;
  assign n36665 = \m3_data_i[12]_pad  & ~n14271 ;
  assign n36666 = n14279 & n36665 ;
  assign n36667 = ~n36664 & ~n36666 ;
  assign n36668 = \m1_data_i[12]_pad  & ~n14271 ;
  assign n36669 = n14296 & n36668 ;
  assign n36670 = \m2_data_i[12]_pad  & n14271 ;
  assign n36671 = n14279 & n36670 ;
  assign n36672 = ~n36669 & ~n36671 ;
  assign n36673 = n36667 & n36672 ;
  assign n36674 = n36662 & n36673 ;
  assign n36675 = \m3_data_i[13]_pad  & ~n14271 ;
  assign n36676 = n14279 & n36675 ;
  assign n36677 = \m4_data_i[13]_pad  & n14271 ;
  assign n36678 = n14288 & n36677 ;
  assign n36679 = ~n36676 & ~n36678 ;
  assign n36680 = \m0_data_i[13]_pad  & n14271 ;
  assign n36681 = n14296 & n36680 ;
  assign n36682 = \m5_data_i[13]_pad  & ~n14271 ;
  assign n36683 = n14288 & n36682 ;
  assign n36684 = ~n36681 & ~n36683 ;
  assign n36685 = n36679 & n36684 ;
  assign n36686 = \m7_data_i[13]_pad  & ~n14271 ;
  assign n36687 = n14264 & n36686 ;
  assign n36688 = \m6_data_i[13]_pad  & n14271 ;
  assign n36689 = n14264 & n36688 ;
  assign n36690 = ~n36687 & ~n36689 ;
  assign n36691 = \m1_data_i[13]_pad  & ~n14271 ;
  assign n36692 = n14296 & n36691 ;
  assign n36693 = \m2_data_i[13]_pad  & n14271 ;
  assign n36694 = n14279 & n36693 ;
  assign n36695 = ~n36692 & ~n36694 ;
  assign n36696 = n36690 & n36695 ;
  assign n36697 = n36685 & n36696 ;
  assign n36698 = \m6_data_i[14]_pad  & n14271 ;
  assign n36699 = n14264 & n36698 ;
  assign n36700 = \m5_data_i[14]_pad  & ~n14271 ;
  assign n36701 = n14288 & n36700 ;
  assign n36702 = ~n36699 & ~n36701 ;
  assign n36703 = \m1_data_i[14]_pad  & ~n14271 ;
  assign n36704 = n14296 & n36703 ;
  assign n36705 = \m4_data_i[14]_pad  & n14271 ;
  assign n36706 = n14288 & n36705 ;
  assign n36707 = ~n36704 & ~n36706 ;
  assign n36708 = n36702 & n36707 ;
  assign n36709 = \m2_data_i[14]_pad  & n14271 ;
  assign n36710 = n14279 & n36709 ;
  assign n36711 = \m3_data_i[14]_pad  & ~n14271 ;
  assign n36712 = n14279 & n36711 ;
  assign n36713 = ~n36710 & ~n36712 ;
  assign n36714 = \m0_data_i[14]_pad  & n14271 ;
  assign n36715 = n14296 & n36714 ;
  assign n36716 = \m7_data_i[14]_pad  & ~n14271 ;
  assign n36717 = n14264 & n36716 ;
  assign n36718 = ~n36715 & ~n36717 ;
  assign n36719 = n36713 & n36718 ;
  assign n36720 = n36708 & n36719 ;
  assign n36721 = \m3_data_i[15]_pad  & ~n14271 ;
  assign n36722 = n14279 & n36721 ;
  assign n36723 = \m4_data_i[15]_pad  & n14271 ;
  assign n36724 = n14288 & n36723 ;
  assign n36725 = ~n36722 & ~n36724 ;
  assign n36726 = \m0_data_i[15]_pad  & n14271 ;
  assign n36727 = n14296 & n36726 ;
  assign n36728 = \m2_data_i[15]_pad  & n14271 ;
  assign n36729 = n14279 & n36728 ;
  assign n36730 = ~n36727 & ~n36729 ;
  assign n36731 = n36725 & n36730 ;
  assign n36732 = \m7_data_i[15]_pad  & ~n14271 ;
  assign n36733 = n14264 & n36732 ;
  assign n36734 = \m1_data_i[15]_pad  & ~n14271 ;
  assign n36735 = n14296 & n36734 ;
  assign n36736 = ~n36733 & ~n36735 ;
  assign n36737 = \m6_data_i[15]_pad  & n14271 ;
  assign n36738 = n14264 & n36737 ;
  assign n36739 = \m5_data_i[15]_pad  & ~n14271 ;
  assign n36740 = n14288 & n36739 ;
  assign n36741 = ~n36738 & ~n36740 ;
  assign n36742 = n36736 & n36741 ;
  assign n36743 = n36731 & n36742 ;
  assign n36744 = \m1_data_i[16]_pad  & ~n14271 ;
  assign n36745 = n14296 & n36744 ;
  assign n36746 = \m2_data_i[16]_pad  & n14271 ;
  assign n36747 = n14279 & n36746 ;
  assign n36748 = ~n36745 & ~n36747 ;
  assign n36749 = \m0_data_i[16]_pad  & n14271 ;
  assign n36750 = n14296 & n36749 ;
  assign n36751 = \m5_data_i[16]_pad  & ~n14271 ;
  assign n36752 = n14288 & n36751 ;
  assign n36753 = ~n36750 & ~n36752 ;
  assign n36754 = n36748 & n36753 ;
  assign n36755 = \m7_data_i[16]_pad  & ~n14271 ;
  assign n36756 = n14264 & n36755 ;
  assign n36757 = \m6_data_i[16]_pad  & n14271 ;
  assign n36758 = n14264 & n36757 ;
  assign n36759 = ~n36756 & ~n36758 ;
  assign n36760 = \m3_data_i[16]_pad  & ~n14271 ;
  assign n36761 = n14279 & n36760 ;
  assign n36762 = \m4_data_i[16]_pad  & n14271 ;
  assign n36763 = n14288 & n36762 ;
  assign n36764 = ~n36761 & ~n36763 ;
  assign n36765 = n36759 & n36764 ;
  assign n36766 = n36754 & n36765 ;
  assign n36767 = \m3_data_i[17]_pad  & ~n14271 ;
  assign n36768 = n14279 & n36767 ;
  assign n36769 = \m4_data_i[17]_pad  & n14271 ;
  assign n36770 = n14288 & n36769 ;
  assign n36771 = ~n36768 & ~n36770 ;
  assign n36772 = \m0_data_i[17]_pad  & n14271 ;
  assign n36773 = n14296 & n36772 ;
  assign n36774 = \m2_data_i[17]_pad  & n14271 ;
  assign n36775 = n14279 & n36774 ;
  assign n36776 = ~n36773 & ~n36775 ;
  assign n36777 = n36771 & n36776 ;
  assign n36778 = \m7_data_i[17]_pad  & ~n14271 ;
  assign n36779 = n14264 & n36778 ;
  assign n36780 = \m1_data_i[17]_pad  & ~n14271 ;
  assign n36781 = n14296 & n36780 ;
  assign n36782 = ~n36779 & ~n36781 ;
  assign n36783 = \m6_data_i[17]_pad  & n14271 ;
  assign n36784 = n14264 & n36783 ;
  assign n36785 = \m5_data_i[17]_pad  & ~n14271 ;
  assign n36786 = n14288 & n36785 ;
  assign n36787 = ~n36784 & ~n36786 ;
  assign n36788 = n36782 & n36787 ;
  assign n36789 = n36777 & n36788 ;
  assign n36790 = \m3_data_i[18]_pad  & ~n14271 ;
  assign n36791 = n14279 & n36790 ;
  assign n36792 = \m4_data_i[18]_pad  & n14271 ;
  assign n36793 = n14288 & n36792 ;
  assign n36794 = ~n36791 & ~n36793 ;
  assign n36795 = \m0_data_i[18]_pad  & n14271 ;
  assign n36796 = n14296 & n36795 ;
  assign n36797 = \m2_data_i[18]_pad  & n14271 ;
  assign n36798 = n14279 & n36797 ;
  assign n36799 = ~n36796 & ~n36798 ;
  assign n36800 = n36794 & n36799 ;
  assign n36801 = \m7_data_i[18]_pad  & ~n14271 ;
  assign n36802 = n14264 & n36801 ;
  assign n36803 = \m1_data_i[18]_pad  & ~n14271 ;
  assign n36804 = n14296 & n36803 ;
  assign n36805 = ~n36802 & ~n36804 ;
  assign n36806 = \m6_data_i[18]_pad  & n14271 ;
  assign n36807 = n14264 & n36806 ;
  assign n36808 = \m5_data_i[18]_pad  & ~n14271 ;
  assign n36809 = n14288 & n36808 ;
  assign n36810 = ~n36807 & ~n36809 ;
  assign n36811 = n36805 & n36810 ;
  assign n36812 = n36800 & n36811 ;
  assign n36813 = \m3_data_i[19]_pad  & ~n14271 ;
  assign n36814 = n14279 & n36813 ;
  assign n36815 = \m4_data_i[19]_pad  & n14271 ;
  assign n36816 = n14288 & n36815 ;
  assign n36817 = ~n36814 & ~n36816 ;
  assign n36818 = \m6_data_i[19]_pad  & n14271 ;
  assign n36819 = n14264 & n36818 ;
  assign n36820 = \m2_data_i[19]_pad  & n14271 ;
  assign n36821 = n14279 & n36820 ;
  assign n36822 = ~n36819 & ~n36821 ;
  assign n36823 = n36817 & n36822 ;
  assign n36824 = \m5_data_i[19]_pad  & ~n14271 ;
  assign n36825 = n14288 & n36824 ;
  assign n36826 = \m1_data_i[19]_pad  & ~n14271 ;
  assign n36827 = n14296 & n36826 ;
  assign n36828 = ~n36825 & ~n36827 ;
  assign n36829 = \m0_data_i[19]_pad  & n14271 ;
  assign n36830 = n14296 & n36829 ;
  assign n36831 = \m7_data_i[19]_pad  & ~n14271 ;
  assign n36832 = n14264 & n36831 ;
  assign n36833 = ~n36830 & ~n36832 ;
  assign n36834 = n36828 & n36833 ;
  assign n36835 = n36823 & n36834 ;
  assign n36836 = \m3_data_i[1]_pad  & ~n14271 ;
  assign n36837 = n14279 & n36836 ;
  assign n36838 = \m4_data_i[1]_pad  & n14271 ;
  assign n36839 = n14288 & n36838 ;
  assign n36840 = ~n36837 & ~n36839 ;
  assign n36841 = \m1_data_i[1]_pad  & ~n14271 ;
  assign n36842 = n14296 & n36841 ;
  assign n36843 = \m5_data_i[1]_pad  & ~n14271 ;
  assign n36844 = n14288 & n36843 ;
  assign n36845 = ~n36842 & ~n36844 ;
  assign n36846 = n36840 & n36845 ;
  assign n36847 = \m2_data_i[1]_pad  & n14271 ;
  assign n36848 = n14279 & n36847 ;
  assign n36849 = \m6_data_i[1]_pad  & n14271 ;
  assign n36850 = n14264 & n36849 ;
  assign n36851 = ~n36848 & ~n36850 ;
  assign n36852 = \m0_data_i[1]_pad  & n14271 ;
  assign n36853 = n14296 & n36852 ;
  assign n36854 = \m7_data_i[1]_pad  & ~n14271 ;
  assign n36855 = n14264 & n36854 ;
  assign n36856 = ~n36853 & ~n36855 ;
  assign n36857 = n36851 & n36856 ;
  assign n36858 = n36846 & n36857 ;
  assign n36859 = \m3_data_i[20]_pad  & ~n14271 ;
  assign n36860 = n14279 & n36859 ;
  assign n36861 = \m4_data_i[20]_pad  & n14271 ;
  assign n36862 = n14288 & n36861 ;
  assign n36863 = ~n36860 & ~n36862 ;
  assign n36864 = \m1_data_i[20]_pad  & ~n14271 ;
  assign n36865 = n14296 & n36864 ;
  assign n36866 = \m5_data_i[20]_pad  & ~n14271 ;
  assign n36867 = n14288 & n36866 ;
  assign n36868 = ~n36865 & ~n36867 ;
  assign n36869 = n36863 & n36868 ;
  assign n36870 = \m2_data_i[20]_pad  & n14271 ;
  assign n36871 = n14279 & n36870 ;
  assign n36872 = \m6_data_i[20]_pad  & n14271 ;
  assign n36873 = n14264 & n36872 ;
  assign n36874 = ~n36871 & ~n36873 ;
  assign n36875 = \m0_data_i[20]_pad  & n14271 ;
  assign n36876 = n14296 & n36875 ;
  assign n36877 = \m7_data_i[20]_pad  & ~n14271 ;
  assign n36878 = n14264 & n36877 ;
  assign n36879 = ~n36876 & ~n36878 ;
  assign n36880 = n36874 & n36879 ;
  assign n36881 = n36869 & n36880 ;
  assign n36882 = \m6_data_i[21]_pad  & n14271 ;
  assign n36883 = n14264 & n36882 ;
  assign n36884 = \m5_data_i[21]_pad  & ~n14271 ;
  assign n36885 = n14288 & n36884 ;
  assign n36886 = ~n36883 & ~n36885 ;
  assign n36887 = \m0_data_i[21]_pad  & n14271 ;
  assign n36888 = n14296 & n36887 ;
  assign n36889 = \m4_data_i[21]_pad  & n14271 ;
  assign n36890 = n14288 & n36889 ;
  assign n36891 = ~n36888 & ~n36890 ;
  assign n36892 = n36886 & n36891 ;
  assign n36893 = \m7_data_i[21]_pad  & ~n14271 ;
  assign n36894 = n14264 & n36893 ;
  assign n36895 = \m3_data_i[21]_pad  & ~n14271 ;
  assign n36896 = n14279 & n36895 ;
  assign n36897 = ~n36894 & ~n36896 ;
  assign n36898 = \m1_data_i[21]_pad  & ~n14271 ;
  assign n36899 = n14296 & n36898 ;
  assign n36900 = \m2_data_i[21]_pad  & n14271 ;
  assign n36901 = n14279 & n36900 ;
  assign n36902 = ~n36899 & ~n36901 ;
  assign n36903 = n36897 & n36902 ;
  assign n36904 = n36892 & n36903 ;
  assign n36905 = \m3_data_i[22]_pad  & ~n14271 ;
  assign n36906 = n14279 & n36905 ;
  assign n36907 = \m4_data_i[22]_pad  & n14271 ;
  assign n36908 = n14288 & n36907 ;
  assign n36909 = ~n36906 & ~n36908 ;
  assign n36910 = \m6_data_i[22]_pad  & n14271 ;
  assign n36911 = n14264 & n36910 ;
  assign n36912 = \m2_data_i[22]_pad  & n14271 ;
  assign n36913 = n14279 & n36912 ;
  assign n36914 = ~n36911 & ~n36913 ;
  assign n36915 = n36909 & n36914 ;
  assign n36916 = \m5_data_i[22]_pad  & ~n14271 ;
  assign n36917 = n14288 & n36916 ;
  assign n36918 = \m1_data_i[22]_pad  & ~n14271 ;
  assign n36919 = n14296 & n36918 ;
  assign n36920 = ~n36917 & ~n36919 ;
  assign n36921 = \m0_data_i[22]_pad  & n14271 ;
  assign n36922 = n14296 & n36921 ;
  assign n36923 = \m7_data_i[22]_pad  & ~n14271 ;
  assign n36924 = n14264 & n36923 ;
  assign n36925 = ~n36922 & ~n36924 ;
  assign n36926 = n36920 & n36925 ;
  assign n36927 = n36915 & n36926 ;
  assign n36928 = \m0_data_i[23]_pad  & n14271 ;
  assign n36929 = n14296 & n36928 ;
  assign n36930 = \m7_data_i[23]_pad  & ~n14271 ;
  assign n36931 = n14264 & n36930 ;
  assign n36932 = ~n36929 & ~n36931 ;
  assign n36933 = \m1_data_i[23]_pad  & ~n14271 ;
  assign n36934 = n14296 & n36933 ;
  assign n36935 = \m5_data_i[23]_pad  & ~n14271 ;
  assign n36936 = n14288 & n36935 ;
  assign n36937 = ~n36934 & ~n36936 ;
  assign n36938 = n36932 & n36937 ;
  assign n36939 = \m2_data_i[23]_pad  & n14271 ;
  assign n36940 = n14279 & n36939 ;
  assign n36941 = \m6_data_i[23]_pad  & n14271 ;
  assign n36942 = n14264 & n36941 ;
  assign n36943 = ~n36940 & ~n36942 ;
  assign n36944 = \m3_data_i[23]_pad  & ~n14271 ;
  assign n36945 = n14279 & n36944 ;
  assign n36946 = \m4_data_i[23]_pad  & n14271 ;
  assign n36947 = n14288 & n36946 ;
  assign n36948 = ~n36945 & ~n36947 ;
  assign n36949 = n36943 & n36948 ;
  assign n36950 = n36938 & n36949 ;
  assign n36951 = \m1_data_i[24]_pad  & ~n14271 ;
  assign n36952 = n14296 & n36951 ;
  assign n36953 = \m2_data_i[24]_pad  & n14271 ;
  assign n36954 = n14279 & n36953 ;
  assign n36955 = ~n36952 & ~n36954 ;
  assign n36956 = \m6_data_i[24]_pad  & n14271 ;
  assign n36957 = n14264 & n36956 ;
  assign n36958 = \m4_data_i[24]_pad  & n14271 ;
  assign n36959 = n14288 & n36958 ;
  assign n36960 = ~n36957 & ~n36959 ;
  assign n36961 = n36955 & n36960 ;
  assign n36962 = \m5_data_i[24]_pad  & ~n14271 ;
  assign n36963 = n14288 & n36962 ;
  assign n36964 = \m3_data_i[24]_pad  & ~n14271 ;
  assign n36965 = n14279 & n36964 ;
  assign n36966 = ~n36963 & ~n36965 ;
  assign n36967 = \m0_data_i[24]_pad  & n14271 ;
  assign n36968 = n14296 & n36967 ;
  assign n36969 = \m7_data_i[24]_pad  & ~n14271 ;
  assign n36970 = n14264 & n36969 ;
  assign n36971 = ~n36968 & ~n36970 ;
  assign n36972 = n36966 & n36971 ;
  assign n36973 = n36961 & n36972 ;
  assign n36974 = \m6_data_i[25]_pad  & n14271 ;
  assign n36975 = n14264 & n36974 ;
  assign n36976 = \m5_data_i[25]_pad  & ~n14271 ;
  assign n36977 = n14288 & n36976 ;
  assign n36978 = ~n36975 & ~n36977 ;
  assign n36979 = \m0_data_i[25]_pad  & n14271 ;
  assign n36980 = n14296 & n36979 ;
  assign n36981 = \m4_data_i[25]_pad  & n14271 ;
  assign n36982 = n14288 & n36981 ;
  assign n36983 = ~n36980 & ~n36982 ;
  assign n36984 = n36978 & n36983 ;
  assign n36985 = \m7_data_i[25]_pad  & ~n14271 ;
  assign n36986 = n14264 & n36985 ;
  assign n36987 = \m3_data_i[25]_pad  & ~n14271 ;
  assign n36988 = n14279 & n36987 ;
  assign n36989 = ~n36986 & ~n36988 ;
  assign n36990 = \m1_data_i[25]_pad  & ~n14271 ;
  assign n36991 = n14296 & n36990 ;
  assign n36992 = \m2_data_i[25]_pad  & n14271 ;
  assign n36993 = n14279 & n36992 ;
  assign n36994 = ~n36991 & ~n36993 ;
  assign n36995 = n36989 & n36994 ;
  assign n36996 = n36984 & n36995 ;
  assign n36997 = \m1_data_i[26]_pad  & ~n14271 ;
  assign n36998 = n14296 & n36997 ;
  assign n36999 = \m2_data_i[26]_pad  & n14271 ;
  assign n37000 = n14279 & n36999 ;
  assign n37001 = ~n36998 & ~n37000 ;
  assign n37002 = \m3_data_i[26]_pad  & ~n14271 ;
  assign n37003 = n14279 & n37002 ;
  assign n37004 = \m5_data_i[26]_pad  & ~n14271 ;
  assign n37005 = n14288 & n37004 ;
  assign n37006 = ~n37003 & ~n37005 ;
  assign n37007 = n37001 & n37006 ;
  assign n37008 = \m4_data_i[26]_pad  & n14271 ;
  assign n37009 = n14288 & n37008 ;
  assign n37010 = \m6_data_i[26]_pad  & n14271 ;
  assign n37011 = n14264 & n37010 ;
  assign n37012 = ~n37009 & ~n37011 ;
  assign n37013 = \m0_data_i[26]_pad  & n14271 ;
  assign n37014 = n14296 & n37013 ;
  assign n37015 = \m7_data_i[26]_pad  & ~n14271 ;
  assign n37016 = n14264 & n37015 ;
  assign n37017 = ~n37014 & ~n37016 ;
  assign n37018 = n37012 & n37017 ;
  assign n37019 = n37007 & n37018 ;
  assign n37020 = \m0_data_i[27]_pad  & n14271 ;
  assign n37021 = n14296 & n37020 ;
  assign n37022 = \m7_data_i[27]_pad  & ~n14271 ;
  assign n37023 = n14264 & n37022 ;
  assign n37024 = ~n37021 & ~n37023 ;
  assign n37025 = \m3_data_i[27]_pad  & ~n14271 ;
  assign n37026 = n14279 & n37025 ;
  assign n37027 = \m2_data_i[27]_pad  & n14271 ;
  assign n37028 = n14279 & n37027 ;
  assign n37029 = ~n37026 & ~n37028 ;
  assign n37030 = n37024 & n37029 ;
  assign n37031 = \m4_data_i[27]_pad  & n14271 ;
  assign n37032 = n14288 & n37031 ;
  assign n37033 = \m1_data_i[27]_pad  & ~n14271 ;
  assign n37034 = n14296 & n37033 ;
  assign n37035 = ~n37032 & ~n37034 ;
  assign n37036 = \m6_data_i[27]_pad  & n14271 ;
  assign n37037 = n14264 & n37036 ;
  assign n37038 = \m5_data_i[27]_pad  & ~n14271 ;
  assign n37039 = n14288 & n37038 ;
  assign n37040 = ~n37037 & ~n37039 ;
  assign n37041 = n37035 & n37040 ;
  assign n37042 = n37030 & n37041 ;
  assign n37043 = \m1_data_i[28]_pad  & ~n14271 ;
  assign n37044 = n14296 & n37043 ;
  assign n37045 = \m2_data_i[28]_pad  & n14271 ;
  assign n37046 = n14279 & n37045 ;
  assign n37047 = ~n37044 & ~n37046 ;
  assign n37048 = \m0_data_i[28]_pad  & n14271 ;
  assign n37049 = n14296 & n37048 ;
  assign n37050 = \m5_data_i[28]_pad  & ~n14271 ;
  assign n37051 = n14288 & n37050 ;
  assign n37052 = ~n37049 & ~n37051 ;
  assign n37053 = n37047 & n37052 ;
  assign n37054 = \m7_data_i[28]_pad  & ~n14271 ;
  assign n37055 = n14264 & n37054 ;
  assign n37056 = \m6_data_i[28]_pad  & n14271 ;
  assign n37057 = n14264 & n37056 ;
  assign n37058 = ~n37055 & ~n37057 ;
  assign n37059 = \m3_data_i[28]_pad  & ~n14271 ;
  assign n37060 = n14279 & n37059 ;
  assign n37061 = \m4_data_i[28]_pad  & n14271 ;
  assign n37062 = n14288 & n37061 ;
  assign n37063 = ~n37060 & ~n37062 ;
  assign n37064 = n37058 & n37063 ;
  assign n37065 = n37053 & n37064 ;
  assign n37066 = \m1_data_i[29]_pad  & ~n14271 ;
  assign n37067 = n14296 & n37066 ;
  assign n37068 = \m2_data_i[29]_pad  & n14271 ;
  assign n37069 = n14279 & n37068 ;
  assign n37070 = ~n37067 & ~n37069 ;
  assign n37071 = \m0_data_i[29]_pad  & n14271 ;
  assign n37072 = n14296 & n37071 ;
  assign n37073 = \m4_data_i[29]_pad  & n14271 ;
  assign n37074 = n14288 & n37073 ;
  assign n37075 = ~n37072 & ~n37074 ;
  assign n37076 = n37070 & n37075 ;
  assign n37077 = \m7_data_i[29]_pad  & ~n14271 ;
  assign n37078 = n14264 & n37077 ;
  assign n37079 = \m3_data_i[29]_pad  & ~n14271 ;
  assign n37080 = n14279 & n37079 ;
  assign n37081 = ~n37078 & ~n37080 ;
  assign n37082 = \m6_data_i[29]_pad  & n14271 ;
  assign n37083 = n14264 & n37082 ;
  assign n37084 = \m5_data_i[29]_pad  & ~n14271 ;
  assign n37085 = n14288 & n37084 ;
  assign n37086 = ~n37083 & ~n37085 ;
  assign n37087 = n37081 & n37086 ;
  assign n37088 = n37076 & n37087 ;
  assign n37089 = \m6_data_i[2]_pad  & n14271 ;
  assign n37090 = n14264 & n37089 ;
  assign n37091 = \m5_data_i[2]_pad  & ~n14271 ;
  assign n37092 = n14288 & n37091 ;
  assign n37093 = ~n37090 & ~n37092 ;
  assign n37094 = \m3_data_i[2]_pad  & ~n14271 ;
  assign n37095 = n14279 & n37094 ;
  assign n37096 = \m7_data_i[2]_pad  & ~n14271 ;
  assign n37097 = n14264 & n37096 ;
  assign n37098 = ~n37095 & ~n37097 ;
  assign n37099 = n37093 & n37098 ;
  assign n37100 = \m4_data_i[2]_pad  & n14271 ;
  assign n37101 = n14288 & n37100 ;
  assign n37102 = \m0_data_i[2]_pad  & n14271 ;
  assign n37103 = n14296 & n37102 ;
  assign n37104 = ~n37101 & ~n37103 ;
  assign n37105 = \m1_data_i[2]_pad  & ~n14271 ;
  assign n37106 = n14296 & n37105 ;
  assign n37107 = \m2_data_i[2]_pad  & n14271 ;
  assign n37108 = n14279 & n37107 ;
  assign n37109 = ~n37106 & ~n37108 ;
  assign n37110 = n37104 & n37109 ;
  assign n37111 = n37099 & n37110 ;
  assign n37112 = \m1_data_i[30]_pad  & ~n14271 ;
  assign n37113 = n14296 & n37112 ;
  assign n37114 = \m2_data_i[30]_pad  & n14271 ;
  assign n37115 = n14279 & n37114 ;
  assign n37116 = ~n37113 & ~n37115 ;
  assign n37117 = \m0_data_i[30]_pad  & n14271 ;
  assign n37118 = n14296 & n37117 ;
  assign n37119 = \m4_data_i[30]_pad  & n14271 ;
  assign n37120 = n14288 & n37119 ;
  assign n37121 = ~n37118 & ~n37120 ;
  assign n37122 = n37116 & n37121 ;
  assign n37123 = \m7_data_i[30]_pad  & ~n14271 ;
  assign n37124 = n14264 & n37123 ;
  assign n37125 = \m3_data_i[30]_pad  & ~n14271 ;
  assign n37126 = n14279 & n37125 ;
  assign n37127 = ~n37124 & ~n37126 ;
  assign n37128 = \m6_data_i[30]_pad  & n14271 ;
  assign n37129 = n14264 & n37128 ;
  assign n37130 = \m5_data_i[30]_pad  & ~n14271 ;
  assign n37131 = n14288 & n37130 ;
  assign n37132 = ~n37129 & ~n37131 ;
  assign n37133 = n37127 & n37132 ;
  assign n37134 = n37122 & n37133 ;
  assign n37135 = \m0_data_i[31]_pad  & n14271 ;
  assign n37136 = n14296 & n37135 ;
  assign n37137 = \m7_data_i[31]_pad  & ~n14271 ;
  assign n37138 = n14264 & n37137 ;
  assign n37139 = ~n37136 & ~n37138 ;
  assign n37140 = \m1_data_i[31]_pad  & ~n14271 ;
  assign n37141 = n14296 & n37140 ;
  assign n37142 = \m4_data_i[31]_pad  & n14271 ;
  assign n37143 = n14288 & n37142 ;
  assign n37144 = ~n37141 & ~n37143 ;
  assign n37145 = n37139 & n37144 ;
  assign n37146 = \m2_data_i[31]_pad  & n14271 ;
  assign n37147 = n14279 & n37146 ;
  assign n37148 = \m3_data_i[31]_pad  & ~n14271 ;
  assign n37149 = n14279 & n37148 ;
  assign n37150 = ~n37147 & ~n37149 ;
  assign n37151 = \m6_data_i[31]_pad  & n14271 ;
  assign n37152 = n14264 & n37151 ;
  assign n37153 = \m5_data_i[31]_pad  & ~n14271 ;
  assign n37154 = n14288 & n37153 ;
  assign n37155 = ~n37152 & ~n37154 ;
  assign n37156 = n37150 & n37155 ;
  assign n37157 = n37145 & n37156 ;
  assign n37158 = \m1_data_i[3]_pad  & ~n14271 ;
  assign n37159 = n14296 & n37158 ;
  assign n37160 = \m2_data_i[3]_pad  & n14271 ;
  assign n37161 = n14279 & n37160 ;
  assign n37162 = ~n37159 & ~n37161 ;
  assign n37163 = \m0_data_i[3]_pad  & n14271 ;
  assign n37164 = n14296 & n37163 ;
  assign n37165 = \m5_data_i[3]_pad  & ~n14271 ;
  assign n37166 = n14288 & n37165 ;
  assign n37167 = ~n37164 & ~n37166 ;
  assign n37168 = n37162 & n37167 ;
  assign n37169 = \m7_data_i[3]_pad  & ~n14271 ;
  assign n37170 = n14264 & n37169 ;
  assign n37171 = \m6_data_i[3]_pad  & n14271 ;
  assign n37172 = n14264 & n37171 ;
  assign n37173 = ~n37170 & ~n37172 ;
  assign n37174 = \m3_data_i[3]_pad  & ~n14271 ;
  assign n37175 = n14279 & n37174 ;
  assign n37176 = \m4_data_i[3]_pad  & n14271 ;
  assign n37177 = n14288 & n37176 ;
  assign n37178 = ~n37175 & ~n37177 ;
  assign n37179 = n37173 & n37178 ;
  assign n37180 = n37168 & n37179 ;
  assign n37181 = \m3_data_i[4]_pad  & ~n14271 ;
  assign n37182 = n14279 & n37181 ;
  assign n37183 = \m4_data_i[4]_pad  & n14271 ;
  assign n37184 = n14288 & n37183 ;
  assign n37185 = ~n37182 & ~n37184 ;
  assign n37186 = \m1_data_i[4]_pad  & ~n14271 ;
  assign n37187 = n14296 & n37186 ;
  assign n37188 = \m5_data_i[4]_pad  & ~n14271 ;
  assign n37189 = n14288 & n37188 ;
  assign n37190 = ~n37187 & ~n37189 ;
  assign n37191 = n37185 & n37190 ;
  assign n37192 = \m2_data_i[4]_pad  & n14271 ;
  assign n37193 = n14279 & n37192 ;
  assign n37194 = \m6_data_i[4]_pad  & n14271 ;
  assign n37195 = n14264 & n37194 ;
  assign n37196 = ~n37193 & ~n37195 ;
  assign n37197 = \m0_data_i[4]_pad  & n14271 ;
  assign n37198 = n14296 & n37197 ;
  assign n37199 = \m7_data_i[4]_pad  & ~n14271 ;
  assign n37200 = n14264 & n37199 ;
  assign n37201 = ~n37198 & ~n37200 ;
  assign n37202 = n37196 & n37201 ;
  assign n37203 = n37191 & n37202 ;
  assign n37204 = \m6_data_i[5]_pad  & n14271 ;
  assign n37205 = n14264 & n37204 ;
  assign n37206 = \m5_data_i[5]_pad  & ~n14271 ;
  assign n37207 = n14288 & n37206 ;
  assign n37208 = ~n37205 & ~n37207 ;
  assign n37209 = \m0_data_i[5]_pad  & n14271 ;
  assign n37210 = n14296 & n37209 ;
  assign n37211 = \m4_data_i[5]_pad  & n14271 ;
  assign n37212 = n14288 & n37211 ;
  assign n37213 = ~n37210 & ~n37212 ;
  assign n37214 = n37208 & n37213 ;
  assign n37215 = \m7_data_i[5]_pad  & ~n14271 ;
  assign n37216 = n14264 & n37215 ;
  assign n37217 = \m3_data_i[5]_pad  & ~n14271 ;
  assign n37218 = n14279 & n37217 ;
  assign n37219 = ~n37216 & ~n37218 ;
  assign n37220 = \m1_data_i[5]_pad  & ~n14271 ;
  assign n37221 = n14296 & n37220 ;
  assign n37222 = \m2_data_i[5]_pad  & n14271 ;
  assign n37223 = n14279 & n37222 ;
  assign n37224 = ~n37221 & ~n37223 ;
  assign n37225 = n37219 & n37224 ;
  assign n37226 = n37214 & n37225 ;
  assign n37227 = \m1_data_i[6]_pad  & ~n14271 ;
  assign n37228 = n14296 & n37227 ;
  assign n37229 = \m2_data_i[6]_pad  & n14271 ;
  assign n37230 = n14279 & n37229 ;
  assign n37231 = ~n37228 & ~n37230 ;
  assign n37232 = \m3_data_i[6]_pad  & ~n14271 ;
  assign n37233 = n14279 & n37232 ;
  assign n37234 = \m5_data_i[6]_pad  & ~n14271 ;
  assign n37235 = n14288 & n37234 ;
  assign n37236 = ~n37233 & ~n37235 ;
  assign n37237 = n37231 & n37236 ;
  assign n37238 = \m4_data_i[6]_pad  & n14271 ;
  assign n37239 = n14288 & n37238 ;
  assign n37240 = \m6_data_i[6]_pad  & n14271 ;
  assign n37241 = n14264 & n37240 ;
  assign n37242 = ~n37239 & ~n37241 ;
  assign n37243 = \m0_data_i[6]_pad  & n14271 ;
  assign n37244 = n14296 & n37243 ;
  assign n37245 = \m7_data_i[6]_pad  & ~n14271 ;
  assign n37246 = n14264 & n37245 ;
  assign n37247 = ~n37244 & ~n37246 ;
  assign n37248 = n37242 & n37247 ;
  assign n37249 = n37237 & n37248 ;
  assign n37250 = \m6_data_i[7]_pad  & n14271 ;
  assign n37251 = n14264 & n37250 ;
  assign n37252 = \m5_data_i[7]_pad  & ~n14271 ;
  assign n37253 = n14288 & n37252 ;
  assign n37254 = ~n37251 & ~n37253 ;
  assign n37255 = \m3_data_i[7]_pad  & ~n14271 ;
  assign n37256 = n14279 & n37255 ;
  assign n37257 = \m2_data_i[7]_pad  & n14271 ;
  assign n37258 = n14279 & n37257 ;
  assign n37259 = ~n37256 & ~n37258 ;
  assign n37260 = n37254 & n37259 ;
  assign n37261 = \m4_data_i[7]_pad  & n14271 ;
  assign n37262 = n14288 & n37261 ;
  assign n37263 = \m1_data_i[7]_pad  & ~n14271 ;
  assign n37264 = n14296 & n37263 ;
  assign n37265 = ~n37262 & ~n37264 ;
  assign n37266 = \m0_data_i[7]_pad  & n14271 ;
  assign n37267 = n14296 & n37266 ;
  assign n37268 = \m7_data_i[7]_pad  & ~n14271 ;
  assign n37269 = n14264 & n37268 ;
  assign n37270 = ~n37267 & ~n37269 ;
  assign n37271 = n37265 & n37270 ;
  assign n37272 = n37260 & n37271 ;
  assign n37273 = \m6_data_i[8]_pad  & n14271 ;
  assign n37274 = n14264 & n37273 ;
  assign n37275 = \m5_data_i[8]_pad  & ~n14271 ;
  assign n37276 = n14288 & n37275 ;
  assign n37277 = ~n37274 & ~n37276 ;
  assign n37278 = \m3_data_i[8]_pad  & ~n14271 ;
  assign n37279 = n14279 & n37278 ;
  assign n37280 = \m7_data_i[8]_pad  & ~n14271 ;
  assign n37281 = n14264 & n37280 ;
  assign n37282 = ~n37279 & ~n37281 ;
  assign n37283 = n37277 & n37282 ;
  assign n37284 = \m4_data_i[8]_pad  & n14271 ;
  assign n37285 = n14288 & n37284 ;
  assign n37286 = \m0_data_i[8]_pad  & n14271 ;
  assign n37287 = n14296 & n37286 ;
  assign n37288 = ~n37285 & ~n37287 ;
  assign n37289 = \m1_data_i[8]_pad  & ~n14271 ;
  assign n37290 = n14296 & n37289 ;
  assign n37291 = \m2_data_i[8]_pad  & n14271 ;
  assign n37292 = n14279 & n37291 ;
  assign n37293 = ~n37290 & ~n37292 ;
  assign n37294 = n37288 & n37293 ;
  assign n37295 = n37283 & n37294 ;
  assign n37296 = \m6_data_i[9]_pad  & n14271 ;
  assign n37297 = n14264 & n37296 ;
  assign n37298 = \m5_data_i[9]_pad  & ~n14271 ;
  assign n37299 = n14288 & n37298 ;
  assign n37300 = ~n37297 & ~n37299 ;
  assign n37301 = \m1_data_i[9]_pad  & ~n14271 ;
  assign n37302 = n14296 & n37301 ;
  assign n37303 = \m7_data_i[9]_pad  & ~n14271 ;
  assign n37304 = n14264 & n37303 ;
  assign n37305 = ~n37302 & ~n37304 ;
  assign n37306 = n37300 & n37305 ;
  assign n37307 = \m2_data_i[9]_pad  & n14271 ;
  assign n37308 = n14279 & n37307 ;
  assign n37309 = \m0_data_i[9]_pad  & n14271 ;
  assign n37310 = n14296 & n37309 ;
  assign n37311 = ~n37308 & ~n37310 ;
  assign n37312 = \m3_data_i[9]_pad  & ~n14271 ;
  assign n37313 = n14279 & n37312 ;
  assign n37314 = \m4_data_i[9]_pad  & n14271 ;
  assign n37315 = n14288 & n37314 ;
  assign n37316 = ~n37313 & ~n37315 ;
  assign n37317 = n37311 & n37316 ;
  assign n37318 = n37306 & n37317 ;
  assign n37319 = \m3_sel_i[0]_pad  & ~n14271 ;
  assign n37320 = n14279 & n37319 ;
  assign n37321 = \m4_sel_i[0]_pad  & n14271 ;
  assign n37322 = n14288 & n37321 ;
  assign n37323 = ~n37320 & ~n37322 ;
  assign n37324 = \m6_sel_i[0]_pad  & n14271 ;
  assign n37325 = n14264 & n37324 ;
  assign n37326 = \m2_sel_i[0]_pad  & n14271 ;
  assign n37327 = n14279 & n37326 ;
  assign n37328 = ~n37325 & ~n37327 ;
  assign n37329 = n37323 & n37328 ;
  assign n37330 = \m5_sel_i[0]_pad  & ~n14271 ;
  assign n37331 = n14288 & n37330 ;
  assign n37332 = \m1_sel_i[0]_pad  & ~n14271 ;
  assign n37333 = n14296 & n37332 ;
  assign n37334 = ~n37331 & ~n37333 ;
  assign n37335 = \m0_sel_i[0]_pad  & n14271 ;
  assign n37336 = n14296 & n37335 ;
  assign n37337 = \m7_sel_i[0]_pad  & ~n14271 ;
  assign n37338 = n14264 & n37337 ;
  assign n37339 = ~n37336 & ~n37338 ;
  assign n37340 = n37334 & n37339 ;
  assign n37341 = n37329 & n37340 ;
  assign n37342 = \m0_sel_i[1]_pad  & n14271 ;
  assign n37343 = n14296 & n37342 ;
  assign n37344 = \m7_sel_i[1]_pad  & ~n14271 ;
  assign n37345 = n14264 & n37344 ;
  assign n37346 = ~n37343 & ~n37345 ;
  assign n37347 = \m6_sel_i[1]_pad  & n14271 ;
  assign n37348 = n14264 & n37347 ;
  assign n37349 = \m2_sel_i[1]_pad  & n14271 ;
  assign n37350 = n14279 & n37349 ;
  assign n37351 = ~n37348 & ~n37350 ;
  assign n37352 = n37346 & n37351 ;
  assign n37353 = \m5_sel_i[1]_pad  & ~n14271 ;
  assign n37354 = n14288 & n37353 ;
  assign n37355 = \m1_sel_i[1]_pad  & ~n14271 ;
  assign n37356 = n14296 & n37355 ;
  assign n37357 = ~n37354 & ~n37356 ;
  assign n37358 = \m3_sel_i[1]_pad  & ~n14271 ;
  assign n37359 = n14279 & n37358 ;
  assign n37360 = \m4_sel_i[1]_pad  & n14271 ;
  assign n37361 = n14288 & n37360 ;
  assign n37362 = ~n37359 & ~n37361 ;
  assign n37363 = n37357 & n37362 ;
  assign n37364 = n37352 & n37363 ;
  assign n37365 = \m1_sel_i[2]_pad  & ~n14271 ;
  assign n37366 = n14296 & n37365 ;
  assign n37367 = \m2_sel_i[2]_pad  & n14271 ;
  assign n37368 = n14279 & n37367 ;
  assign n37369 = ~n37366 & ~n37368 ;
  assign n37370 = \m3_sel_i[2]_pad  & ~n14271 ;
  assign n37371 = n14279 & n37370 ;
  assign n37372 = \m7_sel_i[2]_pad  & ~n14271 ;
  assign n37373 = n14264 & n37372 ;
  assign n37374 = ~n37371 & ~n37373 ;
  assign n37375 = n37369 & n37374 ;
  assign n37376 = \m4_sel_i[2]_pad  & n14271 ;
  assign n37377 = n14288 & n37376 ;
  assign n37378 = \m0_sel_i[2]_pad  & n14271 ;
  assign n37379 = n14296 & n37378 ;
  assign n37380 = ~n37377 & ~n37379 ;
  assign n37381 = \m6_sel_i[2]_pad  & n14271 ;
  assign n37382 = n14264 & n37381 ;
  assign n37383 = \m5_sel_i[2]_pad  & ~n14271 ;
  assign n37384 = n14288 & n37383 ;
  assign n37385 = ~n37382 & ~n37384 ;
  assign n37386 = n37380 & n37385 ;
  assign n37387 = n37375 & n37386 ;
  assign n37388 = \m3_sel_i[3]_pad  & ~n14271 ;
  assign n37389 = n14279 & n37388 ;
  assign n37390 = \m4_sel_i[3]_pad  & n14271 ;
  assign n37391 = n14288 & n37390 ;
  assign n37392 = ~n37389 & ~n37391 ;
  assign n37393 = \m6_sel_i[3]_pad  & n14271 ;
  assign n37394 = n14264 & n37393 ;
  assign n37395 = \m2_sel_i[3]_pad  & n14271 ;
  assign n37396 = n14279 & n37395 ;
  assign n37397 = ~n37394 & ~n37396 ;
  assign n37398 = n37392 & n37397 ;
  assign n37399 = \m5_sel_i[3]_pad  & ~n14271 ;
  assign n37400 = n14288 & n37399 ;
  assign n37401 = \m1_sel_i[3]_pad  & ~n14271 ;
  assign n37402 = n14296 & n37401 ;
  assign n37403 = ~n37400 & ~n37402 ;
  assign n37404 = \m0_sel_i[3]_pad  & n14271 ;
  assign n37405 = n14296 & n37404 ;
  assign n37406 = \m7_sel_i[3]_pad  & ~n14271 ;
  assign n37407 = n14264 & n37406 ;
  assign n37408 = ~n37405 & ~n37407 ;
  assign n37409 = n37403 & n37408 ;
  assign n37410 = n37398 & n37409 ;
  assign n37411 = \m1_stb_i_pad  & n14658 ;
  assign n37412 = ~n14271 & n37411 ;
  assign n37413 = n14296 & n37412 ;
  assign n37414 = \m6_stb_i_pad  & n14640 ;
  assign n37415 = n14271 & n37414 ;
  assign n37416 = n14264 & n37415 ;
  assign n37417 = ~n37413 & ~n37416 ;
  assign n37418 = \m2_stb_i_pad  & n14596 ;
  assign n37419 = n14271 & n37418 ;
  assign n37420 = n14279 & n37419 ;
  assign n37421 = \m3_stb_i_pad  & n14609 ;
  assign n37422 = ~n14271 & n37421 ;
  assign n37423 = n14279 & n37422 ;
  assign n37424 = ~n37420 & ~n37423 ;
  assign n37425 = n37417 & n37424 ;
  assign n37426 = \m0_stb_i_pad  & n14575 ;
  assign n37427 = n14271 & n37426 ;
  assign n37428 = n14296 & n37427 ;
  assign n37429 = \m5_stb_i_pad  & n14561 ;
  assign n37430 = ~n14271 & n37429 ;
  assign n37431 = n14288 & n37430 ;
  assign n37432 = ~n37428 & ~n37431 ;
  assign n37433 = \m4_stb_i_pad  & n14622 ;
  assign n37434 = n14271 & n37433 ;
  assign n37435 = n14288 & n37434 ;
  assign n37436 = \m7_stb_i_pad  & n14653 ;
  assign n37437 = ~n14271 & n37436 ;
  assign n37438 = n14264 & n37437 ;
  assign n37439 = ~n37435 & ~n37438 ;
  assign n37440 = n37432 & n37439 ;
  assign n37441 = n37425 & n37440 ;
  assign n37442 = \m3_we_i_pad  & ~n14271 ;
  assign n37443 = n14279 & n37442 ;
  assign n37444 = \m4_we_i_pad  & n14271 ;
  assign n37445 = n14288 & n37444 ;
  assign n37446 = ~n37443 & ~n37445 ;
  assign n37447 = \m6_we_i_pad  & n14271 ;
  assign n37448 = n14264 & n37447 ;
  assign n37449 = \m2_we_i_pad  & n14271 ;
  assign n37450 = n14279 & n37449 ;
  assign n37451 = ~n37448 & ~n37450 ;
  assign n37452 = n37446 & n37451 ;
  assign n37453 = \m5_we_i_pad  & ~n14271 ;
  assign n37454 = n14288 & n37453 ;
  assign n37455 = \m1_we_i_pad  & ~n14271 ;
  assign n37456 = n14296 & n37455 ;
  assign n37457 = ~n37454 & ~n37456 ;
  assign n37458 = \m0_we_i_pad  & n14271 ;
  assign n37459 = n14296 & n37458 ;
  assign n37460 = \m7_we_i_pad  & ~n14271 ;
  assign n37461 = n14264 & n37460 ;
  assign n37462 = ~n37459 & ~n37461 ;
  assign n37463 = n37457 & n37462 ;
  assign n37464 = n37452 & n37463 ;
  assign n37465 = \m3_addr_i[0]_pad  & ~n14391 ;
  assign n37466 = n14416 & n37465 ;
  assign n37467 = \m4_addr_i[0]_pad  & n14391 ;
  assign n37468 = n14384 & n37467 ;
  assign n37469 = ~n37466 & ~n37468 ;
  assign n37470 = \m6_addr_i[0]_pad  & n14391 ;
  assign n37471 = n14408 & n37470 ;
  assign n37472 = \m2_addr_i[0]_pad  & n14391 ;
  assign n37473 = n14416 & n37472 ;
  assign n37474 = ~n37471 & ~n37473 ;
  assign n37475 = n37469 & n37474 ;
  assign n37476 = \m5_addr_i[0]_pad  & ~n14391 ;
  assign n37477 = n14384 & n37476 ;
  assign n37478 = \m1_addr_i[0]_pad  & ~n14391 ;
  assign n37479 = n14399 & n37478 ;
  assign n37480 = ~n37477 & ~n37479 ;
  assign n37481 = \m0_addr_i[0]_pad  & n14391 ;
  assign n37482 = n14399 & n37481 ;
  assign n37483 = \m7_addr_i[0]_pad  & ~n14391 ;
  assign n37484 = n14408 & n37483 ;
  assign n37485 = ~n37482 & ~n37484 ;
  assign n37486 = n37480 & n37485 ;
  assign n37487 = n37475 & n37486 ;
  assign n37488 = \m3_addr_i[10]_pad  & ~n14391 ;
  assign n37489 = n14416 & n37488 ;
  assign n37490 = \m4_addr_i[10]_pad  & n14391 ;
  assign n37491 = n14384 & n37490 ;
  assign n37492 = ~n37489 & ~n37491 ;
  assign n37493 = \m6_addr_i[10]_pad  & n14391 ;
  assign n37494 = n14408 & n37493 ;
  assign n37495 = \m2_addr_i[10]_pad  & n14391 ;
  assign n37496 = n14416 & n37495 ;
  assign n37497 = ~n37494 & ~n37496 ;
  assign n37498 = n37492 & n37497 ;
  assign n37499 = \m5_addr_i[10]_pad  & ~n14391 ;
  assign n37500 = n14384 & n37499 ;
  assign n37501 = \m1_addr_i[10]_pad  & ~n14391 ;
  assign n37502 = n14399 & n37501 ;
  assign n37503 = ~n37500 & ~n37502 ;
  assign n37504 = \m0_addr_i[10]_pad  & n14391 ;
  assign n37505 = n14399 & n37504 ;
  assign n37506 = \m7_addr_i[10]_pad  & ~n14391 ;
  assign n37507 = n14408 & n37506 ;
  assign n37508 = ~n37505 & ~n37507 ;
  assign n37509 = n37503 & n37508 ;
  assign n37510 = n37498 & n37509 ;
  assign n37511 = \m3_addr_i[11]_pad  & ~n14391 ;
  assign n37512 = n14416 & n37511 ;
  assign n37513 = \m4_addr_i[11]_pad  & n14391 ;
  assign n37514 = n14384 & n37513 ;
  assign n37515 = ~n37512 & ~n37514 ;
  assign n37516 = \m6_addr_i[11]_pad  & n14391 ;
  assign n37517 = n14408 & n37516 ;
  assign n37518 = \m2_addr_i[11]_pad  & n14391 ;
  assign n37519 = n14416 & n37518 ;
  assign n37520 = ~n37517 & ~n37519 ;
  assign n37521 = n37515 & n37520 ;
  assign n37522 = \m5_addr_i[11]_pad  & ~n14391 ;
  assign n37523 = n14384 & n37522 ;
  assign n37524 = \m1_addr_i[11]_pad  & ~n14391 ;
  assign n37525 = n14399 & n37524 ;
  assign n37526 = ~n37523 & ~n37525 ;
  assign n37527 = \m0_addr_i[11]_pad  & n14391 ;
  assign n37528 = n14399 & n37527 ;
  assign n37529 = \m7_addr_i[11]_pad  & ~n14391 ;
  assign n37530 = n14408 & n37529 ;
  assign n37531 = ~n37528 & ~n37530 ;
  assign n37532 = n37526 & n37531 ;
  assign n37533 = n37521 & n37532 ;
  assign n37534 = \m3_addr_i[12]_pad  & ~n14391 ;
  assign n37535 = n14416 & n37534 ;
  assign n37536 = \m4_addr_i[12]_pad  & n14391 ;
  assign n37537 = n14384 & n37536 ;
  assign n37538 = ~n37535 & ~n37537 ;
  assign n37539 = \m6_addr_i[12]_pad  & n14391 ;
  assign n37540 = n14408 & n37539 ;
  assign n37541 = \m2_addr_i[12]_pad  & n14391 ;
  assign n37542 = n14416 & n37541 ;
  assign n37543 = ~n37540 & ~n37542 ;
  assign n37544 = n37538 & n37543 ;
  assign n37545 = \m5_addr_i[12]_pad  & ~n14391 ;
  assign n37546 = n14384 & n37545 ;
  assign n37547 = \m1_addr_i[12]_pad  & ~n14391 ;
  assign n37548 = n14399 & n37547 ;
  assign n37549 = ~n37546 & ~n37548 ;
  assign n37550 = \m0_addr_i[12]_pad  & n14391 ;
  assign n37551 = n14399 & n37550 ;
  assign n37552 = \m7_addr_i[12]_pad  & ~n14391 ;
  assign n37553 = n14408 & n37552 ;
  assign n37554 = ~n37551 & ~n37553 ;
  assign n37555 = n37549 & n37554 ;
  assign n37556 = n37544 & n37555 ;
  assign n37557 = \m3_addr_i[13]_pad  & ~n14391 ;
  assign n37558 = n14416 & n37557 ;
  assign n37559 = \m4_addr_i[13]_pad  & n14391 ;
  assign n37560 = n14384 & n37559 ;
  assign n37561 = ~n37558 & ~n37560 ;
  assign n37562 = \m6_addr_i[13]_pad  & n14391 ;
  assign n37563 = n14408 & n37562 ;
  assign n37564 = \m2_addr_i[13]_pad  & n14391 ;
  assign n37565 = n14416 & n37564 ;
  assign n37566 = ~n37563 & ~n37565 ;
  assign n37567 = n37561 & n37566 ;
  assign n37568 = \m5_addr_i[13]_pad  & ~n14391 ;
  assign n37569 = n14384 & n37568 ;
  assign n37570 = \m1_addr_i[13]_pad  & ~n14391 ;
  assign n37571 = n14399 & n37570 ;
  assign n37572 = ~n37569 & ~n37571 ;
  assign n37573 = \m0_addr_i[13]_pad  & n14391 ;
  assign n37574 = n14399 & n37573 ;
  assign n37575 = \m7_addr_i[13]_pad  & ~n14391 ;
  assign n37576 = n14408 & n37575 ;
  assign n37577 = ~n37574 & ~n37576 ;
  assign n37578 = n37572 & n37577 ;
  assign n37579 = n37567 & n37578 ;
  assign n37580 = \m3_addr_i[14]_pad  & ~n14391 ;
  assign n37581 = n14416 & n37580 ;
  assign n37582 = \m4_addr_i[14]_pad  & n14391 ;
  assign n37583 = n14384 & n37582 ;
  assign n37584 = ~n37581 & ~n37583 ;
  assign n37585 = \m6_addr_i[14]_pad  & n14391 ;
  assign n37586 = n14408 & n37585 ;
  assign n37587 = \m2_addr_i[14]_pad  & n14391 ;
  assign n37588 = n14416 & n37587 ;
  assign n37589 = ~n37586 & ~n37588 ;
  assign n37590 = n37584 & n37589 ;
  assign n37591 = \m5_addr_i[14]_pad  & ~n14391 ;
  assign n37592 = n14384 & n37591 ;
  assign n37593 = \m1_addr_i[14]_pad  & ~n14391 ;
  assign n37594 = n14399 & n37593 ;
  assign n37595 = ~n37592 & ~n37594 ;
  assign n37596 = \m0_addr_i[14]_pad  & n14391 ;
  assign n37597 = n14399 & n37596 ;
  assign n37598 = \m7_addr_i[14]_pad  & ~n14391 ;
  assign n37599 = n14408 & n37598 ;
  assign n37600 = ~n37597 & ~n37599 ;
  assign n37601 = n37595 & n37600 ;
  assign n37602 = n37590 & n37601 ;
  assign n37603 = \m3_addr_i[15]_pad  & ~n14391 ;
  assign n37604 = n14416 & n37603 ;
  assign n37605 = \m4_addr_i[15]_pad  & n14391 ;
  assign n37606 = n14384 & n37605 ;
  assign n37607 = ~n37604 & ~n37606 ;
  assign n37608 = \m6_addr_i[15]_pad  & n14391 ;
  assign n37609 = n14408 & n37608 ;
  assign n37610 = \m2_addr_i[15]_pad  & n14391 ;
  assign n37611 = n14416 & n37610 ;
  assign n37612 = ~n37609 & ~n37611 ;
  assign n37613 = n37607 & n37612 ;
  assign n37614 = \m5_addr_i[15]_pad  & ~n14391 ;
  assign n37615 = n14384 & n37614 ;
  assign n37616 = \m1_addr_i[15]_pad  & ~n14391 ;
  assign n37617 = n14399 & n37616 ;
  assign n37618 = ~n37615 & ~n37617 ;
  assign n37619 = \m0_addr_i[15]_pad  & n14391 ;
  assign n37620 = n14399 & n37619 ;
  assign n37621 = \m7_addr_i[15]_pad  & ~n14391 ;
  assign n37622 = n14408 & n37621 ;
  assign n37623 = ~n37620 & ~n37622 ;
  assign n37624 = n37618 & n37623 ;
  assign n37625 = n37613 & n37624 ;
  assign n37626 = \m3_addr_i[16]_pad  & ~n14391 ;
  assign n37627 = n14416 & n37626 ;
  assign n37628 = \m4_addr_i[16]_pad  & n14391 ;
  assign n37629 = n14384 & n37628 ;
  assign n37630 = ~n37627 & ~n37629 ;
  assign n37631 = \m6_addr_i[16]_pad  & n14391 ;
  assign n37632 = n14408 & n37631 ;
  assign n37633 = \m2_addr_i[16]_pad  & n14391 ;
  assign n37634 = n14416 & n37633 ;
  assign n37635 = ~n37632 & ~n37634 ;
  assign n37636 = n37630 & n37635 ;
  assign n37637 = \m5_addr_i[16]_pad  & ~n14391 ;
  assign n37638 = n14384 & n37637 ;
  assign n37639 = \m1_addr_i[16]_pad  & ~n14391 ;
  assign n37640 = n14399 & n37639 ;
  assign n37641 = ~n37638 & ~n37640 ;
  assign n37642 = \m0_addr_i[16]_pad  & n14391 ;
  assign n37643 = n14399 & n37642 ;
  assign n37644 = \m7_addr_i[16]_pad  & ~n14391 ;
  assign n37645 = n14408 & n37644 ;
  assign n37646 = ~n37643 & ~n37645 ;
  assign n37647 = n37641 & n37646 ;
  assign n37648 = n37636 & n37647 ;
  assign n37649 = \m3_addr_i[17]_pad  & ~n14391 ;
  assign n37650 = n14416 & n37649 ;
  assign n37651 = \m4_addr_i[17]_pad  & n14391 ;
  assign n37652 = n14384 & n37651 ;
  assign n37653 = ~n37650 & ~n37652 ;
  assign n37654 = \m6_addr_i[17]_pad  & n14391 ;
  assign n37655 = n14408 & n37654 ;
  assign n37656 = \m2_addr_i[17]_pad  & n14391 ;
  assign n37657 = n14416 & n37656 ;
  assign n37658 = ~n37655 & ~n37657 ;
  assign n37659 = n37653 & n37658 ;
  assign n37660 = \m5_addr_i[17]_pad  & ~n14391 ;
  assign n37661 = n14384 & n37660 ;
  assign n37662 = \m1_addr_i[17]_pad  & ~n14391 ;
  assign n37663 = n14399 & n37662 ;
  assign n37664 = ~n37661 & ~n37663 ;
  assign n37665 = \m0_addr_i[17]_pad  & n14391 ;
  assign n37666 = n14399 & n37665 ;
  assign n37667 = \m7_addr_i[17]_pad  & ~n14391 ;
  assign n37668 = n14408 & n37667 ;
  assign n37669 = ~n37666 & ~n37668 ;
  assign n37670 = n37664 & n37669 ;
  assign n37671 = n37659 & n37670 ;
  assign n37672 = \m3_addr_i[18]_pad  & ~n14391 ;
  assign n37673 = n14416 & n37672 ;
  assign n37674 = \m4_addr_i[18]_pad  & n14391 ;
  assign n37675 = n14384 & n37674 ;
  assign n37676 = ~n37673 & ~n37675 ;
  assign n37677 = \m6_addr_i[18]_pad  & n14391 ;
  assign n37678 = n14408 & n37677 ;
  assign n37679 = \m2_addr_i[18]_pad  & n14391 ;
  assign n37680 = n14416 & n37679 ;
  assign n37681 = ~n37678 & ~n37680 ;
  assign n37682 = n37676 & n37681 ;
  assign n37683 = \m5_addr_i[18]_pad  & ~n14391 ;
  assign n37684 = n14384 & n37683 ;
  assign n37685 = \m1_addr_i[18]_pad  & ~n14391 ;
  assign n37686 = n14399 & n37685 ;
  assign n37687 = ~n37684 & ~n37686 ;
  assign n37688 = \m0_addr_i[18]_pad  & n14391 ;
  assign n37689 = n14399 & n37688 ;
  assign n37690 = \m7_addr_i[18]_pad  & ~n14391 ;
  assign n37691 = n14408 & n37690 ;
  assign n37692 = ~n37689 & ~n37691 ;
  assign n37693 = n37687 & n37692 ;
  assign n37694 = n37682 & n37693 ;
  assign n37695 = \m3_addr_i[19]_pad  & ~n14391 ;
  assign n37696 = n14416 & n37695 ;
  assign n37697 = \m4_addr_i[19]_pad  & n14391 ;
  assign n37698 = n14384 & n37697 ;
  assign n37699 = ~n37696 & ~n37698 ;
  assign n37700 = \m6_addr_i[19]_pad  & n14391 ;
  assign n37701 = n14408 & n37700 ;
  assign n37702 = \m2_addr_i[19]_pad  & n14391 ;
  assign n37703 = n14416 & n37702 ;
  assign n37704 = ~n37701 & ~n37703 ;
  assign n37705 = n37699 & n37704 ;
  assign n37706 = \m5_addr_i[19]_pad  & ~n14391 ;
  assign n37707 = n14384 & n37706 ;
  assign n37708 = \m1_addr_i[19]_pad  & ~n14391 ;
  assign n37709 = n14399 & n37708 ;
  assign n37710 = ~n37707 & ~n37709 ;
  assign n37711 = \m0_addr_i[19]_pad  & n14391 ;
  assign n37712 = n14399 & n37711 ;
  assign n37713 = \m7_addr_i[19]_pad  & ~n14391 ;
  assign n37714 = n14408 & n37713 ;
  assign n37715 = ~n37712 & ~n37714 ;
  assign n37716 = n37710 & n37715 ;
  assign n37717 = n37705 & n37716 ;
  assign n37718 = \m3_addr_i[1]_pad  & ~n14391 ;
  assign n37719 = n14416 & n37718 ;
  assign n37720 = \m4_addr_i[1]_pad  & n14391 ;
  assign n37721 = n14384 & n37720 ;
  assign n37722 = ~n37719 & ~n37721 ;
  assign n37723 = \m6_addr_i[1]_pad  & n14391 ;
  assign n37724 = n14408 & n37723 ;
  assign n37725 = \m2_addr_i[1]_pad  & n14391 ;
  assign n37726 = n14416 & n37725 ;
  assign n37727 = ~n37724 & ~n37726 ;
  assign n37728 = n37722 & n37727 ;
  assign n37729 = \m5_addr_i[1]_pad  & ~n14391 ;
  assign n37730 = n14384 & n37729 ;
  assign n37731 = \m1_addr_i[1]_pad  & ~n14391 ;
  assign n37732 = n14399 & n37731 ;
  assign n37733 = ~n37730 & ~n37732 ;
  assign n37734 = \m0_addr_i[1]_pad  & n14391 ;
  assign n37735 = n14399 & n37734 ;
  assign n37736 = \m7_addr_i[1]_pad  & ~n14391 ;
  assign n37737 = n14408 & n37736 ;
  assign n37738 = ~n37735 & ~n37737 ;
  assign n37739 = n37733 & n37738 ;
  assign n37740 = n37728 & n37739 ;
  assign n37741 = \m3_addr_i[20]_pad  & ~n14391 ;
  assign n37742 = n14416 & n37741 ;
  assign n37743 = \m4_addr_i[20]_pad  & n14391 ;
  assign n37744 = n14384 & n37743 ;
  assign n37745 = ~n37742 & ~n37744 ;
  assign n37746 = \m6_addr_i[20]_pad  & n14391 ;
  assign n37747 = n14408 & n37746 ;
  assign n37748 = \m2_addr_i[20]_pad  & n14391 ;
  assign n37749 = n14416 & n37748 ;
  assign n37750 = ~n37747 & ~n37749 ;
  assign n37751 = n37745 & n37750 ;
  assign n37752 = \m5_addr_i[20]_pad  & ~n14391 ;
  assign n37753 = n14384 & n37752 ;
  assign n37754 = \m1_addr_i[20]_pad  & ~n14391 ;
  assign n37755 = n14399 & n37754 ;
  assign n37756 = ~n37753 & ~n37755 ;
  assign n37757 = \m0_addr_i[20]_pad  & n14391 ;
  assign n37758 = n14399 & n37757 ;
  assign n37759 = \m7_addr_i[20]_pad  & ~n14391 ;
  assign n37760 = n14408 & n37759 ;
  assign n37761 = ~n37758 & ~n37760 ;
  assign n37762 = n37756 & n37761 ;
  assign n37763 = n37751 & n37762 ;
  assign n37764 = \m3_addr_i[21]_pad  & ~n14391 ;
  assign n37765 = n14416 & n37764 ;
  assign n37766 = \m4_addr_i[21]_pad  & n14391 ;
  assign n37767 = n14384 & n37766 ;
  assign n37768 = ~n37765 & ~n37767 ;
  assign n37769 = \m6_addr_i[21]_pad  & n14391 ;
  assign n37770 = n14408 & n37769 ;
  assign n37771 = \m2_addr_i[21]_pad  & n14391 ;
  assign n37772 = n14416 & n37771 ;
  assign n37773 = ~n37770 & ~n37772 ;
  assign n37774 = n37768 & n37773 ;
  assign n37775 = \m5_addr_i[21]_pad  & ~n14391 ;
  assign n37776 = n14384 & n37775 ;
  assign n37777 = \m1_addr_i[21]_pad  & ~n14391 ;
  assign n37778 = n14399 & n37777 ;
  assign n37779 = ~n37776 & ~n37778 ;
  assign n37780 = \m0_addr_i[21]_pad  & n14391 ;
  assign n37781 = n14399 & n37780 ;
  assign n37782 = \m7_addr_i[21]_pad  & ~n14391 ;
  assign n37783 = n14408 & n37782 ;
  assign n37784 = ~n37781 & ~n37783 ;
  assign n37785 = n37779 & n37784 ;
  assign n37786 = n37774 & n37785 ;
  assign n37787 = \m3_addr_i[22]_pad  & ~n14391 ;
  assign n37788 = n14416 & n37787 ;
  assign n37789 = \m4_addr_i[22]_pad  & n14391 ;
  assign n37790 = n14384 & n37789 ;
  assign n37791 = ~n37788 & ~n37790 ;
  assign n37792 = \m6_addr_i[22]_pad  & n14391 ;
  assign n37793 = n14408 & n37792 ;
  assign n37794 = \m2_addr_i[22]_pad  & n14391 ;
  assign n37795 = n14416 & n37794 ;
  assign n37796 = ~n37793 & ~n37795 ;
  assign n37797 = n37791 & n37796 ;
  assign n37798 = \m5_addr_i[22]_pad  & ~n14391 ;
  assign n37799 = n14384 & n37798 ;
  assign n37800 = \m1_addr_i[22]_pad  & ~n14391 ;
  assign n37801 = n14399 & n37800 ;
  assign n37802 = ~n37799 & ~n37801 ;
  assign n37803 = \m0_addr_i[22]_pad  & n14391 ;
  assign n37804 = n14399 & n37803 ;
  assign n37805 = \m7_addr_i[22]_pad  & ~n14391 ;
  assign n37806 = n14408 & n37805 ;
  assign n37807 = ~n37804 & ~n37806 ;
  assign n37808 = n37802 & n37807 ;
  assign n37809 = n37797 & n37808 ;
  assign n37810 = \m3_addr_i[23]_pad  & ~n14391 ;
  assign n37811 = n14416 & n37810 ;
  assign n37812 = \m4_addr_i[23]_pad  & n14391 ;
  assign n37813 = n14384 & n37812 ;
  assign n37814 = ~n37811 & ~n37813 ;
  assign n37815 = \m6_addr_i[23]_pad  & n14391 ;
  assign n37816 = n14408 & n37815 ;
  assign n37817 = \m2_addr_i[23]_pad  & n14391 ;
  assign n37818 = n14416 & n37817 ;
  assign n37819 = ~n37816 & ~n37818 ;
  assign n37820 = n37814 & n37819 ;
  assign n37821 = \m5_addr_i[23]_pad  & ~n14391 ;
  assign n37822 = n14384 & n37821 ;
  assign n37823 = \m1_addr_i[23]_pad  & ~n14391 ;
  assign n37824 = n14399 & n37823 ;
  assign n37825 = ~n37822 & ~n37824 ;
  assign n37826 = \m0_addr_i[23]_pad  & n14391 ;
  assign n37827 = n14399 & n37826 ;
  assign n37828 = \m7_addr_i[23]_pad  & ~n14391 ;
  assign n37829 = n14408 & n37828 ;
  assign n37830 = ~n37827 & ~n37829 ;
  assign n37831 = n37825 & n37830 ;
  assign n37832 = n37820 & n37831 ;
  assign n37833 = \m3_addr_i[24]_pad  & ~n14391 ;
  assign n37834 = n14416 & n37833 ;
  assign n37835 = \m4_addr_i[24]_pad  & n14391 ;
  assign n37836 = n14384 & n37835 ;
  assign n37837 = ~n37834 & ~n37836 ;
  assign n37838 = \m5_addr_i[24]_pad  & ~n14391 ;
  assign n37839 = n14384 & n37838 ;
  assign n37840 = \m2_addr_i[24]_pad  & n14391 ;
  assign n37841 = n14416 & n37840 ;
  assign n37842 = ~n37839 & ~n37841 ;
  assign n37843 = n37837 & n37842 ;
  assign n37844 = \m6_addr_i[24]_pad  & n14391 ;
  assign n37845 = n14408 & n37844 ;
  assign n37846 = \m1_addr_i[24]_pad  & ~n14391 ;
  assign n37847 = n14399 & n37846 ;
  assign n37848 = ~n37845 & ~n37847 ;
  assign n37849 = \m0_addr_i[24]_pad  & n14391 ;
  assign n37850 = n14399 & n37849 ;
  assign n37851 = \m7_addr_i[24]_pad  & ~n14391 ;
  assign n37852 = n14408 & n37851 ;
  assign n37853 = ~n37850 & ~n37852 ;
  assign n37854 = n37848 & n37853 ;
  assign n37855 = n37843 & n37854 ;
  assign n37856 = \m3_addr_i[25]_pad  & ~n14391 ;
  assign n37857 = n14416 & n37856 ;
  assign n37858 = \m4_addr_i[25]_pad  & n14391 ;
  assign n37859 = n14384 & n37858 ;
  assign n37860 = ~n37857 & ~n37859 ;
  assign n37861 = \m5_addr_i[25]_pad  & ~n14391 ;
  assign n37862 = n14384 & n37861 ;
  assign n37863 = \m2_addr_i[25]_pad  & n14391 ;
  assign n37864 = n14416 & n37863 ;
  assign n37865 = ~n37862 & ~n37864 ;
  assign n37866 = n37860 & n37865 ;
  assign n37867 = \m6_addr_i[25]_pad  & n14391 ;
  assign n37868 = n14408 & n37867 ;
  assign n37869 = \m1_addr_i[25]_pad  & ~n14391 ;
  assign n37870 = n14399 & n37869 ;
  assign n37871 = ~n37868 & ~n37870 ;
  assign n37872 = \m0_addr_i[25]_pad  & n14391 ;
  assign n37873 = n14399 & n37872 ;
  assign n37874 = \m7_addr_i[25]_pad  & ~n14391 ;
  assign n37875 = n14408 & n37874 ;
  assign n37876 = ~n37873 & ~n37875 ;
  assign n37877 = n37871 & n37876 ;
  assign n37878 = n37866 & n37877 ;
  assign n37879 = \m3_addr_i[26]_pad  & ~n14391 ;
  assign n37880 = n14416 & n37879 ;
  assign n37881 = \m4_addr_i[26]_pad  & n14391 ;
  assign n37882 = n14384 & n37881 ;
  assign n37883 = ~n37880 & ~n37882 ;
  assign n37884 = \m5_addr_i[26]_pad  & ~n14391 ;
  assign n37885 = n14384 & n37884 ;
  assign n37886 = \m2_addr_i[26]_pad  & n14391 ;
  assign n37887 = n14416 & n37886 ;
  assign n37888 = ~n37885 & ~n37887 ;
  assign n37889 = n37883 & n37888 ;
  assign n37890 = \m6_addr_i[26]_pad  & n14391 ;
  assign n37891 = n14408 & n37890 ;
  assign n37892 = \m1_addr_i[26]_pad  & ~n14391 ;
  assign n37893 = n14399 & n37892 ;
  assign n37894 = ~n37891 & ~n37893 ;
  assign n37895 = \m0_addr_i[26]_pad  & n14391 ;
  assign n37896 = n14399 & n37895 ;
  assign n37897 = \m7_addr_i[26]_pad  & ~n14391 ;
  assign n37898 = n14408 & n37897 ;
  assign n37899 = ~n37896 & ~n37898 ;
  assign n37900 = n37894 & n37899 ;
  assign n37901 = n37889 & n37900 ;
  assign n37902 = \m3_addr_i[27]_pad  & ~n14391 ;
  assign n37903 = n14416 & n37902 ;
  assign n37904 = \m4_addr_i[27]_pad  & n14391 ;
  assign n37905 = n14384 & n37904 ;
  assign n37906 = ~n37903 & ~n37905 ;
  assign n37907 = \m5_addr_i[27]_pad  & ~n14391 ;
  assign n37908 = n14384 & n37907 ;
  assign n37909 = \m2_addr_i[27]_pad  & n14391 ;
  assign n37910 = n14416 & n37909 ;
  assign n37911 = ~n37908 & ~n37910 ;
  assign n37912 = n37906 & n37911 ;
  assign n37913 = \m6_addr_i[27]_pad  & n14391 ;
  assign n37914 = n14408 & n37913 ;
  assign n37915 = \m1_addr_i[27]_pad  & ~n14391 ;
  assign n37916 = n14399 & n37915 ;
  assign n37917 = ~n37914 & ~n37916 ;
  assign n37918 = \m0_addr_i[27]_pad  & n14391 ;
  assign n37919 = n14399 & n37918 ;
  assign n37920 = \m7_addr_i[27]_pad  & ~n14391 ;
  assign n37921 = n14408 & n37920 ;
  assign n37922 = ~n37919 & ~n37921 ;
  assign n37923 = n37917 & n37922 ;
  assign n37924 = n37912 & n37923 ;
  assign n37925 = \m3_addr_i[28]_pad  & ~n14391 ;
  assign n37926 = n14416 & n37925 ;
  assign n37927 = \m4_addr_i[28]_pad  & n14391 ;
  assign n37928 = n14384 & n37927 ;
  assign n37929 = ~n37926 & ~n37928 ;
  assign n37930 = \m5_addr_i[28]_pad  & ~n14391 ;
  assign n37931 = n14384 & n37930 ;
  assign n37932 = \m2_addr_i[28]_pad  & n14391 ;
  assign n37933 = n14416 & n37932 ;
  assign n37934 = ~n37931 & ~n37933 ;
  assign n37935 = n37929 & n37934 ;
  assign n37936 = \m6_addr_i[28]_pad  & n14391 ;
  assign n37937 = n14408 & n37936 ;
  assign n37938 = \m1_addr_i[28]_pad  & ~n14391 ;
  assign n37939 = n14399 & n37938 ;
  assign n37940 = ~n37937 & ~n37939 ;
  assign n37941 = \m0_addr_i[28]_pad  & n14391 ;
  assign n37942 = n14399 & n37941 ;
  assign n37943 = \m7_addr_i[28]_pad  & ~n14391 ;
  assign n37944 = n14408 & n37943 ;
  assign n37945 = ~n37942 & ~n37944 ;
  assign n37946 = n37940 & n37945 ;
  assign n37947 = n37935 & n37946 ;
  assign n37948 = \m3_addr_i[29]_pad  & ~n14391 ;
  assign n37949 = n14416 & n37948 ;
  assign n37950 = \m4_addr_i[29]_pad  & n14391 ;
  assign n37951 = n14384 & n37950 ;
  assign n37952 = ~n37949 & ~n37951 ;
  assign n37953 = \m5_addr_i[29]_pad  & ~n14391 ;
  assign n37954 = n14384 & n37953 ;
  assign n37955 = \m2_addr_i[29]_pad  & n14391 ;
  assign n37956 = n14416 & n37955 ;
  assign n37957 = ~n37954 & ~n37956 ;
  assign n37958 = n37952 & n37957 ;
  assign n37959 = \m6_addr_i[29]_pad  & n14391 ;
  assign n37960 = n14408 & n37959 ;
  assign n37961 = \m1_addr_i[29]_pad  & ~n14391 ;
  assign n37962 = n14399 & n37961 ;
  assign n37963 = ~n37960 & ~n37962 ;
  assign n37964 = \m0_addr_i[29]_pad  & n14391 ;
  assign n37965 = n14399 & n37964 ;
  assign n37966 = \m7_addr_i[29]_pad  & ~n14391 ;
  assign n37967 = n14408 & n37966 ;
  assign n37968 = ~n37965 & ~n37967 ;
  assign n37969 = n37963 & n37968 ;
  assign n37970 = n37958 & n37969 ;
  assign n37971 = \m3_addr_i[2]_pad  & ~n14391 ;
  assign n37972 = n14416 & n37971 ;
  assign n37973 = \m4_addr_i[2]_pad  & n14391 ;
  assign n37974 = n14384 & n37973 ;
  assign n37975 = ~n37972 & ~n37974 ;
  assign n37976 = \m6_addr_i[2]_pad  & n14391 ;
  assign n37977 = n14408 & n37976 ;
  assign n37978 = \m2_addr_i[2]_pad  & n14391 ;
  assign n37979 = n14416 & n37978 ;
  assign n37980 = ~n37977 & ~n37979 ;
  assign n37981 = n37975 & n37980 ;
  assign n37982 = \m5_addr_i[2]_pad  & ~n14391 ;
  assign n37983 = n14384 & n37982 ;
  assign n37984 = \m1_addr_i[2]_pad  & ~n14391 ;
  assign n37985 = n14399 & n37984 ;
  assign n37986 = ~n37983 & ~n37985 ;
  assign n37987 = \m0_addr_i[2]_pad  & n14391 ;
  assign n37988 = n14399 & n37987 ;
  assign n37989 = \m7_addr_i[2]_pad  & ~n14391 ;
  assign n37990 = n14408 & n37989 ;
  assign n37991 = ~n37988 & ~n37990 ;
  assign n37992 = n37986 & n37991 ;
  assign n37993 = n37981 & n37992 ;
  assign n37994 = \m3_addr_i[30]_pad  & ~n14391 ;
  assign n37995 = n14416 & n37994 ;
  assign n37996 = \m4_addr_i[30]_pad  & n14391 ;
  assign n37997 = n14384 & n37996 ;
  assign n37998 = ~n37995 & ~n37997 ;
  assign n37999 = \m5_addr_i[30]_pad  & ~n14391 ;
  assign n38000 = n14384 & n37999 ;
  assign n38001 = \m2_addr_i[30]_pad  & n14391 ;
  assign n38002 = n14416 & n38001 ;
  assign n38003 = ~n38000 & ~n38002 ;
  assign n38004 = n37998 & n38003 ;
  assign n38005 = \m6_addr_i[30]_pad  & n14391 ;
  assign n38006 = n14408 & n38005 ;
  assign n38007 = \m1_addr_i[30]_pad  & ~n14391 ;
  assign n38008 = n14399 & n38007 ;
  assign n38009 = ~n38006 & ~n38008 ;
  assign n38010 = \m0_addr_i[30]_pad  & n14391 ;
  assign n38011 = n14399 & n38010 ;
  assign n38012 = \m7_addr_i[30]_pad  & ~n14391 ;
  assign n38013 = n14408 & n38012 ;
  assign n38014 = ~n38011 & ~n38013 ;
  assign n38015 = n38009 & n38014 ;
  assign n38016 = n38004 & n38015 ;
  assign n38017 = \m3_addr_i[31]_pad  & ~n14391 ;
  assign n38018 = n14416 & n38017 ;
  assign n38019 = \m4_addr_i[31]_pad  & n14391 ;
  assign n38020 = n14384 & n38019 ;
  assign n38021 = ~n38018 & ~n38020 ;
  assign n38022 = \m5_addr_i[31]_pad  & ~n14391 ;
  assign n38023 = n14384 & n38022 ;
  assign n38024 = \m2_addr_i[31]_pad  & n14391 ;
  assign n38025 = n14416 & n38024 ;
  assign n38026 = ~n38023 & ~n38025 ;
  assign n38027 = n38021 & n38026 ;
  assign n38028 = \m6_addr_i[31]_pad  & n14391 ;
  assign n38029 = n14408 & n38028 ;
  assign n38030 = \m1_addr_i[31]_pad  & ~n14391 ;
  assign n38031 = n14399 & n38030 ;
  assign n38032 = ~n38029 & ~n38031 ;
  assign n38033 = \m0_addr_i[31]_pad  & n14391 ;
  assign n38034 = n14399 & n38033 ;
  assign n38035 = \m7_addr_i[31]_pad  & ~n14391 ;
  assign n38036 = n14408 & n38035 ;
  assign n38037 = ~n38034 & ~n38036 ;
  assign n38038 = n38032 & n38037 ;
  assign n38039 = n38027 & n38038 ;
  assign n38040 = \m3_addr_i[3]_pad  & ~n14391 ;
  assign n38041 = n14416 & n38040 ;
  assign n38042 = \m4_addr_i[3]_pad  & n14391 ;
  assign n38043 = n14384 & n38042 ;
  assign n38044 = ~n38041 & ~n38043 ;
  assign n38045 = \m6_addr_i[3]_pad  & n14391 ;
  assign n38046 = n14408 & n38045 ;
  assign n38047 = \m2_addr_i[3]_pad  & n14391 ;
  assign n38048 = n14416 & n38047 ;
  assign n38049 = ~n38046 & ~n38048 ;
  assign n38050 = n38044 & n38049 ;
  assign n38051 = \m5_addr_i[3]_pad  & ~n14391 ;
  assign n38052 = n14384 & n38051 ;
  assign n38053 = \m1_addr_i[3]_pad  & ~n14391 ;
  assign n38054 = n14399 & n38053 ;
  assign n38055 = ~n38052 & ~n38054 ;
  assign n38056 = \m0_addr_i[3]_pad  & n14391 ;
  assign n38057 = n14399 & n38056 ;
  assign n38058 = \m7_addr_i[3]_pad  & ~n14391 ;
  assign n38059 = n14408 & n38058 ;
  assign n38060 = ~n38057 & ~n38059 ;
  assign n38061 = n38055 & n38060 ;
  assign n38062 = n38050 & n38061 ;
  assign n38063 = \m3_addr_i[4]_pad  & ~n14391 ;
  assign n38064 = n14416 & n38063 ;
  assign n38065 = \m4_addr_i[4]_pad  & n14391 ;
  assign n38066 = n14384 & n38065 ;
  assign n38067 = ~n38064 & ~n38066 ;
  assign n38068 = \m6_addr_i[4]_pad  & n14391 ;
  assign n38069 = n14408 & n38068 ;
  assign n38070 = \m2_addr_i[4]_pad  & n14391 ;
  assign n38071 = n14416 & n38070 ;
  assign n38072 = ~n38069 & ~n38071 ;
  assign n38073 = n38067 & n38072 ;
  assign n38074 = \m5_addr_i[4]_pad  & ~n14391 ;
  assign n38075 = n14384 & n38074 ;
  assign n38076 = \m1_addr_i[4]_pad  & ~n14391 ;
  assign n38077 = n14399 & n38076 ;
  assign n38078 = ~n38075 & ~n38077 ;
  assign n38079 = \m0_addr_i[4]_pad  & n14391 ;
  assign n38080 = n14399 & n38079 ;
  assign n38081 = \m7_addr_i[4]_pad  & ~n14391 ;
  assign n38082 = n14408 & n38081 ;
  assign n38083 = ~n38080 & ~n38082 ;
  assign n38084 = n38078 & n38083 ;
  assign n38085 = n38073 & n38084 ;
  assign n38086 = \m3_addr_i[5]_pad  & ~n14391 ;
  assign n38087 = n14416 & n38086 ;
  assign n38088 = \m4_addr_i[5]_pad  & n14391 ;
  assign n38089 = n14384 & n38088 ;
  assign n38090 = ~n38087 & ~n38089 ;
  assign n38091 = \m6_addr_i[5]_pad  & n14391 ;
  assign n38092 = n14408 & n38091 ;
  assign n38093 = \m2_addr_i[5]_pad  & n14391 ;
  assign n38094 = n14416 & n38093 ;
  assign n38095 = ~n38092 & ~n38094 ;
  assign n38096 = n38090 & n38095 ;
  assign n38097 = \m5_addr_i[5]_pad  & ~n14391 ;
  assign n38098 = n14384 & n38097 ;
  assign n38099 = \m1_addr_i[5]_pad  & ~n14391 ;
  assign n38100 = n14399 & n38099 ;
  assign n38101 = ~n38098 & ~n38100 ;
  assign n38102 = \m0_addr_i[5]_pad  & n14391 ;
  assign n38103 = n14399 & n38102 ;
  assign n38104 = \m7_addr_i[5]_pad  & ~n14391 ;
  assign n38105 = n14408 & n38104 ;
  assign n38106 = ~n38103 & ~n38105 ;
  assign n38107 = n38101 & n38106 ;
  assign n38108 = n38096 & n38107 ;
  assign n38109 = \m3_addr_i[6]_pad  & ~n14391 ;
  assign n38110 = n14416 & n38109 ;
  assign n38111 = \m4_addr_i[6]_pad  & n14391 ;
  assign n38112 = n14384 & n38111 ;
  assign n38113 = ~n38110 & ~n38112 ;
  assign n38114 = \m6_addr_i[6]_pad  & n14391 ;
  assign n38115 = n14408 & n38114 ;
  assign n38116 = \m2_addr_i[6]_pad  & n14391 ;
  assign n38117 = n14416 & n38116 ;
  assign n38118 = ~n38115 & ~n38117 ;
  assign n38119 = n38113 & n38118 ;
  assign n38120 = \m5_addr_i[6]_pad  & ~n14391 ;
  assign n38121 = n14384 & n38120 ;
  assign n38122 = \m1_addr_i[6]_pad  & ~n14391 ;
  assign n38123 = n14399 & n38122 ;
  assign n38124 = ~n38121 & ~n38123 ;
  assign n38125 = \m0_addr_i[6]_pad  & n14391 ;
  assign n38126 = n14399 & n38125 ;
  assign n38127 = \m7_addr_i[6]_pad  & ~n14391 ;
  assign n38128 = n14408 & n38127 ;
  assign n38129 = ~n38126 & ~n38128 ;
  assign n38130 = n38124 & n38129 ;
  assign n38131 = n38119 & n38130 ;
  assign n38132 = \m3_addr_i[7]_pad  & ~n14391 ;
  assign n38133 = n14416 & n38132 ;
  assign n38134 = \m4_addr_i[7]_pad  & n14391 ;
  assign n38135 = n14384 & n38134 ;
  assign n38136 = ~n38133 & ~n38135 ;
  assign n38137 = \m6_addr_i[7]_pad  & n14391 ;
  assign n38138 = n14408 & n38137 ;
  assign n38139 = \m2_addr_i[7]_pad  & n14391 ;
  assign n38140 = n14416 & n38139 ;
  assign n38141 = ~n38138 & ~n38140 ;
  assign n38142 = n38136 & n38141 ;
  assign n38143 = \m5_addr_i[7]_pad  & ~n14391 ;
  assign n38144 = n14384 & n38143 ;
  assign n38145 = \m1_addr_i[7]_pad  & ~n14391 ;
  assign n38146 = n14399 & n38145 ;
  assign n38147 = ~n38144 & ~n38146 ;
  assign n38148 = \m0_addr_i[7]_pad  & n14391 ;
  assign n38149 = n14399 & n38148 ;
  assign n38150 = \m7_addr_i[7]_pad  & ~n14391 ;
  assign n38151 = n14408 & n38150 ;
  assign n38152 = ~n38149 & ~n38151 ;
  assign n38153 = n38147 & n38152 ;
  assign n38154 = n38142 & n38153 ;
  assign n38155 = \m3_addr_i[8]_pad  & ~n14391 ;
  assign n38156 = n14416 & n38155 ;
  assign n38157 = \m4_addr_i[8]_pad  & n14391 ;
  assign n38158 = n14384 & n38157 ;
  assign n38159 = ~n38156 & ~n38158 ;
  assign n38160 = \m6_addr_i[8]_pad  & n14391 ;
  assign n38161 = n14408 & n38160 ;
  assign n38162 = \m2_addr_i[8]_pad  & n14391 ;
  assign n38163 = n14416 & n38162 ;
  assign n38164 = ~n38161 & ~n38163 ;
  assign n38165 = n38159 & n38164 ;
  assign n38166 = \m5_addr_i[8]_pad  & ~n14391 ;
  assign n38167 = n14384 & n38166 ;
  assign n38168 = \m1_addr_i[8]_pad  & ~n14391 ;
  assign n38169 = n14399 & n38168 ;
  assign n38170 = ~n38167 & ~n38169 ;
  assign n38171 = \m0_addr_i[8]_pad  & n14391 ;
  assign n38172 = n14399 & n38171 ;
  assign n38173 = \m7_addr_i[8]_pad  & ~n14391 ;
  assign n38174 = n14408 & n38173 ;
  assign n38175 = ~n38172 & ~n38174 ;
  assign n38176 = n38170 & n38175 ;
  assign n38177 = n38165 & n38176 ;
  assign n38178 = \m3_addr_i[9]_pad  & ~n14391 ;
  assign n38179 = n14416 & n38178 ;
  assign n38180 = \m4_addr_i[9]_pad  & n14391 ;
  assign n38181 = n14384 & n38180 ;
  assign n38182 = ~n38179 & ~n38181 ;
  assign n38183 = \m6_addr_i[9]_pad  & n14391 ;
  assign n38184 = n14408 & n38183 ;
  assign n38185 = \m2_addr_i[9]_pad  & n14391 ;
  assign n38186 = n14416 & n38185 ;
  assign n38187 = ~n38184 & ~n38186 ;
  assign n38188 = n38182 & n38187 ;
  assign n38189 = \m5_addr_i[9]_pad  & ~n14391 ;
  assign n38190 = n14384 & n38189 ;
  assign n38191 = \m1_addr_i[9]_pad  & ~n14391 ;
  assign n38192 = n14399 & n38191 ;
  assign n38193 = ~n38190 & ~n38192 ;
  assign n38194 = \m0_addr_i[9]_pad  & n14391 ;
  assign n38195 = n14399 & n38194 ;
  assign n38196 = \m7_addr_i[9]_pad  & ~n14391 ;
  assign n38197 = n14408 & n38196 ;
  assign n38198 = ~n38195 & ~n38197 ;
  assign n38199 = n38193 & n38198 ;
  assign n38200 = n38188 & n38199 ;
  assign n38201 = \m3_data_i[0]_pad  & ~n14391 ;
  assign n38202 = n14416 & n38201 ;
  assign n38203 = \m4_data_i[0]_pad  & n14391 ;
  assign n38204 = n14384 & n38203 ;
  assign n38205 = ~n38202 & ~n38204 ;
  assign n38206 = \m6_data_i[0]_pad  & n14391 ;
  assign n38207 = n14408 & n38206 ;
  assign n38208 = \m2_data_i[0]_pad  & n14391 ;
  assign n38209 = n14416 & n38208 ;
  assign n38210 = ~n38207 & ~n38209 ;
  assign n38211 = n38205 & n38210 ;
  assign n38212 = \m5_data_i[0]_pad  & ~n14391 ;
  assign n38213 = n14384 & n38212 ;
  assign n38214 = \m1_data_i[0]_pad  & ~n14391 ;
  assign n38215 = n14399 & n38214 ;
  assign n38216 = ~n38213 & ~n38215 ;
  assign n38217 = \m0_data_i[0]_pad  & n14391 ;
  assign n38218 = n14399 & n38217 ;
  assign n38219 = \m7_data_i[0]_pad  & ~n14391 ;
  assign n38220 = n14408 & n38219 ;
  assign n38221 = ~n38218 & ~n38220 ;
  assign n38222 = n38216 & n38221 ;
  assign n38223 = n38211 & n38222 ;
  assign n38224 = \m3_data_i[10]_pad  & ~n14391 ;
  assign n38225 = n14416 & n38224 ;
  assign n38226 = \m4_data_i[10]_pad  & n14391 ;
  assign n38227 = n14384 & n38226 ;
  assign n38228 = ~n38225 & ~n38227 ;
  assign n38229 = \m6_data_i[10]_pad  & n14391 ;
  assign n38230 = n14408 & n38229 ;
  assign n38231 = \m2_data_i[10]_pad  & n14391 ;
  assign n38232 = n14416 & n38231 ;
  assign n38233 = ~n38230 & ~n38232 ;
  assign n38234 = n38228 & n38233 ;
  assign n38235 = \m5_data_i[10]_pad  & ~n14391 ;
  assign n38236 = n14384 & n38235 ;
  assign n38237 = \m1_data_i[10]_pad  & ~n14391 ;
  assign n38238 = n14399 & n38237 ;
  assign n38239 = ~n38236 & ~n38238 ;
  assign n38240 = \m0_data_i[10]_pad  & n14391 ;
  assign n38241 = n14399 & n38240 ;
  assign n38242 = \m7_data_i[10]_pad  & ~n14391 ;
  assign n38243 = n14408 & n38242 ;
  assign n38244 = ~n38241 & ~n38243 ;
  assign n38245 = n38239 & n38244 ;
  assign n38246 = n38234 & n38245 ;
  assign n38247 = \m3_data_i[11]_pad  & ~n14391 ;
  assign n38248 = n14416 & n38247 ;
  assign n38249 = \m4_data_i[11]_pad  & n14391 ;
  assign n38250 = n14384 & n38249 ;
  assign n38251 = ~n38248 & ~n38250 ;
  assign n38252 = \m6_data_i[11]_pad  & n14391 ;
  assign n38253 = n14408 & n38252 ;
  assign n38254 = \m2_data_i[11]_pad  & n14391 ;
  assign n38255 = n14416 & n38254 ;
  assign n38256 = ~n38253 & ~n38255 ;
  assign n38257 = n38251 & n38256 ;
  assign n38258 = \m5_data_i[11]_pad  & ~n14391 ;
  assign n38259 = n14384 & n38258 ;
  assign n38260 = \m1_data_i[11]_pad  & ~n14391 ;
  assign n38261 = n14399 & n38260 ;
  assign n38262 = ~n38259 & ~n38261 ;
  assign n38263 = \m0_data_i[11]_pad  & n14391 ;
  assign n38264 = n14399 & n38263 ;
  assign n38265 = \m7_data_i[11]_pad  & ~n14391 ;
  assign n38266 = n14408 & n38265 ;
  assign n38267 = ~n38264 & ~n38266 ;
  assign n38268 = n38262 & n38267 ;
  assign n38269 = n38257 & n38268 ;
  assign n38270 = \m3_data_i[12]_pad  & ~n14391 ;
  assign n38271 = n14416 & n38270 ;
  assign n38272 = \m4_data_i[12]_pad  & n14391 ;
  assign n38273 = n14384 & n38272 ;
  assign n38274 = ~n38271 & ~n38273 ;
  assign n38275 = \m6_data_i[12]_pad  & n14391 ;
  assign n38276 = n14408 & n38275 ;
  assign n38277 = \m2_data_i[12]_pad  & n14391 ;
  assign n38278 = n14416 & n38277 ;
  assign n38279 = ~n38276 & ~n38278 ;
  assign n38280 = n38274 & n38279 ;
  assign n38281 = \m5_data_i[12]_pad  & ~n14391 ;
  assign n38282 = n14384 & n38281 ;
  assign n38283 = \m1_data_i[12]_pad  & ~n14391 ;
  assign n38284 = n14399 & n38283 ;
  assign n38285 = ~n38282 & ~n38284 ;
  assign n38286 = \m0_data_i[12]_pad  & n14391 ;
  assign n38287 = n14399 & n38286 ;
  assign n38288 = \m7_data_i[12]_pad  & ~n14391 ;
  assign n38289 = n14408 & n38288 ;
  assign n38290 = ~n38287 & ~n38289 ;
  assign n38291 = n38285 & n38290 ;
  assign n38292 = n38280 & n38291 ;
  assign n38293 = \m3_data_i[13]_pad  & ~n14391 ;
  assign n38294 = n14416 & n38293 ;
  assign n38295 = \m4_data_i[13]_pad  & n14391 ;
  assign n38296 = n14384 & n38295 ;
  assign n38297 = ~n38294 & ~n38296 ;
  assign n38298 = \m6_data_i[13]_pad  & n14391 ;
  assign n38299 = n14408 & n38298 ;
  assign n38300 = \m2_data_i[13]_pad  & n14391 ;
  assign n38301 = n14416 & n38300 ;
  assign n38302 = ~n38299 & ~n38301 ;
  assign n38303 = n38297 & n38302 ;
  assign n38304 = \m5_data_i[13]_pad  & ~n14391 ;
  assign n38305 = n14384 & n38304 ;
  assign n38306 = \m1_data_i[13]_pad  & ~n14391 ;
  assign n38307 = n14399 & n38306 ;
  assign n38308 = ~n38305 & ~n38307 ;
  assign n38309 = \m0_data_i[13]_pad  & n14391 ;
  assign n38310 = n14399 & n38309 ;
  assign n38311 = \m7_data_i[13]_pad  & ~n14391 ;
  assign n38312 = n14408 & n38311 ;
  assign n38313 = ~n38310 & ~n38312 ;
  assign n38314 = n38308 & n38313 ;
  assign n38315 = n38303 & n38314 ;
  assign n38316 = \m3_data_i[14]_pad  & ~n14391 ;
  assign n38317 = n14416 & n38316 ;
  assign n38318 = \m4_data_i[14]_pad  & n14391 ;
  assign n38319 = n14384 & n38318 ;
  assign n38320 = ~n38317 & ~n38319 ;
  assign n38321 = \m6_data_i[14]_pad  & n14391 ;
  assign n38322 = n14408 & n38321 ;
  assign n38323 = \m2_data_i[14]_pad  & n14391 ;
  assign n38324 = n14416 & n38323 ;
  assign n38325 = ~n38322 & ~n38324 ;
  assign n38326 = n38320 & n38325 ;
  assign n38327 = \m5_data_i[14]_pad  & ~n14391 ;
  assign n38328 = n14384 & n38327 ;
  assign n38329 = \m1_data_i[14]_pad  & ~n14391 ;
  assign n38330 = n14399 & n38329 ;
  assign n38331 = ~n38328 & ~n38330 ;
  assign n38332 = \m0_data_i[14]_pad  & n14391 ;
  assign n38333 = n14399 & n38332 ;
  assign n38334 = \m7_data_i[14]_pad  & ~n14391 ;
  assign n38335 = n14408 & n38334 ;
  assign n38336 = ~n38333 & ~n38335 ;
  assign n38337 = n38331 & n38336 ;
  assign n38338 = n38326 & n38337 ;
  assign n38339 = \m3_data_i[15]_pad  & ~n14391 ;
  assign n38340 = n14416 & n38339 ;
  assign n38341 = \m4_data_i[15]_pad  & n14391 ;
  assign n38342 = n14384 & n38341 ;
  assign n38343 = ~n38340 & ~n38342 ;
  assign n38344 = \m6_data_i[15]_pad  & n14391 ;
  assign n38345 = n14408 & n38344 ;
  assign n38346 = \m2_data_i[15]_pad  & n14391 ;
  assign n38347 = n14416 & n38346 ;
  assign n38348 = ~n38345 & ~n38347 ;
  assign n38349 = n38343 & n38348 ;
  assign n38350 = \m5_data_i[15]_pad  & ~n14391 ;
  assign n38351 = n14384 & n38350 ;
  assign n38352 = \m1_data_i[15]_pad  & ~n14391 ;
  assign n38353 = n14399 & n38352 ;
  assign n38354 = ~n38351 & ~n38353 ;
  assign n38355 = \m0_data_i[15]_pad  & n14391 ;
  assign n38356 = n14399 & n38355 ;
  assign n38357 = \m7_data_i[15]_pad  & ~n14391 ;
  assign n38358 = n14408 & n38357 ;
  assign n38359 = ~n38356 & ~n38358 ;
  assign n38360 = n38354 & n38359 ;
  assign n38361 = n38349 & n38360 ;
  assign n38362 = \m3_data_i[16]_pad  & ~n14391 ;
  assign n38363 = n14416 & n38362 ;
  assign n38364 = \m4_data_i[16]_pad  & n14391 ;
  assign n38365 = n14384 & n38364 ;
  assign n38366 = ~n38363 & ~n38365 ;
  assign n38367 = \m6_data_i[16]_pad  & n14391 ;
  assign n38368 = n14408 & n38367 ;
  assign n38369 = \m2_data_i[16]_pad  & n14391 ;
  assign n38370 = n14416 & n38369 ;
  assign n38371 = ~n38368 & ~n38370 ;
  assign n38372 = n38366 & n38371 ;
  assign n38373 = \m5_data_i[16]_pad  & ~n14391 ;
  assign n38374 = n14384 & n38373 ;
  assign n38375 = \m1_data_i[16]_pad  & ~n14391 ;
  assign n38376 = n14399 & n38375 ;
  assign n38377 = ~n38374 & ~n38376 ;
  assign n38378 = \m0_data_i[16]_pad  & n14391 ;
  assign n38379 = n14399 & n38378 ;
  assign n38380 = \m7_data_i[16]_pad  & ~n14391 ;
  assign n38381 = n14408 & n38380 ;
  assign n38382 = ~n38379 & ~n38381 ;
  assign n38383 = n38377 & n38382 ;
  assign n38384 = n38372 & n38383 ;
  assign n38385 = \m3_data_i[17]_pad  & ~n14391 ;
  assign n38386 = n14416 & n38385 ;
  assign n38387 = \m4_data_i[17]_pad  & n14391 ;
  assign n38388 = n14384 & n38387 ;
  assign n38389 = ~n38386 & ~n38388 ;
  assign n38390 = \m6_data_i[17]_pad  & n14391 ;
  assign n38391 = n14408 & n38390 ;
  assign n38392 = \m2_data_i[17]_pad  & n14391 ;
  assign n38393 = n14416 & n38392 ;
  assign n38394 = ~n38391 & ~n38393 ;
  assign n38395 = n38389 & n38394 ;
  assign n38396 = \m5_data_i[17]_pad  & ~n14391 ;
  assign n38397 = n14384 & n38396 ;
  assign n38398 = \m1_data_i[17]_pad  & ~n14391 ;
  assign n38399 = n14399 & n38398 ;
  assign n38400 = ~n38397 & ~n38399 ;
  assign n38401 = \m0_data_i[17]_pad  & n14391 ;
  assign n38402 = n14399 & n38401 ;
  assign n38403 = \m7_data_i[17]_pad  & ~n14391 ;
  assign n38404 = n14408 & n38403 ;
  assign n38405 = ~n38402 & ~n38404 ;
  assign n38406 = n38400 & n38405 ;
  assign n38407 = n38395 & n38406 ;
  assign n38408 = \m3_data_i[18]_pad  & ~n14391 ;
  assign n38409 = n14416 & n38408 ;
  assign n38410 = \m4_data_i[18]_pad  & n14391 ;
  assign n38411 = n14384 & n38410 ;
  assign n38412 = ~n38409 & ~n38411 ;
  assign n38413 = \m6_data_i[18]_pad  & n14391 ;
  assign n38414 = n14408 & n38413 ;
  assign n38415 = \m2_data_i[18]_pad  & n14391 ;
  assign n38416 = n14416 & n38415 ;
  assign n38417 = ~n38414 & ~n38416 ;
  assign n38418 = n38412 & n38417 ;
  assign n38419 = \m5_data_i[18]_pad  & ~n14391 ;
  assign n38420 = n14384 & n38419 ;
  assign n38421 = \m1_data_i[18]_pad  & ~n14391 ;
  assign n38422 = n14399 & n38421 ;
  assign n38423 = ~n38420 & ~n38422 ;
  assign n38424 = \m0_data_i[18]_pad  & n14391 ;
  assign n38425 = n14399 & n38424 ;
  assign n38426 = \m7_data_i[18]_pad  & ~n14391 ;
  assign n38427 = n14408 & n38426 ;
  assign n38428 = ~n38425 & ~n38427 ;
  assign n38429 = n38423 & n38428 ;
  assign n38430 = n38418 & n38429 ;
  assign n38431 = \m3_data_i[19]_pad  & ~n14391 ;
  assign n38432 = n14416 & n38431 ;
  assign n38433 = \m4_data_i[19]_pad  & n14391 ;
  assign n38434 = n14384 & n38433 ;
  assign n38435 = ~n38432 & ~n38434 ;
  assign n38436 = \m6_data_i[19]_pad  & n14391 ;
  assign n38437 = n14408 & n38436 ;
  assign n38438 = \m2_data_i[19]_pad  & n14391 ;
  assign n38439 = n14416 & n38438 ;
  assign n38440 = ~n38437 & ~n38439 ;
  assign n38441 = n38435 & n38440 ;
  assign n38442 = \m5_data_i[19]_pad  & ~n14391 ;
  assign n38443 = n14384 & n38442 ;
  assign n38444 = \m1_data_i[19]_pad  & ~n14391 ;
  assign n38445 = n14399 & n38444 ;
  assign n38446 = ~n38443 & ~n38445 ;
  assign n38447 = \m0_data_i[19]_pad  & n14391 ;
  assign n38448 = n14399 & n38447 ;
  assign n38449 = \m7_data_i[19]_pad  & ~n14391 ;
  assign n38450 = n14408 & n38449 ;
  assign n38451 = ~n38448 & ~n38450 ;
  assign n38452 = n38446 & n38451 ;
  assign n38453 = n38441 & n38452 ;
  assign n38454 = \m3_data_i[1]_pad  & ~n14391 ;
  assign n38455 = n14416 & n38454 ;
  assign n38456 = \m4_data_i[1]_pad  & n14391 ;
  assign n38457 = n14384 & n38456 ;
  assign n38458 = ~n38455 & ~n38457 ;
  assign n38459 = \m6_data_i[1]_pad  & n14391 ;
  assign n38460 = n14408 & n38459 ;
  assign n38461 = \m2_data_i[1]_pad  & n14391 ;
  assign n38462 = n14416 & n38461 ;
  assign n38463 = ~n38460 & ~n38462 ;
  assign n38464 = n38458 & n38463 ;
  assign n38465 = \m5_data_i[1]_pad  & ~n14391 ;
  assign n38466 = n14384 & n38465 ;
  assign n38467 = \m1_data_i[1]_pad  & ~n14391 ;
  assign n38468 = n14399 & n38467 ;
  assign n38469 = ~n38466 & ~n38468 ;
  assign n38470 = \m0_data_i[1]_pad  & n14391 ;
  assign n38471 = n14399 & n38470 ;
  assign n38472 = \m7_data_i[1]_pad  & ~n14391 ;
  assign n38473 = n14408 & n38472 ;
  assign n38474 = ~n38471 & ~n38473 ;
  assign n38475 = n38469 & n38474 ;
  assign n38476 = n38464 & n38475 ;
  assign n38477 = \m3_data_i[20]_pad  & ~n14391 ;
  assign n38478 = n14416 & n38477 ;
  assign n38479 = \m4_data_i[20]_pad  & n14391 ;
  assign n38480 = n14384 & n38479 ;
  assign n38481 = ~n38478 & ~n38480 ;
  assign n38482 = \m6_data_i[20]_pad  & n14391 ;
  assign n38483 = n14408 & n38482 ;
  assign n38484 = \m2_data_i[20]_pad  & n14391 ;
  assign n38485 = n14416 & n38484 ;
  assign n38486 = ~n38483 & ~n38485 ;
  assign n38487 = n38481 & n38486 ;
  assign n38488 = \m5_data_i[20]_pad  & ~n14391 ;
  assign n38489 = n14384 & n38488 ;
  assign n38490 = \m1_data_i[20]_pad  & ~n14391 ;
  assign n38491 = n14399 & n38490 ;
  assign n38492 = ~n38489 & ~n38491 ;
  assign n38493 = \m0_data_i[20]_pad  & n14391 ;
  assign n38494 = n14399 & n38493 ;
  assign n38495 = \m7_data_i[20]_pad  & ~n14391 ;
  assign n38496 = n14408 & n38495 ;
  assign n38497 = ~n38494 & ~n38496 ;
  assign n38498 = n38492 & n38497 ;
  assign n38499 = n38487 & n38498 ;
  assign n38500 = \m3_data_i[21]_pad  & ~n14391 ;
  assign n38501 = n14416 & n38500 ;
  assign n38502 = \m4_data_i[21]_pad  & n14391 ;
  assign n38503 = n14384 & n38502 ;
  assign n38504 = ~n38501 & ~n38503 ;
  assign n38505 = \m6_data_i[21]_pad  & n14391 ;
  assign n38506 = n14408 & n38505 ;
  assign n38507 = \m2_data_i[21]_pad  & n14391 ;
  assign n38508 = n14416 & n38507 ;
  assign n38509 = ~n38506 & ~n38508 ;
  assign n38510 = n38504 & n38509 ;
  assign n38511 = \m5_data_i[21]_pad  & ~n14391 ;
  assign n38512 = n14384 & n38511 ;
  assign n38513 = \m1_data_i[21]_pad  & ~n14391 ;
  assign n38514 = n14399 & n38513 ;
  assign n38515 = ~n38512 & ~n38514 ;
  assign n38516 = \m0_data_i[21]_pad  & n14391 ;
  assign n38517 = n14399 & n38516 ;
  assign n38518 = \m7_data_i[21]_pad  & ~n14391 ;
  assign n38519 = n14408 & n38518 ;
  assign n38520 = ~n38517 & ~n38519 ;
  assign n38521 = n38515 & n38520 ;
  assign n38522 = n38510 & n38521 ;
  assign n38523 = \m3_data_i[22]_pad  & ~n14391 ;
  assign n38524 = n14416 & n38523 ;
  assign n38525 = \m4_data_i[22]_pad  & n14391 ;
  assign n38526 = n14384 & n38525 ;
  assign n38527 = ~n38524 & ~n38526 ;
  assign n38528 = \m6_data_i[22]_pad  & n14391 ;
  assign n38529 = n14408 & n38528 ;
  assign n38530 = \m2_data_i[22]_pad  & n14391 ;
  assign n38531 = n14416 & n38530 ;
  assign n38532 = ~n38529 & ~n38531 ;
  assign n38533 = n38527 & n38532 ;
  assign n38534 = \m5_data_i[22]_pad  & ~n14391 ;
  assign n38535 = n14384 & n38534 ;
  assign n38536 = \m1_data_i[22]_pad  & ~n14391 ;
  assign n38537 = n14399 & n38536 ;
  assign n38538 = ~n38535 & ~n38537 ;
  assign n38539 = \m0_data_i[22]_pad  & n14391 ;
  assign n38540 = n14399 & n38539 ;
  assign n38541 = \m7_data_i[22]_pad  & ~n14391 ;
  assign n38542 = n14408 & n38541 ;
  assign n38543 = ~n38540 & ~n38542 ;
  assign n38544 = n38538 & n38543 ;
  assign n38545 = n38533 & n38544 ;
  assign n38546 = \m3_data_i[23]_pad  & ~n14391 ;
  assign n38547 = n14416 & n38546 ;
  assign n38548 = \m4_data_i[23]_pad  & n14391 ;
  assign n38549 = n14384 & n38548 ;
  assign n38550 = ~n38547 & ~n38549 ;
  assign n38551 = \m6_data_i[23]_pad  & n14391 ;
  assign n38552 = n14408 & n38551 ;
  assign n38553 = \m2_data_i[23]_pad  & n14391 ;
  assign n38554 = n14416 & n38553 ;
  assign n38555 = ~n38552 & ~n38554 ;
  assign n38556 = n38550 & n38555 ;
  assign n38557 = \m5_data_i[23]_pad  & ~n14391 ;
  assign n38558 = n14384 & n38557 ;
  assign n38559 = \m1_data_i[23]_pad  & ~n14391 ;
  assign n38560 = n14399 & n38559 ;
  assign n38561 = ~n38558 & ~n38560 ;
  assign n38562 = \m0_data_i[23]_pad  & n14391 ;
  assign n38563 = n14399 & n38562 ;
  assign n38564 = \m7_data_i[23]_pad  & ~n14391 ;
  assign n38565 = n14408 & n38564 ;
  assign n38566 = ~n38563 & ~n38565 ;
  assign n38567 = n38561 & n38566 ;
  assign n38568 = n38556 & n38567 ;
  assign n38569 = \m3_data_i[24]_pad  & ~n14391 ;
  assign n38570 = n14416 & n38569 ;
  assign n38571 = \m4_data_i[24]_pad  & n14391 ;
  assign n38572 = n14384 & n38571 ;
  assign n38573 = ~n38570 & ~n38572 ;
  assign n38574 = \m6_data_i[24]_pad  & n14391 ;
  assign n38575 = n14408 & n38574 ;
  assign n38576 = \m2_data_i[24]_pad  & n14391 ;
  assign n38577 = n14416 & n38576 ;
  assign n38578 = ~n38575 & ~n38577 ;
  assign n38579 = n38573 & n38578 ;
  assign n38580 = \m5_data_i[24]_pad  & ~n14391 ;
  assign n38581 = n14384 & n38580 ;
  assign n38582 = \m1_data_i[24]_pad  & ~n14391 ;
  assign n38583 = n14399 & n38582 ;
  assign n38584 = ~n38581 & ~n38583 ;
  assign n38585 = \m0_data_i[24]_pad  & n14391 ;
  assign n38586 = n14399 & n38585 ;
  assign n38587 = \m7_data_i[24]_pad  & ~n14391 ;
  assign n38588 = n14408 & n38587 ;
  assign n38589 = ~n38586 & ~n38588 ;
  assign n38590 = n38584 & n38589 ;
  assign n38591 = n38579 & n38590 ;
  assign n38592 = \m3_data_i[25]_pad  & ~n14391 ;
  assign n38593 = n14416 & n38592 ;
  assign n38594 = \m4_data_i[25]_pad  & n14391 ;
  assign n38595 = n14384 & n38594 ;
  assign n38596 = ~n38593 & ~n38595 ;
  assign n38597 = \m6_data_i[25]_pad  & n14391 ;
  assign n38598 = n14408 & n38597 ;
  assign n38599 = \m2_data_i[25]_pad  & n14391 ;
  assign n38600 = n14416 & n38599 ;
  assign n38601 = ~n38598 & ~n38600 ;
  assign n38602 = n38596 & n38601 ;
  assign n38603 = \m5_data_i[25]_pad  & ~n14391 ;
  assign n38604 = n14384 & n38603 ;
  assign n38605 = \m1_data_i[25]_pad  & ~n14391 ;
  assign n38606 = n14399 & n38605 ;
  assign n38607 = ~n38604 & ~n38606 ;
  assign n38608 = \m0_data_i[25]_pad  & n14391 ;
  assign n38609 = n14399 & n38608 ;
  assign n38610 = \m7_data_i[25]_pad  & ~n14391 ;
  assign n38611 = n14408 & n38610 ;
  assign n38612 = ~n38609 & ~n38611 ;
  assign n38613 = n38607 & n38612 ;
  assign n38614 = n38602 & n38613 ;
  assign n38615 = \m0_data_i[26]_pad  & n14391 ;
  assign n38616 = n14399 & n38615 ;
  assign n38617 = \m7_data_i[26]_pad  & ~n14391 ;
  assign n38618 = n14408 & n38617 ;
  assign n38619 = ~n38616 & ~n38618 ;
  assign n38620 = \m1_data_i[26]_pad  & ~n14391 ;
  assign n38621 = n14399 & n38620 ;
  assign n38622 = \m4_data_i[26]_pad  & n14391 ;
  assign n38623 = n14384 & n38622 ;
  assign n38624 = ~n38621 & ~n38623 ;
  assign n38625 = n38619 & n38624 ;
  assign n38626 = \m2_data_i[26]_pad  & n14391 ;
  assign n38627 = n14416 & n38626 ;
  assign n38628 = \m3_data_i[26]_pad  & ~n14391 ;
  assign n38629 = n14416 & n38628 ;
  assign n38630 = ~n38627 & ~n38629 ;
  assign n38631 = \m6_data_i[26]_pad  & n14391 ;
  assign n38632 = n14408 & n38631 ;
  assign n38633 = \m5_data_i[26]_pad  & ~n14391 ;
  assign n38634 = n14384 & n38633 ;
  assign n38635 = ~n38632 & ~n38634 ;
  assign n38636 = n38630 & n38635 ;
  assign n38637 = n38625 & n38636 ;
  assign n38638 = \m1_data_i[27]_pad  & ~n14391 ;
  assign n38639 = n14399 & n38638 ;
  assign n38640 = \m2_data_i[27]_pad  & n14391 ;
  assign n38641 = n14416 & n38640 ;
  assign n38642 = ~n38639 & ~n38641 ;
  assign n38643 = \m6_data_i[27]_pad  & n14391 ;
  assign n38644 = n14408 & n38643 ;
  assign n38645 = \m7_data_i[27]_pad  & ~n14391 ;
  assign n38646 = n14408 & n38645 ;
  assign n38647 = ~n38644 & ~n38646 ;
  assign n38648 = n38642 & n38647 ;
  assign n38649 = \m5_data_i[27]_pad  & ~n14391 ;
  assign n38650 = n14384 & n38649 ;
  assign n38651 = \m0_data_i[27]_pad  & n14391 ;
  assign n38652 = n14399 & n38651 ;
  assign n38653 = ~n38650 & ~n38652 ;
  assign n38654 = \m3_data_i[27]_pad  & ~n14391 ;
  assign n38655 = n14416 & n38654 ;
  assign n38656 = \m4_data_i[27]_pad  & n14391 ;
  assign n38657 = n14384 & n38656 ;
  assign n38658 = ~n38655 & ~n38657 ;
  assign n38659 = n38653 & n38658 ;
  assign n38660 = n38648 & n38659 ;
  assign n38661 = \m1_data_i[28]_pad  & ~n14391 ;
  assign n38662 = n14399 & n38661 ;
  assign n38663 = \m2_data_i[28]_pad  & n14391 ;
  assign n38664 = n14416 & n38663 ;
  assign n38665 = ~n38662 & ~n38664 ;
  assign n38666 = \m0_data_i[28]_pad  & n14391 ;
  assign n38667 = n14399 & n38666 ;
  assign n38668 = \m4_data_i[28]_pad  & n14391 ;
  assign n38669 = n14384 & n38668 ;
  assign n38670 = ~n38667 & ~n38669 ;
  assign n38671 = n38665 & n38670 ;
  assign n38672 = \m7_data_i[28]_pad  & ~n14391 ;
  assign n38673 = n14408 & n38672 ;
  assign n38674 = \m3_data_i[28]_pad  & ~n14391 ;
  assign n38675 = n14416 & n38674 ;
  assign n38676 = ~n38673 & ~n38675 ;
  assign n38677 = \m6_data_i[28]_pad  & n14391 ;
  assign n38678 = n14408 & n38677 ;
  assign n38679 = \m5_data_i[28]_pad  & ~n14391 ;
  assign n38680 = n14384 & n38679 ;
  assign n38681 = ~n38678 & ~n38680 ;
  assign n38682 = n38676 & n38681 ;
  assign n38683 = n38671 & n38682 ;
  assign n38684 = \m3_data_i[29]_pad  & ~n14391 ;
  assign n38685 = n14416 & n38684 ;
  assign n38686 = \m4_data_i[29]_pad  & n14391 ;
  assign n38687 = n14384 & n38686 ;
  assign n38688 = ~n38685 & ~n38687 ;
  assign n38689 = \m6_data_i[29]_pad  & n14391 ;
  assign n38690 = n14408 & n38689 ;
  assign n38691 = \m7_data_i[29]_pad  & ~n14391 ;
  assign n38692 = n14408 & n38691 ;
  assign n38693 = ~n38690 & ~n38692 ;
  assign n38694 = n38688 & n38693 ;
  assign n38695 = \m5_data_i[29]_pad  & ~n14391 ;
  assign n38696 = n14384 & n38695 ;
  assign n38697 = \m0_data_i[29]_pad  & n14391 ;
  assign n38698 = n14399 & n38697 ;
  assign n38699 = ~n38696 & ~n38698 ;
  assign n38700 = \m1_data_i[29]_pad  & ~n14391 ;
  assign n38701 = n14399 & n38700 ;
  assign n38702 = \m2_data_i[29]_pad  & n14391 ;
  assign n38703 = n14416 & n38702 ;
  assign n38704 = ~n38701 & ~n38703 ;
  assign n38705 = n38699 & n38704 ;
  assign n38706 = n38694 & n38705 ;
  assign n38707 = \m3_data_i[2]_pad  & ~n14391 ;
  assign n38708 = n14416 & n38707 ;
  assign n38709 = \m4_data_i[2]_pad  & n14391 ;
  assign n38710 = n14384 & n38709 ;
  assign n38711 = ~n38708 & ~n38710 ;
  assign n38712 = \m6_data_i[2]_pad  & n14391 ;
  assign n38713 = n14408 & n38712 ;
  assign n38714 = \m2_data_i[2]_pad  & n14391 ;
  assign n38715 = n14416 & n38714 ;
  assign n38716 = ~n38713 & ~n38715 ;
  assign n38717 = n38711 & n38716 ;
  assign n38718 = \m5_data_i[2]_pad  & ~n14391 ;
  assign n38719 = n14384 & n38718 ;
  assign n38720 = \m1_data_i[2]_pad  & ~n14391 ;
  assign n38721 = n14399 & n38720 ;
  assign n38722 = ~n38719 & ~n38721 ;
  assign n38723 = \m0_data_i[2]_pad  & n14391 ;
  assign n38724 = n14399 & n38723 ;
  assign n38725 = \m7_data_i[2]_pad  & ~n14391 ;
  assign n38726 = n14408 & n38725 ;
  assign n38727 = ~n38724 & ~n38726 ;
  assign n38728 = n38722 & n38727 ;
  assign n38729 = n38717 & n38728 ;
  assign n38730 = \m1_data_i[30]_pad  & ~n14391 ;
  assign n38731 = n14399 & n38730 ;
  assign n38732 = \m2_data_i[30]_pad  & n14391 ;
  assign n38733 = n14416 & n38732 ;
  assign n38734 = ~n38731 & ~n38733 ;
  assign n38735 = \m3_data_i[30]_pad  & ~n14391 ;
  assign n38736 = n14416 & n38735 ;
  assign n38737 = \m7_data_i[30]_pad  & ~n14391 ;
  assign n38738 = n14408 & n38737 ;
  assign n38739 = ~n38736 & ~n38738 ;
  assign n38740 = n38734 & n38739 ;
  assign n38741 = \m4_data_i[30]_pad  & n14391 ;
  assign n38742 = n14384 & n38741 ;
  assign n38743 = \m0_data_i[30]_pad  & n14391 ;
  assign n38744 = n14399 & n38743 ;
  assign n38745 = ~n38742 & ~n38744 ;
  assign n38746 = \m6_data_i[30]_pad  & n14391 ;
  assign n38747 = n14408 & n38746 ;
  assign n38748 = \m5_data_i[30]_pad  & ~n14391 ;
  assign n38749 = n14384 & n38748 ;
  assign n38750 = ~n38747 & ~n38749 ;
  assign n38751 = n38745 & n38750 ;
  assign n38752 = n38740 & n38751 ;
  assign n38753 = \m1_data_i[31]_pad  & ~n14391 ;
  assign n38754 = n14399 & n38753 ;
  assign n38755 = \m2_data_i[31]_pad  & n14391 ;
  assign n38756 = n14416 & n38755 ;
  assign n38757 = ~n38754 & ~n38756 ;
  assign n38758 = \m6_data_i[31]_pad  & n14391 ;
  assign n38759 = n14408 & n38758 ;
  assign n38760 = \m4_data_i[31]_pad  & n14391 ;
  assign n38761 = n14384 & n38760 ;
  assign n38762 = ~n38759 & ~n38761 ;
  assign n38763 = n38757 & n38762 ;
  assign n38764 = \m5_data_i[31]_pad  & ~n14391 ;
  assign n38765 = n14384 & n38764 ;
  assign n38766 = \m3_data_i[31]_pad  & ~n14391 ;
  assign n38767 = n14416 & n38766 ;
  assign n38768 = ~n38765 & ~n38767 ;
  assign n38769 = \m0_data_i[31]_pad  & n14391 ;
  assign n38770 = n14399 & n38769 ;
  assign n38771 = \m7_data_i[31]_pad  & ~n14391 ;
  assign n38772 = n14408 & n38771 ;
  assign n38773 = ~n38770 & ~n38772 ;
  assign n38774 = n38768 & n38773 ;
  assign n38775 = n38763 & n38774 ;
  assign n38776 = \m3_data_i[3]_pad  & ~n14391 ;
  assign n38777 = n14416 & n38776 ;
  assign n38778 = \m4_data_i[3]_pad  & n14391 ;
  assign n38779 = n14384 & n38778 ;
  assign n38780 = ~n38777 & ~n38779 ;
  assign n38781 = \m6_data_i[3]_pad  & n14391 ;
  assign n38782 = n14408 & n38781 ;
  assign n38783 = \m2_data_i[3]_pad  & n14391 ;
  assign n38784 = n14416 & n38783 ;
  assign n38785 = ~n38782 & ~n38784 ;
  assign n38786 = n38780 & n38785 ;
  assign n38787 = \m5_data_i[3]_pad  & ~n14391 ;
  assign n38788 = n14384 & n38787 ;
  assign n38789 = \m1_data_i[3]_pad  & ~n14391 ;
  assign n38790 = n14399 & n38789 ;
  assign n38791 = ~n38788 & ~n38790 ;
  assign n38792 = \m0_data_i[3]_pad  & n14391 ;
  assign n38793 = n14399 & n38792 ;
  assign n38794 = \m7_data_i[3]_pad  & ~n14391 ;
  assign n38795 = n14408 & n38794 ;
  assign n38796 = ~n38793 & ~n38795 ;
  assign n38797 = n38791 & n38796 ;
  assign n38798 = n38786 & n38797 ;
  assign n38799 = \m3_data_i[4]_pad  & ~n14391 ;
  assign n38800 = n14416 & n38799 ;
  assign n38801 = \m4_data_i[4]_pad  & n14391 ;
  assign n38802 = n14384 & n38801 ;
  assign n38803 = ~n38800 & ~n38802 ;
  assign n38804 = \m6_data_i[4]_pad  & n14391 ;
  assign n38805 = n14408 & n38804 ;
  assign n38806 = \m2_data_i[4]_pad  & n14391 ;
  assign n38807 = n14416 & n38806 ;
  assign n38808 = ~n38805 & ~n38807 ;
  assign n38809 = n38803 & n38808 ;
  assign n38810 = \m5_data_i[4]_pad  & ~n14391 ;
  assign n38811 = n14384 & n38810 ;
  assign n38812 = \m1_data_i[4]_pad  & ~n14391 ;
  assign n38813 = n14399 & n38812 ;
  assign n38814 = ~n38811 & ~n38813 ;
  assign n38815 = \m0_data_i[4]_pad  & n14391 ;
  assign n38816 = n14399 & n38815 ;
  assign n38817 = \m7_data_i[4]_pad  & ~n14391 ;
  assign n38818 = n14408 & n38817 ;
  assign n38819 = ~n38816 & ~n38818 ;
  assign n38820 = n38814 & n38819 ;
  assign n38821 = n38809 & n38820 ;
  assign n38822 = \m3_data_i[5]_pad  & ~n14391 ;
  assign n38823 = n14416 & n38822 ;
  assign n38824 = \m4_data_i[5]_pad  & n14391 ;
  assign n38825 = n14384 & n38824 ;
  assign n38826 = ~n38823 & ~n38825 ;
  assign n38827 = \m6_data_i[5]_pad  & n14391 ;
  assign n38828 = n14408 & n38827 ;
  assign n38829 = \m2_data_i[5]_pad  & n14391 ;
  assign n38830 = n14416 & n38829 ;
  assign n38831 = ~n38828 & ~n38830 ;
  assign n38832 = n38826 & n38831 ;
  assign n38833 = \m5_data_i[5]_pad  & ~n14391 ;
  assign n38834 = n14384 & n38833 ;
  assign n38835 = \m1_data_i[5]_pad  & ~n14391 ;
  assign n38836 = n14399 & n38835 ;
  assign n38837 = ~n38834 & ~n38836 ;
  assign n38838 = \m0_data_i[5]_pad  & n14391 ;
  assign n38839 = n14399 & n38838 ;
  assign n38840 = \m7_data_i[5]_pad  & ~n14391 ;
  assign n38841 = n14408 & n38840 ;
  assign n38842 = ~n38839 & ~n38841 ;
  assign n38843 = n38837 & n38842 ;
  assign n38844 = n38832 & n38843 ;
  assign n38845 = \m3_data_i[6]_pad  & ~n14391 ;
  assign n38846 = n14416 & n38845 ;
  assign n38847 = \m4_data_i[6]_pad  & n14391 ;
  assign n38848 = n14384 & n38847 ;
  assign n38849 = ~n38846 & ~n38848 ;
  assign n38850 = \m6_data_i[6]_pad  & n14391 ;
  assign n38851 = n14408 & n38850 ;
  assign n38852 = \m2_data_i[6]_pad  & n14391 ;
  assign n38853 = n14416 & n38852 ;
  assign n38854 = ~n38851 & ~n38853 ;
  assign n38855 = n38849 & n38854 ;
  assign n38856 = \m5_data_i[6]_pad  & ~n14391 ;
  assign n38857 = n14384 & n38856 ;
  assign n38858 = \m1_data_i[6]_pad  & ~n14391 ;
  assign n38859 = n14399 & n38858 ;
  assign n38860 = ~n38857 & ~n38859 ;
  assign n38861 = \m0_data_i[6]_pad  & n14391 ;
  assign n38862 = n14399 & n38861 ;
  assign n38863 = \m7_data_i[6]_pad  & ~n14391 ;
  assign n38864 = n14408 & n38863 ;
  assign n38865 = ~n38862 & ~n38864 ;
  assign n38866 = n38860 & n38865 ;
  assign n38867 = n38855 & n38866 ;
  assign n38868 = \m3_data_i[7]_pad  & ~n14391 ;
  assign n38869 = n14416 & n38868 ;
  assign n38870 = \m4_data_i[7]_pad  & n14391 ;
  assign n38871 = n14384 & n38870 ;
  assign n38872 = ~n38869 & ~n38871 ;
  assign n38873 = \m6_data_i[7]_pad  & n14391 ;
  assign n38874 = n14408 & n38873 ;
  assign n38875 = \m2_data_i[7]_pad  & n14391 ;
  assign n38876 = n14416 & n38875 ;
  assign n38877 = ~n38874 & ~n38876 ;
  assign n38878 = n38872 & n38877 ;
  assign n38879 = \m5_data_i[7]_pad  & ~n14391 ;
  assign n38880 = n14384 & n38879 ;
  assign n38881 = \m1_data_i[7]_pad  & ~n14391 ;
  assign n38882 = n14399 & n38881 ;
  assign n38883 = ~n38880 & ~n38882 ;
  assign n38884 = \m0_data_i[7]_pad  & n14391 ;
  assign n38885 = n14399 & n38884 ;
  assign n38886 = \m7_data_i[7]_pad  & ~n14391 ;
  assign n38887 = n14408 & n38886 ;
  assign n38888 = ~n38885 & ~n38887 ;
  assign n38889 = n38883 & n38888 ;
  assign n38890 = n38878 & n38889 ;
  assign n38891 = \m3_data_i[8]_pad  & ~n14391 ;
  assign n38892 = n14416 & n38891 ;
  assign n38893 = \m4_data_i[8]_pad  & n14391 ;
  assign n38894 = n14384 & n38893 ;
  assign n38895 = ~n38892 & ~n38894 ;
  assign n38896 = \m6_data_i[8]_pad  & n14391 ;
  assign n38897 = n14408 & n38896 ;
  assign n38898 = \m2_data_i[8]_pad  & n14391 ;
  assign n38899 = n14416 & n38898 ;
  assign n38900 = ~n38897 & ~n38899 ;
  assign n38901 = n38895 & n38900 ;
  assign n38902 = \m5_data_i[8]_pad  & ~n14391 ;
  assign n38903 = n14384 & n38902 ;
  assign n38904 = \m1_data_i[8]_pad  & ~n14391 ;
  assign n38905 = n14399 & n38904 ;
  assign n38906 = ~n38903 & ~n38905 ;
  assign n38907 = \m0_data_i[8]_pad  & n14391 ;
  assign n38908 = n14399 & n38907 ;
  assign n38909 = \m7_data_i[8]_pad  & ~n14391 ;
  assign n38910 = n14408 & n38909 ;
  assign n38911 = ~n38908 & ~n38910 ;
  assign n38912 = n38906 & n38911 ;
  assign n38913 = n38901 & n38912 ;
  assign n38914 = \m3_data_i[9]_pad  & ~n14391 ;
  assign n38915 = n14416 & n38914 ;
  assign n38916 = \m4_data_i[9]_pad  & n14391 ;
  assign n38917 = n14384 & n38916 ;
  assign n38918 = ~n38915 & ~n38917 ;
  assign n38919 = \m6_data_i[9]_pad  & n14391 ;
  assign n38920 = n14408 & n38919 ;
  assign n38921 = \m2_data_i[9]_pad  & n14391 ;
  assign n38922 = n14416 & n38921 ;
  assign n38923 = ~n38920 & ~n38922 ;
  assign n38924 = n38918 & n38923 ;
  assign n38925 = \m5_data_i[9]_pad  & ~n14391 ;
  assign n38926 = n14384 & n38925 ;
  assign n38927 = \m1_data_i[9]_pad  & ~n14391 ;
  assign n38928 = n14399 & n38927 ;
  assign n38929 = ~n38926 & ~n38928 ;
  assign n38930 = \m0_data_i[9]_pad  & n14391 ;
  assign n38931 = n14399 & n38930 ;
  assign n38932 = \m7_data_i[9]_pad  & ~n14391 ;
  assign n38933 = n14408 & n38932 ;
  assign n38934 = ~n38931 & ~n38933 ;
  assign n38935 = n38929 & n38934 ;
  assign n38936 = n38924 & n38935 ;
  assign n38937 = \m3_sel_i[0]_pad  & ~n14391 ;
  assign n38938 = n14416 & n38937 ;
  assign n38939 = \m4_sel_i[0]_pad  & n14391 ;
  assign n38940 = n14384 & n38939 ;
  assign n38941 = ~n38938 & ~n38940 ;
  assign n38942 = \m6_sel_i[0]_pad  & n14391 ;
  assign n38943 = n14408 & n38942 ;
  assign n38944 = \m2_sel_i[0]_pad  & n14391 ;
  assign n38945 = n14416 & n38944 ;
  assign n38946 = ~n38943 & ~n38945 ;
  assign n38947 = n38941 & n38946 ;
  assign n38948 = \m5_sel_i[0]_pad  & ~n14391 ;
  assign n38949 = n14384 & n38948 ;
  assign n38950 = \m1_sel_i[0]_pad  & ~n14391 ;
  assign n38951 = n14399 & n38950 ;
  assign n38952 = ~n38949 & ~n38951 ;
  assign n38953 = \m0_sel_i[0]_pad  & n14391 ;
  assign n38954 = n14399 & n38953 ;
  assign n38955 = \m7_sel_i[0]_pad  & ~n14391 ;
  assign n38956 = n14408 & n38955 ;
  assign n38957 = ~n38954 & ~n38956 ;
  assign n38958 = n38952 & n38957 ;
  assign n38959 = n38947 & n38958 ;
  assign n38960 = \m3_sel_i[1]_pad  & ~n14391 ;
  assign n38961 = n14416 & n38960 ;
  assign n38962 = \m4_sel_i[1]_pad  & n14391 ;
  assign n38963 = n14384 & n38962 ;
  assign n38964 = ~n38961 & ~n38963 ;
  assign n38965 = \m6_sel_i[1]_pad  & n14391 ;
  assign n38966 = n14408 & n38965 ;
  assign n38967 = \m2_sel_i[1]_pad  & n14391 ;
  assign n38968 = n14416 & n38967 ;
  assign n38969 = ~n38966 & ~n38968 ;
  assign n38970 = n38964 & n38969 ;
  assign n38971 = \m5_sel_i[1]_pad  & ~n14391 ;
  assign n38972 = n14384 & n38971 ;
  assign n38973 = \m1_sel_i[1]_pad  & ~n14391 ;
  assign n38974 = n14399 & n38973 ;
  assign n38975 = ~n38972 & ~n38974 ;
  assign n38976 = \m0_sel_i[1]_pad  & n14391 ;
  assign n38977 = n14399 & n38976 ;
  assign n38978 = \m7_sel_i[1]_pad  & ~n14391 ;
  assign n38979 = n14408 & n38978 ;
  assign n38980 = ~n38977 & ~n38979 ;
  assign n38981 = n38975 & n38980 ;
  assign n38982 = n38970 & n38981 ;
  assign n38983 = \m3_sel_i[2]_pad  & ~n14391 ;
  assign n38984 = n14416 & n38983 ;
  assign n38985 = \m4_sel_i[2]_pad  & n14391 ;
  assign n38986 = n14384 & n38985 ;
  assign n38987 = ~n38984 & ~n38986 ;
  assign n38988 = \m6_sel_i[2]_pad  & n14391 ;
  assign n38989 = n14408 & n38988 ;
  assign n38990 = \m2_sel_i[2]_pad  & n14391 ;
  assign n38991 = n14416 & n38990 ;
  assign n38992 = ~n38989 & ~n38991 ;
  assign n38993 = n38987 & n38992 ;
  assign n38994 = \m5_sel_i[2]_pad  & ~n14391 ;
  assign n38995 = n14384 & n38994 ;
  assign n38996 = \m1_sel_i[2]_pad  & ~n14391 ;
  assign n38997 = n14399 & n38996 ;
  assign n38998 = ~n38995 & ~n38997 ;
  assign n38999 = \m0_sel_i[2]_pad  & n14391 ;
  assign n39000 = n14399 & n38999 ;
  assign n39001 = \m7_sel_i[2]_pad  & ~n14391 ;
  assign n39002 = n14408 & n39001 ;
  assign n39003 = ~n39000 & ~n39002 ;
  assign n39004 = n38998 & n39003 ;
  assign n39005 = n38993 & n39004 ;
  assign n39006 = \m3_sel_i[3]_pad  & ~n14391 ;
  assign n39007 = n14416 & n39006 ;
  assign n39008 = \m4_sel_i[3]_pad  & n14391 ;
  assign n39009 = n14384 & n39008 ;
  assign n39010 = ~n39007 & ~n39009 ;
  assign n39011 = \m6_sel_i[3]_pad  & n14391 ;
  assign n39012 = n14408 & n39011 ;
  assign n39013 = \m2_sel_i[3]_pad  & n14391 ;
  assign n39014 = n14416 & n39013 ;
  assign n39015 = ~n39012 & ~n39014 ;
  assign n39016 = n39010 & n39015 ;
  assign n39017 = \m5_sel_i[3]_pad  & ~n14391 ;
  assign n39018 = n14384 & n39017 ;
  assign n39019 = \m1_sel_i[3]_pad  & ~n14391 ;
  assign n39020 = n14399 & n39019 ;
  assign n39021 = ~n39018 & ~n39020 ;
  assign n39022 = \m0_sel_i[3]_pad  & n14391 ;
  assign n39023 = n14399 & n39022 ;
  assign n39024 = \m7_sel_i[3]_pad  & ~n14391 ;
  assign n39025 = n14408 & n39024 ;
  assign n39026 = ~n39023 & ~n39025 ;
  assign n39027 = n39021 & n39026 ;
  assign n39028 = n39016 & n39027 ;
  assign n39029 = \m5_stb_i_pad  & n14975 ;
  assign n39030 = ~n14391 & n39029 ;
  assign n39031 = n14384 & n39030 ;
  assign n39032 = \m4_stb_i_pad  & n14946 ;
  assign n39033 = n14391 & n39032 ;
  assign n39034 = n14384 & n39033 ;
  assign n39035 = ~n39031 & ~n39034 ;
  assign n39036 = \m2_stb_i_pad  & n14866 ;
  assign n39037 = n14391 & n39036 ;
  assign n39038 = n14416 & n39037 ;
  assign n39039 = \m1_stb_i_pad  & n14816 ;
  assign n39040 = ~n14391 & n39039 ;
  assign n39041 = n14399 & n39040 ;
  assign n39042 = ~n39038 & ~n39041 ;
  assign n39043 = n39035 & n39042 ;
  assign n39044 = \m3_stb_i_pad  & n14911 ;
  assign n39045 = ~n14391 & n39044 ;
  assign n39046 = n14416 & n39045 ;
  assign n39047 = \m7_stb_i_pad  & n15066 ;
  assign n39048 = ~n14391 & n39047 ;
  assign n39049 = n14408 & n39048 ;
  assign n39050 = ~n39046 & ~n39049 ;
  assign n39051 = \m6_stb_i_pad  & n15022 ;
  assign n39052 = n14391 & n39051 ;
  assign n39053 = n14408 & n39052 ;
  assign n39054 = \m0_stb_i_pad  & n14770 ;
  assign n39055 = n14391 & n39054 ;
  assign n39056 = n14399 & n39055 ;
  assign n39057 = ~n39053 & ~n39056 ;
  assign n39058 = n39050 & n39057 ;
  assign n39059 = n39043 & n39058 ;
  assign n39060 = \m3_we_i_pad  & ~n14391 ;
  assign n39061 = n14416 & n39060 ;
  assign n39062 = \m4_we_i_pad  & n14391 ;
  assign n39063 = n14384 & n39062 ;
  assign n39064 = ~n39061 & ~n39063 ;
  assign n39065 = \m6_we_i_pad  & n14391 ;
  assign n39066 = n14408 & n39065 ;
  assign n39067 = \m2_we_i_pad  & n14391 ;
  assign n39068 = n14416 & n39067 ;
  assign n39069 = ~n39066 & ~n39068 ;
  assign n39070 = n39064 & n39069 ;
  assign n39071 = \m5_we_i_pad  & ~n14391 ;
  assign n39072 = n14384 & n39071 ;
  assign n39073 = \m1_we_i_pad  & ~n14391 ;
  assign n39074 = n14399 & n39073 ;
  assign n39075 = ~n39072 & ~n39074 ;
  assign n39076 = \m0_we_i_pad  & n14391 ;
  assign n39077 = n14399 & n39076 ;
  assign n39078 = \m7_we_i_pad  & ~n14391 ;
  assign n39079 = n14408 & n39078 ;
  assign n39080 = ~n39077 & ~n39079 ;
  assign n39081 = n39075 & n39080 ;
  assign n39082 = n39070 & n39081 ;
  assign n39083 = \m1_addr_i[0]_pad  & ~n14451 ;
  assign n39084 = n14476 & n39083 ;
  assign n39085 = \m2_addr_i[0]_pad  & n14451 ;
  assign n39086 = n14459 & n39085 ;
  assign n39087 = ~n39084 & ~n39086 ;
  assign n39088 = \m6_addr_i[0]_pad  & n14451 ;
  assign n39089 = n14468 & n39088 ;
  assign n39090 = \m7_addr_i[0]_pad  & ~n14451 ;
  assign n39091 = n14468 & n39090 ;
  assign n39092 = ~n39089 & ~n39091 ;
  assign n39093 = n39087 & n39092 ;
  assign n39094 = \m5_addr_i[0]_pad  & ~n14451 ;
  assign n39095 = n14444 & n39094 ;
  assign n39096 = \m0_addr_i[0]_pad  & n14451 ;
  assign n39097 = n14476 & n39096 ;
  assign n39098 = ~n39095 & ~n39097 ;
  assign n39099 = \m3_addr_i[0]_pad  & ~n14451 ;
  assign n39100 = n14459 & n39099 ;
  assign n39101 = \m4_addr_i[0]_pad  & n14451 ;
  assign n39102 = n14444 & n39101 ;
  assign n39103 = ~n39100 & ~n39102 ;
  assign n39104 = n39098 & n39103 ;
  assign n39105 = n39093 & n39104 ;
  assign n39106 = \m3_addr_i[10]_pad  & ~n14451 ;
  assign n39107 = n14459 & n39106 ;
  assign n39108 = \m4_addr_i[10]_pad  & n14451 ;
  assign n39109 = n14444 & n39108 ;
  assign n39110 = ~n39107 & ~n39109 ;
  assign n39111 = \m6_addr_i[10]_pad  & n14451 ;
  assign n39112 = n14468 & n39111 ;
  assign n39113 = \m2_addr_i[10]_pad  & n14451 ;
  assign n39114 = n14459 & n39113 ;
  assign n39115 = ~n39112 & ~n39114 ;
  assign n39116 = n39110 & n39115 ;
  assign n39117 = \m5_addr_i[10]_pad  & ~n14451 ;
  assign n39118 = n14444 & n39117 ;
  assign n39119 = \m1_addr_i[10]_pad  & ~n14451 ;
  assign n39120 = n14476 & n39119 ;
  assign n39121 = ~n39118 & ~n39120 ;
  assign n39122 = \m0_addr_i[10]_pad  & n14451 ;
  assign n39123 = n14476 & n39122 ;
  assign n39124 = \m7_addr_i[10]_pad  & ~n14451 ;
  assign n39125 = n14468 & n39124 ;
  assign n39126 = ~n39123 & ~n39125 ;
  assign n39127 = n39121 & n39126 ;
  assign n39128 = n39116 & n39127 ;
  assign n39129 = \m3_addr_i[11]_pad  & ~n14451 ;
  assign n39130 = n14459 & n39129 ;
  assign n39131 = \m4_addr_i[11]_pad  & n14451 ;
  assign n39132 = n14444 & n39131 ;
  assign n39133 = ~n39130 & ~n39132 ;
  assign n39134 = \m6_addr_i[11]_pad  & n14451 ;
  assign n39135 = n14468 & n39134 ;
  assign n39136 = \m2_addr_i[11]_pad  & n14451 ;
  assign n39137 = n14459 & n39136 ;
  assign n39138 = ~n39135 & ~n39137 ;
  assign n39139 = n39133 & n39138 ;
  assign n39140 = \m5_addr_i[11]_pad  & ~n14451 ;
  assign n39141 = n14444 & n39140 ;
  assign n39142 = \m1_addr_i[11]_pad  & ~n14451 ;
  assign n39143 = n14476 & n39142 ;
  assign n39144 = ~n39141 & ~n39143 ;
  assign n39145 = \m0_addr_i[11]_pad  & n14451 ;
  assign n39146 = n14476 & n39145 ;
  assign n39147 = \m7_addr_i[11]_pad  & ~n14451 ;
  assign n39148 = n14468 & n39147 ;
  assign n39149 = ~n39146 & ~n39148 ;
  assign n39150 = n39144 & n39149 ;
  assign n39151 = n39139 & n39150 ;
  assign n39152 = \m3_addr_i[12]_pad  & ~n14451 ;
  assign n39153 = n14459 & n39152 ;
  assign n39154 = \m4_addr_i[12]_pad  & n14451 ;
  assign n39155 = n14444 & n39154 ;
  assign n39156 = ~n39153 & ~n39155 ;
  assign n39157 = \m6_addr_i[12]_pad  & n14451 ;
  assign n39158 = n14468 & n39157 ;
  assign n39159 = \m2_addr_i[12]_pad  & n14451 ;
  assign n39160 = n14459 & n39159 ;
  assign n39161 = ~n39158 & ~n39160 ;
  assign n39162 = n39156 & n39161 ;
  assign n39163 = \m5_addr_i[12]_pad  & ~n14451 ;
  assign n39164 = n14444 & n39163 ;
  assign n39165 = \m1_addr_i[12]_pad  & ~n14451 ;
  assign n39166 = n14476 & n39165 ;
  assign n39167 = ~n39164 & ~n39166 ;
  assign n39168 = \m0_addr_i[12]_pad  & n14451 ;
  assign n39169 = n14476 & n39168 ;
  assign n39170 = \m7_addr_i[12]_pad  & ~n14451 ;
  assign n39171 = n14468 & n39170 ;
  assign n39172 = ~n39169 & ~n39171 ;
  assign n39173 = n39167 & n39172 ;
  assign n39174 = n39162 & n39173 ;
  assign n39175 = \m3_addr_i[13]_pad  & ~n14451 ;
  assign n39176 = n14459 & n39175 ;
  assign n39177 = \m4_addr_i[13]_pad  & n14451 ;
  assign n39178 = n14444 & n39177 ;
  assign n39179 = ~n39176 & ~n39178 ;
  assign n39180 = \m6_addr_i[13]_pad  & n14451 ;
  assign n39181 = n14468 & n39180 ;
  assign n39182 = \m2_addr_i[13]_pad  & n14451 ;
  assign n39183 = n14459 & n39182 ;
  assign n39184 = ~n39181 & ~n39183 ;
  assign n39185 = n39179 & n39184 ;
  assign n39186 = \m5_addr_i[13]_pad  & ~n14451 ;
  assign n39187 = n14444 & n39186 ;
  assign n39188 = \m1_addr_i[13]_pad  & ~n14451 ;
  assign n39189 = n14476 & n39188 ;
  assign n39190 = ~n39187 & ~n39189 ;
  assign n39191 = \m0_addr_i[13]_pad  & n14451 ;
  assign n39192 = n14476 & n39191 ;
  assign n39193 = \m7_addr_i[13]_pad  & ~n14451 ;
  assign n39194 = n14468 & n39193 ;
  assign n39195 = ~n39192 & ~n39194 ;
  assign n39196 = n39190 & n39195 ;
  assign n39197 = n39185 & n39196 ;
  assign n39198 = \m3_addr_i[14]_pad  & ~n14451 ;
  assign n39199 = n14459 & n39198 ;
  assign n39200 = \m4_addr_i[14]_pad  & n14451 ;
  assign n39201 = n14444 & n39200 ;
  assign n39202 = ~n39199 & ~n39201 ;
  assign n39203 = \m6_addr_i[14]_pad  & n14451 ;
  assign n39204 = n14468 & n39203 ;
  assign n39205 = \m2_addr_i[14]_pad  & n14451 ;
  assign n39206 = n14459 & n39205 ;
  assign n39207 = ~n39204 & ~n39206 ;
  assign n39208 = n39202 & n39207 ;
  assign n39209 = \m5_addr_i[14]_pad  & ~n14451 ;
  assign n39210 = n14444 & n39209 ;
  assign n39211 = \m1_addr_i[14]_pad  & ~n14451 ;
  assign n39212 = n14476 & n39211 ;
  assign n39213 = ~n39210 & ~n39212 ;
  assign n39214 = \m0_addr_i[14]_pad  & n14451 ;
  assign n39215 = n14476 & n39214 ;
  assign n39216 = \m7_addr_i[14]_pad  & ~n14451 ;
  assign n39217 = n14468 & n39216 ;
  assign n39218 = ~n39215 & ~n39217 ;
  assign n39219 = n39213 & n39218 ;
  assign n39220 = n39208 & n39219 ;
  assign n39221 = \m3_addr_i[15]_pad  & ~n14451 ;
  assign n39222 = n14459 & n39221 ;
  assign n39223 = \m4_addr_i[15]_pad  & n14451 ;
  assign n39224 = n14444 & n39223 ;
  assign n39225 = ~n39222 & ~n39224 ;
  assign n39226 = \m6_addr_i[15]_pad  & n14451 ;
  assign n39227 = n14468 & n39226 ;
  assign n39228 = \m2_addr_i[15]_pad  & n14451 ;
  assign n39229 = n14459 & n39228 ;
  assign n39230 = ~n39227 & ~n39229 ;
  assign n39231 = n39225 & n39230 ;
  assign n39232 = \m5_addr_i[15]_pad  & ~n14451 ;
  assign n39233 = n14444 & n39232 ;
  assign n39234 = \m1_addr_i[15]_pad  & ~n14451 ;
  assign n39235 = n14476 & n39234 ;
  assign n39236 = ~n39233 & ~n39235 ;
  assign n39237 = \m0_addr_i[15]_pad  & n14451 ;
  assign n39238 = n14476 & n39237 ;
  assign n39239 = \m7_addr_i[15]_pad  & ~n14451 ;
  assign n39240 = n14468 & n39239 ;
  assign n39241 = ~n39238 & ~n39240 ;
  assign n39242 = n39236 & n39241 ;
  assign n39243 = n39231 & n39242 ;
  assign n39244 = \m3_addr_i[16]_pad  & ~n14451 ;
  assign n39245 = n14459 & n39244 ;
  assign n39246 = \m4_addr_i[16]_pad  & n14451 ;
  assign n39247 = n14444 & n39246 ;
  assign n39248 = ~n39245 & ~n39247 ;
  assign n39249 = \m6_addr_i[16]_pad  & n14451 ;
  assign n39250 = n14468 & n39249 ;
  assign n39251 = \m2_addr_i[16]_pad  & n14451 ;
  assign n39252 = n14459 & n39251 ;
  assign n39253 = ~n39250 & ~n39252 ;
  assign n39254 = n39248 & n39253 ;
  assign n39255 = \m5_addr_i[16]_pad  & ~n14451 ;
  assign n39256 = n14444 & n39255 ;
  assign n39257 = \m1_addr_i[16]_pad  & ~n14451 ;
  assign n39258 = n14476 & n39257 ;
  assign n39259 = ~n39256 & ~n39258 ;
  assign n39260 = \m0_addr_i[16]_pad  & n14451 ;
  assign n39261 = n14476 & n39260 ;
  assign n39262 = \m7_addr_i[16]_pad  & ~n14451 ;
  assign n39263 = n14468 & n39262 ;
  assign n39264 = ~n39261 & ~n39263 ;
  assign n39265 = n39259 & n39264 ;
  assign n39266 = n39254 & n39265 ;
  assign n39267 = \m3_addr_i[17]_pad  & ~n14451 ;
  assign n39268 = n14459 & n39267 ;
  assign n39269 = \m4_addr_i[17]_pad  & n14451 ;
  assign n39270 = n14444 & n39269 ;
  assign n39271 = ~n39268 & ~n39270 ;
  assign n39272 = \m6_addr_i[17]_pad  & n14451 ;
  assign n39273 = n14468 & n39272 ;
  assign n39274 = \m2_addr_i[17]_pad  & n14451 ;
  assign n39275 = n14459 & n39274 ;
  assign n39276 = ~n39273 & ~n39275 ;
  assign n39277 = n39271 & n39276 ;
  assign n39278 = \m5_addr_i[17]_pad  & ~n14451 ;
  assign n39279 = n14444 & n39278 ;
  assign n39280 = \m1_addr_i[17]_pad  & ~n14451 ;
  assign n39281 = n14476 & n39280 ;
  assign n39282 = ~n39279 & ~n39281 ;
  assign n39283 = \m0_addr_i[17]_pad  & n14451 ;
  assign n39284 = n14476 & n39283 ;
  assign n39285 = \m7_addr_i[17]_pad  & ~n14451 ;
  assign n39286 = n14468 & n39285 ;
  assign n39287 = ~n39284 & ~n39286 ;
  assign n39288 = n39282 & n39287 ;
  assign n39289 = n39277 & n39288 ;
  assign n39290 = \m3_addr_i[18]_pad  & ~n14451 ;
  assign n39291 = n14459 & n39290 ;
  assign n39292 = \m4_addr_i[18]_pad  & n14451 ;
  assign n39293 = n14444 & n39292 ;
  assign n39294 = ~n39291 & ~n39293 ;
  assign n39295 = \m6_addr_i[18]_pad  & n14451 ;
  assign n39296 = n14468 & n39295 ;
  assign n39297 = \m2_addr_i[18]_pad  & n14451 ;
  assign n39298 = n14459 & n39297 ;
  assign n39299 = ~n39296 & ~n39298 ;
  assign n39300 = n39294 & n39299 ;
  assign n39301 = \m5_addr_i[18]_pad  & ~n14451 ;
  assign n39302 = n14444 & n39301 ;
  assign n39303 = \m1_addr_i[18]_pad  & ~n14451 ;
  assign n39304 = n14476 & n39303 ;
  assign n39305 = ~n39302 & ~n39304 ;
  assign n39306 = \m0_addr_i[18]_pad  & n14451 ;
  assign n39307 = n14476 & n39306 ;
  assign n39308 = \m7_addr_i[18]_pad  & ~n14451 ;
  assign n39309 = n14468 & n39308 ;
  assign n39310 = ~n39307 & ~n39309 ;
  assign n39311 = n39305 & n39310 ;
  assign n39312 = n39300 & n39311 ;
  assign n39313 = \m3_addr_i[19]_pad  & ~n14451 ;
  assign n39314 = n14459 & n39313 ;
  assign n39315 = \m4_addr_i[19]_pad  & n14451 ;
  assign n39316 = n14444 & n39315 ;
  assign n39317 = ~n39314 & ~n39316 ;
  assign n39318 = \m6_addr_i[19]_pad  & n14451 ;
  assign n39319 = n14468 & n39318 ;
  assign n39320 = \m2_addr_i[19]_pad  & n14451 ;
  assign n39321 = n14459 & n39320 ;
  assign n39322 = ~n39319 & ~n39321 ;
  assign n39323 = n39317 & n39322 ;
  assign n39324 = \m5_addr_i[19]_pad  & ~n14451 ;
  assign n39325 = n14444 & n39324 ;
  assign n39326 = \m1_addr_i[19]_pad  & ~n14451 ;
  assign n39327 = n14476 & n39326 ;
  assign n39328 = ~n39325 & ~n39327 ;
  assign n39329 = \m0_addr_i[19]_pad  & n14451 ;
  assign n39330 = n14476 & n39329 ;
  assign n39331 = \m7_addr_i[19]_pad  & ~n14451 ;
  assign n39332 = n14468 & n39331 ;
  assign n39333 = ~n39330 & ~n39332 ;
  assign n39334 = n39328 & n39333 ;
  assign n39335 = n39323 & n39334 ;
  assign n39336 = \m3_addr_i[1]_pad  & ~n14451 ;
  assign n39337 = n14459 & n39336 ;
  assign n39338 = \m4_addr_i[1]_pad  & n14451 ;
  assign n39339 = n14444 & n39338 ;
  assign n39340 = ~n39337 & ~n39339 ;
  assign n39341 = \m6_addr_i[1]_pad  & n14451 ;
  assign n39342 = n14468 & n39341 ;
  assign n39343 = \m2_addr_i[1]_pad  & n14451 ;
  assign n39344 = n14459 & n39343 ;
  assign n39345 = ~n39342 & ~n39344 ;
  assign n39346 = n39340 & n39345 ;
  assign n39347 = \m5_addr_i[1]_pad  & ~n14451 ;
  assign n39348 = n14444 & n39347 ;
  assign n39349 = \m1_addr_i[1]_pad  & ~n14451 ;
  assign n39350 = n14476 & n39349 ;
  assign n39351 = ~n39348 & ~n39350 ;
  assign n39352 = \m0_addr_i[1]_pad  & n14451 ;
  assign n39353 = n14476 & n39352 ;
  assign n39354 = \m7_addr_i[1]_pad  & ~n14451 ;
  assign n39355 = n14468 & n39354 ;
  assign n39356 = ~n39353 & ~n39355 ;
  assign n39357 = n39351 & n39356 ;
  assign n39358 = n39346 & n39357 ;
  assign n39359 = \m3_addr_i[20]_pad  & ~n14451 ;
  assign n39360 = n14459 & n39359 ;
  assign n39361 = \m4_addr_i[20]_pad  & n14451 ;
  assign n39362 = n14444 & n39361 ;
  assign n39363 = ~n39360 & ~n39362 ;
  assign n39364 = \m6_addr_i[20]_pad  & n14451 ;
  assign n39365 = n14468 & n39364 ;
  assign n39366 = \m2_addr_i[20]_pad  & n14451 ;
  assign n39367 = n14459 & n39366 ;
  assign n39368 = ~n39365 & ~n39367 ;
  assign n39369 = n39363 & n39368 ;
  assign n39370 = \m5_addr_i[20]_pad  & ~n14451 ;
  assign n39371 = n14444 & n39370 ;
  assign n39372 = \m1_addr_i[20]_pad  & ~n14451 ;
  assign n39373 = n14476 & n39372 ;
  assign n39374 = ~n39371 & ~n39373 ;
  assign n39375 = \m0_addr_i[20]_pad  & n14451 ;
  assign n39376 = n14476 & n39375 ;
  assign n39377 = \m7_addr_i[20]_pad  & ~n14451 ;
  assign n39378 = n14468 & n39377 ;
  assign n39379 = ~n39376 & ~n39378 ;
  assign n39380 = n39374 & n39379 ;
  assign n39381 = n39369 & n39380 ;
  assign n39382 = \m3_addr_i[21]_pad  & ~n14451 ;
  assign n39383 = n14459 & n39382 ;
  assign n39384 = \m4_addr_i[21]_pad  & n14451 ;
  assign n39385 = n14444 & n39384 ;
  assign n39386 = ~n39383 & ~n39385 ;
  assign n39387 = \m6_addr_i[21]_pad  & n14451 ;
  assign n39388 = n14468 & n39387 ;
  assign n39389 = \m2_addr_i[21]_pad  & n14451 ;
  assign n39390 = n14459 & n39389 ;
  assign n39391 = ~n39388 & ~n39390 ;
  assign n39392 = n39386 & n39391 ;
  assign n39393 = \m5_addr_i[21]_pad  & ~n14451 ;
  assign n39394 = n14444 & n39393 ;
  assign n39395 = \m1_addr_i[21]_pad  & ~n14451 ;
  assign n39396 = n14476 & n39395 ;
  assign n39397 = ~n39394 & ~n39396 ;
  assign n39398 = \m0_addr_i[21]_pad  & n14451 ;
  assign n39399 = n14476 & n39398 ;
  assign n39400 = \m7_addr_i[21]_pad  & ~n14451 ;
  assign n39401 = n14468 & n39400 ;
  assign n39402 = ~n39399 & ~n39401 ;
  assign n39403 = n39397 & n39402 ;
  assign n39404 = n39392 & n39403 ;
  assign n39405 = \m3_addr_i[22]_pad  & ~n14451 ;
  assign n39406 = n14459 & n39405 ;
  assign n39407 = \m4_addr_i[22]_pad  & n14451 ;
  assign n39408 = n14444 & n39407 ;
  assign n39409 = ~n39406 & ~n39408 ;
  assign n39410 = \m6_addr_i[22]_pad  & n14451 ;
  assign n39411 = n14468 & n39410 ;
  assign n39412 = \m2_addr_i[22]_pad  & n14451 ;
  assign n39413 = n14459 & n39412 ;
  assign n39414 = ~n39411 & ~n39413 ;
  assign n39415 = n39409 & n39414 ;
  assign n39416 = \m5_addr_i[22]_pad  & ~n14451 ;
  assign n39417 = n14444 & n39416 ;
  assign n39418 = \m1_addr_i[22]_pad  & ~n14451 ;
  assign n39419 = n14476 & n39418 ;
  assign n39420 = ~n39417 & ~n39419 ;
  assign n39421 = \m0_addr_i[22]_pad  & n14451 ;
  assign n39422 = n14476 & n39421 ;
  assign n39423 = \m7_addr_i[22]_pad  & ~n14451 ;
  assign n39424 = n14468 & n39423 ;
  assign n39425 = ~n39422 & ~n39424 ;
  assign n39426 = n39420 & n39425 ;
  assign n39427 = n39415 & n39426 ;
  assign n39428 = \m3_addr_i[23]_pad  & ~n14451 ;
  assign n39429 = n14459 & n39428 ;
  assign n39430 = \m4_addr_i[23]_pad  & n14451 ;
  assign n39431 = n14444 & n39430 ;
  assign n39432 = ~n39429 & ~n39431 ;
  assign n39433 = \m6_addr_i[23]_pad  & n14451 ;
  assign n39434 = n14468 & n39433 ;
  assign n39435 = \m2_addr_i[23]_pad  & n14451 ;
  assign n39436 = n14459 & n39435 ;
  assign n39437 = ~n39434 & ~n39436 ;
  assign n39438 = n39432 & n39437 ;
  assign n39439 = \m5_addr_i[23]_pad  & ~n14451 ;
  assign n39440 = n14444 & n39439 ;
  assign n39441 = \m1_addr_i[23]_pad  & ~n14451 ;
  assign n39442 = n14476 & n39441 ;
  assign n39443 = ~n39440 & ~n39442 ;
  assign n39444 = \m0_addr_i[23]_pad  & n14451 ;
  assign n39445 = n14476 & n39444 ;
  assign n39446 = \m7_addr_i[23]_pad  & ~n14451 ;
  assign n39447 = n14468 & n39446 ;
  assign n39448 = ~n39445 & ~n39447 ;
  assign n39449 = n39443 & n39448 ;
  assign n39450 = n39438 & n39449 ;
  assign n39451 = \m3_addr_i[24]_pad  & ~n14451 ;
  assign n39452 = n14459 & n39451 ;
  assign n39453 = \m4_addr_i[24]_pad  & n14451 ;
  assign n39454 = n14444 & n39453 ;
  assign n39455 = ~n39452 & ~n39454 ;
  assign n39456 = \m5_addr_i[24]_pad  & ~n14451 ;
  assign n39457 = n14444 & n39456 ;
  assign n39458 = \m2_addr_i[24]_pad  & n14451 ;
  assign n39459 = n14459 & n39458 ;
  assign n39460 = ~n39457 & ~n39459 ;
  assign n39461 = n39455 & n39460 ;
  assign n39462 = \m6_addr_i[24]_pad  & n14451 ;
  assign n39463 = n14468 & n39462 ;
  assign n39464 = \m1_addr_i[24]_pad  & ~n14451 ;
  assign n39465 = n14476 & n39464 ;
  assign n39466 = ~n39463 & ~n39465 ;
  assign n39467 = \m0_addr_i[24]_pad  & n14451 ;
  assign n39468 = n14476 & n39467 ;
  assign n39469 = \m7_addr_i[24]_pad  & ~n14451 ;
  assign n39470 = n14468 & n39469 ;
  assign n39471 = ~n39468 & ~n39470 ;
  assign n39472 = n39466 & n39471 ;
  assign n39473 = n39461 & n39472 ;
  assign n39474 = \m3_addr_i[25]_pad  & ~n14451 ;
  assign n39475 = n14459 & n39474 ;
  assign n39476 = \m4_addr_i[25]_pad  & n14451 ;
  assign n39477 = n14444 & n39476 ;
  assign n39478 = ~n39475 & ~n39477 ;
  assign n39479 = \m5_addr_i[25]_pad  & ~n14451 ;
  assign n39480 = n14444 & n39479 ;
  assign n39481 = \m2_addr_i[25]_pad  & n14451 ;
  assign n39482 = n14459 & n39481 ;
  assign n39483 = ~n39480 & ~n39482 ;
  assign n39484 = n39478 & n39483 ;
  assign n39485 = \m6_addr_i[25]_pad  & n14451 ;
  assign n39486 = n14468 & n39485 ;
  assign n39487 = \m1_addr_i[25]_pad  & ~n14451 ;
  assign n39488 = n14476 & n39487 ;
  assign n39489 = ~n39486 & ~n39488 ;
  assign n39490 = \m0_addr_i[25]_pad  & n14451 ;
  assign n39491 = n14476 & n39490 ;
  assign n39492 = \m7_addr_i[25]_pad  & ~n14451 ;
  assign n39493 = n14468 & n39492 ;
  assign n39494 = ~n39491 & ~n39493 ;
  assign n39495 = n39489 & n39494 ;
  assign n39496 = n39484 & n39495 ;
  assign n39497 = \m3_addr_i[26]_pad  & ~n14451 ;
  assign n39498 = n14459 & n39497 ;
  assign n39499 = \m4_addr_i[26]_pad  & n14451 ;
  assign n39500 = n14444 & n39499 ;
  assign n39501 = ~n39498 & ~n39500 ;
  assign n39502 = \m5_addr_i[26]_pad  & ~n14451 ;
  assign n39503 = n14444 & n39502 ;
  assign n39504 = \m2_addr_i[26]_pad  & n14451 ;
  assign n39505 = n14459 & n39504 ;
  assign n39506 = ~n39503 & ~n39505 ;
  assign n39507 = n39501 & n39506 ;
  assign n39508 = \m6_addr_i[26]_pad  & n14451 ;
  assign n39509 = n14468 & n39508 ;
  assign n39510 = \m1_addr_i[26]_pad  & ~n14451 ;
  assign n39511 = n14476 & n39510 ;
  assign n39512 = ~n39509 & ~n39511 ;
  assign n39513 = \m0_addr_i[26]_pad  & n14451 ;
  assign n39514 = n14476 & n39513 ;
  assign n39515 = \m7_addr_i[26]_pad  & ~n14451 ;
  assign n39516 = n14468 & n39515 ;
  assign n39517 = ~n39514 & ~n39516 ;
  assign n39518 = n39512 & n39517 ;
  assign n39519 = n39507 & n39518 ;
  assign n39520 = \m3_addr_i[27]_pad  & ~n14451 ;
  assign n39521 = n14459 & n39520 ;
  assign n39522 = \m4_addr_i[27]_pad  & n14451 ;
  assign n39523 = n14444 & n39522 ;
  assign n39524 = ~n39521 & ~n39523 ;
  assign n39525 = \m5_addr_i[27]_pad  & ~n14451 ;
  assign n39526 = n14444 & n39525 ;
  assign n39527 = \m2_addr_i[27]_pad  & n14451 ;
  assign n39528 = n14459 & n39527 ;
  assign n39529 = ~n39526 & ~n39528 ;
  assign n39530 = n39524 & n39529 ;
  assign n39531 = \m6_addr_i[27]_pad  & n14451 ;
  assign n39532 = n14468 & n39531 ;
  assign n39533 = \m1_addr_i[27]_pad  & ~n14451 ;
  assign n39534 = n14476 & n39533 ;
  assign n39535 = ~n39532 & ~n39534 ;
  assign n39536 = \m0_addr_i[27]_pad  & n14451 ;
  assign n39537 = n14476 & n39536 ;
  assign n39538 = \m7_addr_i[27]_pad  & ~n14451 ;
  assign n39539 = n14468 & n39538 ;
  assign n39540 = ~n39537 & ~n39539 ;
  assign n39541 = n39535 & n39540 ;
  assign n39542 = n39530 & n39541 ;
  assign n39543 = \m3_addr_i[28]_pad  & ~n14451 ;
  assign n39544 = n14459 & n39543 ;
  assign n39545 = \m4_addr_i[28]_pad  & n14451 ;
  assign n39546 = n14444 & n39545 ;
  assign n39547 = ~n39544 & ~n39546 ;
  assign n39548 = \m5_addr_i[28]_pad  & ~n14451 ;
  assign n39549 = n14444 & n39548 ;
  assign n39550 = \m2_addr_i[28]_pad  & n14451 ;
  assign n39551 = n14459 & n39550 ;
  assign n39552 = ~n39549 & ~n39551 ;
  assign n39553 = n39547 & n39552 ;
  assign n39554 = \m6_addr_i[28]_pad  & n14451 ;
  assign n39555 = n14468 & n39554 ;
  assign n39556 = \m1_addr_i[28]_pad  & ~n14451 ;
  assign n39557 = n14476 & n39556 ;
  assign n39558 = ~n39555 & ~n39557 ;
  assign n39559 = \m0_addr_i[28]_pad  & n14451 ;
  assign n39560 = n14476 & n39559 ;
  assign n39561 = \m7_addr_i[28]_pad  & ~n14451 ;
  assign n39562 = n14468 & n39561 ;
  assign n39563 = ~n39560 & ~n39562 ;
  assign n39564 = n39558 & n39563 ;
  assign n39565 = n39553 & n39564 ;
  assign n39566 = \m3_addr_i[29]_pad  & ~n14451 ;
  assign n39567 = n14459 & n39566 ;
  assign n39568 = \m4_addr_i[29]_pad  & n14451 ;
  assign n39569 = n14444 & n39568 ;
  assign n39570 = ~n39567 & ~n39569 ;
  assign n39571 = \m5_addr_i[29]_pad  & ~n14451 ;
  assign n39572 = n14444 & n39571 ;
  assign n39573 = \m2_addr_i[29]_pad  & n14451 ;
  assign n39574 = n14459 & n39573 ;
  assign n39575 = ~n39572 & ~n39574 ;
  assign n39576 = n39570 & n39575 ;
  assign n39577 = \m6_addr_i[29]_pad  & n14451 ;
  assign n39578 = n14468 & n39577 ;
  assign n39579 = \m1_addr_i[29]_pad  & ~n14451 ;
  assign n39580 = n14476 & n39579 ;
  assign n39581 = ~n39578 & ~n39580 ;
  assign n39582 = \m0_addr_i[29]_pad  & n14451 ;
  assign n39583 = n14476 & n39582 ;
  assign n39584 = \m7_addr_i[29]_pad  & ~n14451 ;
  assign n39585 = n14468 & n39584 ;
  assign n39586 = ~n39583 & ~n39585 ;
  assign n39587 = n39581 & n39586 ;
  assign n39588 = n39576 & n39587 ;
  assign n39589 = \m3_addr_i[2]_pad  & ~n14451 ;
  assign n39590 = n14459 & n39589 ;
  assign n39591 = \m4_addr_i[2]_pad  & n14451 ;
  assign n39592 = n14444 & n39591 ;
  assign n39593 = ~n39590 & ~n39592 ;
  assign n39594 = \m6_addr_i[2]_pad  & n14451 ;
  assign n39595 = n14468 & n39594 ;
  assign n39596 = \m2_addr_i[2]_pad  & n14451 ;
  assign n39597 = n14459 & n39596 ;
  assign n39598 = ~n39595 & ~n39597 ;
  assign n39599 = n39593 & n39598 ;
  assign n39600 = \m5_addr_i[2]_pad  & ~n14451 ;
  assign n39601 = n14444 & n39600 ;
  assign n39602 = \m1_addr_i[2]_pad  & ~n14451 ;
  assign n39603 = n14476 & n39602 ;
  assign n39604 = ~n39601 & ~n39603 ;
  assign n39605 = \m0_addr_i[2]_pad  & n14451 ;
  assign n39606 = n14476 & n39605 ;
  assign n39607 = \m7_addr_i[2]_pad  & ~n14451 ;
  assign n39608 = n14468 & n39607 ;
  assign n39609 = ~n39606 & ~n39608 ;
  assign n39610 = n39604 & n39609 ;
  assign n39611 = n39599 & n39610 ;
  assign n39612 = \m3_addr_i[30]_pad  & ~n14451 ;
  assign n39613 = n14459 & n39612 ;
  assign n39614 = \m4_addr_i[30]_pad  & n14451 ;
  assign n39615 = n14444 & n39614 ;
  assign n39616 = ~n39613 & ~n39615 ;
  assign n39617 = \m5_addr_i[30]_pad  & ~n14451 ;
  assign n39618 = n14444 & n39617 ;
  assign n39619 = \m2_addr_i[30]_pad  & n14451 ;
  assign n39620 = n14459 & n39619 ;
  assign n39621 = ~n39618 & ~n39620 ;
  assign n39622 = n39616 & n39621 ;
  assign n39623 = \m6_addr_i[30]_pad  & n14451 ;
  assign n39624 = n14468 & n39623 ;
  assign n39625 = \m1_addr_i[30]_pad  & ~n14451 ;
  assign n39626 = n14476 & n39625 ;
  assign n39627 = ~n39624 & ~n39626 ;
  assign n39628 = \m0_addr_i[30]_pad  & n14451 ;
  assign n39629 = n14476 & n39628 ;
  assign n39630 = \m7_addr_i[30]_pad  & ~n14451 ;
  assign n39631 = n14468 & n39630 ;
  assign n39632 = ~n39629 & ~n39631 ;
  assign n39633 = n39627 & n39632 ;
  assign n39634 = n39622 & n39633 ;
  assign n39635 = \m3_addr_i[31]_pad  & ~n14451 ;
  assign n39636 = n14459 & n39635 ;
  assign n39637 = \m4_addr_i[31]_pad  & n14451 ;
  assign n39638 = n14444 & n39637 ;
  assign n39639 = ~n39636 & ~n39638 ;
  assign n39640 = \m5_addr_i[31]_pad  & ~n14451 ;
  assign n39641 = n14444 & n39640 ;
  assign n39642 = \m2_addr_i[31]_pad  & n14451 ;
  assign n39643 = n14459 & n39642 ;
  assign n39644 = ~n39641 & ~n39643 ;
  assign n39645 = n39639 & n39644 ;
  assign n39646 = \m6_addr_i[31]_pad  & n14451 ;
  assign n39647 = n14468 & n39646 ;
  assign n39648 = \m1_addr_i[31]_pad  & ~n14451 ;
  assign n39649 = n14476 & n39648 ;
  assign n39650 = ~n39647 & ~n39649 ;
  assign n39651 = \m0_addr_i[31]_pad  & n14451 ;
  assign n39652 = n14476 & n39651 ;
  assign n39653 = \m7_addr_i[31]_pad  & ~n14451 ;
  assign n39654 = n14468 & n39653 ;
  assign n39655 = ~n39652 & ~n39654 ;
  assign n39656 = n39650 & n39655 ;
  assign n39657 = n39645 & n39656 ;
  assign n39658 = \m3_addr_i[3]_pad  & ~n14451 ;
  assign n39659 = n14459 & n39658 ;
  assign n39660 = \m4_addr_i[3]_pad  & n14451 ;
  assign n39661 = n14444 & n39660 ;
  assign n39662 = ~n39659 & ~n39661 ;
  assign n39663 = \m6_addr_i[3]_pad  & n14451 ;
  assign n39664 = n14468 & n39663 ;
  assign n39665 = \m2_addr_i[3]_pad  & n14451 ;
  assign n39666 = n14459 & n39665 ;
  assign n39667 = ~n39664 & ~n39666 ;
  assign n39668 = n39662 & n39667 ;
  assign n39669 = \m5_addr_i[3]_pad  & ~n14451 ;
  assign n39670 = n14444 & n39669 ;
  assign n39671 = \m1_addr_i[3]_pad  & ~n14451 ;
  assign n39672 = n14476 & n39671 ;
  assign n39673 = ~n39670 & ~n39672 ;
  assign n39674 = \m0_addr_i[3]_pad  & n14451 ;
  assign n39675 = n14476 & n39674 ;
  assign n39676 = \m7_addr_i[3]_pad  & ~n14451 ;
  assign n39677 = n14468 & n39676 ;
  assign n39678 = ~n39675 & ~n39677 ;
  assign n39679 = n39673 & n39678 ;
  assign n39680 = n39668 & n39679 ;
  assign n39681 = \m3_addr_i[4]_pad  & ~n14451 ;
  assign n39682 = n14459 & n39681 ;
  assign n39683 = \m4_addr_i[4]_pad  & n14451 ;
  assign n39684 = n14444 & n39683 ;
  assign n39685 = ~n39682 & ~n39684 ;
  assign n39686 = \m6_addr_i[4]_pad  & n14451 ;
  assign n39687 = n14468 & n39686 ;
  assign n39688 = \m2_addr_i[4]_pad  & n14451 ;
  assign n39689 = n14459 & n39688 ;
  assign n39690 = ~n39687 & ~n39689 ;
  assign n39691 = n39685 & n39690 ;
  assign n39692 = \m5_addr_i[4]_pad  & ~n14451 ;
  assign n39693 = n14444 & n39692 ;
  assign n39694 = \m1_addr_i[4]_pad  & ~n14451 ;
  assign n39695 = n14476 & n39694 ;
  assign n39696 = ~n39693 & ~n39695 ;
  assign n39697 = \m0_addr_i[4]_pad  & n14451 ;
  assign n39698 = n14476 & n39697 ;
  assign n39699 = \m7_addr_i[4]_pad  & ~n14451 ;
  assign n39700 = n14468 & n39699 ;
  assign n39701 = ~n39698 & ~n39700 ;
  assign n39702 = n39696 & n39701 ;
  assign n39703 = n39691 & n39702 ;
  assign n39704 = \m3_addr_i[5]_pad  & ~n14451 ;
  assign n39705 = n14459 & n39704 ;
  assign n39706 = \m4_addr_i[5]_pad  & n14451 ;
  assign n39707 = n14444 & n39706 ;
  assign n39708 = ~n39705 & ~n39707 ;
  assign n39709 = \m6_addr_i[5]_pad  & n14451 ;
  assign n39710 = n14468 & n39709 ;
  assign n39711 = \m2_addr_i[5]_pad  & n14451 ;
  assign n39712 = n14459 & n39711 ;
  assign n39713 = ~n39710 & ~n39712 ;
  assign n39714 = n39708 & n39713 ;
  assign n39715 = \m5_addr_i[5]_pad  & ~n14451 ;
  assign n39716 = n14444 & n39715 ;
  assign n39717 = \m1_addr_i[5]_pad  & ~n14451 ;
  assign n39718 = n14476 & n39717 ;
  assign n39719 = ~n39716 & ~n39718 ;
  assign n39720 = \m0_addr_i[5]_pad  & n14451 ;
  assign n39721 = n14476 & n39720 ;
  assign n39722 = \m7_addr_i[5]_pad  & ~n14451 ;
  assign n39723 = n14468 & n39722 ;
  assign n39724 = ~n39721 & ~n39723 ;
  assign n39725 = n39719 & n39724 ;
  assign n39726 = n39714 & n39725 ;
  assign n39727 = \m3_addr_i[6]_pad  & ~n14451 ;
  assign n39728 = n14459 & n39727 ;
  assign n39729 = \m4_addr_i[6]_pad  & n14451 ;
  assign n39730 = n14444 & n39729 ;
  assign n39731 = ~n39728 & ~n39730 ;
  assign n39732 = \m6_addr_i[6]_pad  & n14451 ;
  assign n39733 = n14468 & n39732 ;
  assign n39734 = \m2_addr_i[6]_pad  & n14451 ;
  assign n39735 = n14459 & n39734 ;
  assign n39736 = ~n39733 & ~n39735 ;
  assign n39737 = n39731 & n39736 ;
  assign n39738 = \m5_addr_i[6]_pad  & ~n14451 ;
  assign n39739 = n14444 & n39738 ;
  assign n39740 = \m1_addr_i[6]_pad  & ~n14451 ;
  assign n39741 = n14476 & n39740 ;
  assign n39742 = ~n39739 & ~n39741 ;
  assign n39743 = \m0_addr_i[6]_pad  & n14451 ;
  assign n39744 = n14476 & n39743 ;
  assign n39745 = \m7_addr_i[6]_pad  & ~n14451 ;
  assign n39746 = n14468 & n39745 ;
  assign n39747 = ~n39744 & ~n39746 ;
  assign n39748 = n39742 & n39747 ;
  assign n39749 = n39737 & n39748 ;
  assign n39750 = \m3_addr_i[7]_pad  & ~n14451 ;
  assign n39751 = n14459 & n39750 ;
  assign n39752 = \m4_addr_i[7]_pad  & n14451 ;
  assign n39753 = n14444 & n39752 ;
  assign n39754 = ~n39751 & ~n39753 ;
  assign n39755 = \m6_addr_i[7]_pad  & n14451 ;
  assign n39756 = n14468 & n39755 ;
  assign n39757 = \m2_addr_i[7]_pad  & n14451 ;
  assign n39758 = n14459 & n39757 ;
  assign n39759 = ~n39756 & ~n39758 ;
  assign n39760 = n39754 & n39759 ;
  assign n39761 = \m5_addr_i[7]_pad  & ~n14451 ;
  assign n39762 = n14444 & n39761 ;
  assign n39763 = \m1_addr_i[7]_pad  & ~n14451 ;
  assign n39764 = n14476 & n39763 ;
  assign n39765 = ~n39762 & ~n39764 ;
  assign n39766 = \m0_addr_i[7]_pad  & n14451 ;
  assign n39767 = n14476 & n39766 ;
  assign n39768 = \m7_addr_i[7]_pad  & ~n14451 ;
  assign n39769 = n14468 & n39768 ;
  assign n39770 = ~n39767 & ~n39769 ;
  assign n39771 = n39765 & n39770 ;
  assign n39772 = n39760 & n39771 ;
  assign n39773 = \m3_addr_i[8]_pad  & ~n14451 ;
  assign n39774 = n14459 & n39773 ;
  assign n39775 = \m4_addr_i[8]_pad  & n14451 ;
  assign n39776 = n14444 & n39775 ;
  assign n39777 = ~n39774 & ~n39776 ;
  assign n39778 = \m6_addr_i[8]_pad  & n14451 ;
  assign n39779 = n14468 & n39778 ;
  assign n39780 = \m2_addr_i[8]_pad  & n14451 ;
  assign n39781 = n14459 & n39780 ;
  assign n39782 = ~n39779 & ~n39781 ;
  assign n39783 = n39777 & n39782 ;
  assign n39784 = \m5_addr_i[8]_pad  & ~n14451 ;
  assign n39785 = n14444 & n39784 ;
  assign n39786 = \m1_addr_i[8]_pad  & ~n14451 ;
  assign n39787 = n14476 & n39786 ;
  assign n39788 = ~n39785 & ~n39787 ;
  assign n39789 = \m0_addr_i[8]_pad  & n14451 ;
  assign n39790 = n14476 & n39789 ;
  assign n39791 = \m7_addr_i[8]_pad  & ~n14451 ;
  assign n39792 = n14468 & n39791 ;
  assign n39793 = ~n39790 & ~n39792 ;
  assign n39794 = n39788 & n39793 ;
  assign n39795 = n39783 & n39794 ;
  assign n39796 = \m3_addr_i[9]_pad  & ~n14451 ;
  assign n39797 = n14459 & n39796 ;
  assign n39798 = \m4_addr_i[9]_pad  & n14451 ;
  assign n39799 = n14444 & n39798 ;
  assign n39800 = ~n39797 & ~n39799 ;
  assign n39801 = \m6_addr_i[9]_pad  & n14451 ;
  assign n39802 = n14468 & n39801 ;
  assign n39803 = \m2_addr_i[9]_pad  & n14451 ;
  assign n39804 = n14459 & n39803 ;
  assign n39805 = ~n39802 & ~n39804 ;
  assign n39806 = n39800 & n39805 ;
  assign n39807 = \m5_addr_i[9]_pad  & ~n14451 ;
  assign n39808 = n14444 & n39807 ;
  assign n39809 = \m1_addr_i[9]_pad  & ~n14451 ;
  assign n39810 = n14476 & n39809 ;
  assign n39811 = ~n39808 & ~n39810 ;
  assign n39812 = \m0_addr_i[9]_pad  & n14451 ;
  assign n39813 = n14476 & n39812 ;
  assign n39814 = \m7_addr_i[9]_pad  & ~n14451 ;
  assign n39815 = n14468 & n39814 ;
  assign n39816 = ~n39813 & ~n39815 ;
  assign n39817 = n39811 & n39816 ;
  assign n39818 = n39806 & n39817 ;
  assign n39819 = \m3_data_i[0]_pad  & ~n14451 ;
  assign n39820 = n14459 & n39819 ;
  assign n39821 = \m4_data_i[0]_pad  & n14451 ;
  assign n39822 = n14444 & n39821 ;
  assign n39823 = ~n39820 & ~n39822 ;
  assign n39824 = \m6_data_i[0]_pad  & n14451 ;
  assign n39825 = n14468 & n39824 ;
  assign n39826 = \m2_data_i[0]_pad  & n14451 ;
  assign n39827 = n14459 & n39826 ;
  assign n39828 = ~n39825 & ~n39827 ;
  assign n39829 = n39823 & n39828 ;
  assign n39830 = \m5_data_i[0]_pad  & ~n14451 ;
  assign n39831 = n14444 & n39830 ;
  assign n39832 = \m1_data_i[0]_pad  & ~n14451 ;
  assign n39833 = n14476 & n39832 ;
  assign n39834 = ~n39831 & ~n39833 ;
  assign n39835 = \m0_data_i[0]_pad  & n14451 ;
  assign n39836 = n14476 & n39835 ;
  assign n39837 = \m7_data_i[0]_pad  & ~n14451 ;
  assign n39838 = n14468 & n39837 ;
  assign n39839 = ~n39836 & ~n39838 ;
  assign n39840 = n39834 & n39839 ;
  assign n39841 = n39829 & n39840 ;
  assign n39842 = \m3_data_i[10]_pad  & ~n14451 ;
  assign n39843 = n14459 & n39842 ;
  assign n39844 = \m4_data_i[10]_pad  & n14451 ;
  assign n39845 = n14444 & n39844 ;
  assign n39846 = ~n39843 & ~n39845 ;
  assign n39847 = \m6_data_i[10]_pad  & n14451 ;
  assign n39848 = n14468 & n39847 ;
  assign n39849 = \m2_data_i[10]_pad  & n14451 ;
  assign n39850 = n14459 & n39849 ;
  assign n39851 = ~n39848 & ~n39850 ;
  assign n39852 = n39846 & n39851 ;
  assign n39853 = \m5_data_i[10]_pad  & ~n14451 ;
  assign n39854 = n14444 & n39853 ;
  assign n39855 = \m1_data_i[10]_pad  & ~n14451 ;
  assign n39856 = n14476 & n39855 ;
  assign n39857 = ~n39854 & ~n39856 ;
  assign n39858 = \m0_data_i[10]_pad  & n14451 ;
  assign n39859 = n14476 & n39858 ;
  assign n39860 = \m7_data_i[10]_pad  & ~n14451 ;
  assign n39861 = n14468 & n39860 ;
  assign n39862 = ~n39859 & ~n39861 ;
  assign n39863 = n39857 & n39862 ;
  assign n39864 = n39852 & n39863 ;
  assign n39865 = \m3_data_i[11]_pad  & ~n14451 ;
  assign n39866 = n14459 & n39865 ;
  assign n39867 = \m4_data_i[11]_pad  & n14451 ;
  assign n39868 = n14444 & n39867 ;
  assign n39869 = ~n39866 & ~n39868 ;
  assign n39870 = \m6_data_i[11]_pad  & n14451 ;
  assign n39871 = n14468 & n39870 ;
  assign n39872 = \m2_data_i[11]_pad  & n14451 ;
  assign n39873 = n14459 & n39872 ;
  assign n39874 = ~n39871 & ~n39873 ;
  assign n39875 = n39869 & n39874 ;
  assign n39876 = \m5_data_i[11]_pad  & ~n14451 ;
  assign n39877 = n14444 & n39876 ;
  assign n39878 = \m1_data_i[11]_pad  & ~n14451 ;
  assign n39879 = n14476 & n39878 ;
  assign n39880 = ~n39877 & ~n39879 ;
  assign n39881 = \m0_data_i[11]_pad  & n14451 ;
  assign n39882 = n14476 & n39881 ;
  assign n39883 = \m7_data_i[11]_pad  & ~n14451 ;
  assign n39884 = n14468 & n39883 ;
  assign n39885 = ~n39882 & ~n39884 ;
  assign n39886 = n39880 & n39885 ;
  assign n39887 = n39875 & n39886 ;
  assign n39888 = \m3_data_i[12]_pad  & ~n14451 ;
  assign n39889 = n14459 & n39888 ;
  assign n39890 = \m4_data_i[12]_pad  & n14451 ;
  assign n39891 = n14444 & n39890 ;
  assign n39892 = ~n39889 & ~n39891 ;
  assign n39893 = \m6_data_i[12]_pad  & n14451 ;
  assign n39894 = n14468 & n39893 ;
  assign n39895 = \m2_data_i[12]_pad  & n14451 ;
  assign n39896 = n14459 & n39895 ;
  assign n39897 = ~n39894 & ~n39896 ;
  assign n39898 = n39892 & n39897 ;
  assign n39899 = \m5_data_i[12]_pad  & ~n14451 ;
  assign n39900 = n14444 & n39899 ;
  assign n39901 = \m1_data_i[12]_pad  & ~n14451 ;
  assign n39902 = n14476 & n39901 ;
  assign n39903 = ~n39900 & ~n39902 ;
  assign n39904 = \m0_data_i[12]_pad  & n14451 ;
  assign n39905 = n14476 & n39904 ;
  assign n39906 = \m7_data_i[12]_pad  & ~n14451 ;
  assign n39907 = n14468 & n39906 ;
  assign n39908 = ~n39905 & ~n39907 ;
  assign n39909 = n39903 & n39908 ;
  assign n39910 = n39898 & n39909 ;
  assign n39911 = \m3_data_i[13]_pad  & ~n14451 ;
  assign n39912 = n14459 & n39911 ;
  assign n39913 = \m4_data_i[13]_pad  & n14451 ;
  assign n39914 = n14444 & n39913 ;
  assign n39915 = ~n39912 & ~n39914 ;
  assign n39916 = \m6_data_i[13]_pad  & n14451 ;
  assign n39917 = n14468 & n39916 ;
  assign n39918 = \m2_data_i[13]_pad  & n14451 ;
  assign n39919 = n14459 & n39918 ;
  assign n39920 = ~n39917 & ~n39919 ;
  assign n39921 = n39915 & n39920 ;
  assign n39922 = \m5_data_i[13]_pad  & ~n14451 ;
  assign n39923 = n14444 & n39922 ;
  assign n39924 = \m1_data_i[13]_pad  & ~n14451 ;
  assign n39925 = n14476 & n39924 ;
  assign n39926 = ~n39923 & ~n39925 ;
  assign n39927 = \m0_data_i[13]_pad  & n14451 ;
  assign n39928 = n14476 & n39927 ;
  assign n39929 = \m7_data_i[13]_pad  & ~n14451 ;
  assign n39930 = n14468 & n39929 ;
  assign n39931 = ~n39928 & ~n39930 ;
  assign n39932 = n39926 & n39931 ;
  assign n39933 = n39921 & n39932 ;
  assign n39934 = \m3_data_i[14]_pad  & ~n14451 ;
  assign n39935 = n14459 & n39934 ;
  assign n39936 = \m4_data_i[14]_pad  & n14451 ;
  assign n39937 = n14444 & n39936 ;
  assign n39938 = ~n39935 & ~n39937 ;
  assign n39939 = \m6_data_i[14]_pad  & n14451 ;
  assign n39940 = n14468 & n39939 ;
  assign n39941 = \m2_data_i[14]_pad  & n14451 ;
  assign n39942 = n14459 & n39941 ;
  assign n39943 = ~n39940 & ~n39942 ;
  assign n39944 = n39938 & n39943 ;
  assign n39945 = \m5_data_i[14]_pad  & ~n14451 ;
  assign n39946 = n14444 & n39945 ;
  assign n39947 = \m1_data_i[14]_pad  & ~n14451 ;
  assign n39948 = n14476 & n39947 ;
  assign n39949 = ~n39946 & ~n39948 ;
  assign n39950 = \m0_data_i[14]_pad  & n14451 ;
  assign n39951 = n14476 & n39950 ;
  assign n39952 = \m7_data_i[14]_pad  & ~n14451 ;
  assign n39953 = n14468 & n39952 ;
  assign n39954 = ~n39951 & ~n39953 ;
  assign n39955 = n39949 & n39954 ;
  assign n39956 = n39944 & n39955 ;
  assign n39957 = \m3_data_i[15]_pad  & ~n14451 ;
  assign n39958 = n14459 & n39957 ;
  assign n39959 = \m4_data_i[15]_pad  & n14451 ;
  assign n39960 = n14444 & n39959 ;
  assign n39961 = ~n39958 & ~n39960 ;
  assign n39962 = \m6_data_i[15]_pad  & n14451 ;
  assign n39963 = n14468 & n39962 ;
  assign n39964 = \m2_data_i[15]_pad  & n14451 ;
  assign n39965 = n14459 & n39964 ;
  assign n39966 = ~n39963 & ~n39965 ;
  assign n39967 = n39961 & n39966 ;
  assign n39968 = \m5_data_i[15]_pad  & ~n14451 ;
  assign n39969 = n14444 & n39968 ;
  assign n39970 = \m1_data_i[15]_pad  & ~n14451 ;
  assign n39971 = n14476 & n39970 ;
  assign n39972 = ~n39969 & ~n39971 ;
  assign n39973 = \m0_data_i[15]_pad  & n14451 ;
  assign n39974 = n14476 & n39973 ;
  assign n39975 = \m7_data_i[15]_pad  & ~n14451 ;
  assign n39976 = n14468 & n39975 ;
  assign n39977 = ~n39974 & ~n39976 ;
  assign n39978 = n39972 & n39977 ;
  assign n39979 = n39967 & n39978 ;
  assign n39980 = \m3_data_i[16]_pad  & ~n14451 ;
  assign n39981 = n14459 & n39980 ;
  assign n39982 = \m4_data_i[16]_pad  & n14451 ;
  assign n39983 = n14444 & n39982 ;
  assign n39984 = ~n39981 & ~n39983 ;
  assign n39985 = \m6_data_i[16]_pad  & n14451 ;
  assign n39986 = n14468 & n39985 ;
  assign n39987 = \m2_data_i[16]_pad  & n14451 ;
  assign n39988 = n14459 & n39987 ;
  assign n39989 = ~n39986 & ~n39988 ;
  assign n39990 = n39984 & n39989 ;
  assign n39991 = \m5_data_i[16]_pad  & ~n14451 ;
  assign n39992 = n14444 & n39991 ;
  assign n39993 = \m1_data_i[16]_pad  & ~n14451 ;
  assign n39994 = n14476 & n39993 ;
  assign n39995 = ~n39992 & ~n39994 ;
  assign n39996 = \m0_data_i[16]_pad  & n14451 ;
  assign n39997 = n14476 & n39996 ;
  assign n39998 = \m7_data_i[16]_pad  & ~n14451 ;
  assign n39999 = n14468 & n39998 ;
  assign n40000 = ~n39997 & ~n39999 ;
  assign n40001 = n39995 & n40000 ;
  assign n40002 = n39990 & n40001 ;
  assign n40003 = \m3_data_i[17]_pad  & ~n14451 ;
  assign n40004 = n14459 & n40003 ;
  assign n40005 = \m4_data_i[17]_pad  & n14451 ;
  assign n40006 = n14444 & n40005 ;
  assign n40007 = ~n40004 & ~n40006 ;
  assign n40008 = \m6_data_i[17]_pad  & n14451 ;
  assign n40009 = n14468 & n40008 ;
  assign n40010 = \m2_data_i[17]_pad  & n14451 ;
  assign n40011 = n14459 & n40010 ;
  assign n40012 = ~n40009 & ~n40011 ;
  assign n40013 = n40007 & n40012 ;
  assign n40014 = \m5_data_i[17]_pad  & ~n14451 ;
  assign n40015 = n14444 & n40014 ;
  assign n40016 = \m1_data_i[17]_pad  & ~n14451 ;
  assign n40017 = n14476 & n40016 ;
  assign n40018 = ~n40015 & ~n40017 ;
  assign n40019 = \m0_data_i[17]_pad  & n14451 ;
  assign n40020 = n14476 & n40019 ;
  assign n40021 = \m7_data_i[17]_pad  & ~n14451 ;
  assign n40022 = n14468 & n40021 ;
  assign n40023 = ~n40020 & ~n40022 ;
  assign n40024 = n40018 & n40023 ;
  assign n40025 = n40013 & n40024 ;
  assign n40026 = \m3_data_i[18]_pad  & ~n14451 ;
  assign n40027 = n14459 & n40026 ;
  assign n40028 = \m4_data_i[18]_pad  & n14451 ;
  assign n40029 = n14444 & n40028 ;
  assign n40030 = ~n40027 & ~n40029 ;
  assign n40031 = \m6_data_i[18]_pad  & n14451 ;
  assign n40032 = n14468 & n40031 ;
  assign n40033 = \m2_data_i[18]_pad  & n14451 ;
  assign n40034 = n14459 & n40033 ;
  assign n40035 = ~n40032 & ~n40034 ;
  assign n40036 = n40030 & n40035 ;
  assign n40037 = \m5_data_i[18]_pad  & ~n14451 ;
  assign n40038 = n14444 & n40037 ;
  assign n40039 = \m1_data_i[18]_pad  & ~n14451 ;
  assign n40040 = n14476 & n40039 ;
  assign n40041 = ~n40038 & ~n40040 ;
  assign n40042 = \m0_data_i[18]_pad  & n14451 ;
  assign n40043 = n14476 & n40042 ;
  assign n40044 = \m7_data_i[18]_pad  & ~n14451 ;
  assign n40045 = n14468 & n40044 ;
  assign n40046 = ~n40043 & ~n40045 ;
  assign n40047 = n40041 & n40046 ;
  assign n40048 = n40036 & n40047 ;
  assign n40049 = \m3_data_i[19]_pad  & ~n14451 ;
  assign n40050 = n14459 & n40049 ;
  assign n40051 = \m4_data_i[19]_pad  & n14451 ;
  assign n40052 = n14444 & n40051 ;
  assign n40053 = ~n40050 & ~n40052 ;
  assign n40054 = \m6_data_i[19]_pad  & n14451 ;
  assign n40055 = n14468 & n40054 ;
  assign n40056 = \m2_data_i[19]_pad  & n14451 ;
  assign n40057 = n14459 & n40056 ;
  assign n40058 = ~n40055 & ~n40057 ;
  assign n40059 = n40053 & n40058 ;
  assign n40060 = \m5_data_i[19]_pad  & ~n14451 ;
  assign n40061 = n14444 & n40060 ;
  assign n40062 = \m1_data_i[19]_pad  & ~n14451 ;
  assign n40063 = n14476 & n40062 ;
  assign n40064 = ~n40061 & ~n40063 ;
  assign n40065 = \m0_data_i[19]_pad  & n14451 ;
  assign n40066 = n14476 & n40065 ;
  assign n40067 = \m7_data_i[19]_pad  & ~n14451 ;
  assign n40068 = n14468 & n40067 ;
  assign n40069 = ~n40066 & ~n40068 ;
  assign n40070 = n40064 & n40069 ;
  assign n40071 = n40059 & n40070 ;
  assign n40072 = \m3_data_i[1]_pad  & ~n14451 ;
  assign n40073 = n14459 & n40072 ;
  assign n40074 = \m4_data_i[1]_pad  & n14451 ;
  assign n40075 = n14444 & n40074 ;
  assign n40076 = ~n40073 & ~n40075 ;
  assign n40077 = \m6_data_i[1]_pad  & n14451 ;
  assign n40078 = n14468 & n40077 ;
  assign n40079 = \m2_data_i[1]_pad  & n14451 ;
  assign n40080 = n14459 & n40079 ;
  assign n40081 = ~n40078 & ~n40080 ;
  assign n40082 = n40076 & n40081 ;
  assign n40083 = \m5_data_i[1]_pad  & ~n14451 ;
  assign n40084 = n14444 & n40083 ;
  assign n40085 = \m1_data_i[1]_pad  & ~n14451 ;
  assign n40086 = n14476 & n40085 ;
  assign n40087 = ~n40084 & ~n40086 ;
  assign n40088 = \m0_data_i[1]_pad  & n14451 ;
  assign n40089 = n14476 & n40088 ;
  assign n40090 = \m7_data_i[1]_pad  & ~n14451 ;
  assign n40091 = n14468 & n40090 ;
  assign n40092 = ~n40089 & ~n40091 ;
  assign n40093 = n40087 & n40092 ;
  assign n40094 = n40082 & n40093 ;
  assign n40095 = \m3_data_i[20]_pad  & ~n14451 ;
  assign n40096 = n14459 & n40095 ;
  assign n40097 = \m4_data_i[20]_pad  & n14451 ;
  assign n40098 = n14444 & n40097 ;
  assign n40099 = ~n40096 & ~n40098 ;
  assign n40100 = \m6_data_i[20]_pad  & n14451 ;
  assign n40101 = n14468 & n40100 ;
  assign n40102 = \m2_data_i[20]_pad  & n14451 ;
  assign n40103 = n14459 & n40102 ;
  assign n40104 = ~n40101 & ~n40103 ;
  assign n40105 = n40099 & n40104 ;
  assign n40106 = \m5_data_i[20]_pad  & ~n14451 ;
  assign n40107 = n14444 & n40106 ;
  assign n40108 = \m1_data_i[20]_pad  & ~n14451 ;
  assign n40109 = n14476 & n40108 ;
  assign n40110 = ~n40107 & ~n40109 ;
  assign n40111 = \m0_data_i[20]_pad  & n14451 ;
  assign n40112 = n14476 & n40111 ;
  assign n40113 = \m7_data_i[20]_pad  & ~n14451 ;
  assign n40114 = n14468 & n40113 ;
  assign n40115 = ~n40112 & ~n40114 ;
  assign n40116 = n40110 & n40115 ;
  assign n40117 = n40105 & n40116 ;
  assign n40118 = \m3_data_i[21]_pad  & ~n14451 ;
  assign n40119 = n14459 & n40118 ;
  assign n40120 = \m4_data_i[21]_pad  & n14451 ;
  assign n40121 = n14444 & n40120 ;
  assign n40122 = ~n40119 & ~n40121 ;
  assign n40123 = \m6_data_i[21]_pad  & n14451 ;
  assign n40124 = n14468 & n40123 ;
  assign n40125 = \m2_data_i[21]_pad  & n14451 ;
  assign n40126 = n14459 & n40125 ;
  assign n40127 = ~n40124 & ~n40126 ;
  assign n40128 = n40122 & n40127 ;
  assign n40129 = \m5_data_i[21]_pad  & ~n14451 ;
  assign n40130 = n14444 & n40129 ;
  assign n40131 = \m1_data_i[21]_pad  & ~n14451 ;
  assign n40132 = n14476 & n40131 ;
  assign n40133 = ~n40130 & ~n40132 ;
  assign n40134 = \m0_data_i[21]_pad  & n14451 ;
  assign n40135 = n14476 & n40134 ;
  assign n40136 = \m7_data_i[21]_pad  & ~n14451 ;
  assign n40137 = n14468 & n40136 ;
  assign n40138 = ~n40135 & ~n40137 ;
  assign n40139 = n40133 & n40138 ;
  assign n40140 = n40128 & n40139 ;
  assign n40141 = \m3_data_i[22]_pad  & ~n14451 ;
  assign n40142 = n14459 & n40141 ;
  assign n40143 = \m4_data_i[22]_pad  & n14451 ;
  assign n40144 = n14444 & n40143 ;
  assign n40145 = ~n40142 & ~n40144 ;
  assign n40146 = \m6_data_i[22]_pad  & n14451 ;
  assign n40147 = n14468 & n40146 ;
  assign n40148 = \m2_data_i[22]_pad  & n14451 ;
  assign n40149 = n14459 & n40148 ;
  assign n40150 = ~n40147 & ~n40149 ;
  assign n40151 = n40145 & n40150 ;
  assign n40152 = \m5_data_i[22]_pad  & ~n14451 ;
  assign n40153 = n14444 & n40152 ;
  assign n40154 = \m1_data_i[22]_pad  & ~n14451 ;
  assign n40155 = n14476 & n40154 ;
  assign n40156 = ~n40153 & ~n40155 ;
  assign n40157 = \m0_data_i[22]_pad  & n14451 ;
  assign n40158 = n14476 & n40157 ;
  assign n40159 = \m7_data_i[22]_pad  & ~n14451 ;
  assign n40160 = n14468 & n40159 ;
  assign n40161 = ~n40158 & ~n40160 ;
  assign n40162 = n40156 & n40161 ;
  assign n40163 = n40151 & n40162 ;
  assign n40164 = \m3_data_i[23]_pad  & ~n14451 ;
  assign n40165 = n14459 & n40164 ;
  assign n40166 = \m4_data_i[23]_pad  & n14451 ;
  assign n40167 = n14444 & n40166 ;
  assign n40168 = ~n40165 & ~n40167 ;
  assign n40169 = \m6_data_i[23]_pad  & n14451 ;
  assign n40170 = n14468 & n40169 ;
  assign n40171 = \m2_data_i[23]_pad  & n14451 ;
  assign n40172 = n14459 & n40171 ;
  assign n40173 = ~n40170 & ~n40172 ;
  assign n40174 = n40168 & n40173 ;
  assign n40175 = \m5_data_i[23]_pad  & ~n14451 ;
  assign n40176 = n14444 & n40175 ;
  assign n40177 = \m1_data_i[23]_pad  & ~n14451 ;
  assign n40178 = n14476 & n40177 ;
  assign n40179 = ~n40176 & ~n40178 ;
  assign n40180 = \m0_data_i[23]_pad  & n14451 ;
  assign n40181 = n14476 & n40180 ;
  assign n40182 = \m7_data_i[23]_pad  & ~n14451 ;
  assign n40183 = n14468 & n40182 ;
  assign n40184 = ~n40181 & ~n40183 ;
  assign n40185 = n40179 & n40184 ;
  assign n40186 = n40174 & n40185 ;
  assign n40187 = \m3_data_i[24]_pad  & ~n14451 ;
  assign n40188 = n14459 & n40187 ;
  assign n40189 = \m4_data_i[24]_pad  & n14451 ;
  assign n40190 = n14444 & n40189 ;
  assign n40191 = ~n40188 & ~n40190 ;
  assign n40192 = \m6_data_i[24]_pad  & n14451 ;
  assign n40193 = n14468 & n40192 ;
  assign n40194 = \m2_data_i[24]_pad  & n14451 ;
  assign n40195 = n14459 & n40194 ;
  assign n40196 = ~n40193 & ~n40195 ;
  assign n40197 = n40191 & n40196 ;
  assign n40198 = \m5_data_i[24]_pad  & ~n14451 ;
  assign n40199 = n14444 & n40198 ;
  assign n40200 = \m1_data_i[24]_pad  & ~n14451 ;
  assign n40201 = n14476 & n40200 ;
  assign n40202 = ~n40199 & ~n40201 ;
  assign n40203 = \m0_data_i[24]_pad  & n14451 ;
  assign n40204 = n14476 & n40203 ;
  assign n40205 = \m7_data_i[24]_pad  & ~n14451 ;
  assign n40206 = n14468 & n40205 ;
  assign n40207 = ~n40204 & ~n40206 ;
  assign n40208 = n40202 & n40207 ;
  assign n40209 = n40197 & n40208 ;
  assign n40210 = \m3_data_i[25]_pad  & ~n14451 ;
  assign n40211 = n14459 & n40210 ;
  assign n40212 = \m4_data_i[25]_pad  & n14451 ;
  assign n40213 = n14444 & n40212 ;
  assign n40214 = ~n40211 & ~n40213 ;
  assign n40215 = \m6_data_i[25]_pad  & n14451 ;
  assign n40216 = n14468 & n40215 ;
  assign n40217 = \m2_data_i[25]_pad  & n14451 ;
  assign n40218 = n14459 & n40217 ;
  assign n40219 = ~n40216 & ~n40218 ;
  assign n40220 = n40214 & n40219 ;
  assign n40221 = \m5_data_i[25]_pad  & ~n14451 ;
  assign n40222 = n14444 & n40221 ;
  assign n40223 = \m1_data_i[25]_pad  & ~n14451 ;
  assign n40224 = n14476 & n40223 ;
  assign n40225 = ~n40222 & ~n40224 ;
  assign n40226 = \m0_data_i[25]_pad  & n14451 ;
  assign n40227 = n14476 & n40226 ;
  assign n40228 = \m7_data_i[25]_pad  & ~n14451 ;
  assign n40229 = n14468 & n40228 ;
  assign n40230 = ~n40227 & ~n40229 ;
  assign n40231 = n40225 & n40230 ;
  assign n40232 = n40220 & n40231 ;
  assign n40233 = \m3_data_i[26]_pad  & ~n14451 ;
  assign n40234 = n14459 & n40233 ;
  assign n40235 = \m4_data_i[26]_pad  & n14451 ;
  assign n40236 = n14444 & n40235 ;
  assign n40237 = ~n40234 & ~n40236 ;
  assign n40238 = \m6_data_i[26]_pad  & n14451 ;
  assign n40239 = n14468 & n40238 ;
  assign n40240 = \m2_data_i[26]_pad  & n14451 ;
  assign n40241 = n14459 & n40240 ;
  assign n40242 = ~n40239 & ~n40241 ;
  assign n40243 = n40237 & n40242 ;
  assign n40244 = \m5_data_i[26]_pad  & ~n14451 ;
  assign n40245 = n14444 & n40244 ;
  assign n40246 = \m1_data_i[26]_pad  & ~n14451 ;
  assign n40247 = n14476 & n40246 ;
  assign n40248 = ~n40245 & ~n40247 ;
  assign n40249 = \m0_data_i[26]_pad  & n14451 ;
  assign n40250 = n14476 & n40249 ;
  assign n40251 = \m7_data_i[26]_pad  & ~n14451 ;
  assign n40252 = n14468 & n40251 ;
  assign n40253 = ~n40250 & ~n40252 ;
  assign n40254 = n40248 & n40253 ;
  assign n40255 = n40243 & n40254 ;
  assign n40256 = \m3_data_i[27]_pad  & ~n14451 ;
  assign n40257 = n14459 & n40256 ;
  assign n40258 = \m4_data_i[27]_pad  & n14451 ;
  assign n40259 = n14444 & n40258 ;
  assign n40260 = ~n40257 & ~n40259 ;
  assign n40261 = \m6_data_i[27]_pad  & n14451 ;
  assign n40262 = n14468 & n40261 ;
  assign n40263 = \m2_data_i[27]_pad  & n14451 ;
  assign n40264 = n14459 & n40263 ;
  assign n40265 = ~n40262 & ~n40264 ;
  assign n40266 = n40260 & n40265 ;
  assign n40267 = \m5_data_i[27]_pad  & ~n14451 ;
  assign n40268 = n14444 & n40267 ;
  assign n40269 = \m1_data_i[27]_pad  & ~n14451 ;
  assign n40270 = n14476 & n40269 ;
  assign n40271 = ~n40268 & ~n40270 ;
  assign n40272 = \m0_data_i[27]_pad  & n14451 ;
  assign n40273 = n14476 & n40272 ;
  assign n40274 = \m7_data_i[27]_pad  & ~n14451 ;
  assign n40275 = n14468 & n40274 ;
  assign n40276 = ~n40273 & ~n40275 ;
  assign n40277 = n40271 & n40276 ;
  assign n40278 = n40266 & n40277 ;
  assign n40279 = \m3_data_i[28]_pad  & ~n14451 ;
  assign n40280 = n14459 & n40279 ;
  assign n40281 = \m4_data_i[28]_pad  & n14451 ;
  assign n40282 = n14444 & n40281 ;
  assign n40283 = ~n40280 & ~n40282 ;
  assign n40284 = \m6_data_i[28]_pad  & n14451 ;
  assign n40285 = n14468 & n40284 ;
  assign n40286 = \m2_data_i[28]_pad  & n14451 ;
  assign n40287 = n14459 & n40286 ;
  assign n40288 = ~n40285 & ~n40287 ;
  assign n40289 = n40283 & n40288 ;
  assign n40290 = \m5_data_i[28]_pad  & ~n14451 ;
  assign n40291 = n14444 & n40290 ;
  assign n40292 = \m1_data_i[28]_pad  & ~n14451 ;
  assign n40293 = n14476 & n40292 ;
  assign n40294 = ~n40291 & ~n40293 ;
  assign n40295 = \m0_data_i[28]_pad  & n14451 ;
  assign n40296 = n14476 & n40295 ;
  assign n40297 = \m7_data_i[28]_pad  & ~n14451 ;
  assign n40298 = n14468 & n40297 ;
  assign n40299 = ~n40296 & ~n40298 ;
  assign n40300 = n40294 & n40299 ;
  assign n40301 = n40289 & n40300 ;
  assign n40302 = \m3_data_i[29]_pad  & ~n14451 ;
  assign n40303 = n14459 & n40302 ;
  assign n40304 = \m4_data_i[29]_pad  & n14451 ;
  assign n40305 = n14444 & n40304 ;
  assign n40306 = ~n40303 & ~n40305 ;
  assign n40307 = \m6_data_i[29]_pad  & n14451 ;
  assign n40308 = n14468 & n40307 ;
  assign n40309 = \m2_data_i[29]_pad  & n14451 ;
  assign n40310 = n14459 & n40309 ;
  assign n40311 = ~n40308 & ~n40310 ;
  assign n40312 = n40306 & n40311 ;
  assign n40313 = \m5_data_i[29]_pad  & ~n14451 ;
  assign n40314 = n14444 & n40313 ;
  assign n40315 = \m1_data_i[29]_pad  & ~n14451 ;
  assign n40316 = n14476 & n40315 ;
  assign n40317 = ~n40314 & ~n40316 ;
  assign n40318 = \m0_data_i[29]_pad  & n14451 ;
  assign n40319 = n14476 & n40318 ;
  assign n40320 = \m7_data_i[29]_pad  & ~n14451 ;
  assign n40321 = n14468 & n40320 ;
  assign n40322 = ~n40319 & ~n40321 ;
  assign n40323 = n40317 & n40322 ;
  assign n40324 = n40312 & n40323 ;
  assign n40325 = \m3_data_i[2]_pad  & ~n14451 ;
  assign n40326 = n14459 & n40325 ;
  assign n40327 = \m4_data_i[2]_pad  & n14451 ;
  assign n40328 = n14444 & n40327 ;
  assign n40329 = ~n40326 & ~n40328 ;
  assign n40330 = \m6_data_i[2]_pad  & n14451 ;
  assign n40331 = n14468 & n40330 ;
  assign n40332 = \m2_data_i[2]_pad  & n14451 ;
  assign n40333 = n14459 & n40332 ;
  assign n40334 = ~n40331 & ~n40333 ;
  assign n40335 = n40329 & n40334 ;
  assign n40336 = \m5_data_i[2]_pad  & ~n14451 ;
  assign n40337 = n14444 & n40336 ;
  assign n40338 = \m1_data_i[2]_pad  & ~n14451 ;
  assign n40339 = n14476 & n40338 ;
  assign n40340 = ~n40337 & ~n40339 ;
  assign n40341 = \m0_data_i[2]_pad  & n14451 ;
  assign n40342 = n14476 & n40341 ;
  assign n40343 = \m7_data_i[2]_pad  & ~n14451 ;
  assign n40344 = n14468 & n40343 ;
  assign n40345 = ~n40342 & ~n40344 ;
  assign n40346 = n40340 & n40345 ;
  assign n40347 = n40335 & n40346 ;
  assign n40348 = \m3_data_i[30]_pad  & ~n14451 ;
  assign n40349 = n14459 & n40348 ;
  assign n40350 = \m4_data_i[30]_pad  & n14451 ;
  assign n40351 = n14444 & n40350 ;
  assign n40352 = ~n40349 & ~n40351 ;
  assign n40353 = \m6_data_i[30]_pad  & n14451 ;
  assign n40354 = n14468 & n40353 ;
  assign n40355 = \m2_data_i[30]_pad  & n14451 ;
  assign n40356 = n14459 & n40355 ;
  assign n40357 = ~n40354 & ~n40356 ;
  assign n40358 = n40352 & n40357 ;
  assign n40359 = \m5_data_i[30]_pad  & ~n14451 ;
  assign n40360 = n14444 & n40359 ;
  assign n40361 = \m1_data_i[30]_pad  & ~n14451 ;
  assign n40362 = n14476 & n40361 ;
  assign n40363 = ~n40360 & ~n40362 ;
  assign n40364 = \m0_data_i[30]_pad  & n14451 ;
  assign n40365 = n14476 & n40364 ;
  assign n40366 = \m7_data_i[30]_pad  & ~n14451 ;
  assign n40367 = n14468 & n40366 ;
  assign n40368 = ~n40365 & ~n40367 ;
  assign n40369 = n40363 & n40368 ;
  assign n40370 = n40358 & n40369 ;
  assign n40371 = \m3_data_i[31]_pad  & ~n14451 ;
  assign n40372 = n14459 & n40371 ;
  assign n40373 = \m4_data_i[31]_pad  & n14451 ;
  assign n40374 = n14444 & n40373 ;
  assign n40375 = ~n40372 & ~n40374 ;
  assign n40376 = \m6_data_i[31]_pad  & n14451 ;
  assign n40377 = n14468 & n40376 ;
  assign n40378 = \m2_data_i[31]_pad  & n14451 ;
  assign n40379 = n14459 & n40378 ;
  assign n40380 = ~n40377 & ~n40379 ;
  assign n40381 = n40375 & n40380 ;
  assign n40382 = \m5_data_i[31]_pad  & ~n14451 ;
  assign n40383 = n14444 & n40382 ;
  assign n40384 = \m1_data_i[31]_pad  & ~n14451 ;
  assign n40385 = n14476 & n40384 ;
  assign n40386 = ~n40383 & ~n40385 ;
  assign n40387 = \m0_data_i[31]_pad  & n14451 ;
  assign n40388 = n14476 & n40387 ;
  assign n40389 = \m7_data_i[31]_pad  & ~n14451 ;
  assign n40390 = n14468 & n40389 ;
  assign n40391 = ~n40388 & ~n40390 ;
  assign n40392 = n40386 & n40391 ;
  assign n40393 = n40381 & n40392 ;
  assign n40394 = \m3_data_i[3]_pad  & ~n14451 ;
  assign n40395 = n14459 & n40394 ;
  assign n40396 = \m4_data_i[3]_pad  & n14451 ;
  assign n40397 = n14444 & n40396 ;
  assign n40398 = ~n40395 & ~n40397 ;
  assign n40399 = \m6_data_i[3]_pad  & n14451 ;
  assign n40400 = n14468 & n40399 ;
  assign n40401 = \m2_data_i[3]_pad  & n14451 ;
  assign n40402 = n14459 & n40401 ;
  assign n40403 = ~n40400 & ~n40402 ;
  assign n40404 = n40398 & n40403 ;
  assign n40405 = \m5_data_i[3]_pad  & ~n14451 ;
  assign n40406 = n14444 & n40405 ;
  assign n40407 = \m1_data_i[3]_pad  & ~n14451 ;
  assign n40408 = n14476 & n40407 ;
  assign n40409 = ~n40406 & ~n40408 ;
  assign n40410 = \m0_data_i[3]_pad  & n14451 ;
  assign n40411 = n14476 & n40410 ;
  assign n40412 = \m7_data_i[3]_pad  & ~n14451 ;
  assign n40413 = n14468 & n40412 ;
  assign n40414 = ~n40411 & ~n40413 ;
  assign n40415 = n40409 & n40414 ;
  assign n40416 = n40404 & n40415 ;
  assign n40417 = \m3_data_i[4]_pad  & ~n14451 ;
  assign n40418 = n14459 & n40417 ;
  assign n40419 = \m4_data_i[4]_pad  & n14451 ;
  assign n40420 = n14444 & n40419 ;
  assign n40421 = ~n40418 & ~n40420 ;
  assign n40422 = \m6_data_i[4]_pad  & n14451 ;
  assign n40423 = n14468 & n40422 ;
  assign n40424 = \m2_data_i[4]_pad  & n14451 ;
  assign n40425 = n14459 & n40424 ;
  assign n40426 = ~n40423 & ~n40425 ;
  assign n40427 = n40421 & n40426 ;
  assign n40428 = \m5_data_i[4]_pad  & ~n14451 ;
  assign n40429 = n14444 & n40428 ;
  assign n40430 = \m1_data_i[4]_pad  & ~n14451 ;
  assign n40431 = n14476 & n40430 ;
  assign n40432 = ~n40429 & ~n40431 ;
  assign n40433 = \m0_data_i[4]_pad  & n14451 ;
  assign n40434 = n14476 & n40433 ;
  assign n40435 = \m7_data_i[4]_pad  & ~n14451 ;
  assign n40436 = n14468 & n40435 ;
  assign n40437 = ~n40434 & ~n40436 ;
  assign n40438 = n40432 & n40437 ;
  assign n40439 = n40427 & n40438 ;
  assign n40440 = \m3_data_i[5]_pad  & ~n14451 ;
  assign n40441 = n14459 & n40440 ;
  assign n40442 = \m4_data_i[5]_pad  & n14451 ;
  assign n40443 = n14444 & n40442 ;
  assign n40444 = ~n40441 & ~n40443 ;
  assign n40445 = \m6_data_i[5]_pad  & n14451 ;
  assign n40446 = n14468 & n40445 ;
  assign n40447 = \m2_data_i[5]_pad  & n14451 ;
  assign n40448 = n14459 & n40447 ;
  assign n40449 = ~n40446 & ~n40448 ;
  assign n40450 = n40444 & n40449 ;
  assign n40451 = \m5_data_i[5]_pad  & ~n14451 ;
  assign n40452 = n14444 & n40451 ;
  assign n40453 = \m1_data_i[5]_pad  & ~n14451 ;
  assign n40454 = n14476 & n40453 ;
  assign n40455 = ~n40452 & ~n40454 ;
  assign n40456 = \m0_data_i[5]_pad  & n14451 ;
  assign n40457 = n14476 & n40456 ;
  assign n40458 = \m7_data_i[5]_pad  & ~n14451 ;
  assign n40459 = n14468 & n40458 ;
  assign n40460 = ~n40457 & ~n40459 ;
  assign n40461 = n40455 & n40460 ;
  assign n40462 = n40450 & n40461 ;
  assign n40463 = \m3_data_i[6]_pad  & ~n14451 ;
  assign n40464 = n14459 & n40463 ;
  assign n40465 = \m4_data_i[6]_pad  & n14451 ;
  assign n40466 = n14444 & n40465 ;
  assign n40467 = ~n40464 & ~n40466 ;
  assign n40468 = \m6_data_i[6]_pad  & n14451 ;
  assign n40469 = n14468 & n40468 ;
  assign n40470 = \m2_data_i[6]_pad  & n14451 ;
  assign n40471 = n14459 & n40470 ;
  assign n40472 = ~n40469 & ~n40471 ;
  assign n40473 = n40467 & n40472 ;
  assign n40474 = \m5_data_i[6]_pad  & ~n14451 ;
  assign n40475 = n14444 & n40474 ;
  assign n40476 = \m1_data_i[6]_pad  & ~n14451 ;
  assign n40477 = n14476 & n40476 ;
  assign n40478 = ~n40475 & ~n40477 ;
  assign n40479 = \m0_data_i[6]_pad  & n14451 ;
  assign n40480 = n14476 & n40479 ;
  assign n40481 = \m7_data_i[6]_pad  & ~n14451 ;
  assign n40482 = n14468 & n40481 ;
  assign n40483 = ~n40480 & ~n40482 ;
  assign n40484 = n40478 & n40483 ;
  assign n40485 = n40473 & n40484 ;
  assign n40486 = \m3_data_i[7]_pad  & ~n14451 ;
  assign n40487 = n14459 & n40486 ;
  assign n40488 = \m4_data_i[7]_pad  & n14451 ;
  assign n40489 = n14444 & n40488 ;
  assign n40490 = ~n40487 & ~n40489 ;
  assign n40491 = \m6_data_i[7]_pad  & n14451 ;
  assign n40492 = n14468 & n40491 ;
  assign n40493 = \m2_data_i[7]_pad  & n14451 ;
  assign n40494 = n14459 & n40493 ;
  assign n40495 = ~n40492 & ~n40494 ;
  assign n40496 = n40490 & n40495 ;
  assign n40497 = \m5_data_i[7]_pad  & ~n14451 ;
  assign n40498 = n14444 & n40497 ;
  assign n40499 = \m1_data_i[7]_pad  & ~n14451 ;
  assign n40500 = n14476 & n40499 ;
  assign n40501 = ~n40498 & ~n40500 ;
  assign n40502 = \m0_data_i[7]_pad  & n14451 ;
  assign n40503 = n14476 & n40502 ;
  assign n40504 = \m7_data_i[7]_pad  & ~n14451 ;
  assign n40505 = n14468 & n40504 ;
  assign n40506 = ~n40503 & ~n40505 ;
  assign n40507 = n40501 & n40506 ;
  assign n40508 = n40496 & n40507 ;
  assign n40509 = \m3_data_i[8]_pad  & ~n14451 ;
  assign n40510 = n14459 & n40509 ;
  assign n40511 = \m4_data_i[8]_pad  & n14451 ;
  assign n40512 = n14444 & n40511 ;
  assign n40513 = ~n40510 & ~n40512 ;
  assign n40514 = \m6_data_i[8]_pad  & n14451 ;
  assign n40515 = n14468 & n40514 ;
  assign n40516 = \m2_data_i[8]_pad  & n14451 ;
  assign n40517 = n14459 & n40516 ;
  assign n40518 = ~n40515 & ~n40517 ;
  assign n40519 = n40513 & n40518 ;
  assign n40520 = \m5_data_i[8]_pad  & ~n14451 ;
  assign n40521 = n14444 & n40520 ;
  assign n40522 = \m1_data_i[8]_pad  & ~n14451 ;
  assign n40523 = n14476 & n40522 ;
  assign n40524 = ~n40521 & ~n40523 ;
  assign n40525 = \m0_data_i[8]_pad  & n14451 ;
  assign n40526 = n14476 & n40525 ;
  assign n40527 = \m7_data_i[8]_pad  & ~n14451 ;
  assign n40528 = n14468 & n40527 ;
  assign n40529 = ~n40526 & ~n40528 ;
  assign n40530 = n40524 & n40529 ;
  assign n40531 = n40519 & n40530 ;
  assign n40532 = \m3_data_i[9]_pad  & ~n14451 ;
  assign n40533 = n14459 & n40532 ;
  assign n40534 = \m4_data_i[9]_pad  & n14451 ;
  assign n40535 = n14444 & n40534 ;
  assign n40536 = ~n40533 & ~n40535 ;
  assign n40537 = \m6_data_i[9]_pad  & n14451 ;
  assign n40538 = n14468 & n40537 ;
  assign n40539 = \m2_data_i[9]_pad  & n14451 ;
  assign n40540 = n14459 & n40539 ;
  assign n40541 = ~n40538 & ~n40540 ;
  assign n40542 = n40536 & n40541 ;
  assign n40543 = \m5_data_i[9]_pad  & ~n14451 ;
  assign n40544 = n14444 & n40543 ;
  assign n40545 = \m1_data_i[9]_pad  & ~n14451 ;
  assign n40546 = n14476 & n40545 ;
  assign n40547 = ~n40544 & ~n40546 ;
  assign n40548 = \m0_data_i[9]_pad  & n14451 ;
  assign n40549 = n14476 & n40548 ;
  assign n40550 = \m7_data_i[9]_pad  & ~n14451 ;
  assign n40551 = n14468 & n40550 ;
  assign n40552 = ~n40549 & ~n40551 ;
  assign n40553 = n40547 & n40552 ;
  assign n40554 = n40542 & n40553 ;
  assign n40555 = \m3_sel_i[0]_pad  & ~n14451 ;
  assign n40556 = n14459 & n40555 ;
  assign n40557 = \m4_sel_i[0]_pad  & n14451 ;
  assign n40558 = n14444 & n40557 ;
  assign n40559 = ~n40556 & ~n40558 ;
  assign n40560 = \m6_sel_i[0]_pad  & n14451 ;
  assign n40561 = n14468 & n40560 ;
  assign n40562 = \m2_sel_i[0]_pad  & n14451 ;
  assign n40563 = n14459 & n40562 ;
  assign n40564 = ~n40561 & ~n40563 ;
  assign n40565 = n40559 & n40564 ;
  assign n40566 = \m5_sel_i[0]_pad  & ~n14451 ;
  assign n40567 = n14444 & n40566 ;
  assign n40568 = \m1_sel_i[0]_pad  & ~n14451 ;
  assign n40569 = n14476 & n40568 ;
  assign n40570 = ~n40567 & ~n40569 ;
  assign n40571 = \m0_sel_i[0]_pad  & n14451 ;
  assign n40572 = n14476 & n40571 ;
  assign n40573 = \m7_sel_i[0]_pad  & ~n14451 ;
  assign n40574 = n14468 & n40573 ;
  assign n40575 = ~n40572 & ~n40574 ;
  assign n40576 = n40570 & n40575 ;
  assign n40577 = n40565 & n40576 ;
  assign n40578 = \m3_sel_i[1]_pad  & ~n14451 ;
  assign n40579 = n14459 & n40578 ;
  assign n40580 = \m4_sel_i[1]_pad  & n14451 ;
  assign n40581 = n14444 & n40580 ;
  assign n40582 = ~n40579 & ~n40581 ;
  assign n40583 = \m6_sel_i[1]_pad  & n14451 ;
  assign n40584 = n14468 & n40583 ;
  assign n40585 = \m2_sel_i[1]_pad  & n14451 ;
  assign n40586 = n14459 & n40585 ;
  assign n40587 = ~n40584 & ~n40586 ;
  assign n40588 = n40582 & n40587 ;
  assign n40589 = \m5_sel_i[1]_pad  & ~n14451 ;
  assign n40590 = n14444 & n40589 ;
  assign n40591 = \m1_sel_i[1]_pad  & ~n14451 ;
  assign n40592 = n14476 & n40591 ;
  assign n40593 = ~n40590 & ~n40592 ;
  assign n40594 = \m0_sel_i[1]_pad  & n14451 ;
  assign n40595 = n14476 & n40594 ;
  assign n40596 = \m7_sel_i[1]_pad  & ~n14451 ;
  assign n40597 = n14468 & n40596 ;
  assign n40598 = ~n40595 & ~n40597 ;
  assign n40599 = n40593 & n40598 ;
  assign n40600 = n40588 & n40599 ;
  assign n40601 = \m3_sel_i[2]_pad  & ~n14451 ;
  assign n40602 = n14459 & n40601 ;
  assign n40603 = \m4_sel_i[2]_pad  & n14451 ;
  assign n40604 = n14444 & n40603 ;
  assign n40605 = ~n40602 & ~n40604 ;
  assign n40606 = \m6_sel_i[2]_pad  & n14451 ;
  assign n40607 = n14468 & n40606 ;
  assign n40608 = \m2_sel_i[2]_pad  & n14451 ;
  assign n40609 = n14459 & n40608 ;
  assign n40610 = ~n40607 & ~n40609 ;
  assign n40611 = n40605 & n40610 ;
  assign n40612 = \m5_sel_i[2]_pad  & ~n14451 ;
  assign n40613 = n14444 & n40612 ;
  assign n40614 = \m1_sel_i[2]_pad  & ~n14451 ;
  assign n40615 = n14476 & n40614 ;
  assign n40616 = ~n40613 & ~n40615 ;
  assign n40617 = \m0_sel_i[2]_pad  & n14451 ;
  assign n40618 = n14476 & n40617 ;
  assign n40619 = \m7_sel_i[2]_pad  & ~n14451 ;
  assign n40620 = n14468 & n40619 ;
  assign n40621 = ~n40618 & ~n40620 ;
  assign n40622 = n40616 & n40621 ;
  assign n40623 = n40611 & n40622 ;
  assign n40624 = \m3_sel_i[3]_pad  & ~n14451 ;
  assign n40625 = n14459 & n40624 ;
  assign n40626 = \m4_sel_i[3]_pad  & n14451 ;
  assign n40627 = n14444 & n40626 ;
  assign n40628 = ~n40625 & ~n40627 ;
  assign n40629 = \m6_sel_i[3]_pad  & n14451 ;
  assign n40630 = n14468 & n40629 ;
  assign n40631 = \m2_sel_i[3]_pad  & n14451 ;
  assign n40632 = n14459 & n40631 ;
  assign n40633 = ~n40630 & ~n40632 ;
  assign n40634 = n40628 & n40633 ;
  assign n40635 = \m5_sel_i[3]_pad  & ~n14451 ;
  assign n40636 = n14444 & n40635 ;
  assign n40637 = \m1_sel_i[3]_pad  & ~n14451 ;
  assign n40638 = n14476 & n40637 ;
  assign n40639 = ~n40636 & ~n40638 ;
  assign n40640 = \m0_sel_i[3]_pad  & n14451 ;
  assign n40641 = n14476 & n40640 ;
  assign n40642 = \m7_sel_i[3]_pad  & ~n14451 ;
  assign n40643 = n14468 & n40642 ;
  assign n40644 = ~n40641 & ~n40643 ;
  assign n40645 = n40639 & n40644 ;
  assign n40646 = n40634 & n40645 ;
  assign n40647 = \m7_stb_i_pad  & n15070 ;
  assign n40648 = ~n14451 & n40647 ;
  assign n40649 = n14468 & n40648 ;
  assign n40650 = \m6_stb_i_pad  & n15026 ;
  assign n40651 = n14451 & n40650 ;
  assign n40652 = n14468 & n40651 ;
  assign n40653 = ~n40649 & ~n40652 ;
  assign n40654 = \m2_stb_i_pad  & n14870 ;
  assign n40655 = n14451 & n40654 ;
  assign n40656 = n14459 & n40655 ;
  assign n40657 = \m3_stb_i_pad  & n14801 ;
  assign n40658 = ~n14451 & n40657 ;
  assign n40659 = n14459 & n40658 ;
  assign n40660 = ~n40656 & ~n40659 ;
  assign n40661 = n40653 & n40660 ;
  assign n40662 = \m1_stb_i_pad  & n14820 ;
  assign n40663 = ~n14451 & n40662 ;
  assign n40664 = n14476 & n40663 ;
  assign n40665 = \m5_stb_i_pad  & n14704 ;
  assign n40666 = ~n14451 & n40665 ;
  assign n40667 = n14444 & n40666 ;
  assign n40668 = ~n40664 & ~n40667 ;
  assign n40669 = \m4_stb_i_pad  & n14950 ;
  assign n40670 = n14451 & n40669 ;
  assign n40671 = n14444 & n40670 ;
  assign n40672 = \m0_stb_i_pad  & n14774 ;
  assign n40673 = n14451 & n40672 ;
  assign n40674 = n14476 & n40673 ;
  assign n40675 = ~n40671 & ~n40674 ;
  assign n40676 = n40668 & n40675 ;
  assign n40677 = n40661 & n40676 ;
  assign n40678 = \m3_we_i_pad  & ~n14451 ;
  assign n40679 = n14459 & n40678 ;
  assign n40680 = \m4_we_i_pad  & n14451 ;
  assign n40681 = n14444 & n40680 ;
  assign n40682 = ~n40679 & ~n40681 ;
  assign n40683 = \m6_we_i_pad  & n14451 ;
  assign n40684 = n14468 & n40683 ;
  assign n40685 = \m2_we_i_pad  & n14451 ;
  assign n40686 = n14459 & n40685 ;
  assign n40687 = ~n40684 & ~n40686 ;
  assign n40688 = n40682 & n40687 ;
  assign n40689 = \m5_we_i_pad  & ~n14451 ;
  assign n40690 = n14444 & n40689 ;
  assign n40691 = \m1_we_i_pad  & ~n14451 ;
  assign n40692 = n14476 & n40691 ;
  assign n40693 = ~n40690 & ~n40692 ;
  assign n40694 = \m0_we_i_pad  & n14451 ;
  assign n40695 = n14476 & n40694 ;
  assign n40696 = \m7_we_i_pad  & ~n14451 ;
  assign n40697 = n14468 & n40696 ;
  assign n40698 = ~n40695 & ~n40697 ;
  assign n40699 = n40693 & n40698 ;
  assign n40700 = n40688 & n40699 ;
  assign n40701 = \m3_addr_i[0]_pad  & ~n13467 ;
  assign n40702 = n13484 & n40701 ;
  assign n40703 = \m4_addr_i[0]_pad  & n13467 ;
  assign n40704 = n13460 & n40703 ;
  assign n40705 = ~n40702 & ~n40704 ;
  assign n40706 = \m6_addr_i[0]_pad  & n13467 ;
  assign n40707 = n13492 & n40706 ;
  assign n40708 = \m2_addr_i[0]_pad  & n13467 ;
  assign n40709 = n13484 & n40708 ;
  assign n40710 = ~n40707 & ~n40709 ;
  assign n40711 = n40705 & n40710 ;
  assign n40712 = \m5_addr_i[0]_pad  & ~n13467 ;
  assign n40713 = n13460 & n40712 ;
  assign n40714 = \m1_addr_i[0]_pad  & ~n13467 ;
  assign n40715 = n13475 & n40714 ;
  assign n40716 = ~n40713 & ~n40715 ;
  assign n40717 = \m0_addr_i[0]_pad  & n13467 ;
  assign n40718 = n13475 & n40717 ;
  assign n40719 = \m7_addr_i[0]_pad  & ~n13467 ;
  assign n40720 = n13492 & n40719 ;
  assign n40721 = ~n40718 & ~n40720 ;
  assign n40722 = n40716 & n40721 ;
  assign n40723 = n40711 & n40722 ;
  assign n40724 = \m3_addr_i[10]_pad  & ~n13467 ;
  assign n40725 = n13484 & n40724 ;
  assign n40726 = \m4_addr_i[10]_pad  & n13467 ;
  assign n40727 = n13460 & n40726 ;
  assign n40728 = ~n40725 & ~n40727 ;
  assign n40729 = \m6_addr_i[10]_pad  & n13467 ;
  assign n40730 = n13492 & n40729 ;
  assign n40731 = \m2_addr_i[10]_pad  & n13467 ;
  assign n40732 = n13484 & n40731 ;
  assign n40733 = ~n40730 & ~n40732 ;
  assign n40734 = n40728 & n40733 ;
  assign n40735 = \m5_addr_i[10]_pad  & ~n13467 ;
  assign n40736 = n13460 & n40735 ;
  assign n40737 = \m1_addr_i[10]_pad  & ~n13467 ;
  assign n40738 = n13475 & n40737 ;
  assign n40739 = ~n40736 & ~n40738 ;
  assign n40740 = \m0_addr_i[10]_pad  & n13467 ;
  assign n40741 = n13475 & n40740 ;
  assign n40742 = \m7_addr_i[10]_pad  & ~n13467 ;
  assign n40743 = n13492 & n40742 ;
  assign n40744 = ~n40741 & ~n40743 ;
  assign n40745 = n40739 & n40744 ;
  assign n40746 = n40734 & n40745 ;
  assign n40747 = \m3_addr_i[11]_pad  & ~n13467 ;
  assign n40748 = n13484 & n40747 ;
  assign n40749 = \m4_addr_i[11]_pad  & n13467 ;
  assign n40750 = n13460 & n40749 ;
  assign n40751 = ~n40748 & ~n40750 ;
  assign n40752 = \m6_addr_i[11]_pad  & n13467 ;
  assign n40753 = n13492 & n40752 ;
  assign n40754 = \m2_addr_i[11]_pad  & n13467 ;
  assign n40755 = n13484 & n40754 ;
  assign n40756 = ~n40753 & ~n40755 ;
  assign n40757 = n40751 & n40756 ;
  assign n40758 = \m5_addr_i[11]_pad  & ~n13467 ;
  assign n40759 = n13460 & n40758 ;
  assign n40760 = \m1_addr_i[11]_pad  & ~n13467 ;
  assign n40761 = n13475 & n40760 ;
  assign n40762 = ~n40759 & ~n40761 ;
  assign n40763 = \m0_addr_i[11]_pad  & n13467 ;
  assign n40764 = n13475 & n40763 ;
  assign n40765 = \m7_addr_i[11]_pad  & ~n13467 ;
  assign n40766 = n13492 & n40765 ;
  assign n40767 = ~n40764 & ~n40766 ;
  assign n40768 = n40762 & n40767 ;
  assign n40769 = n40757 & n40768 ;
  assign n40770 = \m3_addr_i[12]_pad  & ~n13467 ;
  assign n40771 = n13484 & n40770 ;
  assign n40772 = \m4_addr_i[12]_pad  & n13467 ;
  assign n40773 = n13460 & n40772 ;
  assign n40774 = ~n40771 & ~n40773 ;
  assign n40775 = \m6_addr_i[12]_pad  & n13467 ;
  assign n40776 = n13492 & n40775 ;
  assign n40777 = \m2_addr_i[12]_pad  & n13467 ;
  assign n40778 = n13484 & n40777 ;
  assign n40779 = ~n40776 & ~n40778 ;
  assign n40780 = n40774 & n40779 ;
  assign n40781 = \m5_addr_i[12]_pad  & ~n13467 ;
  assign n40782 = n13460 & n40781 ;
  assign n40783 = \m1_addr_i[12]_pad  & ~n13467 ;
  assign n40784 = n13475 & n40783 ;
  assign n40785 = ~n40782 & ~n40784 ;
  assign n40786 = \m0_addr_i[12]_pad  & n13467 ;
  assign n40787 = n13475 & n40786 ;
  assign n40788 = \m7_addr_i[12]_pad  & ~n13467 ;
  assign n40789 = n13492 & n40788 ;
  assign n40790 = ~n40787 & ~n40789 ;
  assign n40791 = n40785 & n40790 ;
  assign n40792 = n40780 & n40791 ;
  assign n40793 = \m3_addr_i[13]_pad  & ~n13467 ;
  assign n40794 = n13484 & n40793 ;
  assign n40795 = \m4_addr_i[13]_pad  & n13467 ;
  assign n40796 = n13460 & n40795 ;
  assign n40797 = ~n40794 & ~n40796 ;
  assign n40798 = \m6_addr_i[13]_pad  & n13467 ;
  assign n40799 = n13492 & n40798 ;
  assign n40800 = \m2_addr_i[13]_pad  & n13467 ;
  assign n40801 = n13484 & n40800 ;
  assign n40802 = ~n40799 & ~n40801 ;
  assign n40803 = n40797 & n40802 ;
  assign n40804 = \m5_addr_i[13]_pad  & ~n13467 ;
  assign n40805 = n13460 & n40804 ;
  assign n40806 = \m1_addr_i[13]_pad  & ~n13467 ;
  assign n40807 = n13475 & n40806 ;
  assign n40808 = ~n40805 & ~n40807 ;
  assign n40809 = \m0_addr_i[13]_pad  & n13467 ;
  assign n40810 = n13475 & n40809 ;
  assign n40811 = \m7_addr_i[13]_pad  & ~n13467 ;
  assign n40812 = n13492 & n40811 ;
  assign n40813 = ~n40810 & ~n40812 ;
  assign n40814 = n40808 & n40813 ;
  assign n40815 = n40803 & n40814 ;
  assign n40816 = \m3_addr_i[14]_pad  & ~n13467 ;
  assign n40817 = n13484 & n40816 ;
  assign n40818 = \m4_addr_i[14]_pad  & n13467 ;
  assign n40819 = n13460 & n40818 ;
  assign n40820 = ~n40817 & ~n40819 ;
  assign n40821 = \m6_addr_i[14]_pad  & n13467 ;
  assign n40822 = n13492 & n40821 ;
  assign n40823 = \m2_addr_i[14]_pad  & n13467 ;
  assign n40824 = n13484 & n40823 ;
  assign n40825 = ~n40822 & ~n40824 ;
  assign n40826 = n40820 & n40825 ;
  assign n40827 = \m5_addr_i[14]_pad  & ~n13467 ;
  assign n40828 = n13460 & n40827 ;
  assign n40829 = \m1_addr_i[14]_pad  & ~n13467 ;
  assign n40830 = n13475 & n40829 ;
  assign n40831 = ~n40828 & ~n40830 ;
  assign n40832 = \m0_addr_i[14]_pad  & n13467 ;
  assign n40833 = n13475 & n40832 ;
  assign n40834 = \m7_addr_i[14]_pad  & ~n13467 ;
  assign n40835 = n13492 & n40834 ;
  assign n40836 = ~n40833 & ~n40835 ;
  assign n40837 = n40831 & n40836 ;
  assign n40838 = n40826 & n40837 ;
  assign n40839 = \m3_addr_i[15]_pad  & ~n13467 ;
  assign n40840 = n13484 & n40839 ;
  assign n40841 = \m4_addr_i[15]_pad  & n13467 ;
  assign n40842 = n13460 & n40841 ;
  assign n40843 = ~n40840 & ~n40842 ;
  assign n40844 = \m6_addr_i[15]_pad  & n13467 ;
  assign n40845 = n13492 & n40844 ;
  assign n40846 = \m2_addr_i[15]_pad  & n13467 ;
  assign n40847 = n13484 & n40846 ;
  assign n40848 = ~n40845 & ~n40847 ;
  assign n40849 = n40843 & n40848 ;
  assign n40850 = \m5_addr_i[15]_pad  & ~n13467 ;
  assign n40851 = n13460 & n40850 ;
  assign n40852 = \m1_addr_i[15]_pad  & ~n13467 ;
  assign n40853 = n13475 & n40852 ;
  assign n40854 = ~n40851 & ~n40853 ;
  assign n40855 = \m0_addr_i[15]_pad  & n13467 ;
  assign n40856 = n13475 & n40855 ;
  assign n40857 = \m7_addr_i[15]_pad  & ~n13467 ;
  assign n40858 = n13492 & n40857 ;
  assign n40859 = ~n40856 & ~n40858 ;
  assign n40860 = n40854 & n40859 ;
  assign n40861 = n40849 & n40860 ;
  assign n40862 = \m3_addr_i[16]_pad  & ~n13467 ;
  assign n40863 = n13484 & n40862 ;
  assign n40864 = \m4_addr_i[16]_pad  & n13467 ;
  assign n40865 = n13460 & n40864 ;
  assign n40866 = ~n40863 & ~n40865 ;
  assign n40867 = \m6_addr_i[16]_pad  & n13467 ;
  assign n40868 = n13492 & n40867 ;
  assign n40869 = \m2_addr_i[16]_pad  & n13467 ;
  assign n40870 = n13484 & n40869 ;
  assign n40871 = ~n40868 & ~n40870 ;
  assign n40872 = n40866 & n40871 ;
  assign n40873 = \m5_addr_i[16]_pad  & ~n13467 ;
  assign n40874 = n13460 & n40873 ;
  assign n40875 = \m1_addr_i[16]_pad  & ~n13467 ;
  assign n40876 = n13475 & n40875 ;
  assign n40877 = ~n40874 & ~n40876 ;
  assign n40878 = \m0_addr_i[16]_pad  & n13467 ;
  assign n40879 = n13475 & n40878 ;
  assign n40880 = \m7_addr_i[16]_pad  & ~n13467 ;
  assign n40881 = n13492 & n40880 ;
  assign n40882 = ~n40879 & ~n40881 ;
  assign n40883 = n40877 & n40882 ;
  assign n40884 = n40872 & n40883 ;
  assign n40885 = \m3_addr_i[17]_pad  & ~n13467 ;
  assign n40886 = n13484 & n40885 ;
  assign n40887 = \m4_addr_i[17]_pad  & n13467 ;
  assign n40888 = n13460 & n40887 ;
  assign n40889 = ~n40886 & ~n40888 ;
  assign n40890 = \m6_addr_i[17]_pad  & n13467 ;
  assign n40891 = n13492 & n40890 ;
  assign n40892 = \m2_addr_i[17]_pad  & n13467 ;
  assign n40893 = n13484 & n40892 ;
  assign n40894 = ~n40891 & ~n40893 ;
  assign n40895 = n40889 & n40894 ;
  assign n40896 = \m5_addr_i[17]_pad  & ~n13467 ;
  assign n40897 = n13460 & n40896 ;
  assign n40898 = \m1_addr_i[17]_pad  & ~n13467 ;
  assign n40899 = n13475 & n40898 ;
  assign n40900 = ~n40897 & ~n40899 ;
  assign n40901 = \m0_addr_i[17]_pad  & n13467 ;
  assign n40902 = n13475 & n40901 ;
  assign n40903 = \m7_addr_i[17]_pad  & ~n13467 ;
  assign n40904 = n13492 & n40903 ;
  assign n40905 = ~n40902 & ~n40904 ;
  assign n40906 = n40900 & n40905 ;
  assign n40907 = n40895 & n40906 ;
  assign n40908 = \m3_addr_i[18]_pad  & ~n13467 ;
  assign n40909 = n13484 & n40908 ;
  assign n40910 = \m4_addr_i[18]_pad  & n13467 ;
  assign n40911 = n13460 & n40910 ;
  assign n40912 = ~n40909 & ~n40911 ;
  assign n40913 = \m6_addr_i[18]_pad  & n13467 ;
  assign n40914 = n13492 & n40913 ;
  assign n40915 = \m2_addr_i[18]_pad  & n13467 ;
  assign n40916 = n13484 & n40915 ;
  assign n40917 = ~n40914 & ~n40916 ;
  assign n40918 = n40912 & n40917 ;
  assign n40919 = \m5_addr_i[18]_pad  & ~n13467 ;
  assign n40920 = n13460 & n40919 ;
  assign n40921 = \m1_addr_i[18]_pad  & ~n13467 ;
  assign n40922 = n13475 & n40921 ;
  assign n40923 = ~n40920 & ~n40922 ;
  assign n40924 = \m0_addr_i[18]_pad  & n13467 ;
  assign n40925 = n13475 & n40924 ;
  assign n40926 = \m7_addr_i[18]_pad  & ~n13467 ;
  assign n40927 = n13492 & n40926 ;
  assign n40928 = ~n40925 & ~n40927 ;
  assign n40929 = n40923 & n40928 ;
  assign n40930 = n40918 & n40929 ;
  assign n40931 = \m3_addr_i[19]_pad  & ~n13467 ;
  assign n40932 = n13484 & n40931 ;
  assign n40933 = \m4_addr_i[19]_pad  & n13467 ;
  assign n40934 = n13460 & n40933 ;
  assign n40935 = ~n40932 & ~n40934 ;
  assign n40936 = \m6_addr_i[19]_pad  & n13467 ;
  assign n40937 = n13492 & n40936 ;
  assign n40938 = \m2_addr_i[19]_pad  & n13467 ;
  assign n40939 = n13484 & n40938 ;
  assign n40940 = ~n40937 & ~n40939 ;
  assign n40941 = n40935 & n40940 ;
  assign n40942 = \m5_addr_i[19]_pad  & ~n13467 ;
  assign n40943 = n13460 & n40942 ;
  assign n40944 = \m1_addr_i[19]_pad  & ~n13467 ;
  assign n40945 = n13475 & n40944 ;
  assign n40946 = ~n40943 & ~n40945 ;
  assign n40947 = \m0_addr_i[19]_pad  & n13467 ;
  assign n40948 = n13475 & n40947 ;
  assign n40949 = \m7_addr_i[19]_pad  & ~n13467 ;
  assign n40950 = n13492 & n40949 ;
  assign n40951 = ~n40948 & ~n40950 ;
  assign n40952 = n40946 & n40951 ;
  assign n40953 = n40941 & n40952 ;
  assign n40954 = \m3_addr_i[1]_pad  & ~n13467 ;
  assign n40955 = n13484 & n40954 ;
  assign n40956 = \m4_addr_i[1]_pad  & n13467 ;
  assign n40957 = n13460 & n40956 ;
  assign n40958 = ~n40955 & ~n40957 ;
  assign n40959 = \m6_addr_i[1]_pad  & n13467 ;
  assign n40960 = n13492 & n40959 ;
  assign n40961 = \m2_addr_i[1]_pad  & n13467 ;
  assign n40962 = n13484 & n40961 ;
  assign n40963 = ~n40960 & ~n40962 ;
  assign n40964 = n40958 & n40963 ;
  assign n40965 = \m5_addr_i[1]_pad  & ~n13467 ;
  assign n40966 = n13460 & n40965 ;
  assign n40967 = \m1_addr_i[1]_pad  & ~n13467 ;
  assign n40968 = n13475 & n40967 ;
  assign n40969 = ~n40966 & ~n40968 ;
  assign n40970 = \m0_addr_i[1]_pad  & n13467 ;
  assign n40971 = n13475 & n40970 ;
  assign n40972 = \m7_addr_i[1]_pad  & ~n13467 ;
  assign n40973 = n13492 & n40972 ;
  assign n40974 = ~n40971 & ~n40973 ;
  assign n40975 = n40969 & n40974 ;
  assign n40976 = n40964 & n40975 ;
  assign n40977 = \m3_addr_i[20]_pad  & ~n13467 ;
  assign n40978 = n13484 & n40977 ;
  assign n40979 = \m4_addr_i[20]_pad  & n13467 ;
  assign n40980 = n13460 & n40979 ;
  assign n40981 = ~n40978 & ~n40980 ;
  assign n40982 = \m6_addr_i[20]_pad  & n13467 ;
  assign n40983 = n13492 & n40982 ;
  assign n40984 = \m2_addr_i[20]_pad  & n13467 ;
  assign n40985 = n13484 & n40984 ;
  assign n40986 = ~n40983 & ~n40985 ;
  assign n40987 = n40981 & n40986 ;
  assign n40988 = \m5_addr_i[20]_pad  & ~n13467 ;
  assign n40989 = n13460 & n40988 ;
  assign n40990 = \m1_addr_i[20]_pad  & ~n13467 ;
  assign n40991 = n13475 & n40990 ;
  assign n40992 = ~n40989 & ~n40991 ;
  assign n40993 = \m0_addr_i[20]_pad  & n13467 ;
  assign n40994 = n13475 & n40993 ;
  assign n40995 = \m7_addr_i[20]_pad  & ~n13467 ;
  assign n40996 = n13492 & n40995 ;
  assign n40997 = ~n40994 & ~n40996 ;
  assign n40998 = n40992 & n40997 ;
  assign n40999 = n40987 & n40998 ;
  assign n41000 = \m3_addr_i[21]_pad  & ~n13467 ;
  assign n41001 = n13484 & n41000 ;
  assign n41002 = \m4_addr_i[21]_pad  & n13467 ;
  assign n41003 = n13460 & n41002 ;
  assign n41004 = ~n41001 & ~n41003 ;
  assign n41005 = \m6_addr_i[21]_pad  & n13467 ;
  assign n41006 = n13492 & n41005 ;
  assign n41007 = \m2_addr_i[21]_pad  & n13467 ;
  assign n41008 = n13484 & n41007 ;
  assign n41009 = ~n41006 & ~n41008 ;
  assign n41010 = n41004 & n41009 ;
  assign n41011 = \m5_addr_i[21]_pad  & ~n13467 ;
  assign n41012 = n13460 & n41011 ;
  assign n41013 = \m1_addr_i[21]_pad  & ~n13467 ;
  assign n41014 = n13475 & n41013 ;
  assign n41015 = ~n41012 & ~n41014 ;
  assign n41016 = \m0_addr_i[21]_pad  & n13467 ;
  assign n41017 = n13475 & n41016 ;
  assign n41018 = \m7_addr_i[21]_pad  & ~n13467 ;
  assign n41019 = n13492 & n41018 ;
  assign n41020 = ~n41017 & ~n41019 ;
  assign n41021 = n41015 & n41020 ;
  assign n41022 = n41010 & n41021 ;
  assign n41023 = \m3_addr_i[22]_pad  & ~n13467 ;
  assign n41024 = n13484 & n41023 ;
  assign n41025 = \m4_addr_i[22]_pad  & n13467 ;
  assign n41026 = n13460 & n41025 ;
  assign n41027 = ~n41024 & ~n41026 ;
  assign n41028 = \m6_addr_i[22]_pad  & n13467 ;
  assign n41029 = n13492 & n41028 ;
  assign n41030 = \m2_addr_i[22]_pad  & n13467 ;
  assign n41031 = n13484 & n41030 ;
  assign n41032 = ~n41029 & ~n41031 ;
  assign n41033 = n41027 & n41032 ;
  assign n41034 = \m5_addr_i[22]_pad  & ~n13467 ;
  assign n41035 = n13460 & n41034 ;
  assign n41036 = \m1_addr_i[22]_pad  & ~n13467 ;
  assign n41037 = n13475 & n41036 ;
  assign n41038 = ~n41035 & ~n41037 ;
  assign n41039 = \m0_addr_i[22]_pad  & n13467 ;
  assign n41040 = n13475 & n41039 ;
  assign n41041 = \m7_addr_i[22]_pad  & ~n13467 ;
  assign n41042 = n13492 & n41041 ;
  assign n41043 = ~n41040 & ~n41042 ;
  assign n41044 = n41038 & n41043 ;
  assign n41045 = n41033 & n41044 ;
  assign n41046 = \m3_addr_i[23]_pad  & ~n13467 ;
  assign n41047 = n13484 & n41046 ;
  assign n41048 = \m4_addr_i[23]_pad  & n13467 ;
  assign n41049 = n13460 & n41048 ;
  assign n41050 = ~n41047 & ~n41049 ;
  assign n41051 = \m6_addr_i[23]_pad  & n13467 ;
  assign n41052 = n13492 & n41051 ;
  assign n41053 = \m2_addr_i[23]_pad  & n13467 ;
  assign n41054 = n13484 & n41053 ;
  assign n41055 = ~n41052 & ~n41054 ;
  assign n41056 = n41050 & n41055 ;
  assign n41057 = \m5_addr_i[23]_pad  & ~n13467 ;
  assign n41058 = n13460 & n41057 ;
  assign n41059 = \m1_addr_i[23]_pad  & ~n13467 ;
  assign n41060 = n13475 & n41059 ;
  assign n41061 = ~n41058 & ~n41060 ;
  assign n41062 = \m0_addr_i[23]_pad  & n13467 ;
  assign n41063 = n13475 & n41062 ;
  assign n41064 = \m7_addr_i[23]_pad  & ~n13467 ;
  assign n41065 = n13492 & n41064 ;
  assign n41066 = ~n41063 & ~n41065 ;
  assign n41067 = n41061 & n41066 ;
  assign n41068 = n41056 & n41067 ;
  assign n41069 = \m3_addr_i[24]_pad  & ~n13467 ;
  assign n41070 = n13484 & n41069 ;
  assign n41071 = \m4_addr_i[24]_pad  & n13467 ;
  assign n41072 = n13460 & n41071 ;
  assign n41073 = ~n41070 & ~n41072 ;
  assign n41074 = \m5_addr_i[24]_pad  & ~n13467 ;
  assign n41075 = n13460 & n41074 ;
  assign n41076 = \m2_addr_i[24]_pad  & n13467 ;
  assign n41077 = n13484 & n41076 ;
  assign n41078 = ~n41075 & ~n41077 ;
  assign n41079 = n41073 & n41078 ;
  assign n41080 = \m6_addr_i[24]_pad  & n13467 ;
  assign n41081 = n13492 & n41080 ;
  assign n41082 = \m1_addr_i[24]_pad  & ~n13467 ;
  assign n41083 = n13475 & n41082 ;
  assign n41084 = ~n41081 & ~n41083 ;
  assign n41085 = \m0_addr_i[24]_pad  & n13467 ;
  assign n41086 = n13475 & n41085 ;
  assign n41087 = \m7_addr_i[24]_pad  & ~n13467 ;
  assign n41088 = n13492 & n41087 ;
  assign n41089 = ~n41086 & ~n41088 ;
  assign n41090 = n41084 & n41089 ;
  assign n41091 = n41079 & n41090 ;
  assign n41092 = \m3_addr_i[25]_pad  & ~n13467 ;
  assign n41093 = n13484 & n41092 ;
  assign n41094 = \m4_addr_i[25]_pad  & n13467 ;
  assign n41095 = n13460 & n41094 ;
  assign n41096 = ~n41093 & ~n41095 ;
  assign n41097 = \m5_addr_i[25]_pad  & ~n13467 ;
  assign n41098 = n13460 & n41097 ;
  assign n41099 = \m2_addr_i[25]_pad  & n13467 ;
  assign n41100 = n13484 & n41099 ;
  assign n41101 = ~n41098 & ~n41100 ;
  assign n41102 = n41096 & n41101 ;
  assign n41103 = \m6_addr_i[25]_pad  & n13467 ;
  assign n41104 = n13492 & n41103 ;
  assign n41105 = \m1_addr_i[25]_pad  & ~n13467 ;
  assign n41106 = n13475 & n41105 ;
  assign n41107 = ~n41104 & ~n41106 ;
  assign n41108 = \m0_addr_i[25]_pad  & n13467 ;
  assign n41109 = n13475 & n41108 ;
  assign n41110 = \m7_addr_i[25]_pad  & ~n13467 ;
  assign n41111 = n13492 & n41110 ;
  assign n41112 = ~n41109 & ~n41111 ;
  assign n41113 = n41107 & n41112 ;
  assign n41114 = n41102 & n41113 ;
  assign n41115 = \m3_addr_i[26]_pad  & ~n13467 ;
  assign n41116 = n13484 & n41115 ;
  assign n41117 = \m4_addr_i[26]_pad  & n13467 ;
  assign n41118 = n13460 & n41117 ;
  assign n41119 = ~n41116 & ~n41118 ;
  assign n41120 = \m5_addr_i[26]_pad  & ~n13467 ;
  assign n41121 = n13460 & n41120 ;
  assign n41122 = \m2_addr_i[26]_pad  & n13467 ;
  assign n41123 = n13484 & n41122 ;
  assign n41124 = ~n41121 & ~n41123 ;
  assign n41125 = n41119 & n41124 ;
  assign n41126 = \m6_addr_i[26]_pad  & n13467 ;
  assign n41127 = n13492 & n41126 ;
  assign n41128 = \m1_addr_i[26]_pad  & ~n13467 ;
  assign n41129 = n13475 & n41128 ;
  assign n41130 = ~n41127 & ~n41129 ;
  assign n41131 = \m0_addr_i[26]_pad  & n13467 ;
  assign n41132 = n13475 & n41131 ;
  assign n41133 = \m7_addr_i[26]_pad  & ~n13467 ;
  assign n41134 = n13492 & n41133 ;
  assign n41135 = ~n41132 & ~n41134 ;
  assign n41136 = n41130 & n41135 ;
  assign n41137 = n41125 & n41136 ;
  assign n41138 = \m3_addr_i[27]_pad  & ~n13467 ;
  assign n41139 = n13484 & n41138 ;
  assign n41140 = \m4_addr_i[27]_pad  & n13467 ;
  assign n41141 = n13460 & n41140 ;
  assign n41142 = ~n41139 & ~n41141 ;
  assign n41143 = \m5_addr_i[27]_pad  & ~n13467 ;
  assign n41144 = n13460 & n41143 ;
  assign n41145 = \m2_addr_i[27]_pad  & n13467 ;
  assign n41146 = n13484 & n41145 ;
  assign n41147 = ~n41144 & ~n41146 ;
  assign n41148 = n41142 & n41147 ;
  assign n41149 = \m6_addr_i[27]_pad  & n13467 ;
  assign n41150 = n13492 & n41149 ;
  assign n41151 = \m1_addr_i[27]_pad  & ~n13467 ;
  assign n41152 = n13475 & n41151 ;
  assign n41153 = ~n41150 & ~n41152 ;
  assign n41154 = \m0_addr_i[27]_pad  & n13467 ;
  assign n41155 = n13475 & n41154 ;
  assign n41156 = \m7_addr_i[27]_pad  & ~n13467 ;
  assign n41157 = n13492 & n41156 ;
  assign n41158 = ~n41155 & ~n41157 ;
  assign n41159 = n41153 & n41158 ;
  assign n41160 = n41148 & n41159 ;
  assign n41161 = \m3_addr_i[28]_pad  & ~n13467 ;
  assign n41162 = n13484 & n41161 ;
  assign n41163 = \m4_addr_i[28]_pad  & n13467 ;
  assign n41164 = n13460 & n41163 ;
  assign n41165 = ~n41162 & ~n41164 ;
  assign n41166 = \m5_addr_i[28]_pad  & ~n13467 ;
  assign n41167 = n13460 & n41166 ;
  assign n41168 = \m2_addr_i[28]_pad  & n13467 ;
  assign n41169 = n13484 & n41168 ;
  assign n41170 = ~n41167 & ~n41169 ;
  assign n41171 = n41165 & n41170 ;
  assign n41172 = \m6_addr_i[28]_pad  & n13467 ;
  assign n41173 = n13492 & n41172 ;
  assign n41174 = \m1_addr_i[28]_pad  & ~n13467 ;
  assign n41175 = n13475 & n41174 ;
  assign n41176 = ~n41173 & ~n41175 ;
  assign n41177 = \m0_addr_i[28]_pad  & n13467 ;
  assign n41178 = n13475 & n41177 ;
  assign n41179 = \m7_addr_i[28]_pad  & ~n13467 ;
  assign n41180 = n13492 & n41179 ;
  assign n41181 = ~n41178 & ~n41180 ;
  assign n41182 = n41176 & n41181 ;
  assign n41183 = n41171 & n41182 ;
  assign n41184 = \m3_addr_i[29]_pad  & ~n13467 ;
  assign n41185 = n13484 & n41184 ;
  assign n41186 = \m4_addr_i[29]_pad  & n13467 ;
  assign n41187 = n13460 & n41186 ;
  assign n41188 = ~n41185 & ~n41187 ;
  assign n41189 = \m5_addr_i[29]_pad  & ~n13467 ;
  assign n41190 = n13460 & n41189 ;
  assign n41191 = \m2_addr_i[29]_pad  & n13467 ;
  assign n41192 = n13484 & n41191 ;
  assign n41193 = ~n41190 & ~n41192 ;
  assign n41194 = n41188 & n41193 ;
  assign n41195 = \m6_addr_i[29]_pad  & n13467 ;
  assign n41196 = n13492 & n41195 ;
  assign n41197 = \m1_addr_i[29]_pad  & ~n13467 ;
  assign n41198 = n13475 & n41197 ;
  assign n41199 = ~n41196 & ~n41198 ;
  assign n41200 = \m0_addr_i[29]_pad  & n13467 ;
  assign n41201 = n13475 & n41200 ;
  assign n41202 = \m7_addr_i[29]_pad  & ~n13467 ;
  assign n41203 = n13492 & n41202 ;
  assign n41204 = ~n41201 & ~n41203 ;
  assign n41205 = n41199 & n41204 ;
  assign n41206 = n41194 & n41205 ;
  assign n41207 = \m3_addr_i[2]_pad  & ~n13467 ;
  assign n41208 = n13484 & n41207 ;
  assign n41209 = \m4_addr_i[2]_pad  & n13467 ;
  assign n41210 = n13460 & n41209 ;
  assign n41211 = ~n41208 & ~n41210 ;
  assign n41212 = \m6_addr_i[2]_pad  & n13467 ;
  assign n41213 = n13492 & n41212 ;
  assign n41214 = \m2_addr_i[2]_pad  & n13467 ;
  assign n41215 = n13484 & n41214 ;
  assign n41216 = ~n41213 & ~n41215 ;
  assign n41217 = n41211 & n41216 ;
  assign n41218 = \m5_addr_i[2]_pad  & ~n13467 ;
  assign n41219 = n13460 & n41218 ;
  assign n41220 = \m1_addr_i[2]_pad  & ~n13467 ;
  assign n41221 = n13475 & n41220 ;
  assign n41222 = ~n41219 & ~n41221 ;
  assign n41223 = \m0_addr_i[2]_pad  & n13467 ;
  assign n41224 = n13475 & n41223 ;
  assign n41225 = \m7_addr_i[2]_pad  & ~n13467 ;
  assign n41226 = n13492 & n41225 ;
  assign n41227 = ~n41224 & ~n41226 ;
  assign n41228 = n41222 & n41227 ;
  assign n41229 = n41217 & n41228 ;
  assign n41230 = \m3_addr_i[30]_pad  & ~n13467 ;
  assign n41231 = n13484 & n41230 ;
  assign n41232 = \m4_addr_i[30]_pad  & n13467 ;
  assign n41233 = n13460 & n41232 ;
  assign n41234 = ~n41231 & ~n41233 ;
  assign n41235 = \m5_addr_i[30]_pad  & ~n13467 ;
  assign n41236 = n13460 & n41235 ;
  assign n41237 = \m2_addr_i[30]_pad  & n13467 ;
  assign n41238 = n13484 & n41237 ;
  assign n41239 = ~n41236 & ~n41238 ;
  assign n41240 = n41234 & n41239 ;
  assign n41241 = \m6_addr_i[30]_pad  & n13467 ;
  assign n41242 = n13492 & n41241 ;
  assign n41243 = \m1_addr_i[30]_pad  & ~n13467 ;
  assign n41244 = n13475 & n41243 ;
  assign n41245 = ~n41242 & ~n41244 ;
  assign n41246 = \m0_addr_i[30]_pad  & n13467 ;
  assign n41247 = n13475 & n41246 ;
  assign n41248 = \m7_addr_i[30]_pad  & ~n13467 ;
  assign n41249 = n13492 & n41248 ;
  assign n41250 = ~n41247 & ~n41249 ;
  assign n41251 = n41245 & n41250 ;
  assign n41252 = n41240 & n41251 ;
  assign n41253 = \m3_addr_i[31]_pad  & ~n13467 ;
  assign n41254 = n13484 & n41253 ;
  assign n41255 = \m4_addr_i[31]_pad  & n13467 ;
  assign n41256 = n13460 & n41255 ;
  assign n41257 = ~n41254 & ~n41256 ;
  assign n41258 = \m5_addr_i[31]_pad  & ~n13467 ;
  assign n41259 = n13460 & n41258 ;
  assign n41260 = \m2_addr_i[31]_pad  & n13467 ;
  assign n41261 = n13484 & n41260 ;
  assign n41262 = ~n41259 & ~n41261 ;
  assign n41263 = n41257 & n41262 ;
  assign n41264 = \m6_addr_i[31]_pad  & n13467 ;
  assign n41265 = n13492 & n41264 ;
  assign n41266 = \m1_addr_i[31]_pad  & ~n13467 ;
  assign n41267 = n13475 & n41266 ;
  assign n41268 = ~n41265 & ~n41267 ;
  assign n41269 = \m0_addr_i[31]_pad  & n13467 ;
  assign n41270 = n13475 & n41269 ;
  assign n41271 = \m7_addr_i[31]_pad  & ~n13467 ;
  assign n41272 = n13492 & n41271 ;
  assign n41273 = ~n41270 & ~n41272 ;
  assign n41274 = n41268 & n41273 ;
  assign n41275 = n41263 & n41274 ;
  assign n41276 = \m3_addr_i[3]_pad  & ~n13467 ;
  assign n41277 = n13484 & n41276 ;
  assign n41278 = \m4_addr_i[3]_pad  & n13467 ;
  assign n41279 = n13460 & n41278 ;
  assign n41280 = ~n41277 & ~n41279 ;
  assign n41281 = \m6_addr_i[3]_pad  & n13467 ;
  assign n41282 = n13492 & n41281 ;
  assign n41283 = \m2_addr_i[3]_pad  & n13467 ;
  assign n41284 = n13484 & n41283 ;
  assign n41285 = ~n41282 & ~n41284 ;
  assign n41286 = n41280 & n41285 ;
  assign n41287 = \m5_addr_i[3]_pad  & ~n13467 ;
  assign n41288 = n13460 & n41287 ;
  assign n41289 = \m1_addr_i[3]_pad  & ~n13467 ;
  assign n41290 = n13475 & n41289 ;
  assign n41291 = ~n41288 & ~n41290 ;
  assign n41292 = \m0_addr_i[3]_pad  & n13467 ;
  assign n41293 = n13475 & n41292 ;
  assign n41294 = \m7_addr_i[3]_pad  & ~n13467 ;
  assign n41295 = n13492 & n41294 ;
  assign n41296 = ~n41293 & ~n41295 ;
  assign n41297 = n41291 & n41296 ;
  assign n41298 = n41286 & n41297 ;
  assign n41299 = \m3_addr_i[4]_pad  & ~n13467 ;
  assign n41300 = n13484 & n41299 ;
  assign n41301 = \m4_addr_i[4]_pad  & n13467 ;
  assign n41302 = n13460 & n41301 ;
  assign n41303 = ~n41300 & ~n41302 ;
  assign n41304 = \m6_addr_i[4]_pad  & n13467 ;
  assign n41305 = n13492 & n41304 ;
  assign n41306 = \m2_addr_i[4]_pad  & n13467 ;
  assign n41307 = n13484 & n41306 ;
  assign n41308 = ~n41305 & ~n41307 ;
  assign n41309 = n41303 & n41308 ;
  assign n41310 = \m5_addr_i[4]_pad  & ~n13467 ;
  assign n41311 = n13460 & n41310 ;
  assign n41312 = \m1_addr_i[4]_pad  & ~n13467 ;
  assign n41313 = n13475 & n41312 ;
  assign n41314 = ~n41311 & ~n41313 ;
  assign n41315 = \m0_addr_i[4]_pad  & n13467 ;
  assign n41316 = n13475 & n41315 ;
  assign n41317 = \m7_addr_i[4]_pad  & ~n13467 ;
  assign n41318 = n13492 & n41317 ;
  assign n41319 = ~n41316 & ~n41318 ;
  assign n41320 = n41314 & n41319 ;
  assign n41321 = n41309 & n41320 ;
  assign n41322 = \m3_addr_i[5]_pad  & ~n13467 ;
  assign n41323 = n13484 & n41322 ;
  assign n41324 = \m4_addr_i[5]_pad  & n13467 ;
  assign n41325 = n13460 & n41324 ;
  assign n41326 = ~n41323 & ~n41325 ;
  assign n41327 = \m6_addr_i[5]_pad  & n13467 ;
  assign n41328 = n13492 & n41327 ;
  assign n41329 = \m2_addr_i[5]_pad  & n13467 ;
  assign n41330 = n13484 & n41329 ;
  assign n41331 = ~n41328 & ~n41330 ;
  assign n41332 = n41326 & n41331 ;
  assign n41333 = \m5_addr_i[5]_pad  & ~n13467 ;
  assign n41334 = n13460 & n41333 ;
  assign n41335 = \m1_addr_i[5]_pad  & ~n13467 ;
  assign n41336 = n13475 & n41335 ;
  assign n41337 = ~n41334 & ~n41336 ;
  assign n41338 = \m0_addr_i[5]_pad  & n13467 ;
  assign n41339 = n13475 & n41338 ;
  assign n41340 = \m7_addr_i[5]_pad  & ~n13467 ;
  assign n41341 = n13492 & n41340 ;
  assign n41342 = ~n41339 & ~n41341 ;
  assign n41343 = n41337 & n41342 ;
  assign n41344 = n41332 & n41343 ;
  assign n41345 = \m3_addr_i[6]_pad  & ~n13467 ;
  assign n41346 = n13484 & n41345 ;
  assign n41347 = \m4_addr_i[6]_pad  & n13467 ;
  assign n41348 = n13460 & n41347 ;
  assign n41349 = ~n41346 & ~n41348 ;
  assign n41350 = \m6_addr_i[6]_pad  & n13467 ;
  assign n41351 = n13492 & n41350 ;
  assign n41352 = \m2_addr_i[6]_pad  & n13467 ;
  assign n41353 = n13484 & n41352 ;
  assign n41354 = ~n41351 & ~n41353 ;
  assign n41355 = n41349 & n41354 ;
  assign n41356 = \m5_addr_i[6]_pad  & ~n13467 ;
  assign n41357 = n13460 & n41356 ;
  assign n41358 = \m1_addr_i[6]_pad  & ~n13467 ;
  assign n41359 = n13475 & n41358 ;
  assign n41360 = ~n41357 & ~n41359 ;
  assign n41361 = \m0_addr_i[6]_pad  & n13467 ;
  assign n41362 = n13475 & n41361 ;
  assign n41363 = \m7_addr_i[6]_pad  & ~n13467 ;
  assign n41364 = n13492 & n41363 ;
  assign n41365 = ~n41362 & ~n41364 ;
  assign n41366 = n41360 & n41365 ;
  assign n41367 = n41355 & n41366 ;
  assign n41368 = \m3_addr_i[7]_pad  & ~n13467 ;
  assign n41369 = n13484 & n41368 ;
  assign n41370 = \m4_addr_i[7]_pad  & n13467 ;
  assign n41371 = n13460 & n41370 ;
  assign n41372 = ~n41369 & ~n41371 ;
  assign n41373 = \m6_addr_i[7]_pad  & n13467 ;
  assign n41374 = n13492 & n41373 ;
  assign n41375 = \m2_addr_i[7]_pad  & n13467 ;
  assign n41376 = n13484 & n41375 ;
  assign n41377 = ~n41374 & ~n41376 ;
  assign n41378 = n41372 & n41377 ;
  assign n41379 = \m5_addr_i[7]_pad  & ~n13467 ;
  assign n41380 = n13460 & n41379 ;
  assign n41381 = \m1_addr_i[7]_pad  & ~n13467 ;
  assign n41382 = n13475 & n41381 ;
  assign n41383 = ~n41380 & ~n41382 ;
  assign n41384 = \m0_addr_i[7]_pad  & n13467 ;
  assign n41385 = n13475 & n41384 ;
  assign n41386 = \m7_addr_i[7]_pad  & ~n13467 ;
  assign n41387 = n13492 & n41386 ;
  assign n41388 = ~n41385 & ~n41387 ;
  assign n41389 = n41383 & n41388 ;
  assign n41390 = n41378 & n41389 ;
  assign n41391 = \m3_addr_i[8]_pad  & ~n13467 ;
  assign n41392 = n13484 & n41391 ;
  assign n41393 = \m4_addr_i[8]_pad  & n13467 ;
  assign n41394 = n13460 & n41393 ;
  assign n41395 = ~n41392 & ~n41394 ;
  assign n41396 = \m6_addr_i[8]_pad  & n13467 ;
  assign n41397 = n13492 & n41396 ;
  assign n41398 = \m2_addr_i[8]_pad  & n13467 ;
  assign n41399 = n13484 & n41398 ;
  assign n41400 = ~n41397 & ~n41399 ;
  assign n41401 = n41395 & n41400 ;
  assign n41402 = \m5_addr_i[8]_pad  & ~n13467 ;
  assign n41403 = n13460 & n41402 ;
  assign n41404 = \m1_addr_i[8]_pad  & ~n13467 ;
  assign n41405 = n13475 & n41404 ;
  assign n41406 = ~n41403 & ~n41405 ;
  assign n41407 = \m0_addr_i[8]_pad  & n13467 ;
  assign n41408 = n13475 & n41407 ;
  assign n41409 = \m7_addr_i[8]_pad  & ~n13467 ;
  assign n41410 = n13492 & n41409 ;
  assign n41411 = ~n41408 & ~n41410 ;
  assign n41412 = n41406 & n41411 ;
  assign n41413 = n41401 & n41412 ;
  assign n41414 = \m3_addr_i[9]_pad  & ~n13467 ;
  assign n41415 = n13484 & n41414 ;
  assign n41416 = \m4_addr_i[9]_pad  & n13467 ;
  assign n41417 = n13460 & n41416 ;
  assign n41418 = ~n41415 & ~n41417 ;
  assign n41419 = \m6_addr_i[9]_pad  & n13467 ;
  assign n41420 = n13492 & n41419 ;
  assign n41421 = \m2_addr_i[9]_pad  & n13467 ;
  assign n41422 = n13484 & n41421 ;
  assign n41423 = ~n41420 & ~n41422 ;
  assign n41424 = n41418 & n41423 ;
  assign n41425 = \m5_addr_i[9]_pad  & ~n13467 ;
  assign n41426 = n13460 & n41425 ;
  assign n41427 = \m1_addr_i[9]_pad  & ~n13467 ;
  assign n41428 = n13475 & n41427 ;
  assign n41429 = ~n41426 & ~n41428 ;
  assign n41430 = \m0_addr_i[9]_pad  & n13467 ;
  assign n41431 = n13475 & n41430 ;
  assign n41432 = \m7_addr_i[9]_pad  & ~n13467 ;
  assign n41433 = n13492 & n41432 ;
  assign n41434 = ~n41431 & ~n41433 ;
  assign n41435 = n41429 & n41434 ;
  assign n41436 = n41424 & n41435 ;
  assign n41437 = \m3_data_i[0]_pad  & ~n13467 ;
  assign n41438 = n13484 & n41437 ;
  assign n41439 = \m4_data_i[0]_pad  & n13467 ;
  assign n41440 = n13460 & n41439 ;
  assign n41441 = ~n41438 & ~n41440 ;
  assign n41442 = \m6_data_i[0]_pad  & n13467 ;
  assign n41443 = n13492 & n41442 ;
  assign n41444 = \m2_data_i[0]_pad  & n13467 ;
  assign n41445 = n13484 & n41444 ;
  assign n41446 = ~n41443 & ~n41445 ;
  assign n41447 = n41441 & n41446 ;
  assign n41448 = \m5_data_i[0]_pad  & ~n13467 ;
  assign n41449 = n13460 & n41448 ;
  assign n41450 = \m1_data_i[0]_pad  & ~n13467 ;
  assign n41451 = n13475 & n41450 ;
  assign n41452 = ~n41449 & ~n41451 ;
  assign n41453 = \m0_data_i[0]_pad  & n13467 ;
  assign n41454 = n13475 & n41453 ;
  assign n41455 = \m7_data_i[0]_pad  & ~n13467 ;
  assign n41456 = n13492 & n41455 ;
  assign n41457 = ~n41454 & ~n41456 ;
  assign n41458 = n41452 & n41457 ;
  assign n41459 = n41447 & n41458 ;
  assign n41460 = \m3_data_i[10]_pad  & ~n13467 ;
  assign n41461 = n13484 & n41460 ;
  assign n41462 = \m4_data_i[10]_pad  & n13467 ;
  assign n41463 = n13460 & n41462 ;
  assign n41464 = ~n41461 & ~n41463 ;
  assign n41465 = \m6_data_i[10]_pad  & n13467 ;
  assign n41466 = n13492 & n41465 ;
  assign n41467 = \m2_data_i[10]_pad  & n13467 ;
  assign n41468 = n13484 & n41467 ;
  assign n41469 = ~n41466 & ~n41468 ;
  assign n41470 = n41464 & n41469 ;
  assign n41471 = \m5_data_i[10]_pad  & ~n13467 ;
  assign n41472 = n13460 & n41471 ;
  assign n41473 = \m1_data_i[10]_pad  & ~n13467 ;
  assign n41474 = n13475 & n41473 ;
  assign n41475 = ~n41472 & ~n41474 ;
  assign n41476 = \m0_data_i[10]_pad  & n13467 ;
  assign n41477 = n13475 & n41476 ;
  assign n41478 = \m7_data_i[10]_pad  & ~n13467 ;
  assign n41479 = n13492 & n41478 ;
  assign n41480 = ~n41477 & ~n41479 ;
  assign n41481 = n41475 & n41480 ;
  assign n41482 = n41470 & n41481 ;
  assign n41483 = \m3_data_i[11]_pad  & ~n13467 ;
  assign n41484 = n13484 & n41483 ;
  assign n41485 = \m4_data_i[11]_pad  & n13467 ;
  assign n41486 = n13460 & n41485 ;
  assign n41487 = ~n41484 & ~n41486 ;
  assign n41488 = \m6_data_i[11]_pad  & n13467 ;
  assign n41489 = n13492 & n41488 ;
  assign n41490 = \m2_data_i[11]_pad  & n13467 ;
  assign n41491 = n13484 & n41490 ;
  assign n41492 = ~n41489 & ~n41491 ;
  assign n41493 = n41487 & n41492 ;
  assign n41494 = \m5_data_i[11]_pad  & ~n13467 ;
  assign n41495 = n13460 & n41494 ;
  assign n41496 = \m1_data_i[11]_pad  & ~n13467 ;
  assign n41497 = n13475 & n41496 ;
  assign n41498 = ~n41495 & ~n41497 ;
  assign n41499 = \m0_data_i[11]_pad  & n13467 ;
  assign n41500 = n13475 & n41499 ;
  assign n41501 = \m7_data_i[11]_pad  & ~n13467 ;
  assign n41502 = n13492 & n41501 ;
  assign n41503 = ~n41500 & ~n41502 ;
  assign n41504 = n41498 & n41503 ;
  assign n41505 = n41493 & n41504 ;
  assign n41506 = \m3_data_i[12]_pad  & ~n13467 ;
  assign n41507 = n13484 & n41506 ;
  assign n41508 = \m4_data_i[12]_pad  & n13467 ;
  assign n41509 = n13460 & n41508 ;
  assign n41510 = ~n41507 & ~n41509 ;
  assign n41511 = \m6_data_i[12]_pad  & n13467 ;
  assign n41512 = n13492 & n41511 ;
  assign n41513 = \m2_data_i[12]_pad  & n13467 ;
  assign n41514 = n13484 & n41513 ;
  assign n41515 = ~n41512 & ~n41514 ;
  assign n41516 = n41510 & n41515 ;
  assign n41517 = \m5_data_i[12]_pad  & ~n13467 ;
  assign n41518 = n13460 & n41517 ;
  assign n41519 = \m1_data_i[12]_pad  & ~n13467 ;
  assign n41520 = n13475 & n41519 ;
  assign n41521 = ~n41518 & ~n41520 ;
  assign n41522 = \m0_data_i[12]_pad  & n13467 ;
  assign n41523 = n13475 & n41522 ;
  assign n41524 = \m7_data_i[12]_pad  & ~n13467 ;
  assign n41525 = n13492 & n41524 ;
  assign n41526 = ~n41523 & ~n41525 ;
  assign n41527 = n41521 & n41526 ;
  assign n41528 = n41516 & n41527 ;
  assign n41529 = \m3_data_i[13]_pad  & ~n13467 ;
  assign n41530 = n13484 & n41529 ;
  assign n41531 = \m4_data_i[13]_pad  & n13467 ;
  assign n41532 = n13460 & n41531 ;
  assign n41533 = ~n41530 & ~n41532 ;
  assign n41534 = \m6_data_i[13]_pad  & n13467 ;
  assign n41535 = n13492 & n41534 ;
  assign n41536 = \m2_data_i[13]_pad  & n13467 ;
  assign n41537 = n13484 & n41536 ;
  assign n41538 = ~n41535 & ~n41537 ;
  assign n41539 = n41533 & n41538 ;
  assign n41540 = \m5_data_i[13]_pad  & ~n13467 ;
  assign n41541 = n13460 & n41540 ;
  assign n41542 = \m1_data_i[13]_pad  & ~n13467 ;
  assign n41543 = n13475 & n41542 ;
  assign n41544 = ~n41541 & ~n41543 ;
  assign n41545 = \m0_data_i[13]_pad  & n13467 ;
  assign n41546 = n13475 & n41545 ;
  assign n41547 = \m7_data_i[13]_pad  & ~n13467 ;
  assign n41548 = n13492 & n41547 ;
  assign n41549 = ~n41546 & ~n41548 ;
  assign n41550 = n41544 & n41549 ;
  assign n41551 = n41539 & n41550 ;
  assign n41552 = \m3_data_i[14]_pad  & ~n13467 ;
  assign n41553 = n13484 & n41552 ;
  assign n41554 = \m4_data_i[14]_pad  & n13467 ;
  assign n41555 = n13460 & n41554 ;
  assign n41556 = ~n41553 & ~n41555 ;
  assign n41557 = \m6_data_i[14]_pad  & n13467 ;
  assign n41558 = n13492 & n41557 ;
  assign n41559 = \m2_data_i[14]_pad  & n13467 ;
  assign n41560 = n13484 & n41559 ;
  assign n41561 = ~n41558 & ~n41560 ;
  assign n41562 = n41556 & n41561 ;
  assign n41563 = \m5_data_i[14]_pad  & ~n13467 ;
  assign n41564 = n13460 & n41563 ;
  assign n41565 = \m1_data_i[14]_pad  & ~n13467 ;
  assign n41566 = n13475 & n41565 ;
  assign n41567 = ~n41564 & ~n41566 ;
  assign n41568 = \m0_data_i[14]_pad  & n13467 ;
  assign n41569 = n13475 & n41568 ;
  assign n41570 = \m7_data_i[14]_pad  & ~n13467 ;
  assign n41571 = n13492 & n41570 ;
  assign n41572 = ~n41569 & ~n41571 ;
  assign n41573 = n41567 & n41572 ;
  assign n41574 = n41562 & n41573 ;
  assign n41575 = \m3_data_i[15]_pad  & ~n13467 ;
  assign n41576 = n13484 & n41575 ;
  assign n41577 = \m4_data_i[15]_pad  & n13467 ;
  assign n41578 = n13460 & n41577 ;
  assign n41579 = ~n41576 & ~n41578 ;
  assign n41580 = \m6_data_i[15]_pad  & n13467 ;
  assign n41581 = n13492 & n41580 ;
  assign n41582 = \m2_data_i[15]_pad  & n13467 ;
  assign n41583 = n13484 & n41582 ;
  assign n41584 = ~n41581 & ~n41583 ;
  assign n41585 = n41579 & n41584 ;
  assign n41586 = \m5_data_i[15]_pad  & ~n13467 ;
  assign n41587 = n13460 & n41586 ;
  assign n41588 = \m1_data_i[15]_pad  & ~n13467 ;
  assign n41589 = n13475 & n41588 ;
  assign n41590 = ~n41587 & ~n41589 ;
  assign n41591 = \m0_data_i[15]_pad  & n13467 ;
  assign n41592 = n13475 & n41591 ;
  assign n41593 = \m7_data_i[15]_pad  & ~n13467 ;
  assign n41594 = n13492 & n41593 ;
  assign n41595 = ~n41592 & ~n41594 ;
  assign n41596 = n41590 & n41595 ;
  assign n41597 = n41585 & n41596 ;
  assign n41598 = \m3_data_i[16]_pad  & ~n13467 ;
  assign n41599 = n13484 & n41598 ;
  assign n41600 = \m4_data_i[16]_pad  & n13467 ;
  assign n41601 = n13460 & n41600 ;
  assign n41602 = ~n41599 & ~n41601 ;
  assign n41603 = \m6_data_i[16]_pad  & n13467 ;
  assign n41604 = n13492 & n41603 ;
  assign n41605 = \m2_data_i[16]_pad  & n13467 ;
  assign n41606 = n13484 & n41605 ;
  assign n41607 = ~n41604 & ~n41606 ;
  assign n41608 = n41602 & n41607 ;
  assign n41609 = \m5_data_i[16]_pad  & ~n13467 ;
  assign n41610 = n13460 & n41609 ;
  assign n41611 = \m1_data_i[16]_pad  & ~n13467 ;
  assign n41612 = n13475 & n41611 ;
  assign n41613 = ~n41610 & ~n41612 ;
  assign n41614 = \m0_data_i[16]_pad  & n13467 ;
  assign n41615 = n13475 & n41614 ;
  assign n41616 = \m7_data_i[16]_pad  & ~n13467 ;
  assign n41617 = n13492 & n41616 ;
  assign n41618 = ~n41615 & ~n41617 ;
  assign n41619 = n41613 & n41618 ;
  assign n41620 = n41608 & n41619 ;
  assign n41621 = \m3_data_i[17]_pad  & ~n13467 ;
  assign n41622 = n13484 & n41621 ;
  assign n41623 = \m4_data_i[17]_pad  & n13467 ;
  assign n41624 = n13460 & n41623 ;
  assign n41625 = ~n41622 & ~n41624 ;
  assign n41626 = \m6_data_i[17]_pad  & n13467 ;
  assign n41627 = n13492 & n41626 ;
  assign n41628 = \m2_data_i[17]_pad  & n13467 ;
  assign n41629 = n13484 & n41628 ;
  assign n41630 = ~n41627 & ~n41629 ;
  assign n41631 = n41625 & n41630 ;
  assign n41632 = \m5_data_i[17]_pad  & ~n13467 ;
  assign n41633 = n13460 & n41632 ;
  assign n41634 = \m1_data_i[17]_pad  & ~n13467 ;
  assign n41635 = n13475 & n41634 ;
  assign n41636 = ~n41633 & ~n41635 ;
  assign n41637 = \m0_data_i[17]_pad  & n13467 ;
  assign n41638 = n13475 & n41637 ;
  assign n41639 = \m7_data_i[17]_pad  & ~n13467 ;
  assign n41640 = n13492 & n41639 ;
  assign n41641 = ~n41638 & ~n41640 ;
  assign n41642 = n41636 & n41641 ;
  assign n41643 = n41631 & n41642 ;
  assign n41644 = \m3_data_i[18]_pad  & ~n13467 ;
  assign n41645 = n13484 & n41644 ;
  assign n41646 = \m4_data_i[18]_pad  & n13467 ;
  assign n41647 = n13460 & n41646 ;
  assign n41648 = ~n41645 & ~n41647 ;
  assign n41649 = \m6_data_i[18]_pad  & n13467 ;
  assign n41650 = n13492 & n41649 ;
  assign n41651 = \m2_data_i[18]_pad  & n13467 ;
  assign n41652 = n13484 & n41651 ;
  assign n41653 = ~n41650 & ~n41652 ;
  assign n41654 = n41648 & n41653 ;
  assign n41655 = \m5_data_i[18]_pad  & ~n13467 ;
  assign n41656 = n13460 & n41655 ;
  assign n41657 = \m1_data_i[18]_pad  & ~n13467 ;
  assign n41658 = n13475 & n41657 ;
  assign n41659 = ~n41656 & ~n41658 ;
  assign n41660 = \m0_data_i[18]_pad  & n13467 ;
  assign n41661 = n13475 & n41660 ;
  assign n41662 = \m7_data_i[18]_pad  & ~n13467 ;
  assign n41663 = n13492 & n41662 ;
  assign n41664 = ~n41661 & ~n41663 ;
  assign n41665 = n41659 & n41664 ;
  assign n41666 = n41654 & n41665 ;
  assign n41667 = \m3_data_i[19]_pad  & ~n13467 ;
  assign n41668 = n13484 & n41667 ;
  assign n41669 = \m4_data_i[19]_pad  & n13467 ;
  assign n41670 = n13460 & n41669 ;
  assign n41671 = ~n41668 & ~n41670 ;
  assign n41672 = \m6_data_i[19]_pad  & n13467 ;
  assign n41673 = n13492 & n41672 ;
  assign n41674 = \m2_data_i[19]_pad  & n13467 ;
  assign n41675 = n13484 & n41674 ;
  assign n41676 = ~n41673 & ~n41675 ;
  assign n41677 = n41671 & n41676 ;
  assign n41678 = \m5_data_i[19]_pad  & ~n13467 ;
  assign n41679 = n13460 & n41678 ;
  assign n41680 = \m1_data_i[19]_pad  & ~n13467 ;
  assign n41681 = n13475 & n41680 ;
  assign n41682 = ~n41679 & ~n41681 ;
  assign n41683 = \m0_data_i[19]_pad  & n13467 ;
  assign n41684 = n13475 & n41683 ;
  assign n41685 = \m7_data_i[19]_pad  & ~n13467 ;
  assign n41686 = n13492 & n41685 ;
  assign n41687 = ~n41684 & ~n41686 ;
  assign n41688 = n41682 & n41687 ;
  assign n41689 = n41677 & n41688 ;
  assign n41690 = \m3_data_i[1]_pad  & ~n13467 ;
  assign n41691 = n13484 & n41690 ;
  assign n41692 = \m4_data_i[1]_pad  & n13467 ;
  assign n41693 = n13460 & n41692 ;
  assign n41694 = ~n41691 & ~n41693 ;
  assign n41695 = \m6_data_i[1]_pad  & n13467 ;
  assign n41696 = n13492 & n41695 ;
  assign n41697 = \m2_data_i[1]_pad  & n13467 ;
  assign n41698 = n13484 & n41697 ;
  assign n41699 = ~n41696 & ~n41698 ;
  assign n41700 = n41694 & n41699 ;
  assign n41701 = \m5_data_i[1]_pad  & ~n13467 ;
  assign n41702 = n13460 & n41701 ;
  assign n41703 = \m1_data_i[1]_pad  & ~n13467 ;
  assign n41704 = n13475 & n41703 ;
  assign n41705 = ~n41702 & ~n41704 ;
  assign n41706 = \m0_data_i[1]_pad  & n13467 ;
  assign n41707 = n13475 & n41706 ;
  assign n41708 = \m7_data_i[1]_pad  & ~n13467 ;
  assign n41709 = n13492 & n41708 ;
  assign n41710 = ~n41707 & ~n41709 ;
  assign n41711 = n41705 & n41710 ;
  assign n41712 = n41700 & n41711 ;
  assign n41713 = \m3_data_i[20]_pad  & ~n13467 ;
  assign n41714 = n13484 & n41713 ;
  assign n41715 = \m4_data_i[20]_pad  & n13467 ;
  assign n41716 = n13460 & n41715 ;
  assign n41717 = ~n41714 & ~n41716 ;
  assign n41718 = \m6_data_i[20]_pad  & n13467 ;
  assign n41719 = n13492 & n41718 ;
  assign n41720 = \m2_data_i[20]_pad  & n13467 ;
  assign n41721 = n13484 & n41720 ;
  assign n41722 = ~n41719 & ~n41721 ;
  assign n41723 = n41717 & n41722 ;
  assign n41724 = \m5_data_i[20]_pad  & ~n13467 ;
  assign n41725 = n13460 & n41724 ;
  assign n41726 = \m1_data_i[20]_pad  & ~n13467 ;
  assign n41727 = n13475 & n41726 ;
  assign n41728 = ~n41725 & ~n41727 ;
  assign n41729 = \m0_data_i[20]_pad  & n13467 ;
  assign n41730 = n13475 & n41729 ;
  assign n41731 = \m7_data_i[20]_pad  & ~n13467 ;
  assign n41732 = n13492 & n41731 ;
  assign n41733 = ~n41730 & ~n41732 ;
  assign n41734 = n41728 & n41733 ;
  assign n41735 = n41723 & n41734 ;
  assign n41736 = \m3_data_i[21]_pad  & ~n13467 ;
  assign n41737 = n13484 & n41736 ;
  assign n41738 = \m4_data_i[21]_pad  & n13467 ;
  assign n41739 = n13460 & n41738 ;
  assign n41740 = ~n41737 & ~n41739 ;
  assign n41741 = \m6_data_i[21]_pad  & n13467 ;
  assign n41742 = n13492 & n41741 ;
  assign n41743 = \m2_data_i[21]_pad  & n13467 ;
  assign n41744 = n13484 & n41743 ;
  assign n41745 = ~n41742 & ~n41744 ;
  assign n41746 = n41740 & n41745 ;
  assign n41747 = \m5_data_i[21]_pad  & ~n13467 ;
  assign n41748 = n13460 & n41747 ;
  assign n41749 = \m1_data_i[21]_pad  & ~n13467 ;
  assign n41750 = n13475 & n41749 ;
  assign n41751 = ~n41748 & ~n41750 ;
  assign n41752 = \m0_data_i[21]_pad  & n13467 ;
  assign n41753 = n13475 & n41752 ;
  assign n41754 = \m7_data_i[21]_pad  & ~n13467 ;
  assign n41755 = n13492 & n41754 ;
  assign n41756 = ~n41753 & ~n41755 ;
  assign n41757 = n41751 & n41756 ;
  assign n41758 = n41746 & n41757 ;
  assign n41759 = \m3_data_i[22]_pad  & ~n13467 ;
  assign n41760 = n13484 & n41759 ;
  assign n41761 = \m4_data_i[22]_pad  & n13467 ;
  assign n41762 = n13460 & n41761 ;
  assign n41763 = ~n41760 & ~n41762 ;
  assign n41764 = \m6_data_i[22]_pad  & n13467 ;
  assign n41765 = n13492 & n41764 ;
  assign n41766 = \m2_data_i[22]_pad  & n13467 ;
  assign n41767 = n13484 & n41766 ;
  assign n41768 = ~n41765 & ~n41767 ;
  assign n41769 = n41763 & n41768 ;
  assign n41770 = \m5_data_i[22]_pad  & ~n13467 ;
  assign n41771 = n13460 & n41770 ;
  assign n41772 = \m1_data_i[22]_pad  & ~n13467 ;
  assign n41773 = n13475 & n41772 ;
  assign n41774 = ~n41771 & ~n41773 ;
  assign n41775 = \m0_data_i[22]_pad  & n13467 ;
  assign n41776 = n13475 & n41775 ;
  assign n41777 = \m7_data_i[22]_pad  & ~n13467 ;
  assign n41778 = n13492 & n41777 ;
  assign n41779 = ~n41776 & ~n41778 ;
  assign n41780 = n41774 & n41779 ;
  assign n41781 = n41769 & n41780 ;
  assign n41782 = \m3_data_i[23]_pad  & ~n13467 ;
  assign n41783 = n13484 & n41782 ;
  assign n41784 = \m4_data_i[23]_pad  & n13467 ;
  assign n41785 = n13460 & n41784 ;
  assign n41786 = ~n41783 & ~n41785 ;
  assign n41787 = \m6_data_i[23]_pad  & n13467 ;
  assign n41788 = n13492 & n41787 ;
  assign n41789 = \m2_data_i[23]_pad  & n13467 ;
  assign n41790 = n13484 & n41789 ;
  assign n41791 = ~n41788 & ~n41790 ;
  assign n41792 = n41786 & n41791 ;
  assign n41793 = \m5_data_i[23]_pad  & ~n13467 ;
  assign n41794 = n13460 & n41793 ;
  assign n41795 = \m1_data_i[23]_pad  & ~n13467 ;
  assign n41796 = n13475 & n41795 ;
  assign n41797 = ~n41794 & ~n41796 ;
  assign n41798 = \m0_data_i[23]_pad  & n13467 ;
  assign n41799 = n13475 & n41798 ;
  assign n41800 = \m7_data_i[23]_pad  & ~n13467 ;
  assign n41801 = n13492 & n41800 ;
  assign n41802 = ~n41799 & ~n41801 ;
  assign n41803 = n41797 & n41802 ;
  assign n41804 = n41792 & n41803 ;
  assign n41805 = \m3_data_i[24]_pad  & ~n13467 ;
  assign n41806 = n13484 & n41805 ;
  assign n41807 = \m4_data_i[24]_pad  & n13467 ;
  assign n41808 = n13460 & n41807 ;
  assign n41809 = ~n41806 & ~n41808 ;
  assign n41810 = \m6_data_i[24]_pad  & n13467 ;
  assign n41811 = n13492 & n41810 ;
  assign n41812 = \m2_data_i[24]_pad  & n13467 ;
  assign n41813 = n13484 & n41812 ;
  assign n41814 = ~n41811 & ~n41813 ;
  assign n41815 = n41809 & n41814 ;
  assign n41816 = \m5_data_i[24]_pad  & ~n13467 ;
  assign n41817 = n13460 & n41816 ;
  assign n41818 = \m1_data_i[24]_pad  & ~n13467 ;
  assign n41819 = n13475 & n41818 ;
  assign n41820 = ~n41817 & ~n41819 ;
  assign n41821 = \m0_data_i[24]_pad  & n13467 ;
  assign n41822 = n13475 & n41821 ;
  assign n41823 = \m7_data_i[24]_pad  & ~n13467 ;
  assign n41824 = n13492 & n41823 ;
  assign n41825 = ~n41822 & ~n41824 ;
  assign n41826 = n41820 & n41825 ;
  assign n41827 = n41815 & n41826 ;
  assign n41828 = \m3_data_i[25]_pad  & ~n13467 ;
  assign n41829 = n13484 & n41828 ;
  assign n41830 = \m4_data_i[25]_pad  & n13467 ;
  assign n41831 = n13460 & n41830 ;
  assign n41832 = ~n41829 & ~n41831 ;
  assign n41833 = \m6_data_i[25]_pad  & n13467 ;
  assign n41834 = n13492 & n41833 ;
  assign n41835 = \m2_data_i[25]_pad  & n13467 ;
  assign n41836 = n13484 & n41835 ;
  assign n41837 = ~n41834 & ~n41836 ;
  assign n41838 = n41832 & n41837 ;
  assign n41839 = \m5_data_i[25]_pad  & ~n13467 ;
  assign n41840 = n13460 & n41839 ;
  assign n41841 = \m1_data_i[25]_pad  & ~n13467 ;
  assign n41842 = n13475 & n41841 ;
  assign n41843 = ~n41840 & ~n41842 ;
  assign n41844 = \m0_data_i[25]_pad  & n13467 ;
  assign n41845 = n13475 & n41844 ;
  assign n41846 = \m7_data_i[25]_pad  & ~n13467 ;
  assign n41847 = n13492 & n41846 ;
  assign n41848 = ~n41845 & ~n41847 ;
  assign n41849 = n41843 & n41848 ;
  assign n41850 = n41838 & n41849 ;
  assign n41851 = \m3_data_i[26]_pad  & ~n13467 ;
  assign n41852 = n13484 & n41851 ;
  assign n41853 = \m4_data_i[26]_pad  & n13467 ;
  assign n41854 = n13460 & n41853 ;
  assign n41855 = ~n41852 & ~n41854 ;
  assign n41856 = \m6_data_i[26]_pad  & n13467 ;
  assign n41857 = n13492 & n41856 ;
  assign n41858 = \m2_data_i[26]_pad  & n13467 ;
  assign n41859 = n13484 & n41858 ;
  assign n41860 = ~n41857 & ~n41859 ;
  assign n41861 = n41855 & n41860 ;
  assign n41862 = \m5_data_i[26]_pad  & ~n13467 ;
  assign n41863 = n13460 & n41862 ;
  assign n41864 = \m1_data_i[26]_pad  & ~n13467 ;
  assign n41865 = n13475 & n41864 ;
  assign n41866 = ~n41863 & ~n41865 ;
  assign n41867 = \m0_data_i[26]_pad  & n13467 ;
  assign n41868 = n13475 & n41867 ;
  assign n41869 = \m7_data_i[26]_pad  & ~n13467 ;
  assign n41870 = n13492 & n41869 ;
  assign n41871 = ~n41868 & ~n41870 ;
  assign n41872 = n41866 & n41871 ;
  assign n41873 = n41861 & n41872 ;
  assign n41874 = \m3_data_i[27]_pad  & ~n13467 ;
  assign n41875 = n13484 & n41874 ;
  assign n41876 = \m4_data_i[27]_pad  & n13467 ;
  assign n41877 = n13460 & n41876 ;
  assign n41878 = ~n41875 & ~n41877 ;
  assign n41879 = \m6_data_i[27]_pad  & n13467 ;
  assign n41880 = n13492 & n41879 ;
  assign n41881 = \m2_data_i[27]_pad  & n13467 ;
  assign n41882 = n13484 & n41881 ;
  assign n41883 = ~n41880 & ~n41882 ;
  assign n41884 = n41878 & n41883 ;
  assign n41885 = \m5_data_i[27]_pad  & ~n13467 ;
  assign n41886 = n13460 & n41885 ;
  assign n41887 = \m1_data_i[27]_pad  & ~n13467 ;
  assign n41888 = n13475 & n41887 ;
  assign n41889 = ~n41886 & ~n41888 ;
  assign n41890 = \m0_data_i[27]_pad  & n13467 ;
  assign n41891 = n13475 & n41890 ;
  assign n41892 = \m7_data_i[27]_pad  & ~n13467 ;
  assign n41893 = n13492 & n41892 ;
  assign n41894 = ~n41891 & ~n41893 ;
  assign n41895 = n41889 & n41894 ;
  assign n41896 = n41884 & n41895 ;
  assign n41897 = \m3_data_i[28]_pad  & ~n13467 ;
  assign n41898 = n13484 & n41897 ;
  assign n41899 = \m4_data_i[28]_pad  & n13467 ;
  assign n41900 = n13460 & n41899 ;
  assign n41901 = ~n41898 & ~n41900 ;
  assign n41902 = \m6_data_i[28]_pad  & n13467 ;
  assign n41903 = n13492 & n41902 ;
  assign n41904 = \m2_data_i[28]_pad  & n13467 ;
  assign n41905 = n13484 & n41904 ;
  assign n41906 = ~n41903 & ~n41905 ;
  assign n41907 = n41901 & n41906 ;
  assign n41908 = \m5_data_i[28]_pad  & ~n13467 ;
  assign n41909 = n13460 & n41908 ;
  assign n41910 = \m1_data_i[28]_pad  & ~n13467 ;
  assign n41911 = n13475 & n41910 ;
  assign n41912 = ~n41909 & ~n41911 ;
  assign n41913 = \m0_data_i[28]_pad  & n13467 ;
  assign n41914 = n13475 & n41913 ;
  assign n41915 = \m7_data_i[28]_pad  & ~n13467 ;
  assign n41916 = n13492 & n41915 ;
  assign n41917 = ~n41914 & ~n41916 ;
  assign n41918 = n41912 & n41917 ;
  assign n41919 = n41907 & n41918 ;
  assign n41920 = \m3_data_i[29]_pad  & ~n13467 ;
  assign n41921 = n13484 & n41920 ;
  assign n41922 = \m4_data_i[29]_pad  & n13467 ;
  assign n41923 = n13460 & n41922 ;
  assign n41924 = ~n41921 & ~n41923 ;
  assign n41925 = \m6_data_i[29]_pad  & n13467 ;
  assign n41926 = n13492 & n41925 ;
  assign n41927 = \m2_data_i[29]_pad  & n13467 ;
  assign n41928 = n13484 & n41927 ;
  assign n41929 = ~n41926 & ~n41928 ;
  assign n41930 = n41924 & n41929 ;
  assign n41931 = \m5_data_i[29]_pad  & ~n13467 ;
  assign n41932 = n13460 & n41931 ;
  assign n41933 = \m1_data_i[29]_pad  & ~n13467 ;
  assign n41934 = n13475 & n41933 ;
  assign n41935 = ~n41932 & ~n41934 ;
  assign n41936 = \m0_data_i[29]_pad  & n13467 ;
  assign n41937 = n13475 & n41936 ;
  assign n41938 = \m7_data_i[29]_pad  & ~n13467 ;
  assign n41939 = n13492 & n41938 ;
  assign n41940 = ~n41937 & ~n41939 ;
  assign n41941 = n41935 & n41940 ;
  assign n41942 = n41930 & n41941 ;
  assign n41943 = \m3_data_i[2]_pad  & ~n13467 ;
  assign n41944 = n13484 & n41943 ;
  assign n41945 = \m4_data_i[2]_pad  & n13467 ;
  assign n41946 = n13460 & n41945 ;
  assign n41947 = ~n41944 & ~n41946 ;
  assign n41948 = \m6_data_i[2]_pad  & n13467 ;
  assign n41949 = n13492 & n41948 ;
  assign n41950 = \m2_data_i[2]_pad  & n13467 ;
  assign n41951 = n13484 & n41950 ;
  assign n41952 = ~n41949 & ~n41951 ;
  assign n41953 = n41947 & n41952 ;
  assign n41954 = \m5_data_i[2]_pad  & ~n13467 ;
  assign n41955 = n13460 & n41954 ;
  assign n41956 = \m1_data_i[2]_pad  & ~n13467 ;
  assign n41957 = n13475 & n41956 ;
  assign n41958 = ~n41955 & ~n41957 ;
  assign n41959 = \m0_data_i[2]_pad  & n13467 ;
  assign n41960 = n13475 & n41959 ;
  assign n41961 = \m7_data_i[2]_pad  & ~n13467 ;
  assign n41962 = n13492 & n41961 ;
  assign n41963 = ~n41960 & ~n41962 ;
  assign n41964 = n41958 & n41963 ;
  assign n41965 = n41953 & n41964 ;
  assign n41966 = \m3_data_i[30]_pad  & ~n13467 ;
  assign n41967 = n13484 & n41966 ;
  assign n41968 = \m4_data_i[30]_pad  & n13467 ;
  assign n41969 = n13460 & n41968 ;
  assign n41970 = ~n41967 & ~n41969 ;
  assign n41971 = \m6_data_i[30]_pad  & n13467 ;
  assign n41972 = n13492 & n41971 ;
  assign n41973 = \m2_data_i[30]_pad  & n13467 ;
  assign n41974 = n13484 & n41973 ;
  assign n41975 = ~n41972 & ~n41974 ;
  assign n41976 = n41970 & n41975 ;
  assign n41977 = \m5_data_i[30]_pad  & ~n13467 ;
  assign n41978 = n13460 & n41977 ;
  assign n41979 = \m1_data_i[30]_pad  & ~n13467 ;
  assign n41980 = n13475 & n41979 ;
  assign n41981 = ~n41978 & ~n41980 ;
  assign n41982 = \m0_data_i[30]_pad  & n13467 ;
  assign n41983 = n13475 & n41982 ;
  assign n41984 = \m7_data_i[30]_pad  & ~n13467 ;
  assign n41985 = n13492 & n41984 ;
  assign n41986 = ~n41983 & ~n41985 ;
  assign n41987 = n41981 & n41986 ;
  assign n41988 = n41976 & n41987 ;
  assign n41989 = \m3_data_i[31]_pad  & ~n13467 ;
  assign n41990 = n13484 & n41989 ;
  assign n41991 = \m4_data_i[31]_pad  & n13467 ;
  assign n41992 = n13460 & n41991 ;
  assign n41993 = ~n41990 & ~n41992 ;
  assign n41994 = \m6_data_i[31]_pad  & n13467 ;
  assign n41995 = n13492 & n41994 ;
  assign n41996 = \m2_data_i[31]_pad  & n13467 ;
  assign n41997 = n13484 & n41996 ;
  assign n41998 = ~n41995 & ~n41997 ;
  assign n41999 = n41993 & n41998 ;
  assign n42000 = \m5_data_i[31]_pad  & ~n13467 ;
  assign n42001 = n13460 & n42000 ;
  assign n42002 = \m1_data_i[31]_pad  & ~n13467 ;
  assign n42003 = n13475 & n42002 ;
  assign n42004 = ~n42001 & ~n42003 ;
  assign n42005 = \m0_data_i[31]_pad  & n13467 ;
  assign n42006 = n13475 & n42005 ;
  assign n42007 = \m7_data_i[31]_pad  & ~n13467 ;
  assign n42008 = n13492 & n42007 ;
  assign n42009 = ~n42006 & ~n42008 ;
  assign n42010 = n42004 & n42009 ;
  assign n42011 = n41999 & n42010 ;
  assign n42012 = \m3_data_i[3]_pad  & ~n13467 ;
  assign n42013 = n13484 & n42012 ;
  assign n42014 = \m4_data_i[3]_pad  & n13467 ;
  assign n42015 = n13460 & n42014 ;
  assign n42016 = ~n42013 & ~n42015 ;
  assign n42017 = \m6_data_i[3]_pad  & n13467 ;
  assign n42018 = n13492 & n42017 ;
  assign n42019 = \m2_data_i[3]_pad  & n13467 ;
  assign n42020 = n13484 & n42019 ;
  assign n42021 = ~n42018 & ~n42020 ;
  assign n42022 = n42016 & n42021 ;
  assign n42023 = \m5_data_i[3]_pad  & ~n13467 ;
  assign n42024 = n13460 & n42023 ;
  assign n42025 = \m1_data_i[3]_pad  & ~n13467 ;
  assign n42026 = n13475 & n42025 ;
  assign n42027 = ~n42024 & ~n42026 ;
  assign n42028 = \m0_data_i[3]_pad  & n13467 ;
  assign n42029 = n13475 & n42028 ;
  assign n42030 = \m7_data_i[3]_pad  & ~n13467 ;
  assign n42031 = n13492 & n42030 ;
  assign n42032 = ~n42029 & ~n42031 ;
  assign n42033 = n42027 & n42032 ;
  assign n42034 = n42022 & n42033 ;
  assign n42035 = \m3_data_i[4]_pad  & ~n13467 ;
  assign n42036 = n13484 & n42035 ;
  assign n42037 = \m4_data_i[4]_pad  & n13467 ;
  assign n42038 = n13460 & n42037 ;
  assign n42039 = ~n42036 & ~n42038 ;
  assign n42040 = \m6_data_i[4]_pad  & n13467 ;
  assign n42041 = n13492 & n42040 ;
  assign n42042 = \m2_data_i[4]_pad  & n13467 ;
  assign n42043 = n13484 & n42042 ;
  assign n42044 = ~n42041 & ~n42043 ;
  assign n42045 = n42039 & n42044 ;
  assign n42046 = \m5_data_i[4]_pad  & ~n13467 ;
  assign n42047 = n13460 & n42046 ;
  assign n42048 = \m1_data_i[4]_pad  & ~n13467 ;
  assign n42049 = n13475 & n42048 ;
  assign n42050 = ~n42047 & ~n42049 ;
  assign n42051 = \m0_data_i[4]_pad  & n13467 ;
  assign n42052 = n13475 & n42051 ;
  assign n42053 = \m7_data_i[4]_pad  & ~n13467 ;
  assign n42054 = n13492 & n42053 ;
  assign n42055 = ~n42052 & ~n42054 ;
  assign n42056 = n42050 & n42055 ;
  assign n42057 = n42045 & n42056 ;
  assign n42058 = \m3_data_i[5]_pad  & ~n13467 ;
  assign n42059 = n13484 & n42058 ;
  assign n42060 = \m4_data_i[5]_pad  & n13467 ;
  assign n42061 = n13460 & n42060 ;
  assign n42062 = ~n42059 & ~n42061 ;
  assign n42063 = \m6_data_i[5]_pad  & n13467 ;
  assign n42064 = n13492 & n42063 ;
  assign n42065 = \m2_data_i[5]_pad  & n13467 ;
  assign n42066 = n13484 & n42065 ;
  assign n42067 = ~n42064 & ~n42066 ;
  assign n42068 = n42062 & n42067 ;
  assign n42069 = \m5_data_i[5]_pad  & ~n13467 ;
  assign n42070 = n13460 & n42069 ;
  assign n42071 = \m1_data_i[5]_pad  & ~n13467 ;
  assign n42072 = n13475 & n42071 ;
  assign n42073 = ~n42070 & ~n42072 ;
  assign n42074 = \m0_data_i[5]_pad  & n13467 ;
  assign n42075 = n13475 & n42074 ;
  assign n42076 = \m7_data_i[5]_pad  & ~n13467 ;
  assign n42077 = n13492 & n42076 ;
  assign n42078 = ~n42075 & ~n42077 ;
  assign n42079 = n42073 & n42078 ;
  assign n42080 = n42068 & n42079 ;
  assign n42081 = \m3_data_i[6]_pad  & ~n13467 ;
  assign n42082 = n13484 & n42081 ;
  assign n42083 = \m4_data_i[6]_pad  & n13467 ;
  assign n42084 = n13460 & n42083 ;
  assign n42085 = ~n42082 & ~n42084 ;
  assign n42086 = \m6_data_i[6]_pad  & n13467 ;
  assign n42087 = n13492 & n42086 ;
  assign n42088 = \m2_data_i[6]_pad  & n13467 ;
  assign n42089 = n13484 & n42088 ;
  assign n42090 = ~n42087 & ~n42089 ;
  assign n42091 = n42085 & n42090 ;
  assign n42092 = \m5_data_i[6]_pad  & ~n13467 ;
  assign n42093 = n13460 & n42092 ;
  assign n42094 = \m1_data_i[6]_pad  & ~n13467 ;
  assign n42095 = n13475 & n42094 ;
  assign n42096 = ~n42093 & ~n42095 ;
  assign n42097 = \m0_data_i[6]_pad  & n13467 ;
  assign n42098 = n13475 & n42097 ;
  assign n42099 = \m7_data_i[6]_pad  & ~n13467 ;
  assign n42100 = n13492 & n42099 ;
  assign n42101 = ~n42098 & ~n42100 ;
  assign n42102 = n42096 & n42101 ;
  assign n42103 = n42091 & n42102 ;
  assign n42104 = \m3_data_i[7]_pad  & ~n13467 ;
  assign n42105 = n13484 & n42104 ;
  assign n42106 = \m4_data_i[7]_pad  & n13467 ;
  assign n42107 = n13460 & n42106 ;
  assign n42108 = ~n42105 & ~n42107 ;
  assign n42109 = \m6_data_i[7]_pad  & n13467 ;
  assign n42110 = n13492 & n42109 ;
  assign n42111 = \m2_data_i[7]_pad  & n13467 ;
  assign n42112 = n13484 & n42111 ;
  assign n42113 = ~n42110 & ~n42112 ;
  assign n42114 = n42108 & n42113 ;
  assign n42115 = \m5_data_i[7]_pad  & ~n13467 ;
  assign n42116 = n13460 & n42115 ;
  assign n42117 = \m1_data_i[7]_pad  & ~n13467 ;
  assign n42118 = n13475 & n42117 ;
  assign n42119 = ~n42116 & ~n42118 ;
  assign n42120 = \m0_data_i[7]_pad  & n13467 ;
  assign n42121 = n13475 & n42120 ;
  assign n42122 = \m7_data_i[7]_pad  & ~n13467 ;
  assign n42123 = n13492 & n42122 ;
  assign n42124 = ~n42121 & ~n42123 ;
  assign n42125 = n42119 & n42124 ;
  assign n42126 = n42114 & n42125 ;
  assign n42127 = \m3_data_i[8]_pad  & ~n13467 ;
  assign n42128 = n13484 & n42127 ;
  assign n42129 = \m4_data_i[8]_pad  & n13467 ;
  assign n42130 = n13460 & n42129 ;
  assign n42131 = ~n42128 & ~n42130 ;
  assign n42132 = \m6_data_i[8]_pad  & n13467 ;
  assign n42133 = n13492 & n42132 ;
  assign n42134 = \m2_data_i[8]_pad  & n13467 ;
  assign n42135 = n13484 & n42134 ;
  assign n42136 = ~n42133 & ~n42135 ;
  assign n42137 = n42131 & n42136 ;
  assign n42138 = \m5_data_i[8]_pad  & ~n13467 ;
  assign n42139 = n13460 & n42138 ;
  assign n42140 = \m1_data_i[8]_pad  & ~n13467 ;
  assign n42141 = n13475 & n42140 ;
  assign n42142 = ~n42139 & ~n42141 ;
  assign n42143 = \m0_data_i[8]_pad  & n13467 ;
  assign n42144 = n13475 & n42143 ;
  assign n42145 = \m7_data_i[8]_pad  & ~n13467 ;
  assign n42146 = n13492 & n42145 ;
  assign n42147 = ~n42144 & ~n42146 ;
  assign n42148 = n42142 & n42147 ;
  assign n42149 = n42137 & n42148 ;
  assign n42150 = \m3_data_i[9]_pad  & ~n13467 ;
  assign n42151 = n13484 & n42150 ;
  assign n42152 = \m4_data_i[9]_pad  & n13467 ;
  assign n42153 = n13460 & n42152 ;
  assign n42154 = ~n42151 & ~n42153 ;
  assign n42155 = \m6_data_i[9]_pad  & n13467 ;
  assign n42156 = n13492 & n42155 ;
  assign n42157 = \m2_data_i[9]_pad  & n13467 ;
  assign n42158 = n13484 & n42157 ;
  assign n42159 = ~n42156 & ~n42158 ;
  assign n42160 = n42154 & n42159 ;
  assign n42161 = \m5_data_i[9]_pad  & ~n13467 ;
  assign n42162 = n13460 & n42161 ;
  assign n42163 = \m1_data_i[9]_pad  & ~n13467 ;
  assign n42164 = n13475 & n42163 ;
  assign n42165 = ~n42162 & ~n42164 ;
  assign n42166 = \m0_data_i[9]_pad  & n13467 ;
  assign n42167 = n13475 & n42166 ;
  assign n42168 = \m7_data_i[9]_pad  & ~n13467 ;
  assign n42169 = n13492 & n42168 ;
  assign n42170 = ~n42167 & ~n42169 ;
  assign n42171 = n42165 & n42170 ;
  assign n42172 = n42160 & n42171 ;
  assign n42173 = \m3_sel_i[0]_pad  & ~n13467 ;
  assign n42174 = n13484 & n42173 ;
  assign n42175 = \m4_sel_i[0]_pad  & n13467 ;
  assign n42176 = n13460 & n42175 ;
  assign n42177 = ~n42174 & ~n42176 ;
  assign n42178 = \m6_sel_i[0]_pad  & n13467 ;
  assign n42179 = n13492 & n42178 ;
  assign n42180 = \m2_sel_i[0]_pad  & n13467 ;
  assign n42181 = n13484 & n42180 ;
  assign n42182 = ~n42179 & ~n42181 ;
  assign n42183 = n42177 & n42182 ;
  assign n42184 = \m5_sel_i[0]_pad  & ~n13467 ;
  assign n42185 = n13460 & n42184 ;
  assign n42186 = \m1_sel_i[0]_pad  & ~n13467 ;
  assign n42187 = n13475 & n42186 ;
  assign n42188 = ~n42185 & ~n42187 ;
  assign n42189 = \m0_sel_i[0]_pad  & n13467 ;
  assign n42190 = n13475 & n42189 ;
  assign n42191 = \m7_sel_i[0]_pad  & ~n13467 ;
  assign n42192 = n13492 & n42191 ;
  assign n42193 = ~n42190 & ~n42192 ;
  assign n42194 = n42188 & n42193 ;
  assign n42195 = n42183 & n42194 ;
  assign n42196 = \m3_sel_i[1]_pad  & ~n13467 ;
  assign n42197 = n13484 & n42196 ;
  assign n42198 = \m4_sel_i[1]_pad  & n13467 ;
  assign n42199 = n13460 & n42198 ;
  assign n42200 = ~n42197 & ~n42199 ;
  assign n42201 = \m6_sel_i[1]_pad  & n13467 ;
  assign n42202 = n13492 & n42201 ;
  assign n42203 = \m2_sel_i[1]_pad  & n13467 ;
  assign n42204 = n13484 & n42203 ;
  assign n42205 = ~n42202 & ~n42204 ;
  assign n42206 = n42200 & n42205 ;
  assign n42207 = \m5_sel_i[1]_pad  & ~n13467 ;
  assign n42208 = n13460 & n42207 ;
  assign n42209 = \m1_sel_i[1]_pad  & ~n13467 ;
  assign n42210 = n13475 & n42209 ;
  assign n42211 = ~n42208 & ~n42210 ;
  assign n42212 = \m0_sel_i[1]_pad  & n13467 ;
  assign n42213 = n13475 & n42212 ;
  assign n42214 = \m7_sel_i[1]_pad  & ~n13467 ;
  assign n42215 = n13492 & n42214 ;
  assign n42216 = ~n42213 & ~n42215 ;
  assign n42217 = n42211 & n42216 ;
  assign n42218 = n42206 & n42217 ;
  assign n42219 = \m3_sel_i[2]_pad  & ~n13467 ;
  assign n42220 = n13484 & n42219 ;
  assign n42221 = \m4_sel_i[2]_pad  & n13467 ;
  assign n42222 = n13460 & n42221 ;
  assign n42223 = ~n42220 & ~n42222 ;
  assign n42224 = \m6_sel_i[2]_pad  & n13467 ;
  assign n42225 = n13492 & n42224 ;
  assign n42226 = \m2_sel_i[2]_pad  & n13467 ;
  assign n42227 = n13484 & n42226 ;
  assign n42228 = ~n42225 & ~n42227 ;
  assign n42229 = n42223 & n42228 ;
  assign n42230 = \m5_sel_i[2]_pad  & ~n13467 ;
  assign n42231 = n13460 & n42230 ;
  assign n42232 = \m1_sel_i[2]_pad  & ~n13467 ;
  assign n42233 = n13475 & n42232 ;
  assign n42234 = ~n42231 & ~n42233 ;
  assign n42235 = \m0_sel_i[2]_pad  & n13467 ;
  assign n42236 = n13475 & n42235 ;
  assign n42237 = \m7_sel_i[2]_pad  & ~n13467 ;
  assign n42238 = n13492 & n42237 ;
  assign n42239 = ~n42236 & ~n42238 ;
  assign n42240 = n42234 & n42239 ;
  assign n42241 = n42229 & n42240 ;
  assign n42242 = \m3_sel_i[3]_pad  & ~n13467 ;
  assign n42243 = n13484 & n42242 ;
  assign n42244 = \m4_sel_i[3]_pad  & n13467 ;
  assign n42245 = n13460 & n42244 ;
  assign n42246 = ~n42243 & ~n42245 ;
  assign n42247 = \m6_sel_i[3]_pad  & n13467 ;
  assign n42248 = n13492 & n42247 ;
  assign n42249 = \m2_sel_i[3]_pad  & n13467 ;
  assign n42250 = n13484 & n42249 ;
  assign n42251 = ~n42248 & ~n42250 ;
  assign n42252 = n42246 & n42251 ;
  assign n42253 = \m5_sel_i[3]_pad  & ~n13467 ;
  assign n42254 = n13460 & n42253 ;
  assign n42255 = \m1_sel_i[3]_pad  & ~n13467 ;
  assign n42256 = n13475 & n42255 ;
  assign n42257 = ~n42254 & ~n42256 ;
  assign n42258 = \m0_sel_i[3]_pad  & n13467 ;
  assign n42259 = n13475 & n42258 ;
  assign n42260 = \m7_sel_i[3]_pad  & ~n13467 ;
  assign n42261 = n13492 & n42260 ;
  assign n42262 = ~n42259 & ~n42261 ;
  assign n42263 = n42257 & n42262 ;
  assign n42264 = n42252 & n42263 ;
  assign n42265 = \m3_stb_i_pad  & n14919 ;
  assign n42266 = ~n13467 & n42265 ;
  assign n42267 = n13484 & n42266 ;
  assign n42268 = \m2_stb_i_pad  & n14875 ;
  assign n42269 = n13467 & n42268 ;
  assign n42270 = n13484 & n42269 ;
  assign n42271 = ~n42267 & ~n42270 ;
  assign n42272 = \m4_stb_i_pad  & n14727 ;
  assign n42273 = n13467 & n42272 ;
  assign n42274 = n13460 & n42273 ;
  assign n42275 = \m1_stb_i_pad  & n14825 ;
  assign n42276 = ~n13467 & n42275 ;
  assign n42277 = n13475 & n42276 ;
  assign n42278 = ~n42274 & ~n42277 ;
  assign n42279 = n42271 & n42278 ;
  assign n42280 = \m5_stb_i_pad  & n14979 ;
  assign n42281 = ~n13467 & n42280 ;
  assign n42282 = n13460 & n42281 ;
  assign n42283 = \m7_stb_i_pad  & n15074 ;
  assign n42284 = ~n13467 & n42283 ;
  assign n42285 = n13492 & n42284 ;
  assign n42286 = ~n42282 & ~n42285 ;
  assign n42287 = \m6_stb_i_pad  & n15030 ;
  assign n42288 = n13467 & n42287 ;
  assign n42289 = n13492 & n42288 ;
  assign n42290 = \m0_stb_i_pad  & n15114 ;
  assign n42291 = n13467 & n42290 ;
  assign n42292 = n13475 & n42291 ;
  assign n42293 = ~n42289 & ~n42292 ;
  assign n42294 = n42286 & n42293 ;
  assign n42295 = n42279 & n42294 ;
  assign n42296 = \m3_we_i_pad  & ~n13467 ;
  assign n42297 = n13484 & n42296 ;
  assign n42298 = \m4_we_i_pad  & n13467 ;
  assign n42299 = n13460 & n42298 ;
  assign n42300 = ~n42297 & ~n42299 ;
  assign n42301 = \m6_we_i_pad  & n13467 ;
  assign n42302 = n13492 & n42301 ;
  assign n42303 = \m2_we_i_pad  & n13467 ;
  assign n42304 = n13484 & n42303 ;
  assign n42305 = ~n42302 & ~n42304 ;
  assign n42306 = n42300 & n42305 ;
  assign n42307 = \m5_we_i_pad  & ~n13467 ;
  assign n42308 = n13460 & n42307 ;
  assign n42309 = \m1_we_i_pad  & ~n13467 ;
  assign n42310 = n13475 & n42309 ;
  assign n42311 = ~n42308 & ~n42310 ;
  assign n42312 = \m0_we_i_pad  & n13467 ;
  assign n42313 = n13475 & n42312 ;
  assign n42314 = \m7_we_i_pad  & ~n13467 ;
  assign n42315 = n13492 & n42314 ;
  assign n42316 = ~n42313 & ~n42315 ;
  assign n42317 = n42311 & n42316 ;
  assign n42318 = n42306 & n42317 ;
  assign n42319 = \m3_addr_i[0]_pad  & ~n13547 ;
  assign n42320 = n13540 & n42319 ;
  assign n42321 = \m4_addr_i[0]_pad  & n13547 ;
  assign n42322 = n13555 & n42321 ;
  assign n42323 = ~n42320 & ~n42322 ;
  assign n42324 = \m6_addr_i[0]_pad  & n13547 ;
  assign n42325 = n13564 & n42324 ;
  assign n42326 = \m7_addr_i[0]_pad  & ~n13547 ;
  assign n42327 = n13564 & n42326 ;
  assign n42328 = ~n42325 & ~n42327 ;
  assign n42329 = n42323 & n42328 ;
  assign n42330 = \m5_addr_i[0]_pad  & ~n13547 ;
  assign n42331 = n13555 & n42330 ;
  assign n42332 = \m0_addr_i[0]_pad  & n13547 ;
  assign n42333 = n13572 & n42332 ;
  assign n42334 = ~n42331 & ~n42333 ;
  assign n42335 = \m1_addr_i[0]_pad  & ~n13547 ;
  assign n42336 = n13572 & n42335 ;
  assign n42337 = \m2_addr_i[0]_pad  & n13547 ;
  assign n42338 = n13540 & n42337 ;
  assign n42339 = ~n42336 & ~n42338 ;
  assign n42340 = n42334 & n42339 ;
  assign n42341 = n42329 & n42340 ;
  assign n42342 = \m3_addr_i[10]_pad  & ~n13547 ;
  assign n42343 = n13540 & n42342 ;
  assign n42344 = \m4_addr_i[10]_pad  & n13547 ;
  assign n42345 = n13555 & n42344 ;
  assign n42346 = ~n42343 & ~n42345 ;
  assign n42347 = \m6_addr_i[10]_pad  & n13547 ;
  assign n42348 = n13564 & n42347 ;
  assign n42349 = \m2_addr_i[10]_pad  & n13547 ;
  assign n42350 = n13540 & n42349 ;
  assign n42351 = ~n42348 & ~n42350 ;
  assign n42352 = n42346 & n42351 ;
  assign n42353 = \m5_addr_i[10]_pad  & ~n13547 ;
  assign n42354 = n13555 & n42353 ;
  assign n42355 = \m1_addr_i[10]_pad  & ~n13547 ;
  assign n42356 = n13572 & n42355 ;
  assign n42357 = ~n42354 & ~n42356 ;
  assign n42358 = \m0_addr_i[10]_pad  & n13547 ;
  assign n42359 = n13572 & n42358 ;
  assign n42360 = \m7_addr_i[10]_pad  & ~n13547 ;
  assign n42361 = n13564 & n42360 ;
  assign n42362 = ~n42359 & ~n42361 ;
  assign n42363 = n42357 & n42362 ;
  assign n42364 = n42352 & n42363 ;
  assign n42365 = \m3_addr_i[11]_pad  & ~n13547 ;
  assign n42366 = n13540 & n42365 ;
  assign n42367 = \m4_addr_i[11]_pad  & n13547 ;
  assign n42368 = n13555 & n42367 ;
  assign n42369 = ~n42366 & ~n42368 ;
  assign n42370 = \m6_addr_i[11]_pad  & n13547 ;
  assign n42371 = n13564 & n42370 ;
  assign n42372 = \m2_addr_i[11]_pad  & n13547 ;
  assign n42373 = n13540 & n42372 ;
  assign n42374 = ~n42371 & ~n42373 ;
  assign n42375 = n42369 & n42374 ;
  assign n42376 = \m5_addr_i[11]_pad  & ~n13547 ;
  assign n42377 = n13555 & n42376 ;
  assign n42378 = \m1_addr_i[11]_pad  & ~n13547 ;
  assign n42379 = n13572 & n42378 ;
  assign n42380 = ~n42377 & ~n42379 ;
  assign n42381 = \m0_addr_i[11]_pad  & n13547 ;
  assign n42382 = n13572 & n42381 ;
  assign n42383 = \m7_addr_i[11]_pad  & ~n13547 ;
  assign n42384 = n13564 & n42383 ;
  assign n42385 = ~n42382 & ~n42384 ;
  assign n42386 = n42380 & n42385 ;
  assign n42387 = n42375 & n42386 ;
  assign n42388 = \m6_addr_i[12]_pad  & n13547 ;
  assign n42389 = n13564 & n42388 ;
  assign n42390 = \m5_addr_i[12]_pad  & ~n13547 ;
  assign n42391 = n13555 & n42390 ;
  assign n42392 = ~n42389 & ~n42391 ;
  assign n42393 = \m1_addr_i[12]_pad  & ~n13547 ;
  assign n42394 = n13572 & n42393 ;
  assign n42395 = \m4_addr_i[12]_pad  & n13547 ;
  assign n42396 = n13555 & n42395 ;
  assign n42397 = ~n42394 & ~n42396 ;
  assign n42398 = n42392 & n42397 ;
  assign n42399 = \m2_addr_i[12]_pad  & n13547 ;
  assign n42400 = n13540 & n42399 ;
  assign n42401 = \m3_addr_i[12]_pad  & ~n13547 ;
  assign n42402 = n13540 & n42401 ;
  assign n42403 = ~n42400 & ~n42402 ;
  assign n42404 = \m0_addr_i[12]_pad  & n13547 ;
  assign n42405 = n13572 & n42404 ;
  assign n42406 = \m7_addr_i[12]_pad  & ~n13547 ;
  assign n42407 = n13564 & n42406 ;
  assign n42408 = ~n42405 & ~n42407 ;
  assign n42409 = n42403 & n42408 ;
  assign n42410 = n42398 & n42409 ;
  assign n42411 = \m6_addr_i[13]_pad  & n13547 ;
  assign n42412 = n13564 & n42411 ;
  assign n42413 = \m5_addr_i[13]_pad  & ~n13547 ;
  assign n42414 = n13555 & n42413 ;
  assign n42415 = ~n42412 & ~n42414 ;
  assign n42416 = \m0_addr_i[13]_pad  & n13547 ;
  assign n42417 = n13572 & n42416 ;
  assign n42418 = \m4_addr_i[13]_pad  & n13547 ;
  assign n42419 = n13555 & n42418 ;
  assign n42420 = ~n42417 & ~n42419 ;
  assign n42421 = n42415 & n42420 ;
  assign n42422 = \m7_addr_i[13]_pad  & ~n13547 ;
  assign n42423 = n13564 & n42422 ;
  assign n42424 = \m3_addr_i[13]_pad  & ~n13547 ;
  assign n42425 = n13540 & n42424 ;
  assign n42426 = ~n42423 & ~n42425 ;
  assign n42427 = \m1_addr_i[13]_pad  & ~n13547 ;
  assign n42428 = n13572 & n42427 ;
  assign n42429 = \m2_addr_i[13]_pad  & n13547 ;
  assign n42430 = n13540 & n42429 ;
  assign n42431 = ~n42428 & ~n42430 ;
  assign n42432 = n42426 & n42431 ;
  assign n42433 = n42421 & n42432 ;
  assign n42434 = \m3_addr_i[14]_pad  & ~n13547 ;
  assign n42435 = n13540 & n42434 ;
  assign n42436 = \m4_addr_i[14]_pad  & n13547 ;
  assign n42437 = n13555 & n42436 ;
  assign n42438 = ~n42435 & ~n42437 ;
  assign n42439 = \m6_addr_i[14]_pad  & n13547 ;
  assign n42440 = n13564 & n42439 ;
  assign n42441 = \m2_addr_i[14]_pad  & n13547 ;
  assign n42442 = n13540 & n42441 ;
  assign n42443 = ~n42440 & ~n42442 ;
  assign n42444 = n42438 & n42443 ;
  assign n42445 = \m5_addr_i[14]_pad  & ~n13547 ;
  assign n42446 = n13555 & n42445 ;
  assign n42447 = \m1_addr_i[14]_pad  & ~n13547 ;
  assign n42448 = n13572 & n42447 ;
  assign n42449 = ~n42446 & ~n42448 ;
  assign n42450 = \m0_addr_i[14]_pad  & n13547 ;
  assign n42451 = n13572 & n42450 ;
  assign n42452 = \m7_addr_i[14]_pad  & ~n13547 ;
  assign n42453 = n13564 & n42452 ;
  assign n42454 = ~n42451 & ~n42453 ;
  assign n42455 = n42449 & n42454 ;
  assign n42456 = n42444 & n42455 ;
  assign n42457 = \m6_addr_i[15]_pad  & n13547 ;
  assign n42458 = n13564 & n42457 ;
  assign n42459 = \m5_addr_i[15]_pad  & ~n13547 ;
  assign n42460 = n13555 & n42459 ;
  assign n42461 = ~n42458 & ~n42460 ;
  assign n42462 = \m3_addr_i[15]_pad  & ~n13547 ;
  assign n42463 = n13540 & n42462 ;
  assign n42464 = \m2_addr_i[15]_pad  & n13547 ;
  assign n42465 = n13540 & n42464 ;
  assign n42466 = ~n42463 & ~n42465 ;
  assign n42467 = n42461 & n42466 ;
  assign n42468 = \m4_addr_i[15]_pad  & n13547 ;
  assign n42469 = n13555 & n42468 ;
  assign n42470 = \m1_addr_i[15]_pad  & ~n13547 ;
  assign n42471 = n13572 & n42470 ;
  assign n42472 = ~n42469 & ~n42471 ;
  assign n42473 = \m0_addr_i[15]_pad  & n13547 ;
  assign n42474 = n13572 & n42473 ;
  assign n42475 = \m7_addr_i[15]_pad  & ~n13547 ;
  assign n42476 = n13564 & n42475 ;
  assign n42477 = ~n42474 & ~n42476 ;
  assign n42478 = n42472 & n42477 ;
  assign n42479 = n42467 & n42478 ;
  assign n42480 = \m3_addr_i[16]_pad  & ~n13547 ;
  assign n42481 = n13540 & n42480 ;
  assign n42482 = \m4_addr_i[16]_pad  & n13547 ;
  assign n42483 = n13555 & n42482 ;
  assign n42484 = ~n42481 & ~n42483 ;
  assign n42485 = \m6_addr_i[16]_pad  & n13547 ;
  assign n42486 = n13564 & n42485 ;
  assign n42487 = \m2_addr_i[16]_pad  & n13547 ;
  assign n42488 = n13540 & n42487 ;
  assign n42489 = ~n42486 & ~n42488 ;
  assign n42490 = n42484 & n42489 ;
  assign n42491 = \m5_addr_i[16]_pad  & ~n13547 ;
  assign n42492 = n13555 & n42491 ;
  assign n42493 = \m1_addr_i[16]_pad  & ~n13547 ;
  assign n42494 = n13572 & n42493 ;
  assign n42495 = ~n42492 & ~n42494 ;
  assign n42496 = \m0_addr_i[16]_pad  & n13547 ;
  assign n42497 = n13572 & n42496 ;
  assign n42498 = \m7_addr_i[16]_pad  & ~n13547 ;
  assign n42499 = n13564 & n42498 ;
  assign n42500 = ~n42497 & ~n42499 ;
  assign n42501 = n42495 & n42500 ;
  assign n42502 = n42490 & n42501 ;
  assign n42503 = \m6_addr_i[17]_pad  & n13547 ;
  assign n42504 = n13564 & n42503 ;
  assign n42505 = \m5_addr_i[17]_pad  & ~n13547 ;
  assign n42506 = n13555 & n42505 ;
  assign n42507 = ~n42504 & ~n42506 ;
  assign n42508 = \m1_addr_i[17]_pad  & ~n13547 ;
  assign n42509 = n13572 & n42508 ;
  assign n42510 = \m4_addr_i[17]_pad  & n13547 ;
  assign n42511 = n13555 & n42510 ;
  assign n42512 = ~n42509 & ~n42511 ;
  assign n42513 = n42507 & n42512 ;
  assign n42514 = \m2_addr_i[17]_pad  & n13547 ;
  assign n42515 = n13540 & n42514 ;
  assign n42516 = \m3_addr_i[17]_pad  & ~n13547 ;
  assign n42517 = n13540 & n42516 ;
  assign n42518 = ~n42515 & ~n42517 ;
  assign n42519 = \m0_addr_i[17]_pad  & n13547 ;
  assign n42520 = n13572 & n42519 ;
  assign n42521 = \m7_addr_i[17]_pad  & ~n13547 ;
  assign n42522 = n13564 & n42521 ;
  assign n42523 = ~n42520 & ~n42522 ;
  assign n42524 = n42518 & n42523 ;
  assign n42525 = n42513 & n42524 ;
  assign n42526 = \m3_addr_i[18]_pad  & ~n13547 ;
  assign n42527 = n13540 & n42526 ;
  assign n42528 = \m4_addr_i[18]_pad  & n13547 ;
  assign n42529 = n13555 & n42528 ;
  assign n42530 = ~n42527 & ~n42529 ;
  assign n42531 = \m6_addr_i[18]_pad  & n13547 ;
  assign n42532 = n13564 & n42531 ;
  assign n42533 = \m2_addr_i[18]_pad  & n13547 ;
  assign n42534 = n13540 & n42533 ;
  assign n42535 = ~n42532 & ~n42534 ;
  assign n42536 = n42530 & n42535 ;
  assign n42537 = \m5_addr_i[18]_pad  & ~n13547 ;
  assign n42538 = n13555 & n42537 ;
  assign n42539 = \m1_addr_i[18]_pad  & ~n13547 ;
  assign n42540 = n13572 & n42539 ;
  assign n42541 = ~n42538 & ~n42540 ;
  assign n42542 = \m0_addr_i[18]_pad  & n13547 ;
  assign n42543 = n13572 & n42542 ;
  assign n42544 = \m7_addr_i[18]_pad  & ~n13547 ;
  assign n42545 = n13564 & n42544 ;
  assign n42546 = ~n42543 & ~n42545 ;
  assign n42547 = n42541 & n42546 ;
  assign n42548 = n42536 & n42547 ;
  assign n42549 = \m3_addr_i[19]_pad  & ~n13547 ;
  assign n42550 = n13540 & n42549 ;
  assign n42551 = \m4_addr_i[19]_pad  & n13547 ;
  assign n42552 = n13555 & n42551 ;
  assign n42553 = ~n42550 & ~n42552 ;
  assign n42554 = \m6_addr_i[19]_pad  & n13547 ;
  assign n42555 = n13564 & n42554 ;
  assign n42556 = \m2_addr_i[19]_pad  & n13547 ;
  assign n42557 = n13540 & n42556 ;
  assign n42558 = ~n42555 & ~n42557 ;
  assign n42559 = n42553 & n42558 ;
  assign n42560 = \m5_addr_i[19]_pad  & ~n13547 ;
  assign n42561 = n13555 & n42560 ;
  assign n42562 = \m1_addr_i[19]_pad  & ~n13547 ;
  assign n42563 = n13572 & n42562 ;
  assign n42564 = ~n42561 & ~n42563 ;
  assign n42565 = \m0_addr_i[19]_pad  & n13547 ;
  assign n42566 = n13572 & n42565 ;
  assign n42567 = \m7_addr_i[19]_pad  & ~n13547 ;
  assign n42568 = n13564 & n42567 ;
  assign n42569 = ~n42566 & ~n42568 ;
  assign n42570 = n42564 & n42569 ;
  assign n42571 = n42559 & n42570 ;
  assign n42572 = \m3_addr_i[1]_pad  & ~n13547 ;
  assign n42573 = n13540 & n42572 ;
  assign n42574 = \m4_addr_i[1]_pad  & n13547 ;
  assign n42575 = n13555 & n42574 ;
  assign n42576 = ~n42573 & ~n42575 ;
  assign n42577 = \m6_addr_i[1]_pad  & n13547 ;
  assign n42578 = n13564 & n42577 ;
  assign n42579 = \m2_addr_i[1]_pad  & n13547 ;
  assign n42580 = n13540 & n42579 ;
  assign n42581 = ~n42578 & ~n42580 ;
  assign n42582 = n42576 & n42581 ;
  assign n42583 = \m5_addr_i[1]_pad  & ~n13547 ;
  assign n42584 = n13555 & n42583 ;
  assign n42585 = \m1_addr_i[1]_pad  & ~n13547 ;
  assign n42586 = n13572 & n42585 ;
  assign n42587 = ~n42584 & ~n42586 ;
  assign n42588 = \m0_addr_i[1]_pad  & n13547 ;
  assign n42589 = n13572 & n42588 ;
  assign n42590 = \m7_addr_i[1]_pad  & ~n13547 ;
  assign n42591 = n13564 & n42590 ;
  assign n42592 = ~n42589 & ~n42591 ;
  assign n42593 = n42587 & n42592 ;
  assign n42594 = n42582 & n42593 ;
  assign n42595 = \m3_addr_i[20]_pad  & ~n13547 ;
  assign n42596 = n13540 & n42595 ;
  assign n42597 = \m4_addr_i[20]_pad  & n13547 ;
  assign n42598 = n13555 & n42597 ;
  assign n42599 = ~n42596 & ~n42598 ;
  assign n42600 = \m6_addr_i[20]_pad  & n13547 ;
  assign n42601 = n13564 & n42600 ;
  assign n42602 = \m2_addr_i[20]_pad  & n13547 ;
  assign n42603 = n13540 & n42602 ;
  assign n42604 = ~n42601 & ~n42603 ;
  assign n42605 = n42599 & n42604 ;
  assign n42606 = \m5_addr_i[20]_pad  & ~n13547 ;
  assign n42607 = n13555 & n42606 ;
  assign n42608 = \m1_addr_i[20]_pad  & ~n13547 ;
  assign n42609 = n13572 & n42608 ;
  assign n42610 = ~n42607 & ~n42609 ;
  assign n42611 = \m0_addr_i[20]_pad  & n13547 ;
  assign n42612 = n13572 & n42611 ;
  assign n42613 = \m7_addr_i[20]_pad  & ~n13547 ;
  assign n42614 = n13564 & n42613 ;
  assign n42615 = ~n42612 & ~n42614 ;
  assign n42616 = n42610 & n42615 ;
  assign n42617 = n42605 & n42616 ;
  assign n42618 = \m3_addr_i[21]_pad  & ~n13547 ;
  assign n42619 = n13540 & n42618 ;
  assign n42620 = \m4_addr_i[21]_pad  & n13547 ;
  assign n42621 = n13555 & n42620 ;
  assign n42622 = ~n42619 & ~n42621 ;
  assign n42623 = \m6_addr_i[21]_pad  & n13547 ;
  assign n42624 = n13564 & n42623 ;
  assign n42625 = \m2_addr_i[21]_pad  & n13547 ;
  assign n42626 = n13540 & n42625 ;
  assign n42627 = ~n42624 & ~n42626 ;
  assign n42628 = n42622 & n42627 ;
  assign n42629 = \m5_addr_i[21]_pad  & ~n13547 ;
  assign n42630 = n13555 & n42629 ;
  assign n42631 = \m1_addr_i[21]_pad  & ~n13547 ;
  assign n42632 = n13572 & n42631 ;
  assign n42633 = ~n42630 & ~n42632 ;
  assign n42634 = \m0_addr_i[21]_pad  & n13547 ;
  assign n42635 = n13572 & n42634 ;
  assign n42636 = \m7_addr_i[21]_pad  & ~n13547 ;
  assign n42637 = n13564 & n42636 ;
  assign n42638 = ~n42635 & ~n42637 ;
  assign n42639 = n42633 & n42638 ;
  assign n42640 = n42628 & n42639 ;
  assign n42641 = \m0_addr_i[22]_pad  & n13547 ;
  assign n42642 = n13572 & n42641 ;
  assign n42643 = \m7_addr_i[22]_pad  & ~n13547 ;
  assign n42644 = n13564 & n42643 ;
  assign n42645 = ~n42642 & ~n42644 ;
  assign n42646 = \m6_addr_i[22]_pad  & n13547 ;
  assign n42647 = n13564 & n42646 ;
  assign n42648 = \m2_addr_i[22]_pad  & n13547 ;
  assign n42649 = n13540 & n42648 ;
  assign n42650 = ~n42647 & ~n42649 ;
  assign n42651 = n42645 & n42650 ;
  assign n42652 = \m5_addr_i[22]_pad  & ~n13547 ;
  assign n42653 = n13555 & n42652 ;
  assign n42654 = \m1_addr_i[22]_pad  & ~n13547 ;
  assign n42655 = n13572 & n42654 ;
  assign n42656 = ~n42653 & ~n42655 ;
  assign n42657 = \m3_addr_i[22]_pad  & ~n13547 ;
  assign n42658 = n13540 & n42657 ;
  assign n42659 = \m4_addr_i[22]_pad  & n13547 ;
  assign n42660 = n13555 & n42659 ;
  assign n42661 = ~n42658 & ~n42660 ;
  assign n42662 = n42656 & n42661 ;
  assign n42663 = n42651 & n42662 ;
  assign n42664 = \m3_addr_i[23]_pad  & ~n13547 ;
  assign n42665 = n13540 & n42664 ;
  assign n42666 = \m4_addr_i[23]_pad  & n13547 ;
  assign n42667 = n13555 & n42666 ;
  assign n42668 = ~n42665 & ~n42667 ;
  assign n42669 = \m6_addr_i[23]_pad  & n13547 ;
  assign n42670 = n13564 & n42669 ;
  assign n42671 = \m2_addr_i[23]_pad  & n13547 ;
  assign n42672 = n13540 & n42671 ;
  assign n42673 = ~n42670 & ~n42672 ;
  assign n42674 = n42668 & n42673 ;
  assign n42675 = \m5_addr_i[23]_pad  & ~n13547 ;
  assign n42676 = n13555 & n42675 ;
  assign n42677 = \m1_addr_i[23]_pad  & ~n13547 ;
  assign n42678 = n13572 & n42677 ;
  assign n42679 = ~n42676 & ~n42678 ;
  assign n42680 = \m0_addr_i[23]_pad  & n13547 ;
  assign n42681 = n13572 & n42680 ;
  assign n42682 = \m7_addr_i[23]_pad  & ~n13547 ;
  assign n42683 = n13564 & n42682 ;
  assign n42684 = ~n42681 & ~n42683 ;
  assign n42685 = n42679 & n42684 ;
  assign n42686 = n42674 & n42685 ;
  assign n42687 = \m3_addr_i[24]_pad  & ~n13547 ;
  assign n42688 = n13540 & n42687 ;
  assign n42689 = \m4_addr_i[24]_pad  & n13547 ;
  assign n42690 = n13555 & n42689 ;
  assign n42691 = ~n42688 & ~n42690 ;
  assign n42692 = \m5_addr_i[24]_pad  & ~n13547 ;
  assign n42693 = n13555 & n42692 ;
  assign n42694 = \m2_addr_i[24]_pad  & n13547 ;
  assign n42695 = n13540 & n42694 ;
  assign n42696 = ~n42693 & ~n42695 ;
  assign n42697 = n42691 & n42696 ;
  assign n42698 = \m6_addr_i[24]_pad  & n13547 ;
  assign n42699 = n13564 & n42698 ;
  assign n42700 = \m1_addr_i[24]_pad  & ~n13547 ;
  assign n42701 = n13572 & n42700 ;
  assign n42702 = ~n42699 & ~n42701 ;
  assign n42703 = \m0_addr_i[24]_pad  & n13547 ;
  assign n42704 = n13572 & n42703 ;
  assign n42705 = \m7_addr_i[24]_pad  & ~n13547 ;
  assign n42706 = n13564 & n42705 ;
  assign n42707 = ~n42704 & ~n42706 ;
  assign n42708 = n42702 & n42707 ;
  assign n42709 = n42697 & n42708 ;
  assign n42710 = \m5_addr_i[25]_pad  & ~n13547 ;
  assign n42711 = n13555 & n42710 ;
  assign n42712 = \m6_addr_i[25]_pad  & n13547 ;
  assign n42713 = n13564 & n42712 ;
  assign n42714 = ~n42711 & ~n42713 ;
  assign n42715 = \m0_addr_i[25]_pad  & n13547 ;
  assign n42716 = n13572 & n42715 ;
  assign n42717 = \m4_addr_i[25]_pad  & n13547 ;
  assign n42718 = n13555 & n42717 ;
  assign n42719 = ~n42716 & ~n42718 ;
  assign n42720 = n42714 & n42719 ;
  assign n42721 = \m7_addr_i[25]_pad  & ~n13547 ;
  assign n42722 = n13564 & n42721 ;
  assign n42723 = \m3_addr_i[25]_pad  & ~n13547 ;
  assign n42724 = n13540 & n42723 ;
  assign n42725 = ~n42722 & ~n42724 ;
  assign n42726 = \m1_addr_i[25]_pad  & ~n13547 ;
  assign n42727 = n13572 & n42726 ;
  assign n42728 = \m2_addr_i[25]_pad  & n13547 ;
  assign n42729 = n13540 & n42728 ;
  assign n42730 = ~n42727 & ~n42729 ;
  assign n42731 = n42725 & n42730 ;
  assign n42732 = n42720 & n42731 ;
  assign n42733 = \m5_addr_i[26]_pad  & ~n13547 ;
  assign n42734 = n13555 & n42733 ;
  assign n42735 = \m6_addr_i[26]_pad  & n13547 ;
  assign n42736 = n13564 & n42735 ;
  assign n42737 = ~n42734 & ~n42736 ;
  assign n42738 = \m1_addr_i[26]_pad  & ~n13547 ;
  assign n42739 = n13572 & n42738 ;
  assign n42740 = \m4_addr_i[26]_pad  & n13547 ;
  assign n42741 = n13555 & n42740 ;
  assign n42742 = ~n42739 & ~n42741 ;
  assign n42743 = n42737 & n42742 ;
  assign n42744 = \m2_addr_i[26]_pad  & n13547 ;
  assign n42745 = n13540 & n42744 ;
  assign n42746 = \m3_addr_i[26]_pad  & ~n13547 ;
  assign n42747 = n13540 & n42746 ;
  assign n42748 = ~n42745 & ~n42747 ;
  assign n42749 = \m0_addr_i[26]_pad  & n13547 ;
  assign n42750 = n13572 & n42749 ;
  assign n42751 = \m7_addr_i[26]_pad  & ~n13547 ;
  assign n42752 = n13564 & n42751 ;
  assign n42753 = ~n42750 & ~n42752 ;
  assign n42754 = n42748 & n42753 ;
  assign n42755 = n42743 & n42754 ;
  assign n42756 = \m3_addr_i[27]_pad  & ~n13547 ;
  assign n42757 = n13540 & n42756 ;
  assign n42758 = \m4_addr_i[27]_pad  & n13547 ;
  assign n42759 = n13555 & n42758 ;
  assign n42760 = ~n42757 & ~n42759 ;
  assign n42761 = \m0_addr_i[27]_pad  & n13547 ;
  assign n42762 = n13572 & n42761 ;
  assign n42763 = \m6_addr_i[27]_pad  & n13547 ;
  assign n42764 = n13564 & n42763 ;
  assign n42765 = ~n42762 & ~n42764 ;
  assign n42766 = n42760 & n42765 ;
  assign n42767 = \m7_addr_i[27]_pad  & ~n13547 ;
  assign n42768 = n13564 & n42767 ;
  assign n42769 = \m5_addr_i[27]_pad  & ~n13547 ;
  assign n42770 = n13555 & n42769 ;
  assign n42771 = ~n42768 & ~n42770 ;
  assign n42772 = \m1_addr_i[27]_pad  & ~n13547 ;
  assign n42773 = n13572 & n42772 ;
  assign n42774 = \m2_addr_i[27]_pad  & n13547 ;
  assign n42775 = n13540 & n42774 ;
  assign n42776 = ~n42773 & ~n42775 ;
  assign n42777 = n42771 & n42776 ;
  assign n42778 = n42766 & n42777 ;
  assign n42779 = \m3_addr_i[28]_pad  & ~n13547 ;
  assign n42780 = n13540 & n42779 ;
  assign n42781 = \m4_addr_i[28]_pad  & n13547 ;
  assign n42782 = n13555 & n42781 ;
  assign n42783 = ~n42780 & ~n42782 ;
  assign n42784 = \m1_addr_i[28]_pad  & ~n13547 ;
  assign n42785 = n13572 & n42784 ;
  assign n42786 = \m7_addr_i[28]_pad  & ~n13547 ;
  assign n42787 = n13564 & n42786 ;
  assign n42788 = ~n42785 & ~n42787 ;
  assign n42789 = n42783 & n42788 ;
  assign n42790 = \m2_addr_i[28]_pad  & n13547 ;
  assign n42791 = n13540 & n42790 ;
  assign n42792 = \m0_addr_i[28]_pad  & n13547 ;
  assign n42793 = n13572 & n42792 ;
  assign n42794 = ~n42791 & ~n42793 ;
  assign n42795 = \m5_addr_i[28]_pad  & ~n13547 ;
  assign n42796 = n13555 & n42795 ;
  assign n42797 = \m6_addr_i[28]_pad  & n13547 ;
  assign n42798 = n13564 & n42797 ;
  assign n42799 = ~n42796 & ~n42798 ;
  assign n42800 = n42794 & n42799 ;
  assign n42801 = n42789 & n42800 ;
  assign n42802 = \m5_addr_i[29]_pad  & ~n13547 ;
  assign n42803 = n13555 & n42802 ;
  assign n42804 = \m6_addr_i[29]_pad  & n13547 ;
  assign n42805 = n13564 & n42804 ;
  assign n42806 = ~n42803 & ~n42805 ;
  assign n42807 = \m0_addr_i[29]_pad  & n13547 ;
  assign n42808 = n13572 & n42807 ;
  assign n42809 = \m4_addr_i[29]_pad  & n13547 ;
  assign n42810 = n13555 & n42809 ;
  assign n42811 = ~n42808 & ~n42810 ;
  assign n42812 = n42806 & n42811 ;
  assign n42813 = \m7_addr_i[29]_pad  & ~n13547 ;
  assign n42814 = n13564 & n42813 ;
  assign n42815 = \m3_addr_i[29]_pad  & ~n13547 ;
  assign n42816 = n13540 & n42815 ;
  assign n42817 = ~n42814 & ~n42816 ;
  assign n42818 = \m1_addr_i[29]_pad  & ~n13547 ;
  assign n42819 = n13572 & n42818 ;
  assign n42820 = \m2_addr_i[29]_pad  & n13547 ;
  assign n42821 = n13540 & n42820 ;
  assign n42822 = ~n42819 & ~n42821 ;
  assign n42823 = n42817 & n42822 ;
  assign n42824 = n42812 & n42823 ;
  assign n42825 = \m0_addr_i[2]_pad  & n13547 ;
  assign n42826 = n13572 & n42825 ;
  assign n42827 = \m7_addr_i[2]_pad  & ~n13547 ;
  assign n42828 = n13564 & n42827 ;
  assign n42829 = ~n42826 & ~n42828 ;
  assign n42830 = \m1_addr_i[2]_pad  & ~n13547 ;
  assign n42831 = n13572 & n42830 ;
  assign n42832 = \m5_addr_i[2]_pad  & ~n13547 ;
  assign n42833 = n13555 & n42832 ;
  assign n42834 = ~n42831 & ~n42833 ;
  assign n42835 = n42829 & n42834 ;
  assign n42836 = \m2_addr_i[2]_pad  & n13547 ;
  assign n42837 = n13540 & n42836 ;
  assign n42838 = \m6_addr_i[2]_pad  & n13547 ;
  assign n42839 = n13564 & n42838 ;
  assign n42840 = ~n42837 & ~n42839 ;
  assign n42841 = \m3_addr_i[2]_pad  & ~n13547 ;
  assign n42842 = n13540 & n42841 ;
  assign n42843 = \m4_addr_i[2]_pad  & n13547 ;
  assign n42844 = n13555 & n42843 ;
  assign n42845 = ~n42842 & ~n42844 ;
  assign n42846 = n42840 & n42845 ;
  assign n42847 = n42835 & n42846 ;
  assign n42848 = \m5_addr_i[30]_pad  & ~n13547 ;
  assign n42849 = n13555 & n42848 ;
  assign n42850 = \m6_addr_i[30]_pad  & n13547 ;
  assign n42851 = n13564 & n42850 ;
  assign n42852 = ~n42849 & ~n42851 ;
  assign n42853 = \m0_addr_i[30]_pad  & n13547 ;
  assign n42854 = n13572 & n42853 ;
  assign n42855 = \m4_addr_i[30]_pad  & n13547 ;
  assign n42856 = n13555 & n42855 ;
  assign n42857 = ~n42854 & ~n42856 ;
  assign n42858 = n42852 & n42857 ;
  assign n42859 = \m7_addr_i[30]_pad  & ~n13547 ;
  assign n42860 = n13564 & n42859 ;
  assign n42861 = \m3_addr_i[30]_pad  & ~n13547 ;
  assign n42862 = n13540 & n42861 ;
  assign n42863 = ~n42860 & ~n42862 ;
  assign n42864 = \m1_addr_i[30]_pad  & ~n13547 ;
  assign n42865 = n13572 & n42864 ;
  assign n42866 = \m2_addr_i[30]_pad  & n13547 ;
  assign n42867 = n13540 & n42866 ;
  assign n42868 = ~n42865 & ~n42867 ;
  assign n42869 = n42863 & n42868 ;
  assign n42870 = n42858 & n42869 ;
  assign n42871 = \m5_addr_i[31]_pad  & ~n13547 ;
  assign n42872 = n13555 & n42871 ;
  assign n42873 = \m6_addr_i[31]_pad  & n13547 ;
  assign n42874 = n13564 & n42873 ;
  assign n42875 = ~n42872 & ~n42874 ;
  assign n42876 = \m3_addr_i[31]_pad  & ~n13547 ;
  assign n42877 = n13540 & n42876 ;
  assign n42878 = \m2_addr_i[31]_pad  & n13547 ;
  assign n42879 = n13540 & n42878 ;
  assign n42880 = ~n42877 & ~n42879 ;
  assign n42881 = n42875 & n42880 ;
  assign n42882 = \m4_addr_i[31]_pad  & n13547 ;
  assign n42883 = n13555 & n42882 ;
  assign n42884 = \m1_addr_i[31]_pad  & ~n13547 ;
  assign n42885 = n13572 & n42884 ;
  assign n42886 = ~n42883 & ~n42885 ;
  assign n42887 = \m0_addr_i[31]_pad  & n13547 ;
  assign n42888 = n13572 & n42887 ;
  assign n42889 = \m7_addr_i[31]_pad  & ~n13547 ;
  assign n42890 = n13564 & n42889 ;
  assign n42891 = ~n42888 & ~n42890 ;
  assign n42892 = n42886 & n42891 ;
  assign n42893 = n42881 & n42892 ;
  assign n42894 = \m1_addr_i[3]_pad  & ~n13547 ;
  assign n42895 = n13572 & n42894 ;
  assign n42896 = \m2_addr_i[3]_pad  & n13547 ;
  assign n42897 = n13540 & n42896 ;
  assign n42898 = ~n42895 & ~n42897 ;
  assign n42899 = \m0_addr_i[3]_pad  & n13547 ;
  assign n42900 = n13572 & n42899 ;
  assign n42901 = \m4_addr_i[3]_pad  & n13547 ;
  assign n42902 = n13555 & n42901 ;
  assign n42903 = ~n42900 & ~n42902 ;
  assign n42904 = n42898 & n42903 ;
  assign n42905 = \m7_addr_i[3]_pad  & ~n13547 ;
  assign n42906 = n13564 & n42905 ;
  assign n42907 = \m3_addr_i[3]_pad  & ~n13547 ;
  assign n42908 = n13540 & n42907 ;
  assign n42909 = ~n42906 & ~n42908 ;
  assign n42910 = \m6_addr_i[3]_pad  & n13547 ;
  assign n42911 = n13564 & n42910 ;
  assign n42912 = \m5_addr_i[3]_pad  & ~n13547 ;
  assign n42913 = n13555 & n42912 ;
  assign n42914 = ~n42911 & ~n42913 ;
  assign n42915 = n42909 & n42914 ;
  assign n42916 = n42904 & n42915 ;
  assign n42917 = \m6_addr_i[4]_pad  & n13547 ;
  assign n42918 = n13564 & n42917 ;
  assign n42919 = \m5_addr_i[4]_pad  & ~n13547 ;
  assign n42920 = n13555 & n42919 ;
  assign n42921 = ~n42918 & ~n42920 ;
  assign n42922 = \m0_addr_i[4]_pad  & n13547 ;
  assign n42923 = n13572 & n42922 ;
  assign n42924 = \m4_addr_i[4]_pad  & n13547 ;
  assign n42925 = n13555 & n42924 ;
  assign n42926 = ~n42923 & ~n42925 ;
  assign n42927 = n42921 & n42926 ;
  assign n42928 = \m7_addr_i[4]_pad  & ~n13547 ;
  assign n42929 = n13564 & n42928 ;
  assign n42930 = \m3_addr_i[4]_pad  & ~n13547 ;
  assign n42931 = n13540 & n42930 ;
  assign n42932 = ~n42929 & ~n42931 ;
  assign n42933 = \m1_addr_i[4]_pad  & ~n13547 ;
  assign n42934 = n13572 & n42933 ;
  assign n42935 = \m2_addr_i[4]_pad  & n13547 ;
  assign n42936 = n13540 & n42935 ;
  assign n42937 = ~n42934 & ~n42936 ;
  assign n42938 = n42932 & n42937 ;
  assign n42939 = n42927 & n42938 ;
  assign n42940 = \m6_addr_i[5]_pad  & n13547 ;
  assign n42941 = n13564 & n42940 ;
  assign n42942 = \m5_addr_i[5]_pad  & ~n13547 ;
  assign n42943 = n13555 & n42942 ;
  assign n42944 = ~n42941 & ~n42943 ;
  assign n42945 = \m1_addr_i[5]_pad  & ~n13547 ;
  assign n42946 = n13572 & n42945 ;
  assign n42947 = \m4_addr_i[5]_pad  & n13547 ;
  assign n42948 = n13555 & n42947 ;
  assign n42949 = ~n42946 & ~n42948 ;
  assign n42950 = n42944 & n42949 ;
  assign n42951 = \m2_addr_i[5]_pad  & n13547 ;
  assign n42952 = n13540 & n42951 ;
  assign n42953 = \m3_addr_i[5]_pad  & ~n13547 ;
  assign n42954 = n13540 & n42953 ;
  assign n42955 = ~n42952 & ~n42954 ;
  assign n42956 = \m0_addr_i[5]_pad  & n13547 ;
  assign n42957 = n13572 & n42956 ;
  assign n42958 = \m7_addr_i[5]_pad  & ~n13547 ;
  assign n42959 = n13564 & n42958 ;
  assign n42960 = ~n42957 & ~n42959 ;
  assign n42961 = n42955 & n42960 ;
  assign n42962 = n42950 & n42961 ;
  assign n42963 = \m6_addr_i[6]_pad  & n13547 ;
  assign n42964 = n13564 & n42963 ;
  assign n42965 = \m5_addr_i[6]_pad  & ~n13547 ;
  assign n42966 = n13555 & n42965 ;
  assign n42967 = ~n42964 & ~n42966 ;
  assign n42968 = \m0_addr_i[6]_pad  & n13547 ;
  assign n42969 = n13572 & n42968 ;
  assign n42970 = \m4_addr_i[6]_pad  & n13547 ;
  assign n42971 = n13555 & n42970 ;
  assign n42972 = ~n42969 & ~n42971 ;
  assign n42973 = n42967 & n42972 ;
  assign n42974 = \m7_addr_i[6]_pad  & ~n13547 ;
  assign n42975 = n13564 & n42974 ;
  assign n42976 = \m3_addr_i[6]_pad  & ~n13547 ;
  assign n42977 = n13540 & n42976 ;
  assign n42978 = ~n42975 & ~n42977 ;
  assign n42979 = \m1_addr_i[6]_pad  & ~n13547 ;
  assign n42980 = n13572 & n42979 ;
  assign n42981 = \m2_addr_i[6]_pad  & n13547 ;
  assign n42982 = n13540 & n42981 ;
  assign n42983 = ~n42980 & ~n42982 ;
  assign n42984 = n42978 & n42983 ;
  assign n42985 = n42973 & n42984 ;
  assign n42986 = \m3_addr_i[7]_pad  & ~n13547 ;
  assign n42987 = n13540 & n42986 ;
  assign n42988 = \m4_addr_i[7]_pad  & n13547 ;
  assign n42989 = n13555 & n42988 ;
  assign n42990 = ~n42987 & ~n42989 ;
  assign n42991 = \m1_addr_i[7]_pad  & ~n13547 ;
  assign n42992 = n13572 & n42991 ;
  assign n42993 = \m5_addr_i[7]_pad  & ~n13547 ;
  assign n42994 = n13555 & n42993 ;
  assign n42995 = ~n42992 & ~n42994 ;
  assign n42996 = n42990 & n42995 ;
  assign n42997 = \m2_addr_i[7]_pad  & n13547 ;
  assign n42998 = n13540 & n42997 ;
  assign n42999 = \m6_addr_i[7]_pad  & n13547 ;
  assign n43000 = n13564 & n42999 ;
  assign n43001 = ~n42998 & ~n43000 ;
  assign n43002 = \m0_addr_i[7]_pad  & n13547 ;
  assign n43003 = n13572 & n43002 ;
  assign n43004 = \m7_addr_i[7]_pad  & ~n13547 ;
  assign n43005 = n13564 & n43004 ;
  assign n43006 = ~n43003 & ~n43005 ;
  assign n43007 = n43001 & n43006 ;
  assign n43008 = n42996 & n43007 ;
  assign n43009 = \m0_addr_i[8]_pad  & n13547 ;
  assign n43010 = n13572 & n43009 ;
  assign n43011 = \m7_addr_i[8]_pad  & ~n13547 ;
  assign n43012 = n13564 & n43011 ;
  assign n43013 = ~n43010 & ~n43012 ;
  assign n43014 = \m3_addr_i[8]_pad  & ~n13547 ;
  assign n43015 = n13540 & n43014 ;
  assign n43016 = \m5_addr_i[8]_pad  & ~n13547 ;
  assign n43017 = n13555 & n43016 ;
  assign n43018 = ~n43015 & ~n43017 ;
  assign n43019 = n43013 & n43018 ;
  assign n43020 = \m4_addr_i[8]_pad  & n13547 ;
  assign n43021 = n13555 & n43020 ;
  assign n43022 = \m6_addr_i[8]_pad  & n13547 ;
  assign n43023 = n13564 & n43022 ;
  assign n43024 = ~n43021 & ~n43023 ;
  assign n43025 = \m1_addr_i[8]_pad  & ~n13547 ;
  assign n43026 = n13572 & n43025 ;
  assign n43027 = \m2_addr_i[8]_pad  & n13547 ;
  assign n43028 = n13540 & n43027 ;
  assign n43029 = ~n43026 & ~n43028 ;
  assign n43030 = n43024 & n43029 ;
  assign n43031 = n43019 & n43030 ;
  assign n43032 = \m6_addr_i[9]_pad  & n13547 ;
  assign n43033 = n13564 & n43032 ;
  assign n43034 = \m5_addr_i[9]_pad  & ~n13547 ;
  assign n43035 = n13555 & n43034 ;
  assign n43036 = ~n43033 & ~n43035 ;
  assign n43037 = \m0_addr_i[9]_pad  & n13547 ;
  assign n43038 = n13572 & n43037 ;
  assign n43039 = \m4_addr_i[9]_pad  & n13547 ;
  assign n43040 = n13555 & n43039 ;
  assign n43041 = ~n43038 & ~n43040 ;
  assign n43042 = n43036 & n43041 ;
  assign n43043 = \m7_addr_i[9]_pad  & ~n13547 ;
  assign n43044 = n13564 & n43043 ;
  assign n43045 = \m3_addr_i[9]_pad  & ~n13547 ;
  assign n43046 = n13540 & n43045 ;
  assign n43047 = ~n43044 & ~n43046 ;
  assign n43048 = \m1_addr_i[9]_pad  & ~n13547 ;
  assign n43049 = n13572 & n43048 ;
  assign n43050 = \m2_addr_i[9]_pad  & n13547 ;
  assign n43051 = n13540 & n43050 ;
  assign n43052 = ~n43049 & ~n43051 ;
  assign n43053 = n43047 & n43052 ;
  assign n43054 = n43042 & n43053 ;
  assign n43055 = \m3_data_i[0]_pad  & ~n13547 ;
  assign n43056 = n13540 & n43055 ;
  assign n43057 = \m4_data_i[0]_pad  & n13547 ;
  assign n43058 = n13555 & n43057 ;
  assign n43059 = ~n43056 & ~n43058 ;
  assign n43060 = \m0_data_i[0]_pad  & n13547 ;
  assign n43061 = n13572 & n43060 ;
  assign n43062 = \m5_data_i[0]_pad  & ~n13547 ;
  assign n43063 = n13555 & n43062 ;
  assign n43064 = ~n43061 & ~n43063 ;
  assign n43065 = n43059 & n43064 ;
  assign n43066 = \m7_data_i[0]_pad  & ~n13547 ;
  assign n43067 = n13564 & n43066 ;
  assign n43068 = \m6_data_i[0]_pad  & n13547 ;
  assign n43069 = n13564 & n43068 ;
  assign n43070 = ~n43067 & ~n43069 ;
  assign n43071 = \m1_data_i[0]_pad  & ~n13547 ;
  assign n43072 = n13572 & n43071 ;
  assign n43073 = \m2_data_i[0]_pad  & n13547 ;
  assign n43074 = n13540 & n43073 ;
  assign n43075 = ~n43072 & ~n43074 ;
  assign n43076 = n43070 & n43075 ;
  assign n43077 = n43065 & n43076 ;
  assign n43078 = \m3_data_i[10]_pad  & ~n13547 ;
  assign n43079 = n13540 & n43078 ;
  assign n43080 = \m4_data_i[10]_pad  & n13547 ;
  assign n43081 = n13555 & n43080 ;
  assign n43082 = ~n43079 & ~n43081 ;
  assign n43083 = \m6_data_i[10]_pad  & n13547 ;
  assign n43084 = n13564 & n43083 ;
  assign n43085 = \m2_data_i[10]_pad  & n13547 ;
  assign n43086 = n13540 & n43085 ;
  assign n43087 = ~n43084 & ~n43086 ;
  assign n43088 = n43082 & n43087 ;
  assign n43089 = \m5_data_i[10]_pad  & ~n13547 ;
  assign n43090 = n13555 & n43089 ;
  assign n43091 = \m1_data_i[10]_pad  & ~n13547 ;
  assign n43092 = n13572 & n43091 ;
  assign n43093 = ~n43090 & ~n43092 ;
  assign n43094 = \m0_data_i[10]_pad  & n13547 ;
  assign n43095 = n13572 & n43094 ;
  assign n43096 = \m7_data_i[10]_pad  & ~n13547 ;
  assign n43097 = n13564 & n43096 ;
  assign n43098 = ~n43095 & ~n43097 ;
  assign n43099 = n43093 & n43098 ;
  assign n43100 = n43088 & n43099 ;
  assign n43101 = \m3_data_i[11]_pad  & ~n13547 ;
  assign n43102 = n13540 & n43101 ;
  assign n43103 = \m4_data_i[11]_pad  & n13547 ;
  assign n43104 = n13555 & n43103 ;
  assign n43105 = ~n43102 & ~n43104 ;
  assign n43106 = \m6_data_i[11]_pad  & n13547 ;
  assign n43107 = n13564 & n43106 ;
  assign n43108 = \m2_data_i[11]_pad  & n13547 ;
  assign n43109 = n13540 & n43108 ;
  assign n43110 = ~n43107 & ~n43109 ;
  assign n43111 = n43105 & n43110 ;
  assign n43112 = \m5_data_i[11]_pad  & ~n13547 ;
  assign n43113 = n13555 & n43112 ;
  assign n43114 = \m1_data_i[11]_pad  & ~n13547 ;
  assign n43115 = n13572 & n43114 ;
  assign n43116 = ~n43113 & ~n43115 ;
  assign n43117 = \m0_data_i[11]_pad  & n13547 ;
  assign n43118 = n13572 & n43117 ;
  assign n43119 = \m7_data_i[11]_pad  & ~n13547 ;
  assign n43120 = n13564 & n43119 ;
  assign n43121 = ~n43118 & ~n43120 ;
  assign n43122 = n43116 & n43121 ;
  assign n43123 = n43111 & n43122 ;
  assign n43124 = \m3_data_i[12]_pad  & ~n13547 ;
  assign n43125 = n13540 & n43124 ;
  assign n43126 = \m4_data_i[12]_pad  & n13547 ;
  assign n43127 = n13555 & n43126 ;
  assign n43128 = ~n43125 & ~n43127 ;
  assign n43129 = \m6_data_i[12]_pad  & n13547 ;
  assign n43130 = n13564 & n43129 ;
  assign n43131 = \m2_data_i[12]_pad  & n13547 ;
  assign n43132 = n13540 & n43131 ;
  assign n43133 = ~n43130 & ~n43132 ;
  assign n43134 = n43128 & n43133 ;
  assign n43135 = \m5_data_i[12]_pad  & ~n13547 ;
  assign n43136 = n13555 & n43135 ;
  assign n43137 = \m1_data_i[12]_pad  & ~n13547 ;
  assign n43138 = n13572 & n43137 ;
  assign n43139 = ~n43136 & ~n43138 ;
  assign n43140 = \m0_data_i[12]_pad  & n13547 ;
  assign n43141 = n13572 & n43140 ;
  assign n43142 = \m7_data_i[12]_pad  & ~n13547 ;
  assign n43143 = n13564 & n43142 ;
  assign n43144 = ~n43141 & ~n43143 ;
  assign n43145 = n43139 & n43144 ;
  assign n43146 = n43134 & n43145 ;
  assign n43147 = \m3_data_i[13]_pad  & ~n13547 ;
  assign n43148 = n13540 & n43147 ;
  assign n43149 = \m4_data_i[13]_pad  & n13547 ;
  assign n43150 = n13555 & n43149 ;
  assign n43151 = ~n43148 & ~n43150 ;
  assign n43152 = \m6_data_i[13]_pad  & n13547 ;
  assign n43153 = n13564 & n43152 ;
  assign n43154 = \m2_data_i[13]_pad  & n13547 ;
  assign n43155 = n13540 & n43154 ;
  assign n43156 = ~n43153 & ~n43155 ;
  assign n43157 = n43151 & n43156 ;
  assign n43158 = \m5_data_i[13]_pad  & ~n13547 ;
  assign n43159 = n13555 & n43158 ;
  assign n43160 = \m1_data_i[13]_pad  & ~n13547 ;
  assign n43161 = n13572 & n43160 ;
  assign n43162 = ~n43159 & ~n43161 ;
  assign n43163 = \m0_data_i[13]_pad  & n13547 ;
  assign n43164 = n13572 & n43163 ;
  assign n43165 = \m7_data_i[13]_pad  & ~n13547 ;
  assign n43166 = n13564 & n43165 ;
  assign n43167 = ~n43164 & ~n43166 ;
  assign n43168 = n43162 & n43167 ;
  assign n43169 = n43157 & n43168 ;
  assign n43170 = \m3_data_i[14]_pad  & ~n13547 ;
  assign n43171 = n13540 & n43170 ;
  assign n43172 = \m4_data_i[14]_pad  & n13547 ;
  assign n43173 = n13555 & n43172 ;
  assign n43174 = ~n43171 & ~n43173 ;
  assign n43175 = \m6_data_i[14]_pad  & n13547 ;
  assign n43176 = n13564 & n43175 ;
  assign n43177 = \m2_data_i[14]_pad  & n13547 ;
  assign n43178 = n13540 & n43177 ;
  assign n43179 = ~n43176 & ~n43178 ;
  assign n43180 = n43174 & n43179 ;
  assign n43181 = \m5_data_i[14]_pad  & ~n13547 ;
  assign n43182 = n13555 & n43181 ;
  assign n43183 = \m1_data_i[14]_pad  & ~n13547 ;
  assign n43184 = n13572 & n43183 ;
  assign n43185 = ~n43182 & ~n43184 ;
  assign n43186 = \m0_data_i[14]_pad  & n13547 ;
  assign n43187 = n13572 & n43186 ;
  assign n43188 = \m7_data_i[14]_pad  & ~n13547 ;
  assign n43189 = n13564 & n43188 ;
  assign n43190 = ~n43187 & ~n43189 ;
  assign n43191 = n43185 & n43190 ;
  assign n43192 = n43180 & n43191 ;
  assign n43193 = \m3_data_i[15]_pad  & ~n13547 ;
  assign n43194 = n13540 & n43193 ;
  assign n43195 = \m4_data_i[15]_pad  & n13547 ;
  assign n43196 = n13555 & n43195 ;
  assign n43197 = ~n43194 & ~n43196 ;
  assign n43198 = \m6_data_i[15]_pad  & n13547 ;
  assign n43199 = n13564 & n43198 ;
  assign n43200 = \m2_data_i[15]_pad  & n13547 ;
  assign n43201 = n13540 & n43200 ;
  assign n43202 = ~n43199 & ~n43201 ;
  assign n43203 = n43197 & n43202 ;
  assign n43204 = \m5_data_i[15]_pad  & ~n13547 ;
  assign n43205 = n13555 & n43204 ;
  assign n43206 = \m1_data_i[15]_pad  & ~n13547 ;
  assign n43207 = n13572 & n43206 ;
  assign n43208 = ~n43205 & ~n43207 ;
  assign n43209 = \m0_data_i[15]_pad  & n13547 ;
  assign n43210 = n13572 & n43209 ;
  assign n43211 = \m7_data_i[15]_pad  & ~n13547 ;
  assign n43212 = n13564 & n43211 ;
  assign n43213 = ~n43210 & ~n43212 ;
  assign n43214 = n43208 & n43213 ;
  assign n43215 = n43203 & n43214 ;
  assign n43216 = \m3_data_i[16]_pad  & ~n13547 ;
  assign n43217 = n13540 & n43216 ;
  assign n43218 = \m4_data_i[16]_pad  & n13547 ;
  assign n43219 = n13555 & n43218 ;
  assign n43220 = ~n43217 & ~n43219 ;
  assign n43221 = \m6_data_i[16]_pad  & n13547 ;
  assign n43222 = n13564 & n43221 ;
  assign n43223 = \m2_data_i[16]_pad  & n13547 ;
  assign n43224 = n13540 & n43223 ;
  assign n43225 = ~n43222 & ~n43224 ;
  assign n43226 = n43220 & n43225 ;
  assign n43227 = \m5_data_i[16]_pad  & ~n13547 ;
  assign n43228 = n13555 & n43227 ;
  assign n43229 = \m1_data_i[16]_pad  & ~n13547 ;
  assign n43230 = n13572 & n43229 ;
  assign n43231 = ~n43228 & ~n43230 ;
  assign n43232 = \m0_data_i[16]_pad  & n13547 ;
  assign n43233 = n13572 & n43232 ;
  assign n43234 = \m7_data_i[16]_pad  & ~n13547 ;
  assign n43235 = n13564 & n43234 ;
  assign n43236 = ~n43233 & ~n43235 ;
  assign n43237 = n43231 & n43236 ;
  assign n43238 = n43226 & n43237 ;
  assign n43239 = \m3_data_i[17]_pad  & ~n13547 ;
  assign n43240 = n13540 & n43239 ;
  assign n43241 = \m4_data_i[17]_pad  & n13547 ;
  assign n43242 = n13555 & n43241 ;
  assign n43243 = ~n43240 & ~n43242 ;
  assign n43244 = \m6_data_i[17]_pad  & n13547 ;
  assign n43245 = n13564 & n43244 ;
  assign n43246 = \m2_data_i[17]_pad  & n13547 ;
  assign n43247 = n13540 & n43246 ;
  assign n43248 = ~n43245 & ~n43247 ;
  assign n43249 = n43243 & n43248 ;
  assign n43250 = \m5_data_i[17]_pad  & ~n13547 ;
  assign n43251 = n13555 & n43250 ;
  assign n43252 = \m1_data_i[17]_pad  & ~n13547 ;
  assign n43253 = n13572 & n43252 ;
  assign n43254 = ~n43251 & ~n43253 ;
  assign n43255 = \m0_data_i[17]_pad  & n13547 ;
  assign n43256 = n13572 & n43255 ;
  assign n43257 = \m7_data_i[17]_pad  & ~n13547 ;
  assign n43258 = n13564 & n43257 ;
  assign n43259 = ~n43256 & ~n43258 ;
  assign n43260 = n43254 & n43259 ;
  assign n43261 = n43249 & n43260 ;
  assign n43262 = \m3_data_i[18]_pad  & ~n13547 ;
  assign n43263 = n13540 & n43262 ;
  assign n43264 = \m4_data_i[18]_pad  & n13547 ;
  assign n43265 = n13555 & n43264 ;
  assign n43266 = ~n43263 & ~n43265 ;
  assign n43267 = \m6_data_i[18]_pad  & n13547 ;
  assign n43268 = n13564 & n43267 ;
  assign n43269 = \m2_data_i[18]_pad  & n13547 ;
  assign n43270 = n13540 & n43269 ;
  assign n43271 = ~n43268 & ~n43270 ;
  assign n43272 = n43266 & n43271 ;
  assign n43273 = \m5_data_i[18]_pad  & ~n13547 ;
  assign n43274 = n13555 & n43273 ;
  assign n43275 = \m1_data_i[18]_pad  & ~n13547 ;
  assign n43276 = n13572 & n43275 ;
  assign n43277 = ~n43274 & ~n43276 ;
  assign n43278 = \m0_data_i[18]_pad  & n13547 ;
  assign n43279 = n13572 & n43278 ;
  assign n43280 = \m7_data_i[18]_pad  & ~n13547 ;
  assign n43281 = n13564 & n43280 ;
  assign n43282 = ~n43279 & ~n43281 ;
  assign n43283 = n43277 & n43282 ;
  assign n43284 = n43272 & n43283 ;
  assign n43285 = \m3_data_i[19]_pad  & ~n13547 ;
  assign n43286 = n13540 & n43285 ;
  assign n43287 = \m4_data_i[19]_pad  & n13547 ;
  assign n43288 = n13555 & n43287 ;
  assign n43289 = ~n43286 & ~n43288 ;
  assign n43290 = \m6_data_i[19]_pad  & n13547 ;
  assign n43291 = n13564 & n43290 ;
  assign n43292 = \m2_data_i[19]_pad  & n13547 ;
  assign n43293 = n13540 & n43292 ;
  assign n43294 = ~n43291 & ~n43293 ;
  assign n43295 = n43289 & n43294 ;
  assign n43296 = \m5_data_i[19]_pad  & ~n13547 ;
  assign n43297 = n13555 & n43296 ;
  assign n43298 = \m1_data_i[19]_pad  & ~n13547 ;
  assign n43299 = n13572 & n43298 ;
  assign n43300 = ~n43297 & ~n43299 ;
  assign n43301 = \m0_data_i[19]_pad  & n13547 ;
  assign n43302 = n13572 & n43301 ;
  assign n43303 = \m7_data_i[19]_pad  & ~n13547 ;
  assign n43304 = n13564 & n43303 ;
  assign n43305 = ~n43302 & ~n43304 ;
  assign n43306 = n43300 & n43305 ;
  assign n43307 = n43295 & n43306 ;
  assign n43308 = \m1_data_i[1]_pad  & ~n13547 ;
  assign n43309 = n13572 & n43308 ;
  assign n43310 = \m2_data_i[1]_pad  & n13547 ;
  assign n43311 = n13540 & n43310 ;
  assign n43312 = ~n43309 & ~n43311 ;
  assign n43313 = \m6_data_i[1]_pad  & n13547 ;
  assign n43314 = n13564 & n43313 ;
  assign n43315 = \m7_data_i[1]_pad  & ~n13547 ;
  assign n43316 = n13564 & n43315 ;
  assign n43317 = ~n43314 & ~n43316 ;
  assign n43318 = n43312 & n43317 ;
  assign n43319 = \m5_data_i[1]_pad  & ~n13547 ;
  assign n43320 = n13555 & n43319 ;
  assign n43321 = \m0_data_i[1]_pad  & n13547 ;
  assign n43322 = n13572 & n43321 ;
  assign n43323 = ~n43320 & ~n43322 ;
  assign n43324 = \m3_data_i[1]_pad  & ~n13547 ;
  assign n43325 = n13540 & n43324 ;
  assign n43326 = \m4_data_i[1]_pad  & n13547 ;
  assign n43327 = n13555 & n43326 ;
  assign n43328 = ~n43325 & ~n43327 ;
  assign n43329 = n43323 & n43328 ;
  assign n43330 = n43318 & n43329 ;
  assign n43331 = \m3_data_i[20]_pad  & ~n13547 ;
  assign n43332 = n13540 & n43331 ;
  assign n43333 = \m4_data_i[20]_pad  & n13547 ;
  assign n43334 = n13555 & n43333 ;
  assign n43335 = ~n43332 & ~n43334 ;
  assign n43336 = \m6_data_i[20]_pad  & n13547 ;
  assign n43337 = n13564 & n43336 ;
  assign n43338 = \m2_data_i[20]_pad  & n13547 ;
  assign n43339 = n13540 & n43338 ;
  assign n43340 = ~n43337 & ~n43339 ;
  assign n43341 = n43335 & n43340 ;
  assign n43342 = \m5_data_i[20]_pad  & ~n13547 ;
  assign n43343 = n13555 & n43342 ;
  assign n43344 = \m1_data_i[20]_pad  & ~n13547 ;
  assign n43345 = n13572 & n43344 ;
  assign n43346 = ~n43343 & ~n43345 ;
  assign n43347 = \m0_data_i[20]_pad  & n13547 ;
  assign n43348 = n13572 & n43347 ;
  assign n43349 = \m7_data_i[20]_pad  & ~n13547 ;
  assign n43350 = n13564 & n43349 ;
  assign n43351 = ~n43348 & ~n43350 ;
  assign n43352 = n43346 & n43351 ;
  assign n43353 = n43341 & n43352 ;
  assign n43354 = \m3_data_i[21]_pad  & ~n13547 ;
  assign n43355 = n13540 & n43354 ;
  assign n43356 = \m4_data_i[21]_pad  & n13547 ;
  assign n43357 = n13555 & n43356 ;
  assign n43358 = ~n43355 & ~n43357 ;
  assign n43359 = \m6_data_i[21]_pad  & n13547 ;
  assign n43360 = n13564 & n43359 ;
  assign n43361 = \m2_data_i[21]_pad  & n13547 ;
  assign n43362 = n13540 & n43361 ;
  assign n43363 = ~n43360 & ~n43362 ;
  assign n43364 = n43358 & n43363 ;
  assign n43365 = \m5_data_i[21]_pad  & ~n13547 ;
  assign n43366 = n13555 & n43365 ;
  assign n43367 = \m1_data_i[21]_pad  & ~n13547 ;
  assign n43368 = n13572 & n43367 ;
  assign n43369 = ~n43366 & ~n43368 ;
  assign n43370 = \m0_data_i[21]_pad  & n13547 ;
  assign n43371 = n13572 & n43370 ;
  assign n43372 = \m7_data_i[21]_pad  & ~n13547 ;
  assign n43373 = n13564 & n43372 ;
  assign n43374 = ~n43371 & ~n43373 ;
  assign n43375 = n43369 & n43374 ;
  assign n43376 = n43364 & n43375 ;
  assign n43377 = \m3_data_i[22]_pad  & ~n13547 ;
  assign n43378 = n13540 & n43377 ;
  assign n43379 = \m4_data_i[22]_pad  & n13547 ;
  assign n43380 = n13555 & n43379 ;
  assign n43381 = ~n43378 & ~n43380 ;
  assign n43382 = \m6_data_i[22]_pad  & n13547 ;
  assign n43383 = n13564 & n43382 ;
  assign n43384 = \m2_data_i[22]_pad  & n13547 ;
  assign n43385 = n13540 & n43384 ;
  assign n43386 = ~n43383 & ~n43385 ;
  assign n43387 = n43381 & n43386 ;
  assign n43388 = \m5_data_i[22]_pad  & ~n13547 ;
  assign n43389 = n13555 & n43388 ;
  assign n43390 = \m1_data_i[22]_pad  & ~n13547 ;
  assign n43391 = n13572 & n43390 ;
  assign n43392 = ~n43389 & ~n43391 ;
  assign n43393 = \m0_data_i[22]_pad  & n13547 ;
  assign n43394 = n13572 & n43393 ;
  assign n43395 = \m7_data_i[22]_pad  & ~n13547 ;
  assign n43396 = n13564 & n43395 ;
  assign n43397 = ~n43394 & ~n43396 ;
  assign n43398 = n43392 & n43397 ;
  assign n43399 = n43387 & n43398 ;
  assign n43400 = \m6_data_i[23]_pad  & n13547 ;
  assign n43401 = n13564 & n43400 ;
  assign n43402 = \m5_data_i[23]_pad  & ~n13547 ;
  assign n43403 = n13555 & n43402 ;
  assign n43404 = ~n43401 & ~n43403 ;
  assign n43405 = \m0_data_i[23]_pad  & n13547 ;
  assign n43406 = n13572 & n43405 ;
  assign n43407 = \m4_data_i[23]_pad  & n13547 ;
  assign n43408 = n13555 & n43407 ;
  assign n43409 = ~n43406 & ~n43408 ;
  assign n43410 = n43404 & n43409 ;
  assign n43411 = \m7_data_i[23]_pad  & ~n13547 ;
  assign n43412 = n13564 & n43411 ;
  assign n43413 = \m3_data_i[23]_pad  & ~n13547 ;
  assign n43414 = n13540 & n43413 ;
  assign n43415 = ~n43412 & ~n43414 ;
  assign n43416 = \m1_data_i[23]_pad  & ~n13547 ;
  assign n43417 = n13572 & n43416 ;
  assign n43418 = \m2_data_i[23]_pad  & n13547 ;
  assign n43419 = n13540 & n43418 ;
  assign n43420 = ~n43417 & ~n43419 ;
  assign n43421 = n43415 & n43420 ;
  assign n43422 = n43410 & n43421 ;
  assign n43423 = \m3_data_i[24]_pad  & ~n13547 ;
  assign n43424 = n13540 & n43423 ;
  assign n43425 = \m4_data_i[24]_pad  & n13547 ;
  assign n43426 = n13555 & n43425 ;
  assign n43427 = ~n43424 & ~n43426 ;
  assign n43428 = \m6_data_i[24]_pad  & n13547 ;
  assign n43429 = n13564 & n43428 ;
  assign n43430 = \m2_data_i[24]_pad  & n13547 ;
  assign n43431 = n13540 & n43430 ;
  assign n43432 = ~n43429 & ~n43431 ;
  assign n43433 = n43427 & n43432 ;
  assign n43434 = \m5_data_i[24]_pad  & ~n13547 ;
  assign n43435 = n13555 & n43434 ;
  assign n43436 = \m1_data_i[24]_pad  & ~n13547 ;
  assign n43437 = n13572 & n43436 ;
  assign n43438 = ~n43435 & ~n43437 ;
  assign n43439 = \m0_data_i[24]_pad  & n13547 ;
  assign n43440 = n13572 & n43439 ;
  assign n43441 = \m7_data_i[24]_pad  & ~n13547 ;
  assign n43442 = n13564 & n43441 ;
  assign n43443 = ~n43440 & ~n43442 ;
  assign n43444 = n43438 & n43443 ;
  assign n43445 = n43433 & n43444 ;
  assign n43446 = \m3_data_i[25]_pad  & ~n13547 ;
  assign n43447 = n13540 & n43446 ;
  assign n43448 = \m4_data_i[25]_pad  & n13547 ;
  assign n43449 = n13555 & n43448 ;
  assign n43450 = ~n43447 & ~n43449 ;
  assign n43451 = \m6_data_i[25]_pad  & n13547 ;
  assign n43452 = n13564 & n43451 ;
  assign n43453 = \m2_data_i[25]_pad  & n13547 ;
  assign n43454 = n13540 & n43453 ;
  assign n43455 = ~n43452 & ~n43454 ;
  assign n43456 = n43450 & n43455 ;
  assign n43457 = \m5_data_i[25]_pad  & ~n13547 ;
  assign n43458 = n13555 & n43457 ;
  assign n43459 = \m1_data_i[25]_pad  & ~n13547 ;
  assign n43460 = n13572 & n43459 ;
  assign n43461 = ~n43458 & ~n43460 ;
  assign n43462 = \m0_data_i[25]_pad  & n13547 ;
  assign n43463 = n13572 & n43462 ;
  assign n43464 = \m7_data_i[25]_pad  & ~n13547 ;
  assign n43465 = n13564 & n43464 ;
  assign n43466 = ~n43463 & ~n43465 ;
  assign n43467 = n43461 & n43466 ;
  assign n43468 = n43456 & n43467 ;
  assign n43469 = \m3_data_i[26]_pad  & ~n13547 ;
  assign n43470 = n13540 & n43469 ;
  assign n43471 = \m4_data_i[26]_pad  & n13547 ;
  assign n43472 = n13555 & n43471 ;
  assign n43473 = ~n43470 & ~n43472 ;
  assign n43474 = \m6_data_i[26]_pad  & n13547 ;
  assign n43475 = n13564 & n43474 ;
  assign n43476 = \m2_data_i[26]_pad  & n13547 ;
  assign n43477 = n13540 & n43476 ;
  assign n43478 = ~n43475 & ~n43477 ;
  assign n43479 = n43473 & n43478 ;
  assign n43480 = \m5_data_i[26]_pad  & ~n13547 ;
  assign n43481 = n13555 & n43480 ;
  assign n43482 = \m1_data_i[26]_pad  & ~n13547 ;
  assign n43483 = n13572 & n43482 ;
  assign n43484 = ~n43481 & ~n43483 ;
  assign n43485 = \m0_data_i[26]_pad  & n13547 ;
  assign n43486 = n13572 & n43485 ;
  assign n43487 = \m7_data_i[26]_pad  & ~n13547 ;
  assign n43488 = n13564 & n43487 ;
  assign n43489 = ~n43486 & ~n43488 ;
  assign n43490 = n43484 & n43489 ;
  assign n43491 = n43479 & n43490 ;
  assign n43492 = \m3_data_i[27]_pad  & ~n13547 ;
  assign n43493 = n13540 & n43492 ;
  assign n43494 = \m4_data_i[27]_pad  & n13547 ;
  assign n43495 = n13555 & n43494 ;
  assign n43496 = ~n43493 & ~n43495 ;
  assign n43497 = \m6_data_i[27]_pad  & n13547 ;
  assign n43498 = n13564 & n43497 ;
  assign n43499 = \m2_data_i[27]_pad  & n13547 ;
  assign n43500 = n13540 & n43499 ;
  assign n43501 = ~n43498 & ~n43500 ;
  assign n43502 = n43496 & n43501 ;
  assign n43503 = \m5_data_i[27]_pad  & ~n13547 ;
  assign n43504 = n13555 & n43503 ;
  assign n43505 = \m1_data_i[27]_pad  & ~n13547 ;
  assign n43506 = n13572 & n43505 ;
  assign n43507 = ~n43504 & ~n43506 ;
  assign n43508 = \m0_data_i[27]_pad  & n13547 ;
  assign n43509 = n13572 & n43508 ;
  assign n43510 = \m7_data_i[27]_pad  & ~n13547 ;
  assign n43511 = n13564 & n43510 ;
  assign n43512 = ~n43509 & ~n43511 ;
  assign n43513 = n43507 & n43512 ;
  assign n43514 = n43502 & n43513 ;
  assign n43515 = \m3_data_i[28]_pad  & ~n13547 ;
  assign n43516 = n13540 & n43515 ;
  assign n43517 = \m4_data_i[28]_pad  & n13547 ;
  assign n43518 = n13555 & n43517 ;
  assign n43519 = ~n43516 & ~n43518 ;
  assign n43520 = \m6_data_i[28]_pad  & n13547 ;
  assign n43521 = n13564 & n43520 ;
  assign n43522 = \m2_data_i[28]_pad  & n13547 ;
  assign n43523 = n13540 & n43522 ;
  assign n43524 = ~n43521 & ~n43523 ;
  assign n43525 = n43519 & n43524 ;
  assign n43526 = \m5_data_i[28]_pad  & ~n13547 ;
  assign n43527 = n13555 & n43526 ;
  assign n43528 = \m1_data_i[28]_pad  & ~n13547 ;
  assign n43529 = n13572 & n43528 ;
  assign n43530 = ~n43527 & ~n43529 ;
  assign n43531 = \m0_data_i[28]_pad  & n13547 ;
  assign n43532 = n13572 & n43531 ;
  assign n43533 = \m7_data_i[28]_pad  & ~n13547 ;
  assign n43534 = n13564 & n43533 ;
  assign n43535 = ~n43532 & ~n43534 ;
  assign n43536 = n43530 & n43535 ;
  assign n43537 = n43525 & n43536 ;
  assign n43538 = \m3_data_i[29]_pad  & ~n13547 ;
  assign n43539 = n13540 & n43538 ;
  assign n43540 = \m4_data_i[29]_pad  & n13547 ;
  assign n43541 = n13555 & n43540 ;
  assign n43542 = ~n43539 & ~n43541 ;
  assign n43543 = \m6_data_i[29]_pad  & n13547 ;
  assign n43544 = n13564 & n43543 ;
  assign n43545 = \m2_data_i[29]_pad  & n13547 ;
  assign n43546 = n13540 & n43545 ;
  assign n43547 = ~n43544 & ~n43546 ;
  assign n43548 = n43542 & n43547 ;
  assign n43549 = \m5_data_i[29]_pad  & ~n13547 ;
  assign n43550 = n13555 & n43549 ;
  assign n43551 = \m1_data_i[29]_pad  & ~n13547 ;
  assign n43552 = n13572 & n43551 ;
  assign n43553 = ~n43550 & ~n43552 ;
  assign n43554 = \m0_data_i[29]_pad  & n13547 ;
  assign n43555 = n13572 & n43554 ;
  assign n43556 = \m7_data_i[29]_pad  & ~n13547 ;
  assign n43557 = n13564 & n43556 ;
  assign n43558 = ~n43555 & ~n43557 ;
  assign n43559 = n43553 & n43558 ;
  assign n43560 = n43548 & n43559 ;
  assign n43561 = \m3_data_i[2]_pad  & ~n13547 ;
  assign n43562 = n13540 & n43561 ;
  assign n43563 = \m4_data_i[2]_pad  & n13547 ;
  assign n43564 = n13555 & n43563 ;
  assign n43565 = ~n43562 & ~n43564 ;
  assign n43566 = \m0_data_i[2]_pad  & n13547 ;
  assign n43567 = n13572 & n43566 ;
  assign n43568 = \m5_data_i[2]_pad  & ~n13547 ;
  assign n43569 = n13555 & n43568 ;
  assign n43570 = ~n43567 & ~n43569 ;
  assign n43571 = n43565 & n43570 ;
  assign n43572 = \m7_data_i[2]_pad  & ~n13547 ;
  assign n43573 = n13564 & n43572 ;
  assign n43574 = \m6_data_i[2]_pad  & n13547 ;
  assign n43575 = n13564 & n43574 ;
  assign n43576 = ~n43573 & ~n43575 ;
  assign n43577 = \m1_data_i[2]_pad  & ~n13547 ;
  assign n43578 = n13572 & n43577 ;
  assign n43579 = \m2_data_i[2]_pad  & n13547 ;
  assign n43580 = n13540 & n43579 ;
  assign n43581 = ~n43578 & ~n43580 ;
  assign n43582 = n43576 & n43581 ;
  assign n43583 = n43571 & n43582 ;
  assign n43584 = \m3_data_i[30]_pad  & ~n13547 ;
  assign n43585 = n13540 & n43584 ;
  assign n43586 = \m4_data_i[30]_pad  & n13547 ;
  assign n43587 = n13555 & n43586 ;
  assign n43588 = ~n43585 & ~n43587 ;
  assign n43589 = \m6_data_i[30]_pad  & n13547 ;
  assign n43590 = n13564 & n43589 ;
  assign n43591 = \m2_data_i[30]_pad  & n13547 ;
  assign n43592 = n13540 & n43591 ;
  assign n43593 = ~n43590 & ~n43592 ;
  assign n43594 = n43588 & n43593 ;
  assign n43595 = \m5_data_i[30]_pad  & ~n13547 ;
  assign n43596 = n13555 & n43595 ;
  assign n43597 = \m1_data_i[30]_pad  & ~n13547 ;
  assign n43598 = n13572 & n43597 ;
  assign n43599 = ~n43596 & ~n43598 ;
  assign n43600 = \m0_data_i[30]_pad  & n13547 ;
  assign n43601 = n13572 & n43600 ;
  assign n43602 = \m7_data_i[30]_pad  & ~n13547 ;
  assign n43603 = n13564 & n43602 ;
  assign n43604 = ~n43601 & ~n43603 ;
  assign n43605 = n43599 & n43604 ;
  assign n43606 = n43594 & n43605 ;
  assign n43607 = \m3_data_i[31]_pad  & ~n13547 ;
  assign n43608 = n13540 & n43607 ;
  assign n43609 = \m4_data_i[31]_pad  & n13547 ;
  assign n43610 = n13555 & n43609 ;
  assign n43611 = ~n43608 & ~n43610 ;
  assign n43612 = \m6_data_i[31]_pad  & n13547 ;
  assign n43613 = n13564 & n43612 ;
  assign n43614 = \m2_data_i[31]_pad  & n13547 ;
  assign n43615 = n13540 & n43614 ;
  assign n43616 = ~n43613 & ~n43615 ;
  assign n43617 = n43611 & n43616 ;
  assign n43618 = \m5_data_i[31]_pad  & ~n13547 ;
  assign n43619 = n13555 & n43618 ;
  assign n43620 = \m1_data_i[31]_pad  & ~n13547 ;
  assign n43621 = n13572 & n43620 ;
  assign n43622 = ~n43619 & ~n43621 ;
  assign n43623 = \m0_data_i[31]_pad  & n13547 ;
  assign n43624 = n13572 & n43623 ;
  assign n43625 = \m7_data_i[31]_pad  & ~n13547 ;
  assign n43626 = n13564 & n43625 ;
  assign n43627 = ~n43624 & ~n43626 ;
  assign n43628 = n43622 & n43627 ;
  assign n43629 = n43617 & n43628 ;
  assign n43630 = \m3_data_i[3]_pad  & ~n13547 ;
  assign n43631 = n13540 & n43630 ;
  assign n43632 = \m4_data_i[3]_pad  & n13547 ;
  assign n43633 = n13555 & n43632 ;
  assign n43634 = ~n43631 & ~n43633 ;
  assign n43635 = \m1_data_i[3]_pad  & ~n13547 ;
  assign n43636 = n13572 & n43635 ;
  assign n43637 = \m7_data_i[3]_pad  & ~n13547 ;
  assign n43638 = n13564 & n43637 ;
  assign n43639 = ~n43636 & ~n43638 ;
  assign n43640 = n43634 & n43639 ;
  assign n43641 = \m2_data_i[3]_pad  & n13547 ;
  assign n43642 = n13540 & n43641 ;
  assign n43643 = \m0_data_i[3]_pad  & n13547 ;
  assign n43644 = n13572 & n43643 ;
  assign n43645 = ~n43642 & ~n43644 ;
  assign n43646 = \m6_data_i[3]_pad  & n13547 ;
  assign n43647 = n13564 & n43646 ;
  assign n43648 = \m5_data_i[3]_pad  & ~n13547 ;
  assign n43649 = n13555 & n43648 ;
  assign n43650 = ~n43647 & ~n43649 ;
  assign n43651 = n43645 & n43650 ;
  assign n43652 = n43640 & n43651 ;
  assign n43653 = \m3_data_i[4]_pad  & ~n13547 ;
  assign n43654 = n13540 & n43653 ;
  assign n43655 = \m4_data_i[4]_pad  & n13547 ;
  assign n43656 = n13555 & n43655 ;
  assign n43657 = ~n43654 & ~n43656 ;
  assign n43658 = \m1_data_i[4]_pad  & ~n13547 ;
  assign n43659 = n13572 & n43658 ;
  assign n43660 = \m7_data_i[4]_pad  & ~n13547 ;
  assign n43661 = n13564 & n43660 ;
  assign n43662 = ~n43659 & ~n43661 ;
  assign n43663 = n43657 & n43662 ;
  assign n43664 = \m2_data_i[4]_pad  & n13547 ;
  assign n43665 = n13540 & n43664 ;
  assign n43666 = \m0_data_i[4]_pad  & n13547 ;
  assign n43667 = n13572 & n43666 ;
  assign n43668 = ~n43665 & ~n43667 ;
  assign n43669 = \m6_data_i[4]_pad  & n13547 ;
  assign n43670 = n13564 & n43669 ;
  assign n43671 = \m5_data_i[4]_pad  & ~n13547 ;
  assign n43672 = n13555 & n43671 ;
  assign n43673 = ~n43670 & ~n43672 ;
  assign n43674 = n43668 & n43673 ;
  assign n43675 = n43663 & n43674 ;
  assign n43676 = \m3_data_i[5]_pad  & ~n13547 ;
  assign n43677 = n13540 & n43676 ;
  assign n43678 = \m4_data_i[5]_pad  & n13547 ;
  assign n43679 = n13555 & n43678 ;
  assign n43680 = ~n43677 & ~n43679 ;
  assign n43681 = \m6_data_i[5]_pad  & n13547 ;
  assign n43682 = n13564 & n43681 ;
  assign n43683 = \m2_data_i[5]_pad  & n13547 ;
  assign n43684 = n13540 & n43683 ;
  assign n43685 = ~n43682 & ~n43684 ;
  assign n43686 = n43680 & n43685 ;
  assign n43687 = \m5_data_i[5]_pad  & ~n13547 ;
  assign n43688 = n13555 & n43687 ;
  assign n43689 = \m1_data_i[5]_pad  & ~n13547 ;
  assign n43690 = n13572 & n43689 ;
  assign n43691 = ~n43688 & ~n43690 ;
  assign n43692 = \m0_data_i[5]_pad  & n13547 ;
  assign n43693 = n13572 & n43692 ;
  assign n43694 = \m7_data_i[5]_pad  & ~n13547 ;
  assign n43695 = n13564 & n43694 ;
  assign n43696 = ~n43693 & ~n43695 ;
  assign n43697 = n43691 & n43696 ;
  assign n43698 = n43686 & n43697 ;
  assign n43699 = \m3_data_i[6]_pad  & ~n13547 ;
  assign n43700 = n13540 & n43699 ;
  assign n43701 = \m4_data_i[6]_pad  & n13547 ;
  assign n43702 = n13555 & n43701 ;
  assign n43703 = ~n43700 & ~n43702 ;
  assign n43704 = \m6_data_i[6]_pad  & n13547 ;
  assign n43705 = n13564 & n43704 ;
  assign n43706 = \m2_data_i[6]_pad  & n13547 ;
  assign n43707 = n13540 & n43706 ;
  assign n43708 = ~n43705 & ~n43707 ;
  assign n43709 = n43703 & n43708 ;
  assign n43710 = \m5_data_i[6]_pad  & ~n13547 ;
  assign n43711 = n13555 & n43710 ;
  assign n43712 = \m1_data_i[6]_pad  & ~n13547 ;
  assign n43713 = n13572 & n43712 ;
  assign n43714 = ~n43711 & ~n43713 ;
  assign n43715 = \m0_data_i[6]_pad  & n13547 ;
  assign n43716 = n13572 & n43715 ;
  assign n43717 = \m7_data_i[6]_pad  & ~n13547 ;
  assign n43718 = n13564 & n43717 ;
  assign n43719 = ~n43716 & ~n43718 ;
  assign n43720 = n43714 & n43719 ;
  assign n43721 = n43709 & n43720 ;
  assign n43722 = \m3_data_i[7]_pad  & ~n13547 ;
  assign n43723 = n13540 & n43722 ;
  assign n43724 = \m4_data_i[7]_pad  & n13547 ;
  assign n43725 = n13555 & n43724 ;
  assign n43726 = ~n43723 & ~n43725 ;
  assign n43727 = \m6_data_i[7]_pad  & n13547 ;
  assign n43728 = n13564 & n43727 ;
  assign n43729 = \m2_data_i[7]_pad  & n13547 ;
  assign n43730 = n13540 & n43729 ;
  assign n43731 = ~n43728 & ~n43730 ;
  assign n43732 = n43726 & n43731 ;
  assign n43733 = \m5_data_i[7]_pad  & ~n13547 ;
  assign n43734 = n13555 & n43733 ;
  assign n43735 = \m1_data_i[7]_pad  & ~n13547 ;
  assign n43736 = n13572 & n43735 ;
  assign n43737 = ~n43734 & ~n43736 ;
  assign n43738 = \m0_data_i[7]_pad  & n13547 ;
  assign n43739 = n13572 & n43738 ;
  assign n43740 = \m7_data_i[7]_pad  & ~n13547 ;
  assign n43741 = n13564 & n43740 ;
  assign n43742 = ~n43739 & ~n43741 ;
  assign n43743 = n43737 & n43742 ;
  assign n43744 = n43732 & n43743 ;
  assign n43745 = \m3_data_i[8]_pad  & ~n13547 ;
  assign n43746 = n13540 & n43745 ;
  assign n43747 = \m4_data_i[8]_pad  & n13547 ;
  assign n43748 = n13555 & n43747 ;
  assign n43749 = ~n43746 & ~n43748 ;
  assign n43750 = \m6_data_i[8]_pad  & n13547 ;
  assign n43751 = n13564 & n43750 ;
  assign n43752 = \m2_data_i[8]_pad  & n13547 ;
  assign n43753 = n13540 & n43752 ;
  assign n43754 = ~n43751 & ~n43753 ;
  assign n43755 = n43749 & n43754 ;
  assign n43756 = \m5_data_i[8]_pad  & ~n13547 ;
  assign n43757 = n13555 & n43756 ;
  assign n43758 = \m1_data_i[8]_pad  & ~n13547 ;
  assign n43759 = n13572 & n43758 ;
  assign n43760 = ~n43757 & ~n43759 ;
  assign n43761 = \m0_data_i[8]_pad  & n13547 ;
  assign n43762 = n13572 & n43761 ;
  assign n43763 = \m7_data_i[8]_pad  & ~n13547 ;
  assign n43764 = n13564 & n43763 ;
  assign n43765 = ~n43762 & ~n43764 ;
  assign n43766 = n43760 & n43765 ;
  assign n43767 = n43755 & n43766 ;
  assign n43768 = \m3_data_i[9]_pad  & ~n13547 ;
  assign n43769 = n13540 & n43768 ;
  assign n43770 = \m4_data_i[9]_pad  & n13547 ;
  assign n43771 = n13555 & n43770 ;
  assign n43772 = ~n43769 & ~n43771 ;
  assign n43773 = \m6_data_i[9]_pad  & n13547 ;
  assign n43774 = n13564 & n43773 ;
  assign n43775 = \m2_data_i[9]_pad  & n13547 ;
  assign n43776 = n13540 & n43775 ;
  assign n43777 = ~n43774 & ~n43776 ;
  assign n43778 = n43772 & n43777 ;
  assign n43779 = \m5_data_i[9]_pad  & ~n13547 ;
  assign n43780 = n13555 & n43779 ;
  assign n43781 = \m1_data_i[9]_pad  & ~n13547 ;
  assign n43782 = n13572 & n43781 ;
  assign n43783 = ~n43780 & ~n43782 ;
  assign n43784 = \m0_data_i[9]_pad  & n13547 ;
  assign n43785 = n13572 & n43784 ;
  assign n43786 = \m7_data_i[9]_pad  & ~n13547 ;
  assign n43787 = n13564 & n43786 ;
  assign n43788 = ~n43785 & ~n43787 ;
  assign n43789 = n43783 & n43788 ;
  assign n43790 = n43778 & n43789 ;
  assign n43791 = \m1_sel_i[0]_pad  & ~n13547 ;
  assign n43792 = n13572 & n43791 ;
  assign n43793 = \m2_sel_i[0]_pad  & n13547 ;
  assign n43794 = n13540 & n43793 ;
  assign n43795 = ~n43792 & ~n43794 ;
  assign n43796 = \m0_sel_i[0]_pad  & n13547 ;
  assign n43797 = n13572 & n43796 ;
  assign n43798 = \m4_sel_i[0]_pad  & n13547 ;
  assign n43799 = n13555 & n43798 ;
  assign n43800 = ~n43797 & ~n43799 ;
  assign n43801 = n43795 & n43800 ;
  assign n43802 = \m7_sel_i[0]_pad  & ~n13547 ;
  assign n43803 = n13564 & n43802 ;
  assign n43804 = \m3_sel_i[0]_pad  & ~n13547 ;
  assign n43805 = n13540 & n43804 ;
  assign n43806 = ~n43803 & ~n43805 ;
  assign n43807 = \m6_sel_i[0]_pad  & n13547 ;
  assign n43808 = n13564 & n43807 ;
  assign n43809 = \m5_sel_i[0]_pad  & ~n13547 ;
  assign n43810 = n13555 & n43809 ;
  assign n43811 = ~n43808 & ~n43810 ;
  assign n43812 = n43806 & n43811 ;
  assign n43813 = n43801 & n43812 ;
  assign n43814 = \m0_sel_i[1]_pad  & n13547 ;
  assign n43815 = n13572 & n43814 ;
  assign n43816 = \m7_sel_i[1]_pad  & ~n13547 ;
  assign n43817 = n13564 & n43816 ;
  assign n43818 = ~n43815 & ~n43817 ;
  assign n43819 = \m3_sel_i[1]_pad  & ~n13547 ;
  assign n43820 = n13540 & n43819 ;
  assign n43821 = \m2_sel_i[1]_pad  & n13547 ;
  assign n43822 = n13540 & n43821 ;
  assign n43823 = ~n43820 & ~n43822 ;
  assign n43824 = n43818 & n43823 ;
  assign n43825 = \m4_sel_i[1]_pad  & n13547 ;
  assign n43826 = n13555 & n43825 ;
  assign n43827 = \m1_sel_i[1]_pad  & ~n13547 ;
  assign n43828 = n13572 & n43827 ;
  assign n43829 = ~n43826 & ~n43828 ;
  assign n43830 = \m6_sel_i[1]_pad  & n13547 ;
  assign n43831 = n13564 & n43830 ;
  assign n43832 = \m5_sel_i[1]_pad  & ~n13547 ;
  assign n43833 = n13555 & n43832 ;
  assign n43834 = ~n43831 & ~n43833 ;
  assign n43835 = n43829 & n43834 ;
  assign n43836 = n43824 & n43835 ;
  assign n43837 = \m1_sel_i[2]_pad  & ~n13547 ;
  assign n43838 = n13572 & n43837 ;
  assign n43839 = \m2_sel_i[2]_pad  & n13547 ;
  assign n43840 = n13540 & n43839 ;
  assign n43841 = ~n43838 & ~n43840 ;
  assign n43842 = \m0_sel_i[2]_pad  & n13547 ;
  assign n43843 = n13572 & n43842 ;
  assign n43844 = \m4_sel_i[2]_pad  & n13547 ;
  assign n43845 = n13555 & n43844 ;
  assign n43846 = ~n43843 & ~n43845 ;
  assign n43847 = n43841 & n43846 ;
  assign n43848 = \m7_sel_i[2]_pad  & ~n13547 ;
  assign n43849 = n13564 & n43848 ;
  assign n43850 = \m3_sel_i[2]_pad  & ~n13547 ;
  assign n43851 = n13540 & n43850 ;
  assign n43852 = ~n43849 & ~n43851 ;
  assign n43853 = \m6_sel_i[2]_pad  & n13547 ;
  assign n43854 = n13564 & n43853 ;
  assign n43855 = \m5_sel_i[2]_pad  & ~n13547 ;
  assign n43856 = n13555 & n43855 ;
  assign n43857 = ~n43854 & ~n43856 ;
  assign n43858 = n43852 & n43857 ;
  assign n43859 = n43847 & n43858 ;
  assign n43860 = \m0_sel_i[3]_pad  & n13547 ;
  assign n43861 = n13572 & n43860 ;
  assign n43862 = \m7_sel_i[3]_pad  & ~n13547 ;
  assign n43863 = n13564 & n43862 ;
  assign n43864 = ~n43861 & ~n43863 ;
  assign n43865 = \m6_sel_i[3]_pad  & n13547 ;
  assign n43866 = n13564 & n43865 ;
  assign n43867 = \m2_sel_i[3]_pad  & n13547 ;
  assign n43868 = n13540 & n43867 ;
  assign n43869 = ~n43866 & ~n43868 ;
  assign n43870 = n43864 & n43869 ;
  assign n43871 = \m5_sel_i[3]_pad  & ~n13547 ;
  assign n43872 = n13555 & n43871 ;
  assign n43873 = \m1_sel_i[3]_pad  & ~n13547 ;
  assign n43874 = n13572 & n43873 ;
  assign n43875 = ~n43872 & ~n43874 ;
  assign n43876 = \m3_sel_i[3]_pad  & ~n13547 ;
  assign n43877 = n13540 & n43876 ;
  assign n43878 = \m4_sel_i[3]_pad  & n13547 ;
  assign n43879 = n13555 & n43878 ;
  assign n43880 = ~n43877 & ~n43879 ;
  assign n43881 = n43875 & n43880 ;
  assign n43882 = n43870 & n43881 ;
  assign n43883 = \m5_stb_i_pad  & n14983 ;
  assign n43884 = ~n13547 & n43883 ;
  assign n43885 = n13555 & n43884 ;
  assign n43886 = \m4_stb_i_pad  & n14954 ;
  assign n43887 = n13547 & n43886 ;
  assign n43888 = n13555 & n43887 ;
  assign n43889 = ~n43885 & ~n43888 ;
  assign n43890 = \m2_stb_i_pad  & n14879 ;
  assign n43891 = n13547 & n43890 ;
  assign n43892 = n13540 & n43891 ;
  assign n43893 = \m1_stb_i_pad  & n14829 ;
  assign n43894 = ~n13547 & n43893 ;
  assign n43895 = n13572 & n43894 ;
  assign n43896 = ~n43892 & ~n43895 ;
  assign n43897 = n43889 & n43896 ;
  assign n43898 = \m3_stb_i_pad  & n14757 ;
  assign n43899 = ~n13547 & n43898 ;
  assign n43900 = n13540 & n43899 ;
  assign n43901 = \m7_stb_i_pad  & n14675 ;
  assign n43902 = ~n13547 & n43901 ;
  assign n43903 = n13564 & n43902 ;
  assign n43904 = ~n43900 & ~n43903 ;
  assign n43905 = \m6_stb_i_pad  & n15034 ;
  assign n43906 = n13547 & n43905 ;
  assign n43907 = n13564 & n43906 ;
  assign n43908 = \m0_stb_i_pad  & n14778 ;
  assign n43909 = n13547 & n43908 ;
  assign n43910 = n13572 & n43909 ;
  assign n43911 = ~n43907 & ~n43910 ;
  assign n43912 = n43904 & n43911 ;
  assign n43913 = n43897 & n43912 ;
  assign n43914 = \m1_we_i_pad  & ~n13547 ;
  assign n43915 = n13572 & n43914 ;
  assign n43916 = \m2_we_i_pad  & n13547 ;
  assign n43917 = n13540 & n43916 ;
  assign n43918 = ~n43915 & ~n43917 ;
  assign n43919 = \m0_we_i_pad  & n13547 ;
  assign n43920 = n13572 & n43919 ;
  assign n43921 = \m4_we_i_pad  & n13547 ;
  assign n43922 = n13555 & n43921 ;
  assign n43923 = ~n43920 & ~n43922 ;
  assign n43924 = n43918 & n43923 ;
  assign n43925 = \m7_we_i_pad  & ~n13547 ;
  assign n43926 = n13564 & n43925 ;
  assign n43927 = \m3_we_i_pad  & ~n13547 ;
  assign n43928 = n13540 & n43927 ;
  assign n43929 = ~n43926 & ~n43928 ;
  assign n43930 = \m6_we_i_pad  & n13547 ;
  assign n43931 = n13564 & n43930 ;
  assign n43932 = \m5_we_i_pad  & ~n13547 ;
  assign n43933 = n13555 & n43932 ;
  assign n43934 = ~n43931 & ~n43933 ;
  assign n43935 = n43929 & n43934 ;
  assign n43936 = n43924 & n43935 ;
  assign n43937 = \m1_addr_i[0]_pad  & ~n13627 ;
  assign n43938 = n13620 & n43937 ;
  assign n43939 = \m2_addr_i[0]_pad  & n13627 ;
  assign n43940 = n13635 & n43939 ;
  assign n43941 = ~n43938 & ~n43940 ;
  assign n43942 = \m6_addr_i[0]_pad  & n13627 ;
  assign n43943 = n13644 & n43942 ;
  assign n43944 = \m7_addr_i[0]_pad  & ~n13627 ;
  assign n43945 = n13644 & n43944 ;
  assign n43946 = ~n43943 & ~n43945 ;
  assign n43947 = n43941 & n43946 ;
  assign n43948 = \m5_addr_i[0]_pad  & ~n13627 ;
  assign n43949 = n13652 & n43948 ;
  assign n43950 = \m0_addr_i[0]_pad  & n13627 ;
  assign n43951 = n13620 & n43950 ;
  assign n43952 = ~n43949 & ~n43951 ;
  assign n43953 = \m3_addr_i[0]_pad  & ~n13627 ;
  assign n43954 = n13635 & n43953 ;
  assign n43955 = \m4_addr_i[0]_pad  & n13627 ;
  assign n43956 = n13652 & n43955 ;
  assign n43957 = ~n43954 & ~n43956 ;
  assign n43958 = n43952 & n43957 ;
  assign n43959 = n43947 & n43958 ;
  assign n43960 = \m3_addr_i[10]_pad  & ~n13627 ;
  assign n43961 = n13635 & n43960 ;
  assign n43962 = \m4_addr_i[10]_pad  & n13627 ;
  assign n43963 = n13652 & n43962 ;
  assign n43964 = ~n43961 & ~n43963 ;
  assign n43965 = \m6_addr_i[10]_pad  & n13627 ;
  assign n43966 = n13644 & n43965 ;
  assign n43967 = \m2_addr_i[10]_pad  & n13627 ;
  assign n43968 = n13635 & n43967 ;
  assign n43969 = ~n43966 & ~n43968 ;
  assign n43970 = n43964 & n43969 ;
  assign n43971 = \m5_addr_i[10]_pad  & ~n13627 ;
  assign n43972 = n13652 & n43971 ;
  assign n43973 = \m1_addr_i[10]_pad  & ~n13627 ;
  assign n43974 = n13620 & n43973 ;
  assign n43975 = ~n43972 & ~n43974 ;
  assign n43976 = \m0_addr_i[10]_pad  & n13627 ;
  assign n43977 = n13620 & n43976 ;
  assign n43978 = \m7_addr_i[10]_pad  & ~n13627 ;
  assign n43979 = n13644 & n43978 ;
  assign n43980 = ~n43977 & ~n43979 ;
  assign n43981 = n43975 & n43980 ;
  assign n43982 = n43970 & n43981 ;
  assign n43983 = \m3_addr_i[11]_pad  & ~n13627 ;
  assign n43984 = n13635 & n43983 ;
  assign n43985 = \m4_addr_i[11]_pad  & n13627 ;
  assign n43986 = n13652 & n43985 ;
  assign n43987 = ~n43984 & ~n43986 ;
  assign n43988 = \m6_addr_i[11]_pad  & n13627 ;
  assign n43989 = n13644 & n43988 ;
  assign n43990 = \m2_addr_i[11]_pad  & n13627 ;
  assign n43991 = n13635 & n43990 ;
  assign n43992 = ~n43989 & ~n43991 ;
  assign n43993 = n43987 & n43992 ;
  assign n43994 = \m5_addr_i[11]_pad  & ~n13627 ;
  assign n43995 = n13652 & n43994 ;
  assign n43996 = \m1_addr_i[11]_pad  & ~n13627 ;
  assign n43997 = n13620 & n43996 ;
  assign n43998 = ~n43995 & ~n43997 ;
  assign n43999 = \m0_addr_i[11]_pad  & n13627 ;
  assign n44000 = n13620 & n43999 ;
  assign n44001 = \m7_addr_i[11]_pad  & ~n13627 ;
  assign n44002 = n13644 & n44001 ;
  assign n44003 = ~n44000 & ~n44002 ;
  assign n44004 = n43998 & n44003 ;
  assign n44005 = n43993 & n44004 ;
  assign n44006 = \m3_addr_i[12]_pad  & ~n13627 ;
  assign n44007 = n13635 & n44006 ;
  assign n44008 = \m4_addr_i[12]_pad  & n13627 ;
  assign n44009 = n13652 & n44008 ;
  assign n44010 = ~n44007 & ~n44009 ;
  assign n44011 = \m6_addr_i[12]_pad  & n13627 ;
  assign n44012 = n13644 & n44011 ;
  assign n44013 = \m7_addr_i[12]_pad  & ~n13627 ;
  assign n44014 = n13644 & n44013 ;
  assign n44015 = ~n44012 & ~n44014 ;
  assign n44016 = n44010 & n44015 ;
  assign n44017 = \m5_addr_i[12]_pad  & ~n13627 ;
  assign n44018 = n13652 & n44017 ;
  assign n44019 = \m0_addr_i[12]_pad  & n13627 ;
  assign n44020 = n13620 & n44019 ;
  assign n44021 = ~n44018 & ~n44020 ;
  assign n44022 = \m1_addr_i[12]_pad  & ~n13627 ;
  assign n44023 = n13620 & n44022 ;
  assign n44024 = \m2_addr_i[12]_pad  & n13627 ;
  assign n44025 = n13635 & n44024 ;
  assign n44026 = ~n44023 & ~n44025 ;
  assign n44027 = n44021 & n44026 ;
  assign n44028 = n44016 & n44027 ;
  assign n44029 = \m3_addr_i[13]_pad  & ~n13627 ;
  assign n44030 = n13635 & n44029 ;
  assign n44031 = \m4_addr_i[13]_pad  & n13627 ;
  assign n44032 = n13652 & n44031 ;
  assign n44033 = ~n44030 & ~n44032 ;
  assign n44034 = \m6_addr_i[13]_pad  & n13627 ;
  assign n44035 = n13644 & n44034 ;
  assign n44036 = \m2_addr_i[13]_pad  & n13627 ;
  assign n44037 = n13635 & n44036 ;
  assign n44038 = ~n44035 & ~n44037 ;
  assign n44039 = n44033 & n44038 ;
  assign n44040 = \m5_addr_i[13]_pad  & ~n13627 ;
  assign n44041 = n13652 & n44040 ;
  assign n44042 = \m1_addr_i[13]_pad  & ~n13627 ;
  assign n44043 = n13620 & n44042 ;
  assign n44044 = ~n44041 & ~n44043 ;
  assign n44045 = \m0_addr_i[13]_pad  & n13627 ;
  assign n44046 = n13620 & n44045 ;
  assign n44047 = \m7_addr_i[13]_pad  & ~n13627 ;
  assign n44048 = n13644 & n44047 ;
  assign n44049 = ~n44046 & ~n44048 ;
  assign n44050 = n44044 & n44049 ;
  assign n44051 = n44039 & n44050 ;
  assign n44052 = \m3_addr_i[14]_pad  & ~n13627 ;
  assign n44053 = n13635 & n44052 ;
  assign n44054 = \m4_addr_i[14]_pad  & n13627 ;
  assign n44055 = n13652 & n44054 ;
  assign n44056 = ~n44053 & ~n44055 ;
  assign n44057 = \m6_addr_i[14]_pad  & n13627 ;
  assign n44058 = n13644 & n44057 ;
  assign n44059 = \m2_addr_i[14]_pad  & n13627 ;
  assign n44060 = n13635 & n44059 ;
  assign n44061 = ~n44058 & ~n44060 ;
  assign n44062 = n44056 & n44061 ;
  assign n44063 = \m5_addr_i[14]_pad  & ~n13627 ;
  assign n44064 = n13652 & n44063 ;
  assign n44065 = \m1_addr_i[14]_pad  & ~n13627 ;
  assign n44066 = n13620 & n44065 ;
  assign n44067 = ~n44064 & ~n44066 ;
  assign n44068 = \m0_addr_i[14]_pad  & n13627 ;
  assign n44069 = n13620 & n44068 ;
  assign n44070 = \m7_addr_i[14]_pad  & ~n13627 ;
  assign n44071 = n13644 & n44070 ;
  assign n44072 = ~n44069 & ~n44071 ;
  assign n44073 = n44067 & n44072 ;
  assign n44074 = n44062 & n44073 ;
  assign n44075 = \m1_addr_i[15]_pad  & ~n13627 ;
  assign n44076 = n13620 & n44075 ;
  assign n44077 = \m2_addr_i[15]_pad  & n13627 ;
  assign n44078 = n13635 & n44077 ;
  assign n44079 = ~n44076 & ~n44078 ;
  assign n44080 = \m3_addr_i[15]_pad  & ~n13627 ;
  assign n44081 = n13635 & n44080 ;
  assign n44082 = \m7_addr_i[15]_pad  & ~n13627 ;
  assign n44083 = n13644 & n44082 ;
  assign n44084 = ~n44081 & ~n44083 ;
  assign n44085 = n44079 & n44084 ;
  assign n44086 = \m4_addr_i[15]_pad  & n13627 ;
  assign n44087 = n13652 & n44086 ;
  assign n44088 = \m0_addr_i[15]_pad  & n13627 ;
  assign n44089 = n13620 & n44088 ;
  assign n44090 = ~n44087 & ~n44089 ;
  assign n44091 = \m6_addr_i[15]_pad  & n13627 ;
  assign n44092 = n13644 & n44091 ;
  assign n44093 = \m5_addr_i[15]_pad  & ~n13627 ;
  assign n44094 = n13652 & n44093 ;
  assign n44095 = ~n44092 & ~n44094 ;
  assign n44096 = n44090 & n44095 ;
  assign n44097 = n44085 & n44096 ;
  assign n44098 = \m3_addr_i[16]_pad  & ~n13627 ;
  assign n44099 = n13635 & n44098 ;
  assign n44100 = \m4_addr_i[16]_pad  & n13627 ;
  assign n44101 = n13652 & n44100 ;
  assign n44102 = ~n44099 & ~n44101 ;
  assign n44103 = \m6_addr_i[16]_pad  & n13627 ;
  assign n44104 = n13644 & n44103 ;
  assign n44105 = \m2_addr_i[16]_pad  & n13627 ;
  assign n44106 = n13635 & n44105 ;
  assign n44107 = ~n44104 & ~n44106 ;
  assign n44108 = n44102 & n44107 ;
  assign n44109 = \m5_addr_i[16]_pad  & ~n13627 ;
  assign n44110 = n13652 & n44109 ;
  assign n44111 = \m1_addr_i[16]_pad  & ~n13627 ;
  assign n44112 = n13620 & n44111 ;
  assign n44113 = ~n44110 & ~n44112 ;
  assign n44114 = \m0_addr_i[16]_pad  & n13627 ;
  assign n44115 = n13620 & n44114 ;
  assign n44116 = \m7_addr_i[16]_pad  & ~n13627 ;
  assign n44117 = n13644 & n44116 ;
  assign n44118 = ~n44115 & ~n44117 ;
  assign n44119 = n44113 & n44118 ;
  assign n44120 = n44108 & n44119 ;
  assign n44121 = \m3_addr_i[17]_pad  & ~n13627 ;
  assign n44122 = n13635 & n44121 ;
  assign n44123 = \m4_addr_i[17]_pad  & n13627 ;
  assign n44124 = n13652 & n44123 ;
  assign n44125 = ~n44122 & ~n44124 ;
  assign n44126 = \m6_addr_i[17]_pad  & n13627 ;
  assign n44127 = n13644 & n44126 ;
  assign n44128 = \m2_addr_i[17]_pad  & n13627 ;
  assign n44129 = n13635 & n44128 ;
  assign n44130 = ~n44127 & ~n44129 ;
  assign n44131 = n44125 & n44130 ;
  assign n44132 = \m5_addr_i[17]_pad  & ~n13627 ;
  assign n44133 = n13652 & n44132 ;
  assign n44134 = \m1_addr_i[17]_pad  & ~n13627 ;
  assign n44135 = n13620 & n44134 ;
  assign n44136 = ~n44133 & ~n44135 ;
  assign n44137 = \m0_addr_i[17]_pad  & n13627 ;
  assign n44138 = n13620 & n44137 ;
  assign n44139 = \m7_addr_i[17]_pad  & ~n13627 ;
  assign n44140 = n13644 & n44139 ;
  assign n44141 = ~n44138 & ~n44140 ;
  assign n44142 = n44136 & n44141 ;
  assign n44143 = n44131 & n44142 ;
  assign n44144 = \m3_addr_i[18]_pad  & ~n13627 ;
  assign n44145 = n13635 & n44144 ;
  assign n44146 = \m4_addr_i[18]_pad  & n13627 ;
  assign n44147 = n13652 & n44146 ;
  assign n44148 = ~n44145 & ~n44147 ;
  assign n44149 = \m6_addr_i[18]_pad  & n13627 ;
  assign n44150 = n13644 & n44149 ;
  assign n44151 = \m2_addr_i[18]_pad  & n13627 ;
  assign n44152 = n13635 & n44151 ;
  assign n44153 = ~n44150 & ~n44152 ;
  assign n44154 = n44148 & n44153 ;
  assign n44155 = \m5_addr_i[18]_pad  & ~n13627 ;
  assign n44156 = n13652 & n44155 ;
  assign n44157 = \m1_addr_i[18]_pad  & ~n13627 ;
  assign n44158 = n13620 & n44157 ;
  assign n44159 = ~n44156 & ~n44158 ;
  assign n44160 = \m0_addr_i[18]_pad  & n13627 ;
  assign n44161 = n13620 & n44160 ;
  assign n44162 = \m7_addr_i[18]_pad  & ~n13627 ;
  assign n44163 = n13644 & n44162 ;
  assign n44164 = ~n44161 & ~n44163 ;
  assign n44165 = n44159 & n44164 ;
  assign n44166 = n44154 & n44165 ;
  assign n44167 = \m3_addr_i[19]_pad  & ~n13627 ;
  assign n44168 = n13635 & n44167 ;
  assign n44169 = \m4_addr_i[19]_pad  & n13627 ;
  assign n44170 = n13652 & n44169 ;
  assign n44171 = ~n44168 & ~n44170 ;
  assign n44172 = \m6_addr_i[19]_pad  & n13627 ;
  assign n44173 = n13644 & n44172 ;
  assign n44174 = \m2_addr_i[19]_pad  & n13627 ;
  assign n44175 = n13635 & n44174 ;
  assign n44176 = ~n44173 & ~n44175 ;
  assign n44177 = n44171 & n44176 ;
  assign n44178 = \m5_addr_i[19]_pad  & ~n13627 ;
  assign n44179 = n13652 & n44178 ;
  assign n44180 = \m1_addr_i[19]_pad  & ~n13627 ;
  assign n44181 = n13620 & n44180 ;
  assign n44182 = ~n44179 & ~n44181 ;
  assign n44183 = \m0_addr_i[19]_pad  & n13627 ;
  assign n44184 = n13620 & n44183 ;
  assign n44185 = \m7_addr_i[19]_pad  & ~n13627 ;
  assign n44186 = n13644 & n44185 ;
  assign n44187 = ~n44184 & ~n44186 ;
  assign n44188 = n44182 & n44187 ;
  assign n44189 = n44177 & n44188 ;
  assign n44190 = \m3_addr_i[1]_pad  & ~n13627 ;
  assign n44191 = n13635 & n44190 ;
  assign n44192 = \m4_addr_i[1]_pad  & n13627 ;
  assign n44193 = n13652 & n44192 ;
  assign n44194 = ~n44191 & ~n44193 ;
  assign n44195 = \m6_addr_i[1]_pad  & n13627 ;
  assign n44196 = n13644 & n44195 ;
  assign n44197 = \m7_addr_i[1]_pad  & ~n13627 ;
  assign n44198 = n13644 & n44197 ;
  assign n44199 = ~n44196 & ~n44198 ;
  assign n44200 = n44194 & n44199 ;
  assign n44201 = \m5_addr_i[1]_pad  & ~n13627 ;
  assign n44202 = n13652 & n44201 ;
  assign n44203 = \m0_addr_i[1]_pad  & n13627 ;
  assign n44204 = n13620 & n44203 ;
  assign n44205 = ~n44202 & ~n44204 ;
  assign n44206 = \m1_addr_i[1]_pad  & ~n13627 ;
  assign n44207 = n13620 & n44206 ;
  assign n44208 = \m2_addr_i[1]_pad  & n13627 ;
  assign n44209 = n13635 & n44208 ;
  assign n44210 = ~n44207 & ~n44209 ;
  assign n44211 = n44205 & n44210 ;
  assign n44212 = n44200 & n44211 ;
  assign n44213 = \m3_addr_i[20]_pad  & ~n13627 ;
  assign n44214 = n13635 & n44213 ;
  assign n44215 = \m4_addr_i[20]_pad  & n13627 ;
  assign n44216 = n13652 & n44215 ;
  assign n44217 = ~n44214 & ~n44216 ;
  assign n44218 = \m6_addr_i[20]_pad  & n13627 ;
  assign n44219 = n13644 & n44218 ;
  assign n44220 = \m2_addr_i[20]_pad  & n13627 ;
  assign n44221 = n13635 & n44220 ;
  assign n44222 = ~n44219 & ~n44221 ;
  assign n44223 = n44217 & n44222 ;
  assign n44224 = \m5_addr_i[20]_pad  & ~n13627 ;
  assign n44225 = n13652 & n44224 ;
  assign n44226 = \m1_addr_i[20]_pad  & ~n13627 ;
  assign n44227 = n13620 & n44226 ;
  assign n44228 = ~n44225 & ~n44227 ;
  assign n44229 = \m0_addr_i[20]_pad  & n13627 ;
  assign n44230 = n13620 & n44229 ;
  assign n44231 = \m7_addr_i[20]_pad  & ~n13627 ;
  assign n44232 = n13644 & n44231 ;
  assign n44233 = ~n44230 & ~n44232 ;
  assign n44234 = n44228 & n44233 ;
  assign n44235 = n44223 & n44234 ;
  assign n44236 = \m3_addr_i[21]_pad  & ~n13627 ;
  assign n44237 = n13635 & n44236 ;
  assign n44238 = \m4_addr_i[21]_pad  & n13627 ;
  assign n44239 = n13652 & n44238 ;
  assign n44240 = ~n44237 & ~n44239 ;
  assign n44241 = \m6_addr_i[21]_pad  & n13627 ;
  assign n44242 = n13644 & n44241 ;
  assign n44243 = \m2_addr_i[21]_pad  & n13627 ;
  assign n44244 = n13635 & n44243 ;
  assign n44245 = ~n44242 & ~n44244 ;
  assign n44246 = n44240 & n44245 ;
  assign n44247 = \m5_addr_i[21]_pad  & ~n13627 ;
  assign n44248 = n13652 & n44247 ;
  assign n44249 = \m1_addr_i[21]_pad  & ~n13627 ;
  assign n44250 = n13620 & n44249 ;
  assign n44251 = ~n44248 & ~n44250 ;
  assign n44252 = \m0_addr_i[21]_pad  & n13627 ;
  assign n44253 = n13620 & n44252 ;
  assign n44254 = \m7_addr_i[21]_pad  & ~n13627 ;
  assign n44255 = n13644 & n44254 ;
  assign n44256 = ~n44253 & ~n44255 ;
  assign n44257 = n44251 & n44256 ;
  assign n44258 = n44246 & n44257 ;
  assign n44259 = \m1_addr_i[22]_pad  & ~n13627 ;
  assign n44260 = n13620 & n44259 ;
  assign n44261 = \m2_addr_i[22]_pad  & n13627 ;
  assign n44262 = n13635 & n44261 ;
  assign n44263 = ~n44260 & ~n44262 ;
  assign n44264 = \m3_addr_i[22]_pad  & ~n13627 ;
  assign n44265 = n13635 & n44264 ;
  assign n44266 = \m5_addr_i[22]_pad  & ~n13627 ;
  assign n44267 = n13652 & n44266 ;
  assign n44268 = ~n44265 & ~n44267 ;
  assign n44269 = n44263 & n44268 ;
  assign n44270 = \m4_addr_i[22]_pad  & n13627 ;
  assign n44271 = n13652 & n44270 ;
  assign n44272 = \m6_addr_i[22]_pad  & n13627 ;
  assign n44273 = n13644 & n44272 ;
  assign n44274 = ~n44271 & ~n44273 ;
  assign n44275 = \m0_addr_i[22]_pad  & n13627 ;
  assign n44276 = n13620 & n44275 ;
  assign n44277 = \m7_addr_i[22]_pad  & ~n13627 ;
  assign n44278 = n13644 & n44277 ;
  assign n44279 = ~n44276 & ~n44278 ;
  assign n44280 = n44274 & n44279 ;
  assign n44281 = n44269 & n44280 ;
  assign n44282 = \m3_addr_i[23]_pad  & ~n13627 ;
  assign n44283 = n13635 & n44282 ;
  assign n44284 = \m4_addr_i[23]_pad  & n13627 ;
  assign n44285 = n13652 & n44284 ;
  assign n44286 = ~n44283 & ~n44285 ;
  assign n44287 = \m1_addr_i[23]_pad  & ~n13627 ;
  assign n44288 = n13620 & n44287 ;
  assign n44289 = \m5_addr_i[23]_pad  & ~n13627 ;
  assign n44290 = n13652 & n44289 ;
  assign n44291 = ~n44288 & ~n44290 ;
  assign n44292 = n44286 & n44291 ;
  assign n44293 = \m2_addr_i[23]_pad  & n13627 ;
  assign n44294 = n13635 & n44293 ;
  assign n44295 = \m6_addr_i[23]_pad  & n13627 ;
  assign n44296 = n13644 & n44295 ;
  assign n44297 = ~n44294 & ~n44296 ;
  assign n44298 = \m0_addr_i[23]_pad  & n13627 ;
  assign n44299 = n13620 & n44298 ;
  assign n44300 = \m7_addr_i[23]_pad  & ~n13627 ;
  assign n44301 = n13644 & n44300 ;
  assign n44302 = ~n44299 & ~n44301 ;
  assign n44303 = n44297 & n44302 ;
  assign n44304 = n44292 & n44303 ;
  assign n44305 = \m1_addr_i[24]_pad  & ~n13627 ;
  assign n44306 = n13620 & n44305 ;
  assign n44307 = \m2_addr_i[24]_pad  & n13627 ;
  assign n44308 = n13635 & n44307 ;
  assign n44309 = ~n44306 & ~n44308 ;
  assign n44310 = \m3_addr_i[24]_pad  & ~n13627 ;
  assign n44311 = n13635 & n44310 ;
  assign n44312 = \m7_addr_i[24]_pad  & ~n13627 ;
  assign n44313 = n13644 & n44312 ;
  assign n44314 = ~n44311 & ~n44313 ;
  assign n44315 = n44309 & n44314 ;
  assign n44316 = \m4_addr_i[24]_pad  & n13627 ;
  assign n44317 = n13652 & n44316 ;
  assign n44318 = \m0_addr_i[24]_pad  & n13627 ;
  assign n44319 = n13620 & n44318 ;
  assign n44320 = ~n44317 & ~n44319 ;
  assign n44321 = \m5_addr_i[24]_pad  & ~n13627 ;
  assign n44322 = n13652 & n44321 ;
  assign n44323 = \m6_addr_i[24]_pad  & n13627 ;
  assign n44324 = n13644 & n44323 ;
  assign n44325 = ~n44322 & ~n44324 ;
  assign n44326 = n44320 & n44325 ;
  assign n44327 = n44315 & n44326 ;
  assign n44328 = \m3_addr_i[25]_pad  & ~n13627 ;
  assign n44329 = n13635 & n44328 ;
  assign n44330 = \m4_addr_i[25]_pad  & n13627 ;
  assign n44331 = n13652 & n44330 ;
  assign n44332 = ~n44329 & ~n44331 ;
  assign n44333 = \m0_addr_i[25]_pad  & n13627 ;
  assign n44334 = n13620 & n44333 ;
  assign n44335 = \m2_addr_i[25]_pad  & n13627 ;
  assign n44336 = n13635 & n44335 ;
  assign n44337 = ~n44334 & ~n44336 ;
  assign n44338 = n44332 & n44337 ;
  assign n44339 = \m7_addr_i[25]_pad  & ~n13627 ;
  assign n44340 = n13644 & n44339 ;
  assign n44341 = \m1_addr_i[25]_pad  & ~n13627 ;
  assign n44342 = n13620 & n44341 ;
  assign n44343 = ~n44340 & ~n44342 ;
  assign n44344 = \m5_addr_i[25]_pad  & ~n13627 ;
  assign n44345 = n13652 & n44344 ;
  assign n44346 = \m6_addr_i[25]_pad  & n13627 ;
  assign n44347 = n13644 & n44346 ;
  assign n44348 = ~n44345 & ~n44347 ;
  assign n44349 = n44343 & n44348 ;
  assign n44350 = n44338 & n44349 ;
  assign n44351 = \m1_addr_i[26]_pad  & ~n13627 ;
  assign n44352 = n13620 & n44351 ;
  assign n44353 = \m2_addr_i[26]_pad  & n13627 ;
  assign n44354 = n13635 & n44353 ;
  assign n44355 = ~n44352 & ~n44354 ;
  assign n44356 = \m0_addr_i[26]_pad  & n13627 ;
  assign n44357 = n13620 & n44356 ;
  assign n44358 = \m4_addr_i[26]_pad  & n13627 ;
  assign n44359 = n13652 & n44358 ;
  assign n44360 = ~n44357 & ~n44359 ;
  assign n44361 = n44355 & n44360 ;
  assign n44362 = \m7_addr_i[26]_pad  & ~n13627 ;
  assign n44363 = n13644 & n44362 ;
  assign n44364 = \m3_addr_i[26]_pad  & ~n13627 ;
  assign n44365 = n13635 & n44364 ;
  assign n44366 = ~n44363 & ~n44365 ;
  assign n44367 = \m5_addr_i[26]_pad  & ~n13627 ;
  assign n44368 = n13652 & n44367 ;
  assign n44369 = \m6_addr_i[26]_pad  & n13627 ;
  assign n44370 = n13644 & n44369 ;
  assign n44371 = ~n44368 & ~n44370 ;
  assign n44372 = n44366 & n44371 ;
  assign n44373 = n44361 & n44372 ;
  assign n44374 = \m3_addr_i[27]_pad  & ~n13627 ;
  assign n44375 = n13635 & n44374 ;
  assign n44376 = \m4_addr_i[27]_pad  & n13627 ;
  assign n44377 = n13652 & n44376 ;
  assign n44378 = ~n44375 & ~n44377 ;
  assign n44379 = \m0_addr_i[27]_pad  & n13627 ;
  assign n44380 = n13620 & n44379 ;
  assign n44381 = \m6_addr_i[27]_pad  & n13627 ;
  assign n44382 = n13644 & n44381 ;
  assign n44383 = ~n44380 & ~n44382 ;
  assign n44384 = n44378 & n44383 ;
  assign n44385 = \m7_addr_i[27]_pad  & ~n13627 ;
  assign n44386 = n13644 & n44385 ;
  assign n44387 = \m5_addr_i[27]_pad  & ~n13627 ;
  assign n44388 = n13652 & n44387 ;
  assign n44389 = ~n44386 & ~n44388 ;
  assign n44390 = \m1_addr_i[27]_pad  & ~n13627 ;
  assign n44391 = n13620 & n44390 ;
  assign n44392 = \m2_addr_i[27]_pad  & n13627 ;
  assign n44393 = n13635 & n44392 ;
  assign n44394 = ~n44391 & ~n44393 ;
  assign n44395 = n44389 & n44394 ;
  assign n44396 = n44384 & n44395 ;
  assign n44397 = \m1_addr_i[28]_pad  & ~n13627 ;
  assign n44398 = n13620 & n44397 ;
  assign n44399 = \m2_addr_i[28]_pad  & n13627 ;
  assign n44400 = n13635 & n44399 ;
  assign n44401 = ~n44398 & ~n44400 ;
  assign n44402 = \m0_addr_i[28]_pad  & n13627 ;
  assign n44403 = n13620 & n44402 ;
  assign n44404 = \m6_addr_i[28]_pad  & n13627 ;
  assign n44405 = n13644 & n44404 ;
  assign n44406 = ~n44403 & ~n44405 ;
  assign n44407 = n44401 & n44406 ;
  assign n44408 = \m7_addr_i[28]_pad  & ~n13627 ;
  assign n44409 = n13644 & n44408 ;
  assign n44410 = \m5_addr_i[28]_pad  & ~n13627 ;
  assign n44411 = n13652 & n44410 ;
  assign n44412 = ~n44409 & ~n44411 ;
  assign n44413 = \m3_addr_i[28]_pad  & ~n13627 ;
  assign n44414 = n13635 & n44413 ;
  assign n44415 = \m4_addr_i[28]_pad  & n13627 ;
  assign n44416 = n13652 & n44415 ;
  assign n44417 = ~n44414 & ~n44416 ;
  assign n44418 = n44412 & n44417 ;
  assign n44419 = n44407 & n44418 ;
  assign n44420 = \m0_addr_i[29]_pad  & n13627 ;
  assign n44421 = n13620 & n44420 ;
  assign n44422 = \m7_addr_i[29]_pad  & ~n13627 ;
  assign n44423 = n13644 & n44422 ;
  assign n44424 = ~n44421 & ~n44423 ;
  assign n44425 = \m5_addr_i[29]_pad  & ~n13627 ;
  assign n44426 = n13652 & n44425 ;
  assign n44427 = \m2_addr_i[29]_pad  & n13627 ;
  assign n44428 = n13635 & n44427 ;
  assign n44429 = ~n44426 & ~n44428 ;
  assign n44430 = n44424 & n44429 ;
  assign n44431 = \m6_addr_i[29]_pad  & n13627 ;
  assign n44432 = n13644 & n44431 ;
  assign n44433 = \m1_addr_i[29]_pad  & ~n13627 ;
  assign n44434 = n13620 & n44433 ;
  assign n44435 = ~n44432 & ~n44434 ;
  assign n44436 = \m3_addr_i[29]_pad  & ~n13627 ;
  assign n44437 = n13635 & n44436 ;
  assign n44438 = \m4_addr_i[29]_pad  & n13627 ;
  assign n44439 = n13652 & n44438 ;
  assign n44440 = ~n44437 & ~n44439 ;
  assign n44441 = n44435 & n44440 ;
  assign n44442 = n44430 & n44441 ;
  assign n44443 = \m3_addr_i[2]_pad  & ~n13627 ;
  assign n44444 = n13635 & n44443 ;
  assign n44445 = \m4_addr_i[2]_pad  & n13627 ;
  assign n44446 = n13652 & n44445 ;
  assign n44447 = ~n44444 & ~n44446 ;
  assign n44448 = \m6_addr_i[2]_pad  & n13627 ;
  assign n44449 = n13644 & n44448 ;
  assign n44450 = \m2_addr_i[2]_pad  & n13627 ;
  assign n44451 = n13635 & n44450 ;
  assign n44452 = ~n44449 & ~n44451 ;
  assign n44453 = n44447 & n44452 ;
  assign n44454 = \m5_addr_i[2]_pad  & ~n13627 ;
  assign n44455 = n13652 & n44454 ;
  assign n44456 = \m1_addr_i[2]_pad  & ~n13627 ;
  assign n44457 = n13620 & n44456 ;
  assign n44458 = ~n44455 & ~n44457 ;
  assign n44459 = \m0_addr_i[2]_pad  & n13627 ;
  assign n44460 = n13620 & n44459 ;
  assign n44461 = \m7_addr_i[2]_pad  & ~n13627 ;
  assign n44462 = n13644 & n44461 ;
  assign n44463 = ~n44460 & ~n44462 ;
  assign n44464 = n44458 & n44463 ;
  assign n44465 = n44453 & n44464 ;
  assign n44466 = \m1_addr_i[30]_pad  & ~n13627 ;
  assign n44467 = n13620 & n44466 ;
  assign n44468 = \m2_addr_i[30]_pad  & n13627 ;
  assign n44469 = n13635 & n44468 ;
  assign n44470 = ~n44467 & ~n44469 ;
  assign n44471 = \m0_addr_i[30]_pad  & n13627 ;
  assign n44472 = n13620 & n44471 ;
  assign n44473 = \m4_addr_i[30]_pad  & n13627 ;
  assign n44474 = n13652 & n44473 ;
  assign n44475 = ~n44472 & ~n44474 ;
  assign n44476 = n44470 & n44475 ;
  assign n44477 = \m7_addr_i[30]_pad  & ~n13627 ;
  assign n44478 = n13644 & n44477 ;
  assign n44479 = \m3_addr_i[30]_pad  & ~n13627 ;
  assign n44480 = n13635 & n44479 ;
  assign n44481 = ~n44478 & ~n44480 ;
  assign n44482 = \m5_addr_i[30]_pad  & ~n13627 ;
  assign n44483 = n13652 & n44482 ;
  assign n44484 = \m6_addr_i[30]_pad  & n13627 ;
  assign n44485 = n13644 & n44484 ;
  assign n44486 = ~n44483 & ~n44485 ;
  assign n44487 = n44481 & n44486 ;
  assign n44488 = n44476 & n44487 ;
  assign n44489 = \m0_addr_i[31]_pad  & n13627 ;
  assign n44490 = n13620 & n44489 ;
  assign n44491 = \m7_addr_i[31]_pad  & ~n13627 ;
  assign n44492 = n13644 & n44491 ;
  assign n44493 = ~n44490 & ~n44492 ;
  assign n44494 = \m3_addr_i[31]_pad  & ~n13627 ;
  assign n44495 = n13635 & n44494 ;
  assign n44496 = \m2_addr_i[31]_pad  & n13627 ;
  assign n44497 = n13635 & n44496 ;
  assign n44498 = ~n44495 & ~n44497 ;
  assign n44499 = n44493 & n44498 ;
  assign n44500 = \m4_addr_i[31]_pad  & n13627 ;
  assign n44501 = n13652 & n44500 ;
  assign n44502 = \m1_addr_i[31]_pad  & ~n13627 ;
  assign n44503 = n13620 & n44502 ;
  assign n44504 = ~n44501 & ~n44503 ;
  assign n44505 = \m5_addr_i[31]_pad  & ~n13627 ;
  assign n44506 = n13652 & n44505 ;
  assign n44507 = \m6_addr_i[31]_pad  & n13627 ;
  assign n44508 = n13644 & n44507 ;
  assign n44509 = ~n44506 & ~n44508 ;
  assign n44510 = n44504 & n44509 ;
  assign n44511 = n44499 & n44510 ;
  assign n44512 = \m3_addr_i[3]_pad  & ~n13627 ;
  assign n44513 = n13635 & n44512 ;
  assign n44514 = \m4_addr_i[3]_pad  & n13627 ;
  assign n44515 = n13652 & n44514 ;
  assign n44516 = ~n44513 & ~n44515 ;
  assign n44517 = \m6_addr_i[3]_pad  & n13627 ;
  assign n44518 = n13644 & n44517 ;
  assign n44519 = \m2_addr_i[3]_pad  & n13627 ;
  assign n44520 = n13635 & n44519 ;
  assign n44521 = ~n44518 & ~n44520 ;
  assign n44522 = n44516 & n44521 ;
  assign n44523 = \m5_addr_i[3]_pad  & ~n13627 ;
  assign n44524 = n13652 & n44523 ;
  assign n44525 = \m1_addr_i[3]_pad  & ~n13627 ;
  assign n44526 = n13620 & n44525 ;
  assign n44527 = ~n44524 & ~n44526 ;
  assign n44528 = \m0_addr_i[3]_pad  & n13627 ;
  assign n44529 = n13620 & n44528 ;
  assign n44530 = \m7_addr_i[3]_pad  & ~n13627 ;
  assign n44531 = n13644 & n44530 ;
  assign n44532 = ~n44529 & ~n44531 ;
  assign n44533 = n44527 & n44532 ;
  assign n44534 = n44522 & n44533 ;
  assign n44535 = \m3_addr_i[4]_pad  & ~n13627 ;
  assign n44536 = n13635 & n44535 ;
  assign n44537 = \m4_addr_i[4]_pad  & n13627 ;
  assign n44538 = n13652 & n44537 ;
  assign n44539 = ~n44536 & ~n44538 ;
  assign n44540 = \m6_addr_i[4]_pad  & n13627 ;
  assign n44541 = n13644 & n44540 ;
  assign n44542 = \m2_addr_i[4]_pad  & n13627 ;
  assign n44543 = n13635 & n44542 ;
  assign n44544 = ~n44541 & ~n44543 ;
  assign n44545 = n44539 & n44544 ;
  assign n44546 = \m5_addr_i[4]_pad  & ~n13627 ;
  assign n44547 = n13652 & n44546 ;
  assign n44548 = \m1_addr_i[4]_pad  & ~n13627 ;
  assign n44549 = n13620 & n44548 ;
  assign n44550 = ~n44547 & ~n44549 ;
  assign n44551 = \m0_addr_i[4]_pad  & n13627 ;
  assign n44552 = n13620 & n44551 ;
  assign n44553 = \m7_addr_i[4]_pad  & ~n13627 ;
  assign n44554 = n13644 & n44553 ;
  assign n44555 = ~n44552 & ~n44554 ;
  assign n44556 = n44550 & n44555 ;
  assign n44557 = n44545 & n44556 ;
  assign n44558 = \m3_addr_i[5]_pad  & ~n13627 ;
  assign n44559 = n13635 & n44558 ;
  assign n44560 = \m4_addr_i[5]_pad  & n13627 ;
  assign n44561 = n13652 & n44560 ;
  assign n44562 = ~n44559 & ~n44561 ;
  assign n44563 = \m6_addr_i[5]_pad  & n13627 ;
  assign n44564 = n13644 & n44563 ;
  assign n44565 = \m2_addr_i[5]_pad  & n13627 ;
  assign n44566 = n13635 & n44565 ;
  assign n44567 = ~n44564 & ~n44566 ;
  assign n44568 = n44562 & n44567 ;
  assign n44569 = \m5_addr_i[5]_pad  & ~n13627 ;
  assign n44570 = n13652 & n44569 ;
  assign n44571 = \m1_addr_i[5]_pad  & ~n13627 ;
  assign n44572 = n13620 & n44571 ;
  assign n44573 = ~n44570 & ~n44572 ;
  assign n44574 = \m0_addr_i[5]_pad  & n13627 ;
  assign n44575 = n13620 & n44574 ;
  assign n44576 = \m7_addr_i[5]_pad  & ~n13627 ;
  assign n44577 = n13644 & n44576 ;
  assign n44578 = ~n44575 & ~n44577 ;
  assign n44579 = n44573 & n44578 ;
  assign n44580 = n44568 & n44579 ;
  assign n44581 = \m3_addr_i[6]_pad  & ~n13627 ;
  assign n44582 = n13635 & n44581 ;
  assign n44583 = \m4_addr_i[6]_pad  & n13627 ;
  assign n44584 = n13652 & n44583 ;
  assign n44585 = ~n44582 & ~n44584 ;
  assign n44586 = \m6_addr_i[6]_pad  & n13627 ;
  assign n44587 = n13644 & n44586 ;
  assign n44588 = \m2_addr_i[6]_pad  & n13627 ;
  assign n44589 = n13635 & n44588 ;
  assign n44590 = ~n44587 & ~n44589 ;
  assign n44591 = n44585 & n44590 ;
  assign n44592 = \m5_addr_i[6]_pad  & ~n13627 ;
  assign n44593 = n13652 & n44592 ;
  assign n44594 = \m1_addr_i[6]_pad  & ~n13627 ;
  assign n44595 = n13620 & n44594 ;
  assign n44596 = ~n44593 & ~n44595 ;
  assign n44597 = \m0_addr_i[6]_pad  & n13627 ;
  assign n44598 = n13620 & n44597 ;
  assign n44599 = \m7_addr_i[6]_pad  & ~n13627 ;
  assign n44600 = n13644 & n44599 ;
  assign n44601 = ~n44598 & ~n44600 ;
  assign n44602 = n44596 & n44601 ;
  assign n44603 = n44591 & n44602 ;
  assign n44604 = \m3_addr_i[7]_pad  & ~n13627 ;
  assign n44605 = n13635 & n44604 ;
  assign n44606 = \m4_addr_i[7]_pad  & n13627 ;
  assign n44607 = n13652 & n44606 ;
  assign n44608 = ~n44605 & ~n44607 ;
  assign n44609 = \m6_addr_i[7]_pad  & n13627 ;
  assign n44610 = n13644 & n44609 ;
  assign n44611 = \m2_addr_i[7]_pad  & n13627 ;
  assign n44612 = n13635 & n44611 ;
  assign n44613 = ~n44610 & ~n44612 ;
  assign n44614 = n44608 & n44613 ;
  assign n44615 = \m5_addr_i[7]_pad  & ~n13627 ;
  assign n44616 = n13652 & n44615 ;
  assign n44617 = \m1_addr_i[7]_pad  & ~n13627 ;
  assign n44618 = n13620 & n44617 ;
  assign n44619 = ~n44616 & ~n44618 ;
  assign n44620 = \m0_addr_i[7]_pad  & n13627 ;
  assign n44621 = n13620 & n44620 ;
  assign n44622 = \m7_addr_i[7]_pad  & ~n13627 ;
  assign n44623 = n13644 & n44622 ;
  assign n44624 = ~n44621 & ~n44623 ;
  assign n44625 = n44619 & n44624 ;
  assign n44626 = n44614 & n44625 ;
  assign n44627 = \m3_addr_i[8]_pad  & ~n13627 ;
  assign n44628 = n13635 & n44627 ;
  assign n44629 = \m4_addr_i[8]_pad  & n13627 ;
  assign n44630 = n13652 & n44629 ;
  assign n44631 = ~n44628 & ~n44630 ;
  assign n44632 = \m6_addr_i[8]_pad  & n13627 ;
  assign n44633 = n13644 & n44632 ;
  assign n44634 = \m2_addr_i[8]_pad  & n13627 ;
  assign n44635 = n13635 & n44634 ;
  assign n44636 = ~n44633 & ~n44635 ;
  assign n44637 = n44631 & n44636 ;
  assign n44638 = \m5_addr_i[8]_pad  & ~n13627 ;
  assign n44639 = n13652 & n44638 ;
  assign n44640 = \m1_addr_i[8]_pad  & ~n13627 ;
  assign n44641 = n13620 & n44640 ;
  assign n44642 = ~n44639 & ~n44641 ;
  assign n44643 = \m0_addr_i[8]_pad  & n13627 ;
  assign n44644 = n13620 & n44643 ;
  assign n44645 = \m7_addr_i[8]_pad  & ~n13627 ;
  assign n44646 = n13644 & n44645 ;
  assign n44647 = ~n44644 & ~n44646 ;
  assign n44648 = n44642 & n44647 ;
  assign n44649 = n44637 & n44648 ;
  assign n44650 = \m3_addr_i[9]_pad  & ~n13627 ;
  assign n44651 = n13635 & n44650 ;
  assign n44652 = \m4_addr_i[9]_pad  & n13627 ;
  assign n44653 = n13652 & n44652 ;
  assign n44654 = ~n44651 & ~n44653 ;
  assign n44655 = \m6_addr_i[9]_pad  & n13627 ;
  assign n44656 = n13644 & n44655 ;
  assign n44657 = \m2_addr_i[9]_pad  & n13627 ;
  assign n44658 = n13635 & n44657 ;
  assign n44659 = ~n44656 & ~n44658 ;
  assign n44660 = n44654 & n44659 ;
  assign n44661 = \m5_addr_i[9]_pad  & ~n13627 ;
  assign n44662 = n13652 & n44661 ;
  assign n44663 = \m1_addr_i[9]_pad  & ~n13627 ;
  assign n44664 = n13620 & n44663 ;
  assign n44665 = ~n44662 & ~n44664 ;
  assign n44666 = \m0_addr_i[9]_pad  & n13627 ;
  assign n44667 = n13620 & n44666 ;
  assign n44668 = \m7_addr_i[9]_pad  & ~n13627 ;
  assign n44669 = n13644 & n44668 ;
  assign n44670 = ~n44667 & ~n44669 ;
  assign n44671 = n44665 & n44670 ;
  assign n44672 = n44660 & n44671 ;
  assign n44673 = \m0_data_i[0]_pad  & n13627 ;
  assign n44674 = n13620 & n44673 ;
  assign n44675 = \m7_data_i[0]_pad  & ~n13627 ;
  assign n44676 = n13644 & n44675 ;
  assign n44677 = ~n44674 & ~n44676 ;
  assign n44678 = \m6_data_i[0]_pad  & n13627 ;
  assign n44679 = n13644 & n44678 ;
  assign n44680 = \m2_data_i[0]_pad  & n13627 ;
  assign n44681 = n13635 & n44680 ;
  assign n44682 = ~n44679 & ~n44681 ;
  assign n44683 = n44677 & n44682 ;
  assign n44684 = \m5_data_i[0]_pad  & ~n13627 ;
  assign n44685 = n13652 & n44684 ;
  assign n44686 = \m1_data_i[0]_pad  & ~n13627 ;
  assign n44687 = n13620 & n44686 ;
  assign n44688 = ~n44685 & ~n44687 ;
  assign n44689 = \m3_data_i[0]_pad  & ~n13627 ;
  assign n44690 = n13635 & n44689 ;
  assign n44691 = \m4_data_i[0]_pad  & n13627 ;
  assign n44692 = n13652 & n44691 ;
  assign n44693 = ~n44690 & ~n44692 ;
  assign n44694 = n44688 & n44693 ;
  assign n44695 = n44683 & n44694 ;
  assign n44696 = \m0_data_i[10]_pad  & n13627 ;
  assign n44697 = n13620 & n44696 ;
  assign n44698 = \m7_data_i[10]_pad  & ~n13627 ;
  assign n44699 = n13644 & n44698 ;
  assign n44700 = ~n44697 & ~n44699 ;
  assign n44701 = \m6_data_i[10]_pad  & n13627 ;
  assign n44702 = n13644 & n44701 ;
  assign n44703 = \m2_data_i[10]_pad  & n13627 ;
  assign n44704 = n13635 & n44703 ;
  assign n44705 = ~n44702 & ~n44704 ;
  assign n44706 = n44700 & n44705 ;
  assign n44707 = \m5_data_i[10]_pad  & ~n13627 ;
  assign n44708 = n13652 & n44707 ;
  assign n44709 = \m1_data_i[10]_pad  & ~n13627 ;
  assign n44710 = n13620 & n44709 ;
  assign n44711 = ~n44708 & ~n44710 ;
  assign n44712 = \m3_data_i[10]_pad  & ~n13627 ;
  assign n44713 = n13635 & n44712 ;
  assign n44714 = \m4_data_i[10]_pad  & n13627 ;
  assign n44715 = n13652 & n44714 ;
  assign n44716 = ~n44713 & ~n44715 ;
  assign n44717 = n44711 & n44716 ;
  assign n44718 = n44706 & n44717 ;
  assign n44719 = \m3_data_i[11]_pad  & ~n13627 ;
  assign n44720 = n13635 & n44719 ;
  assign n44721 = \m4_data_i[11]_pad  & n13627 ;
  assign n44722 = n13652 & n44721 ;
  assign n44723 = ~n44720 & ~n44722 ;
  assign n44724 = \m6_data_i[11]_pad  & n13627 ;
  assign n44725 = n13644 & n44724 ;
  assign n44726 = \m7_data_i[11]_pad  & ~n13627 ;
  assign n44727 = n13644 & n44726 ;
  assign n44728 = ~n44725 & ~n44727 ;
  assign n44729 = n44723 & n44728 ;
  assign n44730 = \m5_data_i[11]_pad  & ~n13627 ;
  assign n44731 = n13652 & n44730 ;
  assign n44732 = \m0_data_i[11]_pad  & n13627 ;
  assign n44733 = n13620 & n44732 ;
  assign n44734 = ~n44731 & ~n44733 ;
  assign n44735 = \m1_data_i[11]_pad  & ~n13627 ;
  assign n44736 = n13620 & n44735 ;
  assign n44737 = \m2_data_i[11]_pad  & n13627 ;
  assign n44738 = n13635 & n44737 ;
  assign n44739 = ~n44736 & ~n44738 ;
  assign n44740 = n44734 & n44739 ;
  assign n44741 = n44729 & n44740 ;
  assign n44742 = \m3_data_i[12]_pad  & ~n13627 ;
  assign n44743 = n13635 & n44742 ;
  assign n44744 = \m4_data_i[12]_pad  & n13627 ;
  assign n44745 = n13652 & n44744 ;
  assign n44746 = ~n44743 & ~n44745 ;
  assign n44747 = \m6_data_i[12]_pad  & n13627 ;
  assign n44748 = n13644 & n44747 ;
  assign n44749 = \m2_data_i[12]_pad  & n13627 ;
  assign n44750 = n13635 & n44749 ;
  assign n44751 = ~n44748 & ~n44750 ;
  assign n44752 = n44746 & n44751 ;
  assign n44753 = \m5_data_i[12]_pad  & ~n13627 ;
  assign n44754 = n13652 & n44753 ;
  assign n44755 = \m1_data_i[12]_pad  & ~n13627 ;
  assign n44756 = n13620 & n44755 ;
  assign n44757 = ~n44754 & ~n44756 ;
  assign n44758 = \m0_data_i[12]_pad  & n13627 ;
  assign n44759 = n13620 & n44758 ;
  assign n44760 = \m7_data_i[12]_pad  & ~n13627 ;
  assign n44761 = n13644 & n44760 ;
  assign n44762 = ~n44759 & ~n44761 ;
  assign n44763 = n44757 & n44762 ;
  assign n44764 = n44752 & n44763 ;
  assign n44765 = \m0_data_i[13]_pad  & n13627 ;
  assign n44766 = n13620 & n44765 ;
  assign n44767 = \m7_data_i[13]_pad  & ~n13627 ;
  assign n44768 = n13644 & n44767 ;
  assign n44769 = ~n44766 & ~n44768 ;
  assign n44770 = \m6_data_i[13]_pad  & n13627 ;
  assign n44771 = n13644 & n44770 ;
  assign n44772 = \m2_data_i[13]_pad  & n13627 ;
  assign n44773 = n13635 & n44772 ;
  assign n44774 = ~n44771 & ~n44773 ;
  assign n44775 = n44769 & n44774 ;
  assign n44776 = \m5_data_i[13]_pad  & ~n13627 ;
  assign n44777 = n13652 & n44776 ;
  assign n44778 = \m1_data_i[13]_pad  & ~n13627 ;
  assign n44779 = n13620 & n44778 ;
  assign n44780 = ~n44777 & ~n44779 ;
  assign n44781 = \m3_data_i[13]_pad  & ~n13627 ;
  assign n44782 = n13635 & n44781 ;
  assign n44783 = \m4_data_i[13]_pad  & n13627 ;
  assign n44784 = n13652 & n44783 ;
  assign n44785 = ~n44782 & ~n44784 ;
  assign n44786 = n44780 & n44785 ;
  assign n44787 = n44775 & n44786 ;
  assign n44788 = \m0_data_i[14]_pad  & n13627 ;
  assign n44789 = n13620 & n44788 ;
  assign n44790 = \m7_data_i[14]_pad  & ~n13627 ;
  assign n44791 = n13644 & n44790 ;
  assign n44792 = ~n44789 & ~n44791 ;
  assign n44793 = \m6_data_i[14]_pad  & n13627 ;
  assign n44794 = n13644 & n44793 ;
  assign n44795 = \m2_data_i[14]_pad  & n13627 ;
  assign n44796 = n13635 & n44795 ;
  assign n44797 = ~n44794 & ~n44796 ;
  assign n44798 = n44792 & n44797 ;
  assign n44799 = \m5_data_i[14]_pad  & ~n13627 ;
  assign n44800 = n13652 & n44799 ;
  assign n44801 = \m1_data_i[14]_pad  & ~n13627 ;
  assign n44802 = n13620 & n44801 ;
  assign n44803 = ~n44800 & ~n44802 ;
  assign n44804 = \m3_data_i[14]_pad  & ~n13627 ;
  assign n44805 = n13635 & n44804 ;
  assign n44806 = \m4_data_i[14]_pad  & n13627 ;
  assign n44807 = n13652 & n44806 ;
  assign n44808 = ~n44805 & ~n44807 ;
  assign n44809 = n44803 & n44808 ;
  assign n44810 = n44798 & n44809 ;
  assign n44811 = \m3_data_i[15]_pad  & ~n13627 ;
  assign n44812 = n13635 & n44811 ;
  assign n44813 = \m4_data_i[15]_pad  & n13627 ;
  assign n44814 = n13652 & n44813 ;
  assign n44815 = ~n44812 & ~n44814 ;
  assign n44816 = \m6_data_i[15]_pad  & n13627 ;
  assign n44817 = n13644 & n44816 ;
  assign n44818 = \m2_data_i[15]_pad  & n13627 ;
  assign n44819 = n13635 & n44818 ;
  assign n44820 = ~n44817 & ~n44819 ;
  assign n44821 = n44815 & n44820 ;
  assign n44822 = \m5_data_i[15]_pad  & ~n13627 ;
  assign n44823 = n13652 & n44822 ;
  assign n44824 = \m1_data_i[15]_pad  & ~n13627 ;
  assign n44825 = n13620 & n44824 ;
  assign n44826 = ~n44823 & ~n44825 ;
  assign n44827 = \m0_data_i[15]_pad  & n13627 ;
  assign n44828 = n13620 & n44827 ;
  assign n44829 = \m7_data_i[15]_pad  & ~n13627 ;
  assign n44830 = n13644 & n44829 ;
  assign n44831 = ~n44828 & ~n44830 ;
  assign n44832 = n44826 & n44831 ;
  assign n44833 = n44821 & n44832 ;
  assign n44834 = \m3_data_i[16]_pad  & ~n13627 ;
  assign n44835 = n13635 & n44834 ;
  assign n44836 = \m4_data_i[16]_pad  & n13627 ;
  assign n44837 = n13652 & n44836 ;
  assign n44838 = ~n44835 & ~n44837 ;
  assign n44839 = \m6_data_i[16]_pad  & n13627 ;
  assign n44840 = n13644 & n44839 ;
  assign n44841 = \m2_data_i[16]_pad  & n13627 ;
  assign n44842 = n13635 & n44841 ;
  assign n44843 = ~n44840 & ~n44842 ;
  assign n44844 = n44838 & n44843 ;
  assign n44845 = \m5_data_i[16]_pad  & ~n13627 ;
  assign n44846 = n13652 & n44845 ;
  assign n44847 = \m1_data_i[16]_pad  & ~n13627 ;
  assign n44848 = n13620 & n44847 ;
  assign n44849 = ~n44846 & ~n44848 ;
  assign n44850 = \m0_data_i[16]_pad  & n13627 ;
  assign n44851 = n13620 & n44850 ;
  assign n44852 = \m7_data_i[16]_pad  & ~n13627 ;
  assign n44853 = n13644 & n44852 ;
  assign n44854 = ~n44851 & ~n44853 ;
  assign n44855 = n44849 & n44854 ;
  assign n44856 = n44844 & n44855 ;
  assign n44857 = \m3_data_i[17]_pad  & ~n13627 ;
  assign n44858 = n13635 & n44857 ;
  assign n44859 = \m4_data_i[17]_pad  & n13627 ;
  assign n44860 = n13652 & n44859 ;
  assign n44861 = ~n44858 & ~n44860 ;
  assign n44862 = \m6_data_i[17]_pad  & n13627 ;
  assign n44863 = n13644 & n44862 ;
  assign n44864 = \m2_data_i[17]_pad  & n13627 ;
  assign n44865 = n13635 & n44864 ;
  assign n44866 = ~n44863 & ~n44865 ;
  assign n44867 = n44861 & n44866 ;
  assign n44868 = \m5_data_i[17]_pad  & ~n13627 ;
  assign n44869 = n13652 & n44868 ;
  assign n44870 = \m1_data_i[17]_pad  & ~n13627 ;
  assign n44871 = n13620 & n44870 ;
  assign n44872 = ~n44869 & ~n44871 ;
  assign n44873 = \m0_data_i[17]_pad  & n13627 ;
  assign n44874 = n13620 & n44873 ;
  assign n44875 = \m7_data_i[17]_pad  & ~n13627 ;
  assign n44876 = n13644 & n44875 ;
  assign n44877 = ~n44874 & ~n44876 ;
  assign n44878 = n44872 & n44877 ;
  assign n44879 = n44867 & n44878 ;
  assign n44880 = \m1_data_i[18]_pad  & ~n13627 ;
  assign n44881 = n13620 & n44880 ;
  assign n44882 = \m2_data_i[18]_pad  & n13627 ;
  assign n44883 = n13635 & n44882 ;
  assign n44884 = ~n44881 & ~n44883 ;
  assign n44885 = \m6_data_i[18]_pad  & n13627 ;
  assign n44886 = n13644 & n44885 ;
  assign n44887 = \m7_data_i[18]_pad  & ~n13627 ;
  assign n44888 = n13644 & n44887 ;
  assign n44889 = ~n44886 & ~n44888 ;
  assign n44890 = n44884 & n44889 ;
  assign n44891 = \m5_data_i[18]_pad  & ~n13627 ;
  assign n44892 = n13652 & n44891 ;
  assign n44893 = \m0_data_i[18]_pad  & n13627 ;
  assign n44894 = n13620 & n44893 ;
  assign n44895 = ~n44892 & ~n44894 ;
  assign n44896 = \m3_data_i[18]_pad  & ~n13627 ;
  assign n44897 = n13635 & n44896 ;
  assign n44898 = \m4_data_i[18]_pad  & n13627 ;
  assign n44899 = n13652 & n44898 ;
  assign n44900 = ~n44897 & ~n44899 ;
  assign n44901 = n44895 & n44900 ;
  assign n44902 = n44890 & n44901 ;
  assign n44903 = \m3_data_i[19]_pad  & ~n13627 ;
  assign n44904 = n13635 & n44903 ;
  assign n44905 = \m4_data_i[19]_pad  & n13627 ;
  assign n44906 = n13652 & n44905 ;
  assign n44907 = ~n44904 & ~n44906 ;
  assign n44908 = \m6_data_i[19]_pad  & n13627 ;
  assign n44909 = n13644 & n44908 ;
  assign n44910 = \m2_data_i[19]_pad  & n13627 ;
  assign n44911 = n13635 & n44910 ;
  assign n44912 = ~n44909 & ~n44911 ;
  assign n44913 = n44907 & n44912 ;
  assign n44914 = \m5_data_i[19]_pad  & ~n13627 ;
  assign n44915 = n13652 & n44914 ;
  assign n44916 = \m1_data_i[19]_pad  & ~n13627 ;
  assign n44917 = n13620 & n44916 ;
  assign n44918 = ~n44915 & ~n44917 ;
  assign n44919 = \m0_data_i[19]_pad  & n13627 ;
  assign n44920 = n13620 & n44919 ;
  assign n44921 = \m7_data_i[19]_pad  & ~n13627 ;
  assign n44922 = n13644 & n44921 ;
  assign n44923 = ~n44920 & ~n44922 ;
  assign n44924 = n44918 & n44923 ;
  assign n44925 = n44913 & n44924 ;
  assign n44926 = \m1_data_i[1]_pad  & ~n13627 ;
  assign n44927 = n13620 & n44926 ;
  assign n44928 = \m2_data_i[1]_pad  & n13627 ;
  assign n44929 = n13635 & n44928 ;
  assign n44930 = ~n44927 & ~n44929 ;
  assign n44931 = \m0_data_i[1]_pad  & n13627 ;
  assign n44932 = n13620 & n44931 ;
  assign n44933 = \m4_data_i[1]_pad  & n13627 ;
  assign n44934 = n13652 & n44933 ;
  assign n44935 = ~n44932 & ~n44934 ;
  assign n44936 = n44930 & n44935 ;
  assign n44937 = \m7_data_i[1]_pad  & ~n13627 ;
  assign n44938 = n13644 & n44937 ;
  assign n44939 = \m3_data_i[1]_pad  & ~n13627 ;
  assign n44940 = n13635 & n44939 ;
  assign n44941 = ~n44938 & ~n44940 ;
  assign n44942 = \m6_data_i[1]_pad  & n13627 ;
  assign n44943 = n13644 & n44942 ;
  assign n44944 = \m5_data_i[1]_pad  & ~n13627 ;
  assign n44945 = n13652 & n44944 ;
  assign n44946 = ~n44943 & ~n44945 ;
  assign n44947 = n44941 & n44946 ;
  assign n44948 = n44936 & n44947 ;
  assign n44949 = \m3_data_i[20]_pad  & ~n13627 ;
  assign n44950 = n13635 & n44949 ;
  assign n44951 = \m4_data_i[20]_pad  & n13627 ;
  assign n44952 = n13652 & n44951 ;
  assign n44953 = ~n44950 & ~n44952 ;
  assign n44954 = \m6_data_i[20]_pad  & n13627 ;
  assign n44955 = n13644 & n44954 ;
  assign n44956 = \m2_data_i[20]_pad  & n13627 ;
  assign n44957 = n13635 & n44956 ;
  assign n44958 = ~n44955 & ~n44957 ;
  assign n44959 = n44953 & n44958 ;
  assign n44960 = \m5_data_i[20]_pad  & ~n13627 ;
  assign n44961 = n13652 & n44960 ;
  assign n44962 = \m1_data_i[20]_pad  & ~n13627 ;
  assign n44963 = n13620 & n44962 ;
  assign n44964 = ~n44961 & ~n44963 ;
  assign n44965 = \m0_data_i[20]_pad  & n13627 ;
  assign n44966 = n13620 & n44965 ;
  assign n44967 = \m7_data_i[20]_pad  & ~n13627 ;
  assign n44968 = n13644 & n44967 ;
  assign n44969 = ~n44966 & ~n44968 ;
  assign n44970 = n44964 & n44969 ;
  assign n44971 = n44959 & n44970 ;
  assign n44972 = \m3_data_i[21]_pad  & ~n13627 ;
  assign n44973 = n13635 & n44972 ;
  assign n44974 = \m4_data_i[21]_pad  & n13627 ;
  assign n44975 = n13652 & n44974 ;
  assign n44976 = ~n44973 & ~n44975 ;
  assign n44977 = \m6_data_i[21]_pad  & n13627 ;
  assign n44978 = n13644 & n44977 ;
  assign n44979 = \m2_data_i[21]_pad  & n13627 ;
  assign n44980 = n13635 & n44979 ;
  assign n44981 = ~n44978 & ~n44980 ;
  assign n44982 = n44976 & n44981 ;
  assign n44983 = \m5_data_i[21]_pad  & ~n13627 ;
  assign n44984 = n13652 & n44983 ;
  assign n44985 = \m1_data_i[21]_pad  & ~n13627 ;
  assign n44986 = n13620 & n44985 ;
  assign n44987 = ~n44984 & ~n44986 ;
  assign n44988 = \m0_data_i[21]_pad  & n13627 ;
  assign n44989 = n13620 & n44988 ;
  assign n44990 = \m7_data_i[21]_pad  & ~n13627 ;
  assign n44991 = n13644 & n44990 ;
  assign n44992 = ~n44989 & ~n44991 ;
  assign n44993 = n44987 & n44992 ;
  assign n44994 = n44982 & n44993 ;
  assign n44995 = \m3_data_i[22]_pad  & ~n13627 ;
  assign n44996 = n13635 & n44995 ;
  assign n44997 = \m4_data_i[22]_pad  & n13627 ;
  assign n44998 = n13652 & n44997 ;
  assign n44999 = ~n44996 & ~n44998 ;
  assign n45000 = \m6_data_i[22]_pad  & n13627 ;
  assign n45001 = n13644 & n45000 ;
  assign n45002 = \m2_data_i[22]_pad  & n13627 ;
  assign n45003 = n13635 & n45002 ;
  assign n45004 = ~n45001 & ~n45003 ;
  assign n45005 = n44999 & n45004 ;
  assign n45006 = \m5_data_i[22]_pad  & ~n13627 ;
  assign n45007 = n13652 & n45006 ;
  assign n45008 = \m1_data_i[22]_pad  & ~n13627 ;
  assign n45009 = n13620 & n45008 ;
  assign n45010 = ~n45007 & ~n45009 ;
  assign n45011 = \m0_data_i[22]_pad  & n13627 ;
  assign n45012 = n13620 & n45011 ;
  assign n45013 = \m7_data_i[22]_pad  & ~n13627 ;
  assign n45014 = n13644 & n45013 ;
  assign n45015 = ~n45012 & ~n45014 ;
  assign n45016 = n45010 & n45015 ;
  assign n45017 = n45005 & n45016 ;
  assign n45018 = \m0_data_i[23]_pad  & n13627 ;
  assign n45019 = n13620 & n45018 ;
  assign n45020 = \m7_data_i[23]_pad  & ~n13627 ;
  assign n45021 = n13644 & n45020 ;
  assign n45022 = ~n45019 & ~n45021 ;
  assign n45023 = \m3_data_i[23]_pad  & ~n13627 ;
  assign n45024 = n13635 & n45023 ;
  assign n45025 = \m5_data_i[23]_pad  & ~n13627 ;
  assign n45026 = n13652 & n45025 ;
  assign n45027 = ~n45024 & ~n45026 ;
  assign n45028 = n45022 & n45027 ;
  assign n45029 = \m4_data_i[23]_pad  & n13627 ;
  assign n45030 = n13652 & n45029 ;
  assign n45031 = \m6_data_i[23]_pad  & n13627 ;
  assign n45032 = n13644 & n45031 ;
  assign n45033 = ~n45030 & ~n45032 ;
  assign n45034 = \m1_data_i[23]_pad  & ~n13627 ;
  assign n45035 = n13620 & n45034 ;
  assign n45036 = \m2_data_i[23]_pad  & n13627 ;
  assign n45037 = n13635 & n45036 ;
  assign n45038 = ~n45035 & ~n45037 ;
  assign n45039 = n45033 & n45038 ;
  assign n45040 = n45028 & n45039 ;
  assign n45041 = \m3_data_i[24]_pad  & ~n13627 ;
  assign n45042 = n13635 & n45041 ;
  assign n45043 = \m4_data_i[24]_pad  & n13627 ;
  assign n45044 = n13652 & n45043 ;
  assign n45045 = ~n45042 & ~n45044 ;
  assign n45046 = \m6_data_i[24]_pad  & n13627 ;
  assign n45047 = n13644 & n45046 ;
  assign n45048 = \m2_data_i[24]_pad  & n13627 ;
  assign n45049 = n13635 & n45048 ;
  assign n45050 = ~n45047 & ~n45049 ;
  assign n45051 = n45045 & n45050 ;
  assign n45052 = \m5_data_i[24]_pad  & ~n13627 ;
  assign n45053 = n13652 & n45052 ;
  assign n45054 = \m1_data_i[24]_pad  & ~n13627 ;
  assign n45055 = n13620 & n45054 ;
  assign n45056 = ~n45053 & ~n45055 ;
  assign n45057 = \m0_data_i[24]_pad  & n13627 ;
  assign n45058 = n13620 & n45057 ;
  assign n45059 = \m7_data_i[24]_pad  & ~n13627 ;
  assign n45060 = n13644 & n45059 ;
  assign n45061 = ~n45058 & ~n45060 ;
  assign n45062 = n45056 & n45061 ;
  assign n45063 = n45051 & n45062 ;
  assign n45064 = \m3_data_i[25]_pad  & ~n13627 ;
  assign n45065 = n13635 & n45064 ;
  assign n45066 = \m4_data_i[25]_pad  & n13627 ;
  assign n45067 = n13652 & n45066 ;
  assign n45068 = ~n45065 & ~n45067 ;
  assign n45069 = \m6_data_i[25]_pad  & n13627 ;
  assign n45070 = n13644 & n45069 ;
  assign n45071 = \m2_data_i[25]_pad  & n13627 ;
  assign n45072 = n13635 & n45071 ;
  assign n45073 = ~n45070 & ~n45072 ;
  assign n45074 = n45068 & n45073 ;
  assign n45075 = \m5_data_i[25]_pad  & ~n13627 ;
  assign n45076 = n13652 & n45075 ;
  assign n45077 = \m1_data_i[25]_pad  & ~n13627 ;
  assign n45078 = n13620 & n45077 ;
  assign n45079 = ~n45076 & ~n45078 ;
  assign n45080 = \m0_data_i[25]_pad  & n13627 ;
  assign n45081 = n13620 & n45080 ;
  assign n45082 = \m7_data_i[25]_pad  & ~n13627 ;
  assign n45083 = n13644 & n45082 ;
  assign n45084 = ~n45081 & ~n45083 ;
  assign n45085 = n45079 & n45084 ;
  assign n45086 = n45074 & n45085 ;
  assign n45087 = \m3_data_i[26]_pad  & ~n13627 ;
  assign n45088 = n13635 & n45087 ;
  assign n45089 = \m4_data_i[26]_pad  & n13627 ;
  assign n45090 = n13652 & n45089 ;
  assign n45091 = ~n45088 & ~n45090 ;
  assign n45092 = \m6_data_i[26]_pad  & n13627 ;
  assign n45093 = n13644 & n45092 ;
  assign n45094 = \m2_data_i[26]_pad  & n13627 ;
  assign n45095 = n13635 & n45094 ;
  assign n45096 = ~n45093 & ~n45095 ;
  assign n45097 = n45091 & n45096 ;
  assign n45098 = \m5_data_i[26]_pad  & ~n13627 ;
  assign n45099 = n13652 & n45098 ;
  assign n45100 = \m1_data_i[26]_pad  & ~n13627 ;
  assign n45101 = n13620 & n45100 ;
  assign n45102 = ~n45099 & ~n45101 ;
  assign n45103 = \m0_data_i[26]_pad  & n13627 ;
  assign n45104 = n13620 & n45103 ;
  assign n45105 = \m7_data_i[26]_pad  & ~n13627 ;
  assign n45106 = n13644 & n45105 ;
  assign n45107 = ~n45104 & ~n45106 ;
  assign n45108 = n45102 & n45107 ;
  assign n45109 = n45097 & n45108 ;
  assign n45110 = \m3_data_i[27]_pad  & ~n13627 ;
  assign n45111 = n13635 & n45110 ;
  assign n45112 = \m4_data_i[27]_pad  & n13627 ;
  assign n45113 = n13652 & n45112 ;
  assign n45114 = ~n45111 & ~n45113 ;
  assign n45115 = \m6_data_i[27]_pad  & n13627 ;
  assign n45116 = n13644 & n45115 ;
  assign n45117 = \m2_data_i[27]_pad  & n13627 ;
  assign n45118 = n13635 & n45117 ;
  assign n45119 = ~n45116 & ~n45118 ;
  assign n45120 = n45114 & n45119 ;
  assign n45121 = \m5_data_i[27]_pad  & ~n13627 ;
  assign n45122 = n13652 & n45121 ;
  assign n45123 = \m1_data_i[27]_pad  & ~n13627 ;
  assign n45124 = n13620 & n45123 ;
  assign n45125 = ~n45122 & ~n45124 ;
  assign n45126 = \m0_data_i[27]_pad  & n13627 ;
  assign n45127 = n13620 & n45126 ;
  assign n45128 = \m7_data_i[27]_pad  & ~n13627 ;
  assign n45129 = n13644 & n45128 ;
  assign n45130 = ~n45127 & ~n45129 ;
  assign n45131 = n45125 & n45130 ;
  assign n45132 = n45120 & n45131 ;
  assign n45133 = \m1_data_i[28]_pad  & ~n13627 ;
  assign n45134 = n13620 & n45133 ;
  assign n45135 = \m2_data_i[28]_pad  & n13627 ;
  assign n45136 = n13635 & n45135 ;
  assign n45137 = ~n45134 & ~n45136 ;
  assign n45138 = \m0_data_i[28]_pad  & n13627 ;
  assign n45139 = n13620 & n45138 ;
  assign n45140 = \m4_data_i[28]_pad  & n13627 ;
  assign n45141 = n13652 & n45140 ;
  assign n45142 = ~n45139 & ~n45141 ;
  assign n45143 = n45137 & n45142 ;
  assign n45144 = \m7_data_i[28]_pad  & ~n13627 ;
  assign n45145 = n13644 & n45144 ;
  assign n45146 = \m3_data_i[28]_pad  & ~n13627 ;
  assign n45147 = n13635 & n45146 ;
  assign n45148 = ~n45145 & ~n45147 ;
  assign n45149 = \m6_data_i[28]_pad  & n13627 ;
  assign n45150 = n13644 & n45149 ;
  assign n45151 = \m5_data_i[28]_pad  & ~n13627 ;
  assign n45152 = n13652 & n45151 ;
  assign n45153 = ~n45150 & ~n45152 ;
  assign n45154 = n45148 & n45153 ;
  assign n45155 = n45143 & n45154 ;
  assign n45156 = \m3_data_i[29]_pad  & ~n13627 ;
  assign n45157 = n13635 & n45156 ;
  assign n45158 = \m4_data_i[29]_pad  & n13627 ;
  assign n45159 = n13652 & n45158 ;
  assign n45160 = ~n45157 & ~n45159 ;
  assign n45161 = \m6_data_i[29]_pad  & n13627 ;
  assign n45162 = n13644 & n45161 ;
  assign n45163 = \m7_data_i[29]_pad  & ~n13627 ;
  assign n45164 = n13644 & n45163 ;
  assign n45165 = ~n45162 & ~n45164 ;
  assign n45166 = n45160 & n45165 ;
  assign n45167 = \m5_data_i[29]_pad  & ~n13627 ;
  assign n45168 = n13652 & n45167 ;
  assign n45169 = \m0_data_i[29]_pad  & n13627 ;
  assign n45170 = n13620 & n45169 ;
  assign n45171 = ~n45168 & ~n45170 ;
  assign n45172 = \m1_data_i[29]_pad  & ~n13627 ;
  assign n45173 = n13620 & n45172 ;
  assign n45174 = \m2_data_i[29]_pad  & n13627 ;
  assign n45175 = n13635 & n45174 ;
  assign n45176 = ~n45173 & ~n45175 ;
  assign n45177 = n45171 & n45176 ;
  assign n45178 = n45166 & n45177 ;
  assign n45179 = \m1_data_i[2]_pad  & ~n13627 ;
  assign n45180 = n13620 & n45179 ;
  assign n45181 = \m2_data_i[2]_pad  & n13627 ;
  assign n45182 = n13635 & n45181 ;
  assign n45183 = ~n45180 & ~n45182 ;
  assign n45184 = \m0_data_i[2]_pad  & n13627 ;
  assign n45185 = n13620 & n45184 ;
  assign n45186 = \m4_data_i[2]_pad  & n13627 ;
  assign n45187 = n13652 & n45186 ;
  assign n45188 = ~n45185 & ~n45187 ;
  assign n45189 = n45183 & n45188 ;
  assign n45190 = \m7_data_i[2]_pad  & ~n13627 ;
  assign n45191 = n13644 & n45190 ;
  assign n45192 = \m3_data_i[2]_pad  & ~n13627 ;
  assign n45193 = n13635 & n45192 ;
  assign n45194 = ~n45191 & ~n45193 ;
  assign n45195 = \m6_data_i[2]_pad  & n13627 ;
  assign n45196 = n13644 & n45195 ;
  assign n45197 = \m5_data_i[2]_pad  & ~n13627 ;
  assign n45198 = n13652 & n45197 ;
  assign n45199 = ~n45196 & ~n45198 ;
  assign n45200 = n45194 & n45199 ;
  assign n45201 = n45189 & n45200 ;
  assign n45202 = \m3_data_i[30]_pad  & ~n13627 ;
  assign n45203 = n13635 & n45202 ;
  assign n45204 = \m4_data_i[30]_pad  & n13627 ;
  assign n45205 = n13652 & n45204 ;
  assign n45206 = ~n45203 & ~n45205 ;
  assign n45207 = \m6_data_i[30]_pad  & n13627 ;
  assign n45208 = n13644 & n45207 ;
  assign n45209 = \m2_data_i[30]_pad  & n13627 ;
  assign n45210 = n13635 & n45209 ;
  assign n45211 = ~n45208 & ~n45210 ;
  assign n45212 = n45206 & n45211 ;
  assign n45213 = \m5_data_i[30]_pad  & ~n13627 ;
  assign n45214 = n13652 & n45213 ;
  assign n45215 = \m1_data_i[30]_pad  & ~n13627 ;
  assign n45216 = n13620 & n45215 ;
  assign n45217 = ~n45214 & ~n45216 ;
  assign n45218 = \m0_data_i[30]_pad  & n13627 ;
  assign n45219 = n13620 & n45218 ;
  assign n45220 = \m7_data_i[30]_pad  & ~n13627 ;
  assign n45221 = n13644 & n45220 ;
  assign n45222 = ~n45219 & ~n45221 ;
  assign n45223 = n45217 & n45222 ;
  assign n45224 = n45212 & n45223 ;
  assign n45225 = \m0_data_i[31]_pad  & n13627 ;
  assign n45226 = n13620 & n45225 ;
  assign n45227 = \m7_data_i[31]_pad  & ~n13627 ;
  assign n45228 = n13644 & n45227 ;
  assign n45229 = ~n45226 & ~n45228 ;
  assign n45230 = \m1_data_i[31]_pad  & ~n13627 ;
  assign n45231 = n13620 & n45230 ;
  assign n45232 = \m4_data_i[31]_pad  & n13627 ;
  assign n45233 = n13652 & n45232 ;
  assign n45234 = ~n45231 & ~n45233 ;
  assign n45235 = n45229 & n45234 ;
  assign n45236 = \m2_data_i[31]_pad  & n13627 ;
  assign n45237 = n13635 & n45236 ;
  assign n45238 = \m3_data_i[31]_pad  & ~n13627 ;
  assign n45239 = n13635 & n45238 ;
  assign n45240 = ~n45237 & ~n45239 ;
  assign n45241 = \m6_data_i[31]_pad  & n13627 ;
  assign n45242 = n13644 & n45241 ;
  assign n45243 = \m5_data_i[31]_pad  & ~n13627 ;
  assign n45244 = n13652 & n45243 ;
  assign n45245 = ~n45242 & ~n45244 ;
  assign n45246 = n45240 & n45245 ;
  assign n45247 = n45235 & n45246 ;
  assign n45248 = \m1_data_i[3]_pad  & ~n13627 ;
  assign n45249 = n13620 & n45248 ;
  assign n45250 = \m2_data_i[3]_pad  & n13627 ;
  assign n45251 = n13635 & n45250 ;
  assign n45252 = ~n45249 & ~n45251 ;
  assign n45253 = \m0_data_i[3]_pad  & n13627 ;
  assign n45254 = n13620 & n45253 ;
  assign n45255 = \m4_data_i[3]_pad  & n13627 ;
  assign n45256 = n13652 & n45255 ;
  assign n45257 = ~n45254 & ~n45256 ;
  assign n45258 = n45252 & n45257 ;
  assign n45259 = \m7_data_i[3]_pad  & ~n13627 ;
  assign n45260 = n13644 & n45259 ;
  assign n45261 = \m3_data_i[3]_pad  & ~n13627 ;
  assign n45262 = n13635 & n45261 ;
  assign n45263 = ~n45260 & ~n45262 ;
  assign n45264 = \m6_data_i[3]_pad  & n13627 ;
  assign n45265 = n13644 & n45264 ;
  assign n45266 = \m5_data_i[3]_pad  & ~n13627 ;
  assign n45267 = n13652 & n45266 ;
  assign n45268 = ~n45265 & ~n45267 ;
  assign n45269 = n45263 & n45268 ;
  assign n45270 = n45258 & n45269 ;
  assign n45271 = \m0_data_i[4]_pad  & n13627 ;
  assign n45272 = n13620 & n45271 ;
  assign n45273 = \m7_data_i[4]_pad  & ~n13627 ;
  assign n45274 = n13644 & n45273 ;
  assign n45275 = ~n45272 & ~n45274 ;
  assign n45276 = \m6_data_i[4]_pad  & n13627 ;
  assign n45277 = n13644 & n45276 ;
  assign n45278 = \m2_data_i[4]_pad  & n13627 ;
  assign n45279 = n13635 & n45278 ;
  assign n45280 = ~n45277 & ~n45279 ;
  assign n45281 = n45275 & n45280 ;
  assign n45282 = \m5_data_i[4]_pad  & ~n13627 ;
  assign n45283 = n13652 & n45282 ;
  assign n45284 = \m1_data_i[4]_pad  & ~n13627 ;
  assign n45285 = n13620 & n45284 ;
  assign n45286 = ~n45283 & ~n45285 ;
  assign n45287 = \m3_data_i[4]_pad  & ~n13627 ;
  assign n45288 = n13635 & n45287 ;
  assign n45289 = \m4_data_i[4]_pad  & n13627 ;
  assign n45290 = n13652 & n45289 ;
  assign n45291 = ~n45288 & ~n45290 ;
  assign n45292 = n45286 & n45291 ;
  assign n45293 = n45281 & n45292 ;
  assign n45294 = \m1_data_i[5]_pad  & ~n13627 ;
  assign n45295 = n13620 & n45294 ;
  assign n45296 = \m2_data_i[5]_pad  & n13627 ;
  assign n45297 = n13635 & n45296 ;
  assign n45298 = ~n45295 & ~n45297 ;
  assign n45299 = \m0_data_i[5]_pad  & n13627 ;
  assign n45300 = n13620 & n45299 ;
  assign n45301 = \m4_data_i[5]_pad  & n13627 ;
  assign n45302 = n13652 & n45301 ;
  assign n45303 = ~n45300 & ~n45302 ;
  assign n45304 = n45298 & n45303 ;
  assign n45305 = \m7_data_i[5]_pad  & ~n13627 ;
  assign n45306 = n13644 & n45305 ;
  assign n45307 = \m3_data_i[5]_pad  & ~n13627 ;
  assign n45308 = n13635 & n45307 ;
  assign n45309 = ~n45306 & ~n45308 ;
  assign n45310 = \m6_data_i[5]_pad  & n13627 ;
  assign n45311 = n13644 & n45310 ;
  assign n45312 = \m5_data_i[5]_pad  & ~n13627 ;
  assign n45313 = n13652 & n45312 ;
  assign n45314 = ~n45311 & ~n45313 ;
  assign n45315 = n45309 & n45314 ;
  assign n45316 = n45304 & n45315 ;
  assign n45317 = \m6_data_i[6]_pad  & n13627 ;
  assign n45318 = n13644 & n45317 ;
  assign n45319 = \m5_data_i[6]_pad  & ~n13627 ;
  assign n45320 = n13652 & n45319 ;
  assign n45321 = ~n45318 & ~n45320 ;
  assign n45322 = \m0_data_i[6]_pad  & n13627 ;
  assign n45323 = n13620 & n45322 ;
  assign n45324 = \m2_data_i[6]_pad  & n13627 ;
  assign n45325 = n13635 & n45324 ;
  assign n45326 = ~n45323 & ~n45325 ;
  assign n45327 = n45321 & n45326 ;
  assign n45328 = \m7_data_i[6]_pad  & ~n13627 ;
  assign n45329 = n13644 & n45328 ;
  assign n45330 = \m1_data_i[6]_pad  & ~n13627 ;
  assign n45331 = n13620 & n45330 ;
  assign n45332 = ~n45329 & ~n45331 ;
  assign n45333 = \m3_data_i[6]_pad  & ~n13627 ;
  assign n45334 = n13635 & n45333 ;
  assign n45335 = \m4_data_i[6]_pad  & n13627 ;
  assign n45336 = n13652 & n45335 ;
  assign n45337 = ~n45334 & ~n45336 ;
  assign n45338 = n45332 & n45337 ;
  assign n45339 = n45327 & n45338 ;
  assign n45340 = \m3_data_i[7]_pad  & ~n13627 ;
  assign n45341 = n13635 & n45340 ;
  assign n45342 = \m4_data_i[7]_pad  & n13627 ;
  assign n45343 = n13652 & n45342 ;
  assign n45344 = ~n45341 & ~n45343 ;
  assign n45345 = \m6_data_i[7]_pad  & n13627 ;
  assign n45346 = n13644 & n45345 ;
  assign n45347 = \m7_data_i[7]_pad  & ~n13627 ;
  assign n45348 = n13644 & n45347 ;
  assign n45349 = ~n45346 & ~n45348 ;
  assign n45350 = n45344 & n45349 ;
  assign n45351 = \m5_data_i[7]_pad  & ~n13627 ;
  assign n45352 = n13652 & n45351 ;
  assign n45353 = \m0_data_i[7]_pad  & n13627 ;
  assign n45354 = n13620 & n45353 ;
  assign n45355 = ~n45352 & ~n45354 ;
  assign n45356 = \m1_data_i[7]_pad  & ~n13627 ;
  assign n45357 = n13620 & n45356 ;
  assign n45358 = \m2_data_i[7]_pad  & n13627 ;
  assign n45359 = n13635 & n45358 ;
  assign n45360 = ~n45357 & ~n45359 ;
  assign n45361 = n45355 & n45360 ;
  assign n45362 = n45350 & n45361 ;
  assign n45363 = \m1_data_i[8]_pad  & ~n13627 ;
  assign n45364 = n13620 & n45363 ;
  assign n45365 = \m2_data_i[8]_pad  & n13627 ;
  assign n45366 = n13635 & n45365 ;
  assign n45367 = ~n45364 & ~n45366 ;
  assign n45368 = \m0_data_i[8]_pad  & n13627 ;
  assign n45369 = n13620 & n45368 ;
  assign n45370 = \m4_data_i[8]_pad  & n13627 ;
  assign n45371 = n13652 & n45370 ;
  assign n45372 = ~n45369 & ~n45371 ;
  assign n45373 = n45367 & n45372 ;
  assign n45374 = \m7_data_i[8]_pad  & ~n13627 ;
  assign n45375 = n13644 & n45374 ;
  assign n45376 = \m3_data_i[8]_pad  & ~n13627 ;
  assign n45377 = n13635 & n45376 ;
  assign n45378 = ~n45375 & ~n45377 ;
  assign n45379 = \m6_data_i[8]_pad  & n13627 ;
  assign n45380 = n13644 & n45379 ;
  assign n45381 = \m5_data_i[8]_pad  & ~n13627 ;
  assign n45382 = n13652 & n45381 ;
  assign n45383 = ~n45380 & ~n45382 ;
  assign n45384 = n45378 & n45383 ;
  assign n45385 = n45373 & n45384 ;
  assign n45386 = \m1_data_i[9]_pad  & ~n13627 ;
  assign n45387 = n13620 & n45386 ;
  assign n45388 = \m2_data_i[9]_pad  & n13627 ;
  assign n45389 = n13635 & n45388 ;
  assign n45390 = ~n45387 & ~n45389 ;
  assign n45391 = \m0_data_i[9]_pad  & n13627 ;
  assign n45392 = n13620 & n45391 ;
  assign n45393 = \m4_data_i[9]_pad  & n13627 ;
  assign n45394 = n13652 & n45393 ;
  assign n45395 = ~n45392 & ~n45394 ;
  assign n45396 = n45390 & n45395 ;
  assign n45397 = \m7_data_i[9]_pad  & ~n13627 ;
  assign n45398 = n13644 & n45397 ;
  assign n45399 = \m3_data_i[9]_pad  & ~n13627 ;
  assign n45400 = n13635 & n45399 ;
  assign n45401 = ~n45398 & ~n45400 ;
  assign n45402 = \m6_data_i[9]_pad  & n13627 ;
  assign n45403 = n13644 & n45402 ;
  assign n45404 = \m5_data_i[9]_pad  & ~n13627 ;
  assign n45405 = n13652 & n45404 ;
  assign n45406 = ~n45403 & ~n45405 ;
  assign n45407 = n45401 & n45406 ;
  assign n45408 = n45396 & n45407 ;
  assign n45409 = \m3_sel_i[0]_pad  & ~n13627 ;
  assign n45410 = n13635 & n45409 ;
  assign n45411 = \m4_sel_i[0]_pad  & n13627 ;
  assign n45412 = n13652 & n45411 ;
  assign n45413 = ~n45410 & ~n45412 ;
  assign n45414 = \m6_sel_i[0]_pad  & n13627 ;
  assign n45415 = n13644 & n45414 ;
  assign n45416 = \m2_sel_i[0]_pad  & n13627 ;
  assign n45417 = n13635 & n45416 ;
  assign n45418 = ~n45415 & ~n45417 ;
  assign n45419 = n45413 & n45418 ;
  assign n45420 = \m5_sel_i[0]_pad  & ~n13627 ;
  assign n45421 = n13652 & n45420 ;
  assign n45422 = \m1_sel_i[0]_pad  & ~n13627 ;
  assign n45423 = n13620 & n45422 ;
  assign n45424 = ~n45421 & ~n45423 ;
  assign n45425 = \m0_sel_i[0]_pad  & n13627 ;
  assign n45426 = n13620 & n45425 ;
  assign n45427 = \m7_sel_i[0]_pad  & ~n13627 ;
  assign n45428 = n13644 & n45427 ;
  assign n45429 = ~n45426 & ~n45428 ;
  assign n45430 = n45424 & n45429 ;
  assign n45431 = n45419 & n45430 ;
  assign n45432 = \m1_sel_i[1]_pad  & ~n13627 ;
  assign n45433 = n13620 & n45432 ;
  assign n45434 = \m2_sel_i[1]_pad  & n13627 ;
  assign n45435 = n13635 & n45434 ;
  assign n45436 = ~n45433 & ~n45435 ;
  assign n45437 = \m0_sel_i[1]_pad  & n13627 ;
  assign n45438 = n13620 & n45437 ;
  assign n45439 = \m4_sel_i[1]_pad  & n13627 ;
  assign n45440 = n13652 & n45439 ;
  assign n45441 = ~n45438 & ~n45440 ;
  assign n45442 = n45436 & n45441 ;
  assign n45443 = \m7_sel_i[1]_pad  & ~n13627 ;
  assign n45444 = n13644 & n45443 ;
  assign n45445 = \m3_sel_i[1]_pad  & ~n13627 ;
  assign n45446 = n13635 & n45445 ;
  assign n45447 = ~n45444 & ~n45446 ;
  assign n45448 = \m6_sel_i[1]_pad  & n13627 ;
  assign n45449 = n13644 & n45448 ;
  assign n45450 = \m5_sel_i[1]_pad  & ~n13627 ;
  assign n45451 = n13652 & n45450 ;
  assign n45452 = ~n45449 & ~n45451 ;
  assign n45453 = n45447 & n45452 ;
  assign n45454 = n45442 & n45453 ;
  assign n45455 = \m1_sel_i[2]_pad  & ~n13627 ;
  assign n45456 = n13620 & n45455 ;
  assign n45457 = \m2_sel_i[2]_pad  & n13627 ;
  assign n45458 = n13635 & n45457 ;
  assign n45459 = ~n45456 & ~n45458 ;
  assign n45460 = \m0_sel_i[2]_pad  & n13627 ;
  assign n45461 = n13620 & n45460 ;
  assign n45462 = \m4_sel_i[2]_pad  & n13627 ;
  assign n45463 = n13652 & n45462 ;
  assign n45464 = ~n45461 & ~n45463 ;
  assign n45465 = n45459 & n45464 ;
  assign n45466 = \m7_sel_i[2]_pad  & ~n13627 ;
  assign n45467 = n13644 & n45466 ;
  assign n45468 = \m3_sel_i[2]_pad  & ~n13627 ;
  assign n45469 = n13635 & n45468 ;
  assign n45470 = ~n45467 & ~n45469 ;
  assign n45471 = \m6_sel_i[2]_pad  & n13627 ;
  assign n45472 = n13644 & n45471 ;
  assign n45473 = \m5_sel_i[2]_pad  & ~n13627 ;
  assign n45474 = n13652 & n45473 ;
  assign n45475 = ~n45472 & ~n45474 ;
  assign n45476 = n45470 & n45475 ;
  assign n45477 = n45465 & n45476 ;
  assign n45478 = \m0_sel_i[3]_pad  & n13627 ;
  assign n45479 = n13620 & n45478 ;
  assign n45480 = \m7_sel_i[3]_pad  & ~n13627 ;
  assign n45481 = n13644 & n45480 ;
  assign n45482 = ~n45479 & ~n45481 ;
  assign n45483 = \m3_sel_i[3]_pad  & ~n13627 ;
  assign n45484 = n13635 & n45483 ;
  assign n45485 = \m2_sel_i[3]_pad  & n13627 ;
  assign n45486 = n13635 & n45485 ;
  assign n45487 = ~n45484 & ~n45486 ;
  assign n45488 = n45482 & n45487 ;
  assign n45489 = \m4_sel_i[3]_pad  & n13627 ;
  assign n45490 = n13652 & n45489 ;
  assign n45491 = \m1_sel_i[3]_pad  & ~n13627 ;
  assign n45492 = n13620 & n45491 ;
  assign n45493 = ~n45490 & ~n45492 ;
  assign n45494 = \m6_sel_i[3]_pad  & n13627 ;
  assign n45495 = n13644 & n45494 ;
  assign n45496 = \m5_sel_i[3]_pad  & ~n13627 ;
  assign n45497 = n13652 & n45496 ;
  assign n45498 = ~n45495 & ~n45497 ;
  assign n45499 = n45493 & n45498 ;
  assign n45500 = n45488 & n45499 ;
  assign n45501 = \m5_stb_i_pad  & n14987 ;
  assign n45502 = ~n13627 & n45501 ;
  assign n45503 = n13652 & n45502 ;
  assign n45504 = \m4_stb_i_pad  & n14723 ;
  assign n45505 = n13627 & n45504 ;
  assign n45506 = n13652 & n45505 ;
  assign n45507 = ~n45503 & ~n45506 ;
  assign n45508 = \m2_stb_i_pad  & n14883 ;
  assign n45509 = n13627 & n45508 ;
  assign n45510 = n13635 & n45509 ;
  assign n45511 = \m6_stb_i_pad  & n14681 ;
  assign n45512 = n13627 & n45511 ;
  assign n45513 = n13644 & n45512 ;
  assign n45514 = ~n45510 & ~n45513 ;
  assign n45515 = n45507 & n45514 ;
  assign n45516 = \m3_stb_i_pad  & n14745 ;
  assign n45517 = ~n13627 & n45516 ;
  assign n45518 = n13635 & n45517 ;
  assign n45519 = \m7_stb_i_pad  & n15078 ;
  assign n45520 = ~n13627 & n45519 ;
  assign n45521 = n13644 & n45520 ;
  assign n45522 = ~n45518 & ~n45521 ;
  assign n45523 = \m1_stb_i_pad  & n14833 ;
  assign n45524 = ~n13627 & n45523 ;
  assign n45525 = n13620 & n45524 ;
  assign n45526 = \m0_stb_i_pad  & n14782 ;
  assign n45527 = n13627 & n45526 ;
  assign n45528 = n13620 & n45527 ;
  assign n45529 = ~n45525 & ~n45528 ;
  assign n45530 = n45522 & n45529 ;
  assign n45531 = n45515 & n45530 ;
  assign n45532 = \m3_we_i_pad  & ~n13627 ;
  assign n45533 = n13635 & n45532 ;
  assign n45534 = \m4_we_i_pad  & n13627 ;
  assign n45535 = n13652 & n45534 ;
  assign n45536 = ~n45533 & ~n45535 ;
  assign n45537 = \m6_we_i_pad  & n13627 ;
  assign n45538 = n13644 & n45537 ;
  assign n45539 = \m7_we_i_pad  & ~n13627 ;
  assign n45540 = n13644 & n45539 ;
  assign n45541 = ~n45538 & ~n45540 ;
  assign n45542 = n45536 & n45541 ;
  assign n45543 = \m5_we_i_pad  & ~n13627 ;
  assign n45544 = n13652 & n45543 ;
  assign n45545 = \m0_we_i_pad  & n13627 ;
  assign n45546 = n13620 & n45545 ;
  assign n45547 = ~n45544 & ~n45546 ;
  assign n45548 = \m1_we_i_pad  & ~n13627 ;
  assign n45549 = n13620 & n45548 ;
  assign n45550 = \m2_we_i_pad  & n13627 ;
  assign n45551 = n13635 & n45550 ;
  assign n45552 = ~n45549 & ~n45551 ;
  assign n45553 = n45547 & n45552 ;
  assign n45554 = n45542 & n45553 ;
  assign n45555 = \m0_addr_i[0]_pad  & n13697 ;
  assign n45556 = n13705 & n45555 ;
  assign n45557 = \m7_addr_i[0]_pad  & ~n13697 ;
  assign n45558 = n13690 & n45557 ;
  assign n45559 = ~n45556 & ~n45558 ;
  assign n45560 = \m3_addr_i[0]_pad  & ~n13697 ;
  assign n45561 = n13714 & n45560 ;
  assign n45562 = \m5_addr_i[0]_pad  & ~n13697 ;
  assign n45563 = n13722 & n45562 ;
  assign n45564 = ~n45561 & ~n45563 ;
  assign n45565 = n45559 & n45564 ;
  assign n45566 = \m4_addr_i[0]_pad  & n13697 ;
  assign n45567 = n13722 & n45566 ;
  assign n45568 = \m6_addr_i[0]_pad  & n13697 ;
  assign n45569 = n13690 & n45568 ;
  assign n45570 = ~n45567 & ~n45569 ;
  assign n45571 = \m1_addr_i[0]_pad  & ~n13697 ;
  assign n45572 = n13705 & n45571 ;
  assign n45573 = \m2_addr_i[0]_pad  & n13697 ;
  assign n45574 = n13714 & n45573 ;
  assign n45575 = ~n45572 & ~n45574 ;
  assign n45576 = n45570 & n45575 ;
  assign n45577 = n45565 & n45576 ;
  assign n45578 = \m3_addr_i[10]_pad  & ~n13697 ;
  assign n45579 = n13714 & n45578 ;
  assign n45580 = \m4_addr_i[10]_pad  & n13697 ;
  assign n45581 = n13722 & n45580 ;
  assign n45582 = ~n45579 & ~n45581 ;
  assign n45583 = \m6_addr_i[10]_pad  & n13697 ;
  assign n45584 = n13690 & n45583 ;
  assign n45585 = \m7_addr_i[10]_pad  & ~n13697 ;
  assign n45586 = n13690 & n45585 ;
  assign n45587 = ~n45584 & ~n45586 ;
  assign n45588 = n45582 & n45587 ;
  assign n45589 = \m5_addr_i[10]_pad  & ~n13697 ;
  assign n45590 = n13722 & n45589 ;
  assign n45591 = \m0_addr_i[10]_pad  & n13697 ;
  assign n45592 = n13705 & n45591 ;
  assign n45593 = ~n45590 & ~n45592 ;
  assign n45594 = \m1_addr_i[10]_pad  & ~n13697 ;
  assign n45595 = n13705 & n45594 ;
  assign n45596 = \m2_addr_i[10]_pad  & n13697 ;
  assign n45597 = n13714 & n45596 ;
  assign n45598 = ~n45595 & ~n45597 ;
  assign n45599 = n45593 & n45598 ;
  assign n45600 = n45588 & n45599 ;
  assign n45601 = \m1_addr_i[11]_pad  & ~n13697 ;
  assign n45602 = n13705 & n45601 ;
  assign n45603 = \m2_addr_i[11]_pad  & n13697 ;
  assign n45604 = n13714 & n45603 ;
  assign n45605 = ~n45602 & ~n45604 ;
  assign n45606 = \m6_addr_i[11]_pad  & n13697 ;
  assign n45607 = n13690 & n45606 ;
  assign n45608 = \m7_addr_i[11]_pad  & ~n13697 ;
  assign n45609 = n13690 & n45608 ;
  assign n45610 = ~n45607 & ~n45609 ;
  assign n45611 = n45605 & n45610 ;
  assign n45612 = \m5_addr_i[11]_pad  & ~n13697 ;
  assign n45613 = n13722 & n45612 ;
  assign n45614 = \m0_addr_i[11]_pad  & n13697 ;
  assign n45615 = n13705 & n45614 ;
  assign n45616 = ~n45613 & ~n45615 ;
  assign n45617 = \m3_addr_i[11]_pad  & ~n13697 ;
  assign n45618 = n13714 & n45617 ;
  assign n45619 = \m4_addr_i[11]_pad  & n13697 ;
  assign n45620 = n13722 & n45619 ;
  assign n45621 = ~n45618 & ~n45620 ;
  assign n45622 = n45616 & n45621 ;
  assign n45623 = n45611 & n45622 ;
  assign n45624 = \m1_addr_i[12]_pad  & ~n13697 ;
  assign n45625 = n13705 & n45624 ;
  assign n45626 = \m2_addr_i[12]_pad  & n13697 ;
  assign n45627 = n13714 & n45626 ;
  assign n45628 = ~n45625 & ~n45627 ;
  assign n45629 = \m6_addr_i[12]_pad  & n13697 ;
  assign n45630 = n13690 & n45629 ;
  assign n45631 = \m7_addr_i[12]_pad  & ~n13697 ;
  assign n45632 = n13690 & n45631 ;
  assign n45633 = ~n45630 & ~n45632 ;
  assign n45634 = n45628 & n45633 ;
  assign n45635 = \m5_addr_i[12]_pad  & ~n13697 ;
  assign n45636 = n13722 & n45635 ;
  assign n45637 = \m0_addr_i[12]_pad  & n13697 ;
  assign n45638 = n13705 & n45637 ;
  assign n45639 = ~n45636 & ~n45638 ;
  assign n45640 = \m3_addr_i[12]_pad  & ~n13697 ;
  assign n45641 = n13714 & n45640 ;
  assign n45642 = \m4_addr_i[12]_pad  & n13697 ;
  assign n45643 = n13722 & n45642 ;
  assign n45644 = ~n45641 & ~n45643 ;
  assign n45645 = n45639 & n45644 ;
  assign n45646 = n45634 & n45645 ;
  assign n45647 = \m3_addr_i[13]_pad  & ~n13697 ;
  assign n45648 = n13714 & n45647 ;
  assign n45649 = \m4_addr_i[13]_pad  & n13697 ;
  assign n45650 = n13722 & n45649 ;
  assign n45651 = ~n45648 & ~n45650 ;
  assign n45652 = \m6_addr_i[13]_pad  & n13697 ;
  assign n45653 = n13690 & n45652 ;
  assign n45654 = \m2_addr_i[13]_pad  & n13697 ;
  assign n45655 = n13714 & n45654 ;
  assign n45656 = ~n45653 & ~n45655 ;
  assign n45657 = n45651 & n45656 ;
  assign n45658 = \m5_addr_i[13]_pad  & ~n13697 ;
  assign n45659 = n13722 & n45658 ;
  assign n45660 = \m1_addr_i[13]_pad  & ~n13697 ;
  assign n45661 = n13705 & n45660 ;
  assign n45662 = ~n45659 & ~n45661 ;
  assign n45663 = \m0_addr_i[13]_pad  & n13697 ;
  assign n45664 = n13705 & n45663 ;
  assign n45665 = \m7_addr_i[13]_pad  & ~n13697 ;
  assign n45666 = n13690 & n45665 ;
  assign n45667 = ~n45664 & ~n45666 ;
  assign n45668 = n45662 & n45667 ;
  assign n45669 = n45657 & n45668 ;
  assign n45670 = \m3_addr_i[14]_pad  & ~n13697 ;
  assign n45671 = n13714 & n45670 ;
  assign n45672 = \m4_addr_i[14]_pad  & n13697 ;
  assign n45673 = n13722 & n45672 ;
  assign n45674 = ~n45671 & ~n45673 ;
  assign n45675 = \m6_addr_i[14]_pad  & n13697 ;
  assign n45676 = n13690 & n45675 ;
  assign n45677 = \m2_addr_i[14]_pad  & n13697 ;
  assign n45678 = n13714 & n45677 ;
  assign n45679 = ~n45676 & ~n45678 ;
  assign n45680 = n45674 & n45679 ;
  assign n45681 = \m5_addr_i[14]_pad  & ~n13697 ;
  assign n45682 = n13722 & n45681 ;
  assign n45683 = \m1_addr_i[14]_pad  & ~n13697 ;
  assign n45684 = n13705 & n45683 ;
  assign n45685 = ~n45682 & ~n45684 ;
  assign n45686 = \m0_addr_i[14]_pad  & n13697 ;
  assign n45687 = n13705 & n45686 ;
  assign n45688 = \m7_addr_i[14]_pad  & ~n13697 ;
  assign n45689 = n13690 & n45688 ;
  assign n45690 = ~n45687 & ~n45689 ;
  assign n45691 = n45685 & n45690 ;
  assign n45692 = n45680 & n45691 ;
  assign n45693 = \m3_addr_i[15]_pad  & ~n13697 ;
  assign n45694 = n13714 & n45693 ;
  assign n45695 = \m4_addr_i[15]_pad  & n13697 ;
  assign n45696 = n13722 & n45695 ;
  assign n45697 = ~n45694 & ~n45696 ;
  assign n45698 = \m6_addr_i[15]_pad  & n13697 ;
  assign n45699 = n13690 & n45698 ;
  assign n45700 = \m2_addr_i[15]_pad  & n13697 ;
  assign n45701 = n13714 & n45700 ;
  assign n45702 = ~n45699 & ~n45701 ;
  assign n45703 = n45697 & n45702 ;
  assign n45704 = \m5_addr_i[15]_pad  & ~n13697 ;
  assign n45705 = n13722 & n45704 ;
  assign n45706 = \m1_addr_i[15]_pad  & ~n13697 ;
  assign n45707 = n13705 & n45706 ;
  assign n45708 = ~n45705 & ~n45707 ;
  assign n45709 = \m0_addr_i[15]_pad  & n13697 ;
  assign n45710 = n13705 & n45709 ;
  assign n45711 = \m7_addr_i[15]_pad  & ~n13697 ;
  assign n45712 = n13690 & n45711 ;
  assign n45713 = ~n45710 & ~n45712 ;
  assign n45714 = n45708 & n45713 ;
  assign n45715 = n45703 & n45714 ;
  assign n45716 = \m3_addr_i[16]_pad  & ~n13697 ;
  assign n45717 = n13714 & n45716 ;
  assign n45718 = \m4_addr_i[16]_pad  & n13697 ;
  assign n45719 = n13722 & n45718 ;
  assign n45720 = ~n45717 & ~n45719 ;
  assign n45721 = \m6_addr_i[16]_pad  & n13697 ;
  assign n45722 = n13690 & n45721 ;
  assign n45723 = \m2_addr_i[16]_pad  & n13697 ;
  assign n45724 = n13714 & n45723 ;
  assign n45725 = ~n45722 & ~n45724 ;
  assign n45726 = n45720 & n45725 ;
  assign n45727 = \m5_addr_i[16]_pad  & ~n13697 ;
  assign n45728 = n13722 & n45727 ;
  assign n45729 = \m1_addr_i[16]_pad  & ~n13697 ;
  assign n45730 = n13705 & n45729 ;
  assign n45731 = ~n45728 & ~n45730 ;
  assign n45732 = \m0_addr_i[16]_pad  & n13697 ;
  assign n45733 = n13705 & n45732 ;
  assign n45734 = \m7_addr_i[16]_pad  & ~n13697 ;
  assign n45735 = n13690 & n45734 ;
  assign n45736 = ~n45733 & ~n45735 ;
  assign n45737 = n45731 & n45736 ;
  assign n45738 = n45726 & n45737 ;
  assign n45739 = \m1_addr_i[17]_pad  & ~n13697 ;
  assign n45740 = n13705 & n45739 ;
  assign n45741 = \m2_addr_i[17]_pad  & n13697 ;
  assign n45742 = n13714 & n45741 ;
  assign n45743 = ~n45740 & ~n45742 ;
  assign n45744 = \m3_addr_i[17]_pad  & ~n13697 ;
  assign n45745 = n13714 & n45744 ;
  assign n45746 = \m7_addr_i[17]_pad  & ~n13697 ;
  assign n45747 = n13690 & n45746 ;
  assign n45748 = ~n45745 & ~n45747 ;
  assign n45749 = n45743 & n45748 ;
  assign n45750 = \m4_addr_i[17]_pad  & n13697 ;
  assign n45751 = n13722 & n45750 ;
  assign n45752 = \m0_addr_i[17]_pad  & n13697 ;
  assign n45753 = n13705 & n45752 ;
  assign n45754 = ~n45751 & ~n45753 ;
  assign n45755 = \m6_addr_i[17]_pad  & n13697 ;
  assign n45756 = n13690 & n45755 ;
  assign n45757 = \m5_addr_i[17]_pad  & ~n13697 ;
  assign n45758 = n13722 & n45757 ;
  assign n45759 = ~n45756 & ~n45758 ;
  assign n45760 = n45754 & n45759 ;
  assign n45761 = n45749 & n45760 ;
  assign n45762 = \m1_addr_i[18]_pad  & ~n13697 ;
  assign n45763 = n13705 & n45762 ;
  assign n45764 = \m2_addr_i[18]_pad  & n13697 ;
  assign n45765 = n13714 & n45764 ;
  assign n45766 = ~n45763 & ~n45765 ;
  assign n45767 = \m3_addr_i[18]_pad  & ~n13697 ;
  assign n45768 = n13714 & n45767 ;
  assign n45769 = \m7_addr_i[18]_pad  & ~n13697 ;
  assign n45770 = n13690 & n45769 ;
  assign n45771 = ~n45768 & ~n45770 ;
  assign n45772 = n45766 & n45771 ;
  assign n45773 = \m4_addr_i[18]_pad  & n13697 ;
  assign n45774 = n13722 & n45773 ;
  assign n45775 = \m0_addr_i[18]_pad  & n13697 ;
  assign n45776 = n13705 & n45775 ;
  assign n45777 = ~n45774 & ~n45776 ;
  assign n45778 = \m6_addr_i[18]_pad  & n13697 ;
  assign n45779 = n13690 & n45778 ;
  assign n45780 = \m5_addr_i[18]_pad  & ~n13697 ;
  assign n45781 = n13722 & n45780 ;
  assign n45782 = ~n45779 & ~n45781 ;
  assign n45783 = n45777 & n45782 ;
  assign n45784 = n45772 & n45783 ;
  assign n45785 = \m3_addr_i[19]_pad  & ~n13697 ;
  assign n45786 = n13714 & n45785 ;
  assign n45787 = \m4_addr_i[19]_pad  & n13697 ;
  assign n45788 = n13722 & n45787 ;
  assign n45789 = ~n45786 & ~n45788 ;
  assign n45790 = \m6_addr_i[19]_pad  & n13697 ;
  assign n45791 = n13690 & n45790 ;
  assign n45792 = \m7_addr_i[19]_pad  & ~n13697 ;
  assign n45793 = n13690 & n45792 ;
  assign n45794 = ~n45791 & ~n45793 ;
  assign n45795 = n45789 & n45794 ;
  assign n45796 = \m5_addr_i[19]_pad  & ~n13697 ;
  assign n45797 = n13722 & n45796 ;
  assign n45798 = \m0_addr_i[19]_pad  & n13697 ;
  assign n45799 = n13705 & n45798 ;
  assign n45800 = ~n45797 & ~n45799 ;
  assign n45801 = \m1_addr_i[19]_pad  & ~n13697 ;
  assign n45802 = n13705 & n45801 ;
  assign n45803 = \m2_addr_i[19]_pad  & n13697 ;
  assign n45804 = n13714 & n45803 ;
  assign n45805 = ~n45802 & ~n45804 ;
  assign n45806 = n45800 & n45805 ;
  assign n45807 = n45795 & n45806 ;
  assign n45808 = \m3_addr_i[1]_pad  & ~n13697 ;
  assign n45809 = n13714 & n45808 ;
  assign n45810 = \m4_addr_i[1]_pad  & n13697 ;
  assign n45811 = n13722 & n45810 ;
  assign n45812 = ~n45809 & ~n45811 ;
  assign n45813 = \m6_addr_i[1]_pad  & n13697 ;
  assign n45814 = n13690 & n45813 ;
  assign n45815 = \m2_addr_i[1]_pad  & n13697 ;
  assign n45816 = n13714 & n45815 ;
  assign n45817 = ~n45814 & ~n45816 ;
  assign n45818 = n45812 & n45817 ;
  assign n45819 = \m5_addr_i[1]_pad  & ~n13697 ;
  assign n45820 = n13722 & n45819 ;
  assign n45821 = \m1_addr_i[1]_pad  & ~n13697 ;
  assign n45822 = n13705 & n45821 ;
  assign n45823 = ~n45820 & ~n45822 ;
  assign n45824 = \m0_addr_i[1]_pad  & n13697 ;
  assign n45825 = n13705 & n45824 ;
  assign n45826 = \m7_addr_i[1]_pad  & ~n13697 ;
  assign n45827 = n13690 & n45826 ;
  assign n45828 = ~n45825 & ~n45827 ;
  assign n45829 = n45823 & n45828 ;
  assign n45830 = n45818 & n45829 ;
  assign n45831 = \m0_addr_i[20]_pad  & n13697 ;
  assign n45832 = n13705 & n45831 ;
  assign n45833 = \m7_addr_i[20]_pad  & ~n13697 ;
  assign n45834 = n13690 & n45833 ;
  assign n45835 = ~n45832 & ~n45834 ;
  assign n45836 = \m3_addr_i[20]_pad  & ~n13697 ;
  assign n45837 = n13714 & n45836 ;
  assign n45838 = \m2_addr_i[20]_pad  & n13697 ;
  assign n45839 = n13714 & n45838 ;
  assign n45840 = ~n45837 & ~n45839 ;
  assign n45841 = n45835 & n45840 ;
  assign n45842 = \m4_addr_i[20]_pad  & n13697 ;
  assign n45843 = n13722 & n45842 ;
  assign n45844 = \m1_addr_i[20]_pad  & ~n13697 ;
  assign n45845 = n13705 & n45844 ;
  assign n45846 = ~n45843 & ~n45845 ;
  assign n45847 = \m6_addr_i[20]_pad  & n13697 ;
  assign n45848 = n13690 & n45847 ;
  assign n45849 = \m5_addr_i[20]_pad  & ~n13697 ;
  assign n45850 = n13722 & n45849 ;
  assign n45851 = ~n45848 & ~n45850 ;
  assign n45852 = n45846 & n45851 ;
  assign n45853 = n45841 & n45852 ;
  assign n45854 = \m3_addr_i[21]_pad  & ~n13697 ;
  assign n45855 = n13714 & n45854 ;
  assign n45856 = \m4_addr_i[21]_pad  & n13697 ;
  assign n45857 = n13722 & n45856 ;
  assign n45858 = ~n45855 & ~n45857 ;
  assign n45859 = \m6_addr_i[21]_pad  & n13697 ;
  assign n45860 = n13690 & n45859 ;
  assign n45861 = \m7_addr_i[21]_pad  & ~n13697 ;
  assign n45862 = n13690 & n45861 ;
  assign n45863 = ~n45860 & ~n45862 ;
  assign n45864 = n45858 & n45863 ;
  assign n45865 = \m5_addr_i[21]_pad  & ~n13697 ;
  assign n45866 = n13722 & n45865 ;
  assign n45867 = \m0_addr_i[21]_pad  & n13697 ;
  assign n45868 = n13705 & n45867 ;
  assign n45869 = ~n45866 & ~n45868 ;
  assign n45870 = \m1_addr_i[21]_pad  & ~n13697 ;
  assign n45871 = n13705 & n45870 ;
  assign n45872 = \m2_addr_i[21]_pad  & n13697 ;
  assign n45873 = n13714 & n45872 ;
  assign n45874 = ~n45871 & ~n45873 ;
  assign n45875 = n45869 & n45874 ;
  assign n45876 = n45864 & n45875 ;
  assign n45877 = \m1_addr_i[22]_pad  & ~n13697 ;
  assign n45878 = n13705 & n45877 ;
  assign n45879 = \m2_addr_i[22]_pad  & n13697 ;
  assign n45880 = n13714 & n45879 ;
  assign n45881 = ~n45878 & ~n45880 ;
  assign n45882 = \m3_addr_i[22]_pad  & ~n13697 ;
  assign n45883 = n13714 & n45882 ;
  assign n45884 = \m7_addr_i[22]_pad  & ~n13697 ;
  assign n45885 = n13690 & n45884 ;
  assign n45886 = ~n45883 & ~n45885 ;
  assign n45887 = n45881 & n45886 ;
  assign n45888 = \m4_addr_i[22]_pad  & n13697 ;
  assign n45889 = n13722 & n45888 ;
  assign n45890 = \m0_addr_i[22]_pad  & n13697 ;
  assign n45891 = n13705 & n45890 ;
  assign n45892 = ~n45889 & ~n45891 ;
  assign n45893 = \m6_addr_i[22]_pad  & n13697 ;
  assign n45894 = n13690 & n45893 ;
  assign n45895 = \m5_addr_i[22]_pad  & ~n13697 ;
  assign n45896 = n13722 & n45895 ;
  assign n45897 = ~n45894 & ~n45896 ;
  assign n45898 = n45892 & n45897 ;
  assign n45899 = n45887 & n45898 ;
  assign n45900 = \m1_addr_i[23]_pad  & ~n13697 ;
  assign n45901 = n13705 & n45900 ;
  assign n45902 = \m2_addr_i[23]_pad  & n13697 ;
  assign n45903 = n13714 & n45902 ;
  assign n45904 = ~n45901 & ~n45903 ;
  assign n45905 = \m3_addr_i[23]_pad  & ~n13697 ;
  assign n45906 = n13714 & n45905 ;
  assign n45907 = \m5_addr_i[23]_pad  & ~n13697 ;
  assign n45908 = n13722 & n45907 ;
  assign n45909 = ~n45906 & ~n45908 ;
  assign n45910 = n45904 & n45909 ;
  assign n45911 = \m4_addr_i[23]_pad  & n13697 ;
  assign n45912 = n13722 & n45911 ;
  assign n45913 = \m6_addr_i[23]_pad  & n13697 ;
  assign n45914 = n13690 & n45913 ;
  assign n45915 = ~n45912 & ~n45914 ;
  assign n45916 = \m0_addr_i[23]_pad  & n13697 ;
  assign n45917 = n13705 & n45916 ;
  assign n45918 = \m7_addr_i[23]_pad  & ~n13697 ;
  assign n45919 = n13690 & n45918 ;
  assign n45920 = ~n45917 & ~n45919 ;
  assign n45921 = n45915 & n45920 ;
  assign n45922 = n45910 & n45921 ;
  assign n45923 = \m1_addr_i[24]_pad  & ~n13697 ;
  assign n45924 = n13705 & n45923 ;
  assign n45925 = \m2_addr_i[24]_pad  & n13697 ;
  assign n45926 = n13714 & n45925 ;
  assign n45927 = ~n45924 & ~n45926 ;
  assign n45928 = \m5_addr_i[24]_pad  & ~n13697 ;
  assign n45929 = n13722 & n45928 ;
  assign n45930 = \m4_addr_i[24]_pad  & n13697 ;
  assign n45931 = n13722 & n45930 ;
  assign n45932 = ~n45929 & ~n45931 ;
  assign n45933 = n45927 & n45932 ;
  assign n45934 = \m6_addr_i[24]_pad  & n13697 ;
  assign n45935 = n13690 & n45934 ;
  assign n45936 = \m3_addr_i[24]_pad  & ~n13697 ;
  assign n45937 = n13714 & n45936 ;
  assign n45938 = ~n45935 & ~n45937 ;
  assign n45939 = \m0_addr_i[24]_pad  & n13697 ;
  assign n45940 = n13705 & n45939 ;
  assign n45941 = \m7_addr_i[24]_pad  & ~n13697 ;
  assign n45942 = n13690 & n45941 ;
  assign n45943 = ~n45940 & ~n45942 ;
  assign n45944 = n45938 & n45943 ;
  assign n45945 = n45933 & n45944 ;
  assign n45946 = \m3_addr_i[25]_pad  & ~n13697 ;
  assign n45947 = n13714 & n45946 ;
  assign n45948 = \m4_addr_i[25]_pad  & n13697 ;
  assign n45949 = n13722 & n45948 ;
  assign n45950 = ~n45947 & ~n45949 ;
  assign n45951 = \m5_addr_i[25]_pad  & ~n13697 ;
  assign n45952 = n13722 & n45951 ;
  assign n45953 = \m2_addr_i[25]_pad  & n13697 ;
  assign n45954 = n13714 & n45953 ;
  assign n45955 = ~n45952 & ~n45954 ;
  assign n45956 = n45950 & n45955 ;
  assign n45957 = \m6_addr_i[25]_pad  & n13697 ;
  assign n45958 = n13690 & n45957 ;
  assign n45959 = \m1_addr_i[25]_pad  & ~n13697 ;
  assign n45960 = n13705 & n45959 ;
  assign n45961 = ~n45958 & ~n45960 ;
  assign n45962 = \m0_addr_i[25]_pad  & n13697 ;
  assign n45963 = n13705 & n45962 ;
  assign n45964 = \m7_addr_i[25]_pad  & ~n13697 ;
  assign n45965 = n13690 & n45964 ;
  assign n45966 = ~n45963 & ~n45965 ;
  assign n45967 = n45961 & n45966 ;
  assign n45968 = n45956 & n45967 ;
  assign n45969 = \m1_addr_i[26]_pad  & ~n13697 ;
  assign n45970 = n13705 & n45969 ;
  assign n45971 = \m2_addr_i[26]_pad  & n13697 ;
  assign n45972 = n13714 & n45971 ;
  assign n45973 = ~n45970 & ~n45972 ;
  assign n45974 = \m3_addr_i[26]_pad  & ~n13697 ;
  assign n45975 = n13714 & n45974 ;
  assign n45976 = \m7_addr_i[26]_pad  & ~n13697 ;
  assign n45977 = n13690 & n45976 ;
  assign n45978 = ~n45975 & ~n45977 ;
  assign n45979 = n45973 & n45978 ;
  assign n45980 = \m4_addr_i[26]_pad  & n13697 ;
  assign n45981 = n13722 & n45980 ;
  assign n45982 = \m0_addr_i[26]_pad  & n13697 ;
  assign n45983 = n13705 & n45982 ;
  assign n45984 = ~n45981 & ~n45983 ;
  assign n45985 = \m5_addr_i[26]_pad  & ~n13697 ;
  assign n45986 = n13722 & n45985 ;
  assign n45987 = \m6_addr_i[26]_pad  & n13697 ;
  assign n45988 = n13690 & n45987 ;
  assign n45989 = ~n45986 & ~n45988 ;
  assign n45990 = n45984 & n45989 ;
  assign n45991 = n45979 & n45990 ;
  assign n45992 = \m3_addr_i[27]_pad  & ~n13697 ;
  assign n45993 = n13714 & n45992 ;
  assign n45994 = \m4_addr_i[27]_pad  & n13697 ;
  assign n45995 = n13722 & n45994 ;
  assign n45996 = ~n45993 & ~n45995 ;
  assign n45997 = \m5_addr_i[27]_pad  & ~n13697 ;
  assign n45998 = n13722 & n45997 ;
  assign n45999 = \m7_addr_i[27]_pad  & ~n13697 ;
  assign n46000 = n13690 & n45999 ;
  assign n46001 = ~n45998 & ~n46000 ;
  assign n46002 = n45996 & n46001 ;
  assign n46003 = \m6_addr_i[27]_pad  & n13697 ;
  assign n46004 = n13690 & n46003 ;
  assign n46005 = \m0_addr_i[27]_pad  & n13697 ;
  assign n46006 = n13705 & n46005 ;
  assign n46007 = ~n46004 & ~n46006 ;
  assign n46008 = \m1_addr_i[27]_pad  & ~n13697 ;
  assign n46009 = n13705 & n46008 ;
  assign n46010 = \m2_addr_i[27]_pad  & n13697 ;
  assign n46011 = n13714 & n46010 ;
  assign n46012 = ~n46009 & ~n46011 ;
  assign n46013 = n46007 & n46012 ;
  assign n46014 = n46002 & n46013 ;
  assign n46015 = \m1_addr_i[28]_pad  & ~n13697 ;
  assign n46016 = n13705 & n46015 ;
  assign n46017 = \m2_addr_i[28]_pad  & n13697 ;
  assign n46018 = n13714 & n46017 ;
  assign n46019 = ~n46016 & ~n46018 ;
  assign n46020 = \m5_addr_i[28]_pad  & ~n13697 ;
  assign n46021 = n13722 & n46020 ;
  assign n46022 = \m7_addr_i[28]_pad  & ~n13697 ;
  assign n46023 = n13690 & n46022 ;
  assign n46024 = ~n46021 & ~n46023 ;
  assign n46025 = n46019 & n46024 ;
  assign n46026 = \m6_addr_i[28]_pad  & n13697 ;
  assign n46027 = n13690 & n46026 ;
  assign n46028 = \m0_addr_i[28]_pad  & n13697 ;
  assign n46029 = n13705 & n46028 ;
  assign n46030 = ~n46027 & ~n46029 ;
  assign n46031 = \m3_addr_i[28]_pad  & ~n13697 ;
  assign n46032 = n13714 & n46031 ;
  assign n46033 = \m4_addr_i[28]_pad  & n13697 ;
  assign n46034 = n13722 & n46033 ;
  assign n46035 = ~n46032 & ~n46034 ;
  assign n46036 = n46030 & n46035 ;
  assign n46037 = n46025 & n46036 ;
  assign n46038 = \m0_addr_i[29]_pad  & n13697 ;
  assign n46039 = n13705 & n46038 ;
  assign n46040 = \m7_addr_i[29]_pad  & ~n13697 ;
  assign n46041 = n13690 & n46040 ;
  assign n46042 = ~n46039 & ~n46041 ;
  assign n46043 = \m1_addr_i[29]_pad  & ~n13697 ;
  assign n46044 = n13705 & n46043 ;
  assign n46045 = \m4_addr_i[29]_pad  & n13697 ;
  assign n46046 = n13722 & n46045 ;
  assign n46047 = ~n46044 & ~n46046 ;
  assign n46048 = n46042 & n46047 ;
  assign n46049 = \m2_addr_i[29]_pad  & n13697 ;
  assign n46050 = n13714 & n46049 ;
  assign n46051 = \m3_addr_i[29]_pad  & ~n13697 ;
  assign n46052 = n13714 & n46051 ;
  assign n46053 = ~n46050 & ~n46052 ;
  assign n46054 = \m5_addr_i[29]_pad  & ~n13697 ;
  assign n46055 = n13722 & n46054 ;
  assign n46056 = \m6_addr_i[29]_pad  & n13697 ;
  assign n46057 = n13690 & n46056 ;
  assign n46058 = ~n46055 & ~n46057 ;
  assign n46059 = n46053 & n46058 ;
  assign n46060 = n46048 & n46059 ;
  assign n46061 = \m3_addr_i[2]_pad  & ~n13697 ;
  assign n46062 = n13714 & n46061 ;
  assign n46063 = \m4_addr_i[2]_pad  & n13697 ;
  assign n46064 = n13722 & n46063 ;
  assign n46065 = ~n46062 & ~n46064 ;
  assign n46066 = \m6_addr_i[2]_pad  & n13697 ;
  assign n46067 = n13690 & n46066 ;
  assign n46068 = \m7_addr_i[2]_pad  & ~n13697 ;
  assign n46069 = n13690 & n46068 ;
  assign n46070 = ~n46067 & ~n46069 ;
  assign n46071 = n46065 & n46070 ;
  assign n46072 = \m5_addr_i[2]_pad  & ~n13697 ;
  assign n46073 = n13722 & n46072 ;
  assign n46074 = \m0_addr_i[2]_pad  & n13697 ;
  assign n46075 = n13705 & n46074 ;
  assign n46076 = ~n46073 & ~n46075 ;
  assign n46077 = \m1_addr_i[2]_pad  & ~n13697 ;
  assign n46078 = n13705 & n46077 ;
  assign n46079 = \m2_addr_i[2]_pad  & n13697 ;
  assign n46080 = n13714 & n46079 ;
  assign n46081 = ~n46078 & ~n46080 ;
  assign n46082 = n46076 & n46081 ;
  assign n46083 = n46071 & n46082 ;
  assign n46084 = \m1_addr_i[30]_pad  & ~n13697 ;
  assign n46085 = n13705 & n46084 ;
  assign n46086 = \m2_addr_i[30]_pad  & n13697 ;
  assign n46087 = n13714 & n46086 ;
  assign n46088 = ~n46085 & ~n46087 ;
  assign n46089 = \m3_addr_i[30]_pad  & ~n13697 ;
  assign n46090 = n13714 & n46089 ;
  assign n46091 = \m7_addr_i[30]_pad  & ~n13697 ;
  assign n46092 = n13690 & n46091 ;
  assign n46093 = ~n46090 & ~n46092 ;
  assign n46094 = n46088 & n46093 ;
  assign n46095 = \m4_addr_i[30]_pad  & n13697 ;
  assign n46096 = n13722 & n46095 ;
  assign n46097 = \m0_addr_i[30]_pad  & n13697 ;
  assign n46098 = n13705 & n46097 ;
  assign n46099 = ~n46096 & ~n46098 ;
  assign n46100 = \m5_addr_i[30]_pad  & ~n13697 ;
  assign n46101 = n13722 & n46100 ;
  assign n46102 = \m6_addr_i[30]_pad  & n13697 ;
  assign n46103 = n13690 & n46102 ;
  assign n46104 = ~n46101 & ~n46103 ;
  assign n46105 = n46099 & n46104 ;
  assign n46106 = n46094 & n46105 ;
  assign n46107 = \m3_addr_i[31]_pad  & ~n13697 ;
  assign n46108 = n13714 & n46107 ;
  assign n46109 = \m4_addr_i[31]_pad  & n13697 ;
  assign n46110 = n13722 & n46109 ;
  assign n46111 = ~n46108 & ~n46110 ;
  assign n46112 = \m5_addr_i[31]_pad  & ~n13697 ;
  assign n46113 = n13722 & n46112 ;
  assign n46114 = \m2_addr_i[31]_pad  & n13697 ;
  assign n46115 = n13714 & n46114 ;
  assign n46116 = ~n46113 & ~n46115 ;
  assign n46117 = n46111 & n46116 ;
  assign n46118 = \m6_addr_i[31]_pad  & n13697 ;
  assign n46119 = n13690 & n46118 ;
  assign n46120 = \m1_addr_i[31]_pad  & ~n13697 ;
  assign n46121 = n13705 & n46120 ;
  assign n46122 = ~n46119 & ~n46121 ;
  assign n46123 = \m0_addr_i[31]_pad  & n13697 ;
  assign n46124 = n13705 & n46123 ;
  assign n46125 = \m7_addr_i[31]_pad  & ~n13697 ;
  assign n46126 = n13690 & n46125 ;
  assign n46127 = ~n46124 & ~n46126 ;
  assign n46128 = n46122 & n46127 ;
  assign n46129 = n46117 & n46128 ;
  assign n46130 = \m3_addr_i[3]_pad  & ~n13697 ;
  assign n46131 = n13714 & n46130 ;
  assign n46132 = \m4_addr_i[3]_pad  & n13697 ;
  assign n46133 = n13722 & n46132 ;
  assign n46134 = ~n46131 & ~n46133 ;
  assign n46135 = \m6_addr_i[3]_pad  & n13697 ;
  assign n46136 = n13690 & n46135 ;
  assign n46137 = \m2_addr_i[3]_pad  & n13697 ;
  assign n46138 = n13714 & n46137 ;
  assign n46139 = ~n46136 & ~n46138 ;
  assign n46140 = n46134 & n46139 ;
  assign n46141 = \m5_addr_i[3]_pad  & ~n13697 ;
  assign n46142 = n13722 & n46141 ;
  assign n46143 = \m1_addr_i[3]_pad  & ~n13697 ;
  assign n46144 = n13705 & n46143 ;
  assign n46145 = ~n46142 & ~n46144 ;
  assign n46146 = \m0_addr_i[3]_pad  & n13697 ;
  assign n46147 = n13705 & n46146 ;
  assign n46148 = \m7_addr_i[3]_pad  & ~n13697 ;
  assign n46149 = n13690 & n46148 ;
  assign n46150 = ~n46147 & ~n46149 ;
  assign n46151 = n46145 & n46150 ;
  assign n46152 = n46140 & n46151 ;
  assign n46153 = \m3_addr_i[4]_pad  & ~n13697 ;
  assign n46154 = n13714 & n46153 ;
  assign n46155 = \m4_addr_i[4]_pad  & n13697 ;
  assign n46156 = n13722 & n46155 ;
  assign n46157 = ~n46154 & ~n46156 ;
  assign n46158 = \m6_addr_i[4]_pad  & n13697 ;
  assign n46159 = n13690 & n46158 ;
  assign n46160 = \m2_addr_i[4]_pad  & n13697 ;
  assign n46161 = n13714 & n46160 ;
  assign n46162 = ~n46159 & ~n46161 ;
  assign n46163 = n46157 & n46162 ;
  assign n46164 = \m5_addr_i[4]_pad  & ~n13697 ;
  assign n46165 = n13722 & n46164 ;
  assign n46166 = \m1_addr_i[4]_pad  & ~n13697 ;
  assign n46167 = n13705 & n46166 ;
  assign n46168 = ~n46165 & ~n46167 ;
  assign n46169 = \m0_addr_i[4]_pad  & n13697 ;
  assign n46170 = n13705 & n46169 ;
  assign n46171 = \m7_addr_i[4]_pad  & ~n13697 ;
  assign n46172 = n13690 & n46171 ;
  assign n46173 = ~n46170 & ~n46172 ;
  assign n46174 = n46168 & n46173 ;
  assign n46175 = n46163 & n46174 ;
  assign n46176 = \m3_addr_i[5]_pad  & ~n13697 ;
  assign n46177 = n13714 & n46176 ;
  assign n46178 = \m4_addr_i[5]_pad  & n13697 ;
  assign n46179 = n13722 & n46178 ;
  assign n46180 = ~n46177 & ~n46179 ;
  assign n46181 = \m6_addr_i[5]_pad  & n13697 ;
  assign n46182 = n13690 & n46181 ;
  assign n46183 = \m2_addr_i[5]_pad  & n13697 ;
  assign n46184 = n13714 & n46183 ;
  assign n46185 = ~n46182 & ~n46184 ;
  assign n46186 = n46180 & n46185 ;
  assign n46187 = \m5_addr_i[5]_pad  & ~n13697 ;
  assign n46188 = n13722 & n46187 ;
  assign n46189 = \m1_addr_i[5]_pad  & ~n13697 ;
  assign n46190 = n13705 & n46189 ;
  assign n46191 = ~n46188 & ~n46190 ;
  assign n46192 = \m0_addr_i[5]_pad  & n13697 ;
  assign n46193 = n13705 & n46192 ;
  assign n46194 = \m7_addr_i[5]_pad  & ~n13697 ;
  assign n46195 = n13690 & n46194 ;
  assign n46196 = ~n46193 & ~n46195 ;
  assign n46197 = n46191 & n46196 ;
  assign n46198 = n46186 & n46197 ;
  assign n46199 = \m1_addr_i[6]_pad  & ~n13697 ;
  assign n46200 = n13705 & n46199 ;
  assign n46201 = \m2_addr_i[6]_pad  & n13697 ;
  assign n46202 = n13714 & n46201 ;
  assign n46203 = ~n46200 & ~n46202 ;
  assign n46204 = \m6_addr_i[6]_pad  & n13697 ;
  assign n46205 = n13690 & n46204 ;
  assign n46206 = \m7_addr_i[6]_pad  & ~n13697 ;
  assign n46207 = n13690 & n46206 ;
  assign n46208 = ~n46205 & ~n46207 ;
  assign n46209 = n46203 & n46208 ;
  assign n46210 = \m5_addr_i[6]_pad  & ~n13697 ;
  assign n46211 = n13722 & n46210 ;
  assign n46212 = \m0_addr_i[6]_pad  & n13697 ;
  assign n46213 = n13705 & n46212 ;
  assign n46214 = ~n46211 & ~n46213 ;
  assign n46215 = \m3_addr_i[6]_pad  & ~n13697 ;
  assign n46216 = n13714 & n46215 ;
  assign n46217 = \m4_addr_i[6]_pad  & n13697 ;
  assign n46218 = n13722 & n46217 ;
  assign n46219 = ~n46216 & ~n46218 ;
  assign n46220 = n46214 & n46219 ;
  assign n46221 = n46209 & n46220 ;
  assign n46222 = \m1_addr_i[7]_pad  & ~n13697 ;
  assign n46223 = n13705 & n46222 ;
  assign n46224 = \m2_addr_i[7]_pad  & n13697 ;
  assign n46225 = n13714 & n46224 ;
  assign n46226 = ~n46223 & ~n46225 ;
  assign n46227 = \m6_addr_i[7]_pad  & n13697 ;
  assign n46228 = n13690 & n46227 ;
  assign n46229 = \m4_addr_i[7]_pad  & n13697 ;
  assign n46230 = n13722 & n46229 ;
  assign n46231 = ~n46228 & ~n46230 ;
  assign n46232 = n46226 & n46231 ;
  assign n46233 = \m5_addr_i[7]_pad  & ~n13697 ;
  assign n46234 = n13722 & n46233 ;
  assign n46235 = \m3_addr_i[7]_pad  & ~n13697 ;
  assign n46236 = n13714 & n46235 ;
  assign n46237 = ~n46234 & ~n46236 ;
  assign n46238 = \m0_addr_i[7]_pad  & n13697 ;
  assign n46239 = n13705 & n46238 ;
  assign n46240 = \m7_addr_i[7]_pad  & ~n13697 ;
  assign n46241 = n13690 & n46240 ;
  assign n46242 = ~n46239 & ~n46241 ;
  assign n46243 = n46237 & n46242 ;
  assign n46244 = n46232 & n46243 ;
  assign n46245 = \m3_addr_i[8]_pad  & ~n13697 ;
  assign n46246 = n13714 & n46245 ;
  assign n46247 = \m4_addr_i[8]_pad  & n13697 ;
  assign n46248 = n13722 & n46247 ;
  assign n46249 = ~n46246 & ~n46248 ;
  assign n46250 = \m6_addr_i[8]_pad  & n13697 ;
  assign n46251 = n13690 & n46250 ;
  assign n46252 = \m2_addr_i[8]_pad  & n13697 ;
  assign n46253 = n13714 & n46252 ;
  assign n46254 = ~n46251 & ~n46253 ;
  assign n46255 = n46249 & n46254 ;
  assign n46256 = \m5_addr_i[8]_pad  & ~n13697 ;
  assign n46257 = n13722 & n46256 ;
  assign n46258 = \m1_addr_i[8]_pad  & ~n13697 ;
  assign n46259 = n13705 & n46258 ;
  assign n46260 = ~n46257 & ~n46259 ;
  assign n46261 = \m0_addr_i[8]_pad  & n13697 ;
  assign n46262 = n13705 & n46261 ;
  assign n46263 = \m7_addr_i[8]_pad  & ~n13697 ;
  assign n46264 = n13690 & n46263 ;
  assign n46265 = ~n46262 & ~n46264 ;
  assign n46266 = n46260 & n46265 ;
  assign n46267 = n46255 & n46266 ;
  assign n46268 = \m1_addr_i[9]_pad  & ~n13697 ;
  assign n46269 = n13705 & n46268 ;
  assign n46270 = \m2_addr_i[9]_pad  & n13697 ;
  assign n46271 = n13714 & n46270 ;
  assign n46272 = ~n46269 & ~n46271 ;
  assign n46273 = \m6_addr_i[9]_pad  & n13697 ;
  assign n46274 = n13690 & n46273 ;
  assign n46275 = \m7_addr_i[9]_pad  & ~n13697 ;
  assign n46276 = n13690 & n46275 ;
  assign n46277 = ~n46274 & ~n46276 ;
  assign n46278 = n46272 & n46277 ;
  assign n46279 = \m5_addr_i[9]_pad  & ~n13697 ;
  assign n46280 = n13722 & n46279 ;
  assign n46281 = \m0_addr_i[9]_pad  & n13697 ;
  assign n46282 = n13705 & n46281 ;
  assign n46283 = ~n46280 & ~n46282 ;
  assign n46284 = \m3_addr_i[9]_pad  & ~n13697 ;
  assign n46285 = n13714 & n46284 ;
  assign n46286 = \m4_addr_i[9]_pad  & n13697 ;
  assign n46287 = n13722 & n46286 ;
  assign n46288 = ~n46285 & ~n46287 ;
  assign n46289 = n46283 & n46288 ;
  assign n46290 = n46278 & n46289 ;
  assign n46291 = \m3_data_i[0]_pad  & ~n13697 ;
  assign n46292 = n13714 & n46291 ;
  assign n46293 = \m4_data_i[0]_pad  & n13697 ;
  assign n46294 = n13722 & n46293 ;
  assign n46295 = ~n46292 & ~n46294 ;
  assign n46296 = \m6_data_i[0]_pad  & n13697 ;
  assign n46297 = n13690 & n46296 ;
  assign n46298 = \m2_data_i[0]_pad  & n13697 ;
  assign n46299 = n13714 & n46298 ;
  assign n46300 = ~n46297 & ~n46299 ;
  assign n46301 = n46295 & n46300 ;
  assign n46302 = \m5_data_i[0]_pad  & ~n13697 ;
  assign n46303 = n13722 & n46302 ;
  assign n46304 = \m1_data_i[0]_pad  & ~n13697 ;
  assign n46305 = n13705 & n46304 ;
  assign n46306 = ~n46303 & ~n46305 ;
  assign n46307 = \m0_data_i[0]_pad  & n13697 ;
  assign n46308 = n13705 & n46307 ;
  assign n46309 = \m7_data_i[0]_pad  & ~n13697 ;
  assign n46310 = n13690 & n46309 ;
  assign n46311 = ~n46308 & ~n46310 ;
  assign n46312 = n46306 & n46311 ;
  assign n46313 = n46301 & n46312 ;
  assign n46314 = \m1_data_i[10]_pad  & ~n13697 ;
  assign n46315 = n13705 & n46314 ;
  assign n46316 = \m2_data_i[10]_pad  & n13697 ;
  assign n46317 = n13714 & n46316 ;
  assign n46318 = ~n46315 & ~n46317 ;
  assign n46319 = \m3_data_i[10]_pad  & ~n13697 ;
  assign n46320 = n13714 & n46319 ;
  assign n46321 = \m5_data_i[10]_pad  & ~n13697 ;
  assign n46322 = n13722 & n46321 ;
  assign n46323 = ~n46320 & ~n46322 ;
  assign n46324 = n46318 & n46323 ;
  assign n46325 = \m4_data_i[10]_pad  & n13697 ;
  assign n46326 = n13722 & n46325 ;
  assign n46327 = \m6_data_i[10]_pad  & n13697 ;
  assign n46328 = n13690 & n46327 ;
  assign n46329 = ~n46326 & ~n46328 ;
  assign n46330 = \m0_data_i[10]_pad  & n13697 ;
  assign n46331 = n13705 & n46330 ;
  assign n46332 = \m7_data_i[10]_pad  & ~n13697 ;
  assign n46333 = n13690 & n46332 ;
  assign n46334 = ~n46331 & ~n46333 ;
  assign n46335 = n46329 & n46334 ;
  assign n46336 = n46324 & n46335 ;
  assign n46337 = \m6_data_i[11]_pad  & n13697 ;
  assign n46338 = n13690 & n46337 ;
  assign n46339 = \m5_data_i[11]_pad  & ~n13697 ;
  assign n46340 = n13722 & n46339 ;
  assign n46341 = ~n46338 & ~n46340 ;
  assign n46342 = \m3_data_i[11]_pad  & ~n13697 ;
  assign n46343 = n13714 & n46342 ;
  assign n46344 = \m2_data_i[11]_pad  & n13697 ;
  assign n46345 = n13714 & n46344 ;
  assign n46346 = ~n46343 & ~n46345 ;
  assign n46347 = n46341 & n46346 ;
  assign n46348 = \m4_data_i[11]_pad  & n13697 ;
  assign n46349 = n13722 & n46348 ;
  assign n46350 = \m1_data_i[11]_pad  & ~n13697 ;
  assign n46351 = n13705 & n46350 ;
  assign n46352 = ~n46349 & ~n46351 ;
  assign n46353 = \m0_data_i[11]_pad  & n13697 ;
  assign n46354 = n13705 & n46353 ;
  assign n46355 = \m7_data_i[11]_pad  & ~n13697 ;
  assign n46356 = n13690 & n46355 ;
  assign n46357 = ~n46354 & ~n46356 ;
  assign n46358 = n46352 & n46357 ;
  assign n46359 = n46347 & n46358 ;
  assign n46360 = \m1_data_i[12]_pad  & ~n13697 ;
  assign n46361 = n13705 & n46360 ;
  assign n46362 = \m2_data_i[12]_pad  & n13697 ;
  assign n46363 = n13714 & n46362 ;
  assign n46364 = ~n46361 & ~n46363 ;
  assign n46365 = \m0_data_i[12]_pad  & n13697 ;
  assign n46366 = n13705 & n46365 ;
  assign n46367 = \m4_data_i[12]_pad  & n13697 ;
  assign n46368 = n13722 & n46367 ;
  assign n46369 = ~n46366 & ~n46368 ;
  assign n46370 = n46364 & n46369 ;
  assign n46371 = \m7_data_i[12]_pad  & ~n13697 ;
  assign n46372 = n13690 & n46371 ;
  assign n46373 = \m3_data_i[12]_pad  & ~n13697 ;
  assign n46374 = n13714 & n46373 ;
  assign n46375 = ~n46372 & ~n46374 ;
  assign n46376 = \m6_data_i[12]_pad  & n13697 ;
  assign n46377 = n13690 & n46376 ;
  assign n46378 = \m5_data_i[12]_pad  & ~n13697 ;
  assign n46379 = n13722 & n46378 ;
  assign n46380 = ~n46377 & ~n46379 ;
  assign n46381 = n46375 & n46380 ;
  assign n46382 = n46370 & n46381 ;
  assign n46383 = \m1_data_i[13]_pad  & ~n13697 ;
  assign n46384 = n13705 & n46383 ;
  assign n46385 = \m2_data_i[13]_pad  & n13697 ;
  assign n46386 = n13714 & n46385 ;
  assign n46387 = ~n46384 & ~n46386 ;
  assign n46388 = \m0_data_i[13]_pad  & n13697 ;
  assign n46389 = n13705 & n46388 ;
  assign n46390 = \m4_data_i[13]_pad  & n13697 ;
  assign n46391 = n13722 & n46390 ;
  assign n46392 = ~n46389 & ~n46391 ;
  assign n46393 = n46387 & n46392 ;
  assign n46394 = \m7_data_i[13]_pad  & ~n13697 ;
  assign n46395 = n13690 & n46394 ;
  assign n46396 = \m3_data_i[13]_pad  & ~n13697 ;
  assign n46397 = n13714 & n46396 ;
  assign n46398 = ~n46395 & ~n46397 ;
  assign n46399 = \m6_data_i[13]_pad  & n13697 ;
  assign n46400 = n13690 & n46399 ;
  assign n46401 = \m5_data_i[13]_pad  & ~n13697 ;
  assign n46402 = n13722 & n46401 ;
  assign n46403 = ~n46400 & ~n46402 ;
  assign n46404 = n46398 & n46403 ;
  assign n46405 = n46393 & n46404 ;
  assign n46406 = \m1_data_i[14]_pad  & ~n13697 ;
  assign n46407 = n13705 & n46406 ;
  assign n46408 = \m2_data_i[14]_pad  & n13697 ;
  assign n46409 = n13714 & n46408 ;
  assign n46410 = ~n46407 & ~n46409 ;
  assign n46411 = \m0_data_i[14]_pad  & n13697 ;
  assign n46412 = n13705 & n46411 ;
  assign n46413 = \m4_data_i[14]_pad  & n13697 ;
  assign n46414 = n13722 & n46413 ;
  assign n46415 = ~n46412 & ~n46414 ;
  assign n46416 = n46410 & n46415 ;
  assign n46417 = \m7_data_i[14]_pad  & ~n13697 ;
  assign n46418 = n13690 & n46417 ;
  assign n46419 = \m3_data_i[14]_pad  & ~n13697 ;
  assign n46420 = n13714 & n46419 ;
  assign n46421 = ~n46418 & ~n46420 ;
  assign n46422 = \m6_data_i[14]_pad  & n13697 ;
  assign n46423 = n13690 & n46422 ;
  assign n46424 = \m5_data_i[14]_pad  & ~n13697 ;
  assign n46425 = n13722 & n46424 ;
  assign n46426 = ~n46423 & ~n46425 ;
  assign n46427 = n46421 & n46426 ;
  assign n46428 = n46416 & n46427 ;
  assign n46429 = \m1_data_i[15]_pad  & ~n13697 ;
  assign n46430 = n13705 & n46429 ;
  assign n46431 = \m2_data_i[15]_pad  & n13697 ;
  assign n46432 = n13714 & n46431 ;
  assign n46433 = ~n46430 & ~n46432 ;
  assign n46434 = \m0_data_i[15]_pad  & n13697 ;
  assign n46435 = n13705 & n46434 ;
  assign n46436 = \m4_data_i[15]_pad  & n13697 ;
  assign n46437 = n13722 & n46436 ;
  assign n46438 = ~n46435 & ~n46437 ;
  assign n46439 = n46433 & n46438 ;
  assign n46440 = \m7_data_i[15]_pad  & ~n13697 ;
  assign n46441 = n13690 & n46440 ;
  assign n46442 = \m3_data_i[15]_pad  & ~n13697 ;
  assign n46443 = n13714 & n46442 ;
  assign n46444 = ~n46441 & ~n46443 ;
  assign n46445 = \m6_data_i[15]_pad  & n13697 ;
  assign n46446 = n13690 & n46445 ;
  assign n46447 = \m5_data_i[15]_pad  & ~n13697 ;
  assign n46448 = n13722 & n46447 ;
  assign n46449 = ~n46446 & ~n46448 ;
  assign n46450 = n46444 & n46449 ;
  assign n46451 = n46439 & n46450 ;
  assign n46452 = \m3_data_i[16]_pad  & ~n13697 ;
  assign n46453 = n13714 & n46452 ;
  assign n46454 = \m4_data_i[16]_pad  & n13697 ;
  assign n46455 = n13722 & n46454 ;
  assign n46456 = ~n46453 & ~n46455 ;
  assign n46457 = \m0_data_i[16]_pad  & n13697 ;
  assign n46458 = n13705 & n46457 ;
  assign n46459 = \m5_data_i[16]_pad  & ~n13697 ;
  assign n46460 = n13722 & n46459 ;
  assign n46461 = ~n46458 & ~n46460 ;
  assign n46462 = n46456 & n46461 ;
  assign n46463 = \m7_data_i[16]_pad  & ~n13697 ;
  assign n46464 = n13690 & n46463 ;
  assign n46465 = \m6_data_i[16]_pad  & n13697 ;
  assign n46466 = n13690 & n46465 ;
  assign n46467 = ~n46464 & ~n46466 ;
  assign n46468 = \m1_data_i[16]_pad  & ~n13697 ;
  assign n46469 = n13705 & n46468 ;
  assign n46470 = \m2_data_i[16]_pad  & n13697 ;
  assign n46471 = n13714 & n46470 ;
  assign n46472 = ~n46469 & ~n46471 ;
  assign n46473 = n46467 & n46472 ;
  assign n46474 = n46462 & n46473 ;
  assign n46475 = \m1_data_i[17]_pad  & ~n13697 ;
  assign n46476 = n13705 & n46475 ;
  assign n46477 = \m2_data_i[17]_pad  & n13697 ;
  assign n46478 = n13714 & n46477 ;
  assign n46479 = ~n46476 & ~n46478 ;
  assign n46480 = \m6_data_i[17]_pad  & n13697 ;
  assign n46481 = n13690 & n46480 ;
  assign n46482 = \m7_data_i[17]_pad  & ~n13697 ;
  assign n46483 = n13690 & n46482 ;
  assign n46484 = ~n46481 & ~n46483 ;
  assign n46485 = n46479 & n46484 ;
  assign n46486 = \m5_data_i[17]_pad  & ~n13697 ;
  assign n46487 = n13722 & n46486 ;
  assign n46488 = \m0_data_i[17]_pad  & n13697 ;
  assign n46489 = n13705 & n46488 ;
  assign n46490 = ~n46487 & ~n46489 ;
  assign n46491 = \m3_data_i[17]_pad  & ~n13697 ;
  assign n46492 = n13714 & n46491 ;
  assign n46493 = \m4_data_i[17]_pad  & n13697 ;
  assign n46494 = n13722 & n46493 ;
  assign n46495 = ~n46492 & ~n46494 ;
  assign n46496 = n46490 & n46495 ;
  assign n46497 = n46485 & n46496 ;
  assign n46498 = \m3_data_i[18]_pad  & ~n13697 ;
  assign n46499 = n13714 & n46498 ;
  assign n46500 = \m4_data_i[18]_pad  & n13697 ;
  assign n46501 = n13722 & n46500 ;
  assign n46502 = ~n46499 & ~n46501 ;
  assign n46503 = \m6_data_i[18]_pad  & n13697 ;
  assign n46504 = n13690 & n46503 ;
  assign n46505 = \m2_data_i[18]_pad  & n13697 ;
  assign n46506 = n13714 & n46505 ;
  assign n46507 = ~n46504 & ~n46506 ;
  assign n46508 = n46502 & n46507 ;
  assign n46509 = \m5_data_i[18]_pad  & ~n13697 ;
  assign n46510 = n13722 & n46509 ;
  assign n46511 = \m1_data_i[18]_pad  & ~n13697 ;
  assign n46512 = n13705 & n46511 ;
  assign n46513 = ~n46510 & ~n46512 ;
  assign n46514 = \m0_data_i[18]_pad  & n13697 ;
  assign n46515 = n13705 & n46514 ;
  assign n46516 = \m7_data_i[18]_pad  & ~n13697 ;
  assign n46517 = n13690 & n46516 ;
  assign n46518 = ~n46515 & ~n46517 ;
  assign n46519 = n46513 & n46518 ;
  assign n46520 = n46508 & n46519 ;
  assign n46521 = \m1_data_i[19]_pad  & ~n13697 ;
  assign n46522 = n13705 & n46521 ;
  assign n46523 = \m2_data_i[19]_pad  & n13697 ;
  assign n46524 = n13714 & n46523 ;
  assign n46525 = ~n46522 & ~n46524 ;
  assign n46526 = \m3_data_i[19]_pad  & ~n13697 ;
  assign n46527 = n13714 & n46526 ;
  assign n46528 = \m7_data_i[19]_pad  & ~n13697 ;
  assign n46529 = n13690 & n46528 ;
  assign n46530 = ~n46527 & ~n46529 ;
  assign n46531 = n46525 & n46530 ;
  assign n46532 = \m4_data_i[19]_pad  & n13697 ;
  assign n46533 = n13722 & n46532 ;
  assign n46534 = \m0_data_i[19]_pad  & n13697 ;
  assign n46535 = n13705 & n46534 ;
  assign n46536 = ~n46533 & ~n46535 ;
  assign n46537 = \m6_data_i[19]_pad  & n13697 ;
  assign n46538 = n13690 & n46537 ;
  assign n46539 = \m5_data_i[19]_pad  & ~n13697 ;
  assign n46540 = n13722 & n46539 ;
  assign n46541 = ~n46538 & ~n46540 ;
  assign n46542 = n46536 & n46541 ;
  assign n46543 = n46531 & n46542 ;
  assign n46544 = \m0_data_i[1]_pad  & n13697 ;
  assign n46545 = n13705 & n46544 ;
  assign n46546 = \m7_data_i[1]_pad  & ~n13697 ;
  assign n46547 = n13690 & n46546 ;
  assign n46548 = ~n46545 & ~n46547 ;
  assign n46549 = \m1_data_i[1]_pad  & ~n13697 ;
  assign n46550 = n13705 & n46549 ;
  assign n46551 = \m4_data_i[1]_pad  & n13697 ;
  assign n46552 = n13722 & n46551 ;
  assign n46553 = ~n46550 & ~n46552 ;
  assign n46554 = n46548 & n46553 ;
  assign n46555 = \m2_data_i[1]_pad  & n13697 ;
  assign n46556 = n13714 & n46555 ;
  assign n46557 = \m3_data_i[1]_pad  & ~n13697 ;
  assign n46558 = n13714 & n46557 ;
  assign n46559 = ~n46556 & ~n46558 ;
  assign n46560 = \m6_data_i[1]_pad  & n13697 ;
  assign n46561 = n13690 & n46560 ;
  assign n46562 = \m5_data_i[1]_pad  & ~n13697 ;
  assign n46563 = n13722 & n46562 ;
  assign n46564 = ~n46561 & ~n46563 ;
  assign n46565 = n46559 & n46564 ;
  assign n46566 = n46554 & n46565 ;
  assign n46567 = \m1_data_i[20]_pad  & ~n13697 ;
  assign n46568 = n13705 & n46567 ;
  assign n46569 = \m2_data_i[20]_pad  & n13697 ;
  assign n46570 = n13714 & n46569 ;
  assign n46571 = ~n46568 & ~n46570 ;
  assign n46572 = \m0_data_i[20]_pad  & n13697 ;
  assign n46573 = n13705 & n46572 ;
  assign n46574 = \m4_data_i[20]_pad  & n13697 ;
  assign n46575 = n13722 & n46574 ;
  assign n46576 = ~n46573 & ~n46575 ;
  assign n46577 = n46571 & n46576 ;
  assign n46578 = \m7_data_i[20]_pad  & ~n13697 ;
  assign n46579 = n13690 & n46578 ;
  assign n46580 = \m3_data_i[20]_pad  & ~n13697 ;
  assign n46581 = n13714 & n46580 ;
  assign n46582 = ~n46579 & ~n46581 ;
  assign n46583 = \m6_data_i[20]_pad  & n13697 ;
  assign n46584 = n13690 & n46583 ;
  assign n46585 = \m5_data_i[20]_pad  & ~n13697 ;
  assign n46586 = n13722 & n46585 ;
  assign n46587 = ~n46584 & ~n46586 ;
  assign n46588 = n46582 & n46587 ;
  assign n46589 = n46577 & n46588 ;
  assign n46590 = \m6_data_i[21]_pad  & n13697 ;
  assign n46591 = n13690 & n46590 ;
  assign n46592 = \m5_data_i[21]_pad  & ~n13697 ;
  assign n46593 = n13722 & n46592 ;
  assign n46594 = ~n46591 & ~n46593 ;
  assign n46595 = \m1_data_i[21]_pad  & ~n13697 ;
  assign n46596 = n13705 & n46595 ;
  assign n46597 = \m4_data_i[21]_pad  & n13697 ;
  assign n46598 = n13722 & n46597 ;
  assign n46599 = ~n46596 & ~n46598 ;
  assign n46600 = n46594 & n46599 ;
  assign n46601 = \m2_data_i[21]_pad  & n13697 ;
  assign n46602 = n13714 & n46601 ;
  assign n46603 = \m3_data_i[21]_pad  & ~n13697 ;
  assign n46604 = n13714 & n46603 ;
  assign n46605 = ~n46602 & ~n46604 ;
  assign n46606 = \m0_data_i[21]_pad  & n13697 ;
  assign n46607 = n13705 & n46606 ;
  assign n46608 = \m7_data_i[21]_pad  & ~n13697 ;
  assign n46609 = n13690 & n46608 ;
  assign n46610 = ~n46607 & ~n46609 ;
  assign n46611 = n46605 & n46610 ;
  assign n46612 = n46600 & n46611 ;
  assign n46613 = \m3_data_i[22]_pad  & ~n13697 ;
  assign n46614 = n13714 & n46613 ;
  assign n46615 = \m4_data_i[22]_pad  & n13697 ;
  assign n46616 = n13722 & n46615 ;
  assign n46617 = ~n46614 & ~n46616 ;
  assign n46618 = \m6_data_i[22]_pad  & n13697 ;
  assign n46619 = n13690 & n46618 ;
  assign n46620 = \m2_data_i[22]_pad  & n13697 ;
  assign n46621 = n13714 & n46620 ;
  assign n46622 = ~n46619 & ~n46621 ;
  assign n46623 = n46617 & n46622 ;
  assign n46624 = \m5_data_i[22]_pad  & ~n13697 ;
  assign n46625 = n13722 & n46624 ;
  assign n46626 = \m1_data_i[22]_pad  & ~n13697 ;
  assign n46627 = n13705 & n46626 ;
  assign n46628 = ~n46625 & ~n46627 ;
  assign n46629 = \m0_data_i[22]_pad  & n13697 ;
  assign n46630 = n13705 & n46629 ;
  assign n46631 = \m7_data_i[22]_pad  & ~n13697 ;
  assign n46632 = n13690 & n46631 ;
  assign n46633 = ~n46630 & ~n46632 ;
  assign n46634 = n46628 & n46633 ;
  assign n46635 = n46623 & n46634 ;
  assign n46636 = \m6_data_i[23]_pad  & n13697 ;
  assign n46637 = n13690 & n46636 ;
  assign n46638 = \m5_data_i[23]_pad  & ~n13697 ;
  assign n46639 = n13722 & n46638 ;
  assign n46640 = ~n46637 & ~n46639 ;
  assign n46641 = \m1_data_i[23]_pad  & ~n13697 ;
  assign n46642 = n13705 & n46641 ;
  assign n46643 = \m4_data_i[23]_pad  & n13697 ;
  assign n46644 = n13722 & n46643 ;
  assign n46645 = ~n46642 & ~n46644 ;
  assign n46646 = n46640 & n46645 ;
  assign n46647 = \m2_data_i[23]_pad  & n13697 ;
  assign n46648 = n13714 & n46647 ;
  assign n46649 = \m3_data_i[23]_pad  & ~n13697 ;
  assign n46650 = n13714 & n46649 ;
  assign n46651 = ~n46648 & ~n46650 ;
  assign n46652 = \m0_data_i[23]_pad  & n13697 ;
  assign n46653 = n13705 & n46652 ;
  assign n46654 = \m7_data_i[23]_pad  & ~n13697 ;
  assign n46655 = n13690 & n46654 ;
  assign n46656 = ~n46653 & ~n46655 ;
  assign n46657 = n46651 & n46656 ;
  assign n46658 = n46646 & n46657 ;
  assign n46659 = \m1_data_i[24]_pad  & ~n13697 ;
  assign n46660 = n13705 & n46659 ;
  assign n46661 = \m2_data_i[24]_pad  & n13697 ;
  assign n46662 = n13714 & n46661 ;
  assign n46663 = ~n46660 & ~n46662 ;
  assign n46664 = \m0_data_i[24]_pad  & n13697 ;
  assign n46665 = n13705 & n46664 ;
  assign n46666 = \m4_data_i[24]_pad  & n13697 ;
  assign n46667 = n13722 & n46666 ;
  assign n46668 = ~n46665 & ~n46667 ;
  assign n46669 = n46663 & n46668 ;
  assign n46670 = \m7_data_i[24]_pad  & ~n13697 ;
  assign n46671 = n13690 & n46670 ;
  assign n46672 = \m3_data_i[24]_pad  & ~n13697 ;
  assign n46673 = n13714 & n46672 ;
  assign n46674 = ~n46671 & ~n46673 ;
  assign n46675 = \m6_data_i[24]_pad  & n13697 ;
  assign n46676 = n13690 & n46675 ;
  assign n46677 = \m5_data_i[24]_pad  & ~n13697 ;
  assign n46678 = n13722 & n46677 ;
  assign n46679 = ~n46676 & ~n46678 ;
  assign n46680 = n46674 & n46679 ;
  assign n46681 = n46669 & n46680 ;
  assign n46682 = \m1_data_i[25]_pad  & ~n13697 ;
  assign n46683 = n13705 & n46682 ;
  assign n46684 = \m2_data_i[25]_pad  & n13697 ;
  assign n46685 = n13714 & n46684 ;
  assign n46686 = ~n46683 & ~n46685 ;
  assign n46687 = \m0_data_i[25]_pad  & n13697 ;
  assign n46688 = n13705 & n46687 ;
  assign n46689 = \m4_data_i[25]_pad  & n13697 ;
  assign n46690 = n13722 & n46689 ;
  assign n46691 = ~n46688 & ~n46690 ;
  assign n46692 = n46686 & n46691 ;
  assign n46693 = \m7_data_i[25]_pad  & ~n13697 ;
  assign n46694 = n13690 & n46693 ;
  assign n46695 = \m3_data_i[25]_pad  & ~n13697 ;
  assign n46696 = n13714 & n46695 ;
  assign n46697 = ~n46694 & ~n46696 ;
  assign n46698 = \m6_data_i[25]_pad  & n13697 ;
  assign n46699 = n13690 & n46698 ;
  assign n46700 = \m5_data_i[25]_pad  & ~n13697 ;
  assign n46701 = n13722 & n46700 ;
  assign n46702 = ~n46699 & ~n46701 ;
  assign n46703 = n46697 & n46702 ;
  assign n46704 = n46692 & n46703 ;
  assign n46705 = \m1_data_i[26]_pad  & ~n13697 ;
  assign n46706 = n13705 & n46705 ;
  assign n46707 = \m2_data_i[26]_pad  & n13697 ;
  assign n46708 = n13714 & n46707 ;
  assign n46709 = ~n46706 & ~n46708 ;
  assign n46710 = \m6_data_i[26]_pad  & n13697 ;
  assign n46711 = n13690 & n46710 ;
  assign n46712 = \m7_data_i[26]_pad  & ~n13697 ;
  assign n46713 = n13690 & n46712 ;
  assign n46714 = ~n46711 & ~n46713 ;
  assign n46715 = n46709 & n46714 ;
  assign n46716 = \m5_data_i[26]_pad  & ~n13697 ;
  assign n46717 = n13722 & n46716 ;
  assign n46718 = \m0_data_i[26]_pad  & n13697 ;
  assign n46719 = n13705 & n46718 ;
  assign n46720 = ~n46717 & ~n46719 ;
  assign n46721 = \m3_data_i[26]_pad  & ~n13697 ;
  assign n46722 = n13714 & n46721 ;
  assign n46723 = \m4_data_i[26]_pad  & n13697 ;
  assign n46724 = n13722 & n46723 ;
  assign n46725 = ~n46722 & ~n46724 ;
  assign n46726 = n46720 & n46725 ;
  assign n46727 = n46715 & n46726 ;
  assign n46728 = \m1_data_i[27]_pad  & ~n13697 ;
  assign n46729 = n13705 & n46728 ;
  assign n46730 = \m2_data_i[27]_pad  & n13697 ;
  assign n46731 = n13714 & n46730 ;
  assign n46732 = ~n46729 & ~n46731 ;
  assign n46733 = \m6_data_i[27]_pad  & n13697 ;
  assign n46734 = n13690 & n46733 ;
  assign n46735 = \m7_data_i[27]_pad  & ~n13697 ;
  assign n46736 = n13690 & n46735 ;
  assign n46737 = ~n46734 & ~n46736 ;
  assign n46738 = n46732 & n46737 ;
  assign n46739 = \m5_data_i[27]_pad  & ~n13697 ;
  assign n46740 = n13722 & n46739 ;
  assign n46741 = \m0_data_i[27]_pad  & n13697 ;
  assign n46742 = n13705 & n46741 ;
  assign n46743 = ~n46740 & ~n46742 ;
  assign n46744 = \m3_data_i[27]_pad  & ~n13697 ;
  assign n46745 = n13714 & n46744 ;
  assign n46746 = \m4_data_i[27]_pad  & n13697 ;
  assign n46747 = n13722 & n46746 ;
  assign n46748 = ~n46745 & ~n46747 ;
  assign n46749 = n46743 & n46748 ;
  assign n46750 = n46738 & n46749 ;
  assign n46751 = \m3_data_i[28]_pad  & ~n13697 ;
  assign n46752 = n13714 & n46751 ;
  assign n46753 = \m4_data_i[28]_pad  & n13697 ;
  assign n46754 = n13722 & n46753 ;
  assign n46755 = ~n46752 & ~n46754 ;
  assign n46756 = \m6_data_i[28]_pad  & n13697 ;
  assign n46757 = n13690 & n46756 ;
  assign n46758 = \m7_data_i[28]_pad  & ~n13697 ;
  assign n46759 = n13690 & n46758 ;
  assign n46760 = ~n46757 & ~n46759 ;
  assign n46761 = n46755 & n46760 ;
  assign n46762 = \m5_data_i[28]_pad  & ~n13697 ;
  assign n46763 = n13722 & n46762 ;
  assign n46764 = \m0_data_i[28]_pad  & n13697 ;
  assign n46765 = n13705 & n46764 ;
  assign n46766 = ~n46763 & ~n46765 ;
  assign n46767 = \m1_data_i[28]_pad  & ~n13697 ;
  assign n46768 = n13705 & n46767 ;
  assign n46769 = \m2_data_i[28]_pad  & n13697 ;
  assign n46770 = n13714 & n46769 ;
  assign n46771 = ~n46768 & ~n46770 ;
  assign n46772 = n46766 & n46771 ;
  assign n46773 = n46761 & n46772 ;
  assign n46774 = \m1_data_i[29]_pad  & ~n13697 ;
  assign n46775 = n13705 & n46774 ;
  assign n46776 = \m2_data_i[29]_pad  & n13697 ;
  assign n46777 = n13714 & n46776 ;
  assign n46778 = ~n46775 & ~n46777 ;
  assign n46779 = \m3_data_i[29]_pad  & ~n13697 ;
  assign n46780 = n13714 & n46779 ;
  assign n46781 = \m7_data_i[29]_pad  & ~n13697 ;
  assign n46782 = n13690 & n46781 ;
  assign n46783 = ~n46780 & ~n46782 ;
  assign n46784 = n46778 & n46783 ;
  assign n46785 = \m4_data_i[29]_pad  & n13697 ;
  assign n46786 = n13722 & n46785 ;
  assign n46787 = \m0_data_i[29]_pad  & n13697 ;
  assign n46788 = n13705 & n46787 ;
  assign n46789 = ~n46786 & ~n46788 ;
  assign n46790 = \m6_data_i[29]_pad  & n13697 ;
  assign n46791 = n13690 & n46790 ;
  assign n46792 = \m5_data_i[29]_pad  & ~n13697 ;
  assign n46793 = n13722 & n46792 ;
  assign n46794 = ~n46791 & ~n46793 ;
  assign n46795 = n46789 & n46794 ;
  assign n46796 = n46784 & n46795 ;
  assign n46797 = \m1_data_i[2]_pad  & ~n13697 ;
  assign n46798 = n13705 & n46797 ;
  assign n46799 = \m2_data_i[2]_pad  & n13697 ;
  assign n46800 = n13714 & n46799 ;
  assign n46801 = ~n46798 & ~n46800 ;
  assign n46802 = \m0_data_i[2]_pad  & n13697 ;
  assign n46803 = n13705 & n46802 ;
  assign n46804 = \m4_data_i[2]_pad  & n13697 ;
  assign n46805 = n13722 & n46804 ;
  assign n46806 = ~n46803 & ~n46805 ;
  assign n46807 = n46801 & n46806 ;
  assign n46808 = \m7_data_i[2]_pad  & ~n13697 ;
  assign n46809 = n13690 & n46808 ;
  assign n46810 = \m3_data_i[2]_pad  & ~n13697 ;
  assign n46811 = n13714 & n46810 ;
  assign n46812 = ~n46809 & ~n46811 ;
  assign n46813 = \m6_data_i[2]_pad  & n13697 ;
  assign n46814 = n13690 & n46813 ;
  assign n46815 = \m5_data_i[2]_pad  & ~n13697 ;
  assign n46816 = n13722 & n46815 ;
  assign n46817 = ~n46814 & ~n46816 ;
  assign n46818 = n46812 & n46817 ;
  assign n46819 = n46807 & n46818 ;
  assign n46820 = \m3_data_i[30]_pad  & ~n13697 ;
  assign n46821 = n13714 & n46820 ;
  assign n46822 = \m4_data_i[30]_pad  & n13697 ;
  assign n46823 = n13722 & n46822 ;
  assign n46824 = ~n46821 & ~n46823 ;
  assign n46825 = \m6_data_i[30]_pad  & n13697 ;
  assign n46826 = n13690 & n46825 ;
  assign n46827 = \m7_data_i[30]_pad  & ~n13697 ;
  assign n46828 = n13690 & n46827 ;
  assign n46829 = ~n46826 & ~n46828 ;
  assign n46830 = n46824 & n46829 ;
  assign n46831 = \m5_data_i[30]_pad  & ~n13697 ;
  assign n46832 = n13722 & n46831 ;
  assign n46833 = \m0_data_i[30]_pad  & n13697 ;
  assign n46834 = n13705 & n46833 ;
  assign n46835 = ~n46832 & ~n46834 ;
  assign n46836 = \m1_data_i[30]_pad  & ~n13697 ;
  assign n46837 = n13705 & n46836 ;
  assign n46838 = \m2_data_i[30]_pad  & n13697 ;
  assign n46839 = n13714 & n46838 ;
  assign n46840 = ~n46837 & ~n46839 ;
  assign n46841 = n46835 & n46840 ;
  assign n46842 = n46830 & n46841 ;
  assign n46843 = \m3_data_i[31]_pad  & ~n13697 ;
  assign n46844 = n13714 & n46843 ;
  assign n46845 = \m4_data_i[31]_pad  & n13697 ;
  assign n46846 = n13722 & n46845 ;
  assign n46847 = ~n46844 & ~n46846 ;
  assign n46848 = \m6_data_i[31]_pad  & n13697 ;
  assign n46849 = n13690 & n46848 ;
  assign n46850 = \m2_data_i[31]_pad  & n13697 ;
  assign n46851 = n13714 & n46850 ;
  assign n46852 = ~n46849 & ~n46851 ;
  assign n46853 = n46847 & n46852 ;
  assign n46854 = \m5_data_i[31]_pad  & ~n13697 ;
  assign n46855 = n13722 & n46854 ;
  assign n46856 = \m1_data_i[31]_pad  & ~n13697 ;
  assign n46857 = n13705 & n46856 ;
  assign n46858 = ~n46855 & ~n46857 ;
  assign n46859 = \m0_data_i[31]_pad  & n13697 ;
  assign n46860 = n13705 & n46859 ;
  assign n46861 = \m7_data_i[31]_pad  & ~n13697 ;
  assign n46862 = n13690 & n46861 ;
  assign n46863 = ~n46860 & ~n46862 ;
  assign n46864 = n46858 & n46863 ;
  assign n46865 = n46853 & n46864 ;
  assign n46866 = \m3_data_i[3]_pad  & ~n13697 ;
  assign n46867 = n13714 & n46866 ;
  assign n46868 = \m4_data_i[3]_pad  & n13697 ;
  assign n46869 = n13722 & n46868 ;
  assign n46870 = ~n46867 & ~n46869 ;
  assign n46871 = \m6_data_i[3]_pad  & n13697 ;
  assign n46872 = n13690 & n46871 ;
  assign n46873 = \m2_data_i[3]_pad  & n13697 ;
  assign n46874 = n13714 & n46873 ;
  assign n46875 = ~n46872 & ~n46874 ;
  assign n46876 = n46870 & n46875 ;
  assign n46877 = \m5_data_i[3]_pad  & ~n13697 ;
  assign n46878 = n13722 & n46877 ;
  assign n46879 = \m1_data_i[3]_pad  & ~n13697 ;
  assign n46880 = n13705 & n46879 ;
  assign n46881 = ~n46878 & ~n46880 ;
  assign n46882 = \m0_data_i[3]_pad  & n13697 ;
  assign n46883 = n13705 & n46882 ;
  assign n46884 = \m7_data_i[3]_pad  & ~n13697 ;
  assign n46885 = n13690 & n46884 ;
  assign n46886 = ~n46883 & ~n46885 ;
  assign n46887 = n46881 & n46886 ;
  assign n46888 = n46876 & n46887 ;
  assign n46889 = \m1_data_i[4]_pad  & ~n13697 ;
  assign n46890 = n13705 & n46889 ;
  assign n46891 = \m2_data_i[4]_pad  & n13697 ;
  assign n46892 = n13714 & n46891 ;
  assign n46893 = ~n46890 & ~n46892 ;
  assign n46894 = \m6_data_i[4]_pad  & n13697 ;
  assign n46895 = n13690 & n46894 ;
  assign n46896 = \m7_data_i[4]_pad  & ~n13697 ;
  assign n46897 = n13690 & n46896 ;
  assign n46898 = ~n46895 & ~n46897 ;
  assign n46899 = n46893 & n46898 ;
  assign n46900 = \m5_data_i[4]_pad  & ~n13697 ;
  assign n46901 = n13722 & n46900 ;
  assign n46902 = \m0_data_i[4]_pad  & n13697 ;
  assign n46903 = n13705 & n46902 ;
  assign n46904 = ~n46901 & ~n46903 ;
  assign n46905 = \m3_data_i[4]_pad  & ~n13697 ;
  assign n46906 = n13714 & n46905 ;
  assign n46907 = \m4_data_i[4]_pad  & n13697 ;
  assign n46908 = n13722 & n46907 ;
  assign n46909 = ~n46906 & ~n46908 ;
  assign n46910 = n46904 & n46909 ;
  assign n46911 = n46899 & n46910 ;
  assign n46912 = \m1_data_i[5]_pad  & ~n13697 ;
  assign n46913 = n13705 & n46912 ;
  assign n46914 = \m2_data_i[5]_pad  & n13697 ;
  assign n46915 = n13714 & n46914 ;
  assign n46916 = ~n46913 & ~n46915 ;
  assign n46917 = \m0_data_i[5]_pad  & n13697 ;
  assign n46918 = n13705 & n46917 ;
  assign n46919 = \m4_data_i[5]_pad  & n13697 ;
  assign n46920 = n13722 & n46919 ;
  assign n46921 = ~n46918 & ~n46920 ;
  assign n46922 = n46916 & n46921 ;
  assign n46923 = \m7_data_i[5]_pad  & ~n13697 ;
  assign n46924 = n13690 & n46923 ;
  assign n46925 = \m3_data_i[5]_pad  & ~n13697 ;
  assign n46926 = n13714 & n46925 ;
  assign n46927 = ~n46924 & ~n46926 ;
  assign n46928 = \m6_data_i[5]_pad  & n13697 ;
  assign n46929 = n13690 & n46928 ;
  assign n46930 = \m5_data_i[5]_pad  & ~n13697 ;
  assign n46931 = n13722 & n46930 ;
  assign n46932 = ~n46929 & ~n46931 ;
  assign n46933 = n46927 & n46932 ;
  assign n46934 = n46922 & n46933 ;
  assign n46935 = \m6_data_i[6]_pad  & n13697 ;
  assign n46936 = n13690 & n46935 ;
  assign n46937 = \m5_data_i[6]_pad  & ~n13697 ;
  assign n46938 = n13722 & n46937 ;
  assign n46939 = ~n46936 & ~n46938 ;
  assign n46940 = \m3_data_i[6]_pad  & ~n13697 ;
  assign n46941 = n13714 & n46940 ;
  assign n46942 = \m7_data_i[6]_pad  & ~n13697 ;
  assign n46943 = n13690 & n46942 ;
  assign n46944 = ~n46941 & ~n46943 ;
  assign n46945 = n46939 & n46944 ;
  assign n46946 = \m4_data_i[6]_pad  & n13697 ;
  assign n46947 = n13722 & n46946 ;
  assign n46948 = \m0_data_i[6]_pad  & n13697 ;
  assign n46949 = n13705 & n46948 ;
  assign n46950 = ~n46947 & ~n46949 ;
  assign n46951 = \m1_data_i[6]_pad  & ~n13697 ;
  assign n46952 = n13705 & n46951 ;
  assign n46953 = \m2_data_i[6]_pad  & n13697 ;
  assign n46954 = n13714 & n46953 ;
  assign n46955 = ~n46952 & ~n46954 ;
  assign n46956 = n46950 & n46955 ;
  assign n46957 = n46945 & n46956 ;
  assign n46958 = \m1_data_i[7]_pad  & ~n13697 ;
  assign n46959 = n13705 & n46958 ;
  assign n46960 = \m2_data_i[7]_pad  & n13697 ;
  assign n46961 = n13714 & n46960 ;
  assign n46962 = ~n46959 & ~n46961 ;
  assign n46963 = \m6_data_i[7]_pad  & n13697 ;
  assign n46964 = n13690 & n46963 ;
  assign n46965 = \m7_data_i[7]_pad  & ~n13697 ;
  assign n46966 = n13690 & n46965 ;
  assign n46967 = ~n46964 & ~n46966 ;
  assign n46968 = n46962 & n46967 ;
  assign n46969 = \m5_data_i[7]_pad  & ~n13697 ;
  assign n46970 = n13722 & n46969 ;
  assign n46971 = \m0_data_i[7]_pad  & n13697 ;
  assign n46972 = n13705 & n46971 ;
  assign n46973 = ~n46970 & ~n46972 ;
  assign n46974 = \m3_data_i[7]_pad  & ~n13697 ;
  assign n46975 = n13714 & n46974 ;
  assign n46976 = \m4_data_i[7]_pad  & n13697 ;
  assign n46977 = n13722 & n46976 ;
  assign n46978 = ~n46975 & ~n46977 ;
  assign n46979 = n46973 & n46978 ;
  assign n46980 = n46968 & n46979 ;
  assign n46981 = \m1_data_i[8]_pad  & ~n13697 ;
  assign n46982 = n13705 & n46981 ;
  assign n46983 = \m2_data_i[8]_pad  & n13697 ;
  assign n46984 = n13714 & n46983 ;
  assign n46985 = ~n46982 & ~n46984 ;
  assign n46986 = \m3_data_i[8]_pad  & ~n13697 ;
  assign n46987 = n13714 & n46986 ;
  assign n46988 = \m7_data_i[8]_pad  & ~n13697 ;
  assign n46989 = n13690 & n46988 ;
  assign n46990 = ~n46987 & ~n46989 ;
  assign n46991 = n46985 & n46990 ;
  assign n46992 = \m4_data_i[8]_pad  & n13697 ;
  assign n46993 = n13722 & n46992 ;
  assign n46994 = \m0_data_i[8]_pad  & n13697 ;
  assign n46995 = n13705 & n46994 ;
  assign n46996 = ~n46993 & ~n46995 ;
  assign n46997 = \m6_data_i[8]_pad  & n13697 ;
  assign n46998 = n13690 & n46997 ;
  assign n46999 = \m5_data_i[8]_pad  & ~n13697 ;
  assign n47000 = n13722 & n46999 ;
  assign n47001 = ~n46998 & ~n47000 ;
  assign n47002 = n46996 & n47001 ;
  assign n47003 = n46991 & n47002 ;
  assign n47004 = \m0_data_i[9]_pad  & n13697 ;
  assign n47005 = n13705 & n47004 ;
  assign n47006 = \m7_data_i[9]_pad  & ~n13697 ;
  assign n47007 = n13690 & n47006 ;
  assign n47008 = ~n47005 & ~n47007 ;
  assign n47009 = \m3_data_i[9]_pad  & ~n13697 ;
  assign n47010 = n13714 & n47009 ;
  assign n47011 = \m2_data_i[9]_pad  & n13697 ;
  assign n47012 = n13714 & n47011 ;
  assign n47013 = ~n47010 & ~n47012 ;
  assign n47014 = n47008 & n47013 ;
  assign n47015 = \m4_data_i[9]_pad  & n13697 ;
  assign n47016 = n13722 & n47015 ;
  assign n47017 = \m1_data_i[9]_pad  & ~n13697 ;
  assign n47018 = n13705 & n47017 ;
  assign n47019 = ~n47016 & ~n47018 ;
  assign n47020 = \m6_data_i[9]_pad  & n13697 ;
  assign n47021 = n13690 & n47020 ;
  assign n47022 = \m5_data_i[9]_pad  & ~n13697 ;
  assign n47023 = n13722 & n47022 ;
  assign n47024 = ~n47021 & ~n47023 ;
  assign n47025 = n47019 & n47024 ;
  assign n47026 = n47014 & n47025 ;
  assign n47027 = \m3_sel_i[0]_pad  & ~n13697 ;
  assign n47028 = n13714 & n47027 ;
  assign n47029 = \m4_sel_i[0]_pad  & n13697 ;
  assign n47030 = n13722 & n47029 ;
  assign n47031 = ~n47028 & ~n47030 ;
  assign n47032 = \m6_sel_i[0]_pad  & n13697 ;
  assign n47033 = n13690 & n47032 ;
  assign n47034 = \m2_sel_i[0]_pad  & n13697 ;
  assign n47035 = n13714 & n47034 ;
  assign n47036 = ~n47033 & ~n47035 ;
  assign n47037 = n47031 & n47036 ;
  assign n47038 = \m5_sel_i[0]_pad  & ~n13697 ;
  assign n47039 = n13722 & n47038 ;
  assign n47040 = \m1_sel_i[0]_pad  & ~n13697 ;
  assign n47041 = n13705 & n47040 ;
  assign n47042 = ~n47039 & ~n47041 ;
  assign n47043 = \m0_sel_i[0]_pad  & n13697 ;
  assign n47044 = n13705 & n47043 ;
  assign n47045 = \m7_sel_i[0]_pad  & ~n13697 ;
  assign n47046 = n13690 & n47045 ;
  assign n47047 = ~n47044 & ~n47046 ;
  assign n47048 = n47042 & n47047 ;
  assign n47049 = n47037 & n47048 ;
  assign n47050 = \m1_sel_i[1]_pad  & ~n13697 ;
  assign n47051 = n13705 & n47050 ;
  assign n47052 = \m2_sel_i[1]_pad  & n13697 ;
  assign n47053 = n13714 & n47052 ;
  assign n47054 = ~n47051 & ~n47053 ;
  assign n47055 = \m6_sel_i[1]_pad  & n13697 ;
  assign n47056 = n13690 & n47055 ;
  assign n47057 = \m7_sel_i[1]_pad  & ~n13697 ;
  assign n47058 = n13690 & n47057 ;
  assign n47059 = ~n47056 & ~n47058 ;
  assign n47060 = n47054 & n47059 ;
  assign n47061 = \m5_sel_i[1]_pad  & ~n13697 ;
  assign n47062 = n13722 & n47061 ;
  assign n47063 = \m0_sel_i[1]_pad  & n13697 ;
  assign n47064 = n13705 & n47063 ;
  assign n47065 = ~n47062 & ~n47064 ;
  assign n47066 = \m3_sel_i[1]_pad  & ~n13697 ;
  assign n47067 = n13714 & n47066 ;
  assign n47068 = \m4_sel_i[1]_pad  & n13697 ;
  assign n47069 = n13722 & n47068 ;
  assign n47070 = ~n47067 & ~n47069 ;
  assign n47071 = n47065 & n47070 ;
  assign n47072 = n47060 & n47071 ;
  assign n47073 = \m3_sel_i[2]_pad  & ~n13697 ;
  assign n47074 = n13714 & n47073 ;
  assign n47075 = \m4_sel_i[2]_pad  & n13697 ;
  assign n47076 = n13722 & n47075 ;
  assign n47077 = ~n47074 & ~n47076 ;
  assign n47078 = \m6_sel_i[2]_pad  & n13697 ;
  assign n47079 = n13690 & n47078 ;
  assign n47080 = \m2_sel_i[2]_pad  & n13697 ;
  assign n47081 = n13714 & n47080 ;
  assign n47082 = ~n47079 & ~n47081 ;
  assign n47083 = n47077 & n47082 ;
  assign n47084 = \m5_sel_i[2]_pad  & ~n13697 ;
  assign n47085 = n13722 & n47084 ;
  assign n47086 = \m1_sel_i[2]_pad  & ~n13697 ;
  assign n47087 = n13705 & n47086 ;
  assign n47088 = ~n47085 & ~n47087 ;
  assign n47089 = \m0_sel_i[2]_pad  & n13697 ;
  assign n47090 = n13705 & n47089 ;
  assign n47091 = \m7_sel_i[2]_pad  & ~n13697 ;
  assign n47092 = n13690 & n47091 ;
  assign n47093 = ~n47090 & ~n47092 ;
  assign n47094 = n47088 & n47093 ;
  assign n47095 = n47083 & n47094 ;
  assign n47096 = \m3_sel_i[3]_pad  & ~n13697 ;
  assign n47097 = n13714 & n47096 ;
  assign n47098 = \m4_sel_i[3]_pad  & n13697 ;
  assign n47099 = n13722 & n47098 ;
  assign n47100 = ~n47097 & ~n47099 ;
  assign n47101 = \m6_sel_i[3]_pad  & n13697 ;
  assign n47102 = n13690 & n47101 ;
  assign n47103 = \m2_sel_i[3]_pad  & n13697 ;
  assign n47104 = n13714 & n47103 ;
  assign n47105 = ~n47102 & ~n47104 ;
  assign n47106 = n47100 & n47105 ;
  assign n47107 = \m5_sel_i[3]_pad  & ~n13697 ;
  assign n47108 = n13722 & n47107 ;
  assign n47109 = \m1_sel_i[3]_pad  & ~n13697 ;
  assign n47110 = n13705 & n47109 ;
  assign n47111 = ~n47108 & ~n47110 ;
  assign n47112 = \m0_sel_i[3]_pad  & n13697 ;
  assign n47113 = n13705 & n47112 ;
  assign n47114 = \m7_sel_i[3]_pad  & ~n13697 ;
  assign n47115 = n13690 & n47114 ;
  assign n47116 = ~n47113 & ~n47115 ;
  assign n47117 = n47111 & n47116 ;
  assign n47118 = n47106 & n47117 ;
  assign n47119 = \m5_stb_i_pad  & n14695 ;
  assign n47120 = ~n13697 & n47119 ;
  assign n47121 = n13722 & n47120 ;
  assign n47122 = \m4_stb_i_pad  & n14958 ;
  assign n47123 = n13697 & n47122 ;
  assign n47124 = n13722 & n47123 ;
  assign n47125 = ~n47121 & ~n47124 ;
  assign n47126 = \m6_stb_i_pad  & n15038 ;
  assign n47127 = n13697 & n47126 ;
  assign n47128 = n13690 & n47127 ;
  assign n47129 = \m1_stb_i_pad  & n14837 ;
  assign n47130 = ~n13697 & n47129 ;
  assign n47131 = n13705 & n47130 ;
  assign n47132 = ~n47128 & ~n47131 ;
  assign n47133 = n47125 & n47132 ;
  assign n47134 = \m7_stb_i_pad  & n14671 ;
  assign n47135 = ~n13697 & n47134 ;
  assign n47136 = n13690 & n47135 ;
  assign n47137 = \m3_stb_i_pad  & n14740 ;
  assign n47138 = ~n13697 & n47137 ;
  assign n47139 = n13714 & n47138 ;
  assign n47140 = ~n47136 & ~n47139 ;
  assign n47141 = \m2_stb_i_pad  & n15090 ;
  assign n47142 = n13697 & n47141 ;
  assign n47143 = n13714 & n47142 ;
  assign n47144 = \m0_stb_i_pad  & n14786 ;
  assign n47145 = n13697 & n47144 ;
  assign n47146 = n13705 & n47145 ;
  assign n47147 = ~n47143 & ~n47146 ;
  assign n47148 = n47140 & n47147 ;
  assign n47149 = n47133 & n47148 ;
  assign n47150 = \m1_we_i_pad  & ~n13697 ;
  assign n47151 = n13705 & n47150 ;
  assign n47152 = \m2_we_i_pad  & n13697 ;
  assign n47153 = n13714 & n47152 ;
  assign n47154 = ~n47151 & ~n47153 ;
  assign n47155 = \m6_we_i_pad  & n13697 ;
  assign n47156 = n13690 & n47155 ;
  assign n47157 = \m7_we_i_pad  & ~n13697 ;
  assign n47158 = n13690 & n47157 ;
  assign n47159 = ~n47156 & ~n47158 ;
  assign n47160 = n47154 & n47159 ;
  assign n47161 = \m5_we_i_pad  & ~n13697 ;
  assign n47162 = n13722 & n47161 ;
  assign n47163 = \m0_we_i_pad  & n13697 ;
  assign n47164 = n13705 & n47163 ;
  assign n47165 = ~n47162 & ~n47164 ;
  assign n47166 = \m3_we_i_pad  & ~n13697 ;
  assign n47167 = n13714 & n47166 ;
  assign n47168 = \m4_we_i_pad  & n13697 ;
  assign n47169 = n13722 & n47168 ;
  assign n47170 = ~n47167 & ~n47169 ;
  assign n47171 = n47165 & n47170 ;
  assign n47172 = n47160 & n47171 ;
  assign n47173 = \m1_addr_i[0]_pad  & ~n13767 ;
  assign n47174 = n13760 & n47173 ;
  assign n47175 = \m2_addr_i[0]_pad  & n13767 ;
  assign n47176 = n13775 & n47175 ;
  assign n47177 = ~n47174 & ~n47176 ;
  assign n47178 = \m6_addr_i[0]_pad  & n13767 ;
  assign n47179 = n13784 & n47178 ;
  assign n47180 = \m7_addr_i[0]_pad  & ~n13767 ;
  assign n47181 = n13784 & n47180 ;
  assign n47182 = ~n47179 & ~n47181 ;
  assign n47183 = n47177 & n47182 ;
  assign n47184 = \m5_addr_i[0]_pad  & ~n13767 ;
  assign n47185 = n13792 & n47184 ;
  assign n47186 = \m0_addr_i[0]_pad  & n13767 ;
  assign n47187 = n13760 & n47186 ;
  assign n47188 = ~n47185 & ~n47187 ;
  assign n47189 = \m3_addr_i[0]_pad  & ~n13767 ;
  assign n47190 = n13775 & n47189 ;
  assign n47191 = \m4_addr_i[0]_pad  & n13767 ;
  assign n47192 = n13792 & n47191 ;
  assign n47193 = ~n47190 & ~n47192 ;
  assign n47194 = n47188 & n47193 ;
  assign n47195 = n47183 & n47194 ;
  assign n47196 = \m3_addr_i[10]_pad  & ~n13767 ;
  assign n47197 = n13775 & n47196 ;
  assign n47198 = \m4_addr_i[10]_pad  & n13767 ;
  assign n47199 = n13792 & n47198 ;
  assign n47200 = ~n47197 & ~n47199 ;
  assign n47201 = \m6_addr_i[10]_pad  & n13767 ;
  assign n47202 = n13784 & n47201 ;
  assign n47203 = \m7_addr_i[10]_pad  & ~n13767 ;
  assign n47204 = n13784 & n47203 ;
  assign n47205 = ~n47202 & ~n47204 ;
  assign n47206 = n47200 & n47205 ;
  assign n47207 = \m5_addr_i[10]_pad  & ~n13767 ;
  assign n47208 = n13792 & n47207 ;
  assign n47209 = \m0_addr_i[10]_pad  & n13767 ;
  assign n47210 = n13760 & n47209 ;
  assign n47211 = ~n47208 & ~n47210 ;
  assign n47212 = \m1_addr_i[10]_pad  & ~n13767 ;
  assign n47213 = n13760 & n47212 ;
  assign n47214 = \m2_addr_i[10]_pad  & n13767 ;
  assign n47215 = n13775 & n47214 ;
  assign n47216 = ~n47213 & ~n47215 ;
  assign n47217 = n47211 & n47216 ;
  assign n47218 = n47206 & n47217 ;
  assign n47219 = \m3_addr_i[11]_pad  & ~n13767 ;
  assign n47220 = n13775 & n47219 ;
  assign n47221 = \m4_addr_i[11]_pad  & n13767 ;
  assign n47222 = n13792 & n47221 ;
  assign n47223 = ~n47220 & ~n47222 ;
  assign n47224 = \m6_addr_i[11]_pad  & n13767 ;
  assign n47225 = n13784 & n47224 ;
  assign n47226 = \m2_addr_i[11]_pad  & n13767 ;
  assign n47227 = n13775 & n47226 ;
  assign n47228 = ~n47225 & ~n47227 ;
  assign n47229 = n47223 & n47228 ;
  assign n47230 = \m5_addr_i[11]_pad  & ~n13767 ;
  assign n47231 = n13792 & n47230 ;
  assign n47232 = \m1_addr_i[11]_pad  & ~n13767 ;
  assign n47233 = n13760 & n47232 ;
  assign n47234 = ~n47231 & ~n47233 ;
  assign n47235 = \m0_addr_i[11]_pad  & n13767 ;
  assign n47236 = n13760 & n47235 ;
  assign n47237 = \m7_addr_i[11]_pad  & ~n13767 ;
  assign n47238 = n13784 & n47237 ;
  assign n47239 = ~n47236 & ~n47238 ;
  assign n47240 = n47234 & n47239 ;
  assign n47241 = n47229 & n47240 ;
  assign n47242 = \m1_addr_i[12]_pad  & ~n13767 ;
  assign n47243 = n13760 & n47242 ;
  assign n47244 = \m2_addr_i[12]_pad  & n13767 ;
  assign n47245 = n13775 & n47244 ;
  assign n47246 = ~n47243 & ~n47245 ;
  assign n47247 = \m3_addr_i[12]_pad  & ~n13767 ;
  assign n47248 = n13775 & n47247 ;
  assign n47249 = \m7_addr_i[12]_pad  & ~n13767 ;
  assign n47250 = n13784 & n47249 ;
  assign n47251 = ~n47248 & ~n47250 ;
  assign n47252 = n47246 & n47251 ;
  assign n47253 = \m4_addr_i[12]_pad  & n13767 ;
  assign n47254 = n13792 & n47253 ;
  assign n47255 = \m0_addr_i[12]_pad  & n13767 ;
  assign n47256 = n13760 & n47255 ;
  assign n47257 = ~n47254 & ~n47256 ;
  assign n47258 = \m6_addr_i[12]_pad  & n13767 ;
  assign n47259 = n13784 & n47258 ;
  assign n47260 = \m5_addr_i[12]_pad  & ~n13767 ;
  assign n47261 = n13792 & n47260 ;
  assign n47262 = ~n47259 & ~n47261 ;
  assign n47263 = n47257 & n47262 ;
  assign n47264 = n47252 & n47263 ;
  assign n47265 = \m3_addr_i[13]_pad  & ~n13767 ;
  assign n47266 = n13775 & n47265 ;
  assign n47267 = \m4_addr_i[13]_pad  & n13767 ;
  assign n47268 = n13792 & n47267 ;
  assign n47269 = ~n47266 & ~n47268 ;
  assign n47270 = \m6_addr_i[13]_pad  & n13767 ;
  assign n47271 = n13784 & n47270 ;
  assign n47272 = \m2_addr_i[13]_pad  & n13767 ;
  assign n47273 = n13775 & n47272 ;
  assign n47274 = ~n47271 & ~n47273 ;
  assign n47275 = n47269 & n47274 ;
  assign n47276 = \m5_addr_i[13]_pad  & ~n13767 ;
  assign n47277 = n13792 & n47276 ;
  assign n47278 = \m1_addr_i[13]_pad  & ~n13767 ;
  assign n47279 = n13760 & n47278 ;
  assign n47280 = ~n47277 & ~n47279 ;
  assign n47281 = \m0_addr_i[13]_pad  & n13767 ;
  assign n47282 = n13760 & n47281 ;
  assign n47283 = \m7_addr_i[13]_pad  & ~n13767 ;
  assign n47284 = n13784 & n47283 ;
  assign n47285 = ~n47282 & ~n47284 ;
  assign n47286 = n47280 & n47285 ;
  assign n47287 = n47275 & n47286 ;
  assign n47288 = \m3_addr_i[14]_pad  & ~n13767 ;
  assign n47289 = n13775 & n47288 ;
  assign n47290 = \m4_addr_i[14]_pad  & n13767 ;
  assign n47291 = n13792 & n47290 ;
  assign n47292 = ~n47289 & ~n47291 ;
  assign n47293 = \m6_addr_i[14]_pad  & n13767 ;
  assign n47294 = n13784 & n47293 ;
  assign n47295 = \m2_addr_i[14]_pad  & n13767 ;
  assign n47296 = n13775 & n47295 ;
  assign n47297 = ~n47294 & ~n47296 ;
  assign n47298 = n47292 & n47297 ;
  assign n47299 = \m5_addr_i[14]_pad  & ~n13767 ;
  assign n47300 = n13792 & n47299 ;
  assign n47301 = \m1_addr_i[14]_pad  & ~n13767 ;
  assign n47302 = n13760 & n47301 ;
  assign n47303 = ~n47300 & ~n47302 ;
  assign n47304 = \m0_addr_i[14]_pad  & n13767 ;
  assign n47305 = n13760 & n47304 ;
  assign n47306 = \m7_addr_i[14]_pad  & ~n13767 ;
  assign n47307 = n13784 & n47306 ;
  assign n47308 = ~n47305 & ~n47307 ;
  assign n47309 = n47303 & n47308 ;
  assign n47310 = n47298 & n47309 ;
  assign n47311 = \m1_addr_i[15]_pad  & ~n13767 ;
  assign n47312 = n13760 & n47311 ;
  assign n47313 = \m2_addr_i[15]_pad  & n13767 ;
  assign n47314 = n13775 & n47313 ;
  assign n47315 = ~n47312 & ~n47314 ;
  assign n47316 = \m6_addr_i[15]_pad  & n13767 ;
  assign n47317 = n13784 & n47316 ;
  assign n47318 = \m7_addr_i[15]_pad  & ~n13767 ;
  assign n47319 = n13784 & n47318 ;
  assign n47320 = ~n47317 & ~n47319 ;
  assign n47321 = n47315 & n47320 ;
  assign n47322 = \m5_addr_i[15]_pad  & ~n13767 ;
  assign n47323 = n13792 & n47322 ;
  assign n47324 = \m0_addr_i[15]_pad  & n13767 ;
  assign n47325 = n13760 & n47324 ;
  assign n47326 = ~n47323 & ~n47325 ;
  assign n47327 = \m3_addr_i[15]_pad  & ~n13767 ;
  assign n47328 = n13775 & n47327 ;
  assign n47329 = \m4_addr_i[15]_pad  & n13767 ;
  assign n47330 = n13792 & n47329 ;
  assign n47331 = ~n47328 & ~n47330 ;
  assign n47332 = n47326 & n47331 ;
  assign n47333 = n47321 & n47332 ;
  assign n47334 = \m3_addr_i[16]_pad  & ~n13767 ;
  assign n47335 = n13775 & n47334 ;
  assign n47336 = \m4_addr_i[16]_pad  & n13767 ;
  assign n47337 = n13792 & n47336 ;
  assign n47338 = ~n47335 & ~n47337 ;
  assign n47339 = \m6_addr_i[16]_pad  & n13767 ;
  assign n47340 = n13784 & n47339 ;
  assign n47341 = \m7_addr_i[16]_pad  & ~n13767 ;
  assign n47342 = n13784 & n47341 ;
  assign n47343 = ~n47340 & ~n47342 ;
  assign n47344 = n47338 & n47343 ;
  assign n47345 = \m5_addr_i[16]_pad  & ~n13767 ;
  assign n47346 = n13792 & n47345 ;
  assign n47347 = \m0_addr_i[16]_pad  & n13767 ;
  assign n47348 = n13760 & n47347 ;
  assign n47349 = ~n47346 & ~n47348 ;
  assign n47350 = \m1_addr_i[16]_pad  & ~n13767 ;
  assign n47351 = n13760 & n47350 ;
  assign n47352 = \m2_addr_i[16]_pad  & n13767 ;
  assign n47353 = n13775 & n47352 ;
  assign n47354 = ~n47351 & ~n47353 ;
  assign n47355 = n47349 & n47354 ;
  assign n47356 = n47344 & n47355 ;
  assign n47357 = \m0_addr_i[17]_pad  & n13767 ;
  assign n47358 = n13760 & n47357 ;
  assign n47359 = \m7_addr_i[17]_pad  & ~n13767 ;
  assign n47360 = n13784 & n47359 ;
  assign n47361 = ~n47358 & ~n47360 ;
  assign n47362 = \m6_addr_i[17]_pad  & n13767 ;
  assign n47363 = n13784 & n47362 ;
  assign n47364 = \m2_addr_i[17]_pad  & n13767 ;
  assign n47365 = n13775 & n47364 ;
  assign n47366 = ~n47363 & ~n47365 ;
  assign n47367 = n47361 & n47366 ;
  assign n47368 = \m5_addr_i[17]_pad  & ~n13767 ;
  assign n47369 = n13792 & n47368 ;
  assign n47370 = \m1_addr_i[17]_pad  & ~n13767 ;
  assign n47371 = n13760 & n47370 ;
  assign n47372 = ~n47369 & ~n47371 ;
  assign n47373 = \m3_addr_i[17]_pad  & ~n13767 ;
  assign n47374 = n13775 & n47373 ;
  assign n47375 = \m4_addr_i[17]_pad  & n13767 ;
  assign n47376 = n13792 & n47375 ;
  assign n47377 = ~n47374 & ~n47376 ;
  assign n47378 = n47372 & n47377 ;
  assign n47379 = n47367 & n47378 ;
  assign n47380 = \m3_addr_i[18]_pad  & ~n13767 ;
  assign n47381 = n13775 & n47380 ;
  assign n47382 = \m4_addr_i[18]_pad  & n13767 ;
  assign n47383 = n13792 & n47382 ;
  assign n47384 = ~n47381 & ~n47383 ;
  assign n47385 = \m6_addr_i[18]_pad  & n13767 ;
  assign n47386 = n13784 & n47385 ;
  assign n47387 = \m7_addr_i[18]_pad  & ~n13767 ;
  assign n47388 = n13784 & n47387 ;
  assign n47389 = ~n47386 & ~n47388 ;
  assign n47390 = n47384 & n47389 ;
  assign n47391 = \m5_addr_i[18]_pad  & ~n13767 ;
  assign n47392 = n13792 & n47391 ;
  assign n47393 = \m0_addr_i[18]_pad  & n13767 ;
  assign n47394 = n13760 & n47393 ;
  assign n47395 = ~n47392 & ~n47394 ;
  assign n47396 = \m1_addr_i[18]_pad  & ~n13767 ;
  assign n47397 = n13760 & n47396 ;
  assign n47398 = \m2_addr_i[18]_pad  & n13767 ;
  assign n47399 = n13775 & n47398 ;
  assign n47400 = ~n47397 & ~n47399 ;
  assign n47401 = n47395 & n47400 ;
  assign n47402 = n47390 & n47401 ;
  assign n47403 = \m1_addr_i[19]_pad  & ~n13767 ;
  assign n47404 = n13760 & n47403 ;
  assign n47405 = \m2_addr_i[19]_pad  & n13767 ;
  assign n47406 = n13775 & n47405 ;
  assign n47407 = ~n47404 & ~n47406 ;
  assign n47408 = \m3_addr_i[19]_pad  & ~n13767 ;
  assign n47409 = n13775 & n47408 ;
  assign n47410 = \m7_addr_i[19]_pad  & ~n13767 ;
  assign n47411 = n13784 & n47410 ;
  assign n47412 = ~n47409 & ~n47411 ;
  assign n47413 = n47407 & n47412 ;
  assign n47414 = \m4_addr_i[19]_pad  & n13767 ;
  assign n47415 = n13792 & n47414 ;
  assign n47416 = \m0_addr_i[19]_pad  & n13767 ;
  assign n47417 = n13760 & n47416 ;
  assign n47418 = ~n47415 & ~n47417 ;
  assign n47419 = \m6_addr_i[19]_pad  & n13767 ;
  assign n47420 = n13784 & n47419 ;
  assign n47421 = \m5_addr_i[19]_pad  & ~n13767 ;
  assign n47422 = n13792 & n47421 ;
  assign n47423 = ~n47420 & ~n47422 ;
  assign n47424 = n47418 & n47423 ;
  assign n47425 = n47413 & n47424 ;
  assign n47426 = \m3_addr_i[1]_pad  & ~n13767 ;
  assign n47427 = n13775 & n47426 ;
  assign n47428 = \m4_addr_i[1]_pad  & n13767 ;
  assign n47429 = n13792 & n47428 ;
  assign n47430 = ~n47427 & ~n47429 ;
  assign n47431 = \m6_addr_i[1]_pad  & n13767 ;
  assign n47432 = n13784 & n47431 ;
  assign n47433 = \m7_addr_i[1]_pad  & ~n13767 ;
  assign n47434 = n13784 & n47433 ;
  assign n47435 = ~n47432 & ~n47434 ;
  assign n47436 = n47430 & n47435 ;
  assign n47437 = \m5_addr_i[1]_pad  & ~n13767 ;
  assign n47438 = n13792 & n47437 ;
  assign n47439 = \m0_addr_i[1]_pad  & n13767 ;
  assign n47440 = n13760 & n47439 ;
  assign n47441 = ~n47438 & ~n47440 ;
  assign n47442 = \m1_addr_i[1]_pad  & ~n13767 ;
  assign n47443 = n13760 & n47442 ;
  assign n47444 = \m2_addr_i[1]_pad  & n13767 ;
  assign n47445 = n13775 & n47444 ;
  assign n47446 = ~n47443 & ~n47445 ;
  assign n47447 = n47441 & n47446 ;
  assign n47448 = n47436 & n47447 ;
  assign n47449 = \m0_addr_i[20]_pad  & n13767 ;
  assign n47450 = n13760 & n47449 ;
  assign n47451 = \m7_addr_i[20]_pad  & ~n13767 ;
  assign n47452 = n13784 & n47451 ;
  assign n47453 = ~n47450 & ~n47452 ;
  assign n47454 = \m1_addr_i[20]_pad  & ~n13767 ;
  assign n47455 = n13760 & n47454 ;
  assign n47456 = \m4_addr_i[20]_pad  & n13767 ;
  assign n47457 = n13792 & n47456 ;
  assign n47458 = ~n47455 & ~n47457 ;
  assign n47459 = n47453 & n47458 ;
  assign n47460 = \m2_addr_i[20]_pad  & n13767 ;
  assign n47461 = n13775 & n47460 ;
  assign n47462 = \m3_addr_i[20]_pad  & ~n13767 ;
  assign n47463 = n13775 & n47462 ;
  assign n47464 = ~n47461 & ~n47463 ;
  assign n47465 = \m6_addr_i[20]_pad  & n13767 ;
  assign n47466 = n13784 & n47465 ;
  assign n47467 = \m5_addr_i[20]_pad  & ~n13767 ;
  assign n47468 = n13792 & n47467 ;
  assign n47469 = ~n47466 & ~n47468 ;
  assign n47470 = n47464 & n47469 ;
  assign n47471 = n47459 & n47470 ;
  assign n47472 = \m3_addr_i[21]_pad  & ~n13767 ;
  assign n47473 = n13775 & n47472 ;
  assign n47474 = \m4_addr_i[21]_pad  & n13767 ;
  assign n47475 = n13792 & n47474 ;
  assign n47476 = ~n47473 & ~n47475 ;
  assign n47477 = \m6_addr_i[21]_pad  & n13767 ;
  assign n47478 = n13784 & n47477 ;
  assign n47479 = \m2_addr_i[21]_pad  & n13767 ;
  assign n47480 = n13775 & n47479 ;
  assign n47481 = ~n47478 & ~n47480 ;
  assign n47482 = n47476 & n47481 ;
  assign n47483 = \m5_addr_i[21]_pad  & ~n13767 ;
  assign n47484 = n13792 & n47483 ;
  assign n47485 = \m1_addr_i[21]_pad  & ~n13767 ;
  assign n47486 = n13760 & n47485 ;
  assign n47487 = ~n47484 & ~n47486 ;
  assign n47488 = \m0_addr_i[21]_pad  & n13767 ;
  assign n47489 = n13760 & n47488 ;
  assign n47490 = \m7_addr_i[21]_pad  & ~n13767 ;
  assign n47491 = n13784 & n47490 ;
  assign n47492 = ~n47489 & ~n47491 ;
  assign n47493 = n47487 & n47492 ;
  assign n47494 = n47482 & n47493 ;
  assign n47495 = \m1_addr_i[22]_pad  & ~n13767 ;
  assign n47496 = n13760 & n47495 ;
  assign n47497 = \m2_addr_i[22]_pad  & n13767 ;
  assign n47498 = n13775 & n47497 ;
  assign n47499 = ~n47496 & ~n47498 ;
  assign n47500 = \m3_addr_i[22]_pad  & ~n13767 ;
  assign n47501 = n13775 & n47500 ;
  assign n47502 = \m7_addr_i[22]_pad  & ~n13767 ;
  assign n47503 = n13784 & n47502 ;
  assign n47504 = ~n47501 & ~n47503 ;
  assign n47505 = n47499 & n47504 ;
  assign n47506 = \m4_addr_i[22]_pad  & n13767 ;
  assign n47507 = n13792 & n47506 ;
  assign n47508 = \m0_addr_i[22]_pad  & n13767 ;
  assign n47509 = n13760 & n47508 ;
  assign n47510 = ~n47507 & ~n47509 ;
  assign n47511 = \m6_addr_i[22]_pad  & n13767 ;
  assign n47512 = n13784 & n47511 ;
  assign n47513 = \m5_addr_i[22]_pad  & ~n13767 ;
  assign n47514 = n13792 & n47513 ;
  assign n47515 = ~n47512 & ~n47514 ;
  assign n47516 = n47510 & n47515 ;
  assign n47517 = n47505 & n47516 ;
  assign n47518 = \m1_addr_i[23]_pad  & ~n13767 ;
  assign n47519 = n13760 & n47518 ;
  assign n47520 = \m2_addr_i[23]_pad  & n13767 ;
  assign n47521 = n13775 & n47520 ;
  assign n47522 = ~n47519 & ~n47521 ;
  assign n47523 = \m6_addr_i[23]_pad  & n13767 ;
  assign n47524 = n13784 & n47523 ;
  assign n47525 = \m7_addr_i[23]_pad  & ~n13767 ;
  assign n47526 = n13784 & n47525 ;
  assign n47527 = ~n47524 & ~n47526 ;
  assign n47528 = n47522 & n47527 ;
  assign n47529 = \m5_addr_i[23]_pad  & ~n13767 ;
  assign n47530 = n13792 & n47529 ;
  assign n47531 = \m0_addr_i[23]_pad  & n13767 ;
  assign n47532 = n13760 & n47531 ;
  assign n47533 = ~n47530 & ~n47532 ;
  assign n47534 = \m3_addr_i[23]_pad  & ~n13767 ;
  assign n47535 = n13775 & n47534 ;
  assign n47536 = \m4_addr_i[23]_pad  & n13767 ;
  assign n47537 = n13792 & n47536 ;
  assign n47538 = ~n47535 & ~n47537 ;
  assign n47539 = n47533 & n47538 ;
  assign n47540 = n47528 & n47539 ;
  assign n47541 = \m1_addr_i[24]_pad  & ~n13767 ;
  assign n47542 = n13760 & n47541 ;
  assign n47543 = \m2_addr_i[24]_pad  & n13767 ;
  assign n47544 = n13775 & n47543 ;
  assign n47545 = ~n47542 & ~n47544 ;
  assign n47546 = \m3_addr_i[24]_pad  & ~n13767 ;
  assign n47547 = n13775 & n47546 ;
  assign n47548 = \m7_addr_i[24]_pad  & ~n13767 ;
  assign n47549 = n13784 & n47548 ;
  assign n47550 = ~n47547 & ~n47549 ;
  assign n47551 = n47545 & n47550 ;
  assign n47552 = \m4_addr_i[24]_pad  & n13767 ;
  assign n47553 = n13792 & n47552 ;
  assign n47554 = \m0_addr_i[24]_pad  & n13767 ;
  assign n47555 = n13760 & n47554 ;
  assign n47556 = ~n47553 & ~n47555 ;
  assign n47557 = \m5_addr_i[24]_pad  & ~n13767 ;
  assign n47558 = n13792 & n47557 ;
  assign n47559 = \m6_addr_i[24]_pad  & n13767 ;
  assign n47560 = n13784 & n47559 ;
  assign n47561 = ~n47558 & ~n47560 ;
  assign n47562 = n47556 & n47561 ;
  assign n47563 = n47551 & n47562 ;
  assign n47564 = \m3_addr_i[25]_pad  & ~n13767 ;
  assign n47565 = n13775 & n47564 ;
  assign n47566 = \m4_addr_i[25]_pad  & n13767 ;
  assign n47567 = n13792 & n47566 ;
  assign n47568 = ~n47565 & ~n47567 ;
  assign n47569 = \m5_addr_i[25]_pad  & ~n13767 ;
  assign n47570 = n13792 & n47569 ;
  assign n47571 = \m2_addr_i[25]_pad  & n13767 ;
  assign n47572 = n13775 & n47571 ;
  assign n47573 = ~n47570 & ~n47572 ;
  assign n47574 = n47568 & n47573 ;
  assign n47575 = \m6_addr_i[25]_pad  & n13767 ;
  assign n47576 = n13784 & n47575 ;
  assign n47577 = \m1_addr_i[25]_pad  & ~n13767 ;
  assign n47578 = n13760 & n47577 ;
  assign n47579 = ~n47576 & ~n47578 ;
  assign n47580 = \m0_addr_i[25]_pad  & n13767 ;
  assign n47581 = n13760 & n47580 ;
  assign n47582 = \m7_addr_i[25]_pad  & ~n13767 ;
  assign n47583 = n13784 & n47582 ;
  assign n47584 = ~n47581 & ~n47583 ;
  assign n47585 = n47579 & n47584 ;
  assign n47586 = n47574 & n47585 ;
  assign n47587 = \m0_addr_i[26]_pad  & n13767 ;
  assign n47588 = n13760 & n47587 ;
  assign n47589 = \m7_addr_i[26]_pad  & ~n13767 ;
  assign n47590 = n13784 & n47589 ;
  assign n47591 = ~n47588 & ~n47590 ;
  assign n47592 = \m5_addr_i[26]_pad  & ~n13767 ;
  assign n47593 = n13792 & n47592 ;
  assign n47594 = \m2_addr_i[26]_pad  & n13767 ;
  assign n47595 = n13775 & n47594 ;
  assign n47596 = ~n47593 & ~n47595 ;
  assign n47597 = n47591 & n47596 ;
  assign n47598 = \m6_addr_i[26]_pad  & n13767 ;
  assign n47599 = n13784 & n47598 ;
  assign n47600 = \m1_addr_i[26]_pad  & ~n13767 ;
  assign n47601 = n13760 & n47600 ;
  assign n47602 = ~n47599 & ~n47601 ;
  assign n47603 = \m3_addr_i[26]_pad  & ~n13767 ;
  assign n47604 = n13775 & n47603 ;
  assign n47605 = \m4_addr_i[26]_pad  & n13767 ;
  assign n47606 = n13792 & n47605 ;
  assign n47607 = ~n47604 & ~n47606 ;
  assign n47608 = n47602 & n47607 ;
  assign n47609 = n47597 & n47608 ;
  assign n47610 = \m3_addr_i[27]_pad  & ~n13767 ;
  assign n47611 = n13775 & n47610 ;
  assign n47612 = \m4_addr_i[27]_pad  & n13767 ;
  assign n47613 = n13792 & n47612 ;
  assign n47614 = ~n47611 & ~n47613 ;
  assign n47615 = \m5_addr_i[27]_pad  & ~n13767 ;
  assign n47616 = n13792 & n47615 ;
  assign n47617 = \m2_addr_i[27]_pad  & n13767 ;
  assign n47618 = n13775 & n47617 ;
  assign n47619 = ~n47616 & ~n47618 ;
  assign n47620 = n47614 & n47619 ;
  assign n47621 = \m6_addr_i[27]_pad  & n13767 ;
  assign n47622 = n13784 & n47621 ;
  assign n47623 = \m1_addr_i[27]_pad  & ~n13767 ;
  assign n47624 = n13760 & n47623 ;
  assign n47625 = ~n47622 & ~n47624 ;
  assign n47626 = \m0_addr_i[27]_pad  & n13767 ;
  assign n47627 = n13760 & n47626 ;
  assign n47628 = \m7_addr_i[27]_pad  & ~n13767 ;
  assign n47629 = n13784 & n47628 ;
  assign n47630 = ~n47627 & ~n47629 ;
  assign n47631 = n47625 & n47630 ;
  assign n47632 = n47620 & n47631 ;
  assign n47633 = \m3_addr_i[28]_pad  & ~n13767 ;
  assign n47634 = n13775 & n47633 ;
  assign n47635 = \m4_addr_i[28]_pad  & n13767 ;
  assign n47636 = n13792 & n47635 ;
  assign n47637 = ~n47634 & ~n47636 ;
  assign n47638 = \m5_addr_i[28]_pad  & ~n13767 ;
  assign n47639 = n13792 & n47638 ;
  assign n47640 = \m7_addr_i[28]_pad  & ~n13767 ;
  assign n47641 = n13784 & n47640 ;
  assign n47642 = ~n47639 & ~n47641 ;
  assign n47643 = n47637 & n47642 ;
  assign n47644 = \m6_addr_i[28]_pad  & n13767 ;
  assign n47645 = n13784 & n47644 ;
  assign n47646 = \m0_addr_i[28]_pad  & n13767 ;
  assign n47647 = n13760 & n47646 ;
  assign n47648 = ~n47645 & ~n47647 ;
  assign n47649 = \m1_addr_i[28]_pad  & ~n13767 ;
  assign n47650 = n13760 & n47649 ;
  assign n47651 = \m2_addr_i[28]_pad  & n13767 ;
  assign n47652 = n13775 & n47651 ;
  assign n47653 = ~n47650 & ~n47652 ;
  assign n47654 = n47648 & n47653 ;
  assign n47655 = n47643 & n47654 ;
  assign n47656 = \m1_addr_i[29]_pad  & ~n13767 ;
  assign n47657 = n13760 & n47656 ;
  assign n47658 = \m2_addr_i[29]_pad  & n13767 ;
  assign n47659 = n13775 & n47658 ;
  assign n47660 = ~n47657 & ~n47659 ;
  assign n47661 = \m3_addr_i[29]_pad  & ~n13767 ;
  assign n47662 = n13775 & n47661 ;
  assign n47663 = \m6_addr_i[29]_pad  & n13767 ;
  assign n47664 = n13784 & n47663 ;
  assign n47665 = ~n47662 & ~n47664 ;
  assign n47666 = n47660 & n47665 ;
  assign n47667 = \m4_addr_i[29]_pad  & n13767 ;
  assign n47668 = n13792 & n47667 ;
  assign n47669 = \m5_addr_i[29]_pad  & ~n13767 ;
  assign n47670 = n13792 & n47669 ;
  assign n47671 = ~n47668 & ~n47670 ;
  assign n47672 = \m0_addr_i[29]_pad  & n13767 ;
  assign n47673 = n13760 & n47672 ;
  assign n47674 = \m7_addr_i[29]_pad  & ~n13767 ;
  assign n47675 = n13784 & n47674 ;
  assign n47676 = ~n47673 & ~n47675 ;
  assign n47677 = n47671 & n47676 ;
  assign n47678 = n47666 & n47677 ;
  assign n47679 = \m6_addr_i[2]_pad  & n13767 ;
  assign n47680 = n13784 & n47679 ;
  assign n47681 = \m5_addr_i[2]_pad  & ~n13767 ;
  assign n47682 = n13792 & n47681 ;
  assign n47683 = ~n47680 & ~n47682 ;
  assign n47684 = \m1_addr_i[2]_pad  & ~n13767 ;
  assign n47685 = n13760 & n47684 ;
  assign n47686 = \m4_addr_i[2]_pad  & n13767 ;
  assign n47687 = n13792 & n47686 ;
  assign n47688 = ~n47685 & ~n47687 ;
  assign n47689 = n47683 & n47688 ;
  assign n47690 = \m2_addr_i[2]_pad  & n13767 ;
  assign n47691 = n13775 & n47690 ;
  assign n47692 = \m3_addr_i[2]_pad  & ~n13767 ;
  assign n47693 = n13775 & n47692 ;
  assign n47694 = ~n47691 & ~n47693 ;
  assign n47695 = \m0_addr_i[2]_pad  & n13767 ;
  assign n47696 = n13760 & n47695 ;
  assign n47697 = \m7_addr_i[2]_pad  & ~n13767 ;
  assign n47698 = n13784 & n47697 ;
  assign n47699 = ~n47696 & ~n47698 ;
  assign n47700 = n47694 & n47699 ;
  assign n47701 = n47689 & n47700 ;
  assign n47702 = \m3_addr_i[30]_pad  & ~n13767 ;
  assign n47703 = n13775 & n47702 ;
  assign n47704 = \m4_addr_i[30]_pad  & n13767 ;
  assign n47705 = n13792 & n47704 ;
  assign n47706 = ~n47703 & ~n47705 ;
  assign n47707 = \m5_addr_i[30]_pad  & ~n13767 ;
  assign n47708 = n13792 & n47707 ;
  assign n47709 = \m7_addr_i[30]_pad  & ~n13767 ;
  assign n47710 = n13784 & n47709 ;
  assign n47711 = ~n47708 & ~n47710 ;
  assign n47712 = n47706 & n47711 ;
  assign n47713 = \m6_addr_i[30]_pad  & n13767 ;
  assign n47714 = n13784 & n47713 ;
  assign n47715 = \m0_addr_i[30]_pad  & n13767 ;
  assign n47716 = n13760 & n47715 ;
  assign n47717 = ~n47714 & ~n47716 ;
  assign n47718 = \m1_addr_i[30]_pad  & ~n13767 ;
  assign n47719 = n13760 & n47718 ;
  assign n47720 = \m2_addr_i[30]_pad  & n13767 ;
  assign n47721 = n13775 & n47720 ;
  assign n47722 = ~n47719 & ~n47721 ;
  assign n47723 = n47717 & n47722 ;
  assign n47724 = n47712 & n47723 ;
  assign n47725 = \m1_addr_i[31]_pad  & ~n13767 ;
  assign n47726 = n13760 & n47725 ;
  assign n47727 = \m2_addr_i[31]_pad  & n13767 ;
  assign n47728 = n13775 & n47727 ;
  assign n47729 = ~n47726 & ~n47728 ;
  assign n47730 = \m5_addr_i[31]_pad  & ~n13767 ;
  assign n47731 = n13792 & n47730 ;
  assign n47732 = \m7_addr_i[31]_pad  & ~n13767 ;
  assign n47733 = n13784 & n47732 ;
  assign n47734 = ~n47731 & ~n47733 ;
  assign n47735 = n47729 & n47734 ;
  assign n47736 = \m6_addr_i[31]_pad  & n13767 ;
  assign n47737 = n13784 & n47736 ;
  assign n47738 = \m0_addr_i[31]_pad  & n13767 ;
  assign n47739 = n13760 & n47738 ;
  assign n47740 = ~n47737 & ~n47739 ;
  assign n47741 = \m3_addr_i[31]_pad  & ~n13767 ;
  assign n47742 = n13775 & n47741 ;
  assign n47743 = \m4_addr_i[31]_pad  & n13767 ;
  assign n47744 = n13792 & n47743 ;
  assign n47745 = ~n47742 & ~n47744 ;
  assign n47746 = n47740 & n47745 ;
  assign n47747 = n47735 & n47746 ;
  assign n47748 = \m3_addr_i[3]_pad  & ~n13767 ;
  assign n47749 = n13775 & n47748 ;
  assign n47750 = \m4_addr_i[3]_pad  & n13767 ;
  assign n47751 = n13792 & n47750 ;
  assign n47752 = ~n47749 & ~n47751 ;
  assign n47753 = \m6_addr_i[3]_pad  & n13767 ;
  assign n47754 = n13784 & n47753 ;
  assign n47755 = \m2_addr_i[3]_pad  & n13767 ;
  assign n47756 = n13775 & n47755 ;
  assign n47757 = ~n47754 & ~n47756 ;
  assign n47758 = n47752 & n47757 ;
  assign n47759 = \m5_addr_i[3]_pad  & ~n13767 ;
  assign n47760 = n13792 & n47759 ;
  assign n47761 = \m1_addr_i[3]_pad  & ~n13767 ;
  assign n47762 = n13760 & n47761 ;
  assign n47763 = ~n47760 & ~n47762 ;
  assign n47764 = \m0_addr_i[3]_pad  & n13767 ;
  assign n47765 = n13760 & n47764 ;
  assign n47766 = \m7_addr_i[3]_pad  & ~n13767 ;
  assign n47767 = n13784 & n47766 ;
  assign n47768 = ~n47765 & ~n47767 ;
  assign n47769 = n47763 & n47768 ;
  assign n47770 = n47758 & n47769 ;
  assign n47771 = \m1_addr_i[4]_pad  & ~n13767 ;
  assign n47772 = n13760 & n47771 ;
  assign n47773 = \m2_addr_i[4]_pad  & n13767 ;
  assign n47774 = n13775 & n47773 ;
  assign n47775 = ~n47772 & ~n47774 ;
  assign n47776 = \m6_addr_i[4]_pad  & n13767 ;
  assign n47777 = n13784 & n47776 ;
  assign n47778 = \m7_addr_i[4]_pad  & ~n13767 ;
  assign n47779 = n13784 & n47778 ;
  assign n47780 = ~n47777 & ~n47779 ;
  assign n47781 = n47775 & n47780 ;
  assign n47782 = \m5_addr_i[4]_pad  & ~n13767 ;
  assign n47783 = n13792 & n47782 ;
  assign n47784 = \m0_addr_i[4]_pad  & n13767 ;
  assign n47785 = n13760 & n47784 ;
  assign n47786 = ~n47783 & ~n47785 ;
  assign n47787 = \m3_addr_i[4]_pad  & ~n13767 ;
  assign n47788 = n13775 & n47787 ;
  assign n47789 = \m4_addr_i[4]_pad  & n13767 ;
  assign n47790 = n13792 & n47789 ;
  assign n47791 = ~n47788 & ~n47790 ;
  assign n47792 = n47786 & n47791 ;
  assign n47793 = n47781 & n47792 ;
  assign n47794 = \m3_addr_i[5]_pad  & ~n13767 ;
  assign n47795 = n13775 & n47794 ;
  assign n47796 = \m4_addr_i[5]_pad  & n13767 ;
  assign n47797 = n13792 & n47796 ;
  assign n47798 = ~n47795 & ~n47797 ;
  assign n47799 = \m6_addr_i[5]_pad  & n13767 ;
  assign n47800 = n13784 & n47799 ;
  assign n47801 = \m2_addr_i[5]_pad  & n13767 ;
  assign n47802 = n13775 & n47801 ;
  assign n47803 = ~n47800 & ~n47802 ;
  assign n47804 = n47798 & n47803 ;
  assign n47805 = \m5_addr_i[5]_pad  & ~n13767 ;
  assign n47806 = n13792 & n47805 ;
  assign n47807 = \m1_addr_i[5]_pad  & ~n13767 ;
  assign n47808 = n13760 & n47807 ;
  assign n47809 = ~n47806 & ~n47808 ;
  assign n47810 = \m0_addr_i[5]_pad  & n13767 ;
  assign n47811 = n13760 & n47810 ;
  assign n47812 = \m7_addr_i[5]_pad  & ~n13767 ;
  assign n47813 = n13784 & n47812 ;
  assign n47814 = ~n47811 & ~n47813 ;
  assign n47815 = n47809 & n47814 ;
  assign n47816 = n47804 & n47815 ;
  assign n47817 = \m3_addr_i[6]_pad  & ~n13767 ;
  assign n47818 = n13775 & n47817 ;
  assign n47819 = \m4_addr_i[6]_pad  & n13767 ;
  assign n47820 = n13792 & n47819 ;
  assign n47821 = ~n47818 & ~n47820 ;
  assign n47822 = \m6_addr_i[6]_pad  & n13767 ;
  assign n47823 = n13784 & n47822 ;
  assign n47824 = \m2_addr_i[6]_pad  & n13767 ;
  assign n47825 = n13775 & n47824 ;
  assign n47826 = ~n47823 & ~n47825 ;
  assign n47827 = n47821 & n47826 ;
  assign n47828 = \m5_addr_i[6]_pad  & ~n13767 ;
  assign n47829 = n13792 & n47828 ;
  assign n47830 = \m1_addr_i[6]_pad  & ~n13767 ;
  assign n47831 = n13760 & n47830 ;
  assign n47832 = ~n47829 & ~n47831 ;
  assign n47833 = \m0_addr_i[6]_pad  & n13767 ;
  assign n47834 = n13760 & n47833 ;
  assign n47835 = \m7_addr_i[6]_pad  & ~n13767 ;
  assign n47836 = n13784 & n47835 ;
  assign n47837 = ~n47834 & ~n47836 ;
  assign n47838 = n47832 & n47837 ;
  assign n47839 = n47827 & n47838 ;
  assign n47840 = \m3_addr_i[7]_pad  & ~n13767 ;
  assign n47841 = n13775 & n47840 ;
  assign n47842 = \m4_addr_i[7]_pad  & n13767 ;
  assign n47843 = n13792 & n47842 ;
  assign n47844 = ~n47841 & ~n47843 ;
  assign n47845 = \m6_addr_i[7]_pad  & n13767 ;
  assign n47846 = n13784 & n47845 ;
  assign n47847 = \m2_addr_i[7]_pad  & n13767 ;
  assign n47848 = n13775 & n47847 ;
  assign n47849 = ~n47846 & ~n47848 ;
  assign n47850 = n47844 & n47849 ;
  assign n47851 = \m5_addr_i[7]_pad  & ~n13767 ;
  assign n47852 = n13792 & n47851 ;
  assign n47853 = \m1_addr_i[7]_pad  & ~n13767 ;
  assign n47854 = n13760 & n47853 ;
  assign n47855 = ~n47852 & ~n47854 ;
  assign n47856 = \m0_addr_i[7]_pad  & n13767 ;
  assign n47857 = n13760 & n47856 ;
  assign n47858 = \m7_addr_i[7]_pad  & ~n13767 ;
  assign n47859 = n13784 & n47858 ;
  assign n47860 = ~n47857 & ~n47859 ;
  assign n47861 = n47855 & n47860 ;
  assign n47862 = n47850 & n47861 ;
  assign n47863 = \m6_addr_i[8]_pad  & n13767 ;
  assign n47864 = n13784 & n47863 ;
  assign n47865 = \m5_addr_i[8]_pad  & ~n13767 ;
  assign n47866 = n13792 & n47865 ;
  assign n47867 = ~n47864 & ~n47866 ;
  assign n47868 = \m0_addr_i[8]_pad  & n13767 ;
  assign n47869 = n13760 & n47868 ;
  assign n47870 = \m4_addr_i[8]_pad  & n13767 ;
  assign n47871 = n13792 & n47870 ;
  assign n47872 = ~n47869 & ~n47871 ;
  assign n47873 = n47867 & n47872 ;
  assign n47874 = \m7_addr_i[8]_pad  & ~n13767 ;
  assign n47875 = n13784 & n47874 ;
  assign n47876 = \m3_addr_i[8]_pad  & ~n13767 ;
  assign n47877 = n13775 & n47876 ;
  assign n47878 = ~n47875 & ~n47877 ;
  assign n47879 = \m1_addr_i[8]_pad  & ~n13767 ;
  assign n47880 = n13760 & n47879 ;
  assign n47881 = \m2_addr_i[8]_pad  & n13767 ;
  assign n47882 = n13775 & n47881 ;
  assign n47883 = ~n47880 & ~n47882 ;
  assign n47884 = n47878 & n47883 ;
  assign n47885 = n47873 & n47884 ;
  assign n47886 = \m3_addr_i[9]_pad  & ~n13767 ;
  assign n47887 = n13775 & n47886 ;
  assign n47888 = \m4_addr_i[9]_pad  & n13767 ;
  assign n47889 = n13792 & n47888 ;
  assign n47890 = ~n47887 & ~n47889 ;
  assign n47891 = \m6_addr_i[9]_pad  & n13767 ;
  assign n47892 = n13784 & n47891 ;
  assign n47893 = \m2_addr_i[9]_pad  & n13767 ;
  assign n47894 = n13775 & n47893 ;
  assign n47895 = ~n47892 & ~n47894 ;
  assign n47896 = n47890 & n47895 ;
  assign n47897 = \m5_addr_i[9]_pad  & ~n13767 ;
  assign n47898 = n13792 & n47897 ;
  assign n47899 = \m1_addr_i[9]_pad  & ~n13767 ;
  assign n47900 = n13760 & n47899 ;
  assign n47901 = ~n47898 & ~n47900 ;
  assign n47902 = \m0_addr_i[9]_pad  & n13767 ;
  assign n47903 = n13760 & n47902 ;
  assign n47904 = \m7_addr_i[9]_pad  & ~n13767 ;
  assign n47905 = n13784 & n47904 ;
  assign n47906 = ~n47903 & ~n47905 ;
  assign n47907 = n47901 & n47906 ;
  assign n47908 = n47896 & n47907 ;
  assign n47909 = \m1_data_i[0]_pad  & ~n13767 ;
  assign n47910 = n13760 & n47909 ;
  assign n47911 = \m2_data_i[0]_pad  & n13767 ;
  assign n47912 = n13775 & n47911 ;
  assign n47913 = ~n47910 & ~n47912 ;
  assign n47914 = \m3_data_i[0]_pad  & ~n13767 ;
  assign n47915 = n13775 & n47914 ;
  assign n47916 = \m7_data_i[0]_pad  & ~n13767 ;
  assign n47917 = n13784 & n47916 ;
  assign n47918 = ~n47915 & ~n47917 ;
  assign n47919 = n47913 & n47918 ;
  assign n47920 = \m4_data_i[0]_pad  & n13767 ;
  assign n47921 = n13792 & n47920 ;
  assign n47922 = \m0_data_i[0]_pad  & n13767 ;
  assign n47923 = n13760 & n47922 ;
  assign n47924 = ~n47921 & ~n47923 ;
  assign n47925 = \m6_data_i[0]_pad  & n13767 ;
  assign n47926 = n13784 & n47925 ;
  assign n47927 = \m5_data_i[0]_pad  & ~n13767 ;
  assign n47928 = n13792 & n47927 ;
  assign n47929 = ~n47926 & ~n47928 ;
  assign n47930 = n47924 & n47929 ;
  assign n47931 = n47919 & n47930 ;
  assign n47932 = \m3_data_i[10]_pad  & ~n13767 ;
  assign n47933 = n13775 & n47932 ;
  assign n47934 = \m4_data_i[10]_pad  & n13767 ;
  assign n47935 = n13792 & n47934 ;
  assign n47936 = ~n47933 & ~n47935 ;
  assign n47937 = \m6_data_i[10]_pad  & n13767 ;
  assign n47938 = n13784 & n47937 ;
  assign n47939 = \m7_data_i[10]_pad  & ~n13767 ;
  assign n47940 = n13784 & n47939 ;
  assign n47941 = ~n47938 & ~n47940 ;
  assign n47942 = n47936 & n47941 ;
  assign n47943 = \m5_data_i[10]_pad  & ~n13767 ;
  assign n47944 = n13792 & n47943 ;
  assign n47945 = \m0_data_i[10]_pad  & n13767 ;
  assign n47946 = n13760 & n47945 ;
  assign n47947 = ~n47944 & ~n47946 ;
  assign n47948 = \m1_data_i[10]_pad  & ~n13767 ;
  assign n47949 = n13760 & n47948 ;
  assign n47950 = \m2_data_i[10]_pad  & n13767 ;
  assign n47951 = n13775 & n47950 ;
  assign n47952 = ~n47949 & ~n47951 ;
  assign n47953 = n47947 & n47952 ;
  assign n47954 = n47942 & n47953 ;
  assign n47955 = \m3_data_i[11]_pad  & ~n13767 ;
  assign n47956 = n13775 & n47955 ;
  assign n47957 = \m4_data_i[11]_pad  & n13767 ;
  assign n47958 = n13792 & n47957 ;
  assign n47959 = ~n47956 & ~n47958 ;
  assign n47960 = \m6_data_i[11]_pad  & n13767 ;
  assign n47961 = n13784 & n47960 ;
  assign n47962 = \m7_data_i[11]_pad  & ~n13767 ;
  assign n47963 = n13784 & n47962 ;
  assign n47964 = ~n47961 & ~n47963 ;
  assign n47965 = n47959 & n47964 ;
  assign n47966 = \m5_data_i[11]_pad  & ~n13767 ;
  assign n47967 = n13792 & n47966 ;
  assign n47968 = \m0_data_i[11]_pad  & n13767 ;
  assign n47969 = n13760 & n47968 ;
  assign n47970 = ~n47967 & ~n47969 ;
  assign n47971 = \m1_data_i[11]_pad  & ~n13767 ;
  assign n47972 = n13760 & n47971 ;
  assign n47973 = \m2_data_i[11]_pad  & n13767 ;
  assign n47974 = n13775 & n47973 ;
  assign n47975 = ~n47972 & ~n47974 ;
  assign n47976 = n47970 & n47975 ;
  assign n47977 = n47965 & n47976 ;
  assign n47978 = \m3_data_i[12]_pad  & ~n13767 ;
  assign n47979 = n13775 & n47978 ;
  assign n47980 = \m4_data_i[12]_pad  & n13767 ;
  assign n47981 = n13792 & n47980 ;
  assign n47982 = ~n47979 & ~n47981 ;
  assign n47983 = \m6_data_i[12]_pad  & n13767 ;
  assign n47984 = n13784 & n47983 ;
  assign n47985 = \m7_data_i[12]_pad  & ~n13767 ;
  assign n47986 = n13784 & n47985 ;
  assign n47987 = ~n47984 & ~n47986 ;
  assign n47988 = n47982 & n47987 ;
  assign n47989 = \m5_data_i[12]_pad  & ~n13767 ;
  assign n47990 = n13792 & n47989 ;
  assign n47991 = \m0_data_i[12]_pad  & n13767 ;
  assign n47992 = n13760 & n47991 ;
  assign n47993 = ~n47990 & ~n47992 ;
  assign n47994 = \m1_data_i[12]_pad  & ~n13767 ;
  assign n47995 = n13760 & n47994 ;
  assign n47996 = \m2_data_i[12]_pad  & n13767 ;
  assign n47997 = n13775 & n47996 ;
  assign n47998 = ~n47995 & ~n47997 ;
  assign n47999 = n47993 & n47998 ;
  assign n48000 = n47988 & n47999 ;
  assign n48001 = \m3_data_i[13]_pad  & ~n13767 ;
  assign n48002 = n13775 & n48001 ;
  assign n48003 = \m4_data_i[13]_pad  & n13767 ;
  assign n48004 = n13792 & n48003 ;
  assign n48005 = ~n48002 & ~n48004 ;
  assign n48006 = \m6_data_i[13]_pad  & n13767 ;
  assign n48007 = n13784 & n48006 ;
  assign n48008 = \m2_data_i[13]_pad  & n13767 ;
  assign n48009 = n13775 & n48008 ;
  assign n48010 = ~n48007 & ~n48009 ;
  assign n48011 = n48005 & n48010 ;
  assign n48012 = \m5_data_i[13]_pad  & ~n13767 ;
  assign n48013 = n13792 & n48012 ;
  assign n48014 = \m1_data_i[13]_pad  & ~n13767 ;
  assign n48015 = n13760 & n48014 ;
  assign n48016 = ~n48013 & ~n48015 ;
  assign n48017 = \m0_data_i[13]_pad  & n13767 ;
  assign n48018 = n13760 & n48017 ;
  assign n48019 = \m7_data_i[13]_pad  & ~n13767 ;
  assign n48020 = n13784 & n48019 ;
  assign n48021 = ~n48018 & ~n48020 ;
  assign n48022 = n48016 & n48021 ;
  assign n48023 = n48011 & n48022 ;
  assign n48024 = \m1_data_i[14]_pad  & ~n13767 ;
  assign n48025 = n13760 & n48024 ;
  assign n48026 = \m2_data_i[14]_pad  & n13767 ;
  assign n48027 = n13775 & n48026 ;
  assign n48028 = ~n48025 & ~n48027 ;
  assign n48029 = \m6_data_i[14]_pad  & n13767 ;
  assign n48030 = n13784 & n48029 ;
  assign n48031 = \m7_data_i[14]_pad  & ~n13767 ;
  assign n48032 = n13784 & n48031 ;
  assign n48033 = ~n48030 & ~n48032 ;
  assign n48034 = n48028 & n48033 ;
  assign n48035 = \m5_data_i[14]_pad  & ~n13767 ;
  assign n48036 = n13792 & n48035 ;
  assign n48037 = \m0_data_i[14]_pad  & n13767 ;
  assign n48038 = n13760 & n48037 ;
  assign n48039 = ~n48036 & ~n48038 ;
  assign n48040 = \m3_data_i[14]_pad  & ~n13767 ;
  assign n48041 = n13775 & n48040 ;
  assign n48042 = \m4_data_i[14]_pad  & n13767 ;
  assign n48043 = n13792 & n48042 ;
  assign n48044 = ~n48041 & ~n48043 ;
  assign n48045 = n48039 & n48044 ;
  assign n48046 = n48034 & n48045 ;
  assign n48047 = \m3_data_i[15]_pad  & ~n13767 ;
  assign n48048 = n13775 & n48047 ;
  assign n48049 = \m4_data_i[15]_pad  & n13767 ;
  assign n48050 = n13792 & n48049 ;
  assign n48051 = ~n48048 & ~n48050 ;
  assign n48052 = \m6_data_i[15]_pad  & n13767 ;
  assign n48053 = n13784 & n48052 ;
  assign n48054 = \m2_data_i[15]_pad  & n13767 ;
  assign n48055 = n13775 & n48054 ;
  assign n48056 = ~n48053 & ~n48055 ;
  assign n48057 = n48051 & n48056 ;
  assign n48058 = \m5_data_i[15]_pad  & ~n13767 ;
  assign n48059 = n13792 & n48058 ;
  assign n48060 = \m1_data_i[15]_pad  & ~n13767 ;
  assign n48061 = n13760 & n48060 ;
  assign n48062 = ~n48059 & ~n48061 ;
  assign n48063 = \m0_data_i[15]_pad  & n13767 ;
  assign n48064 = n13760 & n48063 ;
  assign n48065 = \m7_data_i[15]_pad  & ~n13767 ;
  assign n48066 = n13784 & n48065 ;
  assign n48067 = ~n48064 & ~n48066 ;
  assign n48068 = n48062 & n48067 ;
  assign n48069 = n48057 & n48068 ;
  assign n48070 = \m3_data_i[16]_pad  & ~n13767 ;
  assign n48071 = n13775 & n48070 ;
  assign n48072 = \m4_data_i[16]_pad  & n13767 ;
  assign n48073 = n13792 & n48072 ;
  assign n48074 = ~n48071 & ~n48073 ;
  assign n48075 = \m6_data_i[16]_pad  & n13767 ;
  assign n48076 = n13784 & n48075 ;
  assign n48077 = \m2_data_i[16]_pad  & n13767 ;
  assign n48078 = n13775 & n48077 ;
  assign n48079 = ~n48076 & ~n48078 ;
  assign n48080 = n48074 & n48079 ;
  assign n48081 = \m5_data_i[16]_pad  & ~n13767 ;
  assign n48082 = n13792 & n48081 ;
  assign n48083 = \m1_data_i[16]_pad  & ~n13767 ;
  assign n48084 = n13760 & n48083 ;
  assign n48085 = ~n48082 & ~n48084 ;
  assign n48086 = \m0_data_i[16]_pad  & n13767 ;
  assign n48087 = n13760 & n48086 ;
  assign n48088 = \m7_data_i[16]_pad  & ~n13767 ;
  assign n48089 = n13784 & n48088 ;
  assign n48090 = ~n48087 & ~n48089 ;
  assign n48091 = n48085 & n48090 ;
  assign n48092 = n48080 & n48091 ;
  assign n48093 = \m3_data_i[17]_pad  & ~n13767 ;
  assign n48094 = n13775 & n48093 ;
  assign n48095 = \m4_data_i[17]_pad  & n13767 ;
  assign n48096 = n13792 & n48095 ;
  assign n48097 = ~n48094 & ~n48096 ;
  assign n48098 = \m6_data_i[17]_pad  & n13767 ;
  assign n48099 = n13784 & n48098 ;
  assign n48100 = \m7_data_i[17]_pad  & ~n13767 ;
  assign n48101 = n13784 & n48100 ;
  assign n48102 = ~n48099 & ~n48101 ;
  assign n48103 = n48097 & n48102 ;
  assign n48104 = \m5_data_i[17]_pad  & ~n13767 ;
  assign n48105 = n13792 & n48104 ;
  assign n48106 = \m0_data_i[17]_pad  & n13767 ;
  assign n48107 = n13760 & n48106 ;
  assign n48108 = ~n48105 & ~n48107 ;
  assign n48109 = \m1_data_i[17]_pad  & ~n13767 ;
  assign n48110 = n13760 & n48109 ;
  assign n48111 = \m2_data_i[17]_pad  & n13767 ;
  assign n48112 = n13775 & n48111 ;
  assign n48113 = ~n48110 & ~n48112 ;
  assign n48114 = n48108 & n48113 ;
  assign n48115 = n48103 & n48114 ;
  assign n48116 = \m1_data_i[18]_pad  & ~n13767 ;
  assign n48117 = n13760 & n48116 ;
  assign n48118 = \m2_data_i[18]_pad  & n13767 ;
  assign n48119 = n13775 & n48118 ;
  assign n48120 = ~n48117 & ~n48119 ;
  assign n48121 = \m3_data_i[18]_pad  & ~n13767 ;
  assign n48122 = n13775 & n48121 ;
  assign n48123 = \m7_data_i[18]_pad  & ~n13767 ;
  assign n48124 = n13784 & n48123 ;
  assign n48125 = ~n48122 & ~n48124 ;
  assign n48126 = n48120 & n48125 ;
  assign n48127 = \m4_data_i[18]_pad  & n13767 ;
  assign n48128 = n13792 & n48127 ;
  assign n48129 = \m0_data_i[18]_pad  & n13767 ;
  assign n48130 = n13760 & n48129 ;
  assign n48131 = ~n48128 & ~n48130 ;
  assign n48132 = \m6_data_i[18]_pad  & n13767 ;
  assign n48133 = n13784 & n48132 ;
  assign n48134 = \m5_data_i[18]_pad  & ~n13767 ;
  assign n48135 = n13792 & n48134 ;
  assign n48136 = ~n48133 & ~n48135 ;
  assign n48137 = n48131 & n48136 ;
  assign n48138 = n48126 & n48137 ;
  assign n48139 = \m1_data_i[19]_pad  & ~n13767 ;
  assign n48140 = n13760 & n48139 ;
  assign n48141 = \m2_data_i[19]_pad  & n13767 ;
  assign n48142 = n13775 & n48141 ;
  assign n48143 = ~n48140 & ~n48142 ;
  assign n48144 = \m6_data_i[19]_pad  & n13767 ;
  assign n48145 = n13784 & n48144 ;
  assign n48146 = \m7_data_i[19]_pad  & ~n13767 ;
  assign n48147 = n13784 & n48146 ;
  assign n48148 = ~n48145 & ~n48147 ;
  assign n48149 = n48143 & n48148 ;
  assign n48150 = \m5_data_i[19]_pad  & ~n13767 ;
  assign n48151 = n13792 & n48150 ;
  assign n48152 = \m0_data_i[19]_pad  & n13767 ;
  assign n48153 = n13760 & n48152 ;
  assign n48154 = ~n48151 & ~n48153 ;
  assign n48155 = \m3_data_i[19]_pad  & ~n13767 ;
  assign n48156 = n13775 & n48155 ;
  assign n48157 = \m4_data_i[19]_pad  & n13767 ;
  assign n48158 = n13792 & n48157 ;
  assign n48159 = ~n48156 & ~n48158 ;
  assign n48160 = n48154 & n48159 ;
  assign n48161 = n48149 & n48160 ;
  assign n48162 = \m0_data_i[1]_pad  & n13767 ;
  assign n48163 = n13760 & n48162 ;
  assign n48164 = \m7_data_i[1]_pad  & ~n13767 ;
  assign n48165 = n13784 & n48164 ;
  assign n48166 = ~n48163 & ~n48165 ;
  assign n48167 = \m3_data_i[1]_pad  & ~n13767 ;
  assign n48168 = n13775 & n48167 ;
  assign n48169 = \m2_data_i[1]_pad  & n13767 ;
  assign n48170 = n13775 & n48169 ;
  assign n48171 = ~n48168 & ~n48170 ;
  assign n48172 = n48166 & n48171 ;
  assign n48173 = \m4_data_i[1]_pad  & n13767 ;
  assign n48174 = n13792 & n48173 ;
  assign n48175 = \m1_data_i[1]_pad  & ~n13767 ;
  assign n48176 = n13760 & n48175 ;
  assign n48177 = ~n48174 & ~n48176 ;
  assign n48178 = \m6_data_i[1]_pad  & n13767 ;
  assign n48179 = n13784 & n48178 ;
  assign n48180 = \m5_data_i[1]_pad  & ~n13767 ;
  assign n48181 = n13792 & n48180 ;
  assign n48182 = ~n48179 & ~n48181 ;
  assign n48183 = n48177 & n48182 ;
  assign n48184 = n48172 & n48183 ;
  assign n48185 = \m0_data_i[20]_pad  & n13767 ;
  assign n48186 = n13760 & n48185 ;
  assign n48187 = \m7_data_i[20]_pad  & ~n13767 ;
  assign n48188 = n13784 & n48187 ;
  assign n48189 = ~n48186 & ~n48188 ;
  assign n48190 = \m3_data_i[20]_pad  & ~n13767 ;
  assign n48191 = n13775 & n48190 ;
  assign n48192 = \m2_data_i[20]_pad  & n13767 ;
  assign n48193 = n13775 & n48192 ;
  assign n48194 = ~n48191 & ~n48193 ;
  assign n48195 = n48189 & n48194 ;
  assign n48196 = \m4_data_i[20]_pad  & n13767 ;
  assign n48197 = n13792 & n48196 ;
  assign n48198 = \m1_data_i[20]_pad  & ~n13767 ;
  assign n48199 = n13760 & n48198 ;
  assign n48200 = ~n48197 & ~n48199 ;
  assign n48201 = \m6_data_i[20]_pad  & n13767 ;
  assign n48202 = n13784 & n48201 ;
  assign n48203 = \m5_data_i[20]_pad  & ~n13767 ;
  assign n48204 = n13792 & n48203 ;
  assign n48205 = ~n48202 & ~n48204 ;
  assign n48206 = n48200 & n48205 ;
  assign n48207 = n48195 & n48206 ;
  assign n48208 = \m1_data_i[21]_pad  & ~n13767 ;
  assign n48209 = n13760 & n48208 ;
  assign n48210 = \m2_data_i[21]_pad  & n13767 ;
  assign n48211 = n13775 & n48210 ;
  assign n48212 = ~n48209 & ~n48211 ;
  assign n48213 = \m3_data_i[21]_pad  & ~n13767 ;
  assign n48214 = n13775 & n48213 ;
  assign n48215 = \m7_data_i[21]_pad  & ~n13767 ;
  assign n48216 = n13784 & n48215 ;
  assign n48217 = ~n48214 & ~n48216 ;
  assign n48218 = n48212 & n48217 ;
  assign n48219 = \m4_data_i[21]_pad  & n13767 ;
  assign n48220 = n13792 & n48219 ;
  assign n48221 = \m0_data_i[21]_pad  & n13767 ;
  assign n48222 = n13760 & n48221 ;
  assign n48223 = ~n48220 & ~n48222 ;
  assign n48224 = \m6_data_i[21]_pad  & n13767 ;
  assign n48225 = n13784 & n48224 ;
  assign n48226 = \m5_data_i[21]_pad  & ~n13767 ;
  assign n48227 = n13792 & n48226 ;
  assign n48228 = ~n48225 & ~n48227 ;
  assign n48229 = n48223 & n48228 ;
  assign n48230 = n48218 & n48229 ;
  assign n48231 = \m1_data_i[22]_pad  & ~n13767 ;
  assign n48232 = n13760 & n48231 ;
  assign n48233 = \m2_data_i[22]_pad  & n13767 ;
  assign n48234 = n13775 & n48233 ;
  assign n48235 = ~n48232 & ~n48234 ;
  assign n48236 = \m6_data_i[22]_pad  & n13767 ;
  assign n48237 = n13784 & n48236 ;
  assign n48238 = \m7_data_i[22]_pad  & ~n13767 ;
  assign n48239 = n13784 & n48238 ;
  assign n48240 = ~n48237 & ~n48239 ;
  assign n48241 = n48235 & n48240 ;
  assign n48242 = \m5_data_i[22]_pad  & ~n13767 ;
  assign n48243 = n13792 & n48242 ;
  assign n48244 = \m0_data_i[22]_pad  & n13767 ;
  assign n48245 = n13760 & n48244 ;
  assign n48246 = ~n48243 & ~n48245 ;
  assign n48247 = \m3_data_i[22]_pad  & ~n13767 ;
  assign n48248 = n13775 & n48247 ;
  assign n48249 = \m4_data_i[22]_pad  & n13767 ;
  assign n48250 = n13792 & n48249 ;
  assign n48251 = ~n48248 & ~n48250 ;
  assign n48252 = n48246 & n48251 ;
  assign n48253 = n48241 & n48252 ;
  assign n48254 = \m3_data_i[23]_pad  & ~n13767 ;
  assign n48255 = n13775 & n48254 ;
  assign n48256 = \m4_data_i[23]_pad  & n13767 ;
  assign n48257 = n13792 & n48256 ;
  assign n48258 = ~n48255 & ~n48257 ;
  assign n48259 = \m6_data_i[23]_pad  & n13767 ;
  assign n48260 = n13784 & n48259 ;
  assign n48261 = \m2_data_i[23]_pad  & n13767 ;
  assign n48262 = n13775 & n48261 ;
  assign n48263 = ~n48260 & ~n48262 ;
  assign n48264 = n48258 & n48263 ;
  assign n48265 = \m5_data_i[23]_pad  & ~n13767 ;
  assign n48266 = n13792 & n48265 ;
  assign n48267 = \m1_data_i[23]_pad  & ~n13767 ;
  assign n48268 = n13760 & n48267 ;
  assign n48269 = ~n48266 & ~n48268 ;
  assign n48270 = \m0_data_i[23]_pad  & n13767 ;
  assign n48271 = n13760 & n48270 ;
  assign n48272 = \m7_data_i[23]_pad  & ~n13767 ;
  assign n48273 = n13784 & n48272 ;
  assign n48274 = ~n48271 & ~n48273 ;
  assign n48275 = n48269 & n48274 ;
  assign n48276 = n48264 & n48275 ;
  assign n48277 = \m1_data_i[24]_pad  & ~n13767 ;
  assign n48278 = n13760 & n48277 ;
  assign n48279 = \m2_data_i[24]_pad  & n13767 ;
  assign n48280 = n13775 & n48279 ;
  assign n48281 = ~n48278 & ~n48280 ;
  assign n48282 = \m3_data_i[24]_pad  & ~n13767 ;
  assign n48283 = n13775 & n48282 ;
  assign n48284 = \m7_data_i[24]_pad  & ~n13767 ;
  assign n48285 = n13784 & n48284 ;
  assign n48286 = ~n48283 & ~n48285 ;
  assign n48287 = n48281 & n48286 ;
  assign n48288 = \m4_data_i[24]_pad  & n13767 ;
  assign n48289 = n13792 & n48288 ;
  assign n48290 = \m0_data_i[24]_pad  & n13767 ;
  assign n48291 = n13760 & n48290 ;
  assign n48292 = ~n48289 & ~n48291 ;
  assign n48293 = \m6_data_i[24]_pad  & n13767 ;
  assign n48294 = n13784 & n48293 ;
  assign n48295 = \m5_data_i[24]_pad  & ~n13767 ;
  assign n48296 = n13792 & n48295 ;
  assign n48297 = ~n48294 & ~n48296 ;
  assign n48298 = n48292 & n48297 ;
  assign n48299 = n48287 & n48298 ;
  assign n48300 = \m3_data_i[25]_pad  & ~n13767 ;
  assign n48301 = n13775 & n48300 ;
  assign n48302 = \m4_data_i[25]_pad  & n13767 ;
  assign n48303 = n13792 & n48302 ;
  assign n48304 = ~n48301 & ~n48303 ;
  assign n48305 = \m6_data_i[25]_pad  & n13767 ;
  assign n48306 = n13784 & n48305 ;
  assign n48307 = \m7_data_i[25]_pad  & ~n13767 ;
  assign n48308 = n13784 & n48307 ;
  assign n48309 = ~n48306 & ~n48308 ;
  assign n48310 = n48304 & n48309 ;
  assign n48311 = \m5_data_i[25]_pad  & ~n13767 ;
  assign n48312 = n13792 & n48311 ;
  assign n48313 = \m0_data_i[25]_pad  & n13767 ;
  assign n48314 = n13760 & n48313 ;
  assign n48315 = ~n48312 & ~n48314 ;
  assign n48316 = \m1_data_i[25]_pad  & ~n13767 ;
  assign n48317 = n13760 & n48316 ;
  assign n48318 = \m2_data_i[25]_pad  & n13767 ;
  assign n48319 = n13775 & n48318 ;
  assign n48320 = ~n48317 & ~n48319 ;
  assign n48321 = n48315 & n48320 ;
  assign n48322 = n48310 & n48321 ;
  assign n48323 = \m0_data_i[26]_pad  & n13767 ;
  assign n48324 = n13760 & n48323 ;
  assign n48325 = \m7_data_i[26]_pad  & ~n13767 ;
  assign n48326 = n13784 & n48325 ;
  assign n48327 = ~n48324 & ~n48326 ;
  assign n48328 = \m3_data_i[26]_pad  & ~n13767 ;
  assign n48329 = n13775 & n48328 ;
  assign n48330 = \m2_data_i[26]_pad  & n13767 ;
  assign n48331 = n13775 & n48330 ;
  assign n48332 = ~n48329 & ~n48331 ;
  assign n48333 = n48327 & n48332 ;
  assign n48334 = \m4_data_i[26]_pad  & n13767 ;
  assign n48335 = n13792 & n48334 ;
  assign n48336 = \m1_data_i[26]_pad  & ~n13767 ;
  assign n48337 = n13760 & n48336 ;
  assign n48338 = ~n48335 & ~n48337 ;
  assign n48339 = \m6_data_i[26]_pad  & n13767 ;
  assign n48340 = n13784 & n48339 ;
  assign n48341 = \m5_data_i[26]_pad  & ~n13767 ;
  assign n48342 = n13792 & n48341 ;
  assign n48343 = ~n48340 & ~n48342 ;
  assign n48344 = n48338 & n48343 ;
  assign n48345 = n48333 & n48344 ;
  assign n48346 = \m3_data_i[27]_pad  & ~n13767 ;
  assign n48347 = n13775 & n48346 ;
  assign n48348 = \m4_data_i[27]_pad  & n13767 ;
  assign n48349 = n13792 & n48348 ;
  assign n48350 = ~n48347 & ~n48349 ;
  assign n48351 = \m6_data_i[27]_pad  & n13767 ;
  assign n48352 = n13784 & n48351 ;
  assign n48353 = \m2_data_i[27]_pad  & n13767 ;
  assign n48354 = n13775 & n48353 ;
  assign n48355 = ~n48352 & ~n48354 ;
  assign n48356 = n48350 & n48355 ;
  assign n48357 = \m5_data_i[27]_pad  & ~n13767 ;
  assign n48358 = n13792 & n48357 ;
  assign n48359 = \m1_data_i[27]_pad  & ~n13767 ;
  assign n48360 = n13760 & n48359 ;
  assign n48361 = ~n48358 & ~n48360 ;
  assign n48362 = \m0_data_i[27]_pad  & n13767 ;
  assign n48363 = n13760 & n48362 ;
  assign n48364 = \m7_data_i[27]_pad  & ~n13767 ;
  assign n48365 = n13784 & n48364 ;
  assign n48366 = ~n48363 & ~n48365 ;
  assign n48367 = n48361 & n48366 ;
  assign n48368 = n48356 & n48367 ;
  assign n48369 = \m1_data_i[28]_pad  & ~n13767 ;
  assign n48370 = n13760 & n48369 ;
  assign n48371 = \m2_data_i[28]_pad  & n13767 ;
  assign n48372 = n13775 & n48371 ;
  assign n48373 = ~n48370 & ~n48372 ;
  assign n48374 = \m6_data_i[28]_pad  & n13767 ;
  assign n48375 = n13784 & n48374 ;
  assign n48376 = \m7_data_i[28]_pad  & ~n13767 ;
  assign n48377 = n13784 & n48376 ;
  assign n48378 = ~n48375 & ~n48377 ;
  assign n48379 = n48373 & n48378 ;
  assign n48380 = \m5_data_i[28]_pad  & ~n13767 ;
  assign n48381 = n13792 & n48380 ;
  assign n48382 = \m0_data_i[28]_pad  & n13767 ;
  assign n48383 = n13760 & n48382 ;
  assign n48384 = ~n48381 & ~n48383 ;
  assign n48385 = \m3_data_i[28]_pad  & ~n13767 ;
  assign n48386 = n13775 & n48385 ;
  assign n48387 = \m4_data_i[28]_pad  & n13767 ;
  assign n48388 = n13792 & n48387 ;
  assign n48389 = ~n48386 & ~n48388 ;
  assign n48390 = n48384 & n48389 ;
  assign n48391 = n48379 & n48390 ;
  assign n48392 = \m3_data_i[29]_pad  & ~n13767 ;
  assign n48393 = n13775 & n48392 ;
  assign n48394 = \m4_data_i[29]_pad  & n13767 ;
  assign n48395 = n13792 & n48394 ;
  assign n48396 = ~n48393 & ~n48395 ;
  assign n48397 = \m6_data_i[29]_pad  & n13767 ;
  assign n48398 = n13784 & n48397 ;
  assign n48399 = \m2_data_i[29]_pad  & n13767 ;
  assign n48400 = n13775 & n48399 ;
  assign n48401 = ~n48398 & ~n48400 ;
  assign n48402 = n48396 & n48401 ;
  assign n48403 = \m5_data_i[29]_pad  & ~n13767 ;
  assign n48404 = n13792 & n48403 ;
  assign n48405 = \m1_data_i[29]_pad  & ~n13767 ;
  assign n48406 = n13760 & n48405 ;
  assign n48407 = ~n48404 & ~n48406 ;
  assign n48408 = \m0_data_i[29]_pad  & n13767 ;
  assign n48409 = n13760 & n48408 ;
  assign n48410 = \m7_data_i[29]_pad  & ~n13767 ;
  assign n48411 = n13784 & n48410 ;
  assign n48412 = ~n48409 & ~n48411 ;
  assign n48413 = n48407 & n48412 ;
  assign n48414 = n48402 & n48413 ;
  assign n48415 = \m3_data_i[2]_pad  & ~n13767 ;
  assign n48416 = n13775 & n48415 ;
  assign n48417 = \m4_data_i[2]_pad  & n13767 ;
  assign n48418 = n13792 & n48417 ;
  assign n48419 = ~n48416 & ~n48418 ;
  assign n48420 = \m6_data_i[2]_pad  & n13767 ;
  assign n48421 = n13784 & n48420 ;
  assign n48422 = \m2_data_i[2]_pad  & n13767 ;
  assign n48423 = n13775 & n48422 ;
  assign n48424 = ~n48421 & ~n48423 ;
  assign n48425 = n48419 & n48424 ;
  assign n48426 = \m5_data_i[2]_pad  & ~n13767 ;
  assign n48427 = n13792 & n48426 ;
  assign n48428 = \m1_data_i[2]_pad  & ~n13767 ;
  assign n48429 = n13760 & n48428 ;
  assign n48430 = ~n48427 & ~n48429 ;
  assign n48431 = \m0_data_i[2]_pad  & n13767 ;
  assign n48432 = n13760 & n48431 ;
  assign n48433 = \m7_data_i[2]_pad  & ~n13767 ;
  assign n48434 = n13784 & n48433 ;
  assign n48435 = ~n48432 & ~n48434 ;
  assign n48436 = n48430 & n48435 ;
  assign n48437 = n48425 & n48436 ;
  assign n48438 = \m0_data_i[30]_pad  & n13767 ;
  assign n48439 = n13760 & n48438 ;
  assign n48440 = \m7_data_i[30]_pad  & ~n13767 ;
  assign n48441 = n13784 & n48440 ;
  assign n48442 = ~n48439 & ~n48441 ;
  assign n48443 = \m3_data_i[30]_pad  & ~n13767 ;
  assign n48444 = n13775 & n48443 ;
  assign n48445 = \m5_data_i[30]_pad  & ~n13767 ;
  assign n48446 = n13792 & n48445 ;
  assign n48447 = ~n48444 & ~n48446 ;
  assign n48448 = n48442 & n48447 ;
  assign n48449 = \m4_data_i[30]_pad  & n13767 ;
  assign n48450 = n13792 & n48449 ;
  assign n48451 = \m6_data_i[30]_pad  & n13767 ;
  assign n48452 = n13784 & n48451 ;
  assign n48453 = ~n48450 & ~n48452 ;
  assign n48454 = \m1_data_i[30]_pad  & ~n13767 ;
  assign n48455 = n13760 & n48454 ;
  assign n48456 = \m2_data_i[30]_pad  & n13767 ;
  assign n48457 = n13775 & n48456 ;
  assign n48458 = ~n48455 & ~n48457 ;
  assign n48459 = n48453 & n48458 ;
  assign n48460 = n48448 & n48459 ;
  assign n48461 = \m1_data_i[31]_pad  & ~n13767 ;
  assign n48462 = n13760 & n48461 ;
  assign n48463 = \m2_data_i[31]_pad  & n13767 ;
  assign n48464 = n13775 & n48463 ;
  assign n48465 = ~n48462 & ~n48464 ;
  assign n48466 = \m3_data_i[31]_pad  & ~n13767 ;
  assign n48467 = n13775 & n48466 ;
  assign n48468 = \m7_data_i[31]_pad  & ~n13767 ;
  assign n48469 = n13784 & n48468 ;
  assign n48470 = ~n48467 & ~n48469 ;
  assign n48471 = n48465 & n48470 ;
  assign n48472 = \m4_data_i[31]_pad  & n13767 ;
  assign n48473 = n13792 & n48472 ;
  assign n48474 = \m0_data_i[31]_pad  & n13767 ;
  assign n48475 = n13760 & n48474 ;
  assign n48476 = ~n48473 & ~n48475 ;
  assign n48477 = \m6_data_i[31]_pad  & n13767 ;
  assign n48478 = n13784 & n48477 ;
  assign n48479 = \m5_data_i[31]_pad  & ~n13767 ;
  assign n48480 = n13792 & n48479 ;
  assign n48481 = ~n48478 & ~n48480 ;
  assign n48482 = n48476 & n48481 ;
  assign n48483 = n48471 & n48482 ;
  assign n48484 = \m1_data_i[3]_pad  & ~n13767 ;
  assign n48485 = n13760 & n48484 ;
  assign n48486 = \m2_data_i[3]_pad  & n13767 ;
  assign n48487 = n13775 & n48486 ;
  assign n48488 = ~n48485 & ~n48487 ;
  assign n48489 = \m6_data_i[3]_pad  & n13767 ;
  assign n48490 = n13784 & n48489 ;
  assign n48491 = \m7_data_i[3]_pad  & ~n13767 ;
  assign n48492 = n13784 & n48491 ;
  assign n48493 = ~n48490 & ~n48492 ;
  assign n48494 = n48488 & n48493 ;
  assign n48495 = \m5_data_i[3]_pad  & ~n13767 ;
  assign n48496 = n13792 & n48495 ;
  assign n48497 = \m0_data_i[3]_pad  & n13767 ;
  assign n48498 = n13760 & n48497 ;
  assign n48499 = ~n48496 & ~n48498 ;
  assign n48500 = \m3_data_i[3]_pad  & ~n13767 ;
  assign n48501 = n13775 & n48500 ;
  assign n48502 = \m4_data_i[3]_pad  & n13767 ;
  assign n48503 = n13792 & n48502 ;
  assign n48504 = ~n48501 & ~n48503 ;
  assign n48505 = n48499 & n48504 ;
  assign n48506 = n48494 & n48505 ;
  assign n48507 = \m0_data_i[4]_pad  & n13767 ;
  assign n48508 = n13760 & n48507 ;
  assign n48509 = \m7_data_i[4]_pad  & ~n13767 ;
  assign n48510 = n13784 & n48509 ;
  assign n48511 = ~n48508 & ~n48510 ;
  assign n48512 = \m3_data_i[4]_pad  & ~n13767 ;
  assign n48513 = n13775 & n48512 ;
  assign n48514 = \m2_data_i[4]_pad  & n13767 ;
  assign n48515 = n13775 & n48514 ;
  assign n48516 = ~n48513 & ~n48515 ;
  assign n48517 = n48511 & n48516 ;
  assign n48518 = \m4_data_i[4]_pad  & n13767 ;
  assign n48519 = n13792 & n48518 ;
  assign n48520 = \m1_data_i[4]_pad  & ~n13767 ;
  assign n48521 = n13760 & n48520 ;
  assign n48522 = ~n48519 & ~n48521 ;
  assign n48523 = \m6_data_i[4]_pad  & n13767 ;
  assign n48524 = n13784 & n48523 ;
  assign n48525 = \m5_data_i[4]_pad  & ~n13767 ;
  assign n48526 = n13792 & n48525 ;
  assign n48527 = ~n48524 & ~n48526 ;
  assign n48528 = n48522 & n48527 ;
  assign n48529 = n48517 & n48528 ;
  assign n48530 = \m3_data_i[5]_pad  & ~n13767 ;
  assign n48531 = n13775 & n48530 ;
  assign n48532 = \m4_data_i[5]_pad  & n13767 ;
  assign n48533 = n13792 & n48532 ;
  assign n48534 = ~n48531 & ~n48533 ;
  assign n48535 = \m6_data_i[5]_pad  & n13767 ;
  assign n48536 = n13784 & n48535 ;
  assign n48537 = \m2_data_i[5]_pad  & n13767 ;
  assign n48538 = n13775 & n48537 ;
  assign n48539 = ~n48536 & ~n48538 ;
  assign n48540 = n48534 & n48539 ;
  assign n48541 = \m5_data_i[5]_pad  & ~n13767 ;
  assign n48542 = n13792 & n48541 ;
  assign n48543 = \m1_data_i[5]_pad  & ~n13767 ;
  assign n48544 = n13760 & n48543 ;
  assign n48545 = ~n48542 & ~n48544 ;
  assign n48546 = \m0_data_i[5]_pad  & n13767 ;
  assign n48547 = n13760 & n48546 ;
  assign n48548 = \m7_data_i[5]_pad  & ~n13767 ;
  assign n48549 = n13784 & n48548 ;
  assign n48550 = ~n48547 & ~n48549 ;
  assign n48551 = n48545 & n48550 ;
  assign n48552 = n48540 & n48551 ;
  assign n48553 = \m3_data_i[6]_pad  & ~n13767 ;
  assign n48554 = n13775 & n48553 ;
  assign n48555 = \m4_data_i[6]_pad  & n13767 ;
  assign n48556 = n13792 & n48555 ;
  assign n48557 = ~n48554 & ~n48556 ;
  assign n48558 = \m6_data_i[6]_pad  & n13767 ;
  assign n48559 = n13784 & n48558 ;
  assign n48560 = \m7_data_i[6]_pad  & ~n13767 ;
  assign n48561 = n13784 & n48560 ;
  assign n48562 = ~n48559 & ~n48561 ;
  assign n48563 = n48557 & n48562 ;
  assign n48564 = \m5_data_i[6]_pad  & ~n13767 ;
  assign n48565 = n13792 & n48564 ;
  assign n48566 = \m0_data_i[6]_pad  & n13767 ;
  assign n48567 = n13760 & n48566 ;
  assign n48568 = ~n48565 & ~n48567 ;
  assign n48569 = \m1_data_i[6]_pad  & ~n13767 ;
  assign n48570 = n13760 & n48569 ;
  assign n48571 = \m2_data_i[6]_pad  & n13767 ;
  assign n48572 = n13775 & n48571 ;
  assign n48573 = ~n48570 & ~n48572 ;
  assign n48574 = n48568 & n48573 ;
  assign n48575 = n48563 & n48574 ;
  assign n48576 = \m3_data_i[7]_pad  & ~n13767 ;
  assign n48577 = n13775 & n48576 ;
  assign n48578 = \m4_data_i[7]_pad  & n13767 ;
  assign n48579 = n13792 & n48578 ;
  assign n48580 = ~n48577 & ~n48579 ;
  assign n48581 = \m6_data_i[7]_pad  & n13767 ;
  assign n48582 = n13784 & n48581 ;
  assign n48583 = \m2_data_i[7]_pad  & n13767 ;
  assign n48584 = n13775 & n48583 ;
  assign n48585 = ~n48582 & ~n48584 ;
  assign n48586 = n48580 & n48585 ;
  assign n48587 = \m5_data_i[7]_pad  & ~n13767 ;
  assign n48588 = n13792 & n48587 ;
  assign n48589 = \m1_data_i[7]_pad  & ~n13767 ;
  assign n48590 = n13760 & n48589 ;
  assign n48591 = ~n48588 & ~n48590 ;
  assign n48592 = \m0_data_i[7]_pad  & n13767 ;
  assign n48593 = n13760 & n48592 ;
  assign n48594 = \m7_data_i[7]_pad  & ~n13767 ;
  assign n48595 = n13784 & n48594 ;
  assign n48596 = ~n48593 & ~n48595 ;
  assign n48597 = n48591 & n48596 ;
  assign n48598 = n48586 & n48597 ;
  assign n48599 = \m1_data_i[8]_pad  & ~n13767 ;
  assign n48600 = n13760 & n48599 ;
  assign n48601 = \m2_data_i[8]_pad  & n13767 ;
  assign n48602 = n13775 & n48601 ;
  assign n48603 = ~n48600 & ~n48602 ;
  assign n48604 = \m3_data_i[8]_pad  & ~n13767 ;
  assign n48605 = n13775 & n48604 ;
  assign n48606 = \m7_data_i[8]_pad  & ~n13767 ;
  assign n48607 = n13784 & n48606 ;
  assign n48608 = ~n48605 & ~n48607 ;
  assign n48609 = n48603 & n48608 ;
  assign n48610 = \m4_data_i[8]_pad  & n13767 ;
  assign n48611 = n13792 & n48610 ;
  assign n48612 = \m0_data_i[8]_pad  & n13767 ;
  assign n48613 = n13760 & n48612 ;
  assign n48614 = ~n48611 & ~n48613 ;
  assign n48615 = \m6_data_i[8]_pad  & n13767 ;
  assign n48616 = n13784 & n48615 ;
  assign n48617 = \m5_data_i[8]_pad  & ~n13767 ;
  assign n48618 = n13792 & n48617 ;
  assign n48619 = ~n48616 & ~n48618 ;
  assign n48620 = n48614 & n48619 ;
  assign n48621 = n48609 & n48620 ;
  assign n48622 = \m3_data_i[9]_pad  & ~n13767 ;
  assign n48623 = n13775 & n48622 ;
  assign n48624 = \m4_data_i[9]_pad  & n13767 ;
  assign n48625 = n13792 & n48624 ;
  assign n48626 = ~n48623 & ~n48625 ;
  assign n48627 = \m6_data_i[9]_pad  & n13767 ;
  assign n48628 = n13784 & n48627 ;
  assign n48629 = \m7_data_i[9]_pad  & ~n13767 ;
  assign n48630 = n13784 & n48629 ;
  assign n48631 = ~n48628 & ~n48630 ;
  assign n48632 = n48626 & n48631 ;
  assign n48633 = \m5_data_i[9]_pad  & ~n13767 ;
  assign n48634 = n13792 & n48633 ;
  assign n48635 = \m0_data_i[9]_pad  & n13767 ;
  assign n48636 = n13760 & n48635 ;
  assign n48637 = ~n48634 & ~n48636 ;
  assign n48638 = \m1_data_i[9]_pad  & ~n13767 ;
  assign n48639 = n13760 & n48638 ;
  assign n48640 = \m2_data_i[9]_pad  & n13767 ;
  assign n48641 = n13775 & n48640 ;
  assign n48642 = ~n48639 & ~n48641 ;
  assign n48643 = n48637 & n48642 ;
  assign n48644 = n48632 & n48643 ;
  assign n48645 = \m1_sel_i[0]_pad  & ~n13767 ;
  assign n48646 = n13760 & n48645 ;
  assign n48647 = \m2_sel_i[0]_pad  & n13767 ;
  assign n48648 = n13775 & n48647 ;
  assign n48649 = ~n48646 & ~n48648 ;
  assign n48650 = \m6_sel_i[0]_pad  & n13767 ;
  assign n48651 = n13784 & n48650 ;
  assign n48652 = \m7_sel_i[0]_pad  & ~n13767 ;
  assign n48653 = n13784 & n48652 ;
  assign n48654 = ~n48651 & ~n48653 ;
  assign n48655 = n48649 & n48654 ;
  assign n48656 = \m5_sel_i[0]_pad  & ~n13767 ;
  assign n48657 = n13792 & n48656 ;
  assign n48658 = \m0_sel_i[0]_pad  & n13767 ;
  assign n48659 = n13760 & n48658 ;
  assign n48660 = ~n48657 & ~n48659 ;
  assign n48661 = \m3_sel_i[0]_pad  & ~n13767 ;
  assign n48662 = n13775 & n48661 ;
  assign n48663 = \m4_sel_i[0]_pad  & n13767 ;
  assign n48664 = n13792 & n48663 ;
  assign n48665 = ~n48662 & ~n48664 ;
  assign n48666 = n48660 & n48665 ;
  assign n48667 = n48655 & n48666 ;
  assign n48668 = \m3_sel_i[1]_pad  & ~n13767 ;
  assign n48669 = n13775 & n48668 ;
  assign n48670 = \m4_sel_i[1]_pad  & n13767 ;
  assign n48671 = n13792 & n48670 ;
  assign n48672 = ~n48669 & ~n48671 ;
  assign n48673 = \m6_sel_i[1]_pad  & n13767 ;
  assign n48674 = n13784 & n48673 ;
  assign n48675 = \m7_sel_i[1]_pad  & ~n13767 ;
  assign n48676 = n13784 & n48675 ;
  assign n48677 = ~n48674 & ~n48676 ;
  assign n48678 = n48672 & n48677 ;
  assign n48679 = \m5_sel_i[1]_pad  & ~n13767 ;
  assign n48680 = n13792 & n48679 ;
  assign n48681 = \m0_sel_i[1]_pad  & n13767 ;
  assign n48682 = n13760 & n48681 ;
  assign n48683 = ~n48680 & ~n48682 ;
  assign n48684 = \m1_sel_i[1]_pad  & ~n13767 ;
  assign n48685 = n13760 & n48684 ;
  assign n48686 = \m2_sel_i[1]_pad  & n13767 ;
  assign n48687 = n13775 & n48686 ;
  assign n48688 = ~n48685 & ~n48687 ;
  assign n48689 = n48683 & n48688 ;
  assign n48690 = n48678 & n48689 ;
  assign n48691 = \m0_sel_i[2]_pad  & n13767 ;
  assign n48692 = n13760 & n48691 ;
  assign n48693 = \m7_sel_i[2]_pad  & ~n13767 ;
  assign n48694 = n13784 & n48693 ;
  assign n48695 = ~n48692 & ~n48694 ;
  assign n48696 = \m3_sel_i[2]_pad  & ~n13767 ;
  assign n48697 = n13775 & n48696 ;
  assign n48698 = \m2_sel_i[2]_pad  & n13767 ;
  assign n48699 = n13775 & n48698 ;
  assign n48700 = ~n48697 & ~n48699 ;
  assign n48701 = n48695 & n48700 ;
  assign n48702 = \m4_sel_i[2]_pad  & n13767 ;
  assign n48703 = n13792 & n48702 ;
  assign n48704 = \m1_sel_i[2]_pad  & ~n13767 ;
  assign n48705 = n13760 & n48704 ;
  assign n48706 = ~n48703 & ~n48705 ;
  assign n48707 = \m6_sel_i[2]_pad  & n13767 ;
  assign n48708 = n13784 & n48707 ;
  assign n48709 = \m5_sel_i[2]_pad  & ~n13767 ;
  assign n48710 = n13792 & n48709 ;
  assign n48711 = ~n48708 & ~n48710 ;
  assign n48712 = n48706 & n48711 ;
  assign n48713 = n48701 & n48712 ;
  assign n48714 = \m1_sel_i[3]_pad  & ~n13767 ;
  assign n48715 = n13760 & n48714 ;
  assign n48716 = \m2_sel_i[3]_pad  & n13767 ;
  assign n48717 = n13775 & n48716 ;
  assign n48718 = ~n48715 & ~n48717 ;
  assign n48719 = \m3_sel_i[3]_pad  & ~n13767 ;
  assign n48720 = n13775 & n48719 ;
  assign n48721 = \m7_sel_i[3]_pad  & ~n13767 ;
  assign n48722 = n13784 & n48721 ;
  assign n48723 = ~n48720 & ~n48722 ;
  assign n48724 = n48718 & n48723 ;
  assign n48725 = \m4_sel_i[3]_pad  & n13767 ;
  assign n48726 = n13792 & n48725 ;
  assign n48727 = \m0_sel_i[3]_pad  & n13767 ;
  assign n48728 = n13760 & n48727 ;
  assign n48729 = ~n48726 & ~n48728 ;
  assign n48730 = \m6_sel_i[3]_pad  & n13767 ;
  assign n48731 = n13784 & n48730 ;
  assign n48732 = \m5_sel_i[3]_pad  & ~n13767 ;
  assign n48733 = n13792 & n48732 ;
  assign n48734 = ~n48731 & ~n48733 ;
  assign n48735 = n48729 & n48734 ;
  assign n48736 = n48724 & n48735 ;
  assign n48737 = \m5_stb_i_pad  & n14991 ;
  assign n48738 = ~n13767 & n48737 ;
  assign n48739 = n13792 & n48738 ;
  assign n48740 = \m4_stb_i_pad  & n14717 ;
  assign n48741 = n13767 & n48740 ;
  assign n48742 = n13792 & n48741 ;
  assign n48743 = ~n48739 & ~n48742 ;
  assign n48744 = \m6_stb_i_pad  & n14690 ;
  assign n48745 = n13767 & n48744 ;
  assign n48746 = n13784 & n48745 ;
  assign n48747 = \m1_stb_i_pad  & n14841 ;
  assign n48748 = ~n13767 & n48747 ;
  assign n48749 = n13760 & n48748 ;
  assign n48750 = ~n48746 & ~n48749 ;
  assign n48751 = n48743 & n48750 ;
  assign n48752 = \m7_stb_i_pad  & n15086 ;
  assign n48753 = ~n13767 & n48752 ;
  assign n48754 = n13784 & n48753 ;
  assign n48755 = \m3_stb_i_pad  & n14923 ;
  assign n48756 = ~n13767 & n48755 ;
  assign n48757 = n13775 & n48756 ;
  assign n48758 = ~n48754 & ~n48757 ;
  assign n48759 = \m2_stb_i_pad  & n15082 ;
  assign n48760 = n13767 & n48759 ;
  assign n48761 = n13775 & n48760 ;
  assign n48762 = \m0_stb_i_pad  & n14791 ;
  assign n48763 = n13767 & n48762 ;
  assign n48764 = n13760 & n48763 ;
  assign n48765 = ~n48761 & ~n48764 ;
  assign n48766 = n48758 & n48765 ;
  assign n48767 = n48751 & n48766 ;
  assign n48768 = \m6_we_i_pad  & n13767 ;
  assign n48769 = n13784 & n48768 ;
  assign n48770 = \m5_we_i_pad  & ~n13767 ;
  assign n48771 = n13792 & n48770 ;
  assign n48772 = ~n48769 & ~n48771 ;
  assign n48773 = \m3_we_i_pad  & ~n13767 ;
  assign n48774 = n13775 & n48773 ;
  assign n48775 = \m2_we_i_pad  & n13767 ;
  assign n48776 = n13775 & n48775 ;
  assign n48777 = ~n48774 & ~n48776 ;
  assign n48778 = n48772 & n48777 ;
  assign n48779 = \m4_we_i_pad  & n13767 ;
  assign n48780 = n13792 & n48779 ;
  assign n48781 = \m1_we_i_pad  & ~n13767 ;
  assign n48782 = n13760 & n48781 ;
  assign n48783 = ~n48780 & ~n48782 ;
  assign n48784 = \m0_we_i_pad  & n13767 ;
  assign n48785 = n13760 & n48784 ;
  assign n48786 = \m7_we_i_pad  & ~n13767 ;
  assign n48787 = n13784 & n48786 ;
  assign n48788 = ~n48785 & ~n48787 ;
  assign n48789 = n48783 & n48788 ;
  assign n48790 = n48778 & n48789 ;
  assign n48791 = \m3_addr_i[0]_pad  & ~n13847 ;
  assign n48792 = n13840 & n48791 ;
  assign n48793 = \m4_addr_i[0]_pad  & n13847 ;
  assign n48794 = n13872 & n48793 ;
  assign n48795 = ~n48792 & ~n48794 ;
  assign n48796 = \m6_addr_i[0]_pad  & n13847 ;
  assign n48797 = n13864 & n48796 ;
  assign n48798 = \m2_addr_i[0]_pad  & n13847 ;
  assign n48799 = n13840 & n48798 ;
  assign n48800 = ~n48797 & ~n48799 ;
  assign n48801 = n48795 & n48800 ;
  assign n48802 = \m5_addr_i[0]_pad  & ~n13847 ;
  assign n48803 = n13872 & n48802 ;
  assign n48804 = \m1_addr_i[0]_pad  & ~n13847 ;
  assign n48805 = n13855 & n48804 ;
  assign n48806 = ~n48803 & ~n48805 ;
  assign n48807 = \m0_addr_i[0]_pad  & n13847 ;
  assign n48808 = n13855 & n48807 ;
  assign n48809 = \m7_addr_i[0]_pad  & ~n13847 ;
  assign n48810 = n13864 & n48809 ;
  assign n48811 = ~n48808 & ~n48810 ;
  assign n48812 = n48806 & n48811 ;
  assign n48813 = n48801 & n48812 ;
  assign n48814 = \m3_addr_i[10]_pad  & ~n13847 ;
  assign n48815 = n13840 & n48814 ;
  assign n48816 = \m4_addr_i[10]_pad  & n13847 ;
  assign n48817 = n13872 & n48816 ;
  assign n48818 = ~n48815 & ~n48817 ;
  assign n48819 = \m1_addr_i[10]_pad  & ~n13847 ;
  assign n48820 = n13855 & n48819 ;
  assign n48821 = \m5_addr_i[10]_pad  & ~n13847 ;
  assign n48822 = n13872 & n48821 ;
  assign n48823 = ~n48820 & ~n48822 ;
  assign n48824 = n48818 & n48823 ;
  assign n48825 = \m2_addr_i[10]_pad  & n13847 ;
  assign n48826 = n13840 & n48825 ;
  assign n48827 = \m6_addr_i[10]_pad  & n13847 ;
  assign n48828 = n13864 & n48827 ;
  assign n48829 = ~n48826 & ~n48828 ;
  assign n48830 = \m0_addr_i[10]_pad  & n13847 ;
  assign n48831 = n13855 & n48830 ;
  assign n48832 = \m7_addr_i[10]_pad  & ~n13847 ;
  assign n48833 = n13864 & n48832 ;
  assign n48834 = ~n48831 & ~n48833 ;
  assign n48835 = n48829 & n48834 ;
  assign n48836 = n48824 & n48835 ;
  assign n48837 = \m3_addr_i[11]_pad  & ~n13847 ;
  assign n48838 = n13840 & n48837 ;
  assign n48839 = \m4_addr_i[11]_pad  & n13847 ;
  assign n48840 = n13872 & n48839 ;
  assign n48841 = ~n48838 & ~n48840 ;
  assign n48842 = \m1_addr_i[11]_pad  & ~n13847 ;
  assign n48843 = n13855 & n48842 ;
  assign n48844 = \m5_addr_i[11]_pad  & ~n13847 ;
  assign n48845 = n13872 & n48844 ;
  assign n48846 = ~n48843 & ~n48845 ;
  assign n48847 = n48841 & n48846 ;
  assign n48848 = \m2_addr_i[11]_pad  & n13847 ;
  assign n48849 = n13840 & n48848 ;
  assign n48850 = \m6_addr_i[11]_pad  & n13847 ;
  assign n48851 = n13864 & n48850 ;
  assign n48852 = ~n48849 & ~n48851 ;
  assign n48853 = \m0_addr_i[11]_pad  & n13847 ;
  assign n48854 = n13855 & n48853 ;
  assign n48855 = \m7_addr_i[11]_pad  & ~n13847 ;
  assign n48856 = n13864 & n48855 ;
  assign n48857 = ~n48854 & ~n48856 ;
  assign n48858 = n48852 & n48857 ;
  assign n48859 = n48847 & n48858 ;
  assign n48860 = \m1_addr_i[12]_pad  & ~n13847 ;
  assign n48861 = n13855 & n48860 ;
  assign n48862 = \m2_addr_i[12]_pad  & n13847 ;
  assign n48863 = n13840 & n48862 ;
  assign n48864 = ~n48861 & ~n48863 ;
  assign n48865 = \m0_addr_i[12]_pad  & n13847 ;
  assign n48866 = n13855 & n48865 ;
  assign n48867 = \m4_addr_i[12]_pad  & n13847 ;
  assign n48868 = n13872 & n48867 ;
  assign n48869 = ~n48866 & ~n48868 ;
  assign n48870 = n48864 & n48869 ;
  assign n48871 = \m7_addr_i[12]_pad  & ~n13847 ;
  assign n48872 = n13864 & n48871 ;
  assign n48873 = \m3_addr_i[12]_pad  & ~n13847 ;
  assign n48874 = n13840 & n48873 ;
  assign n48875 = ~n48872 & ~n48874 ;
  assign n48876 = \m6_addr_i[12]_pad  & n13847 ;
  assign n48877 = n13864 & n48876 ;
  assign n48878 = \m5_addr_i[12]_pad  & ~n13847 ;
  assign n48879 = n13872 & n48878 ;
  assign n48880 = ~n48877 & ~n48879 ;
  assign n48881 = n48875 & n48880 ;
  assign n48882 = n48870 & n48881 ;
  assign n48883 = \m0_addr_i[13]_pad  & n13847 ;
  assign n48884 = n13855 & n48883 ;
  assign n48885 = \m7_addr_i[13]_pad  & ~n13847 ;
  assign n48886 = n13864 & n48885 ;
  assign n48887 = ~n48884 & ~n48886 ;
  assign n48888 = \m1_addr_i[13]_pad  & ~n13847 ;
  assign n48889 = n13855 & n48888 ;
  assign n48890 = \m5_addr_i[13]_pad  & ~n13847 ;
  assign n48891 = n13872 & n48890 ;
  assign n48892 = ~n48889 & ~n48891 ;
  assign n48893 = n48887 & n48892 ;
  assign n48894 = \m2_addr_i[13]_pad  & n13847 ;
  assign n48895 = n13840 & n48894 ;
  assign n48896 = \m6_addr_i[13]_pad  & n13847 ;
  assign n48897 = n13864 & n48896 ;
  assign n48898 = ~n48895 & ~n48897 ;
  assign n48899 = \m3_addr_i[13]_pad  & ~n13847 ;
  assign n48900 = n13840 & n48899 ;
  assign n48901 = \m4_addr_i[13]_pad  & n13847 ;
  assign n48902 = n13872 & n48901 ;
  assign n48903 = ~n48900 & ~n48902 ;
  assign n48904 = n48898 & n48903 ;
  assign n48905 = n48893 & n48904 ;
  assign n48906 = \m6_addr_i[14]_pad  & n13847 ;
  assign n48907 = n13864 & n48906 ;
  assign n48908 = \m5_addr_i[14]_pad  & ~n13847 ;
  assign n48909 = n13872 & n48908 ;
  assign n48910 = ~n48907 & ~n48909 ;
  assign n48911 = \m3_addr_i[14]_pad  & ~n13847 ;
  assign n48912 = n13840 & n48911 ;
  assign n48913 = \m7_addr_i[14]_pad  & ~n13847 ;
  assign n48914 = n13864 & n48913 ;
  assign n48915 = ~n48912 & ~n48914 ;
  assign n48916 = n48910 & n48915 ;
  assign n48917 = \m4_addr_i[14]_pad  & n13847 ;
  assign n48918 = n13872 & n48917 ;
  assign n48919 = \m0_addr_i[14]_pad  & n13847 ;
  assign n48920 = n13855 & n48919 ;
  assign n48921 = ~n48918 & ~n48920 ;
  assign n48922 = \m1_addr_i[14]_pad  & ~n13847 ;
  assign n48923 = n13855 & n48922 ;
  assign n48924 = \m2_addr_i[14]_pad  & n13847 ;
  assign n48925 = n13840 & n48924 ;
  assign n48926 = ~n48923 & ~n48925 ;
  assign n48927 = n48921 & n48926 ;
  assign n48928 = n48916 & n48927 ;
  assign n48929 = \m1_addr_i[15]_pad  & ~n13847 ;
  assign n48930 = n13855 & n48929 ;
  assign n48931 = \m2_addr_i[15]_pad  & n13847 ;
  assign n48932 = n13840 & n48931 ;
  assign n48933 = ~n48930 & ~n48932 ;
  assign n48934 = \m0_addr_i[15]_pad  & n13847 ;
  assign n48935 = n13855 & n48934 ;
  assign n48936 = \m4_addr_i[15]_pad  & n13847 ;
  assign n48937 = n13872 & n48936 ;
  assign n48938 = ~n48935 & ~n48937 ;
  assign n48939 = n48933 & n48938 ;
  assign n48940 = \m7_addr_i[15]_pad  & ~n13847 ;
  assign n48941 = n13864 & n48940 ;
  assign n48942 = \m3_addr_i[15]_pad  & ~n13847 ;
  assign n48943 = n13840 & n48942 ;
  assign n48944 = ~n48941 & ~n48943 ;
  assign n48945 = \m6_addr_i[15]_pad  & n13847 ;
  assign n48946 = n13864 & n48945 ;
  assign n48947 = \m5_addr_i[15]_pad  & ~n13847 ;
  assign n48948 = n13872 & n48947 ;
  assign n48949 = ~n48946 & ~n48948 ;
  assign n48950 = n48944 & n48949 ;
  assign n48951 = n48939 & n48950 ;
  assign n48952 = \m1_addr_i[16]_pad  & ~n13847 ;
  assign n48953 = n13855 & n48952 ;
  assign n48954 = \m2_addr_i[16]_pad  & n13847 ;
  assign n48955 = n13840 & n48954 ;
  assign n48956 = ~n48953 & ~n48955 ;
  assign n48957 = \m0_addr_i[16]_pad  & n13847 ;
  assign n48958 = n13855 & n48957 ;
  assign n48959 = \m5_addr_i[16]_pad  & ~n13847 ;
  assign n48960 = n13872 & n48959 ;
  assign n48961 = ~n48958 & ~n48960 ;
  assign n48962 = n48956 & n48961 ;
  assign n48963 = \m7_addr_i[16]_pad  & ~n13847 ;
  assign n48964 = n13864 & n48963 ;
  assign n48965 = \m6_addr_i[16]_pad  & n13847 ;
  assign n48966 = n13864 & n48965 ;
  assign n48967 = ~n48964 & ~n48966 ;
  assign n48968 = \m3_addr_i[16]_pad  & ~n13847 ;
  assign n48969 = n13840 & n48968 ;
  assign n48970 = \m4_addr_i[16]_pad  & n13847 ;
  assign n48971 = n13872 & n48970 ;
  assign n48972 = ~n48969 & ~n48971 ;
  assign n48973 = n48967 & n48972 ;
  assign n48974 = n48962 & n48973 ;
  assign n48975 = \m1_addr_i[17]_pad  & ~n13847 ;
  assign n48976 = n13855 & n48975 ;
  assign n48977 = \m2_addr_i[17]_pad  & n13847 ;
  assign n48978 = n13840 & n48977 ;
  assign n48979 = ~n48976 & ~n48978 ;
  assign n48980 = \m0_addr_i[17]_pad  & n13847 ;
  assign n48981 = n13855 & n48980 ;
  assign n48982 = \m5_addr_i[17]_pad  & ~n13847 ;
  assign n48983 = n13872 & n48982 ;
  assign n48984 = ~n48981 & ~n48983 ;
  assign n48985 = n48979 & n48984 ;
  assign n48986 = \m7_addr_i[17]_pad  & ~n13847 ;
  assign n48987 = n13864 & n48986 ;
  assign n48988 = \m6_addr_i[17]_pad  & n13847 ;
  assign n48989 = n13864 & n48988 ;
  assign n48990 = ~n48987 & ~n48989 ;
  assign n48991 = \m3_addr_i[17]_pad  & ~n13847 ;
  assign n48992 = n13840 & n48991 ;
  assign n48993 = \m4_addr_i[17]_pad  & n13847 ;
  assign n48994 = n13872 & n48993 ;
  assign n48995 = ~n48992 & ~n48994 ;
  assign n48996 = n48990 & n48995 ;
  assign n48997 = n48985 & n48996 ;
  assign n48998 = \m6_addr_i[18]_pad  & n13847 ;
  assign n48999 = n13864 & n48998 ;
  assign n49000 = \m5_addr_i[18]_pad  & ~n13847 ;
  assign n49001 = n13872 & n49000 ;
  assign n49002 = ~n48999 & ~n49001 ;
  assign n49003 = \m1_addr_i[18]_pad  & ~n13847 ;
  assign n49004 = n13855 & n49003 ;
  assign n49005 = \m4_addr_i[18]_pad  & n13847 ;
  assign n49006 = n13872 & n49005 ;
  assign n49007 = ~n49004 & ~n49006 ;
  assign n49008 = n49002 & n49007 ;
  assign n49009 = \m2_addr_i[18]_pad  & n13847 ;
  assign n49010 = n13840 & n49009 ;
  assign n49011 = \m3_addr_i[18]_pad  & ~n13847 ;
  assign n49012 = n13840 & n49011 ;
  assign n49013 = ~n49010 & ~n49012 ;
  assign n49014 = \m0_addr_i[18]_pad  & n13847 ;
  assign n49015 = n13855 & n49014 ;
  assign n49016 = \m7_addr_i[18]_pad  & ~n13847 ;
  assign n49017 = n13864 & n49016 ;
  assign n49018 = ~n49015 & ~n49017 ;
  assign n49019 = n49013 & n49018 ;
  assign n49020 = n49008 & n49019 ;
  assign n49021 = \m3_addr_i[19]_pad  & ~n13847 ;
  assign n49022 = n13840 & n49021 ;
  assign n49023 = \m4_addr_i[19]_pad  & n13847 ;
  assign n49024 = n13872 & n49023 ;
  assign n49025 = ~n49022 & ~n49024 ;
  assign n49026 = \m0_addr_i[19]_pad  & n13847 ;
  assign n49027 = n13855 & n49026 ;
  assign n49028 = \m5_addr_i[19]_pad  & ~n13847 ;
  assign n49029 = n13872 & n49028 ;
  assign n49030 = ~n49027 & ~n49029 ;
  assign n49031 = n49025 & n49030 ;
  assign n49032 = \m7_addr_i[19]_pad  & ~n13847 ;
  assign n49033 = n13864 & n49032 ;
  assign n49034 = \m6_addr_i[19]_pad  & n13847 ;
  assign n49035 = n13864 & n49034 ;
  assign n49036 = ~n49033 & ~n49035 ;
  assign n49037 = \m1_addr_i[19]_pad  & ~n13847 ;
  assign n49038 = n13855 & n49037 ;
  assign n49039 = \m2_addr_i[19]_pad  & n13847 ;
  assign n49040 = n13840 & n49039 ;
  assign n49041 = ~n49038 & ~n49040 ;
  assign n49042 = n49036 & n49041 ;
  assign n49043 = n49031 & n49042 ;
  assign n49044 = \m3_addr_i[1]_pad  & ~n13847 ;
  assign n49045 = n13840 & n49044 ;
  assign n49046 = \m4_addr_i[1]_pad  & n13847 ;
  assign n49047 = n13872 & n49046 ;
  assign n49048 = ~n49045 & ~n49047 ;
  assign n49049 = \m6_addr_i[1]_pad  & n13847 ;
  assign n49050 = n13864 & n49049 ;
  assign n49051 = \m2_addr_i[1]_pad  & n13847 ;
  assign n49052 = n13840 & n49051 ;
  assign n49053 = ~n49050 & ~n49052 ;
  assign n49054 = n49048 & n49053 ;
  assign n49055 = \m5_addr_i[1]_pad  & ~n13847 ;
  assign n49056 = n13872 & n49055 ;
  assign n49057 = \m1_addr_i[1]_pad  & ~n13847 ;
  assign n49058 = n13855 & n49057 ;
  assign n49059 = ~n49056 & ~n49058 ;
  assign n49060 = \m0_addr_i[1]_pad  & n13847 ;
  assign n49061 = n13855 & n49060 ;
  assign n49062 = \m7_addr_i[1]_pad  & ~n13847 ;
  assign n49063 = n13864 & n49062 ;
  assign n49064 = ~n49061 & ~n49063 ;
  assign n49065 = n49059 & n49064 ;
  assign n49066 = n49054 & n49065 ;
  assign n49067 = \m0_addr_i[20]_pad  & n13847 ;
  assign n49068 = n13855 & n49067 ;
  assign n49069 = \m7_addr_i[20]_pad  & ~n13847 ;
  assign n49070 = n13864 & n49069 ;
  assign n49071 = ~n49068 & ~n49070 ;
  assign n49072 = \m1_addr_i[20]_pad  & ~n13847 ;
  assign n49073 = n13855 & n49072 ;
  assign n49074 = \m5_addr_i[20]_pad  & ~n13847 ;
  assign n49075 = n13872 & n49074 ;
  assign n49076 = ~n49073 & ~n49075 ;
  assign n49077 = n49071 & n49076 ;
  assign n49078 = \m2_addr_i[20]_pad  & n13847 ;
  assign n49079 = n13840 & n49078 ;
  assign n49080 = \m6_addr_i[20]_pad  & n13847 ;
  assign n49081 = n13864 & n49080 ;
  assign n49082 = ~n49079 & ~n49081 ;
  assign n49083 = \m3_addr_i[20]_pad  & ~n13847 ;
  assign n49084 = n13840 & n49083 ;
  assign n49085 = \m4_addr_i[20]_pad  & n13847 ;
  assign n49086 = n13872 & n49085 ;
  assign n49087 = ~n49084 & ~n49086 ;
  assign n49088 = n49082 & n49087 ;
  assign n49089 = n49077 & n49088 ;
  assign n49090 = \m6_addr_i[21]_pad  & n13847 ;
  assign n49091 = n13864 & n49090 ;
  assign n49092 = \m5_addr_i[21]_pad  & ~n13847 ;
  assign n49093 = n13872 & n49092 ;
  assign n49094 = ~n49091 & ~n49093 ;
  assign n49095 = \m3_addr_i[21]_pad  & ~n13847 ;
  assign n49096 = n13840 & n49095 ;
  assign n49097 = \m2_addr_i[21]_pad  & n13847 ;
  assign n49098 = n13840 & n49097 ;
  assign n49099 = ~n49096 & ~n49098 ;
  assign n49100 = n49094 & n49099 ;
  assign n49101 = \m4_addr_i[21]_pad  & n13847 ;
  assign n49102 = n13872 & n49101 ;
  assign n49103 = \m1_addr_i[21]_pad  & ~n13847 ;
  assign n49104 = n13855 & n49103 ;
  assign n49105 = ~n49102 & ~n49104 ;
  assign n49106 = \m0_addr_i[21]_pad  & n13847 ;
  assign n49107 = n13855 & n49106 ;
  assign n49108 = \m7_addr_i[21]_pad  & ~n13847 ;
  assign n49109 = n13864 & n49108 ;
  assign n49110 = ~n49107 & ~n49109 ;
  assign n49111 = n49105 & n49110 ;
  assign n49112 = n49100 & n49111 ;
  assign n49113 = \m1_addr_i[22]_pad  & ~n13847 ;
  assign n49114 = n13855 & n49113 ;
  assign n49115 = \m2_addr_i[22]_pad  & n13847 ;
  assign n49116 = n13840 & n49115 ;
  assign n49117 = ~n49114 & ~n49116 ;
  assign n49118 = \m0_addr_i[22]_pad  & n13847 ;
  assign n49119 = n13855 & n49118 ;
  assign n49120 = \m5_addr_i[22]_pad  & ~n13847 ;
  assign n49121 = n13872 & n49120 ;
  assign n49122 = ~n49119 & ~n49121 ;
  assign n49123 = n49117 & n49122 ;
  assign n49124 = \m7_addr_i[22]_pad  & ~n13847 ;
  assign n49125 = n13864 & n49124 ;
  assign n49126 = \m6_addr_i[22]_pad  & n13847 ;
  assign n49127 = n13864 & n49126 ;
  assign n49128 = ~n49125 & ~n49127 ;
  assign n49129 = \m3_addr_i[22]_pad  & ~n13847 ;
  assign n49130 = n13840 & n49129 ;
  assign n49131 = \m4_addr_i[22]_pad  & n13847 ;
  assign n49132 = n13872 & n49131 ;
  assign n49133 = ~n49130 & ~n49132 ;
  assign n49134 = n49128 & n49133 ;
  assign n49135 = n49123 & n49134 ;
  assign n49136 = \m6_addr_i[23]_pad  & n13847 ;
  assign n49137 = n13864 & n49136 ;
  assign n49138 = \m5_addr_i[23]_pad  & ~n13847 ;
  assign n49139 = n13872 & n49138 ;
  assign n49140 = ~n49137 & ~n49139 ;
  assign n49141 = \m3_addr_i[23]_pad  & ~n13847 ;
  assign n49142 = n13840 & n49141 ;
  assign n49143 = \m7_addr_i[23]_pad  & ~n13847 ;
  assign n49144 = n13864 & n49143 ;
  assign n49145 = ~n49142 & ~n49144 ;
  assign n49146 = n49140 & n49145 ;
  assign n49147 = \m4_addr_i[23]_pad  & n13847 ;
  assign n49148 = n13872 & n49147 ;
  assign n49149 = \m0_addr_i[23]_pad  & n13847 ;
  assign n49150 = n13855 & n49149 ;
  assign n49151 = ~n49148 & ~n49150 ;
  assign n49152 = \m1_addr_i[23]_pad  & ~n13847 ;
  assign n49153 = n13855 & n49152 ;
  assign n49154 = \m2_addr_i[23]_pad  & n13847 ;
  assign n49155 = n13840 & n49154 ;
  assign n49156 = ~n49153 & ~n49155 ;
  assign n49157 = n49151 & n49156 ;
  assign n49158 = n49146 & n49157 ;
  assign n49159 = \m0_addr_i[24]_pad  & n13847 ;
  assign n49160 = n13855 & n49159 ;
  assign n49161 = \m7_addr_i[24]_pad  & ~n13847 ;
  assign n49162 = n13864 & n49161 ;
  assign n49163 = ~n49160 & ~n49162 ;
  assign n49164 = \m1_addr_i[24]_pad  & ~n13847 ;
  assign n49165 = n13855 & n49164 ;
  assign n49166 = \m6_addr_i[24]_pad  & n13847 ;
  assign n49167 = n13864 & n49166 ;
  assign n49168 = ~n49165 & ~n49167 ;
  assign n49169 = n49163 & n49168 ;
  assign n49170 = \m2_addr_i[24]_pad  & n13847 ;
  assign n49171 = n13840 & n49170 ;
  assign n49172 = \m5_addr_i[24]_pad  & ~n13847 ;
  assign n49173 = n13872 & n49172 ;
  assign n49174 = ~n49171 & ~n49173 ;
  assign n49175 = \m3_addr_i[24]_pad  & ~n13847 ;
  assign n49176 = n13840 & n49175 ;
  assign n49177 = \m4_addr_i[24]_pad  & n13847 ;
  assign n49178 = n13872 & n49177 ;
  assign n49179 = ~n49176 & ~n49178 ;
  assign n49180 = n49174 & n49179 ;
  assign n49181 = n49169 & n49180 ;
  assign n49182 = \m0_addr_i[25]_pad  & n13847 ;
  assign n49183 = n13855 & n49182 ;
  assign n49184 = \m7_addr_i[25]_pad  & ~n13847 ;
  assign n49185 = n13864 & n49184 ;
  assign n49186 = ~n49183 & ~n49185 ;
  assign n49187 = \m5_addr_i[25]_pad  & ~n13847 ;
  assign n49188 = n13872 & n49187 ;
  assign n49189 = \m2_addr_i[25]_pad  & n13847 ;
  assign n49190 = n13840 & n49189 ;
  assign n49191 = ~n49188 & ~n49190 ;
  assign n49192 = n49186 & n49191 ;
  assign n49193 = \m6_addr_i[25]_pad  & n13847 ;
  assign n49194 = n13864 & n49193 ;
  assign n49195 = \m1_addr_i[25]_pad  & ~n13847 ;
  assign n49196 = n13855 & n49195 ;
  assign n49197 = ~n49194 & ~n49196 ;
  assign n49198 = \m3_addr_i[25]_pad  & ~n13847 ;
  assign n49199 = n13840 & n49198 ;
  assign n49200 = \m4_addr_i[25]_pad  & n13847 ;
  assign n49201 = n13872 & n49200 ;
  assign n49202 = ~n49199 & ~n49201 ;
  assign n49203 = n49197 & n49202 ;
  assign n49204 = n49192 & n49203 ;
  assign n49205 = \m1_addr_i[26]_pad  & ~n13847 ;
  assign n49206 = n13855 & n49205 ;
  assign n49207 = \m2_addr_i[26]_pad  & n13847 ;
  assign n49208 = n13840 & n49207 ;
  assign n49209 = ~n49206 & ~n49208 ;
  assign n49210 = \m5_addr_i[26]_pad  & ~n13847 ;
  assign n49211 = n13872 & n49210 ;
  assign n49212 = \m7_addr_i[26]_pad  & ~n13847 ;
  assign n49213 = n13864 & n49212 ;
  assign n49214 = ~n49211 & ~n49213 ;
  assign n49215 = n49209 & n49214 ;
  assign n49216 = \m6_addr_i[26]_pad  & n13847 ;
  assign n49217 = n13864 & n49216 ;
  assign n49218 = \m0_addr_i[26]_pad  & n13847 ;
  assign n49219 = n13855 & n49218 ;
  assign n49220 = ~n49217 & ~n49219 ;
  assign n49221 = \m3_addr_i[26]_pad  & ~n13847 ;
  assign n49222 = n13840 & n49221 ;
  assign n49223 = \m4_addr_i[26]_pad  & n13847 ;
  assign n49224 = n13872 & n49223 ;
  assign n49225 = ~n49222 & ~n49224 ;
  assign n49226 = n49220 & n49225 ;
  assign n49227 = n49215 & n49226 ;
  assign n49228 = \m1_addr_i[27]_pad  & ~n13847 ;
  assign n49229 = n13855 & n49228 ;
  assign n49230 = \m2_addr_i[27]_pad  & n13847 ;
  assign n49231 = n13840 & n49230 ;
  assign n49232 = ~n49229 & ~n49231 ;
  assign n49233 = \m3_addr_i[27]_pad  & ~n13847 ;
  assign n49234 = n13840 & n49233 ;
  assign n49235 = \m7_addr_i[27]_pad  & ~n13847 ;
  assign n49236 = n13864 & n49235 ;
  assign n49237 = ~n49234 & ~n49236 ;
  assign n49238 = n49232 & n49237 ;
  assign n49239 = \m4_addr_i[27]_pad  & n13847 ;
  assign n49240 = n13872 & n49239 ;
  assign n49241 = \m0_addr_i[27]_pad  & n13847 ;
  assign n49242 = n13855 & n49241 ;
  assign n49243 = ~n49240 & ~n49242 ;
  assign n49244 = \m5_addr_i[27]_pad  & ~n13847 ;
  assign n49245 = n13872 & n49244 ;
  assign n49246 = \m6_addr_i[27]_pad  & n13847 ;
  assign n49247 = n13864 & n49246 ;
  assign n49248 = ~n49245 & ~n49247 ;
  assign n49249 = n49243 & n49248 ;
  assign n49250 = n49238 & n49249 ;
  assign n49251 = \m5_addr_i[28]_pad  & ~n13847 ;
  assign n49252 = n13872 & n49251 ;
  assign n49253 = \m6_addr_i[28]_pad  & n13847 ;
  assign n49254 = n13864 & n49253 ;
  assign n49255 = ~n49252 & ~n49254 ;
  assign n49256 = \m3_addr_i[28]_pad  & ~n13847 ;
  assign n49257 = n13840 & n49256 ;
  assign n49258 = \m2_addr_i[28]_pad  & n13847 ;
  assign n49259 = n13840 & n49258 ;
  assign n49260 = ~n49257 & ~n49259 ;
  assign n49261 = n49255 & n49260 ;
  assign n49262 = \m4_addr_i[28]_pad  & n13847 ;
  assign n49263 = n13872 & n49262 ;
  assign n49264 = \m1_addr_i[28]_pad  & ~n13847 ;
  assign n49265 = n13855 & n49264 ;
  assign n49266 = ~n49263 & ~n49265 ;
  assign n49267 = \m0_addr_i[28]_pad  & n13847 ;
  assign n49268 = n13855 & n49267 ;
  assign n49269 = \m7_addr_i[28]_pad  & ~n13847 ;
  assign n49270 = n13864 & n49269 ;
  assign n49271 = ~n49268 & ~n49270 ;
  assign n49272 = n49266 & n49271 ;
  assign n49273 = n49261 & n49272 ;
  assign n49274 = \m1_addr_i[29]_pad  & ~n13847 ;
  assign n49275 = n13855 & n49274 ;
  assign n49276 = \m2_addr_i[29]_pad  & n13847 ;
  assign n49277 = n13840 & n49276 ;
  assign n49278 = ~n49275 & ~n49277 ;
  assign n49279 = \m5_addr_i[29]_pad  & ~n13847 ;
  assign n49280 = n13872 & n49279 ;
  assign n49281 = \m7_addr_i[29]_pad  & ~n13847 ;
  assign n49282 = n13864 & n49281 ;
  assign n49283 = ~n49280 & ~n49282 ;
  assign n49284 = n49278 & n49283 ;
  assign n49285 = \m6_addr_i[29]_pad  & n13847 ;
  assign n49286 = n13864 & n49285 ;
  assign n49287 = \m0_addr_i[29]_pad  & n13847 ;
  assign n49288 = n13855 & n49287 ;
  assign n49289 = ~n49286 & ~n49288 ;
  assign n49290 = \m3_addr_i[29]_pad  & ~n13847 ;
  assign n49291 = n13840 & n49290 ;
  assign n49292 = \m4_addr_i[29]_pad  & n13847 ;
  assign n49293 = n13872 & n49292 ;
  assign n49294 = ~n49291 & ~n49293 ;
  assign n49295 = n49289 & n49294 ;
  assign n49296 = n49284 & n49295 ;
  assign n49297 = \m3_addr_i[2]_pad  & ~n13847 ;
  assign n49298 = n13840 & n49297 ;
  assign n49299 = \m4_addr_i[2]_pad  & n13847 ;
  assign n49300 = n13872 & n49299 ;
  assign n49301 = ~n49298 & ~n49300 ;
  assign n49302 = \m6_addr_i[2]_pad  & n13847 ;
  assign n49303 = n13864 & n49302 ;
  assign n49304 = \m7_addr_i[2]_pad  & ~n13847 ;
  assign n49305 = n13864 & n49304 ;
  assign n49306 = ~n49303 & ~n49305 ;
  assign n49307 = n49301 & n49306 ;
  assign n49308 = \m5_addr_i[2]_pad  & ~n13847 ;
  assign n49309 = n13872 & n49308 ;
  assign n49310 = \m0_addr_i[2]_pad  & n13847 ;
  assign n49311 = n13855 & n49310 ;
  assign n49312 = ~n49309 & ~n49311 ;
  assign n49313 = \m1_addr_i[2]_pad  & ~n13847 ;
  assign n49314 = n13855 & n49313 ;
  assign n49315 = \m2_addr_i[2]_pad  & n13847 ;
  assign n49316 = n13840 & n49315 ;
  assign n49317 = ~n49314 & ~n49316 ;
  assign n49318 = n49312 & n49317 ;
  assign n49319 = n49307 & n49318 ;
  assign n49320 = \m0_addr_i[30]_pad  & n13847 ;
  assign n49321 = n13855 & n49320 ;
  assign n49322 = \m7_addr_i[30]_pad  & ~n13847 ;
  assign n49323 = n13864 & n49322 ;
  assign n49324 = ~n49321 & ~n49323 ;
  assign n49325 = \m3_addr_i[30]_pad  & ~n13847 ;
  assign n49326 = n13840 & n49325 ;
  assign n49327 = \m6_addr_i[30]_pad  & n13847 ;
  assign n49328 = n13864 & n49327 ;
  assign n49329 = ~n49326 & ~n49328 ;
  assign n49330 = n49324 & n49329 ;
  assign n49331 = \m4_addr_i[30]_pad  & n13847 ;
  assign n49332 = n13872 & n49331 ;
  assign n49333 = \m5_addr_i[30]_pad  & ~n13847 ;
  assign n49334 = n13872 & n49333 ;
  assign n49335 = ~n49332 & ~n49334 ;
  assign n49336 = \m1_addr_i[30]_pad  & ~n13847 ;
  assign n49337 = n13855 & n49336 ;
  assign n49338 = \m2_addr_i[30]_pad  & n13847 ;
  assign n49339 = n13840 & n49338 ;
  assign n49340 = ~n49337 & ~n49339 ;
  assign n49341 = n49335 & n49340 ;
  assign n49342 = n49330 & n49341 ;
  assign n49343 = \m1_addr_i[31]_pad  & ~n13847 ;
  assign n49344 = n13855 & n49343 ;
  assign n49345 = \m2_addr_i[31]_pad  & n13847 ;
  assign n49346 = n13840 & n49345 ;
  assign n49347 = ~n49344 & ~n49346 ;
  assign n49348 = \m0_addr_i[31]_pad  & n13847 ;
  assign n49349 = n13855 & n49348 ;
  assign n49350 = \m4_addr_i[31]_pad  & n13847 ;
  assign n49351 = n13872 & n49350 ;
  assign n49352 = ~n49349 & ~n49351 ;
  assign n49353 = n49347 & n49352 ;
  assign n49354 = \m7_addr_i[31]_pad  & ~n13847 ;
  assign n49355 = n13864 & n49354 ;
  assign n49356 = \m3_addr_i[31]_pad  & ~n13847 ;
  assign n49357 = n13840 & n49356 ;
  assign n49358 = ~n49355 & ~n49357 ;
  assign n49359 = \m5_addr_i[31]_pad  & ~n13847 ;
  assign n49360 = n13872 & n49359 ;
  assign n49361 = \m6_addr_i[31]_pad  & n13847 ;
  assign n49362 = n13864 & n49361 ;
  assign n49363 = ~n49360 & ~n49362 ;
  assign n49364 = n49358 & n49363 ;
  assign n49365 = n49353 & n49364 ;
  assign n49366 = \m3_addr_i[3]_pad  & ~n13847 ;
  assign n49367 = n13840 & n49366 ;
  assign n49368 = \m4_addr_i[3]_pad  & n13847 ;
  assign n49369 = n13872 & n49368 ;
  assign n49370 = ~n49367 & ~n49369 ;
  assign n49371 = \m6_addr_i[3]_pad  & n13847 ;
  assign n49372 = n13864 & n49371 ;
  assign n49373 = \m2_addr_i[3]_pad  & n13847 ;
  assign n49374 = n13840 & n49373 ;
  assign n49375 = ~n49372 & ~n49374 ;
  assign n49376 = n49370 & n49375 ;
  assign n49377 = \m5_addr_i[3]_pad  & ~n13847 ;
  assign n49378 = n13872 & n49377 ;
  assign n49379 = \m1_addr_i[3]_pad  & ~n13847 ;
  assign n49380 = n13855 & n49379 ;
  assign n49381 = ~n49378 & ~n49380 ;
  assign n49382 = \m0_addr_i[3]_pad  & n13847 ;
  assign n49383 = n13855 & n49382 ;
  assign n49384 = \m7_addr_i[3]_pad  & ~n13847 ;
  assign n49385 = n13864 & n49384 ;
  assign n49386 = ~n49383 & ~n49385 ;
  assign n49387 = n49381 & n49386 ;
  assign n49388 = n49376 & n49387 ;
  assign n49389 = \m3_addr_i[4]_pad  & ~n13847 ;
  assign n49390 = n13840 & n49389 ;
  assign n49391 = \m4_addr_i[4]_pad  & n13847 ;
  assign n49392 = n13872 & n49391 ;
  assign n49393 = ~n49390 & ~n49392 ;
  assign n49394 = \m6_addr_i[4]_pad  & n13847 ;
  assign n49395 = n13864 & n49394 ;
  assign n49396 = \m2_addr_i[4]_pad  & n13847 ;
  assign n49397 = n13840 & n49396 ;
  assign n49398 = ~n49395 & ~n49397 ;
  assign n49399 = n49393 & n49398 ;
  assign n49400 = \m5_addr_i[4]_pad  & ~n13847 ;
  assign n49401 = n13872 & n49400 ;
  assign n49402 = \m1_addr_i[4]_pad  & ~n13847 ;
  assign n49403 = n13855 & n49402 ;
  assign n49404 = ~n49401 & ~n49403 ;
  assign n49405 = \m0_addr_i[4]_pad  & n13847 ;
  assign n49406 = n13855 & n49405 ;
  assign n49407 = \m7_addr_i[4]_pad  & ~n13847 ;
  assign n49408 = n13864 & n49407 ;
  assign n49409 = ~n49406 & ~n49408 ;
  assign n49410 = n49404 & n49409 ;
  assign n49411 = n49399 & n49410 ;
  assign n49412 = \m1_addr_i[5]_pad  & ~n13847 ;
  assign n49413 = n13855 & n49412 ;
  assign n49414 = \m2_addr_i[5]_pad  & n13847 ;
  assign n49415 = n13840 & n49414 ;
  assign n49416 = ~n49413 & ~n49415 ;
  assign n49417 = \m3_addr_i[5]_pad  & ~n13847 ;
  assign n49418 = n13840 & n49417 ;
  assign n49419 = \m7_addr_i[5]_pad  & ~n13847 ;
  assign n49420 = n13864 & n49419 ;
  assign n49421 = ~n49418 & ~n49420 ;
  assign n49422 = n49416 & n49421 ;
  assign n49423 = \m4_addr_i[5]_pad  & n13847 ;
  assign n49424 = n13872 & n49423 ;
  assign n49425 = \m0_addr_i[5]_pad  & n13847 ;
  assign n49426 = n13855 & n49425 ;
  assign n49427 = ~n49424 & ~n49426 ;
  assign n49428 = \m6_addr_i[5]_pad  & n13847 ;
  assign n49429 = n13864 & n49428 ;
  assign n49430 = \m5_addr_i[5]_pad  & ~n13847 ;
  assign n49431 = n13872 & n49430 ;
  assign n49432 = ~n49429 & ~n49431 ;
  assign n49433 = n49427 & n49432 ;
  assign n49434 = n49422 & n49433 ;
  assign n49435 = \m1_addr_i[6]_pad  & ~n13847 ;
  assign n49436 = n13855 & n49435 ;
  assign n49437 = \m2_addr_i[6]_pad  & n13847 ;
  assign n49438 = n13840 & n49437 ;
  assign n49439 = ~n49436 & ~n49438 ;
  assign n49440 = \m0_addr_i[6]_pad  & n13847 ;
  assign n49441 = n13855 & n49440 ;
  assign n49442 = \m4_addr_i[6]_pad  & n13847 ;
  assign n49443 = n13872 & n49442 ;
  assign n49444 = ~n49441 & ~n49443 ;
  assign n49445 = n49439 & n49444 ;
  assign n49446 = \m7_addr_i[6]_pad  & ~n13847 ;
  assign n49447 = n13864 & n49446 ;
  assign n49448 = \m3_addr_i[6]_pad  & ~n13847 ;
  assign n49449 = n13840 & n49448 ;
  assign n49450 = ~n49447 & ~n49449 ;
  assign n49451 = \m6_addr_i[6]_pad  & n13847 ;
  assign n49452 = n13864 & n49451 ;
  assign n49453 = \m5_addr_i[6]_pad  & ~n13847 ;
  assign n49454 = n13872 & n49453 ;
  assign n49455 = ~n49452 & ~n49454 ;
  assign n49456 = n49450 & n49455 ;
  assign n49457 = n49445 & n49456 ;
  assign n49458 = \m6_addr_i[7]_pad  & n13847 ;
  assign n49459 = n13864 & n49458 ;
  assign n49460 = \m5_addr_i[7]_pad  & ~n13847 ;
  assign n49461 = n13872 & n49460 ;
  assign n49462 = ~n49459 & ~n49461 ;
  assign n49463 = \m1_addr_i[7]_pad  & ~n13847 ;
  assign n49464 = n13855 & n49463 ;
  assign n49465 = \m4_addr_i[7]_pad  & n13847 ;
  assign n49466 = n13872 & n49465 ;
  assign n49467 = ~n49464 & ~n49466 ;
  assign n49468 = n49462 & n49467 ;
  assign n49469 = \m2_addr_i[7]_pad  & n13847 ;
  assign n49470 = n13840 & n49469 ;
  assign n49471 = \m3_addr_i[7]_pad  & ~n13847 ;
  assign n49472 = n13840 & n49471 ;
  assign n49473 = ~n49470 & ~n49472 ;
  assign n49474 = \m0_addr_i[7]_pad  & n13847 ;
  assign n49475 = n13855 & n49474 ;
  assign n49476 = \m7_addr_i[7]_pad  & ~n13847 ;
  assign n49477 = n13864 & n49476 ;
  assign n49478 = ~n49475 & ~n49477 ;
  assign n49479 = n49473 & n49478 ;
  assign n49480 = n49468 & n49479 ;
  assign n49481 = \m1_addr_i[8]_pad  & ~n13847 ;
  assign n49482 = n13855 & n49481 ;
  assign n49483 = \m2_addr_i[8]_pad  & n13847 ;
  assign n49484 = n13840 & n49483 ;
  assign n49485 = ~n49482 & ~n49484 ;
  assign n49486 = \m3_addr_i[8]_pad  & ~n13847 ;
  assign n49487 = n13840 & n49486 ;
  assign n49488 = \m7_addr_i[8]_pad  & ~n13847 ;
  assign n49489 = n13864 & n49488 ;
  assign n49490 = ~n49487 & ~n49489 ;
  assign n49491 = n49485 & n49490 ;
  assign n49492 = \m4_addr_i[8]_pad  & n13847 ;
  assign n49493 = n13872 & n49492 ;
  assign n49494 = \m0_addr_i[8]_pad  & n13847 ;
  assign n49495 = n13855 & n49494 ;
  assign n49496 = ~n49493 & ~n49495 ;
  assign n49497 = \m6_addr_i[8]_pad  & n13847 ;
  assign n49498 = n13864 & n49497 ;
  assign n49499 = \m5_addr_i[8]_pad  & ~n13847 ;
  assign n49500 = n13872 & n49499 ;
  assign n49501 = ~n49498 & ~n49500 ;
  assign n49502 = n49496 & n49501 ;
  assign n49503 = n49491 & n49502 ;
  assign n49504 = \m0_addr_i[9]_pad  & n13847 ;
  assign n49505 = n13855 & n49504 ;
  assign n49506 = \m7_addr_i[9]_pad  & ~n13847 ;
  assign n49507 = n13864 & n49506 ;
  assign n49508 = ~n49505 & ~n49507 ;
  assign n49509 = \m1_addr_i[9]_pad  & ~n13847 ;
  assign n49510 = n13855 & n49509 ;
  assign n49511 = \m4_addr_i[9]_pad  & n13847 ;
  assign n49512 = n13872 & n49511 ;
  assign n49513 = ~n49510 & ~n49512 ;
  assign n49514 = n49508 & n49513 ;
  assign n49515 = \m2_addr_i[9]_pad  & n13847 ;
  assign n49516 = n13840 & n49515 ;
  assign n49517 = \m3_addr_i[9]_pad  & ~n13847 ;
  assign n49518 = n13840 & n49517 ;
  assign n49519 = ~n49516 & ~n49518 ;
  assign n49520 = \m6_addr_i[9]_pad  & n13847 ;
  assign n49521 = n13864 & n49520 ;
  assign n49522 = \m5_addr_i[9]_pad  & ~n13847 ;
  assign n49523 = n13872 & n49522 ;
  assign n49524 = ~n49521 & ~n49523 ;
  assign n49525 = n49519 & n49524 ;
  assign n49526 = n49514 & n49525 ;
  assign n49527 = \m0_data_i[0]_pad  & n13847 ;
  assign n49528 = n13855 & n49527 ;
  assign n49529 = \m7_data_i[0]_pad  & ~n13847 ;
  assign n49530 = n13864 & n49529 ;
  assign n49531 = ~n49528 & ~n49530 ;
  assign n49532 = \m6_data_i[0]_pad  & n13847 ;
  assign n49533 = n13864 & n49532 ;
  assign n49534 = \m2_data_i[0]_pad  & n13847 ;
  assign n49535 = n13840 & n49534 ;
  assign n49536 = ~n49533 & ~n49535 ;
  assign n49537 = n49531 & n49536 ;
  assign n49538 = \m5_data_i[0]_pad  & ~n13847 ;
  assign n49539 = n13872 & n49538 ;
  assign n49540 = \m1_data_i[0]_pad  & ~n13847 ;
  assign n49541 = n13855 & n49540 ;
  assign n49542 = ~n49539 & ~n49541 ;
  assign n49543 = \m3_data_i[0]_pad  & ~n13847 ;
  assign n49544 = n13840 & n49543 ;
  assign n49545 = \m4_data_i[0]_pad  & n13847 ;
  assign n49546 = n13872 & n49545 ;
  assign n49547 = ~n49544 & ~n49546 ;
  assign n49548 = n49542 & n49547 ;
  assign n49549 = n49537 & n49548 ;
  assign n49550 = \m6_data_i[10]_pad  & n13847 ;
  assign n49551 = n13864 & n49550 ;
  assign n49552 = \m5_data_i[10]_pad  & ~n13847 ;
  assign n49553 = n13872 & n49552 ;
  assign n49554 = ~n49551 & ~n49553 ;
  assign n49555 = \m1_data_i[10]_pad  & ~n13847 ;
  assign n49556 = n13855 & n49555 ;
  assign n49557 = \m7_data_i[10]_pad  & ~n13847 ;
  assign n49558 = n13864 & n49557 ;
  assign n49559 = ~n49556 & ~n49558 ;
  assign n49560 = n49554 & n49559 ;
  assign n49561 = \m2_data_i[10]_pad  & n13847 ;
  assign n49562 = n13840 & n49561 ;
  assign n49563 = \m0_data_i[10]_pad  & n13847 ;
  assign n49564 = n13855 & n49563 ;
  assign n49565 = ~n49562 & ~n49564 ;
  assign n49566 = \m3_data_i[10]_pad  & ~n13847 ;
  assign n49567 = n13840 & n49566 ;
  assign n49568 = \m4_data_i[10]_pad  & n13847 ;
  assign n49569 = n13872 & n49568 ;
  assign n49570 = ~n49567 & ~n49569 ;
  assign n49571 = n49565 & n49570 ;
  assign n49572 = n49560 & n49571 ;
  assign n49573 = \m1_data_i[11]_pad  & ~n13847 ;
  assign n49574 = n13855 & n49573 ;
  assign n49575 = \m2_data_i[11]_pad  & n13847 ;
  assign n49576 = n13840 & n49575 ;
  assign n49577 = ~n49574 & ~n49576 ;
  assign n49578 = \m6_data_i[11]_pad  & n13847 ;
  assign n49579 = n13864 & n49578 ;
  assign n49580 = \m4_data_i[11]_pad  & n13847 ;
  assign n49581 = n13872 & n49580 ;
  assign n49582 = ~n49579 & ~n49581 ;
  assign n49583 = n49577 & n49582 ;
  assign n49584 = \m5_data_i[11]_pad  & ~n13847 ;
  assign n49585 = n13872 & n49584 ;
  assign n49586 = \m3_data_i[11]_pad  & ~n13847 ;
  assign n49587 = n13840 & n49586 ;
  assign n49588 = ~n49585 & ~n49587 ;
  assign n49589 = \m0_data_i[11]_pad  & n13847 ;
  assign n49590 = n13855 & n49589 ;
  assign n49591 = \m7_data_i[11]_pad  & ~n13847 ;
  assign n49592 = n13864 & n49591 ;
  assign n49593 = ~n49590 & ~n49592 ;
  assign n49594 = n49588 & n49593 ;
  assign n49595 = n49583 & n49594 ;
  assign n49596 = \m1_data_i[12]_pad  & ~n13847 ;
  assign n49597 = n13855 & n49596 ;
  assign n49598 = \m2_data_i[12]_pad  & n13847 ;
  assign n49599 = n13840 & n49598 ;
  assign n49600 = ~n49597 & ~n49599 ;
  assign n49601 = \m6_data_i[12]_pad  & n13847 ;
  assign n49602 = n13864 & n49601 ;
  assign n49603 = \m7_data_i[12]_pad  & ~n13847 ;
  assign n49604 = n13864 & n49603 ;
  assign n49605 = ~n49602 & ~n49604 ;
  assign n49606 = n49600 & n49605 ;
  assign n49607 = \m5_data_i[12]_pad  & ~n13847 ;
  assign n49608 = n13872 & n49607 ;
  assign n49609 = \m0_data_i[12]_pad  & n13847 ;
  assign n49610 = n13855 & n49609 ;
  assign n49611 = ~n49608 & ~n49610 ;
  assign n49612 = \m3_data_i[12]_pad  & ~n13847 ;
  assign n49613 = n13840 & n49612 ;
  assign n49614 = \m4_data_i[12]_pad  & n13847 ;
  assign n49615 = n13872 & n49614 ;
  assign n49616 = ~n49613 & ~n49615 ;
  assign n49617 = n49611 & n49616 ;
  assign n49618 = n49606 & n49617 ;
  assign n49619 = \m1_data_i[13]_pad  & ~n13847 ;
  assign n49620 = n13855 & n49619 ;
  assign n49621 = \m2_data_i[13]_pad  & n13847 ;
  assign n49622 = n13840 & n49621 ;
  assign n49623 = ~n49620 & ~n49622 ;
  assign n49624 = \m6_data_i[13]_pad  & n13847 ;
  assign n49625 = n13864 & n49624 ;
  assign n49626 = \m7_data_i[13]_pad  & ~n13847 ;
  assign n49627 = n13864 & n49626 ;
  assign n49628 = ~n49625 & ~n49627 ;
  assign n49629 = n49623 & n49628 ;
  assign n49630 = \m5_data_i[13]_pad  & ~n13847 ;
  assign n49631 = n13872 & n49630 ;
  assign n49632 = \m0_data_i[13]_pad  & n13847 ;
  assign n49633 = n13855 & n49632 ;
  assign n49634 = ~n49631 & ~n49633 ;
  assign n49635 = \m3_data_i[13]_pad  & ~n13847 ;
  assign n49636 = n13840 & n49635 ;
  assign n49637 = \m4_data_i[13]_pad  & n13847 ;
  assign n49638 = n13872 & n49637 ;
  assign n49639 = ~n49636 & ~n49638 ;
  assign n49640 = n49634 & n49639 ;
  assign n49641 = n49629 & n49640 ;
  assign n49642 = \m3_data_i[14]_pad  & ~n13847 ;
  assign n49643 = n13840 & n49642 ;
  assign n49644 = \m4_data_i[14]_pad  & n13847 ;
  assign n49645 = n13872 & n49644 ;
  assign n49646 = ~n49643 & ~n49645 ;
  assign n49647 = \m6_data_i[14]_pad  & n13847 ;
  assign n49648 = n13864 & n49647 ;
  assign n49649 = \m7_data_i[14]_pad  & ~n13847 ;
  assign n49650 = n13864 & n49649 ;
  assign n49651 = ~n49648 & ~n49650 ;
  assign n49652 = n49646 & n49651 ;
  assign n49653 = \m5_data_i[14]_pad  & ~n13847 ;
  assign n49654 = n13872 & n49653 ;
  assign n49655 = \m0_data_i[14]_pad  & n13847 ;
  assign n49656 = n13855 & n49655 ;
  assign n49657 = ~n49654 & ~n49656 ;
  assign n49658 = \m1_data_i[14]_pad  & ~n13847 ;
  assign n49659 = n13855 & n49658 ;
  assign n49660 = \m2_data_i[14]_pad  & n13847 ;
  assign n49661 = n13840 & n49660 ;
  assign n49662 = ~n49659 & ~n49661 ;
  assign n49663 = n49657 & n49662 ;
  assign n49664 = n49652 & n49663 ;
  assign n49665 = \m6_data_i[15]_pad  & n13847 ;
  assign n49666 = n13864 & n49665 ;
  assign n49667 = \m5_data_i[15]_pad  & ~n13847 ;
  assign n49668 = n13872 & n49667 ;
  assign n49669 = ~n49666 & ~n49668 ;
  assign n49670 = \m3_data_i[15]_pad  & ~n13847 ;
  assign n49671 = n13840 & n49670 ;
  assign n49672 = \m2_data_i[15]_pad  & n13847 ;
  assign n49673 = n13840 & n49672 ;
  assign n49674 = ~n49671 & ~n49673 ;
  assign n49675 = n49669 & n49674 ;
  assign n49676 = \m4_data_i[15]_pad  & n13847 ;
  assign n49677 = n13872 & n49676 ;
  assign n49678 = \m1_data_i[15]_pad  & ~n13847 ;
  assign n49679 = n13855 & n49678 ;
  assign n49680 = ~n49677 & ~n49679 ;
  assign n49681 = \m0_data_i[15]_pad  & n13847 ;
  assign n49682 = n13855 & n49681 ;
  assign n49683 = \m7_data_i[15]_pad  & ~n13847 ;
  assign n49684 = n13864 & n49683 ;
  assign n49685 = ~n49682 & ~n49684 ;
  assign n49686 = n49680 & n49685 ;
  assign n49687 = n49675 & n49686 ;
  assign n49688 = \m1_data_i[16]_pad  & ~n13847 ;
  assign n49689 = n13855 & n49688 ;
  assign n49690 = \m2_data_i[16]_pad  & n13847 ;
  assign n49691 = n13840 & n49690 ;
  assign n49692 = ~n49689 & ~n49691 ;
  assign n49693 = \m0_data_i[16]_pad  & n13847 ;
  assign n49694 = n13855 & n49693 ;
  assign n49695 = \m4_data_i[16]_pad  & n13847 ;
  assign n49696 = n13872 & n49695 ;
  assign n49697 = ~n49694 & ~n49696 ;
  assign n49698 = n49692 & n49697 ;
  assign n49699 = \m7_data_i[16]_pad  & ~n13847 ;
  assign n49700 = n13864 & n49699 ;
  assign n49701 = \m3_data_i[16]_pad  & ~n13847 ;
  assign n49702 = n13840 & n49701 ;
  assign n49703 = ~n49700 & ~n49702 ;
  assign n49704 = \m6_data_i[16]_pad  & n13847 ;
  assign n49705 = n13864 & n49704 ;
  assign n49706 = \m5_data_i[16]_pad  & ~n13847 ;
  assign n49707 = n13872 & n49706 ;
  assign n49708 = ~n49705 & ~n49707 ;
  assign n49709 = n49703 & n49708 ;
  assign n49710 = n49698 & n49709 ;
  assign n49711 = \m3_data_i[17]_pad  & ~n13847 ;
  assign n49712 = n13840 & n49711 ;
  assign n49713 = \m4_data_i[17]_pad  & n13847 ;
  assign n49714 = n13872 & n49713 ;
  assign n49715 = ~n49712 & ~n49714 ;
  assign n49716 = \m0_data_i[17]_pad  & n13847 ;
  assign n49717 = n13855 & n49716 ;
  assign n49718 = \m5_data_i[17]_pad  & ~n13847 ;
  assign n49719 = n13872 & n49718 ;
  assign n49720 = ~n49717 & ~n49719 ;
  assign n49721 = n49715 & n49720 ;
  assign n49722 = \m7_data_i[17]_pad  & ~n13847 ;
  assign n49723 = n13864 & n49722 ;
  assign n49724 = \m6_data_i[17]_pad  & n13847 ;
  assign n49725 = n13864 & n49724 ;
  assign n49726 = ~n49723 & ~n49725 ;
  assign n49727 = \m1_data_i[17]_pad  & ~n13847 ;
  assign n49728 = n13855 & n49727 ;
  assign n49729 = \m2_data_i[17]_pad  & n13847 ;
  assign n49730 = n13840 & n49729 ;
  assign n49731 = ~n49728 & ~n49730 ;
  assign n49732 = n49726 & n49731 ;
  assign n49733 = n49721 & n49732 ;
  assign n49734 = \m3_data_i[18]_pad  & ~n13847 ;
  assign n49735 = n13840 & n49734 ;
  assign n49736 = \m4_data_i[18]_pad  & n13847 ;
  assign n49737 = n13872 & n49736 ;
  assign n49738 = ~n49735 & ~n49737 ;
  assign n49739 = \m6_data_i[18]_pad  & n13847 ;
  assign n49740 = n13864 & n49739 ;
  assign n49741 = \m2_data_i[18]_pad  & n13847 ;
  assign n49742 = n13840 & n49741 ;
  assign n49743 = ~n49740 & ~n49742 ;
  assign n49744 = n49738 & n49743 ;
  assign n49745 = \m5_data_i[18]_pad  & ~n13847 ;
  assign n49746 = n13872 & n49745 ;
  assign n49747 = \m1_data_i[18]_pad  & ~n13847 ;
  assign n49748 = n13855 & n49747 ;
  assign n49749 = ~n49746 & ~n49748 ;
  assign n49750 = \m0_data_i[18]_pad  & n13847 ;
  assign n49751 = n13855 & n49750 ;
  assign n49752 = \m7_data_i[18]_pad  & ~n13847 ;
  assign n49753 = n13864 & n49752 ;
  assign n49754 = ~n49751 & ~n49753 ;
  assign n49755 = n49749 & n49754 ;
  assign n49756 = n49744 & n49755 ;
  assign n49757 = \m0_data_i[19]_pad  & n13847 ;
  assign n49758 = n13855 & n49757 ;
  assign n49759 = \m7_data_i[19]_pad  & ~n13847 ;
  assign n49760 = n13864 & n49759 ;
  assign n49761 = ~n49758 & ~n49760 ;
  assign n49762 = \m1_data_i[19]_pad  & ~n13847 ;
  assign n49763 = n13855 & n49762 ;
  assign n49764 = \m4_data_i[19]_pad  & n13847 ;
  assign n49765 = n13872 & n49764 ;
  assign n49766 = ~n49763 & ~n49765 ;
  assign n49767 = n49761 & n49766 ;
  assign n49768 = \m2_data_i[19]_pad  & n13847 ;
  assign n49769 = n13840 & n49768 ;
  assign n49770 = \m3_data_i[19]_pad  & ~n13847 ;
  assign n49771 = n13840 & n49770 ;
  assign n49772 = ~n49769 & ~n49771 ;
  assign n49773 = \m6_data_i[19]_pad  & n13847 ;
  assign n49774 = n13864 & n49773 ;
  assign n49775 = \m5_data_i[19]_pad  & ~n13847 ;
  assign n49776 = n13872 & n49775 ;
  assign n49777 = ~n49774 & ~n49776 ;
  assign n49778 = n49772 & n49777 ;
  assign n49779 = n49767 & n49778 ;
  assign n49780 = \m3_data_i[1]_pad  & ~n13847 ;
  assign n49781 = n13840 & n49780 ;
  assign n49782 = \m4_data_i[1]_pad  & n13847 ;
  assign n49783 = n13872 & n49782 ;
  assign n49784 = ~n49781 & ~n49783 ;
  assign n49785 = \m6_data_i[1]_pad  & n13847 ;
  assign n49786 = n13864 & n49785 ;
  assign n49787 = \m2_data_i[1]_pad  & n13847 ;
  assign n49788 = n13840 & n49787 ;
  assign n49789 = ~n49786 & ~n49788 ;
  assign n49790 = n49784 & n49789 ;
  assign n49791 = \m5_data_i[1]_pad  & ~n13847 ;
  assign n49792 = n13872 & n49791 ;
  assign n49793 = \m1_data_i[1]_pad  & ~n13847 ;
  assign n49794 = n13855 & n49793 ;
  assign n49795 = ~n49792 & ~n49794 ;
  assign n49796 = \m0_data_i[1]_pad  & n13847 ;
  assign n49797 = n13855 & n49796 ;
  assign n49798 = \m7_data_i[1]_pad  & ~n13847 ;
  assign n49799 = n13864 & n49798 ;
  assign n49800 = ~n49797 & ~n49799 ;
  assign n49801 = n49795 & n49800 ;
  assign n49802 = n49790 & n49801 ;
  assign n49803 = \m3_data_i[20]_pad  & ~n13847 ;
  assign n49804 = n13840 & n49803 ;
  assign n49805 = \m4_data_i[20]_pad  & n13847 ;
  assign n49806 = n13872 & n49805 ;
  assign n49807 = ~n49804 & ~n49806 ;
  assign n49808 = \m6_data_i[20]_pad  & n13847 ;
  assign n49809 = n13864 & n49808 ;
  assign n49810 = \m2_data_i[20]_pad  & n13847 ;
  assign n49811 = n13840 & n49810 ;
  assign n49812 = ~n49809 & ~n49811 ;
  assign n49813 = n49807 & n49812 ;
  assign n49814 = \m5_data_i[20]_pad  & ~n13847 ;
  assign n49815 = n13872 & n49814 ;
  assign n49816 = \m1_data_i[20]_pad  & ~n13847 ;
  assign n49817 = n13855 & n49816 ;
  assign n49818 = ~n49815 & ~n49817 ;
  assign n49819 = \m0_data_i[20]_pad  & n13847 ;
  assign n49820 = n13855 & n49819 ;
  assign n49821 = \m7_data_i[20]_pad  & ~n13847 ;
  assign n49822 = n13864 & n49821 ;
  assign n49823 = ~n49820 & ~n49822 ;
  assign n49824 = n49818 & n49823 ;
  assign n49825 = n49813 & n49824 ;
  assign n49826 = \m1_data_i[21]_pad  & ~n13847 ;
  assign n49827 = n13855 & n49826 ;
  assign n49828 = \m2_data_i[21]_pad  & n13847 ;
  assign n49829 = n13840 & n49828 ;
  assign n49830 = ~n49827 & ~n49829 ;
  assign n49831 = \m6_data_i[21]_pad  & n13847 ;
  assign n49832 = n13864 & n49831 ;
  assign n49833 = \m7_data_i[21]_pad  & ~n13847 ;
  assign n49834 = n13864 & n49833 ;
  assign n49835 = ~n49832 & ~n49834 ;
  assign n49836 = n49830 & n49835 ;
  assign n49837 = \m5_data_i[21]_pad  & ~n13847 ;
  assign n49838 = n13872 & n49837 ;
  assign n49839 = \m0_data_i[21]_pad  & n13847 ;
  assign n49840 = n13855 & n49839 ;
  assign n49841 = ~n49838 & ~n49840 ;
  assign n49842 = \m3_data_i[21]_pad  & ~n13847 ;
  assign n49843 = n13840 & n49842 ;
  assign n49844 = \m4_data_i[21]_pad  & n13847 ;
  assign n49845 = n13872 & n49844 ;
  assign n49846 = ~n49843 & ~n49845 ;
  assign n49847 = n49841 & n49846 ;
  assign n49848 = n49836 & n49847 ;
  assign n49849 = \m3_data_i[22]_pad  & ~n13847 ;
  assign n49850 = n13840 & n49849 ;
  assign n49851 = \m4_data_i[22]_pad  & n13847 ;
  assign n49852 = n13872 & n49851 ;
  assign n49853 = ~n49850 & ~n49852 ;
  assign n49854 = \m6_data_i[22]_pad  & n13847 ;
  assign n49855 = n13864 & n49854 ;
  assign n49856 = \m2_data_i[22]_pad  & n13847 ;
  assign n49857 = n13840 & n49856 ;
  assign n49858 = ~n49855 & ~n49857 ;
  assign n49859 = n49853 & n49858 ;
  assign n49860 = \m5_data_i[22]_pad  & ~n13847 ;
  assign n49861 = n13872 & n49860 ;
  assign n49862 = \m1_data_i[22]_pad  & ~n13847 ;
  assign n49863 = n13855 & n49862 ;
  assign n49864 = ~n49861 & ~n49863 ;
  assign n49865 = \m0_data_i[22]_pad  & n13847 ;
  assign n49866 = n13855 & n49865 ;
  assign n49867 = \m7_data_i[22]_pad  & ~n13847 ;
  assign n49868 = n13864 & n49867 ;
  assign n49869 = ~n49866 & ~n49868 ;
  assign n49870 = n49864 & n49869 ;
  assign n49871 = n49859 & n49870 ;
  assign n49872 = \m3_data_i[23]_pad  & ~n13847 ;
  assign n49873 = n13840 & n49872 ;
  assign n49874 = \m4_data_i[23]_pad  & n13847 ;
  assign n49875 = n13872 & n49874 ;
  assign n49876 = ~n49873 & ~n49875 ;
  assign n49877 = \m6_data_i[23]_pad  & n13847 ;
  assign n49878 = n13864 & n49877 ;
  assign n49879 = \m2_data_i[23]_pad  & n13847 ;
  assign n49880 = n13840 & n49879 ;
  assign n49881 = ~n49878 & ~n49880 ;
  assign n49882 = n49876 & n49881 ;
  assign n49883 = \m5_data_i[23]_pad  & ~n13847 ;
  assign n49884 = n13872 & n49883 ;
  assign n49885 = \m1_data_i[23]_pad  & ~n13847 ;
  assign n49886 = n13855 & n49885 ;
  assign n49887 = ~n49884 & ~n49886 ;
  assign n49888 = \m0_data_i[23]_pad  & n13847 ;
  assign n49889 = n13855 & n49888 ;
  assign n49890 = \m7_data_i[23]_pad  & ~n13847 ;
  assign n49891 = n13864 & n49890 ;
  assign n49892 = ~n49889 & ~n49891 ;
  assign n49893 = n49887 & n49892 ;
  assign n49894 = n49882 & n49893 ;
  assign n49895 = \m3_data_i[24]_pad  & ~n13847 ;
  assign n49896 = n13840 & n49895 ;
  assign n49897 = \m4_data_i[24]_pad  & n13847 ;
  assign n49898 = n13872 & n49897 ;
  assign n49899 = ~n49896 & ~n49898 ;
  assign n49900 = \m6_data_i[24]_pad  & n13847 ;
  assign n49901 = n13864 & n49900 ;
  assign n49902 = \m2_data_i[24]_pad  & n13847 ;
  assign n49903 = n13840 & n49902 ;
  assign n49904 = ~n49901 & ~n49903 ;
  assign n49905 = n49899 & n49904 ;
  assign n49906 = \m5_data_i[24]_pad  & ~n13847 ;
  assign n49907 = n13872 & n49906 ;
  assign n49908 = \m1_data_i[24]_pad  & ~n13847 ;
  assign n49909 = n13855 & n49908 ;
  assign n49910 = ~n49907 & ~n49909 ;
  assign n49911 = \m0_data_i[24]_pad  & n13847 ;
  assign n49912 = n13855 & n49911 ;
  assign n49913 = \m7_data_i[24]_pad  & ~n13847 ;
  assign n49914 = n13864 & n49913 ;
  assign n49915 = ~n49912 & ~n49914 ;
  assign n49916 = n49910 & n49915 ;
  assign n49917 = n49905 & n49916 ;
  assign n49918 = \m3_data_i[25]_pad  & ~n13847 ;
  assign n49919 = n13840 & n49918 ;
  assign n49920 = \m4_data_i[25]_pad  & n13847 ;
  assign n49921 = n13872 & n49920 ;
  assign n49922 = ~n49919 & ~n49921 ;
  assign n49923 = \m6_data_i[25]_pad  & n13847 ;
  assign n49924 = n13864 & n49923 ;
  assign n49925 = \m7_data_i[25]_pad  & ~n13847 ;
  assign n49926 = n13864 & n49925 ;
  assign n49927 = ~n49924 & ~n49926 ;
  assign n49928 = n49922 & n49927 ;
  assign n49929 = \m5_data_i[25]_pad  & ~n13847 ;
  assign n49930 = n13872 & n49929 ;
  assign n49931 = \m0_data_i[25]_pad  & n13847 ;
  assign n49932 = n13855 & n49931 ;
  assign n49933 = ~n49930 & ~n49932 ;
  assign n49934 = \m1_data_i[25]_pad  & ~n13847 ;
  assign n49935 = n13855 & n49934 ;
  assign n49936 = \m2_data_i[25]_pad  & n13847 ;
  assign n49937 = n13840 & n49936 ;
  assign n49938 = ~n49935 & ~n49937 ;
  assign n49939 = n49933 & n49938 ;
  assign n49940 = n49928 & n49939 ;
  assign n49941 = \m1_data_i[26]_pad  & ~n13847 ;
  assign n49942 = n13855 & n49941 ;
  assign n49943 = \m2_data_i[26]_pad  & n13847 ;
  assign n49944 = n13840 & n49943 ;
  assign n49945 = ~n49942 & ~n49944 ;
  assign n49946 = \m0_data_i[26]_pad  & n13847 ;
  assign n49947 = n13855 & n49946 ;
  assign n49948 = \m4_data_i[26]_pad  & n13847 ;
  assign n49949 = n13872 & n49948 ;
  assign n49950 = ~n49947 & ~n49949 ;
  assign n49951 = n49945 & n49950 ;
  assign n49952 = \m7_data_i[26]_pad  & ~n13847 ;
  assign n49953 = n13864 & n49952 ;
  assign n49954 = \m3_data_i[26]_pad  & ~n13847 ;
  assign n49955 = n13840 & n49954 ;
  assign n49956 = ~n49953 & ~n49955 ;
  assign n49957 = \m6_data_i[26]_pad  & n13847 ;
  assign n49958 = n13864 & n49957 ;
  assign n49959 = \m5_data_i[26]_pad  & ~n13847 ;
  assign n49960 = n13872 & n49959 ;
  assign n49961 = ~n49958 & ~n49960 ;
  assign n49962 = n49956 & n49961 ;
  assign n49963 = n49951 & n49962 ;
  assign n49964 = \m3_data_i[27]_pad  & ~n13847 ;
  assign n49965 = n13840 & n49964 ;
  assign n49966 = \m4_data_i[27]_pad  & n13847 ;
  assign n49967 = n13872 & n49966 ;
  assign n49968 = ~n49965 & ~n49967 ;
  assign n49969 = \m0_data_i[27]_pad  & n13847 ;
  assign n49970 = n13855 & n49969 ;
  assign n49971 = \m2_data_i[27]_pad  & n13847 ;
  assign n49972 = n13840 & n49971 ;
  assign n49973 = ~n49970 & ~n49972 ;
  assign n49974 = n49968 & n49973 ;
  assign n49975 = \m7_data_i[27]_pad  & ~n13847 ;
  assign n49976 = n13864 & n49975 ;
  assign n49977 = \m1_data_i[27]_pad  & ~n13847 ;
  assign n49978 = n13855 & n49977 ;
  assign n49979 = ~n49976 & ~n49978 ;
  assign n49980 = \m6_data_i[27]_pad  & n13847 ;
  assign n49981 = n13864 & n49980 ;
  assign n49982 = \m5_data_i[27]_pad  & ~n13847 ;
  assign n49983 = n13872 & n49982 ;
  assign n49984 = ~n49981 & ~n49983 ;
  assign n49985 = n49979 & n49984 ;
  assign n49986 = n49974 & n49985 ;
  assign n49987 = \m3_data_i[28]_pad  & ~n13847 ;
  assign n49988 = n13840 & n49987 ;
  assign n49989 = \m4_data_i[28]_pad  & n13847 ;
  assign n49990 = n13872 & n49989 ;
  assign n49991 = ~n49988 & ~n49990 ;
  assign n49992 = \m0_data_i[28]_pad  & n13847 ;
  assign n49993 = n13855 & n49992 ;
  assign n49994 = \m5_data_i[28]_pad  & ~n13847 ;
  assign n49995 = n13872 & n49994 ;
  assign n49996 = ~n49993 & ~n49995 ;
  assign n49997 = n49991 & n49996 ;
  assign n49998 = \m7_data_i[28]_pad  & ~n13847 ;
  assign n49999 = n13864 & n49998 ;
  assign n50000 = \m6_data_i[28]_pad  & n13847 ;
  assign n50001 = n13864 & n50000 ;
  assign n50002 = ~n49999 & ~n50001 ;
  assign n50003 = \m1_data_i[28]_pad  & ~n13847 ;
  assign n50004 = n13855 & n50003 ;
  assign n50005 = \m2_data_i[28]_pad  & n13847 ;
  assign n50006 = n13840 & n50005 ;
  assign n50007 = ~n50004 & ~n50006 ;
  assign n50008 = n50002 & n50007 ;
  assign n50009 = n49997 & n50008 ;
  assign n50010 = \m1_data_i[29]_pad  & ~n13847 ;
  assign n50011 = n13855 & n50010 ;
  assign n50012 = \m2_data_i[29]_pad  & n13847 ;
  assign n50013 = n13840 & n50012 ;
  assign n50014 = ~n50011 & ~n50013 ;
  assign n50015 = \m3_data_i[29]_pad  & ~n13847 ;
  assign n50016 = n13840 & n50015 ;
  assign n50017 = \m5_data_i[29]_pad  & ~n13847 ;
  assign n50018 = n13872 & n50017 ;
  assign n50019 = ~n50016 & ~n50018 ;
  assign n50020 = n50014 & n50019 ;
  assign n50021 = \m4_data_i[29]_pad  & n13847 ;
  assign n50022 = n13872 & n50021 ;
  assign n50023 = \m6_data_i[29]_pad  & n13847 ;
  assign n50024 = n13864 & n50023 ;
  assign n50025 = ~n50022 & ~n50024 ;
  assign n50026 = \m0_data_i[29]_pad  & n13847 ;
  assign n50027 = n13855 & n50026 ;
  assign n50028 = \m7_data_i[29]_pad  & ~n13847 ;
  assign n50029 = n13864 & n50028 ;
  assign n50030 = ~n50027 & ~n50029 ;
  assign n50031 = n50025 & n50030 ;
  assign n50032 = n50020 & n50031 ;
  assign n50033 = \m1_data_i[2]_pad  & ~n13847 ;
  assign n50034 = n13855 & n50033 ;
  assign n50035 = \m2_data_i[2]_pad  & n13847 ;
  assign n50036 = n13840 & n50035 ;
  assign n50037 = ~n50034 & ~n50036 ;
  assign n50038 = \m6_data_i[2]_pad  & n13847 ;
  assign n50039 = n13864 & n50038 ;
  assign n50040 = \m7_data_i[2]_pad  & ~n13847 ;
  assign n50041 = n13864 & n50040 ;
  assign n50042 = ~n50039 & ~n50041 ;
  assign n50043 = n50037 & n50042 ;
  assign n50044 = \m5_data_i[2]_pad  & ~n13847 ;
  assign n50045 = n13872 & n50044 ;
  assign n50046 = \m0_data_i[2]_pad  & n13847 ;
  assign n50047 = n13855 & n50046 ;
  assign n50048 = ~n50045 & ~n50047 ;
  assign n50049 = \m3_data_i[2]_pad  & ~n13847 ;
  assign n50050 = n13840 & n50049 ;
  assign n50051 = \m4_data_i[2]_pad  & n13847 ;
  assign n50052 = n13872 & n50051 ;
  assign n50053 = ~n50050 & ~n50052 ;
  assign n50054 = n50048 & n50053 ;
  assign n50055 = n50043 & n50054 ;
  assign n50056 = \m0_data_i[30]_pad  & n13847 ;
  assign n50057 = n13855 & n50056 ;
  assign n50058 = \m7_data_i[30]_pad  & ~n13847 ;
  assign n50059 = n13864 & n50058 ;
  assign n50060 = ~n50057 & ~n50059 ;
  assign n50061 = \m3_data_i[30]_pad  & ~n13847 ;
  assign n50062 = n13840 & n50061 ;
  assign n50063 = \m2_data_i[30]_pad  & n13847 ;
  assign n50064 = n13840 & n50063 ;
  assign n50065 = ~n50062 & ~n50064 ;
  assign n50066 = n50060 & n50065 ;
  assign n50067 = \m4_data_i[30]_pad  & n13847 ;
  assign n50068 = n13872 & n50067 ;
  assign n50069 = \m1_data_i[30]_pad  & ~n13847 ;
  assign n50070 = n13855 & n50069 ;
  assign n50071 = ~n50068 & ~n50070 ;
  assign n50072 = \m6_data_i[30]_pad  & n13847 ;
  assign n50073 = n13864 & n50072 ;
  assign n50074 = \m5_data_i[30]_pad  & ~n13847 ;
  assign n50075 = n13872 & n50074 ;
  assign n50076 = ~n50073 & ~n50075 ;
  assign n50077 = n50071 & n50076 ;
  assign n50078 = n50066 & n50077 ;
  assign n50079 = \m0_data_i[31]_pad  & n13847 ;
  assign n50080 = n13855 & n50079 ;
  assign n50081 = \m7_data_i[31]_pad  & ~n13847 ;
  assign n50082 = n13864 & n50081 ;
  assign n50083 = ~n50080 & ~n50082 ;
  assign n50084 = \m1_data_i[31]_pad  & ~n13847 ;
  assign n50085 = n13855 & n50084 ;
  assign n50086 = \m5_data_i[31]_pad  & ~n13847 ;
  assign n50087 = n13872 & n50086 ;
  assign n50088 = ~n50085 & ~n50087 ;
  assign n50089 = n50083 & n50088 ;
  assign n50090 = \m2_data_i[31]_pad  & n13847 ;
  assign n50091 = n13840 & n50090 ;
  assign n50092 = \m6_data_i[31]_pad  & n13847 ;
  assign n50093 = n13864 & n50092 ;
  assign n50094 = ~n50091 & ~n50093 ;
  assign n50095 = \m3_data_i[31]_pad  & ~n13847 ;
  assign n50096 = n13840 & n50095 ;
  assign n50097 = \m4_data_i[31]_pad  & n13847 ;
  assign n50098 = n13872 & n50097 ;
  assign n50099 = ~n50096 & ~n50098 ;
  assign n50100 = n50094 & n50099 ;
  assign n50101 = n50089 & n50100 ;
  assign n50102 = \m0_data_i[3]_pad  & n13847 ;
  assign n50103 = n13855 & n50102 ;
  assign n50104 = \m7_data_i[3]_pad  & ~n13847 ;
  assign n50105 = n13864 & n50104 ;
  assign n50106 = ~n50103 & ~n50105 ;
  assign n50107 = \m3_data_i[3]_pad  & ~n13847 ;
  assign n50108 = n13840 & n50107 ;
  assign n50109 = \m5_data_i[3]_pad  & ~n13847 ;
  assign n50110 = n13872 & n50109 ;
  assign n50111 = ~n50108 & ~n50110 ;
  assign n50112 = n50106 & n50111 ;
  assign n50113 = \m4_data_i[3]_pad  & n13847 ;
  assign n50114 = n13872 & n50113 ;
  assign n50115 = \m6_data_i[3]_pad  & n13847 ;
  assign n50116 = n13864 & n50115 ;
  assign n50117 = ~n50114 & ~n50116 ;
  assign n50118 = \m1_data_i[3]_pad  & ~n13847 ;
  assign n50119 = n13855 & n50118 ;
  assign n50120 = \m2_data_i[3]_pad  & n13847 ;
  assign n50121 = n13840 & n50120 ;
  assign n50122 = ~n50119 & ~n50121 ;
  assign n50123 = n50117 & n50122 ;
  assign n50124 = n50112 & n50123 ;
  assign n50125 = \m1_data_i[4]_pad  & ~n13847 ;
  assign n50126 = n13855 & n50125 ;
  assign n50127 = \m2_data_i[4]_pad  & n13847 ;
  assign n50128 = n13840 & n50127 ;
  assign n50129 = ~n50126 & ~n50128 ;
  assign n50130 = \m6_data_i[4]_pad  & n13847 ;
  assign n50131 = n13864 & n50130 ;
  assign n50132 = \m4_data_i[4]_pad  & n13847 ;
  assign n50133 = n13872 & n50132 ;
  assign n50134 = ~n50131 & ~n50133 ;
  assign n50135 = n50129 & n50134 ;
  assign n50136 = \m5_data_i[4]_pad  & ~n13847 ;
  assign n50137 = n13872 & n50136 ;
  assign n50138 = \m3_data_i[4]_pad  & ~n13847 ;
  assign n50139 = n13840 & n50138 ;
  assign n50140 = ~n50137 & ~n50139 ;
  assign n50141 = \m0_data_i[4]_pad  & n13847 ;
  assign n50142 = n13855 & n50141 ;
  assign n50143 = \m7_data_i[4]_pad  & ~n13847 ;
  assign n50144 = n13864 & n50143 ;
  assign n50145 = ~n50142 & ~n50144 ;
  assign n50146 = n50140 & n50145 ;
  assign n50147 = n50135 & n50146 ;
  assign n50148 = \m1_data_i[5]_pad  & ~n13847 ;
  assign n50149 = n13855 & n50148 ;
  assign n50150 = \m2_data_i[5]_pad  & n13847 ;
  assign n50151 = n13840 & n50150 ;
  assign n50152 = ~n50149 & ~n50151 ;
  assign n50153 = \m0_data_i[5]_pad  & n13847 ;
  assign n50154 = n13855 & n50153 ;
  assign n50155 = \m5_data_i[5]_pad  & ~n13847 ;
  assign n50156 = n13872 & n50155 ;
  assign n50157 = ~n50154 & ~n50156 ;
  assign n50158 = n50152 & n50157 ;
  assign n50159 = \m7_data_i[5]_pad  & ~n13847 ;
  assign n50160 = n13864 & n50159 ;
  assign n50161 = \m6_data_i[5]_pad  & n13847 ;
  assign n50162 = n13864 & n50161 ;
  assign n50163 = ~n50160 & ~n50162 ;
  assign n50164 = \m3_data_i[5]_pad  & ~n13847 ;
  assign n50165 = n13840 & n50164 ;
  assign n50166 = \m4_data_i[5]_pad  & n13847 ;
  assign n50167 = n13872 & n50166 ;
  assign n50168 = ~n50165 & ~n50167 ;
  assign n50169 = n50163 & n50168 ;
  assign n50170 = n50158 & n50169 ;
  assign n50171 = \m6_data_i[6]_pad  & n13847 ;
  assign n50172 = n13864 & n50171 ;
  assign n50173 = \m5_data_i[6]_pad  & ~n13847 ;
  assign n50174 = n13872 & n50173 ;
  assign n50175 = ~n50172 & ~n50174 ;
  assign n50176 = \m0_data_i[6]_pad  & n13847 ;
  assign n50177 = n13855 & n50176 ;
  assign n50178 = \m2_data_i[6]_pad  & n13847 ;
  assign n50179 = n13840 & n50178 ;
  assign n50180 = ~n50177 & ~n50179 ;
  assign n50181 = n50175 & n50180 ;
  assign n50182 = \m7_data_i[6]_pad  & ~n13847 ;
  assign n50183 = n13864 & n50182 ;
  assign n50184 = \m1_data_i[6]_pad  & ~n13847 ;
  assign n50185 = n13855 & n50184 ;
  assign n50186 = ~n50183 & ~n50185 ;
  assign n50187 = \m3_data_i[6]_pad  & ~n13847 ;
  assign n50188 = n13840 & n50187 ;
  assign n50189 = \m4_data_i[6]_pad  & n13847 ;
  assign n50190 = n13872 & n50189 ;
  assign n50191 = ~n50188 & ~n50190 ;
  assign n50192 = n50186 & n50191 ;
  assign n50193 = n50181 & n50192 ;
  assign n50194 = \m6_data_i[7]_pad  & n13847 ;
  assign n50195 = n13864 & n50194 ;
  assign n50196 = \m5_data_i[7]_pad  & ~n13847 ;
  assign n50197 = n13872 & n50196 ;
  assign n50198 = ~n50195 & ~n50197 ;
  assign n50199 = \m1_data_i[7]_pad  & ~n13847 ;
  assign n50200 = n13855 & n50199 ;
  assign n50201 = \m7_data_i[7]_pad  & ~n13847 ;
  assign n50202 = n13864 & n50201 ;
  assign n50203 = ~n50200 & ~n50202 ;
  assign n50204 = n50198 & n50203 ;
  assign n50205 = \m2_data_i[7]_pad  & n13847 ;
  assign n50206 = n13840 & n50205 ;
  assign n50207 = \m0_data_i[7]_pad  & n13847 ;
  assign n50208 = n13855 & n50207 ;
  assign n50209 = ~n50206 & ~n50208 ;
  assign n50210 = \m3_data_i[7]_pad  & ~n13847 ;
  assign n50211 = n13840 & n50210 ;
  assign n50212 = \m4_data_i[7]_pad  & n13847 ;
  assign n50213 = n13872 & n50212 ;
  assign n50214 = ~n50211 & ~n50213 ;
  assign n50215 = n50209 & n50214 ;
  assign n50216 = n50204 & n50215 ;
  assign n50217 = \m3_data_i[8]_pad  & ~n13847 ;
  assign n50218 = n13840 & n50217 ;
  assign n50219 = \m4_data_i[8]_pad  & n13847 ;
  assign n50220 = n13872 & n50219 ;
  assign n50221 = ~n50218 & ~n50220 ;
  assign n50222 = \m6_data_i[8]_pad  & n13847 ;
  assign n50223 = n13864 & n50222 ;
  assign n50224 = \m7_data_i[8]_pad  & ~n13847 ;
  assign n50225 = n13864 & n50224 ;
  assign n50226 = ~n50223 & ~n50225 ;
  assign n50227 = n50221 & n50226 ;
  assign n50228 = \m5_data_i[8]_pad  & ~n13847 ;
  assign n50229 = n13872 & n50228 ;
  assign n50230 = \m0_data_i[8]_pad  & n13847 ;
  assign n50231 = n13855 & n50230 ;
  assign n50232 = ~n50229 & ~n50231 ;
  assign n50233 = \m1_data_i[8]_pad  & ~n13847 ;
  assign n50234 = n13855 & n50233 ;
  assign n50235 = \m2_data_i[8]_pad  & n13847 ;
  assign n50236 = n13840 & n50235 ;
  assign n50237 = ~n50234 & ~n50236 ;
  assign n50238 = n50232 & n50237 ;
  assign n50239 = n50227 & n50238 ;
  assign n50240 = \m3_data_i[9]_pad  & ~n13847 ;
  assign n50241 = n13840 & n50240 ;
  assign n50242 = \m4_data_i[9]_pad  & n13847 ;
  assign n50243 = n13872 & n50242 ;
  assign n50244 = ~n50241 & ~n50243 ;
  assign n50245 = \m6_data_i[9]_pad  & n13847 ;
  assign n50246 = n13864 & n50245 ;
  assign n50247 = \m2_data_i[9]_pad  & n13847 ;
  assign n50248 = n13840 & n50247 ;
  assign n50249 = ~n50246 & ~n50248 ;
  assign n50250 = n50244 & n50249 ;
  assign n50251 = \m5_data_i[9]_pad  & ~n13847 ;
  assign n50252 = n13872 & n50251 ;
  assign n50253 = \m1_data_i[9]_pad  & ~n13847 ;
  assign n50254 = n13855 & n50253 ;
  assign n50255 = ~n50252 & ~n50254 ;
  assign n50256 = \m0_data_i[9]_pad  & n13847 ;
  assign n50257 = n13855 & n50256 ;
  assign n50258 = \m7_data_i[9]_pad  & ~n13847 ;
  assign n50259 = n13864 & n50258 ;
  assign n50260 = ~n50257 & ~n50259 ;
  assign n50261 = n50255 & n50260 ;
  assign n50262 = n50250 & n50261 ;
  assign n50263 = \m1_sel_i[0]_pad  & ~n13847 ;
  assign n50264 = n13855 & n50263 ;
  assign n50265 = \m2_sel_i[0]_pad  & n13847 ;
  assign n50266 = n13840 & n50265 ;
  assign n50267 = ~n50264 & ~n50266 ;
  assign n50268 = \m6_sel_i[0]_pad  & n13847 ;
  assign n50269 = n13864 & n50268 ;
  assign n50270 = \m4_sel_i[0]_pad  & n13847 ;
  assign n50271 = n13872 & n50270 ;
  assign n50272 = ~n50269 & ~n50271 ;
  assign n50273 = n50267 & n50272 ;
  assign n50274 = \m5_sel_i[0]_pad  & ~n13847 ;
  assign n50275 = n13872 & n50274 ;
  assign n50276 = \m3_sel_i[0]_pad  & ~n13847 ;
  assign n50277 = n13840 & n50276 ;
  assign n50278 = ~n50275 & ~n50277 ;
  assign n50279 = \m0_sel_i[0]_pad  & n13847 ;
  assign n50280 = n13855 & n50279 ;
  assign n50281 = \m7_sel_i[0]_pad  & ~n13847 ;
  assign n50282 = n13864 & n50281 ;
  assign n50283 = ~n50280 & ~n50282 ;
  assign n50284 = n50278 & n50283 ;
  assign n50285 = n50273 & n50284 ;
  assign n50286 = \m1_sel_i[1]_pad  & ~n13847 ;
  assign n50287 = n13855 & n50286 ;
  assign n50288 = \m2_sel_i[1]_pad  & n13847 ;
  assign n50289 = n13840 & n50288 ;
  assign n50290 = ~n50287 & ~n50289 ;
  assign n50291 = \m6_sel_i[1]_pad  & n13847 ;
  assign n50292 = n13864 & n50291 ;
  assign n50293 = \m7_sel_i[1]_pad  & ~n13847 ;
  assign n50294 = n13864 & n50293 ;
  assign n50295 = ~n50292 & ~n50294 ;
  assign n50296 = n50290 & n50295 ;
  assign n50297 = \m5_sel_i[1]_pad  & ~n13847 ;
  assign n50298 = n13872 & n50297 ;
  assign n50299 = \m0_sel_i[1]_pad  & n13847 ;
  assign n50300 = n13855 & n50299 ;
  assign n50301 = ~n50298 & ~n50300 ;
  assign n50302 = \m3_sel_i[1]_pad  & ~n13847 ;
  assign n50303 = n13840 & n50302 ;
  assign n50304 = \m4_sel_i[1]_pad  & n13847 ;
  assign n50305 = n13872 & n50304 ;
  assign n50306 = ~n50303 & ~n50305 ;
  assign n50307 = n50301 & n50306 ;
  assign n50308 = n50296 & n50307 ;
  assign n50309 = \m0_sel_i[2]_pad  & n13847 ;
  assign n50310 = n13855 & n50309 ;
  assign n50311 = \m7_sel_i[2]_pad  & ~n13847 ;
  assign n50312 = n13864 & n50311 ;
  assign n50313 = ~n50310 & ~n50312 ;
  assign n50314 = \m6_sel_i[2]_pad  & n13847 ;
  assign n50315 = n13864 & n50314 ;
  assign n50316 = \m4_sel_i[2]_pad  & n13847 ;
  assign n50317 = n13872 & n50316 ;
  assign n50318 = ~n50315 & ~n50317 ;
  assign n50319 = n50313 & n50318 ;
  assign n50320 = \m5_sel_i[2]_pad  & ~n13847 ;
  assign n50321 = n13872 & n50320 ;
  assign n50322 = \m3_sel_i[2]_pad  & ~n13847 ;
  assign n50323 = n13840 & n50322 ;
  assign n50324 = ~n50321 & ~n50323 ;
  assign n50325 = \m1_sel_i[2]_pad  & ~n13847 ;
  assign n50326 = n13855 & n50325 ;
  assign n50327 = \m2_sel_i[2]_pad  & n13847 ;
  assign n50328 = n13840 & n50327 ;
  assign n50329 = ~n50326 & ~n50328 ;
  assign n50330 = n50324 & n50329 ;
  assign n50331 = n50319 & n50330 ;
  assign n50332 = \m1_sel_i[3]_pad  & ~n13847 ;
  assign n50333 = n13855 & n50332 ;
  assign n50334 = \m2_sel_i[3]_pad  & n13847 ;
  assign n50335 = n13840 & n50334 ;
  assign n50336 = ~n50333 & ~n50335 ;
  assign n50337 = \m0_sel_i[3]_pad  & n13847 ;
  assign n50338 = n13855 & n50337 ;
  assign n50339 = \m4_sel_i[3]_pad  & n13847 ;
  assign n50340 = n13872 & n50339 ;
  assign n50341 = ~n50338 & ~n50340 ;
  assign n50342 = n50336 & n50341 ;
  assign n50343 = \m7_sel_i[3]_pad  & ~n13847 ;
  assign n50344 = n13864 & n50343 ;
  assign n50345 = \m3_sel_i[3]_pad  & ~n13847 ;
  assign n50346 = n13840 & n50345 ;
  assign n50347 = ~n50344 & ~n50346 ;
  assign n50348 = \m6_sel_i[3]_pad  & n13847 ;
  assign n50349 = n13864 & n50348 ;
  assign n50350 = \m5_sel_i[3]_pad  & ~n13847 ;
  assign n50351 = n13872 & n50350 ;
  assign n50352 = ~n50349 & ~n50351 ;
  assign n50353 = n50347 & n50352 ;
  assign n50354 = n50342 & n50353 ;
  assign n50355 = \m3_stb_i_pad  & n14927 ;
  assign n50356 = ~n13847 & n50355 ;
  assign n50357 = n13840 & n50356 ;
  assign n50358 = \m2_stb_i_pad  & n14887 ;
  assign n50359 = n13847 & n50358 ;
  assign n50360 = n13840 & n50359 ;
  assign n50361 = ~n50357 & ~n50360 ;
  assign n50362 = \m6_stb_i_pad  & n15042 ;
  assign n50363 = n13847 & n50362 ;
  assign n50364 = n13864 & n50363 ;
  assign n50365 = \m1_stb_i_pad  & n14845 ;
  assign n50366 = ~n13847 & n50365 ;
  assign n50367 = n13855 & n50366 ;
  assign n50368 = ~n50364 & ~n50367 ;
  assign n50369 = n50361 & n50368 ;
  assign n50370 = \m7_stb_i_pad  & n14666 ;
  assign n50371 = ~n13847 & n50370 ;
  assign n50372 = n13864 & n50371 ;
  assign n50373 = \m5_stb_i_pad  & n14995 ;
  assign n50374 = ~n13847 & n50373 ;
  assign n50375 = n13872 & n50374 ;
  assign n50376 = ~n50372 & ~n50375 ;
  assign n50377 = \m4_stb_i_pad  & n14713 ;
  assign n50378 = n13847 & n50377 ;
  assign n50379 = n13872 & n50378 ;
  assign n50380 = \m0_stb_i_pad  & n15110 ;
  assign n50381 = n13847 & n50380 ;
  assign n50382 = n13855 & n50381 ;
  assign n50383 = ~n50379 & ~n50382 ;
  assign n50384 = n50376 & n50383 ;
  assign n50385 = n50369 & n50384 ;
  assign n50386 = \m3_we_i_pad  & ~n13847 ;
  assign n50387 = n13840 & n50386 ;
  assign n50388 = \m4_we_i_pad  & n13847 ;
  assign n50389 = n13872 & n50388 ;
  assign n50390 = ~n50387 & ~n50389 ;
  assign n50391 = \m6_we_i_pad  & n13847 ;
  assign n50392 = n13864 & n50391 ;
  assign n50393 = \m2_we_i_pad  & n13847 ;
  assign n50394 = n13840 & n50393 ;
  assign n50395 = ~n50392 & ~n50394 ;
  assign n50396 = n50390 & n50395 ;
  assign n50397 = \m5_we_i_pad  & ~n13847 ;
  assign n50398 = n13872 & n50397 ;
  assign n50399 = \m1_we_i_pad  & ~n13847 ;
  assign n50400 = n13855 & n50399 ;
  assign n50401 = ~n50398 & ~n50400 ;
  assign n50402 = \m0_we_i_pad  & n13847 ;
  assign n50403 = n13855 & n50402 ;
  assign n50404 = \m7_we_i_pad  & ~n13847 ;
  assign n50405 = n13864 & n50404 ;
  assign n50406 = ~n50403 & ~n50405 ;
  assign n50407 = n50401 & n50406 ;
  assign n50408 = n50396 & n50407 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g106655/_1_  = n2259 ;
  assign \g106703/_1_  = ~n1998 ;
  assign \g69412/_0_  = n2291 ;
  assign \g69413/_0_  = n2323 ;
  assign \g69417/_1_  = n2355 ;
  assign \g69418/_0_  = n2387 ;
  assign \g69420/_1_  = n2419 ;
  assign \g69421/_0_  = n2451 ;
  assign \g69423/_1_  = n2483 ;
  assign \g69424/_0_  = n2515 ;
  assign \g69426/_1_  = n2547 ;
  assign \g69428/_1_  = n2579 ;
  assign \g69430/_1_  = n2611 ;
  assign \g69432/_1_  = n2643 ;
  assign \g69434/_1_  = n2675 ;
  assign \g69436/_1_  = n2707 ;
  assign \g69438/_1_  = n2739 ;
  assign \g69757/_2_  = ~n2801 ;
  assign \g69758/_2_  = ~n2863 ;
  assign \g69759/_2_  = ~n2925 ;
  assign \g69760/_2_  = ~n2987 ;
  assign \g69761/_0_  = ~n3058 ;
  assign \g69762/_2_  = ~n3120 ;
  assign \g69763/_2_  = ~n3182 ;
  assign \g69764/_2_  = ~n3244 ;
  assign \g69765/_2_  = ~n3306 ;
  assign \g69766/_2_  = ~n3368 ;
  assign \g69767/_0_  = ~n3431 ;
  assign \g69768/_0_  = ~n3494 ;
  assign \g69769/_0_  = ~n3557 ;
  assign \g69770/_0_  = ~n3620 ;
  assign \g69771/_0_  = ~n3683 ;
  assign \g69772/_0_  = ~n3746 ;
  assign \g70206/_0_  = n3806 ;
  assign \g70392/_0_  = ~n3827 ;
  assign \g70393/_0_  = n3847 ;
  assign \g70394/_0_  = n3901 ;
  assign \g70395/_0_  = n3947 ;
  assign \g70396/_0_  = n4001 ;
  assign \g70397/_0_  = ~n4036 ;
  assign \g70398/_0_  = ~n4087 ;
  assign \g70399/_0_  = ~n4122 ;
  assign \g70400/_0_  = ~n4157 ;
  assign \g70401/_0_  = ~n4192 ;
  assign \g70402/_0_  = n4246 ;
  assign \g70403/_0_  = ~n4281 ;
  assign \g70404/_0_  = ~n4332 ;
  assign \g70405/_0_  = n4386 ;
  assign \g70406/_0_  = ~n4437 ;
  assign \g70407/_0_  = ~n4472 ;
  assign \g70408/_0_  = ~n4523 ;
  assign \g70409/_0_  = ~n4574 ;
  assign \g70410/_0_  = ~n4609 ;
  assign \g70411/_0_  = n4663 ;
  assign \g70412/_0_  = n4717 ;
  assign \g70413/_0_  = n4771 ;
  assign \g70414/_0_  = ~n4822 ;
  assign \g70415/_0_  = n4876 ;
  assign \g70416/_0_  = ~n4910 ;
  assign \g70417/_0_  = ~n4962 ;
  assign \g70418/_0_  = n4998 ;
  assign \g70419/_0_  = ~n5032 ;
  assign \g70420/_0_  = ~n5071 ;
  assign \g70421/_0_  = ~n5110 ;
  assign \g70422/_0_  = ~n5144 ;
  assign \g70423/_0_  = ~n5186 ;
  assign \g70424/_0_  = ~n5225 ;
  assign \g70425/_0_  = ~n5268 ;
  assign \g70426/_0_  = ~n5311 ;
  assign \g70427/_0_  = n5349 ;
  assign \g70428/_0_  = ~n5392 ;
  assign \g70429/_0_  = ~n5443 ;
  assign \g70430/_0_  = ~n5486 ;
  assign \g70431/_0_  = ~n5559 ;
  assign \g70432/_0_  = n5641 ;
  assign \g70433/_0_  = ~n5705 ;
  assign \g70434/_0_  = ~n5783 ;
  assign \g70435/_0_  = ~n5834 ;
  assign \g70436/_0_  = ~n5897 ;
  assign \g70437/_0_  = ~n5968 ;
  assign \g70438/_0_  = ~n6046 ;
  assign \g70439/_0_  = n6094 ;
  assign \g70440/_0_  = n6176 ;
  assign \g70441/_0_  = ~n6240 ;
  assign \g70442/_0_  = ~n6318 ;
  assign \g70443/_0_  = ~n6391 ;
  assign \g70444/_0_  = ~n6470 ;
  assign \g70445/_0_  = ~n6534 ;
  assign \g70446/_0_  = ~n6612 ;
  assign \g70447/_0_  = ~n6678 ;
  assign \g70448/_0_  = ~n6742 ;
  assign \g70449/_0_  = ~n6813 ;
  assign \g70450/_0_  = ~n6866 ;
  assign \g70451/_0_  = ~n6940 ;
  assign \g70452/_0_  = ~n6960 ;
  assign \g70453/_0_  = ~n7025 ;
  assign \g70454/_0_  = ~n7094 ;
  assign \g70455/_0_  = ~n7160 ;
  assign \g70456/_0_  = ~n7223 ;
  assign \g70457/_0_  = ~n7294 ;
  assign \g70458/_0_  = ~n7363 ;
  assign \g70459/_0_  = ~n7436 ;
  assign \g70460/_0_  = ~n7515 ;
  assign \g70461/_0_  = ~n7579 ;
  assign \g70462/_0_  = ~n7657 ;
  assign \g70463/_0_  = ~n7727 ;
  assign \g70464/_0_  = ~n7790 ;
  assign \g70465/_0_  = ~n7861 ;
  assign \g70466/_0_  = ~n7939 ;
  assign \g70467/_0_  = ~n8005 ;
  assign \g70468/_0_  = ~n8084 ;
  assign \g70469/_0_  = ~n8155 ;
  assign \g70470/_0_  = ~n8233 ;
  assign \g70471/_0_  = ~n8283 ;
  assign \g70472/_0_  = ~n8346 ;
  assign \g70473/_0_  = ~n8410 ;
  assign \g70474/_0_  = ~n8488 ;
  assign \g70475/_0_  = ~n8537 ;
  assign \g70476/_0_  = ~n8600 ;
  assign \g70477/_0_  = ~n8664 ;
  assign \g70478/_0_  = ~n8733 ;
  assign \g70479/_0_  = n8804 ;
  assign \g70480/_0_  = n8886 ;
  assign \g70481/_0_  = ~n8950 ;
  assign \g70482/_0_  = ~n9028 ;
  assign \g70483/_0_  = ~n9077 ;
  assign \g70484/_0_  = ~n9140 ;
  assign \g70485/_0_  = ~n9211 ;
  assign \g70486/_0_  = ~n9280 ;
  assign \g70487/_0_  = ~n9329 ;
  assign \g70488/_0_  = n9411 ;
  assign \g70489/_0_  = ~n9490 ;
  assign \g70490/_0_  = ~n9559 ;
  assign \g70491/_0_  = ~n9608 ;
  assign \g70492/_0_  = ~n9671 ;
  assign \g70493/_0_  = ~n9735 ;
  assign \g70494/_0_  = ~n9804 ;
  assign \g70495/_0_  = ~n9839 ;
  assign \g70496/_0_  = ~n9874 ;
  assign \g70497/_0_  = ~n9901 ;
  assign \g70498/_0_  = ~n9928 ;
  assign \g70499/_0_  = ~n9955 ;
  assign \g70500/_0_  = ~n9990 ;
  assign \g70501/_0_  = ~n10025 ;
  assign \g70502/_0_  = ~n10052 ;
  assign \g70503/_0_  = ~n10070 ;
  assign \g70504/_0_  = ~n10106 ;
  assign \g70505/_0_  = ~n10141 ;
  assign \g70506/_0_  = ~n10176 ;
  assign \g70507/_0_  = ~n10211 ;
  assign \g70508/_0_  = ~n10293 ;
  assign \g70509/_0_  = ~n10325 ;
  assign \g70510/_0_  = ~n10348 ;
  assign \g70511/_0_  = ~n10372 ;
  assign \g70513/_0_  = ~n10390 ;
  assign \g70515/_0_  = ~n10408 ;
  assign \g70516/_0_  = ~n10443 ;
  assign \g70517/_0_  = ~n10478 ;
  assign \g70518/_0_  = ~n10513 ;
  assign \g70519/_0_  = ~n10548 ;
  assign \g70521/_0_  = ~n10566 ;
  assign \g70522/_0_  = ~n10602 ;
  assign \g70524/_0_  = ~n10620 ;
  assign \g70557/_0_  = ~n10638 ;
  assign \g70559/_0_  = ~n10677 ;
  assign \g70560/_0_  = ~n10711 ;
  assign \g70561/_0_  = ~n10752 ;
  assign \g70562/_0_  = ~n10791 ;
  assign \g70563/_0_  = ~n10830 ;
  assign \g70564/_0_  = ~n10863 ;
  assign \g70565/_0_  = ~n10901 ;
  assign \g70566/_0_  = ~n10934 ;
  assign \g70567/_0_  = ~n10967 ;
  assign \g70568/_0_  = ~n11006 ;
  assign \g70569/_0_  = ~n11047 ;
  assign \g70570/_0_  = ~n11086 ;
  assign \g70571/_0_  = ~n11124 ;
  assign \g70572/_0_  = ~n11157 ;
  assign \g70573/_0_  = ~n11198 ;
  assign \g70574/_0_  = ~n11237 ;
  assign \g70575/_0_  = ~n11275 ;
  assign \g70576/_0_  = ~n11314 ;
  assign \g70577/_0_  = ~n11355 ;
  assign \g70578/_0_  = ~n11388 ;
  assign \g70579/_0_  = ~n11429 ;
  assign \g70580/_0_  = ~n11463 ;
  assign \g70581/_0_  = ~n11502 ;
  assign \g70582/_0_  = ~n11535 ;
  assign \g70583/_0_  = ~n11576 ;
  assign \g70584/_0_  = ~n11615 ;
  assign \g70585/_0_  = ~n11654 ;
  assign \g70586/_0_  = ~n11692 ;
  assign \g70587/_0_  = ~n11733 ;
  assign \g70588/_0_  = ~n11766 ;
  assign \g70589/_0_  = ~n11803 ;
  assign \g70590/_0_  = ~n11832 ;
  assign \g70591/_0_  = ~n11865 ;
  assign \g70592/_0_  = ~n11902 ;
  assign \g70593/_0_  = ~n11933 ;
  assign \g70594/_0_  = ~n11973 ;
  assign \g70595/_0_  = ~n12004 ;
  assign \g70596/_0_  = ~n12041 ;
  assign \g70597/_0_  = ~n12078 ;
  assign \g70598/_0_  = ~n12109 ;
  assign \g70599/_0_  = ~n12130 ;
  assign \g70600/_0_  = ~n12151 ;
  assign \g70601/_0_  = n12178 ;
  assign \g70602/_0_  = ~n12199 ;
  assign \g70603/_0_  = ~n12220 ;
  assign \g70604/_0_  = ~n12241 ;
  assign \g70605/_0_  = n12245 ;
  assign \g70606/_0_  = ~n12273 ;
  assign \g70607/_0_  = ~n12300 ;
  assign \g70608/_0_  = ~n12327 ;
  assign \g70609/_0_  = ~n12354 ;
  assign \g70610/_0_  = ~n12381 ;
  assign \g70611/_0_  = ~n12408 ;
  assign \g70612/_0_  = ~n12435 ;
  assign \g70613/_0_  = ~n12462 ;
  assign \g70614/_0_  = ~n12489 ;
  assign \g70615/_0_  = ~n12516 ;
  assign \g70616/_0_  = ~n12543 ;
  assign \g70617/_0_  = ~n12570 ;
  assign \g70618/_0_  = ~n12597 ;
  assign \g70619/_0_  = ~n12624 ;
  assign \g70620/_0_  = ~n12651 ;
  assign \g70621/_0_  = ~n12678 ;
  assign \g70622/_0_  = ~n12682 ;
  assign \g70623/_0_  = ~n12685 ;
  assign \g70624/_0_  = ~n12688 ;
  assign \g70625/_0_  = ~n12691 ;
  assign \g70626/_0_  = ~n12694 ;
  assign \g70627/_0_  = ~n12697 ;
  assign \g70628/_0_  = ~n12700 ;
  assign \g70629/_0_  = ~n12703 ;
  assign \g70630/_0_  = ~n12706 ;
  assign \g70631/_0_  = ~n12709 ;
  assign \g70632/_0_  = ~n12712 ;
  assign \g70633/_0_  = ~n12715 ;
  assign \g70634/_0_  = ~n12718 ;
  assign \g70635/_0_  = ~n12721 ;
  assign \g70636/_0_  = ~n12724 ;
  assign \g70637/_0_  = ~n12727 ;
  assign \g70638/_0_  = ~n12731 ;
  assign \g70639/_0_  = ~n12734 ;
  assign \g70640/_0_  = ~n12737 ;
  assign \g70641/_0_  = ~n12740 ;
  assign \g70642/_0_  = ~n12743 ;
  assign \g70643/_0_  = ~n12746 ;
  assign \g70644/_0_  = ~n12749 ;
  assign \g70645/_0_  = ~n12752 ;
  assign \g70646/_0_  = ~n12755 ;
  assign \g70647/_0_  = ~n12758 ;
  assign \g70648/_0_  = ~n12761 ;
  assign \g70649/_0_  = ~n12764 ;
  assign \g70650/_0_  = ~n12767 ;
  assign \g70651/_0_  = ~n12770 ;
  assign \g70652/_0_  = ~n12773 ;
  assign \g70653/_0_  = ~n12776 ;
  assign \g70654/_0_  = ~n12780 ;
  assign \g70655/_0_  = ~n12783 ;
  assign \g70656/_0_  = ~n12786 ;
  assign \g70657/_0_  = ~n12789 ;
  assign \g70658/_0_  = ~n12792 ;
  assign \g70659/_0_  = ~n12795 ;
  assign \g70660/_0_  = ~n12798 ;
  assign \g70661/_0_  = ~n12801 ;
  assign \g70662/_0_  = ~n12804 ;
  assign \g70663/_0_  = ~n12807 ;
  assign \g70664/_0_  = ~n12810 ;
  assign \g70665/_0_  = ~n12813 ;
  assign \g70666/_0_  = ~n12816 ;
  assign \g70667/_0_  = ~n12819 ;
  assign \g70668/_0_  = ~n12822 ;
  assign \g70669/_0_  = ~n12825 ;
  assign \g70670/_0_  = ~n12829 ;
  assign \g70671/_0_  = ~n12832 ;
  assign \g70672/_0_  = ~n12835 ;
  assign \g70673/_0_  = ~n12838 ;
  assign \g70674/_0_  = ~n12841 ;
  assign \g70675/_0_  = ~n12844 ;
  assign \g70676/_0_  = ~n12847 ;
  assign \g70677/_0_  = ~n12850 ;
  assign \g70678/_0_  = ~n12853 ;
  assign \g70679/_0_  = ~n12856 ;
  assign \g70680/_0_  = ~n12859 ;
  assign \g70681/_0_  = ~n12862 ;
  assign \g70682/_0_  = ~n12865 ;
  assign \g70683/_0_  = ~n12868 ;
  assign \g70684/_0_  = ~n12871 ;
  assign \g70685/_0_  = ~n12874 ;
  assign \g70686/_0_  = ~n12878 ;
  assign \g70687/_0_  = ~n12881 ;
  assign \g70688/_0_  = ~n12884 ;
  assign \g70689/_0_  = ~n12887 ;
  assign \g70690/_0_  = ~n12890 ;
  assign \g70691/_0_  = ~n12893 ;
  assign \g70692/_0_  = ~n12896 ;
  assign \g70693/_0_  = ~n12899 ;
  assign \g70694/_0_  = ~n12902 ;
  assign \g70695/_0_  = ~n12905 ;
  assign \g70696/_0_  = ~n12908 ;
  assign \g70697/_0_  = ~n12911 ;
  assign \g70698/_0_  = ~n12914 ;
  assign \g70699/_0_  = ~n12917 ;
  assign \g70700/_0_  = ~n12920 ;
  assign \g70701/_0_  = ~n12923 ;
  assign \g70702/_0_  = ~n12927 ;
  assign \g70703/_0_  = ~n12930 ;
  assign \g70704/_0_  = ~n12933 ;
  assign \g70705/_0_  = ~n12936 ;
  assign \g70706/_0_  = ~n12939 ;
  assign \g70707/_0_  = ~n12942 ;
  assign \g70708/_0_  = ~n12945 ;
  assign \g70709/_0_  = ~n12948 ;
  assign \g70710/_0_  = ~n12951 ;
  assign \g70711/_0_  = ~n12954 ;
  assign \g70712/_0_  = ~n12957 ;
  assign \g70713/_0_  = ~n12960 ;
  assign \g70714/_0_  = ~n12963 ;
  assign \g70715/_0_  = ~n12966 ;
  assign \g70716/_0_  = ~n12969 ;
  assign \g70717/_0_  = ~n12972 ;
  assign \g70718/_0_  = ~n12976 ;
  assign \g70719/_0_  = ~n12979 ;
  assign \g70720/_0_  = ~n12982 ;
  assign \g70721/_0_  = ~n12985 ;
  assign \g70722/_0_  = ~n12988 ;
  assign \g70723/_0_  = ~n12991 ;
  assign \g70724/_0_  = ~n12994 ;
  assign \g70725/_0_  = ~n12997 ;
  assign \g70726/_0_  = ~n13000 ;
  assign \g70727/_0_  = ~n13003 ;
  assign \g70728/_0_  = ~n13006 ;
  assign \g70729/_0_  = ~n13009 ;
  assign \g70730/_0_  = ~n13012 ;
  assign \g70731/_0_  = ~n13015 ;
  assign \g70732/_0_  = ~n13018 ;
  assign \g70733/_0_  = ~n13021 ;
  assign \g70734/_0_  = ~n13025 ;
  assign \g70735/_0_  = ~n13028 ;
  assign \g70736/_0_  = ~n13031 ;
  assign \g70737/_0_  = ~n13034 ;
  assign \g70738/_0_  = ~n13037 ;
  assign \g70739/_0_  = ~n13040 ;
  assign \g70740/_0_  = ~n13043 ;
  assign \g70741/_0_  = ~n13046 ;
  assign \g70742/_0_  = ~n13049 ;
  assign \g70743/_0_  = ~n13052 ;
  assign \g70744/_0_  = ~n13055 ;
  assign \g70745/_0_  = ~n13058 ;
  assign \g70746/_0_  = ~n13061 ;
  assign \g70747/_0_  = ~n13064 ;
  assign \g70748/_0_  = ~n13067 ;
  assign \g70749/_0_  = ~n13070 ;
  assign \g70750/_0_  = ~n13074 ;
  assign \g70751/_0_  = ~n13077 ;
  assign \g70752/_0_  = ~n13080 ;
  assign \g70753/_0_  = ~n13083 ;
  assign \g70754/_0_  = ~n13086 ;
  assign \g70755/_0_  = ~n13089 ;
  assign \g70756/_0_  = ~n13092 ;
  assign \g70757/_0_  = ~n13095 ;
  assign \g70758/_0_  = ~n13098 ;
  assign \g70759/_0_  = ~n13101 ;
  assign \g70760/_0_  = ~n13104 ;
  assign \g70761/_0_  = ~n13107 ;
  assign \g70762/_0_  = ~n13110 ;
  assign \g70763/_0_  = ~n13113 ;
  assign \g70764/_0_  = ~n13116 ;
  assign \g70765/_0_  = ~n13119 ;
  assign \g70766/_0_  = ~n13123 ;
  assign \g70767/_0_  = ~n13126 ;
  assign \g70768/_0_  = ~n13129 ;
  assign \g70769/_0_  = ~n13132 ;
  assign \g70770/_0_  = ~n13135 ;
  assign \g70771/_0_  = ~n13138 ;
  assign \g70772/_0_  = ~n13141 ;
  assign \g70773/_0_  = ~n13144 ;
  assign \g70774/_0_  = ~n13147 ;
  assign \g70775/_0_  = ~n13150 ;
  assign \g70776/_0_  = ~n13153 ;
  assign \g70777/_0_  = ~n13156 ;
  assign \g70778/_0_  = ~n13159 ;
  assign \g70779/_0_  = ~n13162 ;
  assign \g70780/_0_  = ~n13165 ;
  assign \g70781/_0_  = ~n13168 ;
  assign \g70782/_0_  = ~n13172 ;
  assign \g70783/_0_  = ~n13175 ;
  assign \g70784/_0_  = ~n13178 ;
  assign \g70785/_0_  = ~n13181 ;
  assign \g70786/_0_  = ~n13184 ;
  assign \g70787/_0_  = ~n13187 ;
  assign \g70788/_0_  = ~n13190 ;
  assign \g70789/_0_  = ~n13193 ;
  assign \g70790/_0_  = ~n13196 ;
  assign \g70791/_0_  = ~n13199 ;
  assign \g70792/_0_  = ~n13202 ;
  assign \g70793/_0_  = ~n13205 ;
  assign \g70794/_0_  = ~n13208 ;
  assign \g70795/_0_  = ~n13211 ;
  assign \g70796/_0_  = ~n13214 ;
  assign \g70797/_0_  = ~n13217 ;
  assign \g70798/_0_  = ~n13221 ;
  assign \g70799/_0_  = ~n13224 ;
  assign \g70800/_0_  = ~n13227 ;
  assign \g70801/_0_  = ~n13230 ;
  assign \g70802/_0_  = ~n13233 ;
  assign \g70803/_0_  = ~n13236 ;
  assign \g70804/_0_  = ~n13239 ;
  assign \g70805/_0_  = ~n13242 ;
  assign \g70806/_0_  = ~n13245 ;
  assign \g70807/_0_  = ~n13248 ;
  assign \g70808/_0_  = ~n13251 ;
  assign \g70809/_0_  = ~n13254 ;
  assign \g70810/_0_  = ~n13257 ;
  assign \g70811/_0_  = ~n13260 ;
  assign \g70812/_0_  = ~n13263 ;
  assign \g70813/_0_  = ~n13266 ;
  assign \g70814/_0_  = ~n13270 ;
  assign \g70815/_0_  = ~n13273 ;
  assign \g70816/_0_  = ~n13276 ;
  assign \g70817/_0_  = ~n13279 ;
  assign \g70818/_0_  = ~n13282 ;
  assign \g70819/_0_  = ~n13285 ;
  assign \g70820/_0_  = ~n13288 ;
  assign \g70821/_0_  = ~n13291 ;
  assign \g70822/_0_  = ~n13294 ;
  assign \g70823/_0_  = ~n13297 ;
  assign \g70824/_0_  = ~n13300 ;
  assign \g70825/_0_  = ~n13303 ;
  assign \g70826/_0_  = ~n13306 ;
  assign \g70827/_0_  = ~n13309 ;
  assign \g70828/_0_  = ~n13312 ;
  assign \g70829/_0_  = ~n13315 ;
  assign \g70830/_0_  = ~n13319 ;
  assign \g70831/_0_  = ~n13322 ;
  assign \g70832/_0_  = ~n13325 ;
  assign \g70833/_0_  = ~n13328 ;
  assign \g70834/_0_  = ~n13331 ;
  assign \g70835/_0_  = ~n13334 ;
  assign \g70836/_0_  = ~n13337 ;
  assign \g70837/_0_  = ~n13340 ;
  assign \g70838/_0_  = ~n13343 ;
  assign \g70839/_0_  = ~n13346 ;
  assign \g70840/_0_  = ~n13349 ;
  assign \g70841/_0_  = ~n13352 ;
  assign \g70842/_0_  = ~n13355 ;
  assign \g70843/_0_  = ~n13358 ;
  assign \g70844/_0_  = ~n13361 ;
  assign \g70845/_0_  = ~n13364 ;
  assign \g70846/_0_  = ~n13368 ;
  assign \g70847/_0_  = ~n13371 ;
  assign \g70848/_0_  = ~n13374 ;
  assign \g70849/_0_  = ~n13377 ;
  assign \g70850/_0_  = ~n13380 ;
  assign \g70851/_0_  = ~n13383 ;
  assign \g70852/_0_  = ~n13386 ;
  assign \g70853/_0_  = ~n13389 ;
  assign \g70854/_0_  = ~n13392 ;
  assign \g70855/_0_  = ~n13395 ;
  assign \g70856/_0_  = ~n13398 ;
  assign \g70857/_0_  = ~n13401 ;
  assign \g70858/_0_  = ~n13404 ;
  assign \g70859/_0_  = ~n13407 ;
  assign \g70860/_0_  = ~n13410 ;
  assign \g70861/_0_  = ~n13413 ;
  assign \g71404/_0_  = n13416 ;
  assign \g71407/_0_  = n13441 ;
  assign \g72631/_0_  = n13501 ;
  assign \g72631/_1_  = ~n13501 ;
  assign \g72633/_0_  = n13511 ;
  assign \g72642/_0_  = n13521 ;
  assign \g72649/_0_  = n13581 ;
  assign \g72649/_1_  = ~n13581 ;
  assign \g72652/_0_  = n13591 ;
  assign \g72660/_0_  = n13601 ;
  assign \g72666/_0_  = n13661 ;
  assign \g72666/_1_  = ~n13661 ;
  assign \g72671/_0_  = n13671 ;
  assign \g72681/_0_  = n13731 ;
  assign \g72681/_1_  = ~n13731 ;
  assign \g72689/_0_  = n13741 ;
  assign \g72696/_0_  = n13801 ;
  assign \g72696/_1_  = ~n13801 ;
  assign \g72698/_0_  = n13811 ;
  assign \g72707/_0_  = n13821 ;
  assign \g72715/_0_  = n13881 ;
  assign \g72715/_1_  = ~n13881 ;
  assign \g72718/_0_  = n13891 ;
  assign \g72726/_0_  = n13902 ;
  assign \g72732/_0_  = n13962 ;
  assign \g72732/_1_  = ~n13962 ;
  assign \g72736/_0_  = n13973 ;
  assign \g72743/_0_  = n13983 ;
  assign \g72745/_0_  = n14043 ;
  assign \g72745/_1_  = ~n14043 ;
  assign \g72752/_0_  = n14103 ;
  assign \g72752/_1_  = ~n14103 ;
  assign \g72756/_0_  = n14114 ;
  assign \g72763/_0_  = n14174 ;
  assign \g72763/_1_  = ~n14174 ;
  assign \g72765/_0_  = n14185 ;
  assign \g72767/_0_  = n14245 ;
  assign \g72767/_1_  = ~n14245 ;
  assign \g72769/_0_  = n14305 ;
  assign \g72769/_1_  = ~n14305 ;
  assign \g72772/_0_  = n14365 ;
  assign \g72772/_1_  = ~n14365 ;
  assign \g72774/_0_  = n14425 ;
  assign \g72774/_1_  = ~n14425 ;
  assign \g72790/_0_  = n14485 ;
  assign \g72790/_1_  = ~n14485 ;
  assign \g72797/_0_  = n14496 ;
  assign \g73807/_0_  = n14500 ;
  assign \g73820/_0_  = n14504 ;
  assign \g73832/_0_  = n14508 ;
  assign \g73844/_0_  = n14512 ;
  assign \g73856/_0_  = n14516 ;
  assign \g73871/_0_  = n14520 ;
  assign \g73883/_0_  = n14524 ;
  assign \g73895/_0_  = n14528 ;
  assign \g73905/_3_  = n2106 ;
  assign \g73910/_0_  = n14532 ;
  assign \g73922/_0_  = n14536 ;
  assign \g73934/_0_  = n14540 ;
  assign \g73946/_0_  = n14544 ;
  assign \g73958/_0_  = n14548 ;
  assign \g73970/_0_  = n14552 ;
  assign \g73982/_0_  = n14556 ;
  assign \g87036/_0_  = ~n14564 ;
  assign \g87042/_0_  = ~n14572 ;
  assign \g87043/_0_  = ~n14577 ;
  assign \g87044/_0_  = ~n14585 ;
  assign \g87045/_0_  = ~n14593 ;
  assign \g87046/_0_  = ~n14598 ;
  assign \g87047/_0_  = ~n14606 ;
  assign \g87048/_0_  = ~n14611 ;
  assign \g87049/_0_  = ~n14619 ;
  assign \g87050/_0_  = ~n14624 ;
  assign \g87051/_0_  = ~n14629 ;
  assign \g87052/_0_  = ~n14637 ;
  assign \g87053/_0_  = ~n14642 ;
  assign \g87054/_0_  = ~n14650 ;
  assign \g87055/_0_  = ~n14655 ;
  assign \g87062/_0_  = ~n14660 ;
  assign \g88572/_0_  = ~n14663 ;
  assign \g88681/_0_  = ~n14668 ;
  assign \g88682/_0_  = ~n14673 ;
  assign \g88683/_0_  = ~n14677 ;
  assign \g88684/_0_  = ~n14683 ;
  assign \g88685/_0_  = ~n14687 ;
  assign \g88686/_0_  = ~n14692 ;
  assign \g88687/_0_  = ~n14697 ;
  assign \g88688/_0_  = ~n14702 ;
  assign \g88689/_0_  = ~n14706 ;
  assign \g88690/_0_  = ~n14710 ;
  assign \g88691/_0_  = ~n14715 ;
  assign \g88692/_0_  = ~n14719 ;
  assign \g88693/_0_  = ~n14725 ;
  assign \g88695/_0_  = ~n14729 ;
  assign \g88697/_0_  = ~n14733 ;
  assign \g88698/_0_  = ~n14737 ;
  assign \g88700/_0_  = ~n14742 ;
  assign \g88701/_0_  = ~n14747 ;
  assign \g88703/_0_  = ~n14751 ;
  assign \g88704/_0_  = ~n14755 ;
  assign \g88705/_0_  = ~n14759 ;
  assign \g88706/_0_  = ~n14764 ;
  assign \g88707/_0_  = ~n14767 ;
  assign \g88709/_0_  = ~n14772 ;
  assign \g88710/_0_  = ~n14776 ;
  assign \g88711/_0_  = ~n14780 ;
  assign \g88712/_0_  = ~n14784 ;
  assign \g88713/_0_  = ~n14788 ;
  assign \g88714/_0_  = ~n14793 ;
  assign \g88716/_0_  = ~n14799 ;
  assign \g88717/_0_  = ~n14803 ;
  assign \g88718/_0_  = ~n14807 ;
  assign \g88719/_0_  = ~n14811 ;
  assign \g88720/_0_  = ~n14814 ;
  assign \g88722/_0_  = ~n14818 ;
  assign \g88723/_0_  = ~n14822 ;
  assign \g88724/_0_  = ~n14827 ;
  assign \g88725/_0_  = ~n14831 ;
  assign \g88726/_0_  = ~n14835 ;
  assign \g88727/_0_  = ~n14839 ;
  assign \g88728/_0_  = ~n14843 ;
  assign \g88729/_0_  = ~n14847 ;
  assign \g88731/_0_  = ~n14853 ;
  assign \g88732/_0_  = ~n14857 ;
  assign \g88733/_0_  = ~n14861 ;
  assign \g88734/_0_  = ~n14864 ;
  assign \g88736/_0_  = ~n14868 ;
  assign \g88737/_0_  = ~n14872 ;
  assign \g88738/_0_  = ~n14877 ;
  assign \g88739/_0_  = ~n14881 ;
  assign \g88740/_0_  = ~n14885 ;
  assign \g88741/_0_  = ~n14889 ;
  assign \g88742/_0_  = ~n14894 ;
  assign \g88743/_0_  = ~n14898 ;
  assign \g88744/_0_  = ~n14902 ;
  assign \g88745/_0_  = ~n14906 ;
  assign \g88746/_0_  = ~n14909 ;
  assign \g88748/_0_  = ~n14913 ;
  assign \g88749/_0_  = ~n14917 ;
  assign \g88750/_0_  = ~n14921 ;
  assign \g88752/_0_  = ~n14925 ;
  assign \g88753/_0_  = ~n14929 ;
  assign \g88754/_0_  = ~n14933 ;
  assign \g88755/_0_  = ~n14937 ;
  assign \g88756/_0_  = ~n14941 ;
  assign \g88757/_0_  = ~n14944 ;
  assign \g88759/_0_  = ~n14948 ;
  assign \g88760/_0_  = ~n14952 ;
  assign \g88761/_0_  = ~n14956 ;
  assign \g88762/_0_  = ~n14960 ;
  assign \g88764/_0_  = ~n14965 ;
  assign \g88765/_0_  = ~n14969 ;
  assign \g88766/_0_  = ~n14973 ;
  assign \g88768/_0_  = ~n14977 ;
  assign \g88769/_0_  = ~n14981 ;
  assign \g88770/_0_  = ~n14985 ;
  assign \g88771/_0_  = ~n14989 ;
  assign \g88772/_0_  = ~n14993 ;
  assign \g88773/_0_  = ~n14997 ;
  assign \g88775/_0_  = ~n15001 ;
  assign \g88776/_0_  = ~n15005 ;
  assign \g88777/_0_  = ~n15009 ;
  assign \g88778/_0_  = ~n15013 ;
  assign \g88779/_0_  = ~n15017 ;
  assign \g88780/_0_  = ~n15020 ;
  assign \g88782/_0_  = ~n15024 ;
  assign \g88783/_0_  = ~n15028 ;
  assign \g88784/_0_  = ~n15032 ;
  assign \g88785/_0_  = ~n15036 ;
  assign \g88786/_0_  = ~n15040 ;
  assign \g88787/_0_  = ~n15044 ;
  assign \g88789/_0_  = ~n15049 ;
  assign \g88790/_0_  = ~n15053 ;
  assign \g88791/_0_  = ~n15057 ;
  assign \g88792/_0_  = ~n15061 ;
  assign \g88793/_0_  = ~n15064 ;
  assign \g88795/_0_  = ~n15068 ;
  assign \g88796/_0_  = ~n15072 ;
  assign \g88797/_0_  = ~n15076 ;
  assign \g88799/_0_  = ~n15080 ;
  assign \g88800/_0_  = ~n15084 ;
  assign \g88801/_0_  = ~n15088 ;
  assign \g88802/_0_  = ~n15092 ;
  assign \g88806/_0_  = ~n15096 ;
  assign \g88807/_0_  = ~n15100 ;
  assign \g88808/_0_  = ~n15104 ;
  assign \g88809/_0_  = ~n15108 ;
  assign \g88810/_0_  = ~n15112 ;
  assign \g88813/_0_  = ~n15116 ;
  assign \g88814/_0_  = ~n15120 ;
  assign \g88815/_0_  = ~n15124 ;
  assign \m0_ack_o_pad  = ~n15189 ;
  assign \m0_data_o[0]_pad  = ~n15226 ;
  assign \m0_data_o[10]_pad  = ~n15263 ;
  assign \m0_data_o[11]_pad  = ~n15300 ;
  assign \m0_data_o[12]_pad  = ~n15337 ;
  assign \m0_data_o[13]_pad  = ~n15374 ;
  assign \m0_data_o[14]_pad  = ~n15411 ;
  assign \m0_data_o[15]_pad  = ~n15448 ;
  assign \m0_data_o[16]_pad  = ~n15480 ;
  assign \m0_data_o[17]_pad  = ~n15512 ;
  assign \m0_data_o[18]_pad  = ~n15544 ;
  assign \m0_data_o[19]_pad  = ~n15576 ;
  assign \m0_data_o[1]_pad  = ~n15613 ;
  assign \m0_data_o[20]_pad  = ~n15645 ;
  assign \m0_data_o[21]_pad  = ~n15677 ;
  assign \m0_data_o[22]_pad  = ~n15709 ;
  assign \m0_data_o[23]_pad  = ~n15741 ;
  assign \m0_data_o[24]_pad  = ~n15773 ;
  assign \m0_data_o[25]_pad  = ~n15805 ;
  assign \m0_data_o[26]_pad  = ~n15837 ;
  assign \m0_data_o[27]_pad  = ~n15869 ;
  assign \m0_data_o[28]_pad  = ~n15901 ;
  assign \m0_data_o[29]_pad  = ~n15933 ;
  assign \m0_data_o[2]_pad  = ~n15970 ;
  assign \m0_data_o[30]_pad  = ~n16002 ;
  assign \m0_data_o[31]_pad  = ~n16034 ;
  assign \m0_data_o[3]_pad  = ~n16071 ;
  assign \m0_data_o[4]_pad  = ~n16108 ;
  assign \m0_data_o[5]_pad  = ~n16145 ;
  assign \m0_data_o[6]_pad  = ~n16182 ;
  assign \m0_data_o[7]_pad  = ~n16219 ;
  assign \m0_data_o[8]_pad  = ~n16256 ;
  assign \m0_data_o[9]_pad  = ~n16293 ;
  assign \m0_err_o_pad  = ~n16355 ;
  assign \m0_rty_o_pad  = ~n16417 ;
  assign \m1_ack_o_pad  = ~n16481 ;
  assign \m1_data_o[0]_pad  = ~n16515 ;
  assign \m1_data_o[10]_pad  = ~n16549 ;
  assign \m1_data_o[11]_pad  = ~n16583 ;
  assign \m1_data_o[12]_pad  = ~n16617 ;
  assign \m1_data_o[13]_pad  = ~n16651 ;
  assign \m1_data_o[14]_pad  = ~n16685 ;
  assign \m1_data_o[15]_pad  = ~n16719 ;
  assign \m1_data_o[16]_pad  = ~n16751 ;
  assign \m1_data_o[17]_pad  = ~n16783 ;
  assign \m1_data_o[18]_pad  = ~n16815 ;
  assign \m1_data_o[19]_pad  = ~n16847 ;
  assign \m1_data_o[1]_pad  = ~n16881 ;
  assign \m1_data_o[20]_pad  = ~n16913 ;
  assign \m1_data_o[21]_pad  = ~n16945 ;
  assign \m1_data_o[22]_pad  = ~n16977 ;
  assign \m1_data_o[23]_pad  = ~n17009 ;
  assign \m1_data_o[24]_pad  = ~n17041 ;
  assign \m1_data_o[25]_pad  = ~n17073 ;
  assign \m1_data_o[26]_pad  = ~n17105 ;
  assign \m1_data_o[27]_pad  = ~n17137 ;
  assign \m1_data_o[28]_pad  = ~n17169 ;
  assign \m1_data_o[29]_pad  = ~n17201 ;
  assign \m1_data_o[2]_pad  = ~n17235 ;
  assign \m1_data_o[30]_pad  = ~n17267 ;
  assign \m1_data_o[31]_pad  = ~n17299 ;
  assign \m1_data_o[3]_pad  = ~n17333 ;
  assign \m1_data_o[4]_pad  = ~n17367 ;
  assign \m1_data_o[5]_pad  = ~n17401 ;
  assign \m1_data_o[6]_pad  = ~n17435 ;
  assign \m1_data_o[7]_pad  = ~n17469 ;
  assign \m1_data_o[8]_pad  = ~n17503 ;
  assign \m1_data_o[9]_pad  = ~n17537 ;
  assign \m1_err_o_pad  = ~n17599 ;
  assign \m1_rty_o_pad  = ~n17661 ;
  assign \m2_ack_o_pad  = ~n17725 ;
  assign \m2_data_o[0]_pad  = ~n17759 ;
  assign \m2_data_o[10]_pad  = ~n17793 ;
  assign \m2_data_o[11]_pad  = ~n17827 ;
  assign \m2_data_o[12]_pad  = ~n17861 ;
  assign \m2_data_o[13]_pad  = ~n17895 ;
  assign \m2_data_o[14]_pad  = ~n17929 ;
  assign \m2_data_o[15]_pad  = ~n17963 ;
  assign \m2_data_o[16]_pad  = ~n17995 ;
  assign \m2_data_o[17]_pad  = ~n18027 ;
  assign \m2_data_o[18]_pad  = ~n18059 ;
  assign \m2_data_o[19]_pad  = ~n18091 ;
  assign \m2_data_o[1]_pad  = ~n18125 ;
  assign \m2_data_o[20]_pad  = ~n18157 ;
  assign \m2_data_o[21]_pad  = ~n18189 ;
  assign \m2_data_o[22]_pad  = ~n18221 ;
  assign \m2_data_o[23]_pad  = ~n18253 ;
  assign \m2_data_o[24]_pad  = ~n18285 ;
  assign \m2_data_o[25]_pad  = ~n18317 ;
  assign \m2_data_o[26]_pad  = ~n18349 ;
  assign \m2_data_o[27]_pad  = ~n18381 ;
  assign \m2_data_o[28]_pad  = ~n18413 ;
  assign \m2_data_o[29]_pad  = ~n18445 ;
  assign \m2_data_o[2]_pad  = ~n18479 ;
  assign \m2_data_o[30]_pad  = ~n18511 ;
  assign \m2_data_o[31]_pad  = ~n18543 ;
  assign \m2_data_o[3]_pad  = ~n18577 ;
  assign \m2_data_o[4]_pad  = ~n18611 ;
  assign \m2_data_o[5]_pad  = ~n18645 ;
  assign \m2_data_o[6]_pad  = ~n18679 ;
  assign \m2_data_o[7]_pad  = ~n18713 ;
  assign \m2_data_o[8]_pad  = ~n18747 ;
  assign \m2_data_o[9]_pad  = ~n18781 ;
  assign \m2_err_o_pad  = ~n18843 ;
  assign \m2_rty_o_pad  = ~n18905 ;
  assign \m3_ack_o_pad  = ~n18969 ;
  assign \m3_data_o[0]_pad  = ~n19003 ;
  assign \m3_data_o[10]_pad  = ~n19037 ;
  assign \m3_data_o[11]_pad  = ~n19071 ;
  assign \m3_data_o[12]_pad  = ~n19105 ;
  assign \m3_data_o[13]_pad  = ~n19139 ;
  assign \m3_data_o[14]_pad  = ~n19173 ;
  assign \m3_data_o[15]_pad  = ~n19207 ;
  assign \m3_data_o[16]_pad  = ~n19239 ;
  assign \m3_data_o[17]_pad  = ~n19271 ;
  assign \m3_data_o[18]_pad  = ~n19303 ;
  assign \m3_data_o[19]_pad  = ~n19335 ;
  assign \m3_data_o[1]_pad  = ~n19369 ;
  assign \m3_data_o[20]_pad  = ~n19401 ;
  assign \m3_data_o[21]_pad  = ~n19433 ;
  assign \m3_data_o[22]_pad  = ~n19465 ;
  assign \m3_data_o[23]_pad  = ~n19497 ;
  assign \m3_data_o[24]_pad  = ~n19529 ;
  assign \m3_data_o[25]_pad  = ~n19561 ;
  assign \m3_data_o[26]_pad  = ~n19593 ;
  assign \m3_data_o[27]_pad  = ~n19625 ;
  assign \m3_data_o[28]_pad  = ~n19657 ;
  assign \m3_data_o[29]_pad  = ~n19689 ;
  assign \m3_data_o[2]_pad  = ~n19723 ;
  assign \m3_data_o[30]_pad  = ~n19755 ;
  assign \m3_data_o[31]_pad  = ~n19787 ;
  assign \m3_data_o[3]_pad  = ~n19821 ;
  assign \m3_data_o[4]_pad  = ~n19855 ;
  assign \m3_data_o[5]_pad  = ~n19889 ;
  assign \m3_data_o[6]_pad  = ~n19923 ;
  assign \m3_data_o[7]_pad  = ~n19957 ;
  assign \m3_data_o[8]_pad  = ~n19991 ;
  assign \m3_data_o[9]_pad  = ~n20025 ;
  assign \m3_err_o_pad  = ~n20087 ;
  assign \m3_rty_o_pad  = ~n20149 ;
  assign \m4_ack_o_pad  = ~n20213 ;
  assign \m4_data_o[0]_pad  = ~n20247 ;
  assign \m4_data_o[10]_pad  = ~n20281 ;
  assign \m4_data_o[11]_pad  = ~n20315 ;
  assign \m4_data_o[12]_pad  = ~n20349 ;
  assign \m4_data_o[13]_pad  = ~n20383 ;
  assign \m4_data_o[14]_pad  = ~n20417 ;
  assign \m4_data_o[15]_pad  = ~n20451 ;
  assign \m4_data_o[16]_pad  = ~n20483 ;
  assign \m4_data_o[17]_pad  = ~n20515 ;
  assign \m4_data_o[18]_pad  = ~n20547 ;
  assign \m4_data_o[19]_pad  = ~n20579 ;
  assign \m4_data_o[1]_pad  = ~n20613 ;
  assign \m4_data_o[20]_pad  = ~n20645 ;
  assign \m4_data_o[21]_pad  = ~n20677 ;
  assign \m4_data_o[22]_pad  = ~n20709 ;
  assign \m4_data_o[23]_pad  = ~n20741 ;
  assign \m4_data_o[24]_pad  = ~n20773 ;
  assign \m4_data_o[25]_pad  = ~n20805 ;
  assign \m4_data_o[26]_pad  = ~n20837 ;
  assign \m4_data_o[27]_pad  = ~n20869 ;
  assign \m4_data_o[28]_pad  = ~n20901 ;
  assign \m4_data_o[29]_pad  = ~n20933 ;
  assign \m4_data_o[2]_pad  = ~n20967 ;
  assign \m4_data_o[30]_pad  = ~n20999 ;
  assign \m4_data_o[31]_pad  = ~n21031 ;
  assign \m4_data_o[3]_pad  = ~n21065 ;
  assign \m4_data_o[4]_pad  = ~n21099 ;
  assign \m4_data_o[5]_pad  = ~n21133 ;
  assign \m4_data_o[6]_pad  = ~n21167 ;
  assign \m4_data_o[7]_pad  = ~n21201 ;
  assign \m4_data_o[8]_pad  = ~n21235 ;
  assign \m4_data_o[9]_pad  = ~n21269 ;
  assign \m4_err_o_pad  = ~n21331 ;
  assign \m4_rty_o_pad  = ~n21393 ;
  assign \m5_ack_o_pad  = ~n21457 ;
  assign \m5_data_o[0]_pad  = ~n21491 ;
  assign \m5_data_o[10]_pad  = ~n21525 ;
  assign \m5_data_o[11]_pad  = ~n21559 ;
  assign \m5_data_o[12]_pad  = ~n21593 ;
  assign \m5_data_o[13]_pad  = ~n21627 ;
  assign \m5_data_o[14]_pad  = ~n21661 ;
  assign \m5_data_o[15]_pad  = ~n21695 ;
  assign \m5_data_o[16]_pad  = ~n21727 ;
  assign \m5_data_o[17]_pad  = ~n21759 ;
  assign \m5_data_o[18]_pad  = ~n21791 ;
  assign \m5_data_o[19]_pad  = ~n21823 ;
  assign \m5_data_o[1]_pad  = ~n21857 ;
  assign \m5_data_o[20]_pad  = ~n21889 ;
  assign \m5_data_o[21]_pad  = ~n21921 ;
  assign \m5_data_o[22]_pad  = ~n21953 ;
  assign \m5_data_o[23]_pad  = ~n21985 ;
  assign \m5_data_o[24]_pad  = ~n22017 ;
  assign \m5_data_o[25]_pad  = ~n22049 ;
  assign \m5_data_o[26]_pad  = ~n22081 ;
  assign \m5_data_o[27]_pad  = ~n22113 ;
  assign \m5_data_o[28]_pad  = ~n22145 ;
  assign \m5_data_o[29]_pad  = ~n22177 ;
  assign \m5_data_o[2]_pad  = ~n22211 ;
  assign \m5_data_o[30]_pad  = ~n22243 ;
  assign \m5_data_o[31]_pad  = ~n22275 ;
  assign \m5_data_o[3]_pad  = ~n22309 ;
  assign \m5_data_o[4]_pad  = ~n22343 ;
  assign \m5_data_o[5]_pad  = ~n22377 ;
  assign \m5_data_o[6]_pad  = ~n22411 ;
  assign \m5_data_o[7]_pad  = ~n22445 ;
  assign \m5_data_o[8]_pad  = ~n22479 ;
  assign \m5_data_o[9]_pad  = ~n22513 ;
  assign \m5_err_o_pad  = ~n22575 ;
  assign \m5_rty_o_pad  = ~n22637 ;
  assign \m6_ack_o_pad  = ~n22701 ;
  assign \m6_data_o[0]_pad  = ~n22735 ;
  assign \m6_data_o[10]_pad  = ~n22769 ;
  assign \m6_data_o[11]_pad  = ~n22803 ;
  assign \m6_data_o[12]_pad  = ~n22837 ;
  assign \m6_data_o[13]_pad  = ~n22871 ;
  assign \m6_data_o[14]_pad  = ~n22905 ;
  assign \m6_data_o[15]_pad  = ~n22939 ;
  assign \m6_data_o[16]_pad  = ~n22971 ;
  assign \m6_data_o[17]_pad  = ~n23003 ;
  assign \m6_data_o[18]_pad  = ~n23035 ;
  assign \m6_data_o[19]_pad  = ~n23067 ;
  assign \m6_data_o[1]_pad  = ~n23101 ;
  assign \m6_data_o[20]_pad  = ~n23133 ;
  assign \m6_data_o[21]_pad  = ~n23165 ;
  assign \m6_data_o[22]_pad  = ~n23197 ;
  assign \m6_data_o[23]_pad  = ~n23229 ;
  assign \m6_data_o[24]_pad  = ~n23261 ;
  assign \m6_data_o[25]_pad  = ~n23293 ;
  assign \m6_data_o[26]_pad  = ~n23325 ;
  assign \m6_data_o[27]_pad  = ~n23357 ;
  assign \m6_data_o[28]_pad  = ~n23389 ;
  assign \m6_data_o[29]_pad  = ~n23421 ;
  assign \m6_data_o[2]_pad  = ~n23455 ;
  assign \m6_data_o[30]_pad  = ~n23487 ;
  assign \m6_data_o[31]_pad  = ~n23519 ;
  assign \m6_data_o[3]_pad  = ~n23553 ;
  assign \m6_data_o[4]_pad  = ~n23587 ;
  assign \m6_data_o[5]_pad  = ~n23621 ;
  assign \m6_data_o[6]_pad  = ~n23655 ;
  assign \m6_data_o[7]_pad  = ~n23689 ;
  assign \m6_data_o[8]_pad  = ~n23723 ;
  assign \m6_data_o[9]_pad  = ~n23757 ;
  assign \m6_err_o_pad  = ~n23819 ;
  assign \m6_rty_o_pad  = ~n23881 ;
  assign \m7_ack_o_pad  = ~n23945 ;
  assign \m7_data_o[0]_pad  = ~n23979 ;
  assign \m7_data_o[10]_pad  = ~n24013 ;
  assign \m7_data_o[11]_pad  = ~n24047 ;
  assign \m7_data_o[12]_pad  = ~n24081 ;
  assign \m7_data_o[13]_pad  = ~n24115 ;
  assign \m7_data_o[14]_pad  = ~n24149 ;
  assign \m7_data_o[15]_pad  = ~n24183 ;
  assign \m7_data_o[16]_pad  = ~n24215 ;
  assign \m7_data_o[17]_pad  = ~n24247 ;
  assign \m7_data_o[18]_pad  = ~n24279 ;
  assign \m7_data_o[19]_pad  = ~n24311 ;
  assign \m7_data_o[1]_pad  = ~n24345 ;
  assign \m7_data_o[20]_pad  = ~n24377 ;
  assign \m7_data_o[21]_pad  = ~n24409 ;
  assign \m7_data_o[22]_pad  = ~n24441 ;
  assign \m7_data_o[23]_pad  = ~n24473 ;
  assign \m7_data_o[24]_pad  = ~n24505 ;
  assign \m7_data_o[25]_pad  = ~n24537 ;
  assign \m7_data_o[26]_pad  = ~n24569 ;
  assign \m7_data_o[27]_pad  = ~n24601 ;
  assign \m7_data_o[28]_pad  = ~n24633 ;
  assign \m7_data_o[29]_pad  = ~n24665 ;
  assign \m7_data_o[2]_pad  = ~n24699 ;
  assign \m7_data_o[30]_pad  = ~n24731 ;
  assign \m7_data_o[31]_pad  = ~n24763 ;
  assign \m7_data_o[3]_pad  = ~n24797 ;
  assign \m7_data_o[4]_pad  = ~n24831 ;
  assign \m7_data_o[5]_pad  = ~n24865 ;
  assign \m7_data_o[6]_pad  = ~n24899 ;
  assign \m7_data_o[7]_pad  = ~n24933 ;
  assign \m7_data_o[8]_pad  = ~n24967 ;
  assign \m7_data_o[9]_pad  = ~n25001 ;
  assign \m7_err_o_pad  = ~n25063 ;
  assign \m7_rty_o_pad  = ~n25125 ;
  assign \s0_addr_o[0]_pad  = ~n25148 ;
  assign \s0_addr_o[10]_pad  = ~n25171 ;
  assign \s0_addr_o[11]_pad  = ~n25194 ;
  assign \s0_addr_o[12]_pad  = ~n25217 ;
  assign \s0_addr_o[13]_pad  = ~n25240 ;
  assign \s0_addr_o[14]_pad  = ~n25263 ;
  assign \s0_addr_o[15]_pad  = ~n25286 ;
  assign \s0_addr_o[16]_pad  = ~n25309 ;
  assign \s0_addr_o[17]_pad  = ~n25332 ;
  assign \s0_addr_o[18]_pad  = ~n25355 ;
  assign \s0_addr_o[19]_pad  = ~n25378 ;
  assign \s0_addr_o[1]_pad  = ~n25401 ;
  assign \s0_addr_o[20]_pad  = ~n25424 ;
  assign \s0_addr_o[21]_pad  = ~n25447 ;
  assign \s0_addr_o[22]_pad  = ~n25470 ;
  assign \s0_addr_o[23]_pad  = ~n25493 ;
  assign \s0_addr_o[24]_pad  = ~n25516 ;
  assign \s0_addr_o[25]_pad  = ~n25539 ;
  assign \s0_addr_o[26]_pad  = ~n25562 ;
  assign \s0_addr_o[27]_pad  = ~n25585 ;
  assign \s0_addr_o[28]_pad  = ~n25608 ;
  assign \s0_addr_o[29]_pad  = ~n25631 ;
  assign \s0_addr_o[2]_pad  = ~n25654 ;
  assign \s0_addr_o[30]_pad  = ~n25677 ;
  assign \s0_addr_o[31]_pad  = ~n25700 ;
  assign \s0_addr_o[3]_pad  = ~n25723 ;
  assign \s0_addr_o[4]_pad  = ~n25746 ;
  assign \s0_addr_o[5]_pad  = ~n25769 ;
  assign \s0_addr_o[6]_pad  = ~n25792 ;
  assign \s0_addr_o[7]_pad  = ~n25815 ;
  assign \s0_addr_o[8]_pad  = ~n25838 ;
  assign \s0_addr_o[9]_pad  = ~n25861 ;
  assign \s0_data_o[0]_pad  = ~n25884 ;
  assign \s0_data_o[10]_pad  = ~n25907 ;
  assign \s0_data_o[11]_pad  = ~n25930 ;
  assign \s0_data_o[12]_pad  = ~n25953 ;
  assign \s0_data_o[13]_pad  = ~n25976 ;
  assign \s0_data_o[14]_pad  = ~n25999 ;
  assign \s0_data_o[15]_pad  = ~n26022 ;
  assign \s0_data_o[16]_pad  = ~n26045 ;
  assign \s0_data_o[17]_pad  = ~n26068 ;
  assign \s0_data_o[18]_pad  = ~n26091 ;
  assign \s0_data_o[19]_pad  = ~n26114 ;
  assign \s0_data_o[1]_pad  = ~n26137 ;
  assign \s0_data_o[20]_pad  = ~n26160 ;
  assign \s0_data_o[21]_pad  = ~n26183 ;
  assign \s0_data_o[22]_pad  = ~n26206 ;
  assign \s0_data_o[23]_pad  = ~n26229 ;
  assign \s0_data_o[24]_pad  = ~n26252 ;
  assign \s0_data_o[25]_pad  = ~n26275 ;
  assign \s0_data_o[26]_pad  = ~n26298 ;
  assign \s0_data_o[27]_pad  = ~n26321 ;
  assign \s0_data_o[28]_pad  = ~n26344 ;
  assign \s0_data_o[29]_pad  = ~n26367 ;
  assign \s0_data_o[2]_pad  = ~n26390 ;
  assign \s0_data_o[30]_pad  = ~n26413 ;
  assign \s0_data_o[31]_pad  = ~n26436 ;
  assign \s0_data_o[3]_pad  = ~n26459 ;
  assign \s0_data_o[4]_pad  = ~n26482 ;
  assign \s0_data_o[5]_pad  = ~n26505 ;
  assign \s0_data_o[6]_pad  = ~n26528 ;
  assign \s0_data_o[7]_pad  = ~n26551 ;
  assign \s0_data_o[8]_pad  = ~n26574 ;
  assign \s0_data_o[9]_pad  = ~n26597 ;
  assign \s0_sel_o[0]_pad  = ~n26620 ;
  assign \s0_sel_o[1]_pad  = ~n26643 ;
  assign \s0_sel_o[2]_pad  = ~n26666 ;
  assign \s0_sel_o[3]_pad  = ~n26689 ;
  assign \s0_stb_o_pad  = ~n26720 ;
  assign \s0_we_o_pad  = ~n26743 ;
  assign \s10_addr_o[0]_pad  = ~n26766 ;
  assign \s10_addr_o[10]_pad  = ~n26789 ;
  assign \s10_addr_o[11]_pad  = ~n26812 ;
  assign \s10_addr_o[12]_pad  = ~n26835 ;
  assign \s10_addr_o[13]_pad  = ~n26858 ;
  assign \s10_addr_o[14]_pad  = ~n26881 ;
  assign \s10_addr_o[15]_pad  = ~n26904 ;
  assign \s10_addr_o[16]_pad  = ~n26927 ;
  assign \s10_addr_o[17]_pad  = ~n26950 ;
  assign \s10_addr_o[18]_pad  = ~n26973 ;
  assign \s10_addr_o[19]_pad  = ~n26996 ;
  assign \s10_addr_o[1]_pad  = ~n27019 ;
  assign \s10_addr_o[20]_pad  = ~n27042 ;
  assign \s10_addr_o[21]_pad  = ~n27065 ;
  assign \s10_addr_o[22]_pad  = ~n27088 ;
  assign \s10_addr_o[23]_pad  = ~n27111 ;
  assign \s10_addr_o[24]_pad  = ~n27134 ;
  assign \s10_addr_o[25]_pad  = ~n27157 ;
  assign \s10_addr_o[26]_pad  = ~n27180 ;
  assign \s10_addr_o[27]_pad  = ~n27203 ;
  assign \s10_addr_o[28]_pad  = ~n27226 ;
  assign \s10_addr_o[29]_pad  = ~n27249 ;
  assign \s10_addr_o[2]_pad  = ~n27272 ;
  assign \s10_addr_o[30]_pad  = ~n27295 ;
  assign \s10_addr_o[31]_pad  = ~n27318 ;
  assign \s10_addr_o[3]_pad  = ~n27341 ;
  assign \s10_addr_o[4]_pad  = ~n27364 ;
  assign \s10_addr_o[5]_pad  = ~n27387 ;
  assign \s10_addr_o[6]_pad  = ~n27410 ;
  assign \s10_addr_o[7]_pad  = ~n27433 ;
  assign \s10_addr_o[8]_pad  = ~n27456 ;
  assign \s10_addr_o[9]_pad  = ~n27479 ;
  assign \s10_data_o[0]_pad  = ~n27502 ;
  assign \s10_data_o[10]_pad  = ~n27525 ;
  assign \s10_data_o[11]_pad  = ~n27548 ;
  assign \s10_data_o[12]_pad  = ~n27571 ;
  assign \s10_data_o[13]_pad  = ~n27594 ;
  assign \s10_data_o[14]_pad  = ~n27617 ;
  assign \s10_data_o[15]_pad  = ~n27640 ;
  assign \s10_data_o[16]_pad  = ~n27663 ;
  assign \s10_data_o[17]_pad  = ~n27686 ;
  assign \s10_data_o[18]_pad  = ~n27709 ;
  assign \s10_data_o[19]_pad  = ~n27732 ;
  assign \s10_data_o[1]_pad  = ~n27755 ;
  assign \s10_data_o[20]_pad  = ~n27778 ;
  assign \s10_data_o[21]_pad  = ~n27801 ;
  assign \s10_data_o[22]_pad  = ~n27824 ;
  assign \s10_data_o[23]_pad  = ~n27847 ;
  assign \s10_data_o[24]_pad  = ~n27870 ;
  assign \s10_data_o[25]_pad  = ~n27893 ;
  assign \s10_data_o[26]_pad  = ~n27916 ;
  assign \s10_data_o[27]_pad  = ~n27939 ;
  assign \s10_data_o[28]_pad  = ~n27962 ;
  assign \s10_data_o[29]_pad  = ~n27985 ;
  assign \s10_data_o[2]_pad  = ~n28008 ;
  assign \s10_data_o[30]_pad  = ~n28031 ;
  assign \s10_data_o[31]_pad  = ~n28054 ;
  assign \s10_data_o[3]_pad  = ~n28077 ;
  assign \s10_data_o[4]_pad  = ~n28100 ;
  assign \s10_data_o[5]_pad  = ~n28123 ;
  assign \s10_data_o[6]_pad  = ~n28146 ;
  assign \s10_data_o[7]_pad  = ~n28169 ;
  assign \s10_data_o[8]_pad  = ~n28192 ;
  assign \s10_data_o[9]_pad  = ~n28215 ;
  assign \s10_sel_o[0]_pad  = ~n28238 ;
  assign \s10_sel_o[1]_pad  = ~n28261 ;
  assign \s10_sel_o[2]_pad  = ~n28284 ;
  assign \s10_sel_o[3]_pad  = ~n28307 ;
  assign \s10_stb_o_pad  = ~n28338 ;
  assign \s10_we_o_pad  = ~n28361 ;
  assign \s11_addr_o[0]_pad  = ~n28384 ;
  assign \s11_addr_o[10]_pad  = ~n28407 ;
  assign \s11_addr_o[11]_pad  = ~n28430 ;
  assign \s11_addr_o[12]_pad  = ~n28453 ;
  assign \s11_addr_o[13]_pad  = ~n28476 ;
  assign \s11_addr_o[14]_pad  = ~n28499 ;
  assign \s11_addr_o[15]_pad  = ~n28522 ;
  assign \s11_addr_o[16]_pad  = ~n28545 ;
  assign \s11_addr_o[17]_pad  = ~n28568 ;
  assign \s11_addr_o[18]_pad  = ~n28591 ;
  assign \s11_addr_o[19]_pad  = ~n28614 ;
  assign \s11_addr_o[1]_pad  = ~n28637 ;
  assign \s11_addr_o[20]_pad  = ~n28660 ;
  assign \s11_addr_o[21]_pad  = ~n28683 ;
  assign \s11_addr_o[22]_pad  = ~n28706 ;
  assign \s11_addr_o[23]_pad  = ~n28729 ;
  assign \s11_addr_o[24]_pad  = ~n28752 ;
  assign \s11_addr_o[25]_pad  = ~n28775 ;
  assign \s11_addr_o[26]_pad  = ~n28798 ;
  assign \s11_addr_o[27]_pad  = ~n28821 ;
  assign \s11_addr_o[28]_pad  = ~n28844 ;
  assign \s11_addr_o[29]_pad  = ~n28867 ;
  assign \s11_addr_o[2]_pad  = ~n28890 ;
  assign \s11_addr_o[30]_pad  = ~n28913 ;
  assign \s11_addr_o[31]_pad  = ~n28936 ;
  assign \s11_addr_o[3]_pad  = ~n28959 ;
  assign \s11_addr_o[4]_pad  = ~n28982 ;
  assign \s11_addr_o[5]_pad  = ~n29005 ;
  assign \s11_addr_o[6]_pad  = ~n29028 ;
  assign \s11_addr_o[7]_pad  = ~n29051 ;
  assign \s11_addr_o[8]_pad  = ~n29074 ;
  assign \s11_addr_o[9]_pad  = ~n29097 ;
  assign \s11_data_o[0]_pad  = ~n29120 ;
  assign \s11_data_o[10]_pad  = ~n29143 ;
  assign \s11_data_o[11]_pad  = ~n29166 ;
  assign \s11_data_o[12]_pad  = ~n29189 ;
  assign \s11_data_o[13]_pad  = ~n29212 ;
  assign \s11_data_o[14]_pad  = ~n29235 ;
  assign \s11_data_o[15]_pad  = ~n29258 ;
  assign \s11_data_o[16]_pad  = ~n29281 ;
  assign \s11_data_o[17]_pad  = ~n29304 ;
  assign \s11_data_o[18]_pad  = ~n29327 ;
  assign \s11_data_o[19]_pad  = ~n29350 ;
  assign \s11_data_o[1]_pad  = ~n29373 ;
  assign \s11_data_o[20]_pad  = ~n29396 ;
  assign \s11_data_o[21]_pad  = ~n29419 ;
  assign \s11_data_o[22]_pad  = ~n29442 ;
  assign \s11_data_o[23]_pad  = ~n29465 ;
  assign \s11_data_o[24]_pad  = ~n29488 ;
  assign \s11_data_o[25]_pad  = ~n29511 ;
  assign \s11_data_o[26]_pad  = ~n29534 ;
  assign \s11_data_o[27]_pad  = ~n29557 ;
  assign \s11_data_o[28]_pad  = ~n29580 ;
  assign \s11_data_o[29]_pad  = ~n29603 ;
  assign \s11_data_o[2]_pad  = ~n29626 ;
  assign \s11_data_o[30]_pad  = ~n29649 ;
  assign \s11_data_o[31]_pad  = ~n29672 ;
  assign \s11_data_o[3]_pad  = ~n29695 ;
  assign \s11_data_o[4]_pad  = ~n29718 ;
  assign \s11_data_o[5]_pad  = ~n29741 ;
  assign \s11_data_o[6]_pad  = ~n29764 ;
  assign \s11_data_o[7]_pad  = ~n29787 ;
  assign \s11_data_o[8]_pad  = ~n29810 ;
  assign \s11_data_o[9]_pad  = ~n29833 ;
  assign \s11_sel_o[0]_pad  = ~n29856 ;
  assign \s11_sel_o[1]_pad  = ~n29879 ;
  assign \s11_sel_o[2]_pad  = ~n29902 ;
  assign \s11_sel_o[3]_pad  = ~n29925 ;
  assign \s11_stb_o_pad  = ~n29956 ;
  assign \s11_we_o_pad  = ~n29979 ;
  assign \s12_addr_o[0]_pad  = ~n30002 ;
  assign \s12_addr_o[10]_pad  = ~n30025 ;
  assign \s12_addr_o[11]_pad  = ~n30048 ;
  assign \s12_addr_o[12]_pad  = ~n30071 ;
  assign \s12_addr_o[13]_pad  = ~n30094 ;
  assign \s12_addr_o[14]_pad  = ~n30117 ;
  assign \s12_addr_o[15]_pad  = ~n30140 ;
  assign \s12_addr_o[16]_pad  = ~n30163 ;
  assign \s12_addr_o[17]_pad  = ~n30186 ;
  assign \s12_addr_o[18]_pad  = ~n30209 ;
  assign \s12_addr_o[19]_pad  = ~n30232 ;
  assign \s12_addr_o[1]_pad  = ~n30255 ;
  assign \s12_addr_o[20]_pad  = ~n30278 ;
  assign \s12_addr_o[21]_pad  = ~n30301 ;
  assign \s12_addr_o[22]_pad  = ~n30324 ;
  assign \s12_addr_o[23]_pad  = ~n30347 ;
  assign \s12_addr_o[24]_pad  = ~n30370 ;
  assign \s12_addr_o[25]_pad  = ~n30393 ;
  assign \s12_addr_o[26]_pad  = ~n30416 ;
  assign \s12_addr_o[27]_pad  = ~n30439 ;
  assign \s12_addr_o[28]_pad  = ~n30462 ;
  assign \s12_addr_o[29]_pad  = ~n30485 ;
  assign \s12_addr_o[2]_pad  = ~n30508 ;
  assign \s12_addr_o[30]_pad  = ~n30531 ;
  assign \s12_addr_o[31]_pad  = ~n30554 ;
  assign \s12_addr_o[3]_pad  = ~n30577 ;
  assign \s12_addr_o[4]_pad  = ~n30600 ;
  assign \s12_addr_o[5]_pad  = ~n30623 ;
  assign \s12_addr_o[6]_pad  = ~n30646 ;
  assign \s12_addr_o[7]_pad  = ~n30669 ;
  assign \s12_addr_o[8]_pad  = ~n30692 ;
  assign \s12_addr_o[9]_pad  = ~n30715 ;
  assign \s12_data_o[0]_pad  = ~n30738 ;
  assign \s12_data_o[10]_pad  = ~n30761 ;
  assign \s12_data_o[11]_pad  = ~n30784 ;
  assign \s12_data_o[12]_pad  = ~n30807 ;
  assign \s12_data_o[13]_pad  = ~n30830 ;
  assign \s12_data_o[14]_pad  = ~n30853 ;
  assign \s12_data_o[15]_pad  = ~n30876 ;
  assign \s12_data_o[16]_pad  = ~n30899 ;
  assign \s12_data_o[17]_pad  = ~n30922 ;
  assign \s12_data_o[18]_pad  = ~n30945 ;
  assign \s12_data_o[19]_pad  = ~n30968 ;
  assign \s12_data_o[1]_pad  = ~n30991 ;
  assign \s12_data_o[20]_pad  = ~n31014 ;
  assign \s12_data_o[21]_pad  = ~n31037 ;
  assign \s12_data_o[22]_pad  = ~n31060 ;
  assign \s12_data_o[23]_pad  = ~n31083 ;
  assign \s12_data_o[24]_pad  = ~n31106 ;
  assign \s12_data_o[25]_pad  = ~n31129 ;
  assign \s12_data_o[26]_pad  = ~n31152 ;
  assign \s12_data_o[27]_pad  = ~n31175 ;
  assign \s12_data_o[28]_pad  = ~n31198 ;
  assign \s12_data_o[29]_pad  = ~n31221 ;
  assign \s12_data_o[2]_pad  = ~n31244 ;
  assign \s12_data_o[30]_pad  = ~n31267 ;
  assign \s12_data_o[31]_pad  = ~n31290 ;
  assign \s12_data_o[3]_pad  = ~n31313 ;
  assign \s12_data_o[4]_pad  = ~n31336 ;
  assign \s12_data_o[5]_pad  = ~n31359 ;
  assign \s12_data_o[6]_pad  = ~n31382 ;
  assign \s12_data_o[7]_pad  = ~n31405 ;
  assign \s12_data_o[8]_pad  = ~n31428 ;
  assign \s12_data_o[9]_pad  = ~n31451 ;
  assign \s12_sel_o[0]_pad  = ~n31474 ;
  assign \s12_sel_o[1]_pad  = ~n31497 ;
  assign \s12_sel_o[2]_pad  = ~n31520 ;
  assign \s12_sel_o[3]_pad  = ~n31543 ;
  assign \s12_stb_o_pad  = ~n31574 ;
  assign \s12_we_o_pad  = ~n31597 ;
  assign \s13_addr_o[0]_pad  = ~n31620 ;
  assign \s13_addr_o[10]_pad  = ~n31643 ;
  assign \s13_addr_o[11]_pad  = ~n31666 ;
  assign \s13_addr_o[12]_pad  = ~n31689 ;
  assign \s13_addr_o[13]_pad  = ~n31712 ;
  assign \s13_addr_o[14]_pad  = ~n31735 ;
  assign \s13_addr_o[15]_pad  = ~n31758 ;
  assign \s13_addr_o[16]_pad  = ~n31781 ;
  assign \s13_addr_o[17]_pad  = ~n31804 ;
  assign \s13_addr_o[18]_pad  = ~n31827 ;
  assign \s13_addr_o[19]_pad  = ~n31850 ;
  assign \s13_addr_o[1]_pad  = ~n31873 ;
  assign \s13_addr_o[20]_pad  = ~n31896 ;
  assign \s13_addr_o[21]_pad  = ~n31919 ;
  assign \s13_addr_o[22]_pad  = ~n31942 ;
  assign \s13_addr_o[23]_pad  = ~n31965 ;
  assign \s13_addr_o[24]_pad  = ~n31988 ;
  assign \s13_addr_o[25]_pad  = ~n32011 ;
  assign \s13_addr_o[26]_pad  = ~n32034 ;
  assign \s13_addr_o[27]_pad  = ~n32057 ;
  assign \s13_addr_o[28]_pad  = ~n32080 ;
  assign \s13_addr_o[29]_pad  = ~n32103 ;
  assign \s13_addr_o[2]_pad  = ~n32126 ;
  assign \s13_addr_o[30]_pad  = ~n32149 ;
  assign \s13_addr_o[31]_pad  = ~n32172 ;
  assign \s13_addr_o[3]_pad  = ~n32195 ;
  assign \s13_addr_o[4]_pad  = ~n32218 ;
  assign \s13_addr_o[5]_pad  = ~n32241 ;
  assign \s13_addr_o[6]_pad  = ~n32264 ;
  assign \s13_addr_o[7]_pad  = ~n32287 ;
  assign \s13_addr_o[8]_pad  = ~n32310 ;
  assign \s13_addr_o[9]_pad  = ~n32333 ;
  assign \s13_data_o[0]_pad  = ~n32356 ;
  assign \s13_data_o[10]_pad  = ~n32379 ;
  assign \s13_data_o[11]_pad  = ~n32402 ;
  assign \s13_data_o[12]_pad  = ~n32425 ;
  assign \s13_data_o[13]_pad  = ~n32448 ;
  assign \s13_data_o[14]_pad  = ~n32471 ;
  assign \s13_data_o[15]_pad  = ~n32494 ;
  assign \s13_data_o[16]_pad  = ~n32517 ;
  assign \s13_data_o[17]_pad  = ~n32540 ;
  assign \s13_data_o[18]_pad  = ~n32563 ;
  assign \s13_data_o[19]_pad  = ~n32586 ;
  assign \s13_data_o[1]_pad  = ~n32609 ;
  assign \s13_data_o[20]_pad  = ~n32632 ;
  assign \s13_data_o[21]_pad  = ~n32655 ;
  assign \s13_data_o[22]_pad  = ~n32678 ;
  assign \s13_data_o[23]_pad  = ~n32701 ;
  assign \s13_data_o[24]_pad  = ~n32724 ;
  assign \s13_data_o[25]_pad  = ~n32747 ;
  assign \s13_data_o[26]_pad  = ~n32770 ;
  assign \s13_data_o[27]_pad  = ~n32793 ;
  assign \s13_data_o[28]_pad  = ~n32816 ;
  assign \s13_data_o[29]_pad  = ~n32839 ;
  assign \s13_data_o[2]_pad  = ~n32862 ;
  assign \s13_data_o[30]_pad  = ~n32885 ;
  assign \s13_data_o[31]_pad  = ~n32908 ;
  assign \s13_data_o[3]_pad  = ~n32931 ;
  assign \s13_data_o[4]_pad  = ~n32954 ;
  assign \s13_data_o[5]_pad  = ~n32977 ;
  assign \s13_data_o[6]_pad  = ~n33000 ;
  assign \s13_data_o[7]_pad  = ~n33023 ;
  assign \s13_data_o[8]_pad  = ~n33046 ;
  assign \s13_data_o[9]_pad  = ~n33069 ;
  assign \s13_sel_o[0]_pad  = ~n33092 ;
  assign \s13_sel_o[1]_pad  = ~n33115 ;
  assign \s13_sel_o[2]_pad  = ~n33138 ;
  assign \s13_sel_o[3]_pad  = ~n33161 ;
  assign \s13_stb_o_pad  = ~n33192 ;
  assign \s13_we_o_pad  = ~n33215 ;
  assign \s14_addr_o[0]_pad  = ~n33238 ;
  assign \s14_addr_o[10]_pad  = ~n33261 ;
  assign \s14_addr_o[11]_pad  = ~n33284 ;
  assign \s14_addr_o[12]_pad  = ~n33307 ;
  assign \s14_addr_o[13]_pad  = ~n33330 ;
  assign \s14_addr_o[14]_pad  = ~n33353 ;
  assign \s14_addr_o[15]_pad  = ~n33376 ;
  assign \s14_addr_o[16]_pad  = ~n33399 ;
  assign \s14_addr_o[17]_pad  = ~n33422 ;
  assign \s14_addr_o[18]_pad  = ~n33445 ;
  assign \s14_addr_o[19]_pad  = ~n33468 ;
  assign \s14_addr_o[1]_pad  = ~n33491 ;
  assign \s14_addr_o[20]_pad  = ~n33514 ;
  assign \s14_addr_o[21]_pad  = ~n33537 ;
  assign \s14_addr_o[22]_pad  = ~n33560 ;
  assign \s14_addr_o[23]_pad  = ~n33583 ;
  assign \s14_addr_o[24]_pad  = ~n33606 ;
  assign \s14_addr_o[25]_pad  = ~n33629 ;
  assign \s14_addr_o[26]_pad  = ~n33652 ;
  assign \s14_addr_o[27]_pad  = ~n33675 ;
  assign \s14_addr_o[28]_pad  = ~n33698 ;
  assign \s14_addr_o[29]_pad  = ~n33721 ;
  assign \s14_addr_o[2]_pad  = ~n33744 ;
  assign \s14_addr_o[30]_pad  = ~n33767 ;
  assign \s14_addr_o[31]_pad  = ~n33790 ;
  assign \s14_addr_o[3]_pad  = ~n33813 ;
  assign \s14_addr_o[4]_pad  = ~n33836 ;
  assign \s14_addr_o[5]_pad  = ~n33859 ;
  assign \s14_addr_o[6]_pad  = ~n33882 ;
  assign \s14_addr_o[7]_pad  = ~n33905 ;
  assign \s14_addr_o[8]_pad  = ~n33928 ;
  assign \s14_addr_o[9]_pad  = ~n33951 ;
  assign \s14_data_o[0]_pad  = ~n33974 ;
  assign \s14_data_o[10]_pad  = ~n33997 ;
  assign \s14_data_o[11]_pad  = ~n34020 ;
  assign \s14_data_o[12]_pad  = ~n34043 ;
  assign \s14_data_o[13]_pad  = ~n34066 ;
  assign \s14_data_o[14]_pad  = ~n34089 ;
  assign \s14_data_o[15]_pad  = ~n34112 ;
  assign \s14_data_o[16]_pad  = ~n34135 ;
  assign \s14_data_o[17]_pad  = ~n34158 ;
  assign \s14_data_o[18]_pad  = ~n34181 ;
  assign \s14_data_o[19]_pad  = ~n34204 ;
  assign \s14_data_o[1]_pad  = ~n34227 ;
  assign \s14_data_o[20]_pad  = ~n34250 ;
  assign \s14_data_o[21]_pad  = ~n34273 ;
  assign \s14_data_o[22]_pad  = ~n34296 ;
  assign \s14_data_o[23]_pad  = ~n34319 ;
  assign \s14_data_o[24]_pad  = ~n34342 ;
  assign \s14_data_o[25]_pad  = ~n34365 ;
  assign \s14_data_o[26]_pad  = ~n34388 ;
  assign \s14_data_o[27]_pad  = ~n34411 ;
  assign \s14_data_o[28]_pad  = ~n34434 ;
  assign \s14_data_o[29]_pad  = ~n34457 ;
  assign \s14_data_o[2]_pad  = ~n34480 ;
  assign \s14_data_o[30]_pad  = ~n34503 ;
  assign \s14_data_o[31]_pad  = ~n34526 ;
  assign \s14_data_o[3]_pad  = ~n34549 ;
  assign \s14_data_o[4]_pad  = ~n34572 ;
  assign \s14_data_o[5]_pad  = ~n34595 ;
  assign \s14_data_o[6]_pad  = ~n34618 ;
  assign \s14_data_o[7]_pad  = ~n34641 ;
  assign \s14_data_o[8]_pad  = ~n34664 ;
  assign \s14_data_o[9]_pad  = ~n34687 ;
  assign \s14_sel_o[0]_pad  = ~n34710 ;
  assign \s14_sel_o[1]_pad  = ~n34733 ;
  assign \s14_sel_o[2]_pad  = ~n34756 ;
  assign \s14_sel_o[3]_pad  = ~n34779 ;
  assign \s14_stb_o_pad  = ~n34810 ;
  assign \s14_we_o_pad  = ~n34833 ;
  assign \s15_addr_o[0]_pad  = ~n34856 ;
  assign \s15_addr_o[10]_pad  = ~n34879 ;
  assign \s15_addr_o[11]_pad  = ~n34902 ;
  assign \s15_addr_o[12]_pad  = ~n34925 ;
  assign \s15_addr_o[13]_pad  = ~n34948 ;
  assign \s15_addr_o[14]_pad  = ~n34971 ;
  assign \s15_addr_o[15]_pad  = ~n34994 ;
  assign \s15_addr_o[16]_pad  = ~n35017 ;
  assign \s15_addr_o[17]_pad  = ~n35040 ;
  assign \s15_addr_o[18]_pad  = ~n35063 ;
  assign \s15_addr_o[19]_pad  = ~n35086 ;
  assign \s15_addr_o[1]_pad  = ~n35109 ;
  assign \s15_addr_o[20]_pad  = ~n35132 ;
  assign \s15_addr_o[21]_pad  = ~n35155 ;
  assign \s15_addr_o[22]_pad  = ~n35178 ;
  assign \s15_addr_o[23]_pad  = ~n35201 ;
  assign \s15_addr_o[24]_pad  = ~n2152 ;
  assign \s15_addr_o[25]_pad  = ~n2232 ;
  assign \s15_addr_o[26]_pad  = ~n2255 ;
  assign \s15_addr_o[27]_pad  = ~n2129 ;
  assign \s15_addr_o[28]_pad  = ~n35224 ;
  assign \s15_addr_o[29]_pad  = ~n35247 ;
  assign \s15_addr_o[2]_pad  = ~n1951 ;
  assign \s15_addr_o[30]_pad  = ~n35270 ;
  assign \s15_addr_o[31]_pad  = ~n35293 ;
  assign \s15_addr_o[3]_pad  = ~n1974 ;
  assign \s15_addr_o[4]_pad  = ~n2021 ;
  assign \s15_addr_o[6]_pad  = ~n35316 ;
  assign \s15_addr_o[7]_pad  = ~n35339 ;
  assign \s15_addr_o[8]_pad  = ~n35362 ;
  assign \s15_addr_o[9]_pad  = ~n35385 ;
  assign \s15_cyc_o_pad  = n35386 ;
  assign \s15_data_o[0]_pad  = ~n12268 ;
  assign \s15_data_o[10]_pad  = ~n12296 ;
  assign \s15_data_o[11]_pad  = ~n12323 ;
  assign \s15_data_o[12]_pad  = ~n12350 ;
  assign \s15_data_o[13]_pad  = ~n12377 ;
  assign \s15_data_o[14]_pad  = ~n12404 ;
  assign \s15_data_o[15]_pad  = ~n12431 ;
  assign \s15_data_o[16]_pad  = ~n35409 ;
  assign \s15_data_o[17]_pad  = ~n35432 ;
  assign \s15_data_o[18]_pad  = ~n35455 ;
  assign \s15_data_o[19]_pad  = ~n35478 ;
  assign \s15_data_o[1]_pad  = ~n12458 ;
  assign \s15_data_o[20]_pad  = ~n35501 ;
  assign \s15_data_o[21]_pad  = ~n35524 ;
  assign \s15_data_o[22]_pad  = ~n35547 ;
  assign \s15_data_o[23]_pad  = ~n35570 ;
  assign \s15_data_o[24]_pad  = ~n35593 ;
  assign \s15_data_o[25]_pad  = ~n35616 ;
  assign \s15_data_o[26]_pad  = ~n35639 ;
  assign \s15_data_o[27]_pad  = ~n35662 ;
  assign \s15_data_o[28]_pad  = ~n35685 ;
  assign \s15_data_o[29]_pad  = ~n35708 ;
  assign \s15_data_o[2]_pad  = ~n12485 ;
  assign \s15_data_o[30]_pad  = ~n35731 ;
  assign \s15_data_o[31]_pad  = ~n35754 ;
  assign \s15_data_o[3]_pad  = ~n12512 ;
  assign \s15_data_o[4]_pad  = ~n12539 ;
  assign \s15_data_o[5]_pad  = ~n12566 ;
  assign \s15_data_o[6]_pad  = ~n12593 ;
  assign \s15_data_o[7]_pad  = ~n12620 ;
  assign \s15_data_o[8]_pad  = ~n12647 ;
  assign \s15_data_o[9]_pad  = ~n12674 ;
  assign \s15_sel_o[0]_pad  = ~n35777 ;
  assign \s15_sel_o[1]_pad  = ~n35800 ;
  assign \s15_sel_o[2]_pad  = ~n35823 ;
  assign \s15_sel_o[3]_pad  = ~n35846 ;
  assign \s15_stb_o_pad  = ~n2209 ;
  assign \s15_we_o_pad  = ~n13439 ;
  assign \s1_addr_o[0]_pad  = ~n35869 ;
  assign \s1_addr_o[10]_pad  = ~n35892 ;
  assign \s1_addr_o[11]_pad  = ~n35915 ;
  assign \s1_addr_o[12]_pad  = ~n35938 ;
  assign \s1_addr_o[13]_pad  = ~n35961 ;
  assign \s1_addr_o[14]_pad  = ~n35984 ;
  assign \s1_addr_o[15]_pad  = ~n36007 ;
  assign \s1_addr_o[16]_pad  = ~n36030 ;
  assign \s1_addr_o[17]_pad  = ~n36053 ;
  assign \s1_addr_o[18]_pad  = ~n36076 ;
  assign \s1_addr_o[19]_pad  = ~n36099 ;
  assign \s1_addr_o[1]_pad  = ~n36122 ;
  assign \s1_addr_o[20]_pad  = ~n36145 ;
  assign \s1_addr_o[21]_pad  = ~n36168 ;
  assign \s1_addr_o[22]_pad  = ~n36191 ;
  assign \s1_addr_o[23]_pad  = ~n36214 ;
  assign \s1_addr_o[24]_pad  = ~n36237 ;
  assign \s1_addr_o[25]_pad  = ~n36260 ;
  assign \s1_addr_o[26]_pad  = ~n36283 ;
  assign \s1_addr_o[27]_pad  = ~n36306 ;
  assign \s1_addr_o[28]_pad  = ~n36329 ;
  assign \s1_addr_o[29]_pad  = ~n36352 ;
  assign \s1_addr_o[2]_pad  = ~n36375 ;
  assign \s1_addr_o[30]_pad  = ~n36398 ;
  assign \s1_addr_o[31]_pad  = ~n36421 ;
  assign \s1_addr_o[3]_pad  = ~n36444 ;
  assign \s1_addr_o[4]_pad  = ~n36467 ;
  assign \s1_addr_o[5]_pad  = ~n36490 ;
  assign \s1_addr_o[6]_pad  = ~n36513 ;
  assign \s1_addr_o[7]_pad  = ~n36536 ;
  assign \s1_addr_o[8]_pad  = ~n36559 ;
  assign \s1_addr_o[9]_pad  = ~n36582 ;
  assign \s1_data_o[0]_pad  = ~n36605 ;
  assign \s1_data_o[10]_pad  = ~n36628 ;
  assign \s1_data_o[11]_pad  = ~n36651 ;
  assign \s1_data_o[12]_pad  = ~n36674 ;
  assign \s1_data_o[13]_pad  = ~n36697 ;
  assign \s1_data_o[14]_pad  = ~n36720 ;
  assign \s1_data_o[15]_pad  = ~n36743 ;
  assign \s1_data_o[16]_pad  = ~n36766 ;
  assign \s1_data_o[17]_pad  = ~n36789 ;
  assign \s1_data_o[18]_pad  = ~n36812 ;
  assign \s1_data_o[19]_pad  = ~n36835 ;
  assign \s1_data_o[1]_pad  = ~n36858 ;
  assign \s1_data_o[20]_pad  = ~n36881 ;
  assign \s1_data_o[21]_pad  = ~n36904 ;
  assign \s1_data_o[22]_pad  = ~n36927 ;
  assign \s1_data_o[23]_pad  = ~n36950 ;
  assign \s1_data_o[24]_pad  = ~n36973 ;
  assign \s1_data_o[25]_pad  = ~n36996 ;
  assign \s1_data_o[26]_pad  = ~n37019 ;
  assign \s1_data_o[27]_pad  = ~n37042 ;
  assign \s1_data_o[28]_pad  = ~n37065 ;
  assign \s1_data_o[29]_pad  = ~n37088 ;
  assign \s1_data_o[2]_pad  = ~n37111 ;
  assign \s1_data_o[30]_pad  = ~n37134 ;
  assign \s1_data_o[31]_pad  = ~n37157 ;
  assign \s1_data_o[3]_pad  = ~n37180 ;
  assign \s1_data_o[4]_pad  = ~n37203 ;
  assign \s1_data_o[5]_pad  = ~n37226 ;
  assign \s1_data_o[6]_pad  = ~n37249 ;
  assign \s1_data_o[7]_pad  = ~n37272 ;
  assign \s1_data_o[8]_pad  = ~n37295 ;
  assign \s1_data_o[9]_pad  = ~n37318 ;
  assign \s1_sel_o[0]_pad  = ~n37341 ;
  assign \s1_sel_o[1]_pad  = ~n37364 ;
  assign \s1_sel_o[2]_pad  = ~n37387 ;
  assign \s1_sel_o[3]_pad  = ~n37410 ;
  assign \s1_stb_o_pad  = ~n37441 ;
  assign \s1_we_o_pad  = ~n37464 ;
  assign \s2_addr_o[0]_pad  = ~n37487 ;
  assign \s2_addr_o[10]_pad  = ~n37510 ;
  assign \s2_addr_o[11]_pad  = ~n37533 ;
  assign \s2_addr_o[12]_pad  = ~n37556 ;
  assign \s2_addr_o[13]_pad  = ~n37579 ;
  assign \s2_addr_o[14]_pad  = ~n37602 ;
  assign \s2_addr_o[15]_pad  = ~n37625 ;
  assign \s2_addr_o[16]_pad  = ~n37648 ;
  assign \s2_addr_o[17]_pad  = ~n37671 ;
  assign \s2_addr_o[18]_pad  = ~n37694 ;
  assign \s2_addr_o[19]_pad  = ~n37717 ;
  assign \s2_addr_o[1]_pad  = ~n37740 ;
  assign \s2_addr_o[20]_pad  = ~n37763 ;
  assign \s2_addr_o[21]_pad  = ~n37786 ;
  assign \s2_addr_o[22]_pad  = ~n37809 ;
  assign \s2_addr_o[23]_pad  = ~n37832 ;
  assign \s2_addr_o[24]_pad  = ~n37855 ;
  assign \s2_addr_o[25]_pad  = ~n37878 ;
  assign \s2_addr_o[26]_pad  = ~n37901 ;
  assign \s2_addr_o[27]_pad  = ~n37924 ;
  assign \s2_addr_o[28]_pad  = ~n37947 ;
  assign \s2_addr_o[29]_pad  = ~n37970 ;
  assign \s2_addr_o[2]_pad  = ~n37993 ;
  assign \s2_addr_o[30]_pad  = ~n38016 ;
  assign \s2_addr_o[31]_pad  = ~n38039 ;
  assign \s2_addr_o[3]_pad  = ~n38062 ;
  assign \s2_addr_o[4]_pad  = ~n38085 ;
  assign \s2_addr_o[5]_pad  = ~n38108 ;
  assign \s2_addr_o[6]_pad  = ~n38131 ;
  assign \s2_addr_o[7]_pad  = ~n38154 ;
  assign \s2_addr_o[8]_pad  = ~n38177 ;
  assign \s2_addr_o[9]_pad  = ~n38200 ;
  assign \s2_data_o[0]_pad  = ~n38223 ;
  assign \s2_data_o[10]_pad  = ~n38246 ;
  assign \s2_data_o[11]_pad  = ~n38269 ;
  assign \s2_data_o[12]_pad  = ~n38292 ;
  assign \s2_data_o[13]_pad  = ~n38315 ;
  assign \s2_data_o[14]_pad  = ~n38338 ;
  assign \s2_data_o[15]_pad  = ~n38361 ;
  assign \s2_data_o[16]_pad  = ~n38384 ;
  assign \s2_data_o[17]_pad  = ~n38407 ;
  assign \s2_data_o[18]_pad  = ~n38430 ;
  assign \s2_data_o[19]_pad  = ~n38453 ;
  assign \s2_data_o[1]_pad  = ~n38476 ;
  assign \s2_data_o[20]_pad  = ~n38499 ;
  assign \s2_data_o[21]_pad  = ~n38522 ;
  assign \s2_data_o[22]_pad  = ~n38545 ;
  assign \s2_data_o[23]_pad  = ~n38568 ;
  assign \s2_data_o[24]_pad  = ~n38591 ;
  assign \s2_data_o[25]_pad  = ~n38614 ;
  assign \s2_data_o[26]_pad  = ~n38637 ;
  assign \s2_data_o[27]_pad  = ~n38660 ;
  assign \s2_data_o[28]_pad  = ~n38683 ;
  assign \s2_data_o[29]_pad  = ~n38706 ;
  assign \s2_data_o[2]_pad  = ~n38729 ;
  assign \s2_data_o[30]_pad  = ~n38752 ;
  assign \s2_data_o[31]_pad  = ~n38775 ;
  assign \s2_data_o[3]_pad  = ~n38798 ;
  assign \s2_data_o[4]_pad  = ~n38821 ;
  assign \s2_data_o[5]_pad  = ~n38844 ;
  assign \s2_data_o[6]_pad  = ~n38867 ;
  assign \s2_data_o[7]_pad  = ~n38890 ;
  assign \s2_data_o[8]_pad  = ~n38913 ;
  assign \s2_data_o[9]_pad  = ~n38936 ;
  assign \s2_sel_o[0]_pad  = ~n38959 ;
  assign \s2_sel_o[1]_pad  = ~n38982 ;
  assign \s2_sel_o[2]_pad  = ~n39005 ;
  assign \s2_sel_o[3]_pad  = ~n39028 ;
  assign \s2_stb_o_pad  = ~n39059 ;
  assign \s2_we_o_pad  = ~n39082 ;
  assign \s3_addr_o[0]_pad  = ~n39105 ;
  assign \s3_addr_o[10]_pad  = ~n39128 ;
  assign \s3_addr_o[11]_pad  = ~n39151 ;
  assign \s3_addr_o[12]_pad  = ~n39174 ;
  assign \s3_addr_o[13]_pad  = ~n39197 ;
  assign \s3_addr_o[14]_pad  = ~n39220 ;
  assign \s3_addr_o[15]_pad  = ~n39243 ;
  assign \s3_addr_o[16]_pad  = ~n39266 ;
  assign \s3_addr_o[17]_pad  = ~n39289 ;
  assign \s3_addr_o[18]_pad  = ~n39312 ;
  assign \s3_addr_o[19]_pad  = ~n39335 ;
  assign \s3_addr_o[1]_pad  = ~n39358 ;
  assign \s3_addr_o[20]_pad  = ~n39381 ;
  assign \s3_addr_o[21]_pad  = ~n39404 ;
  assign \s3_addr_o[22]_pad  = ~n39427 ;
  assign \s3_addr_o[23]_pad  = ~n39450 ;
  assign \s3_addr_o[24]_pad  = ~n39473 ;
  assign \s3_addr_o[25]_pad  = ~n39496 ;
  assign \s3_addr_o[26]_pad  = ~n39519 ;
  assign \s3_addr_o[27]_pad  = ~n39542 ;
  assign \s3_addr_o[28]_pad  = ~n39565 ;
  assign \s3_addr_o[29]_pad  = ~n39588 ;
  assign \s3_addr_o[2]_pad  = ~n39611 ;
  assign \s3_addr_o[30]_pad  = ~n39634 ;
  assign \s3_addr_o[31]_pad  = ~n39657 ;
  assign \s3_addr_o[3]_pad  = ~n39680 ;
  assign \s3_addr_o[4]_pad  = ~n39703 ;
  assign \s3_addr_o[5]_pad  = ~n39726 ;
  assign \s3_addr_o[6]_pad  = ~n39749 ;
  assign \s3_addr_o[7]_pad  = ~n39772 ;
  assign \s3_addr_o[8]_pad  = ~n39795 ;
  assign \s3_addr_o[9]_pad  = ~n39818 ;
  assign \s3_data_o[0]_pad  = ~n39841 ;
  assign \s3_data_o[10]_pad  = ~n39864 ;
  assign \s3_data_o[11]_pad  = ~n39887 ;
  assign \s3_data_o[12]_pad  = ~n39910 ;
  assign \s3_data_o[13]_pad  = ~n39933 ;
  assign \s3_data_o[14]_pad  = ~n39956 ;
  assign \s3_data_o[15]_pad  = ~n39979 ;
  assign \s3_data_o[16]_pad  = ~n40002 ;
  assign \s3_data_o[17]_pad  = ~n40025 ;
  assign \s3_data_o[18]_pad  = ~n40048 ;
  assign \s3_data_o[19]_pad  = ~n40071 ;
  assign \s3_data_o[1]_pad  = ~n40094 ;
  assign \s3_data_o[20]_pad  = ~n40117 ;
  assign \s3_data_o[21]_pad  = ~n40140 ;
  assign \s3_data_o[22]_pad  = ~n40163 ;
  assign \s3_data_o[23]_pad  = ~n40186 ;
  assign \s3_data_o[24]_pad  = ~n40209 ;
  assign \s3_data_o[25]_pad  = ~n40232 ;
  assign \s3_data_o[26]_pad  = ~n40255 ;
  assign \s3_data_o[27]_pad  = ~n40278 ;
  assign \s3_data_o[28]_pad  = ~n40301 ;
  assign \s3_data_o[29]_pad  = ~n40324 ;
  assign \s3_data_o[2]_pad  = ~n40347 ;
  assign \s3_data_o[30]_pad  = ~n40370 ;
  assign \s3_data_o[31]_pad  = ~n40393 ;
  assign \s3_data_o[3]_pad  = ~n40416 ;
  assign \s3_data_o[4]_pad  = ~n40439 ;
  assign \s3_data_o[5]_pad  = ~n40462 ;
  assign \s3_data_o[6]_pad  = ~n40485 ;
  assign \s3_data_o[7]_pad  = ~n40508 ;
  assign \s3_data_o[8]_pad  = ~n40531 ;
  assign \s3_data_o[9]_pad  = ~n40554 ;
  assign \s3_sel_o[0]_pad  = ~n40577 ;
  assign \s3_sel_o[1]_pad  = ~n40600 ;
  assign \s3_sel_o[2]_pad  = ~n40623 ;
  assign \s3_sel_o[3]_pad  = ~n40646 ;
  assign \s3_stb_o_pad  = ~n40677 ;
  assign \s3_we_o_pad  = ~n40700 ;
  assign \s4_addr_o[0]_pad  = ~n40723 ;
  assign \s4_addr_o[10]_pad  = ~n40746 ;
  assign \s4_addr_o[11]_pad  = ~n40769 ;
  assign \s4_addr_o[12]_pad  = ~n40792 ;
  assign \s4_addr_o[13]_pad  = ~n40815 ;
  assign \s4_addr_o[14]_pad  = ~n40838 ;
  assign \s4_addr_o[15]_pad  = ~n40861 ;
  assign \s4_addr_o[16]_pad  = ~n40884 ;
  assign \s4_addr_o[17]_pad  = ~n40907 ;
  assign \s4_addr_o[18]_pad  = ~n40930 ;
  assign \s4_addr_o[19]_pad  = ~n40953 ;
  assign \s4_addr_o[1]_pad  = ~n40976 ;
  assign \s4_addr_o[20]_pad  = ~n40999 ;
  assign \s4_addr_o[21]_pad  = ~n41022 ;
  assign \s4_addr_o[22]_pad  = ~n41045 ;
  assign \s4_addr_o[23]_pad  = ~n41068 ;
  assign \s4_addr_o[24]_pad  = ~n41091 ;
  assign \s4_addr_o[25]_pad  = ~n41114 ;
  assign \s4_addr_o[26]_pad  = ~n41137 ;
  assign \s4_addr_o[27]_pad  = ~n41160 ;
  assign \s4_addr_o[28]_pad  = ~n41183 ;
  assign \s4_addr_o[29]_pad  = ~n41206 ;
  assign \s4_addr_o[2]_pad  = ~n41229 ;
  assign \s4_addr_o[30]_pad  = ~n41252 ;
  assign \s4_addr_o[31]_pad  = ~n41275 ;
  assign \s4_addr_o[3]_pad  = ~n41298 ;
  assign \s4_addr_o[4]_pad  = ~n41321 ;
  assign \s4_addr_o[5]_pad  = ~n41344 ;
  assign \s4_addr_o[6]_pad  = ~n41367 ;
  assign \s4_addr_o[7]_pad  = ~n41390 ;
  assign \s4_addr_o[8]_pad  = ~n41413 ;
  assign \s4_addr_o[9]_pad  = ~n41436 ;
  assign \s4_data_o[0]_pad  = ~n41459 ;
  assign \s4_data_o[10]_pad  = ~n41482 ;
  assign \s4_data_o[11]_pad  = ~n41505 ;
  assign \s4_data_o[12]_pad  = ~n41528 ;
  assign \s4_data_o[13]_pad  = ~n41551 ;
  assign \s4_data_o[14]_pad  = ~n41574 ;
  assign \s4_data_o[15]_pad  = ~n41597 ;
  assign \s4_data_o[16]_pad  = ~n41620 ;
  assign \s4_data_o[17]_pad  = ~n41643 ;
  assign \s4_data_o[18]_pad  = ~n41666 ;
  assign \s4_data_o[19]_pad  = ~n41689 ;
  assign \s4_data_o[1]_pad  = ~n41712 ;
  assign \s4_data_o[20]_pad  = ~n41735 ;
  assign \s4_data_o[21]_pad  = ~n41758 ;
  assign \s4_data_o[22]_pad  = ~n41781 ;
  assign \s4_data_o[23]_pad  = ~n41804 ;
  assign \s4_data_o[24]_pad  = ~n41827 ;
  assign \s4_data_o[25]_pad  = ~n41850 ;
  assign \s4_data_o[26]_pad  = ~n41873 ;
  assign \s4_data_o[27]_pad  = ~n41896 ;
  assign \s4_data_o[28]_pad  = ~n41919 ;
  assign \s4_data_o[29]_pad  = ~n41942 ;
  assign \s4_data_o[2]_pad  = ~n41965 ;
  assign \s4_data_o[30]_pad  = ~n41988 ;
  assign \s4_data_o[31]_pad  = ~n42011 ;
  assign \s4_data_o[3]_pad  = ~n42034 ;
  assign \s4_data_o[4]_pad  = ~n42057 ;
  assign \s4_data_o[5]_pad  = ~n42080 ;
  assign \s4_data_o[6]_pad  = ~n42103 ;
  assign \s4_data_o[7]_pad  = ~n42126 ;
  assign \s4_data_o[8]_pad  = ~n42149 ;
  assign \s4_data_o[9]_pad  = ~n42172 ;
  assign \s4_sel_o[0]_pad  = ~n42195 ;
  assign \s4_sel_o[1]_pad  = ~n42218 ;
  assign \s4_sel_o[2]_pad  = ~n42241 ;
  assign \s4_sel_o[3]_pad  = ~n42264 ;
  assign \s4_stb_o_pad  = ~n42295 ;
  assign \s4_we_o_pad  = ~n42318 ;
  assign \s5_addr_o[0]_pad  = ~n42341 ;
  assign \s5_addr_o[10]_pad  = ~n42364 ;
  assign \s5_addr_o[11]_pad  = ~n42387 ;
  assign \s5_addr_o[12]_pad  = ~n42410 ;
  assign \s5_addr_o[13]_pad  = ~n42433 ;
  assign \s5_addr_o[14]_pad  = ~n42456 ;
  assign \s5_addr_o[15]_pad  = ~n42479 ;
  assign \s5_addr_o[16]_pad  = ~n42502 ;
  assign \s5_addr_o[17]_pad  = ~n42525 ;
  assign \s5_addr_o[18]_pad  = ~n42548 ;
  assign \s5_addr_o[19]_pad  = ~n42571 ;
  assign \s5_addr_o[1]_pad  = ~n42594 ;
  assign \s5_addr_o[20]_pad  = ~n42617 ;
  assign \s5_addr_o[21]_pad  = ~n42640 ;
  assign \s5_addr_o[22]_pad  = ~n42663 ;
  assign \s5_addr_o[23]_pad  = ~n42686 ;
  assign \s5_addr_o[24]_pad  = ~n42709 ;
  assign \s5_addr_o[25]_pad  = ~n42732 ;
  assign \s5_addr_o[26]_pad  = ~n42755 ;
  assign \s5_addr_o[27]_pad  = ~n42778 ;
  assign \s5_addr_o[28]_pad  = ~n42801 ;
  assign \s5_addr_o[29]_pad  = ~n42824 ;
  assign \s5_addr_o[2]_pad  = ~n42847 ;
  assign \s5_addr_o[30]_pad  = ~n42870 ;
  assign \s5_addr_o[31]_pad  = ~n42893 ;
  assign \s5_addr_o[3]_pad  = ~n42916 ;
  assign \s5_addr_o[4]_pad  = ~n42939 ;
  assign \s5_addr_o[5]_pad  = ~n42962 ;
  assign \s5_addr_o[6]_pad  = ~n42985 ;
  assign \s5_addr_o[7]_pad  = ~n43008 ;
  assign \s5_addr_o[8]_pad  = ~n43031 ;
  assign \s5_addr_o[9]_pad  = ~n43054 ;
  assign \s5_data_o[0]_pad  = ~n43077 ;
  assign \s5_data_o[10]_pad  = ~n43100 ;
  assign \s5_data_o[11]_pad  = ~n43123 ;
  assign \s5_data_o[12]_pad  = ~n43146 ;
  assign \s5_data_o[13]_pad  = ~n43169 ;
  assign \s5_data_o[14]_pad  = ~n43192 ;
  assign \s5_data_o[15]_pad  = ~n43215 ;
  assign \s5_data_o[16]_pad  = ~n43238 ;
  assign \s5_data_o[17]_pad  = ~n43261 ;
  assign \s5_data_o[18]_pad  = ~n43284 ;
  assign \s5_data_o[19]_pad  = ~n43307 ;
  assign \s5_data_o[1]_pad  = ~n43330 ;
  assign \s5_data_o[20]_pad  = ~n43353 ;
  assign \s5_data_o[21]_pad  = ~n43376 ;
  assign \s5_data_o[22]_pad  = ~n43399 ;
  assign \s5_data_o[23]_pad  = ~n43422 ;
  assign \s5_data_o[24]_pad  = ~n43445 ;
  assign \s5_data_o[25]_pad  = ~n43468 ;
  assign \s5_data_o[26]_pad  = ~n43491 ;
  assign \s5_data_o[27]_pad  = ~n43514 ;
  assign \s5_data_o[28]_pad  = ~n43537 ;
  assign \s5_data_o[29]_pad  = ~n43560 ;
  assign \s5_data_o[2]_pad  = ~n43583 ;
  assign \s5_data_o[30]_pad  = ~n43606 ;
  assign \s5_data_o[31]_pad  = ~n43629 ;
  assign \s5_data_o[3]_pad  = ~n43652 ;
  assign \s5_data_o[4]_pad  = ~n43675 ;
  assign \s5_data_o[5]_pad  = ~n43698 ;
  assign \s5_data_o[6]_pad  = ~n43721 ;
  assign \s5_data_o[7]_pad  = ~n43744 ;
  assign \s5_data_o[8]_pad  = ~n43767 ;
  assign \s5_data_o[9]_pad  = ~n43790 ;
  assign \s5_sel_o[0]_pad  = ~n43813 ;
  assign \s5_sel_o[1]_pad  = ~n43836 ;
  assign \s5_sel_o[2]_pad  = ~n43859 ;
  assign \s5_sel_o[3]_pad  = ~n43882 ;
  assign \s5_stb_o_pad  = ~n43913 ;
  assign \s5_we_o_pad  = ~n43936 ;
  assign \s6_addr_o[0]_pad  = ~n43959 ;
  assign \s6_addr_o[10]_pad  = ~n43982 ;
  assign \s6_addr_o[11]_pad  = ~n44005 ;
  assign \s6_addr_o[12]_pad  = ~n44028 ;
  assign \s6_addr_o[13]_pad  = ~n44051 ;
  assign \s6_addr_o[14]_pad  = ~n44074 ;
  assign \s6_addr_o[15]_pad  = ~n44097 ;
  assign \s6_addr_o[16]_pad  = ~n44120 ;
  assign \s6_addr_o[17]_pad  = ~n44143 ;
  assign \s6_addr_o[18]_pad  = ~n44166 ;
  assign \s6_addr_o[19]_pad  = ~n44189 ;
  assign \s6_addr_o[1]_pad  = ~n44212 ;
  assign \s6_addr_o[20]_pad  = ~n44235 ;
  assign \s6_addr_o[21]_pad  = ~n44258 ;
  assign \s6_addr_o[22]_pad  = ~n44281 ;
  assign \s6_addr_o[23]_pad  = ~n44304 ;
  assign \s6_addr_o[24]_pad  = ~n44327 ;
  assign \s6_addr_o[25]_pad  = ~n44350 ;
  assign \s6_addr_o[26]_pad  = ~n44373 ;
  assign \s6_addr_o[27]_pad  = ~n44396 ;
  assign \s6_addr_o[28]_pad  = ~n44419 ;
  assign \s6_addr_o[29]_pad  = ~n44442 ;
  assign \s6_addr_o[2]_pad  = ~n44465 ;
  assign \s6_addr_o[30]_pad  = ~n44488 ;
  assign \s6_addr_o[31]_pad  = ~n44511 ;
  assign \s6_addr_o[3]_pad  = ~n44534 ;
  assign \s6_addr_o[4]_pad  = ~n44557 ;
  assign \s6_addr_o[5]_pad  = ~n44580 ;
  assign \s6_addr_o[6]_pad  = ~n44603 ;
  assign \s6_addr_o[7]_pad  = ~n44626 ;
  assign \s6_addr_o[8]_pad  = ~n44649 ;
  assign \s6_addr_o[9]_pad  = ~n44672 ;
  assign \s6_data_o[0]_pad  = ~n44695 ;
  assign \s6_data_o[10]_pad  = ~n44718 ;
  assign \s6_data_o[11]_pad  = ~n44741 ;
  assign \s6_data_o[12]_pad  = ~n44764 ;
  assign \s6_data_o[13]_pad  = ~n44787 ;
  assign \s6_data_o[14]_pad  = ~n44810 ;
  assign \s6_data_o[15]_pad  = ~n44833 ;
  assign \s6_data_o[16]_pad  = ~n44856 ;
  assign \s6_data_o[17]_pad  = ~n44879 ;
  assign \s6_data_o[18]_pad  = ~n44902 ;
  assign \s6_data_o[19]_pad  = ~n44925 ;
  assign \s6_data_o[1]_pad  = ~n44948 ;
  assign \s6_data_o[20]_pad  = ~n44971 ;
  assign \s6_data_o[21]_pad  = ~n44994 ;
  assign \s6_data_o[22]_pad  = ~n45017 ;
  assign \s6_data_o[23]_pad  = ~n45040 ;
  assign \s6_data_o[24]_pad  = ~n45063 ;
  assign \s6_data_o[25]_pad  = ~n45086 ;
  assign \s6_data_o[26]_pad  = ~n45109 ;
  assign \s6_data_o[27]_pad  = ~n45132 ;
  assign \s6_data_o[28]_pad  = ~n45155 ;
  assign \s6_data_o[29]_pad  = ~n45178 ;
  assign \s6_data_o[2]_pad  = ~n45201 ;
  assign \s6_data_o[30]_pad  = ~n45224 ;
  assign \s6_data_o[31]_pad  = ~n45247 ;
  assign \s6_data_o[3]_pad  = ~n45270 ;
  assign \s6_data_o[4]_pad  = ~n45293 ;
  assign \s6_data_o[5]_pad  = ~n45316 ;
  assign \s6_data_o[6]_pad  = ~n45339 ;
  assign \s6_data_o[7]_pad  = ~n45362 ;
  assign \s6_data_o[8]_pad  = ~n45385 ;
  assign \s6_data_o[9]_pad  = ~n45408 ;
  assign \s6_sel_o[0]_pad  = ~n45431 ;
  assign \s6_sel_o[1]_pad  = ~n45454 ;
  assign \s6_sel_o[2]_pad  = ~n45477 ;
  assign \s6_sel_o[3]_pad  = ~n45500 ;
  assign \s6_stb_o_pad  = ~n45531 ;
  assign \s6_we_o_pad  = ~n45554 ;
  assign \s7_addr_o[0]_pad  = ~n45577 ;
  assign \s7_addr_o[10]_pad  = ~n45600 ;
  assign \s7_addr_o[11]_pad  = ~n45623 ;
  assign \s7_addr_o[12]_pad  = ~n45646 ;
  assign \s7_addr_o[13]_pad  = ~n45669 ;
  assign \s7_addr_o[14]_pad  = ~n45692 ;
  assign \s7_addr_o[15]_pad  = ~n45715 ;
  assign \s7_addr_o[16]_pad  = ~n45738 ;
  assign \s7_addr_o[17]_pad  = ~n45761 ;
  assign \s7_addr_o[18]_pad  = ~n45784 ;
  assign \s7_addr_o[19]_pad  = ~n45807 ;
  assign \s7_addr_o[1]_pad  = ~n45830 ;
  assign \s7_addr_o[20]_pad  = ~n45853 ;
  assign \s7_addr_o[21]_pad  = ~n45876 ;
  assign \s7_addr_o[22]_pad  = ~n45899 ;
  assign \s7_addr_o[23]_pad  = ~n45922 ;
  assign \s7_addr_o[24]_pad  = ~n45945 ;
  assign \s7_addr_o[25]_pad  = ~n45968 ;
  assign \s7_addr_o[26]_pad  = ~n45991 ;
  assign \s7_addr_o[27]_pad  = ~n46014 ;
  assign \s7_addr_o[28]_pad  = ~n46037 ;
  assign \s7_addr_o[29]_pad  = ~n46060 ;
  assign \s7_addr_o[2]_pad  = ~n46083 ;
  assign \s7_addr_o[30]_pad  = ~n46106 ;
  assign \s7_addr_o[31]_pad  = ~n46129 ;
  assign \s7_addr_o[3]_pad  = ~n46152 ;
  assign \s7_addr_o[4]_pad  = ~n46175 ;
  assign \s7_addr_o[5]_pad  = ~n46198 ;
  assign \s7_addr_o[6]_pad  = ~n46221 ;
  assign \s7_addr_o[7]_pad  = ~n46244 ;
  assign \s7_addr_o[8]_pad  = ~n46267 ;
  assign \s7_addr_o[9]_pad  = ~n46290 ;
  assign \s7_data_o[0]_pad  = ~n46313 ;
  assign \s7_data_o[10]_pad  = ~n46336 ;
  assign \s7_data_o[11]_pad  = ~n46359 ;
  assign \s7_data_o[12]_pad  = ~n46382 ;
  assign \s7_data_o[13]_pad  = ~n46405 ;
  assign \s7_data_o[14]_pad  = ~n46428 ;
  assign \s7_data_o[15]_pad  = ~n46451 ;
  assign \s7_data_o[16]_pad  = ~n46474 ;
  assign \s7_data_o[17]_pad  = ~n46497 ;
  assign \s7_data_o[18]_pad  = ~n46520 ;
  assign \s7_data_o[19]_pad  = ~n46543 ;
  assign \s7_data_o[1]_pad  = ~n46566 ;
  assign \s7_data_o[20]_pad  = ~n46589 ;
  assign \s7_data_o[21]_pad  = ~n46612 ;
  assign \s7_data_o[22]_pad  = ~n46635 ;
  assign \s7_data_o[23]_pad  = ~n46658 ;
  assign \s7_data_o[24]_pad  = ~n46681 ;
  assign \s7_data_o[25]_pad  = ~n46704 ;
  assign \s7_data_o[26]_pad  = ~n46727 ;
  assign \s7_data_o[27]_pad  = ~n46750 ;
  assign \s7_data_o[28]_pad  = ~n46773 ;
  assign \s7_data_o[29]_pad  = ~n46796 ;
  assign \s7_data_o[2]_pad  = ~n46819 ;
  assign \s7_data_o[30]_pad  = ~n46842 ;
  assign \s7_data_o[31]_pad  = ~n46865 ;
  assign \s7_data_o[3]_pad  = ~n46888 ;
  assign \s7_data_o[4]_pad  = ~n46911 ;
  assign \s7_data_o[5]_pad  = ~n46934 ;
  assign \s7_data_o[6]_pad  = ~n46957 ;
  assign \s7_data_o[7]_pad  = ~n46980 ;
  assign \s7_data_o[8]_pad  = ~n47003 ;
  assign \s7_data_o[9]_pad  = ~n47026 ;
  assign \s7_sel_o[0]_pad  = ~n47049 ;
  assign \s7_sel_o[1]_pad  = ~n47072 ;
  assign \s7_sel_o[2]_pad  = ~n47095 ;
  assign \s7_sel_o[3]_pad  = ~n47118 ;
  assign \s7_stb_o_pad  = ~n47149 ;
  assign \s7_we_o_pad  = ~n47172 ;
  assign \s8_addr_o[0]_pad  = ~n47195 ;
  assign \s8_addr_o[10]_pad  = ~n47218 ;
  assign \s8_addr_o[11]_pad  = ~n47241 ;
  assign \s8_addr_o[12]_pad  = ~n47264 ;
  assign \s8_addr_o[13]_pad  = ~n47287 ;
  assign \s8_addr_o[14]_pad  = ~n47310 ;
  assign \s8_addr_o[15]_pad  = ~n47333 ;
  assign \s8_addr_o[16]_pad  = ~n47356 ;
  assign \s8_addr_o[17]_pad  = ~n47379 ;
  assign \s8_addr_o[18]_pad  = ~n47402 ;
  assign \s8_addr_o[19]_pad  = ~n47425 ;
  assign \s8_addr_o[1]_pad  = ~n47448 ;
  assign \s8_addr_o[20]_pad  = ~n47471 ;
  assign \s8_addr_o[21]_pad  = ~n47494 ;
  assign \s8_addr_o[22]_pad  = ~n47517 ;
  assign \s8_addr_o[23]_pad  = ~n47540 ;
  assign \s8_addr_o[24]_pad  = ~n47563 ;
  assign \s8_addr_o[25]_pad  = ~n47586 ;
  assign \s8_addr_o[26]_pad  = ~n47609 ;
  assign \s8_addr_o[27]_pad  = ~n47632 ;
  assign \s8_addr_o[28]_pad  = ~n47655 ;
  assign \s8_addr_o[29]_pad  = ~n47678 ;
  assign \s8_addr_o[2]_pad  = ~n47701 ;
  assign \s8_addr_o[30]_pad  = ~n47724 ;
  assign \s8_addr_o[31]_pad  = ~n47747 ;
  assign \s8_addr_o[3]_pad  = ~n47770 ;
  assign \s8_addr_o[4]_pad  = ~n47793 ;
  assign \s8_addr_o[5]_pad  = ~n47816 ;
  assign \s8_addr_o[6]_pad  = ~n47839 ;
  assign \s8_addr_o[7]_pad  = ~n47862 ;
  assign \s8_addr_o[8]_pad  = ~n47885 ;
  assign \s8_addr_o[9]_pad  = ~n47908 ;
  assign \s8_data_o[0]_pad  = ~n47931 ;
  assign \s8_data_o[10]_pad  = ~n47954 ;
  assign \s8_data_o[11]_pad  = ~n47977 ;
  assign \s8_data_o[12]_pad  = ~n48000 ;
  assign \s8_data_o[13]_pad  = ~n48023 ;
  assign \s8_data_o[14]_pad  = ~n48046 ;
  assign \s8_data_o[15]_pad  = ~n48069 ;
  assign \s8_data_o[16]_pad  = ~n48092 ;
  assign \s8_data_o[17]_pad  = ~n48115 ;
  assign \s8_data_o[18]_pad  = ~n48138 ;
  assign \s8_data_o[19]_pad  = ~n48161 ;
  assign \s8_data_o[1]_pad  = ~n48184 ;
  assign \s8_data_o[20]_pad  = ~n48207 ;
  assign \s8_data_o[21]_pad  = ~n48230 ;
  assign \s8_data_o[22]_pad  = ~n48253 ;
  assign \s8_data_o[23]_pad  = ~n48276 ;
  assign \s8_data_o[24]_pad  = ~n48299 ;
  assign \s8_data_o[25]_pad  = ~n48322 ;
  assign \s8_data_o[26]_pad  = ~n48345 ;
  assign \s8_data_o[27]_pad  = ~n48368 ;
  assign \s8_data_o[28]_pad  = ~n48391 ;
  assign \s8_data_o[29]_pad  = ~n48414 ;
  assign \s8_data_o[2]_pad  = ~n48437 ;
  assign \s8_data_o[30]_pad  = ~n48460 ;
  assign \s8_data_o[31]_pad  = ~n48483 ;
  assign \s8_data_o[3]_pad  = ~n48506 ;
  assign \s8_data_o[4]_pad  = ~n48529 ;
  assign \s8_data_o[5]_pad  = ~n48552 ;
  assign \s8_data_o[6]_pad  = ~n48575 ;
  assign \s8_data_o[7]_pad  = ~n48598 ;
  assign \s8_data_o[8]_pad  = ~n48621 ;
  assign \s8_data_o[9]_pad  = ~n48644 ;
  assign \s8_sel_o[0]_pad  = ~n48667 ;
  assign \s8_sel_o[1]_pad  = ~n48690 ;
  assign \s8_sel_o[2]_pad  = ~n48713 ;
  assign \s8_sel_o[3]_pad  = ~n48736 ;
  assign \s8_stb_o_pad  = ~n48767 ;
  assign \s8_we_o_pad  = ~n48790 ;
  assign \s9_addr_o[0]_pad  = ~n48813 ;
  assign \s9_addr_o[10]_pad  = ~n48836 ;
  assign \s9_addr_o[11]_pad  = ~n48859 ;
  assign \s9_addr_o[12]_pad  = ~n48882 ;
  assign \s9_addr_o[13]_pad  = ~n48905 ;
  assign \s9_addr_o[14]_pad  = ~n48928 ;
  assign \s9_addr_o[15]_pad  = ~n48951 ;
  assign \s9_addr_o[16]_pad  = ~n48974 ;
  assign \s9_addr_o[17]_pad  = ~n48997 ;
  assign \s9_addr_o[18]_pad  = ~n49020 ;
  assign \s9_addr_o[19]_pad  = ~n49043 ;
  assign \s9_addr_o[1]_pad  = ~n49066 ;
  assign \s9_addr_o[20]_pad  = ~n49089 ;
  assign \s9_addr_o[21]_pad  = ~n49112 ;
  assign \s9_addr_o[22]_pad  = ~n49135 ;
  assign \s9_addr_o[23]_pad  = ~n49158 ;
  assign \s9_addr_o[24]_pad  = ~n49181 ;
  assign \s9_addr_o[25]_pad  = ~n49204 ;
  assign \s9_addr_o[26]_pad  = ~n49227 ;
  assign \s9_addr_o[27]_pad  = ~n49250 ;
  assign \s9_addr_o[28]_pad  = ~n49273 ;
  assign \s9_addr_o[29]_pad  = ~n49296 ;
  assign \s9_addr_o[2]_pad  = ~n49319 ;
  assign \s9_addr_o[30]_pad  = ~n49342 ;
  assign \s9_addr_o[31]_pad  = ~n49365 ;
  assign \s9_addr_o[3]_pad  = ~n49388 ;
  assign \s9_addr_o[4]_pad  = ~n49411 ;
  assign \s9_addr_o[5]_pad  = ~n49434 ;
  assign \s9_addr_o[6]_pad  = ~n49457 ;
  assign \s9_addr_o[7]_pad  = ~n49480 ;
  assign \s9_addr_o[8]_pad  = ~n49503 ;
  assign \s9_addr_o[9]_pad  = ~n49526 ;
  assign \s9_data_o[0]_pad  = ~n49549 ;
  assign \s9_data_o[10]_pad  = ~n49572 ;
  assign \s9_data_o[11]_pad  = ~n49595 ;
  assign \s9_data_o[12]_pad  = ~n49618 ;
  assign \s9_data_o[13]_pad  = ~n49641 ;
  assign \s9_data_o[14]_pad  = ~n49664 ;
  assign \s9_data_o[15]_pad  = ~n49687 ;
  assign \s9_data_o[16]_pad  = ~n49710 ;
  assign \s9_data_o[17]_pad  = ~n49733 ;
  assign \s9_data_o[18]_pad  = ~n49756 ;
  assign \s9_data_o[19]_pad  = ~n49779 ;
  assign \s9_data_o[1]_pad  = ~n49802 ;
  assign \s9_data_o[20]_pad  = ~n49825 ;
  assign \s9_data_o[21]_pad  = ~n49848 ;
  assign \s9_data_o[22]_pad  = ~n49871 ;
  assign \s9_data_o[23]_pad  = ~n49894 ;
  assign \s9_data_o[24]_pad  = ~n49917 ;
  assign \s9_data_o[25]_pad  = ~n49940 ;
  assign \s9_data_o[26]_pad  = ~n49963 ;
  assign \s9_data_o[27]_pad  = ~n49986 ;
  assign \s9_data_o[28]_pad  = ~n50009 ;
  assign \s9_data_o[29]_pad  = ~n50032 ;
  assign \s9_data_o[2]_pad  = ~n50055 ;
  assign \s9_data_o[30]_pad  = ~n50078 ;
  assign \s9_data_o[31]_pad  = ~n50101 ;
  assign \s9_data_o[3]_pad  = ~n50124 ;
  assign \s9_data_o[4]_pad  = ~n50147 ;
  assign \s9_data_o[5]_pad  = ~n50170 ;
  assign \s9_data_o[6]_pad  = ~n50193 ;
  assign \s9_data_o[7]_pad  = ~n50216 ;
  assign \s9_data_o[8]_pad  = ~n50239 ;
  assign \s9_data_o[9]_pad  = ~n50262 ;
  assign \s9_sel_o[0]_pad  = ~n50285 ;
  assign \s9_sel_o[1]_pad  = ~n50308 ;
  assign \s9_sel_o[2]_pad  = ~n50331 ;
  assign \s9_sel_o[3]_pad  = ~n50354 ;
  assign \s9_stb_o_pad  = ~n50385 ;
  assign \s9_we_o_pad  = ~n50408 ;
endmodule
