module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, \j0_pad , j_pad, \k0_pad , k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \a1_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u0_pad , \v0_pad , \w0_pad , \x0_pad , \y0_pad , \z0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \a1_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u0_pad  ;
	output \v0_pad  ;
	output \w0_pad  ;
	output \x0_pad  ;
	output \y0_pad  ;
	output \z0_pad  ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\k0_pad ,
		u_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		s_pad,
		u_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		m_pad,
		t_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\d0_pad ,
		t_pad,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		_w38_,
		_w39_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w37_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		u_pad,
		v_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		d_pad,
		t_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		t_pad,
		w_pad,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		_w38_,
		_w45_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w44_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		u_pad,
		w_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		c_pad,
		t_pad,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		t_pad,
		x_pad,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		_w38_,
		_w51_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w50_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		u_pad,
		x_pad,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		b_pad,
		t_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		t_pad,
		y_pad,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		_w38_,
		_w57_,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w56_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		u_pad,
		y_pad,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		a_pad,
		t_pad,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		q_pad,
		t_pad,
		_w64_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		_w38_,
		_w63_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		_w64_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w62_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		u_pad,
		z_pad,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		h_pad,
		t_pad,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\a0_pad ,
		t_pad,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		_w38_,
		_w69_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w68_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\a0_pad ,
		u_pad,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		g_pad,
		t_pad,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\b0_pad ,
		t_pad,
		_w76_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		_w38_,
		_w75_,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w74_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\b0_pad ,
		u_pad,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		f_pad,
		t_pad,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\c0_pad ,
		t_pad,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		_w38_,
		_w81_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w80_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\c0_pad ,
		u_pad,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		e_pad,
		t_pad,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		t_pad,
		v_pad,
		_w88_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		_w38_,
		_w87_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w88_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w86_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		\d0_pad ,
		u_pad,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		l_pad,
		t_pad,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\e0_pad ,
		t_pad,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		_w38_,
		_w93_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w92_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\e0_pad ,
		u_pad,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		k_pad,
		t_pad,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\f0_pad ,
		t_pad,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		_w38_,
		_w99_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w98_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\f0_pad ,
		u_pad,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		j_pad,
		t_pad,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\g0_pad ,
		t_pad,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		_w38_,
		_w105_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w104_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\g0_pad ,
		u_pad,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		i_pad,
		t_pad,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		t_pad,
		z_pad,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		_w38_,
		_w111_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w112_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w110_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\h0_pad ,
		u_pad,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		p_pad,
		t_pad,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\i0_pad ,
		t_pad,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w38_,
		_w117_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w116_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		\i0_pad ,
		u_pad,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		o_pad,
		t_pad,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\j0_pad ,
		t_pad,
		_w124_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w38_,
		_w123_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w124_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w122_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\j0_pad ,
		u_pad,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		n_pad,
		t_pad,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\k0_pad ,
		t_pad,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		_w38_,
		_w129_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w128_,
		_w132_,
		_w133_
	);
	assign \a1_pad  = _w43_ ;
	assign \l0_pad  = _w49_ ;
	assign \m0_pad  = _w55_ ;
	assign \n0_pad  = _w61_ ;
	assign \o0_pad  = _w67_ ;
	assign \p0_pad  = _w73_ ;
	assign \q0_pad  = _w79_ ;
	assign \r0_pad  = _w85_ ;
	assign \s0_pad  = _w91_ ;
	assign \t0_pad  = _w97_ ;
	assign \u0_pad  = _w103_ ;
	assign \v0_pad  = _w109_ ;
	assign \w0_pad  = _w115_ ;
	assign \x0_pad  = _w121_ ;
	assign \y0_pad  = _w127_ ;
	assign \z0_pad  = _w133_ ;
endmodule;