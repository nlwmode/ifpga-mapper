module top (\g108_reg/NET0131 , \g109_pad , \g1212_reg/NET0131 , \g1218_reg/NET0131 , \g1223_reg/NET0131 , \g1227_reg/NET0131 , \g1231_reg/NET0131 , \g1235_reg/NET0131 , \g1240_reg/NET0131 , \g1245_reg/NET0131 , \g1250_reg/NET0131 , \g1255_reg/NET0131 , \g1260_reg/NET0131 , \g1265_reg/NET0131 , \g1270_reg/NET0131 , \g1275_reg/NET0131 , \g1280_reg/NET0131 , \g1284_reg/NET0131 , \g1289_reg/NET0131 , \g1292_reg/NET0131 , \g1296_reg/NET0131 , \g1300_reg/NET0131 , \g1304_reg/NET0131 , \g1336_reg/NET0131 , \g1341_reg/NET0131 , \g1346_reg/NET0131 , \g1351_reg/NET0131 , \g1361_reg/NET0131 , \g1362_reg/NET0131 , \g1365_reg/NET0131 , \g1368_reg/NET0131 , \g1371_reg/NET0131 , \g1374_reg/NET0131 , \g1377_reg/NET0131 , \g1380_reg/NET0131 , \g1383_reg/NET0131 , \g1386_reg/NET0131 , \g1389_reg/NET0131 , \g1397_reg/NET0131 , \g1400_reg/NET0131 , \g1615_reg/NET0131 , \g1618_reg/NET0131 , \g1621_reg/NET0131 , \g1624_reg/NET0131 , \g1627_reg/NET0131 , \g1630_reg/NET0131 , \g1633_reg/NET0131 , \g1636_reg/NET0131 , \g1718_reg/NET0131 , \g186_reg/NET0131 , \g192_reg/NET0131 , \g197_reg/NET0131 , \g201_reg/NET0131 , \g207_reg/NET0131 , \g213_reg/NET0131 , \g219_reg/NET0131 , \g225_reg/NET0131 , \g231_reg/NET0131 , \g2355_pad , \g237_reg/NET0131 , \g243_reg/NET0131 , \g248_reg/NET0131 , \g3007_pad , \g305_reg/NET0131 , \g3069_pad , \g309_reg/NET0131 , \g312_reg/NET0131 , \g315_reg/NET0131 , \g318_reg/NET0131 , \g321_reg/NET0131 , \g324_reg/NET0131 , \g327_reg/NET0131 , \g330_reg/NET0131 , \g333_reg/NET0131 , \g369_reg/NET0131 , \g374_reg/NET0131 , \g378_reg/NET0131 , \g382_reg/NET0131 , \g386_reg/NET0131 , \g391_reg/NET0131 , \g396_reg/NET0131 , \g401_reg/NET0131 , \g406_reg/NET0131 , \g411_reg/NET0131 , \g416_reg/NET0131 , \g4173_pad , \g4174_pad , \g4175_pad , \g4176_pad , \g4177_pad , \g4178_pad , \g4179_pad , \g4180_pad , \g4181_pad , \g421_reg/NET0131 , \g426_reg/NET0131 , \g431_reg/NET0131 , \g435_reg/NET0131 , \g440_reg/NET0131 , \g444_reg/NET0131 , \g448_reg/NET0131 , \g452_reg/NET0131 , \g546_reg/NET0131 , \g549_reg/NET0131 , \g554_reg/NET0131 , \g557_reg/NET0131 , \g560_reg/NET0131 , \g563_reg/NET0131 , \g566_reg/NET0131 , \g569_reg/NET0131 , \g572_reg/NET0131 , \g575_reg/NET0131 , \g741_pad , \g742_pad , \g743_pad , \g744_pad , \g757_reg/NET0131 , \g876_reg/NET0131 , \g971_reg/NET0131 , \g976_reg/NET0131 , \g981_reg/NET0131 , \g986_reg/NET0131 , \g21280/_0_ , \g21281/_0_ , \g21282/_0_ , \g21307/_0_ , \g21322/_0_ , \g21333/_0_ , \g21334/_0_ , \g21338/_0_ , \g21350/_0_ , \g21355/_0_ , \g21356/_0_ , \g21357/_0_ , \g21358/_1_ , \g21359/_0_ , \g21370/_0_ , \g21371/_0_ , \g21378/_0_ , \g21379/_0_ , \g21380/_1_ , \g21381/_0_ , \g21390/_0_ , \g21394/_0_ , \g21396/_0_ , \g21397/_0_ , \g21398/_1_ , \g21412/_0_ , \g21413/_0_ , \g21419/_0_ , \g21420/_00_ , \g21421/_00_ , \g21424/_0_ , \g21425/_0_ , \g21426/_1_ , \g21437/_0_ , \g21444/_0_ , \g21450/_0_ , \g21455/_0_ , \g21457/_0_ , \g21458/_1_ , \g21459/_0_ , \g21470/_0_ , \g21486/_0_ , \g21487/_0_ , \g21495/_0_ , \g21498/_1_ , \g21499/_0_ , \g21500/_0_ , \g21502/_0_ , \g21503/_0_ , \g21508/_0_ , \g21509/_0_ , \g21510/_0_ , \g21511/_0_ , \g21515/_0_ , \g21520/_0_ , \g21523/_0_ , \g21524/_0_ , \g21525/_0_ , \g21538/_0_ , \g21544/_0_ , \g21550/_1_ , \g21562/_0_ , \g21563/_0_ , \g21584/_0_ , \g21591/_0_ , \g21593/_0_ , \g21601/_3_ , \g21603/_3_ , \g21605/_3_ , \g21607/_3_ , \g21609/_3_ , \g21611/_3_ , \g21613/_3_ , \g21615/_3_ , \g21617/_3_ , \g21619/_3_ , \g21621/_3_ , \g21623/_3_ , \g21625/_3_ , \g21627/_3_ , \g21640/_0_ , \g21641/_0_ , \g21642/_0_ , \g21693/_0_ , \g21694/_0_ , \g21735/_2_ , \g21745/_2_ , \g21796/_0_ , \g21799/_0_ , \g21803/_0_ , \g21812/_0_ , \g21814/_0_ , \g21816/_0_ , \g21828/_0_ , \g22203/_0_ , \g22260/_1_ , \g22317/_0_ , \g22339/_0_ , \g22392/_0_ , \g22395/_1_ , \g2601_pad , \g27_dup/_0_ , \g5816_pad );
	input \g108_reg/NET0131  ;
	input \g109_pad  ;
	input \g1212_reg/NET0131  ;
	input \g1218_reg/NET0131  ;
	input \g1223_reg/NET0131  ;
	input \g1227_reg/NET0131  ;
	input \g1231_reg/NET0131  ;
	input \g1235_reg/NET0131  ;
	input \g1240_reg/NET0131  ;
	input \g1245_reg/NET0131  ;
	input \g1250_reg/NET0131  ;
	input \g1255_reg/NET0131  ;
	input \g1260_reg/NET0131  ;
	input \g1265_reg/NET0131  ;
	input \g1270_reg/NET0131  ;
	input \g1275_reg/NET0131  ;
	input \g1280_reg/NET0131  ;
	input \g1284_reg/NET0131  ;
	input \g1289_reg/NET0131  ;
	input \g1292_reg/NET0131  ;
	input \g1296_reg/NET0131  ;
	input \g1300_reg/NET0131  ;
	input \g1304_reg/NET0131  ;
	input \g1336_reg/NET0131  ;
	input \g1341_reg/NET0131  ;
	input \g1346_reg/NET0131  ;
	input \g1351_reg/NET0131  ;
	input \g1361_reg/NET0131  ;
	input \g1362_reg/NET0131  ;
	input \g1365_reg/NET0131  ;
	input \g1368_reg/NET0131  ;
	input \g1371_reg/NET0131  ;
	input \g1374_reg/NET0131  ;
	input \g1377_reg/NET0131  ;
	input \g1380_reg/NET0131  ;
	input \g1383_reg/NET0131  ;
	input \g1386_reg/NET0131  ;
	input \g1389_reg/NET0131  ;
	input \g1397_reg/NET0131  ;
	input \g1400_reg/NET0131  ;
	input \g1615_reg/NET0131  ;
	input \g1618_reg/NET0131  ;
	input \g1621_reg/NET0131  ;
	input \g1624_reg/NET0131  ;
	input \g1627_reg/NET0131  ;
	input \g1630_reg/NET0131  ;
	input \g1633_reg/NET0131  ;
	input \g1636_reg/NET0131  ;
	input \g1718_reg/NET0131  ;
	input \g186_reg/NET0131  ;
	input \g192_reg/NET0131  ;
	input \g197_reg/NET0131  ;
	input \g201_reg/NET0131  ;
	input \g207_reg/NET0131  ;
	input \g213_reg/NET0131  ;
	input \g219_reg/NET0131  ;
	input \g225_reg/NET0131  ;
	input \g231_reg/NET0131  ;
	input \g2355_pad  ;
	input \g237_reg/NET0131  ;
	input \g243_reg/NET0131  ;
	input \g248_reg/NET0131  ;
	input \g3007_pad  ;
	input \g305_reg/NET0131  ;
	input \g3069_pad  ;
	input \g309_reg/NET0131  ;
	input \g312_reg/NET0131  ;
	input \g315_reg/NET0131  ;
	input \g318_reg/NET0131  ;
	input \g321_reg/NET0131  ;
	input \g324_reg/NET0131  ;
	input \g327_reg/NET0131  ;
	input \g330_reg/NET0131  ;
	input \g333_reg/NET0131  ;
	input \g369_reg/NET0131  ;
	input \g374_reg/NET0131  ;
	input \g378_reg/NET0131  ;
	input \g382_reg/NET0131  ;
	input \g386_reg/NET0131  ;
	input \g391_reg/NET0131  ;
	input \g396_reg/NET0131  ;
	input \g401_reg/NET0131  ;
	input \g406_reg/NET0131  ;
	input \g411_reg/NET0131  ;
	input \g416_reg/NET0131  ;
	input \g4173_pad  ;
	input \g4174_pad  ;
	input \g4175_pad  ;
	input \g4176_pad  ;
	input \g4177_pad  ;
	input \g4178_pad  ;
	input \g4179_pad  ;
	input \g4180_pad  ;
	input \g4181_pad  ;
	input \g421_reg/NET0131  ;
	input \g426_reg/NET0131  ;
	input \g431_reg/NET0131  ;
	input \g435_reg/NET0131  ;
	input \g440_reg/NET0131  ;
	input \g444_reg/NET0131  ;
	input \g448_reg/NET0131  ;
	input \g452_reg/NET0131  ;
	input \g546_reg/NET0131  ;
	input \g549_reg/NET0131  ;
	input \g554_reg/NET0131  ;
	input \g557_reg/NET0131  ;
	input \g560_reg/NET0131  ;
	input \g563_reg/NET0131  ;
	input \g566_reg/NET0131  ;
	input \g569_reg/NET0131  ;
	input \g572_reg/NET0131  ;
	input \g575_reg/NET0131  ;
	input \g741_pad  ;
	input \g742_pad  ;
	input \g743_pad  ;
	input \g744_pad  ;
	input \g757_reg/NET0131  ;
	input \g876_reg/NET0131  ;
	input \g971_reg/NET0131  ;
	input \g976_reg/NET0131  ;
	input \g981_reg/NET0131  ;
	input \g986_reg/NET0131  ;
	output \g21280/_0_  ;
	output \g21281/_0_  ;
	output \g21282/_0_  ;
	output \g21307/_0_  ;
	output \g21322/_0_  ;
	output \g21333/_0_  ;
	output \g21334/_0_  ;
	output \g21338/_0_  ;
	output \g21350/_0_  ;
	output \g21355/_0_  ;
	output \g21356/_0_  ;
	output \g21357/_0_  ;
	output \g21358/_1_  ;
	output \g21359/_0_  ;
	output \g21370/_0_  ;
	output \g21371/_0_  ;
	output \g21378/_0_  ;
	output \g21379/_0_  ;
	output \g21380/_1_  ;
	output \g21381/_0_  ;
	output \g21390/_0_  ;
	output \g21394/_0_  ;
	output \g21396/_0_  ;
	output \g21397/_0_  ;
	output \g21398/_1_  ;
	output \g21412/_0_  ;
	output \g21413/_0_  ;
	output \g21419/_0_  ;
	output \g21420/_00_  ;
	output \g21421/_00_  ;
	output \g21424/_0_  ;
	output \g21425/_0_  ;
	output \g21426/_1_  ;
	output \g21437/_0_  ;
	output \g21444/_0_  ;
	output \g21450/_0_  ;
	output \g21455/_0_  ;
	output \g21457/_0_  ;
	output \g21458/_1_  ;
	output \g21459/_0_  ;
	output \g21470/_0_  ;
	output \g21486/_0_  ;
	output \g21487/_0_  ;
	output \g21495/_0_  ;
	output \g21498/_1_  ;
	output \g21499/_0_  ;
	output \g21500/_0_  ;
	output \g21502/_0_  ;
	output \g21503/_0_  ;
	output \g21508/_0_  ;
	output \g21509/_0_  ;
	output \g21510/_0_  ;
	output \g21511/_0_  ;
	output \g21515/_0_  ;
	output \g21520/_0_  ;
	output \g21523/_0_  ;
	output \g21524/_0_  ;
	output \g21525/_0_  ;
	output \g21538/_0_  ;
	output \g21544/_0_  ;
	output \g21550/_1_  ;
	output \g21562/_0_  ;
	output \g21563/_0_  ;
	output \g21584/_0_  ;
	output \g21591/_0_  ;
	output \g21593/_0_  ;
	output \g21601/_3_  ;
	output \g21603/_3_  ;
	output \g21605/_3_  ;
	output \g21607/_3_  ;
	output \g21609/_3_  ;
	output \g21611/_3_  ;
	output \g21613/_3_  ;
	output \g21615/_3_  ;
	output \g21617/_3_  ;
	output \g21619/_3_  ;
	output \g21621/_3_  ;
	output \g21623/_3_  ;
	output \g21625/_3_  ;
	output \g21627/_3_  ;
	output \g21640/_0_  ;
	output \g21641/_0_  ;
	output \g21642/_0_  ;
	output \g21693/_0_  ;
	output \g21694/_0_  ;
	output \g21735/_2_  ;
	output \g21745/_2_  ;
	output \g21796/_0_  ;
	output \g21799/_0_  ;
	output \g21803/_0_  ;
	output \g21812/_0_  ;
	output \g21814/_0_  ;
	output \g21816/_0_  ;
	output \g21828/_0_  ;
	output \g22203/_0_  ;
	output \g22260/_1_  ;
	output \g22317/_0_  ;
	output \g22339/_0_  ;
	output \g22392/_0_  ;
	output \g22395/_1_  ;
	output \g2601_pad  ;
	output \g27_dup/_0_  ;
	output \g5816_pad  ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\g378_reg/NET0131 ,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\g382_reg/NET0131 ,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\g309_reg/NET0131 ,
		\g416_reg/NET0131 ,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\g333_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\g321_reg/NET0131 ,
		\g391_reg/NET0131 ,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\g333_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w129_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\g309_reg/NET0131 ,
		\g416_reg/NET0131 ,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\g327_reg/NET0131 ,
		\g401_reg/NET0131 ,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\g327_reg/NET0131 ,
		\g401_reg/NET0131 ,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w131_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\g324_reg/NET0131 ,
		\g396_reg/NET0131 ,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\g324_reg/NET0131 ,
		\g396_reg/NET0131 ,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w134_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\g312_reg/NET0131 ,
		\g421_reg/NET0131 ,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\g312_reg/NET0131 ,
		\g421_reg/NET0131 ,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\g330_reg/NET0131 ,
		\g406_reg/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\g330_reg/NET0131 ,
		\g406_reg/NET0131 ,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\g315_reg/NET0131 ,
		\g426_reg/NET0131 ,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\g315_reg/NET0131 ,
		\g426_reg/NET0131 ,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\g318_reg/NET0131 ,
		\g386_reg/NET0131 ,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		\g318_reg/NET0131 ,
		\g386_reg/NET0131 ,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\g321_reg/NET0131 ,
		\g391_reg/NET0131 ,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\g431_reg/NET0131 ,
		\g435_reg/NET0131 ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\g386_reg/NET0131 ,
		\g391_reg/NET0131 ,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\g396_reg/NET0131 ,
		\g401_reg/NET0131 ,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\g406_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\g416_reg/NET0131 ,
		\g421_reg/NET0131 ,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\g426_reg/NET0131 ,
		\g440_reg/NET0131 ,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\g444_reg/NET0131 ,
		\g448_reg/NET0131 ,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\g452_reg/NET0131 ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w152_,
		_w153_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w150_,
		_w151_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w148_,
		_w149_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w155_,
		_w156_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\g431_reg/NET0131 ,
		\g435_reg/NET0131 ,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w148_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w161_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\g305_reg/NET0131 ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\g305_reg/NET0131 ,
		_w164_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w126_,
		_w127_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w128_,
		_w129_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w130_,
		_w140_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w141_,
		_w145_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w146_,
		_w147_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w168_,
		_w169_,
		_w173_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w133_,
		_w167_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w136_,
		_w139_,
		_w175_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w144_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w173_,
		_w174_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w172_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w176_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		_w165_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w166_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w125_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\g3007_pad ,
		\g876_reg/NET0131 ,
		_w183_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\g1212_reg/NET0131 ,
		\g757_reg/NET0131 ,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w183_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\g109_pad ,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w182_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\g976_reg/NET0131 ,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\g971_reg/NET0131 ,
		\g976_reg/NET0131 ,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\g971_reg/NET0131 ,
		\g976_reg/NET0131 ,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w186_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w182_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w188_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\g981_reg/NET0131 ,
		_w187_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\g981_reg/NET0131 ,
		_w189_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\g981_reg/NET0131 ,
		_w189_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w196_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w186_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w182_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w195_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\g986_reg/NET0131 ,
		_w187_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\g986_reg/NET0131 ,
		_w196_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\g986_reg/NET0131 ,
		_w196_,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w186_,
		_w203_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w182_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w202_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\g1386_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\g1386_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\g197_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\g197_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\g1362_reg/NET0131 ,
		\g1365_reg/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\g1368_reg/NET0131 ,
		\g1371_reg/NET0131 ,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		\g1374_reg/NET0131 ,
		\g1377_reg/NET0131 ,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\g1380_reg/NET0131 ,
		\g1383_reg/NET0131 ,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\g1397_reg/NET0131 ,
		\g1400_reg/NET0131 ,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\g186_reg/NET0131 ,
		\g192_reg/NET0131 ,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		\g207_reg/NET0131 ,
		\g213_reg/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\g219_reg/NET0131 ,
		\g225_reg/NET0131 ,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\g231_reg/NET0131 ,
		\g237_reg/NET0131 ,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\g243_reg/NET0131 ,
		\g248_reg/NET0131 ,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w221_,
		_w222_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		_w219_,
		_w220_,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w217_,
		_w218_,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w215_,
		_w216_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w209_,
		_w212_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w229_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w227_,
		_w228_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w225_,
		_w226_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w231_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w211_,
		_w214_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w235_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w211_,
		_w214_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\g109_pad ,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w237_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\g2355_pad ,
		\g557_reg/NET0131 ,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\g213_reg/NET0131 ,
		\g2355_pad ,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w241_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		\g2355_pad ,
		\g546_reg/NET0131 ,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\g186_reg/NET0131 ,
		\g2355_pad ,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\g1615_reg/NET0131 ,
		\g2355_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w242_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\g1718_reg/NET0131 ,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\g2355_pad ,
		\g560_reg/NET0131 ,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\g219_reg/NET0131 ,
		\g2355_pad ,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\g1618_reg/NET0131 ,
		\g2355_pad ,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w245_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		\g1718_reg/NET0131 ,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		\g2355_pad ,
		\g554_reg/NET0131 ,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\g207_reg/NET0131 ,
		\g2355_pad ,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\g1621_reg/NET0131 ,
		\g2355_pad ,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w251_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\g1718_reg/NET0131 ,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\g109_pad ,
		\g186_reg/NET0131 ,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		\g2355_pad ,
		\g563_reg/NET0131 ,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\g225_reg/NET0131 ,
		\g2355_pad ,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\g109_pad ,
		\g1383_reg/NET0131 ,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\g1718_reg/NET0131 ,
		_w257_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\g1624_reg/NET0131 ,
		\g2355_pad ,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w264_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		\g1718_reg/NET0131 ,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\g109_pad ,
		\g207_reg/NET0131 ,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		\g2355_pad ,
		\g566_reg/NET0131 ,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		\g231_reg/NET0131 ,
		\g2355_pad ,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\g109_pad ,
		\g1380_reg/NET0131 ,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\g1627_reg/NET0131 ,
		\g2355_pad ,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w273_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\g1718_reg/NET0131 ,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\g2355_pad ,
		\g569_reg/NET0131 ,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\g2355_pad ,
		\g237_reg/NET0131 ,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\g109_pad ,
		\g213_reg/NET0131 ,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\g4173_pad ,
		\g4174_pad ,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\g4175_pad ,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\g4176_pad ,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\g4177_pad ,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\g4178_pad ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\g4179_pad ,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\g4180_pad ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\g4181_pad ,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\g4181_pad ,
		_w289_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		\g1718_reg/NET0131 ,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		\g109_pad ,
		_w290_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w292_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\g109_pad ,
		\g1377_reg/NET0131 ,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\g1630_reg/NET0131 ,
		\g2355_pad ,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w280_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\g1718_reg/NET0131 ,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\g1235_reg/NET0131 ,
		\g1250_reg/NET0131 ,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\g1265_reg/NET0131 ,
		\g1275_reg/NET0131 ,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\g1240_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\g1255_reg/NET0131 ,
		\g1260_reg/NET0131 ,
		_w303_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		\g1270_reg/NET0131 ,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w302_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\g1292_reg/NET0131 ,
		\g1296_reg/NET0131 ,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		\g1300_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w301_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w305_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\g1280_reg/NET0131 ,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\g1284_reg/NET0131 ,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		\g1280_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w312_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		_w301_,
		_w305_,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\g1218_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\g1227_reg/NET0131 ,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w317_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\g1231_reg/NET0131 ,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w316_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		\g1361_reg/NET0131 ,
		\g3069_pad ,
		_w323_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		\g108_reg/NET0131 ,
		\g1212_reg/NET0131 ,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		_w323_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\g109_pad ,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w322_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\g1346_reg/NET0131 ,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w322_,
		_w326_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\g1336_reg/NET0131 ,
		\g1341_reg/NET0131 ,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		\g1346_reg/NET0131 ,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		\g1346_reg/NET0131 ,
		_w330_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w331_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		_w329_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w328_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\g1351_reg/NET0131 ,
		_w327_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\g1351_reg/NET0131 ,
		_w332_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\g1351_reg/NET0131 ,
		_w332_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w337_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w329_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w336_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		\g2355_pad ,
		\g572_reg/NET0131 ,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\g2355_pad ,
		\g243_reg/NET0131 ,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		\g109_pad ,
		\g219_reg/NET0131 ,
		_w345_
	);
	LUT2 #(
		.INIT('h2)
	) name223 (
		\g109_pad ,
		\g1718_reg/NET0131 ,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		\g4180_pad ,
		_w288_,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w289_,
		_w346_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w347_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		\g109_pad ,
		\g1371_reg/NET0131 ,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		\g1633_reg/NET0131 ,
		\g2355_pad ,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		\g1718_reg/NET0131 ,
		_w343_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\g109_pad ,
		\g225_reg/NET0131 ,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		\g4179_pad ,
		_w287_,
		_w355_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w288_,
		_w346_,
		_w356_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		\g2355_pad ,
		\g575_reg/NET0131 ,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		\g2355_pad ,
		\g248_reg/NET0131 ,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w358_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\g109_pad ,
		\g1368_reg/NET0131 ,
		_w361_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		\g1636_reg/NET0131 ,
		\g2355_pad ,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		\g1718_reg/NET0131 ,
		_w359_,
		_w363_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		\g4178_pad ,
		_w286_,
		_w365_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w287_,
		_w346_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w365_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		\g109_pad ,
		\g231_reg/NET0131 ,
		_w368_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\g109_pad ,
		\g1212_reg/NET0131 ,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\g1231_reg/NET0131 ,
		_w319_,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		_w317_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\g1218_reg/NET0131 ,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		\g1218_reg/NET0131 ,
		_w371_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w369_,
		_w372_,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w373_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		\g1223_reg/NET0131 ,
		_w372_,
		_w376_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\g1223_reg/NET0131 ,
		_w372_,
		_w377_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		_w369_,
		_w376_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		_w377_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		\g1227_reg/NET0131 ,
		_w318_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name258 (
		\g109_pad ,
		_w319_,
		_w381_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w380_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w371_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\g1227_reg/NET0131 ,
		_w369_,
		_w384_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w371_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w383_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		\g1231_reg/NET0131 ,
		_w320_,
		_w387_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		_w369_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		\g369_reg/NET0131 ,
		_w125_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		_w369_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\g369_reg/NET0131 ,
		\g374_reg/NET0131 ,
		_w391_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w123_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w125_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		_w369_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		\g382_reg/NET0131 ,
		_w124_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		\g378_reg/NET0131 ,
		_w123_,
		_w396_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		_w369_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w395_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		\g382_reg/NET0131 ,
		_w124_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		_w369_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		\g109_pad ,
		_w317_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		\g1275_reg/NET0131 ,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w314_,
		_w321_,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w402_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		\g4177_pad ,
		_w285_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w286_,
		_w346_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w405_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		\g109_pad ,
		\g1365_reg/NET0131 ,
		_w408_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		\g2355_pad ,
		\g549_reg/NET0131 ,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\g192_reg/NET0131 ,
		\g2355_pad ,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w409_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		\g201_reg/NET0131 ,
		\g2355_pad ,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\g109_pad ,
		\g237_reg/NET0131 ,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		\g4176_pad ,
		_w284_,
		_w414_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		_w285_,
		_w346_,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		_w414_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		\g1718_reg/NET0131 ,
		_w410_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		\g109_pad ,
		\g1362_reg/NET0131 ,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		\g4173_pad ,
		\g4174_pad ,
		_w419_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w283_,
		_w346_,
		_w420_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w419_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		\g1275_reg/NET0131 ,
		_w317_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		\g1235_reg/NET0131 ,
		_w401_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		\g1235_reg/NET0131 ,
		_w317_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		\g1240_reg/NET0131 ,
		_w401_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		\g1240_reg/NET0131 ,
		_w317_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\g1245_reg/NET0131 ,
		_w401_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		\g1245_reg/NET0131 ,
		_w317_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		\g1250_reg/NET0131 ,
		_w401_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w431_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		\g1250_reg/NET0131 ,
		_w317_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		\g1255_reg/NET0131 ,
		_w401_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w434_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\g1255_reg/NET0131 ,
		_w317_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		\g1260_reg/NET0131 ,
		_w401_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w437_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		\g1260_reg/NET0131 ,
		_w317_,
		_w440_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\g1265_reg/NET0131 ,
		_w401_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		_w440_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		\g1265_reg/NET0131 ,
		_w317_,
		_w443_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\g1270_reg/NET0131 ,
		_w401_,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w443_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\g1284_reg/NET0131 ,
		_w317_,
		_w446_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		\g1280_reg/NET0131 ,
		_w401_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w446_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\g1292_reg/NET0131 ,
		_w317_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		\g1284_reg/NET0131 ,
		_w401_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w449_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\g1296_reg/NET0131 ,
		_w317_,
		_w452_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\g1292_reg/NET0131 ,
		_w401_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w452_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		\g1300_reg/NET0131 ,
		_w317_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		\g1296_reg/NET0131 ,
		_w401_,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w455_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\g1304_reg/NET0131 ,
		_w317_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		\g1300_reg/NET0131 ,
		_w401_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w458_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		\g1270_reg/NET0131 ,
		_w317_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\g1304_reg/NET0131 ,
		_w401_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w461_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\g109_pad ,
		\g243_reg/NET0131 ,
		_w464_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\g4173_pad ,
		_w346_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		\g4175_pad ,
		_w283_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w284_,
		_w346_,
		_w467_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		\g109_pad ,
		\g1400_reg/NET0131 ,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\g1212_reg/NET0131 ,
		\g1289_reg/NET0131 ,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		\g109_pad ,
		\g741_pad ,
		_w471_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\g742_pad ,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		\g109_pad ,
		\g743_pad ,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\g744_pad ,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		\g109_pad ,
		\g1374_reg/NET0131 ,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		\g109_pad ,
		\g197_reg/NET0131 ,
		_w476_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		\g109_pad ,
		\g201_reg/NET0131 ,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		\g109_pad ,
		\g1389_reg/NET0131 ,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\g109_pad ,
		\g1397_reg/NET0131 ,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\g109_pad ,
		\g192_reg/NET0131 ,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\g109_pad ,
		\g248_reg/NET0131 ,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		\g1718_reg/NET0131 ,
		_w291_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w292_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		\g971_reg/NET0131 ,
		_w182_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		\g971_reg/NET0131 ,
		_w182_,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name363 (
		_w186_,
		_w484_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name364 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		\g1336_reg/NET0131 ,
		_w329_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		\g1336_reg/NET0131 ,
		_w327_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w488_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		\g1341_reg/NET0131 ,
		_w327_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		\g1336_reg/NET0131 ,
		\g1341_reg/NET0131 ,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w330_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		_w329_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w491_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		_w125_,
		_w164_,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		\g305_reg/NET0131 ,
		_w125_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		_w496_,
		_w497_,
		_w498_
	);
	assign \g21280/_0_  = _w194_ ;
	assign \g21281/_0_  = _w201_ ;
	assign \g21282/_0_  = _w208_ ;
	assign \g21307/_0_  = _w240_ ;
	assign \g21322/_0_  = _w243_ ;
	assign \g21333/_0_  = _w246_ ;
	assign \g21334/_0_  = _w249_ ;
	assign \g21338/_0_  = _w252_ ;
	assign \g21350/_0_  = _w255_ ;
	assign \g21355/_0_  = _w258_ ;
	assign \g21356/_0_  = _w261_ ;
	assign \g21357/_0_  = _w262_ ;
	assign \g21358/_1_  = _w245_ ;
	assign \g21359/_0_  = _w265_ ;
	assign \g21370/_0_  = _w266_ ;
	assign \g21371/_0_  = _w267_ ;
	assign \g21378/_0_  = _w270_ ;
	assign \g21379/_0_  = _w271_ ;
	assign \g21380/_1_  = _w257_ ;
	assign \g21381/_0_  = _w274_ ;
	assign \g21390/_0_  = _w275_ ;
	assign \g21394/_0_  = _w278_ ;
	assign \g21396/_0_  = _w281_ ;
	assign \g21397/_0_  = _w282_ ;
	assign \g21398/_1_  = _w242_ ;
	assign \g21412/_0_  = _w294_ ;
	assign \g21413/_0_  = _w295_ ;
	assign \g21419/_0_  = _w298_ ;
	assign \g21420/_00_  = _w335_ ;
	assign \g21421/_00_  = _w341_ ;
	assign \g21424/_0_  = _w344_ ;
	assign \g21425/_0_  = _w345_ ;
	assign \g21426/_1_  = _w251_ ;
	assign \g21437/_0_  = _w349_ ;
	assign \g21444/_0_  = _w350_ ;
	assign \g21450/_0_  = _w353_ ;
	assign \g21455/_0_  = _w354_ ;
	assign \g21457/_0_  = _w357_ ;
	assign \g21458/_1_  = _w264_ ;
	assign \g21459/_0_  = _w360_ ;
	assign \g21470/_0_  = _w361_ ;
	assign \g21486/_0_  = _w364_ ;
	assign \g21487/_0_  = _w367_ ;
	assign \g21495/_0_  = _w368_ ;
	assign \g21498/_1_  = _w273_ ;
	assign \g21499/_0_  = _w375_ ;
	assign \g21500/_0_  = _w379_ ;
	assign \g21502/_0_  = _w386_ ;
	assign \g21503/_0_  = _w388_ ;
	assign \g21508/_0_  = _w390_ ;
	assign \g21509/_0_  = _w394_ ;
	assign \g21510/_0_  = _w398_ ;
	assign \g21511/_0_  = _w400_ ;
	assign \g21515/_0_  = _w404_ ;
	assign \g21520/_0_  = _w407_ ;
	assign \g21523/_0_  = _w408_ ;
	assign \g21524/_0_  = _w411_ ;
	assign \g21525/_0_  = _w412_ ;
	assign \g21538/_0_  = _w280_ ;
	assign \g21544/_0_  = _w413_ ;
	assign \g21550/_1_  = _w204_ ;
	assign \g21562/_0_  = _w416_ ;
	assign \g21563/_0_  = _w417_ ;
	assign \g21584/_0_  = _w338_ ;
	assign \g21591/_0_  = _w418_ ;
	assign \g21593/_0_  = _w421_ ;
	assign \g21601/_3_  = _w424_ ;
	assign \g21603/_3_  = _w427_ ;
	assign \g21605/_3_  = _w430_ ;
	assign \g21607/_3_  = _w433_ ;
	assign \g21609/_3_  = _w436_ ;
	assign \g21611/_3_  = _w439_ ;
	assign \g21613/_3_  = _w442_ ;
	assign \g21615/_3_  = _w445_ ;
	assign \g21617/_3_  = _w448_ ;
	assign \g21619/_3_  = _w451_ ;
	assign \g21621/_3_  = _w454_ ;
	assign \g21623/_3_  = _w457_ ;
	assign \g21625/_3_  = _w460_ ;
	assign \g21627/_3_  = _w463_ ;
	assign \g21640/_0_  = _w464_ ;
	assign \g21641/_0_  = _w465_ ;
	assign \g21642/_0_  = _w468_ ;
	assign \g21693/_0_  = _w469_ ;
	assign \g21694/_0_  = _w470_ ;
	assign \g21735/_2_  = _w472_ ;
	assign \g21745/_2_  = _w474_ ;
	assign \g21796/_0_  = _w475_ ;
	assign \g21799/_0_  = _w476_ ;
	assign \g21803/_0_  = _w477_ ;
	assign \g21812/_0_  = _w478_ ;
	assign \g21814/_0_  = _w479_ ;
	assign \g21816/_0_  = _w480_ ;
	assign \g21828/_0_  = _w481_ ;
	assign \g22203/_0_  = _w483_ ;
	assign \g22260/_1_  = _w182_ ;
	assign \g22317/_0_  = _w487_ ;
	assign \g22339/_0_  = _w490_ ;
	assign \g22392/_0_  = _w495_ ;
	assign \g22395/_1_  = _w322_ ;
	assign \g2601_pad  = 1'b0;
	assign \g27_dup/_0_  = _w498_ ;
	assign \g5816_pad  = 1'b0;
endmodule;