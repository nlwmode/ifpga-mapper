module top (\G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G19_pad , \G20_pad , \G22_pad , \G23_pad , \G24_pad , \G25_pad , \G26_pad , \G28_pad , \G2_pad , \G30_pad , \G31_pad , \G32_pad , \G33_pad , \G34_pad , \G35_pad , \G3_pad , \G4_pad , \G5_pad , \G64_reg/NET0131 , \G65_reg/NET0131 , \G66_reg/NET0131 , \G69_reg/NET0131 , \G6_pad , \G70_reg/NET0131 , \G71_reg/NET0131 , \G72_reg/NET0131 , \G73_reg/NET0131 , \G74_reg/NET0131 , \G75_reg/NET0131 , \G76_reg/NET0131 , \G77_reg/NET0131 , \G79_reg/NET0131 , \G81_reg/NET0131 , \G8_pad , \G9_pad , \G100BF_pad , \G103BF_pad , \G104BF_pad , \G105BF_pad , \G107_pad , \G83_pad , \G84_pad , \G86BF_pad , \G89BF_pad , \G95BF_pad , \G96BF_pad , \G97BF_pad , \G98BF_pad , \G99BF_pad , \_al_n0 , \_al_n1 , \g1017/_3_ , \g1150/_0_ , \g1168/_0_ , \g1308/_1_ , \g1318/_0_ , \g1337/_2_ , \g1339/_1_ , \g16/_0_ , \g26/_2_ , \g27/_0_ , \g29/_0_ , \g867/_3_ , \g875/_0_ , \g898/_0_ , \g931/_0_ , \g938/_0_ , \g967/_0_ , \g987/_0_ );
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G19_pad  ;
	input \G20_pad  ;
	input \G22_pad  ;
	input \G23_pad  ;
	input \G24_pad  ;
	input \G25_pad  ;
	input \G26_pad  ;
	input \G28_pad  ;
	input \G2_pad  ;
	input \G30_pad  ;
	input \G31_pad  ;
	input \G32_pad  ;
	input \G33_pad  ;
	input \G34_pad  ;
	input \G35_pad  ;
	input \G3_pad  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G64_reg/NET0131  ;
	input \G65_reg/NET0131  ;
	input \G66_reg/NET0131  ;
	input \G69_reg/NET0131  ;
	input \G6_pad  ;
	input \G70_reg/NET0131  ;
	input \G71_reg/NET0131  ;
	input \G72_reg/NET0131  ;
	input \G73_reg/NET0131  ;
	input \G74_reg/NET0131  ;
	input \G75_reg/NET0131  ;
	input \G76_reg/NET0131  ;
	input \G77_reg/NET0131  ;
	input \G79_reg/NET0131  ;
	input \G81_reg/NET0131  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G100BF_pad  ;
	output \G103BF_pad  ;
	output \G104BF_pad  ;
	output \G105BF_pad  ;
	output \G107_pad  ;
	output \G83_pad  ;
	output \G84_pad  ;
	output \G86BF_pad  ;
	output \G89BF_pad  ;
	output \G95BF_pad  ;
	output \G96BF_pad  ;
	output \G97BF_pad  ;
	output \G98BF_pad  ;
	output \G99BF_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1017/_3_  ;
	output \g1150/_0_  ;
	output \g1168/_0_  ;
	output \g1308/_1_  ;
	output \g1318/_0_  ;
	output \g1337/_2_  ;
	output \g1339/_1_  ;
	output \g16/_0_  ;
	output \g26/_2_  ;
	output \g27/_0_  ;
	output \g29/_0_  ;
	output \g867/_3_  ;
	output \g875/_0_  ;
	output \g898/_0_  ;
	output \g931/_0_  ;
	output \g938/_0_  ;
	output \g967/_0_  ;
	output \g987/_0_  ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\G4_pad ,
		\G69_reg/NET0131 ,
		_w45_
	);
	LUT3 #(
		.INIT('hdf)
	) name1 (
		\G35_pad ,
		\G4_pad ,
		\G69_reg/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\G3_pad ,
		\G75_reg/NET0131 ,
		_w47_
	);
	LUT3 #(
		.INIT('h80)
	) name3 (
		\G14_pad ,
		\G3_pad ,
		\G75_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\G3_pad ,
		\G77_reg/NET0131 ,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\G11_pad ,
		\G3_pad ,
		_w50_
	);
	LUT3 #(
		.INIT('h8a)
	) name6 (
		\G24_pad ,
		\G2_pad ,
		\G66_reg/NET0131 ,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\G10_pad ,
		\G13_pad ,
		_w52_
	);
	LUT4 #(
		.INIT('h0100)
	) name8 (
		\G10_pad ,
		\G13_pad ,
		\G3_pad ,
		\G9_pad ,
		_w53_
	);
	LUT4 #(
		.INIT('h0020)
	) name9 (
		\G77_reg/NET0131 ,
		_w50_,
		_w51_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w49_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('he)
	) name11 (
		_w49_,
		_w54_,
		_w56_
	);
	LUT3 #(
		.INIT('h04)
	) name12 (
		\G2_pad ,
		\G64_reg/NET0131 ,
		\G76_reg/NET0131 ,
		_w57_
	);
	LUT4 #(
		.INIT('h0002)
	) name13 (
		\G10_pad ,
		\G13_pad ,
		\G3_pad ,
		\G9_pad ,
		_w58_
	);
	LUT4 #(
		.INIT('h00c8)
	) name14 (
		\G11_pad ,
		\G23_pad ,
		\G3_pad ,
		\G65_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('hb)
	) name15 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT3 #(
		.INIT('h10)
	) name16 (
		\G2_pad ,
		\G3_pad ,
		\G64_reg/NET0131 ,
		_w61_
	);
	LUT4 #(
		.INIT('h1055)
	) name17 (
		_w57_,
		_w58_,
		_w59_,
		_w61_,
		_w62_
	);
	LUT4 #(
		.INIT('h0001)
	) name18 (
		\G10_pad ,
		\G13_pad ,
		\G3_pad ,
		\G9_pad ,
		_w63_
	);
	LUT4 #(
		.INIT('hc800)
	) name19 (
		\G11_pad ,
		\G22_pad ,
		\G3_pad ,
		\G75_reg/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w63_,
		_w64_,
		_w65_
	);
	LUT3 #(
		.INIT('h20)
	) name21 (
		\G14_pad ,
		_w63_,
		_w64_,
		_w66_
	);
	LUT4 #(
		.INIT('hfe00)
	) name22 (
		_w49_,
		_w54_,
		_w62_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w48_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\G15_pad ,
		\G76_reg/NET0131 ,
		_w69_
	);
	LUT4 #(
		.INIT('h45ff)
	) name25 (
		\G3_pad ,
		_w58_,
		_w59_,
		_w69_,
		_w70_
	);
	LUT3 #(
		.INIT('h57)
	) name26 (
		\G16_pad ,
		_w49_,
		_w54_,
		_w71_
	);
	LUT3 #(
		.INIT('h20)
	) name27 (
		\G18_pad ,
		\G4_pad ,
		\G79_reg/NET0131 ,
		_w72_
	);
	LUT3 #(
		.INIT('h20)
	) name28 (
		\G19_pad ,
		\G4_pad ,
		\G65_reg/NET0131 ,
		_w73_
	);
	LUT3 #(
		.INIT('h20)
	) name29 (
		\G20_pad ,
		\G4_pad ,
		\G81_reg/NET0131 ,
		_w74_
	);
	LUT3 #(
		.INIT('hc8)
	) name30 (
		\G11_pad ,
		\G22_pad ,
		\G3_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w63_,
		_w75_,
		_w76_
	);
	LUT4 #(
		.INIT('hfe00)
	) name32 (
		_w49_,
		_w54_,
		_w62_,
		_w76_,
		_w77_
	);
	LUT4 #(
		.INIT('h01ff)
	) name33 (
		_w49_,
		_w54_,
		_w62_,
		_w76_,
		_w78_
	);
	LUT4 #(
		.INIT('h0200)
	) name34 (
		\G10_pad ,
		\G13_pad ,
		\G3_pad ,
		\G9_pad ,
		_w79_
	);
	LUT3 #(
		.INIT('hc8)
	) name35 (
		\G11_pad ,
		\G25_pad ,
		\G3_pad ,
		_w80_
	);
	LUT2 #(
		.INIT('hb)
	) name36 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\G30_pad ,
		\G74_reg/NET0131 ,
		_w82_
	);
	LUT3 #(
		.INIT('h40)
	) name38 (
		_w63_,
		_w75_,
		_w82_,
		_w83_
	);
	LUT4 #(
		.INIT('h01ff)
	) name39 (
		_w49_,
		_w54_,
		_w62_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\G4_pad ,
		\G73_reg/NET0131 ,
		_w85_
	);
	LUT3 #(
		.INIT('hdf)
	) name41 (
		\G31_pad ,
		\G4_pad ,
		\G73_reg/NET0131 ,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\G32_pad ,
		\G72_reg/NET0131 ,
		_w87_
	);
	LUT3 #(
		.INIT('hbf)
	) name43 (
		_w58_,
		_w59_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\G4_pad ,
		\G71_reg/NET0131 ,
		_w89_
	);
	LUT3 #(
		.INIT('hdf)
	) name45 (
		\G33_pad ,
		\G4_pad ,
		\G71_reg/NET0131 ,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\G34_pad ,
		\G70_reg/NET0131 ,
		_w91_
	);
	LUT4 #(
		.INIT('hfbff)
	) name47 (
		_w50_,
		_w51_,
		_w53_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('h8000)
	) name48 (
		\G11_pad ,
		\G12_pad ,
		\G13_pad ,
		\G28_pad ,
		_w93_
	);
	LUT4 #(
		.INIT('hc800)
	) name49 (
		\G11_pad ,
		\G22_pad ,
		\G3_pad ,
		\G74_reg/NET0131 ,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w63_,
		_w94_,
		_w95_
	);
	LUT4 #(
		.INIT('hfe00)
	) name51 (
		_w49_,
		_w54_,
		_w62_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('hd)
	) name52 (
		_w85_,
		_w96_,
		_w97_
	);
	LUT3 #(
		.INIT('hd0)
	) name53 (
		\G2_pad ,
		\G5_pad ,
		\G76_reg/NET0131 ,
		_w98_
	);
	LUT4 #(
		.INIT('hba00)
	) name54 (
		\G3_pad ,
		_w58_,
		_w59_,
		_w98_,
		_w99_
	);
	LUT4 #(
		.INIT('hfe00)
	) name55 (
		_w49_,
		_w54_,
		_w62_,
		_w65_,
		_w100_
	);
	LUT4 #(
		.INIT('h4000)
	) name56 (
		\G4_pad ,
		\G5_pad ,
		\G71_reg/NET0131 ,
		\G72_reg/NET0131 ,
		_w101_
	);
	LUT3 #(
		.INIT('h40)
	) name57 (
		_w58_,
		_w59_,
		_w101_,
		_w102_
	);
	LUT4 #(
		.INIT('h0100)
	) name58 (
		_w47_,
		_w49_,
		_w54_,
		_w102_,
		_w103_
	);
	LUT3 #(
		.INIT('hba)
	) name59 (
		_w99_,
		_w100_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('he)
	) name60 (
		_w47_,
		_w100_,
		_w105_
	);
	LUT3 #(
		.INIT('hfb)
	) name61 (
		_w50_,
		_w51_,
		_w53_,
		_w106_
	);
	LUT3 #(
		.INIT('h54)
	) name62 (
		\G2_pad ,
		_w49_,
		_w54_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\G2_pad ,
		\G76_reg/NET0131 ,
		_w108_
	);
	LUT4 #(
		.INIT('hba00)
	) name64 (
		\G3_pad ,
		_w58_,
		_w59_,
		_w108_,
		_w109_
	);
	LUT3 #(
		.INIT('h10)
	) name65 (
		_w49_,
		_w54_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\G2_pad ,
		\G76_reg/NET0131 ,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\G2_pad ,
		\G3_pad ,
		_w112_
	);
	LUT4 #(
		.INIT('h040f)
	) name68 (
		_w58_,
		_w59_,
		_w111_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w47_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		_w65_,
		_w113_,
		_w115_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name71 (
		_w55_,
		_w62_,
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\G2_pad ,
		\G8_pad ,
		_w117_
	);
	LUT4 #(
		.INIT('hc040)
	) name73 (
		\G2_pad ,
		\G3_pad ,
		\G75_reg/NET0131 ,
		\G8_pad ,
		_w118_
	);
	LUT3 #(
		.INIT('h04)
	) name74 (
		_w63_,
		_w64_,
		_w117_,
		_w119_
	);
	LUT4 #(
		.INIT('hfe00)
	) name75 (
		_w49_,
		_w54_,
		_w62_,
		_w119_,
		_w120_
	);
	LUT3 #(
		.INIT('h10)
	) name76 (
		_w49_,
		_w54_,
		_w95_,
		_w121_
	);
	LUT4 #(
		.INIT('h0400)
	) name77 (
		\G4_pad ,
		\G73_reg/NET0131 ,
		\G76_reg/NET0131 ,
		\G8_pad ,
		_w122_
	);
	LUT4 #(
		.INIT('h1000)
	) name78 (
		\G3_pad ,
		\G4_pad ,
		\G73_reg/NET0131 ,
		\G8_pad ,
		_w123_
	);
	LUT4 #(
		.INIT('h040f)
	) name79 (
		_w58_,
		_w59_,
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		_w62_,
		_w124_,
		_w125_
	);
	LUT4 #(
		.INIT('hfeee)
	) name81 (
		_w118_,
		_w120_,
		_w121_,
		_w125_,
		_w126_
	);
	LUT4 #(
		.INIT('h0020)
	) name82 (
		\G10_pad ,
		\G13_pad ,
		\G72_reg/NET0131 ,
		\G9_pad ,
		_w127_
	);
	LUT4 #(
		.INIT('h4000)
	) name83 (
		_w58_,
		_w59_,
		_w89_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\G12_pad ,
		\G26_pad ,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT4 #(
		.INIT('h0e00)
	) name86 (
		\G11_pad ,
		\G3_pad ,
		\G4_pad ,
		\G69_reg/NET0131 ,
		_w131_
	);
	LUT4 #(
		.INIT('h0800)
	) name87 (
		\G70_reg/NET0131 ,
		_w51_,
		_w53_,
		_w131_,
		_w132_
	);
	LUT3 #(
		.INIT('h80)
	) name88 (
		\G9_pad ,
		_w52_,
		_w132_,
		_w133_
	);
	LUT4 #(
		.INIT('h0040)
	) name89 (
		\G4_pad ,
		\G73_reg/NET0131 ,
		\G74_reg/NET0131 ,
		\G9_pad ,
		_w134_
	);
	LUT4 #(
		.INIT('h2000)
	) name90 (
		_w52_,
		_w63_,
		_w75_,
		_w134_,
		_w135_
	);
	LUT4 #(
		.INIT('hfe00)
	) name91 (
		_w49_,
		_w54_,
		_w62_,
		_w135_,
		_w136_
	);
	LUT3 #(
		.INIT('h02)
	) name92 (
		_w130_,
		_w133_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\G2_pad ,
		\G6_pad ,
		_w138_
	);
	LUT3 #(
		.INIT('h0e)
	) name94 (
		_w49_,
		_w54_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\G6_pad ,
		\G76_reg/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		\G3_pad ,
		\G6_pad ,
		_w141_
	);
	LUT4 #(
		.INIT('h040f)
	) name97 (
		_w58_,
		_w59_,
		_w140_,
		_w141_,
		_w142_
	);
	LUT3 #(
		.INIT('h04)
	) name98 (
		_w47_,
		_w132_,
		_w142_,
		_w143_
	);
	LUT3 #(
		.INIT('hdc)
	) name99 (
		_w100_,
		_w139_,
		_w143_,
		_w144_
	);
	LUT3 #(
		.INIT('hf4)
	) name100 (
		_w77_,
		_w85_,
		_w96_,
		_w145_
	);
	LUT4 #(
		.INIT('h0020)
	) name101 (
		\G70_reg/NET0131 ,
		_w50_,
		_w51_,
		_w53_,
		_w146_
	);
	LUT2 #(
		.INIT('hd)
	) name102 (
		_w45_,
		_w146_,
		_w147_
	);
	LUT4 #(
		.INIT('haa8a)
	) name103 (
		_w45_,
		_w50_,
		_w51_,
		_w53_,
		_w148_
	);
	LUT2 #(
		.INIT('he)
	) name104 (
		_w146_,
		_w148_,
		_w149_
	);
	LUT4 #(
		.INIT('h20ff)
	) name105 (
		\G72_reg/NET0131 ,
		_w58_,
		_w59_,
		_w89_,
		_w150_
	);
	LUT4 #(
		.INIT('hef20)
	) name106 (
		\G72_reg/NET0131 ,
		_w58_,
		_w59_,
		_w89_,
		_w151_
	);
	assign \G100BF_pad  = _w46_ ;
	assign \G103BF_pad  = _w68_ ;
	assign \G104BF_pad  = _w70_ ;
	assign \G105BF_pad  = _w71_ ;
	assign \G107_pad  = _w72_ ;
	assign \G83_pad  = _w73_ ;
	assign \G84_pad  = _w74_ ;
	assign \G86BF_pad  = _w78_ ;
	assign \G89BF_pad  = _w81_ ;
	assign \G95BF_pad  = _w84_ ;
	assign \G96BF_pad  = _w86_ ;
	assign \G97BF_pad  = _w88_ ;
	assign \G98BF_pad  = _w90_ ;
	assign \G99BF_pad  = _w92_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1017/_3_  = _w93_ ;
	assign \g1150/_0_  = _w97_ ;
	assign \g1168/_0_  = _w104_ ;
	assign \g1308/_1_  = _w105_ ;
	assign \g1318/_0_  = _w106_ ;
	assign \g1337/_2_  = _w107_ ;
	assign \g1339/_1_  = _w56_ ;
	assign \g16/_0_  = _w110_ ;
	assign \g26/_2_  = _w116_ ;
	assign \g27/_0_  = _w126_ ;
	assign \g29/_0_  = _w60_ ;
	assign \g867/_3_  = _w137_ ;
	assign \g875/_0_  = _w144_ ;
	assign \g898/_0_  = _w145_ ;
	assign \g931/_0_  = _w147_ ;
	assign \g938/_0_  = _w149_ ;
	assign \g967/_0_  = _w150_ ;
	assign \g987/_0_  = _w151_ ;
endmodule;