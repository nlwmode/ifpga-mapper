module top( ADS_n_pad , \Address[0]_pad  , \Address[10]_pad  , \Address[11]_pad  , \Address[12]_pad  , \Address[13]_pad  , \Address[14]_pad  , \Address[15]_pad  , \Address[16]_pad  , \Address[17]_pad  , \Address[18]_pad  , \Address[19]_pad  , \Address[1]_pad  , \Address[20]_pad  , \Address[21]_pad  , \Address[22]_pad  , \Address[23]_pad  , \Address[24]_pad  , \Address[25]_pad  , \Address[26]_pad  , \Address[27]_pad  , \Address[28]_pad  , \Address[29]_pad  , \Address[2]_pad  , \Address[3]_pad  , \Address[4]_pad  , \Address[5]_pad  , \Address[6]_pad  , \Address[7]_pad  , \Address[8]_pad  , \Address[9]_pad  , \BE_n[0]_pad  , \BE_n[1]_pad  , \BE_n[2]_pad  , \BE_n[3]_pad  , \BS16_n_pad  , \ByteEnable_reg[0]/NET0131  , \ByteEnable_reg[1]/NET0131  , \ByteEnable_reg[2]/NET0131  , \ByteEnable_reg[3]/NET0131  , \CodeFetch_reg/NET0131  , D_C_n_pad , \DataWidth_reg[0]/NET0131  , \DataWidth_reg[1]/NET0131  , \Datai[0]_pad  , \Datai[10]_pad  , \Datai[11]_pad  , \Datai[12]_pad  , \Datai[13]_pad  , \Datai[14]_pad  , \Datai[15]_pad  , \Datai[16]_pad  , \Datai[17]_pad  , \Datai[18]_pad  , \Datai[19]_pad  , \Datai[1]_pad  , \Datai[20]_pad  , \Datai[21]_pad  , \Datai[22]_pad  , \Datai[23]_pad  , \Datai[24]_pad  , \Datai[25]_pad  , \Datai[26]_pad  , \Datai[27]_pad  , \Datai[28]_pad  , \Datai[29]_pad  , \Datai[2]_pad  , \Datai[30]_pad  , \Datai[31]_pad  , \Datai[3]_pad  , \Datai[4]_pad  , \Datai[5]_pad  , \Datai[6]_pad  , \Datai[7]_pad  , \Datai[8]_pad  , \Datai[9]_pad  , \Datao[0]_pad  , \Datao[10]_pad  , \Datao[11]_pad  , \Datao[12]_pad  , \Datao[13]_pad  , \Datao[14]_pad  , \Datao[15]_pad  , \Datao[16]_pad  , \Datao[17]_pad  , \Datao[18]_pad  , \Datao[19]_pad  , \Datao[1]_pad  , \Datao[20]_pad  , \Datao[21]_pad  , \Datao[23]_pad  , \Datao[24]_pad  , \Datao[25]_pad  , \Datao[26]_pad  , \Datao[27]_pad  , \Datao[28]_pad  , \Datao[29]_pad  , \Datao[2]_pad  , \Datao[30]_pad  , \Datao[3]_pad  , \Datao[4]_pad  , \Datao[5]_pad  , \Datao[6]_pad  , \Datao[7]_pad  , \Datao[8]_pad  , \Datao[9]_pad  , \Datao_reg[22]/NET0131  , \EAX_reg[0]/NET0131  , \EAX_reg[10]/NET0131  , \EAX_reg[11]/NET0131  , \EAX_reg[12]/NET0131  , \EAX_reg[13]/NET0131  , \EAX_reg[14]/NET0131  , \EAX_reg[15]/NET0131  , \EAX_reg[16]/NET0131  , \EAX_reg[17]/NET0131  , \EAX_reg[18]/NET0131  , \EAX_reg[19]/NET0131  , \EAX_reg[1]/NET0131  , \EAX_reg[20]/NET0131  , \EAX_reg[21]/NET0131  , \EAX_reg[22]/NET0131  , \EAX_reg[23]/NET0131  , \EAX_reg[24]/NET0131  , \EAX_reg[25]/NET0131  , \EAX_reg[26]/NET0131  , \EAX_reg[27]/NET0131  , \EAX_reg[28]/NET0131  , \EAX_reg[29]/NET0131  , \EAX_reg[2]/NET0131  , \EAX_reg[30]/NET0131  , \EAX_reg[31]/NET0131  , \EAX_reg[3]/NET0131  , \EAX_reg[4]/NET0131  , \EAX_reg[5]/NET0131  , \EAX_reg[6]/NET0131  , \EAX_reg[7]/NET0131  , \EAX_reg[8]/NET0131  , \EAX_reg[9]/NET0131  , \EBX_reg[0]/NET0131  , \EBX_reg[10]/NET0131  , \EBX_reg[11]/NET0131  , \EBX_reg[12]/NET0131  , \EBX_reg[13]/NET0131  , \EBX_reg[14]/NET0131  , \EBX_reg[15]/NET0131  , \EBX_reg[16]/NET0131  , \EBX_reg[17]/NET0131  , \EBX_reg[18]/NET0131  , \EBX_reg[19]/NET0131  , \EBX_reg[1]/NET0131  , \EBX_reg[20]/NET0131  , \EBX_reg[21]/NET0131  , \EBX_reg[22]/NET0131  , \EBX_reg[23]/NET0131  , \EBX_reg[24]/NET0131  , \EBX_reg[25]/NET0131  , \EBX_reg[26]/NET0131  , \EBX_reg[27]/NET0131  , \EBX_reg[28]/NET0131  , \EBX_reg[29]/NET0131  , \EBX_reg[2]/NET0131  , \EBX_reg[30]/NET0131  , \EBX_reg[31]/NET0131  , \EBX_reg[3]/NET0131  , \EBX_reg[4]/NET0131  , \EBX_reg[5]/NET0131  , \EBX_reg[6]/NET0131  , \EBX_reg[7]/NET0131  , \EBX_reg[8]/NET0131  , \EBX_reg[9]/NET0131  , \Flush_reg/NET0131  , HOLD_pad , \InstAddrPointer_reg[0]/NET0131  , \InstAddrPointer_reg[10]/NET0131  , \InstAddrPointer_reg[11]/NET0131  , \InstAddrPointer_reg[12]/NET0131  , \InstAddrPointer_reg[13]/NET0131  , \InstAddrPointer_reg[14]/NET0131  , \InstAddrPointer_reg[15]/NET0131  , \InstAddrPointer_reg[16]/NET0131  , \InstAddrPointer_reg[17]/NET0131  , \InstAddrPointer_reg[18]/NET0131  , \InstAddrPointer_reg[19]/NET0131  , \InstAddrPointer_reg[1]/NET0131  , \InstAddrPointer_reg[20]/NET0131  , \InstAddrPointer_reg[21]/NET0131  , \InstAddrPointer_reg[22]/NET0131  , \InstAddrPointer_reg[23]/NET0131  , \InstAddrPointer_reg[24]/NET0131  , \InstAddrPointer_reg[25]/NET0131  , \InstAddrPointer_reg[26]/NET0131  , \InstAddrPointer_reg[27]/NET0131  , \InstAddrPointer_reg[28]/NET0131  , \InstAddrPointer_reg[29]/NET0131  , \InstAddrPointer_reg[2]/NET0131  , \InstAddrPointer_reg[30]/NET0131  , \InstAddrPointer_reg[31]/NET0131  , \InstAddrPointer_reg[3]/NET0131  , \InstAddrPointer_reg[4]/NET0131  , \InstAddrPointer_reg[5]/NET0131  , \InstAddrPointer_reg[6]/NET0131  , \InstAddrPointer_reg[7]/NET0131  , \InstAddrPointer_reg[8]/NET0131  , \InstAddrPointer_reg[9]/NET0131  , \InstQueueRd_Addr_reg[0]/NET0131  , \InstQueueRd_Addr_reg[1]/NET0131  , \InstQueueRd_Addr_reg[2]/NET0131  , \InstQueueRd_Addr_reg[3]/NET0131  , \InstQueueWr_Addr_reg[0]/NET0131  , \InstQueueWr_Addr_reg[1]/NET0131  , \InstQueueWr_Addr_reg[2]/NET0131  , \InstQueueWr_Addr_reg[3]/NET0131  , \InstQueue_reg[0][0]/NET0131  , \InstQueue_reg[0][1]/NET0131  , \InstQueue_reg[0][2]/NET0131  , \InstQueue_reg[0][3]/NET0131  , \InstQueue_reg[0][4]/NET0131  , \InstQueue_reg[0][5]/NET0131  , \InstQueue_reg[0][6]/NET0131  , \InstQueue_reg[0][7]/NET0131  , \InstQueue_reg[10][0]/NET0131  , \InstQueue_reg[10][1]/NET0131  , \InstQueue_reg[10][2]/NET0131  , \InstQueue_reg[10][3]/NET0131  , \InstQueue_reg[10][4]/NET0131  , \InstQueue_reg[10][5]/NET0131  , \InstQueue_reg[10][6]/NET0131  , \InstQueue_reg[10][7]/NET0131  , \InstQueue_reg[11][0]/NET0131  , \InstQueue_reg[11][1]/NET0131  , \InstQueue_reg[11][2]/NET0131  , \InstQueue_reg[11][3]/NET0131  , \InstQueue_reg[11][4]/NET0131  , \InstQueue_reg[11][5]/NET0131  , \InstQueue_reg[11][6]/NET0131  , \InstQueue_reg[11][7]/NET0131  , \InstQueue_reg[12][0]/NET0131  , \InstQueue_reg[12][1]/NET0131  , \InstQueue_reg[12][2]/NET0131  , \InstQueue_reg[12][3]/NET0131  , \InstQueue_reg[12][4]/NET0131  , \InstQueue_reg[12][5]/NET0131  , \InstQueue_reg[12][6]/NET0131  , \InstQueue_reg[12][7]/NET0131  , \InstQueue_reg[13][0]/NET0131  , \InstQueue_reg[13][1]/NET0131  , \InstQueue_reg[13][2]/NET0131  , \InstQueue_reg[13][3]/NET0131  , \InstQueue_reg[13][4]/NET0131  , \InstQueue_reg[13][5]/NET0131  , \InstQueue_reg[13][6]/NET0131  , \InstQueue_reg[13][7]/NET0131  , \InstQueue_reg[14][0]/NET0131  , \InstQueue_reg[14][1]/NET0131  , \InstQueue_reg[14][2]/NET0131  , \InstQueue_reg[14][3]/NET0131  , \InstQueue_reg[14][4]/NET0131  , \InstQueue_reg[14][5]/NET0131  , \InstQueue_reg[14][6]/NET0131  , \InstQueue_reg[14][7]/NET0131  , \InstQueue_reg[15][0]/NET0131  , \InstQueue_reg[15][1]/NET0131  , \InstQueue_reg[15][2]/NET0131  , \InstQueue_reg[15][3]/NET0131  , \InstQueue_reg[15][4]/NET0131  , \InstQueue_reg[15][5]/NET0131  , \InstQueue_reg[15][6]/NET0131  , \InstQueue_reg[15][7]/NET0131  , \InstQueue_reg[1][0]/NET0131  , \InstQueue_reg[1][1]/NET0131  , \InstQueue_reg[1][2]/NET0131  , \InstQueue_reg[1][3]/NET0131  , \InstQueue_reg[1][4]/NET0131  , \InstQueue_reg[1][5]/NET0131  , \InstQueue_reg[1][6]/NET0131  , \InstQueue_reg[1][7]/NET0131  , \InstQueue_reg[2][0]/NET0131  , \InstQueue_reg[2][1]/NET0131  , \InstQueue_reg[2][2]/NET0131  , \InstQueue_reg[2][3]/NET0131  , \InstQueue_reg[2][4]/NET0131  , \InstQueue_reg[2][5]/NET0131  , \InstQueue_reg[2][6]/NET0131  , \InstQueue_reg[2][7]/NET0131  , \InstQueue_reg[3][0]/NET0131  , \InstQueue_reg[3][1]/NET0131  , \InstQueue_reg[3][2]/NET0131  , \InstQueue_reg[3][3]/NET0131  , \InstQueue_reg[3][4]/NET0131  , \InstQueue_reg[3][5]/NET0131  , \InstQueue_reg[3][6]/NET0131  , \InstQueue_reg[3][7]/NET0131  , \InstQueue_reg[4][0]/NET0131  , \InstQueue_reg[4][1]/NET0131  , \InstQueue_reg[4][2]/NET0131  , \InstQueue_reg[4][3]/NET0131  , \InstQueue_reg[4][4]/NET0131  , \InstQueue_reg[4][5]/NET0131  , \InstQueue_reg[4][6]/NET0131  , \InstQueue_reg[4][7]/NET0131  , \InstQueue_reg[5][0]/NET0131  , \InstQueue_reg[5][1]/NET0131  , \InstQueue_reg[5][2]/NET0131  , \InstQueue_reg[5][3]/NET0131  , \InstQueue_reg[5][4]/NET0131  , \InstQueue_reg[5][5]/NET0131  , \InstQueue_reg[5][6]/NET0131  , \InstQueue_reg[5][7]/NET0131  , \InstQueue_reg[6][0]/NET0131  , \InstQueue_reg[6][1]/NET0131  , \InstQueue_reg[6][2]/NET0131  , \InstQueue_reg[6][3]/NET0131  , \InstQueue_reg[6][4]/NET0131  , \InstQueue_reg[6][5]/NET0131  , \InstQueue_reg[6][6]/NET0131  , \InstQueue_reg[6][7]/NET0131  , \InstQueue_reg[7][0]/NET0131  , \InstQueue_reg[7][1]/NET0131  , \InstQueue_reg[7][2]/NET0131  , \InstQueue_reg[7][3]/NET0131  , \InstQueue_reg[7][4]/NET0131  , \InstQueue_reg[7][5]/NET0131  , \InstQueue_reg[7][6]/NET0131  , \InstQueue_reg[7][7]/NET0131  , \InstQueue_reg[8][0]/NET0131  , \InstQueue_reg[8][1]/NET0131  , \InstQueue_reg[8][2]/NET0131  , \InstQueue_reg[8][3]/NET0131  , \InstQueue_reg[8][4]/NET0131  , \InstQueue_reg[8][5]/NET0131  , \InstQueue_reg[8][6]/NET0131  , \InstQueue_reg[8][7]/NET0131  , \InstQueue_reg[9][0]/NET0131  , \InstQueue_reg[9][1]/NET0131  , \InstQueue_reg[9][2]/NET0131  , \InstQueue_reg[9][3]/NET0131  , \InstQueue_reg[9][4]/NET0131  , \InstQueue_reg[9][5]/NET0131  , \InstQueue_reg[9][6]/NET0131  , \InstQueue_reg[9][7]/NET0131  , M_IO_n_pad , \MemoryFetch_reg/NET0131  , \More_reg/NET0131  , NA_n_pad , \PhyAddrPointer_reg[0]/NET0131  , \PhyAddrPointer_reg[10]/NET0131  , \PhyAddrPointer_reg[11]/NET0131  , \PhyAddrPointer_reg[12]/NET0131  , \PhyAddrPointer_reg[13]/NET0131  , \PhyAddrPointer_reg[14]/NET0131  , \PhyAddrPointer_reg[15]/NET0131  , \PhyAddrPointer_reg[16]/NET0131  , \PhyAddrPointer_reg[17]/NET0131  , \PhyAddrPointer_reg[18]/NET0131  , \PhyAddrPointer_reg[19]/NET0131  , \PhyAddrPointer_reg[1]/NET0131  , \PhyAddrPointer_reg[20]/NET0131  , \PhyAddrPointer_reg[21]/NET0131  , \PhyAddrPointer_reg[22]/NET0131  , \PhyAddrPointer_reg[23]/NET0131  , \PhyAddrPointer_reg[24]/NET0131  , \PhyAddrPointer_reg[25]/NET0131  , \PhyAddrPointer_reg[26]/NET0131  , \PhyAddrPointer_reg[27]/NET0131  , \PhyAddrPointer_reg[28]/NET0131  , \PhyAddrPointer_reg[29]/NET0131  , \PhyAddrPointer_reg[2]/NET0131  , \PhyAddrPointer_reg[30]/NET0131  , \PhyAddrPointer_reg[31]/NET0131  , \PhyAddrPointer_reg[3]/NET0131  , \PhyAddrPointer_reg[4]/NET0131  , \PhyAddrPointer_reg[5]/NET0131  , \PhyAddrPointer_reg[6]/NET0131  , \PhyAddrPointer_reg[7]/NET0131  , \PhyAddrPointer_reg[8]/NET0131  , \PhyAddrPointer_reg[9]/NET0131  , READY_n_pad , \ReadRequest_reg/NET0131  , \RequestPending_reg/NET0131  , \State2_reg[0]/NET0131  , \State2_reg[1]/NET0131  , \State2_reg[2]/NET0131  , \State2_reg[3]/NET0131  , \State_reg[0]/NET0131  , \State_reg[1]/NET0131  , \State_reg[2]/NET0131  , W_R_n_pad , \lWord_reg[0]/NET0131  , \lWord_reg[10]/NET0131  , \lWord_reg[11]/NET0131  , \lWord_reg[12]/NET0131  , \lWord_reg[13]/NET0131  , \lWord_reg[14]/NET0131  , \lWord_reg[15]/NET0131  , \lWord_reg[1]/NET0131  , \lWord_reg[2]/NET0131  , \lWord_reg[3]/NET0131  , \lWord_reg[4]/NET0131  , \lWord_reg[5]/NET0131  , \lWord_reg[6]/NET0131  , \lWord_reg[7]/NET0131  , \lWord_reg[8]/NET0131  , \lWord_reg[9]/NET0131  , \rEIP_reg[0]/NET0131  , \rEIP_reg[10]/NET0131  , \rEIP_reg[11]/NET0131  , \rEIP_reg[12]/NET0131  , \rEIP_reg[13]/NET0131  , \rEIP_reg[14]/NET0131  , \rEIP_reg[15]/NET0131  , \rEIP_reg[16]/NET0131  , \rEIP_reg[17]/NET0131  , \rEIP_reg[18]/NET0131  , \rEIP_reg[19]/NET0131  , \rEIP_reg[1]/NET0131  , \rEIP_reg[20]/NET0131  , \rEIP_reg[21]/NET0131  , \rEIP_reg[22]/NET0131  , \rEIP_reg[23]/NET0131  , \rEIP_reg[24]/NET0131  , \rEIP_reg[25]/NET0131  , \rEIP_reg[26]/NET0131  , \rEIP_reg[27]/NET0131  , \rEIP_reg[28]/NET0131  , \rEIP_reg[29]/NET0131  , \rEIP_reg[2]/NET0131  , \rEIP_reg[30]/NET0131  , \rEIP_reg[31]/NET0131  , \rEIP_reg[3]/NET0131  , \rEIP_reg[4]/NET0131  , \rEIP_reg[5]/NET0131  , \rEIP_reg[6]/NET0131  , \rEIP_reg[7]/NET0131  , \rEIP_reg[8]/NET0131  , \rEIP_reg[9]/NET0131  , \uWord_reg[0]/NET0131  , \uWord_reg[10]/NET0131  , \uWord_reg[11]/NET0131  , \uWord_reg[12]/NET0131  , \uWord_reg[13]/NET0131  , \uWord_reg[14]/NET0131  , \uWord_reg[1]/NET0131  , \uWord_reg[2]/NET0131  , \uWord_reg[3]/NET0131  , \uWord_reg[4]/NET0131  , \uWord_reg[5]/NET0131  , \uWord_reg[6]/NET0131  , \uWord_reg[7]/NET0131  , \uWord_reg[8]/NET0131  , \uWord_reg[9]/NET0131  , \_al_n0  , \_al_n1  , \g47521/_2_  , \g47523/_0_  , \g47526/_0_  , \g47529/_0_  , \g47533/_0_  , \g47540/_0_  , \g47551/_0_  , \g47552/_0_  , \g47553/_0_  , \g47563/_2_  , \g47566/_0_  , \g47567/_0_  , \g47568/_0_  , \g47569/_0_  , \g47583/_2_  , \g47584/_0_  , \g47585/_0_  , \g47589/_0_  , \g47602/_0_  , \g47603/_0_  , \g47604/_2_  , \g47605/_0_  , \g47606/_2_  , \g47609/_0_  , \g47611/_0_  , \g47631/_0_  , \g47632/_0_  , \g47633/_0_  , \g47635/_0_  , \g47636/_0_  , \g47637/_0_  , \g47638/_2_  , \g47643/_0_  , \g47665/_2_  , \g47666/_0_  , \g47667/_0_  , \g47670/_0_  , \g47672/_0_  , \g47677/_0_  , \g47678/_0_  , \g47706/_0_  , \g47711/_0_  , \g47717/_0_  , \g47718/_0_  , \g47721/_0_  , \g47722/_0_  , \g47751/_0_  , \g47755/_0_  , \g47756/_0_  , \g47757/_0_  , \g47759/_0_  , \g47789/_0_  , \g47793/_0_  , \g47797/_0_  , \g47798/_0_  , \g47799/_0_  , \g47802/_0_  , \g47804/_0_  , \g47807/_0_  , \g47809/_0_  , \g47862/_0_  , \g47863/_0_  , \g47864/_0_  , \g47869/_0_  , \g47870/_0_  , \g47924/_0_  , \g47925/_0_  , \g47926/_0_  , \g47927/_0_  , \g47928/_0_  , \g47930/_0_  , \g47932/_0_  , \g47933/_0_  , \g47934/_0_  , \g47935/_0_  , \g47936/_0_  , \g47937/_0_  , \g47938/_0_  , \g47939/_0_  , \g47940/_0_  , \g47941/_0_  , \g47957/_0_  , \g47970/_0_  , \g47973/_0_  , \g47975/_0_  , \g48058/_0_  , \g48059/_0_  , \g48060/_0_  , \g48061/_0_  , \g48062/_0_  , \g48064/_0_  , \g48065/_0_  , \g48066/_0_  , \g48067/_0_  , \g48068/_0_  , \g48069/_0_  , \g48070/_0_  , \g48071/_0_  , \g48072/_0_  , \g48073/_0_  , \g48074/_0_  , \g48087/_0_  , \g48110/_0_  , \g48117/_0_  , \g48118/_0_  , \g48119/_0_  , \g48120/_0_  , \g48121/_0_  , \g48122/_0_  , \g48124/_0_  , \g48125/_0_  , \g48126/_0_  , \g48127/_0_  , \g48128/_0_  , \g48129/_0_  , \g48130/_0_  , \g48131/_0_  , \g48132/_0_  , \g48133/_0_  , \g48134/_0_  , \g48168/_0_  , \g48169/_0_  , \g48170/_0_  , \g48171/_0_  , \g48172/_0_  , \g48173/_0_  , \g48174/_0_  , \g48175/_0_  , \g48177/_0_  , \g48178/_0_  , \g48179/_0_  , \g48180/_0_  , \g48181/_0_  , \g48182/_0_  , \g48183/_0_  , \g48184/_0_  , \g48185/_0_  , \g48186/_0_  , \g48187/_0_  , \g48188/_0_  , \g48189/_0_  , \g48192/_0_  , \g48193/_0_  , \g48194/_0_  , \g48195/_0_  , \g48196/_0_  , \g48197/_0_  , \g48198/_0_  , \g48199/_0_  , \g48200/_0_  , \g48201/_0_  , \g48202/_0_  , \g48203/_0_  , \g48213/_0_  , \g48214/_0_  , \g48215/_0_  , \g48216/_0_  , \g48217/_0_  , \g48218/_0_  , \g48219/_0_  , \g48220/_0_  , \g48221/_0_  , \g48222/_0_  , \g48223/_0_  , \g48224/_0_  , \g48225/_0_  , \g48226/_0_  , \g48227/_0_  , \g48228/_0_  , \g48229/_0_  , \g48230/_0_  , \g48231/_0_  , \g48232/_0_  , \g48234/_0_  , \g48236/_0_  , \g48237/_0_  , \g48238/_0_  , \g48239/_0_  , \g48240/_0_  , \g48241/_0_  , \g48243/_0_  , \g48244/_0_  , \g48245/_0_  , \g48246/_0_  , \g48263/_0_  , \g48270/_0_  , \g48273/_0_  , \g48276/_0_  , \g48277/_0_  , \g48370/_0_  , \g48377/_0_  , \g48391/_0_  , \g48423/_0_  , \g48428/_0_  , \g48429/_0_  , \g48431/_0_  , \g48433/_0_  , \g48434/_0_  , \g48435/_0_  , \g48436/_0_  , \g48437/_0_  , \g48438/_0_  , \g48439/_0_  , \g48440/_0_  , \g48441/_0_  , \g48442/_0_  , \g48443/_0_  , \g48610/_0_  , \g48634/_0_  , \g48635/_0_  , \g48636/_0_  , \g48637/_0_  , \g48638/_0_  , \g48639/_0_  , \g48640/_0_  , \g48642/_0_  , \g48643/_0_  , \g48644/_0_  , \g48645/_0_  , \g48646/_0_  , \g48647/_0_  , \g48648/_0_  , \g48649/_0_  , \g48650/_0_  , \g48651/_0_  , \g48652/_0_  , \g48653/_0_  , \g48654/_0_  , \g48655/_0_  , \g48656/_0_  , \g48657/_0_  , \g48658/_0_  , \g48659/_0_  , \g48660/_0_  , \g48662/_0_  , \g48663/_0_  , \g48664/_0_  , \g48665/_0_  , \g48666/_0_  , \g48667/_0_  , \g48668/_0_  , \g48669/_0_  , \g48750/_0_  , \g48753/_0_  , \g48756/_0_  , \g48759/_0_  , \g48763/_0_  , \g48766/_0_  , \g48769/_0_  , \g48772/_0_  , \g48775/_0_  , \g48778/_0_  , \g48781/_0_  , \g48785/_0_  , \g48789/_0_  , \g48792/_0_  , \g48796/_0_  , \g48799/_0_  , \g48937/_0_  , \g48958/_0_  , \g48959/_0_  , \g48964/_0_  , \g48965/_0_  , \g48966/_0_  , \g48967/_0_  , \g48968/_0_  , \g48969/_0_  , \g48970/_0_  , \g48971/_0_  , \g48972/_0_  , \g48973/_0_  , \g48974/_0_  , \g48975/_0_  , \g48976/_0_  , \g48977/_0_  , \g48978/_0_  , \g48979/_0_  , \g49/_0_  , \g49069/_0_  , \g49070/_0_  , \g49071/_0_  , \g49073/_0_  , \g49074/_0_  , \g49076/_0_  , \g49078/_0_  , \g49081/_0_  , \g49083/_0_  , \g49085/_0_  , \g49087/_0_  , \g49088/_0_  , \g49090/_0_  , \g49092/_0_  , \g49095/_0_  , \g49098/_0_  , \g49125/_0_  , \g49162/_0_  , \g49202/_0_  , \g49203/_0_  , \g49206/_0_  , \g49340/_0_  , \g49457/_0_  , \g49512/_0_  , \g49513/_0_  , \g49514/_0_  , \g49515/_0_  , \g49516/_0_  , \g49517/_0_  , \g49518/_0_  , \g49519/_0_  , \g49520/_0_  , \g49521/_0_  , \g49522/_0_  , \g49523/_0_  , \g49524/_0_  , \g49525/_0_  , \g49526/_0_  , \g49527/_0_  , \g49534/_0_  , \g49551/_0_  , \g49573/_0_  , \g49574/_0_  , \g49578/_0_  , \g49582/_0_  , \g49584/_0_  , \g49592/_0_  , \g49600/_0_  , \g49604/_0_  , \g49608/_0_  , \g49612/_0_  , \g49616/_0_  , \g49619/_0_  , \g49620/_0_  , \g49623/_0_  , \g49627/_0_  , \g49630/_0_  , \g49634/_0_  , \g49635/_0_  , \g49639/_0_  , \g49645/_0_  , \g49744/_0_  , \g49766/_0_  , \g50098/_0_  , \g50124/_0_  , \g50195/_0_  , \g50198/_0_  , \g50201/_0_  , \g50203/_0_  , \g50205/_0_  , \g50207/_0_  , \g50209/_0_  , \g50213/_0_  , \g50222/_0_  , \g50228/_0_  , \g50231/_0_  , \g50237/_0_  , \g50240/_0_  , \g50335/_0_  , \g50477/_0_  , \g50478/_0_  , \g50671/_0_  , \g50757/_0_  , \g50938/_0_  , \g50998/_0_  , \g51008/_0_  , \g51579/_0_  , \g51637/_0_  , \g51662/_0_  , \g52424/_0_  , \g53184/_0_  , \g53206/_0_  , \g53270/_0_  , \g53730/_0_  , \g53754/_0_  , \g54176/_0_  , \g54214/_0_  , \g54229/_0_  , \g54392/_0_  , \g54400/_0_  , \g54415/_0_  , \g54421/_0_  , \g54604/_0_  , \g54607/_0_  , \g54638/_0_  , \g54694/_0_  , \g54759/_0_  , \g55607/_0_  , \g55863/_1_  , \g56073/_0_  , \g56292/_0_  , \g56320/_0_  , \g56527/_0_  , \g56531/_0_  , \g56533/_0_  , \g56562/_0_  , \g56615/_0_  , \g56720/_0_  , \g57044/_0_  , \g60635/_1_  , \g62873/_0_  , \g62886/_0_  , \g63001/_0_  , \g63101/_0_  , \g63129/_0_  , \g63198/_0_  , \g63449/_0_  , \g63471/_0_  , \g63493/_0_  , \g63626/_0_  , \g63688/_0_  , \g63800/_0_  , \g63934/_0_  , \g63954/_0_  , \g64060/_0_  , \g64375/_0_  , \g65/_0_  , \g67/_0_  );
  input ADS_n_pad ;
  input \Address[0]_pad  ;
  input \Address[10]_pad  ;
  input \Address[11]_pad  ;
  input \Address[12]_pad  ;
  input \Address[13]_pad  ;
  input \Address[14]_pad  ;
  input \Address[15]_pad  ;
  input \Address[16]_pad  ;
  input \Address[17]_pad  ;
  input \Address[18]_pad  ;
  input \Address[19]_pad  ;
  input \Address[1]_pad  ;
  input \Address[20]_pad  ;
  input \Address[21]_pad  ;
  input \Address[22]_pad  ;
  input \Address[23]_pad  ;
  input \Address[24]_pad  ;
  input \Address[25]_pad  ;
  input \Address[26]_pad  ;
  input \Address[27]_pad  ;
  input \Address[28]_pad  ;
  input \Address[29]_pad  ;
  input \Address[2]_pad  ;
  input \Address[3]_pad  ;
  input \Address[4]_pad  ;
  input \Address[5]_pad  ;
  input \Address[6]_pad  ;
  input \Address[7]_pad  ;
  input \Address[8]_pad  ;
  input \Address[9]_pad  ;
  input \BE_n[0]_pad  ;
  input \BE_n[1]_pad  ;
  input \BE_n[2]_pad  ;
  input \BE_n[3]_pad  ;
  input \BS16_n_pad  ;
  input \ByteEnable_reg[0]/NET0131  ;
  input \ByteEnable_reg[1]/NET0131  ;
  input \ByteEnable_reg[2]/NET0131  ;
  input \ByteEnable_reg[3]/NET0131  ;
  input \CodeFetch_reg/NET0131  ;
  input D_C_n_pad ;
  input \DataWidth_reg[0]/NET0131  ;
  input \DataWidth_reg[1]/NET0131  ;
  input \Datai[0]_pad  ;
  input \Datai[10]_pad  ;
  input \Datai[11]_pad  ;
  input \Datai[12]_pad  ;
  input \Datai[13]_pad  ;
  input \Datai[14]_pad  ;
  input \Datai[15]_pad  ;
  input \Datai[16]_pad  ;
  input \Datai[17]_pad  ;
  input \Datai[18]_pad  ;
  input \Datai[19]_pad  ;
  input \Datai[1]_pad  ;
  input \Datai[20]_pad  ;
  input \Datai[21]_pad  ;
  input \Datai[22]_pad  ;
  input \Datai[23]_pad  ;
  input \Datai[24]_pad  ;
  input \Datai[25]_pad  ;
  input \Datai[26]_pad  ;
  input \Datai[27]_pad  ;
  input \Datai[28]_pad  ;
  input \Datai[29]_pad  ;
  input \Datai[2]_pad  ;
  input \Datai[30]_pad  ;
  input \Datai[31]_pad  ;
  input \Datai[3]_pad  ;
  input \Datai[4]_pad  ;
  input \Datai[5]_pad  ;
  input \Datai[6]_pad  ;
  input \Datai[7]_pad  ;
  input \Datai[8]_pad  ;
  input \Datai[9]_pad  ;
  input \Datao[0]_pad  ;
  input \Datao[10]_pad  ;
  input \Datao[11]_pad  ;
  input \Datao[12]_pad  ;
  input \Datao[13]_pad  ;
  input \Datao[14]_pad  ;
  input \Datao[15]_pad  ;
  input \Datao[16]_pad  ;
  input \Datao[17]_pad  ;
  input \Datao[18]_pad  ;
  input \Datao[19]_pad  ;
  input \Datao[1]_pad  ;
  input \Datao[20]_pad  ;
  input \Datao[21]_pad  ;
  input \Datao[23]_pad  ;
  input \Datao[24]_pad  ;
  input \Datao[25]_pad  ;
  input \Datao[26]_pad  ;
  input \Datao[27]_pad  ;
  input \Datao[28]_pad  ;
  input \Datao[29]_pad  ;
  input \Datao[2]_pad  ;
  input \Datao[30]_pad  ;
  input \Datao[3]_pad  ;
  input \Datao[4]_pad  ;
  input \Datao[5]_pad  ;
  input \Datao[6]_pad  ;
  input \Datao[7]_pad  ;
  input \Datao[8]_pad  ;
  input \Datao[9]_pad  ;
  input \Datao_reg[22]/NET0131  ;
  input \EAX_reg[0]/NET0131  ;
  input \EAX_reg[10]/NET0131  ;
  input \EAX_reg[11]/NET0131  ;
  input \EAX_reg[12]/NET0131  ;
  input \EAX_reg[13]/NET0131  ;
  input \EAX_reg[14]/NET0131  ;
  input \EAX_reg[15]/NET0131  ;
  input \EAX_reg[16]/NET0131  ;
  input \EAX_reg[17]/NET0131  ;
  input \EAX_reg[18]/NET0131  ;
  input \EAX_reg[19]/NET0131  ;
  input \EAX_reg[1]/NET0131  ;
  input \EAX_reg[20]/NET0131  ;
  input \EAX_reg[21]/NET0131  ;
  input \EAX_reg[22]/NET0131  ;
  input \EAX_reg[23]/NET0131  ;
  input \EAX_reg[24]/NET0131  ;
  input \EAX_reg[25]/NET0131  ;
  input \EAX_reg[26]/NET0131  ;
  input \EAX_reg[27]/NET0131  ;
  input \EAX_reg[28]/NET0131  ;
  input \EAX_reg[29]/NET0131  ;
  input \EAX_reg[2]/NET0131  ;
  input \EAX_reg[30]/NET0131  ;
  input \EAX_reg[31]/NET0131  ;
  input \EAX_reg[3]/NET0131  ;
  input \EAX_reg[4]/NET0131  ;
  input \EAX_reg[5]/NET0131  ;
  input \EAX_reg[6]/NET0131  ;
  input \EAX_reg[7]/NET0131  ;
  input \EAX_reg[8]/NET0131  ;
  input \EAX_reg[9]/NET0131  ;
  input \EBX_reg[0]/NET0131  ;
  input \EBX_reg[10]/NET0131  ;
  input \EBX_reg[11]/NET0131  ;
  input \EBX_reg[12]/NET0131  ;
  input \EBX_reg[13]/NET0131  ;
  input \EBX_reg[14]/NET0131  ;
  input \EBX_reg[15]/NET0131  ;
  input \EBX_reg[16]/NET0131  ;
  input \EBX_reg[17]/NET0131  ;
  input \EBX_reg[18]/NET0131  ;
  input \EBX_reg[19]/NET0131  ;
  input \EBX_reg[1]/NET0131  ;
  input \EBX_reg[20]/NET0131  ;
  input \EBX_reg[21]/NET0131  ;
  input \EBX_reg[22]/NET0131  ;
  input \EBX_reg[23]/NET0131  ;
  input \EBX_reg[24]/NET0131  ;
  input \EBX_reg[25]/NET0131  ;
  input \EBX_reg[26]/NET0131  ;
  input \EBX_reg[27]/NET0131  ;
  input \EBX_reg[28]/NET0131  ;
  input \EBX_reg[29]/NET0131  ;
  input \EBX_reg[2]/NET0131  ;
  input \EBX_reg[30]/NET0131  ;
  input \EBX_reg[31]/NET0131  ;
  input \EBX_reg[3]/NET0131  ;
  input \EBX_reg[4]/NET0131  ;
  input \EBX_reg[5]/NET0131  ;
  input \EBX_reg[6]/NET0131  ;
  input \EBX_reg[7]/NET0131  ;
  input \EBX_reg[8]/NET0131  ;
  input \EBX_reg[9]/NET0131  ;
  input \Flush_reg/NET0131  ;
  input HOLD_pad ;
  input \InstAddrPointer_reg[0]/NET0131  ;
  input \InstAddrPointer_reg[10]/NET0131  ;
  input \InstAddrPointer_reg[11]/NET0131  ;
  input \InstAddrPointer_reg[12]/NET0131  ;
  input \InstAddrPointer_reg[13]/NET0131  ;
  input \InstAddrPointer_reg[14]/NET0131  ;
  input \InstAddrPointer_reg[15]/NET0131  ;
  input \InstAddrPointer_reg[16]/NET0131  ;
  input \InstAddrPointer_reg[17]/NET0131  ;
  input \InstAddrPointer_reg[18]/NET0131  ;
  input \InstAddrPointer_reg[19]/NET0131  ;
  input \InstAddrPointer_reg[1]/NET0131  ;
  input \InstAddrPointer_reg[20]/NET0131  ;
  input \InstAddrPointer_reg[21]/NET0131  ;
  input \InstAddrPointer_reg[22]/NET0131  ;
  input \InstAddrPointer_reg[23]/NET0131  ;
  input \InstAddrPointer_reg[24]/NET0131  ;
  input \InstAddrPointer_reg[25]/NET0131  ;
  input \InstAddrPointer_reg[26]/NET0131  ;
  input \InstAddrPointer_reg[27]/NET0131  ;
  input \InstAddrPointer_reg[28]/NET0131  ;
  input \InstAddrPointer_reg[29]/NET0131  ;
  input \InstAddrPointer_reg[2]/NET0131  ;
  input \InstAddrPointer_reg[30]/NET0131  ;
  input \InstAddrPointer_reg[31]/NET0131  ;
  input \InstAddrPointer_reg[3]/NET0131  ;
  input \InstAddrPointer_reg[4]/NET0131  ;
  input \InstAddrPointer_reg[5]/NET0131  ;
  input \InstAddrPointer_reg[6]/NET0131  ;
  input \InstAddrPointer_reg[7]/NET0131  ;
  input \InstAddrPointer_reg[8]/NET0131  ;
  input \InstAddrPointer_reg[9]/NET0131  ;
  input \InstQueueRd_Addr_reg[0]/NET0131  ;
  input \InstQueueRd_Addr_reg[1]/NET0131  ;
  input \InstQueueRd_Addr_reg[2]/NET0131  ;
  input \InstQueueRd_Addr_reg[3]/NET0131  ;
  input \InstQueueWr_Addr_reg[0]/NET0131  ;
  input \InstQueueWr_Addr_reg[1]/NET0131  ;
  input \InstQueueWr_Addr_reg[2]/NET0131  ;
  input \InstQueueWr_Addr_reg[3]/NET0131  ;
  input \InstQueue_reg[0][0]/NET0131  ;
  input \InstQueue_reg[0][1]/NET0131  ;
  input \InstQueue_reg[0][2]/NET0131  ;
  input \InstQueue_reg[0][3]/NET0131  ;
  input \InstQueue_reg[0][4]/NET0131  ;
  input \InstQueue_reg[0][5]/NET0131  ;
  input \InstQueue_reg[0][6]/NET0131  ;
  input \InstQueue_reg[0][7]/NET0131  ;
  input \InstQueue_reg[10][0]/NET0131  ;
  input \InstQueue_reg[10][1]/NET0131  ;
  input \InstQueue_reg[10][2]/NET0131  ;
  input \InstQueue_reg[10][3]/NET0131  ;
  input \InstQueue_reg[10][4]/NET0131  ;
  input \InstQueue_reg[10][5]/NET0131  ;
  input \InstQueue_reg[10][6]/NET0131  ;
  input \InstQueue_reg[10][7]/NET0131  ;
  input \InstQueue_reg[11][0]/NET0131  ;
  input \InstQueue_reg[11][1]/NET0131  ;
  input \InstQueue_reg[11][2]/NET0131  ;
  input \InstQueue_reg[11][3]/NET0131  ;
  input \InstQueue_reg[11][4]/NET0131  ;
  input \InstQueue_reg[11][5]/NET0131  ;
  input \InstQueue_reg[11][6]/NET0131  ;
  input \InstQueue_reg[11][7]/NET0131  ;
  input \InstQueue_reg[12][0]/NET0131  ;
  input \InstQueue_reg[12][1]/NET0131  ;
  input \InstQueue_reg[12][2]/NET0131  ;
  input \InstQueue_reg[12][3]/NET0131  ;
  input \InstQueue_reg[12][4]/NET0131  ;
  input \InstQueue_reg[12][5]/NET0131  ;
  input \InstQueue_reg[12][6]/NET0131  ;
  input \InstQueue_reg[12][7]/NET0131  ;
  input \InstQueue_reg[13][0]/NET0131  ;
  input \InstQueue_reg[13][1]/NET0131  ;
  input \InstQueue_reg[13][2]/NET0131  ;
  input \InstQueue_reg[13][3]/NET0131  ;
  input \InstQueue_reg[13][4]/NET0131  ;
  input \InstQueue_reg[13][5]/NET0131  ;
  input \InstQueue_reg[13][6]/NET0131  ;
  input \InstQueue_reg[13][7]/NET0131  ;
  input \InstQueue_reg[14][0]/NET0131  ;
  input \InstQueue_reg[14][1]/NET0131  ;
  input \InstQueue_reg[14][2]/NET0131  ;
  input \InstQueue_reg[14][3]/NET0131  ;
  input \InstQueue_reg[14][4]/NET0131  ;
  input \InstQueue_reg[14][5]/NET0131  ;
  input \InstQueue_reg[14][6]/NET0131  ;
  input \InstQueue_reg[14][7]/NET0131  ;
  input \InstQueue_reg[15][0]/NET0131  ;
  input \InstQueue_reg[15][1]/NET0131  ;
  input \InstQueue_reg[15][2]/NET0131  ;
  input \InstQueue_reg[15][3]/NET0131  ;
  input \InstQueue_reg[15][4]/NET0131  ;
  input \InstQueue_reg[15][5]/NET0131  ;
  input \InstQueue_reg[15][6]/NET0131  ;
  input \InstQueue_reg[15][7]/NET0131  ;
  input \InstQueue_reg[1][0]/NET0131  ;
  input \InstQueue_reg[1][1]/NET0131  ;
  input \InstQueue_reg[1][2]/NET0131  ;
  input \InstQueue_reg[1][3]/NET0131  ;
  input \InstQueue_reg[1][4]/NET0131  ;
  input \InstQueue_reg[1][5]/NET0131  ;
  input \InstQueue_reg[1][6]/NET0131  ;
  input \InstQueue_reg[1][7]/NET0131  ;
  input \InstQueue_reg[2][0]/NET0131  ;
  input \InstQueue_reg[2][1]/NET0131  ;
  input \InstQueue_reg[2][2]/NET0131  ;
  input \InstQueue_reg[2][3]/NET0131  ;
  input \InstQueue_reg[2][4]/NET0131  ;
  input \InstQueue_reg[2][5]/NET0131  ;
  input \InstQueue_reg[2][6]/NET0131  ;
  input \InstQueue_reg[2][7]/NET0131  ;
  input \InstQueue_reg[3][0]/NET0131  ;
  input \InstQueue_reg[3][1]/NET0131  ;
  input \InstQueue_reg[3][2]/NET0131  ;
  input \InstQueue_reg[3][3]/NET0131  ;
  input \InstQueue_reg[3][4]/NET0131  ;
  input \InstQueue_reg[3][5]/NET0131  ;
  input \InstQueue_reg[3][6]/NET0131  ;
  input \InstQueue_reg[3][7]/NET0131  ;
  input \InstQueue_reg[4][0]/NET0131  ;
  input \InstQueue_reg[4][1]/NET0131  ;
  input \InstQueue_reg[4][2]/NET0131  ;
  input \InstQueue_reg[4][3]/NET0131  ;
  input \InstQueue_reg[4][4]/NET0131  ;
  input \InstQueue_reg[4][5]/NET0131  ;
  input \InstQueue_reg[4][6]/NET0131  ;
  input \InstQueue_reg[4][7]/NET0131  ;
  input \InstQueue_reg[5][0]/NET0131  ;
  input \InstQueue_reg[5][1]/NET0131  ;
  input \InstQueue_reg[5][2]/NET0131  ;
  input \InstQueue_reg[5][3]/NET0131  ;
  input \InstQueue_reg[5][4]/NET0131  ;
  input \InstQueue_reg[5][5]/NET0131  ;
  input \InstQueue_reg[5][6]/NET0131  ;
  input \InstQueue_reg[5][7]/NET0131  ;
  input \InstQueue_reg[6][0]/NET0131  ;
  input \InstQueue_reg[6][1]/NET0131  ;
  input \InstQueue_reg[6][2]/NET0131  ;
  input \InstQueue_reg[6][3]/NET0131  ;
  input \InstQueue_reg[6][4]/NET0131  ;
  input \InstQueue_reg[6][5]/NET0131  ;
  input \InstQueue_reg[6][6]/NET0131  ;
  input \InstQueue_reg[6][7]/NET0131  ;
  input \InstQueue_reg[7][0]/NET0131  ;
  input \InstQueue_reg[7][1]/NET0131  ;
  input \InstQueue_reg[7][2]/NET0131  ;
  input \InstQueue_reg[7][3]/NET0131  ;
  input \InstQueue_reg[7][4]/NET0131  ;
  input \InstQueue_reg[7][5]/NET0131  ;
  input \InstQueue_reg[7][6]/NET0131  ;
  input \InstQueue_reg[7][7]/NET0131  ;
  input \InstQueue_reg[8][0]/NET0131  ;
  input \InstQueue_reg[8][1]/NET0131  ;
  input \InstQueue_reg[8][2]/NET0131  ;
  input \InstQueue_reg[8][3]/NET0131  ;
  input \InstQueue_reg[8][4]/NET0131  ;
  input \InstQueue_reg[8][5]/NET0131  ;
  input \InstQueue_reg[8][6]/NET0131  ;
  input \InstQueue_reg[8][7]/NET0131  ;
  input \InstQueue_reg[9][0]/NET0131  ;
  input \InstQueue_reg[9][1]/NET0131  ;
  input \InstQueue_reg[9][2]/NET0131  ;
  input \InstQueue_reg[9][3]/NET0131  ;
  input \InstQueue_reg[9][4]/NET0131  ;
  input \InstQueue_reg[9][5]/NET0131  ;
  input \InstQueue_reg[9][6]/NET0131  ;
  input \InstQueue_reg[9][7]/NET0131  ;
  input M_IO_n_pad ;
  input \MemoryFetch_reg/NET0131  ;
  input \More_reg/NET0131  ;
  input NA_n_pad ;
  input \PhyAddrPointer_reg[0]/NET0131  ;
  input \PhyAddrPointer_reg[10]/NET0131  ;
  input \PhyAddrPointer_reg[11]/NET0131  ;
  input \PhyAddrPointer_reg[12]/NET0131  ;
  input \PhyAddrPointer_reg[13]/NET0131  ;
  input \PhyAddrPointer_reg[14]/NET0131  ;
  input \PhyAddrPointer_reg[15]/NET0131  ;
  input \PhyAddrPointer_reg[16]/NET0131  ;
  input \PhyAddrPointer_reg[17]/NET0131  ;
  input \PhyAddrPointer_reg[18]/NET0131  ;
  input \PhyAddrPointer_reg[19]/NET0131  ;
  input \PhyAddrPointer_reg[1]/NET0131  ;
  input \PhyAddrPointer_reg[20]/NET0131  ;
  input \PhyAddrPointer_reg[21]/NET0131  ;
  input \PhyAddrPointer_reg[22]/NET0131  ;
  input \PhyAddrPointer_reg[23]/NET0131  ;
  input \PhyAddrPointer_reg[24]/NET0131  ;
  input \PhyAddrPointer_reg[25]/NET0131  ;
  input \PhyAddrPointer_reg[26]/NET0131  ;
  input \PhyAddrPointer_reg[27]/NET0131  ;
  input \PhyAddrPointer_reg[28]/NET0131  ;
  input \PhyAddrPointer_reg[29]/NET0131  ;
  input \PhyAddrPointer_reg[2]/NET0131  ;
  input \PhyAddrPointer_reg[30]/NET0131  ;
  input \PhyAddrPointer_reg[31]/NET0131  ;
  input \PhyAddrPointer_reg[3]/NET0131  ;
  input \PhyAddrPointer_reg[4]/NET0131  ;
  input \PhyAddrPointer_reg[5]/NET0131  ;
  input \PhyAddrPointer_reg[6]/NET0131  ;
  input \PhyAddrPointer_reg[7]/NET0131  ;
  input \PhyAddrPointer_reg[8]/NET0131  ;
  input \PhyAddrPointer_reg[9]/NET0131  ;
  input READY_n_pad ;
  input \ReadRequest_reg/NET0131  ;
  input \RequestPending_reg/NET0131  ;
  input \State2_reg[0]/NET0131  ;
  input \State2_reg[1]/NET0131  ;
  input \State2_reg[2]/NET0131  ;
  input \State2_reg[3]/NET0131  ;
  input \State_reg[0]/NET0131  ;
  input \State_reg[1]/NET0131  ;
  input \State_reg[2]/NET0131  ;
  input W_R_n_pad ;
  input \lWord_reg[0]/NET0131  ;
  input \lWord_reg[10]/NET0131  ;
  input \lWord_reg[11]/NET0131  ;
  input \lWord_reg[12]/NET0131  ;
  input \lWord_reg[13]/NET0131  ;
  input \lWord_reg[14]/NET0131  ;
  input \lWord_reg[15]/NET0131  ;
  input \lWord_reg[1]/NET0131  ;
  input \lWord_reg[2]/NET0131  ;
  input \lWord_reg[3]/NET0131  ;
  input \lWord_reg[4]/NET0131  ;
  input \lWord_reg[5]/NET0131  ;
  input \lWord_reg[6]/NET0131  ;
  input \lWord_reg[7]/NET0131  ;
  input \lWord_reg[8]/NET0131  ;
  input \lWord_reg[9]/NET0131  ;
  input \rEIP_reg[0]/NET0131  ;
  input \rEIP_reg[10]/NET0131  ;
  input \rEIP_reg[11]/NET0131  ;
  input \rEIP_reg[12]/NET0131  ;
  input \rEIP_reg[13]/NET0131  ;
  input \rEIP_reg[14]/NET0131  ;
  input \rEIP_reg[15]/NET0131  ;
  input \rEIP_reg[16]/NET0131  ;
  input \rEIP_reg[17]/NET0131  ;
  input \rEIP_reg[18]/NET0131  ;
  input \rEIP_reg[19]/NET0131  ;
  input \rEIP_reg[1]/NET0131  ;
  input \rEIP_reg[20]/NET0131  ;
  input \rEIP_reg[21]/NET0131  ;
  input \rEIP_reg[22]/NET0131  ;
  input \rEIP_reg[23]/NET0131  ;
  input \rEIP_reg[24]/NET0131  ;
  input \rEIP_reg[25]/NET0131  ;
  input \rEIP_reg[26]/NET0131  ;
  input \rEIP_reg[27]/NET0131  ;
  input \rEIP_reg[28]/NET0131  ;
  input \rEIP_reg[29]/NET0131  ;
  input \rEIP_reg[2]/NET0131  ;
  input \rEIP_reg[30]/NET0131  ;
  input \rEIP_reg[31]/NET0131  ;
  input \rEIP_reg[3]/NET0131  ;
  input \rEIP_reg[4]/NET0131  ;
  input \rEIP_reg[5]/NET0131  ;
  input \rEIP_reg[6]/NET0131  ;
  input \rEIP_reg[7]/NET0131  ;
  input \rEIP_reg[8]/NET0131  ;
  input \rEIP_reg[9]/NET0131  ;
  input \uWord_reg[0]/NET0131  ;
  input \uWord_reg[10]/NET0131  ;
  input \uWord_reg[11]/NET0131  ;
  input \uWord_reg[12]/NET0131  ;
  input \uWord_reg[13]/NET0131  ;
  input \uWord_reg[14]/NET0131  ;
  input \uWord_reg[1]/NET0131  ;
  input \uWord_reg[2]/NET0131  ;
  input \uWord_reg[3]/NET0131  ;
  input \uWord_reg[4]/NET0131  ;
  input \uWord_reg[5]/NET0131  ;
  input \uWord_reg[6]/NET0131  ;
  input \uWord_reg[7]/NET0131  ;
  input \uWord_reg[8]/NET0131  ;
  input \uWord_reg[9]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g47521/_2_  ;
  output \g47523/_0_  ;
  output \g47526/_0_  ;
  output \g47529/_0_  ;
  output \g47533/_0_  ;
  output \g47540/_0_  ;
  output \g47551/_0_  ;
  output \g47552/_0_  ;
  output \g47553/_0_  ;
  output \g47563/_2_  ;
  output \g47566/_0_  ;
  output \g47567/_0_  ;
  output \g47568/_0_  ;
  output \g47569/_0_  ;
  output \g47583/_2_  ;
  output \g47584/_0_  ;
  output \g47585/_0_  ;
  output \g47589/_0_  ;
  output \g47602/_0_  ;
  output \g47603/_0_  ;
  output \g47604/_2_  ;
  output \g47605/_0_  ;
  output \g47606/_2_  ;
  output \g47609/_0_  ;
  output \g47611/_0_  ;
  output \g47631/_0_  ;
  output \g47632/_0_  ;
  output \g47633/_0_  ;
  output \g47635/_0_  ;
  output \g47636/_0_  ;
  output \g47637/_0_  ;
  output \g47638/_2_  ;
  output \g47643/_0_  ;
  output \g47665/_2_  ;
  output \g47666/_0_  ;
  output \g47667/_0_  ;
  output \g47670/_0_  ;
  output \g47672/_0_  ;
  output \g47677/_0_  ;
  output \g47678/_0_  ;
  output \g47706/_0_  ;
  output \g47711/_0_  ;
  output \g47717/_0_  ;
  output \g47718/_0_  ;
  output \g47721/_0_  ;
  output \g47722/_0_  ;
  output \g47751/_0_  ;
  output \g47755/_0_  ;
  output \g47756/_0_  ;
  output \g47757/_0_  ;
  output \g47759/_0_  ;
  output \g47789/_0_  ;
  output \g47793/_0_  ;
  output \g47797/_0_  ;
  output \g47798/_0_  ;
  output \g47799/_0_  ;
  output \g47802/_0_  ;
  output \g47804/_0_  ;
  output \g47807/_0_  ;
  output \g47809/_0_  ;
  output \g47862/_0_  ;
  output \g47863/_0_  ;
  output \g47864/_0_  ;
  output \g47869/_0_  ;
  output \g47870/_0_  ;
  output \g47924/_0_  ;
  output \g47925/_0_  ;
  output \g47926/_0_  ;
  output \g47927/_0_  ;
  output \g47928/_0_  ;
  output \g47930/_0_  ;
  output \g47932/_0_  ;
  output \g47933/_0_  ;
  output \g47934/_0_  ;
  output \g47935/_0_  ;
  output \g47936/_0_  ;
  output \g47937/_0_  ;
  output \g47938/_0_  ;
  output \g47939/_0_  ;
  output \g47940/_0_  ;
  output \g47941/_0_  ;
  output \g47957/_0_  ;
  output \g47970/_0_  ;
  output \g47973/_0_  ;
  output \g47975/_0_  ;
  output \g48058/_0_  ;
  output \g48059/_0_  ;
  output \g48060/_0_  ;
  output \g48061/_0_  ;
  output \g48062/_0_  ;
  output \g48064/_0_  ;
  output \g48065/_0_  ;
  output \g48066/_0_  ;
  output \g48067/_0_  ;
  output \g48068/_0_  ;
  output \g48069/_0_  ;
  output \g48070/_0_  ;
  output \g48071/_0_  ;
  output \g48072/_0_  ;
  output \g48073/_0_  ;
  output \g48074/_0_  ;
  output \g48087/_0_  ;
  output \g48110/_0_  ;
  output \g48117/_0_  ;
  output \g48118/_0_  ;
  output \g48119/_0_  ;
  output \g48120/_0_  ;
  output \g48121/_0_  ;
  output \g48122/_0_  ;
  output \g48124/_0_  ;
  output \g48125/_0_  ;
  output \g48126/_0_  ;
  output \g48127/_0_  ;
  output \g48128/_0_  ;
  output \g48129/_0_  ;
  output \g48130/_0_  ;
  output \g48131/_0_  ;
  output \g48132/_0_  ;
  output \g48133/_0_  ;
  output \g48134/_0_  ;
  output \g48168/_0_  ;
  output \g48169/_0_  ;
  output \g48170/_0_  ;
  output \g48171/_0_  ;
  output \g48172/_0_  ;
  output \g48173/_0_  ;
  output \g48174/_0_  ;
  output \g48175/_0_  ;
  output \g48177/_0_  ;
  output \g48178/_0_  ;
  output \g48179/_0_  ;
  output \g48180/_0_  ;
  output \g48181/_0_  ;
  output \g48182/_0_  ;
  output \g48183/_0_  ;
  output \g48184/_0_  ;
  output \g48185/_0_  ;
  output \g48186/_0_  ;
  output \g48187/_0_  ;
  output \g48188/_0_  ;
  output \g48189/_0_  ;
  output \g48192/_0_  ;
  output \g48193/_0_  ;
  output \g48194/_0_  ;
  output \g48195/_0_  ;
  output \g48196/_0_  ;
  output \g48197/_0_  ;
  output \g48198/_0_  ;
  output \g48199/_0_  ;
  output \g48200/_0_  ;
  output \g48201/_0_  ;
  output \g48202/_0_  ;
  output \g48203/_0_  ;
  output \g48213/_0_  ;
  output \g48214/_0_  ;
  output \g48215/_0_  ;
  output \g48216/_0_  ;
  output \g48217/_0_  ;
  output \g48218/_0_  ;
  output \g48219/_0_  ;
  output \g48220/_0_  ;
  output \g48221/_0_  ;
  output \g48222/_0_  ;
  output \g48223/_0_  ;
  output \g48224/_0_  ;
  output \g48225/_0_  ;
  output \g48226/_0_  ;
  output \g48227/_0_  ;
  output \g48228/_0_  ;
  output \g48229/_0_  ;
  output \g48230/_0_  ;
  output \g48231/_0_  ;
  output \g48232/_0_  ;
  output \g48234/_0_  ;
  output \g48236/_0_  ;
  output \g48237/_0_  ;
  output \g48238/_0_  ;
  output \g48239/_0_  ;
  output \g48240/_0_  ;
  output \g48241/_0_  ;
  output \g48243/_0_  ;
  output \g48244/_0_  ;
  output \g48245/_0_  ;
  output \g48246/_0_  ;
  output \g48263/_0_  ;
  output \g48270/_0_  ;
  output \g48273/_0_  ;
  output \g48276/_0_  ;
  output \g48277/_0_  ;
  output \g48370/_0_  ;
  output \g48377/_0_  ;
  output \g48391/_0_  ;
  output \g48423/_0_  ;
  output \g48428/_0_  ;
  output \g48429/_0_  ;
  output \g48431/_0_  ;
  output \g48433/_0_  ;
  output \g48434/_0_  ;
  output \g48435/_0_  ;
  output \g48436/_0_  ;
  output \g48437/_0_  ;
  output \g48438/_0_  ;
  output \g48439/_0_  ;
  output \g48440/_0_  ;
  output \g48441/_0_  ;
  output \g48442/_0_  ;
  output \g48443/_0_  ;
  output \g48610/_0_  ;
  output \g48634/_0_  ;
  output \g48635/_0_  ;
  output \g48636/_0_  ;
  output \g48637/_0_  ;
  output \g48638/_0_  ;
  output \g48639/_0_  ;
  output \g48640/_0_  ;
  output \g48642/_0_  ;
  output \g48643/_0_  ;
  output \g48644/_0_  ;
  output \g48645/_0_  ;
  output \g48646/_0_  ;
  output \g48647/_0_  ;
  output \g48648/_0_  ;
  output \g48649/_0_  ;
  output \g48650/_0_  ;
  output \g48651/_0_  ;
  output \g48652/_0_  ;
  output \g48653/_0_  ;
  output \g48654/_0_  ;
  output \g48655/_0_  ;
  output \g48656/_0_  ;
  output \g48657/_0_  ;
  output \g48658/_0_  ;
  output \g48659/_0_  ;
  output \g48660/_0_  ;
  output \g48662/_0_  ;
  output \g48663/_0_  ;
  output \g48664/_0_  ;
  output \g48665/_0_  ;
  output \g48666/_0_  ;
  output \g48667/_0_  ;
  output \g48668/_0_  ;
  output \g48669/_0_  ;
  output \g48750/_0_  ;
  output \g48753/_0_  ;
  output \g48756/_0_  ;
  output \g48759/_0_  ;
  output \g48763/_0_  ;
  output \g48766/_0_  ;
  output \g48769/_0_  ;
  output \g48772/_0_  ;
  output \g48775/_0_  ;
  output \g48778/_0_  ;
  output \g48781/_0_  ;
  output \g48785/_0_  ;
  output \g48789/_0_  ;
  output \g48792/_0_  ;
  output \g48796/_0_  ;
  output \g48799/_0_  ;
  output \g48937/_0_  ;
  output \g48958/_0_  ;
  output \g48959/_0_  ;
  output \g48964/_0_  ;
  output \g48965/_0_  ;
  output \g48966/_0_  ;
  output \g48967/_0_  ;
  output \g48968/_0_  ;
  output \g48969/_0_  ;
  output \g48970/_0_  ;
  output \g48971/_0_  ;
  output \g48972/_0_  ;
  output \g48973/_0_  ;
  output \g48974/_0_  ;
  output \g48975/_0_  ;
  output \g48976/_0_  ;
  output \g48977/_0_  ;
  output \g48978/_0_  ;
  output \g48979/_0_  ;
  output \g49/_0_  ;
  output \g49069/_0_  ;
  output \g49070/_0_  ;
  output \g49071/_0_  ;
  output \g49073/_0_  ;
  output \g49074/_0_  ;
  output \g49076/_0_  ;
  output \g49078/_0_  ;
  output \g49081/_0_  ;
  output \g49083/_0_  ;
  output \g49085/_0_  ;
  output \g49087/_0_  ;
  output \g49088/_0_  ;
  output \g49090/_0_  ;
  output \g49092/_0_  ;
  output \g49095/_0_  ;
  output \g49098/_0_  ;
  output \g49125/_0_  ;
  output \g49162/_0_  ;
  output \g49202/_0_  ;
  output \g49203/_0_  ;
  output \g49206/_0_  ;
  output \g49340/_0_  ;
  output \g49457/_0_  ;
  output \g49512/_0_  ;
  output \g49513/_0_  ;
  output \g49514/_0_  ;
  output \g49515/_0_  ;
  output \g49516/_0_  ;
  output \g49517/_0_  ;
  output \g49518/_0_  ;
  output \g49519/_0_  ;
  output \g49520/_0_  ;
  output \g49521/_0_  ;
  output \g49522/_0_  ;
  output \g49523/_0_  ;
  output \g49524/_0_  ;
  output \g49525/_0_  ;
  output \g49526/_0_  ;
  output \g49527/_0_  ;
  output \g49534/_0_  ;
  output \g49551/_0_  ;
  output \g49573/_0_  ;
  output \g49574/_0_  ;
  output \g49578/_0_  ;
  output \g49582/_0_  ;
  output \g49584/_0_  ;
  output \g49592/_0_  ;
  output \g49600/_0_  ;
  output \g49604/_0_  ;
  output \g49608/_0_  ;
  output \g49612/_0_  ;
  output \g49616/_0_  ;
  output \g49619/_0_  ;
  output \g49620/_0_  ;
  output \g49623/_0_  ;
  output \g49627/_0_  ;
  output \g49630/_0_  ;
  output \g49634/_0_  ;
  output \g49635/_0_  ;
  output \g49639/_0_  ;
  output \g49645/_0_  ;
  output \g49744/_0_  ;
  output \g49766/_0_  ;
  output \g50098/_0_  ;
  output \g50124/_0_  ;
  output \g50195/_0_  ;
  output \g50198/_0_  ;
  output \g50201/_0_  ;
  output \g50203/_0_  ;
  output \g50205/_0_  ;
  output \g50207/_0_  ;
  output \g50209/_0_  ;
  output \g50213/_0_  ;
  output \g50222/_0_  ;
  output \g50228/_0_  ;
  output \g50231/_0_  ;
  output \g50237/_0_  ;
  output \g50240/_0_  ;
  output \g50335/_0_  ;
  output \g50477/_0_  ;
  output \g50478/_0_  ;
  output \g50671/_0_  ;
  output \g50757/_0_  ;
  output \g50938/_0_  ;
  output \g50998/_0_  ;
  output \g51008/_0_  ;
  output \g51579/_0_  ;
  output \g51637/_0_  ;
  output \g51662/_0_  ;
  output \g52424/_0_  ;
  output \g53184/_0_  ;
  output \g53206/_0_  ;
  output \g53270/_0_  ;
  output \g53730/_0_  ;
  output \g53754/_0_  ;
  output \g54176/_0_  ;
  output \g54214/_0_  ;
  output \g54229/_0_  ;
  output \g54392/_0_  ;
  output \g54400/_0_  ;
  output \g54415/_0_  ;
  output \g54421/_0_  ;
  output \g54604/_0_  ;
  output \g54607/_0_  ;
  output \g54638/_0_  ;
  output \g54694/_0_  ;
  output \g54759/_0_  ;
  output \g55607/_0_  ;
  output \g55863/_1_  ;
  output \g56073/_0_  ;
  output \g56292/_0_  ;
  output \g56320/_0_  ;
  output \g56527/_0_  ;
  output \g56531/_0_  ;
  output \g56533/_0_  ;
  output \g56562/_0_  ;
  output \g56615/_0_  ;
  output \g56720/_0_  ;
  output \g57044/_0_  ;
  output \g60635/_1_  ;
  output \g62873/_0_  ;
  output \g62886/_0_  ;
  output \g63001/_0_  ;
  output \g63101/_0_  ;
  output \g63129/_0_  ;
  output \g63198/_0_  ;
  output \g63449/_0_  ;
  output \g63471/_0_  ;
  output \g63493/_0_  ;
  output \g63626/_0_  ;
  output \g63688/_0_  ;
  output \g63800/_0_  ;
  output \g63934/_0_  ;
  output \g63954/_0_  ;
  output \g64060/_0_  ;
  output \g64375/_0_  ;
  output \g65/_0_  ;
  output \g67/_0_  ;
  wire n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 ;
  assign n459 = ~\InstQueueRd_Addr_reg[2]/NET0131  & ~\InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n465 = \InstQueueRd_Addr_reg[0]/NET0131  & ~\InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n466 = n459 & n465 ;
  assign n467 = \InstQueue_reg[1][7]/NET0131  & n466 ;
  assign n468 = ~\InstQueueRd_Addr_reg[2]/NET0131  & \InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n469 = n465 & n468 ;
  assign n470 = \InstQueue_reg[9][7]/NET0131  & n469 ;
  assign n494 = ~n467 & ~n470 ;
  assign n452 = \InstQueueRd_Addr_reg[2]/NET0131  & \InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n471 = n452 & n465 ;
  assign n472 = \InstQueue_reg[13][7]/NET0131  & n471 ;
  assign n473 = \InstQueueRd_Addr_reg[0]/NET0131  & \InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n474 = n468 & n473 ;
  assign n475 = \InstQueue_reg[11][7]/NET0131  & n474 ;
  assign n495 = ~n472 & ~n475 ;
  assign n502 = n494 & n495 ;
  assign n453 = ~\InstQueueRd_Addr_reg[0]/NET0131  & \InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n454 = n452 & n453 ;
  assign n455 = \InstQueue_reg[14][7]/NET0131  & n454 ;
  assign n456 = \InstQueueRd_Addr_reg[2]/NET0131  & ~\InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n457 = n453 & n456 ;
  assign n458 = \InstQueue_reg[6][7]/NET0131  & n457 ;
  assign n492 = ~n455 & ~n458 ;
  assign n460 = ~\InstQueueRd_Addr_reg[0]/NET0131  & ~\InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n461 = n459 & n460 ;
  assign n462 = \InstQueue_reg[0][7]/NET0131  & n461 ;
  assign n463 = n456 & n460 ;
  assign n464 = \InstQueue_reg[4][7]/NET0131  & n463 ;
  assign n493 = ~n462 & ~n464 ;
  assign n503 = n492 & n493 ;
  assign n504 = n502 & n503 ;
  assign n484 = n456 & n465 ;
  assign n485 = \InstQueue_reg[5][7]/NET0131  & n484 ;
  assign n486 = n460 & n468 ;
  assign n487 = \InstQueue_reg[8][7]/NET0131  & n486 ;
  assign n498 = ~n485 & ~n487 ;
  assign n488 = n452 & n460 ;
  assign n489 = \InstQueue_reg[12][7]/NET0131  & n488 ;
  assign n490 = n453 & n468 ;
  assign n491 = \InstQueue_reg[10][7]/NET0131  & n490 ;
  assign n499 = ~n489 & ~n491 ;
  assign n500 = n498 & n499 ;
  assign n476 = n452 & n473 ;
  assign n477 = \InstQueue_reg[15][7]/NET0131  & n476 ;
  assign n478 = n453 & n459 ;
  assign n479 = \InstQueue_reg[2][7]/NET0131  & n478 ;
  assign n496 = ~n477 & ~n479 ;
  assign n480 = n459 & n473 ;
  assign n481 = \InstQueue_reg[3][7]/NET0131  & n480 ;
  assign n482 = n456 & n473 ;
  assign n483 = \InstQueue_reg[7][7]/NET0131  & n482 ;
  assign n497 = ~n481 & ~n483 ;
  assign n501 = n496 & n497 ;
  assign n505 = n500 & n501 ;
  assign n506 = n504 & n505 ;
  assign n511 = \InstQueue_reg[1][6]/NET0131  & n466 ;
  assign n512 = \InstQueue_reg[0][6]/NET0131  & n461 ;
  assign n525 = ~n511 & ~n512 ;
  assign n513 = \InstQueue_reg[5][6]/NET0131  & n484 ;
  assign n514 = \InstQueue_reg[8][6]/NET0131  & n486 ;
  assign n526 = ~n513 & ~n514 ;
  assign n533 = n525 & n526 ;
  assign n507 = \InstQueue_reg[14][6]/NET0131  & n454 ;
  assign n508 = \InstQueue_reg[11][6]/NET0131  & n474 ;
  assign n523 = ~n507 & ~n508 ;
  assign n509 = \InstQueue_reg[6][6]/NET0131  & n457 ;
  assign n510 = \InstQueue_reg[3][6]/NET0131  & n480 ;
  assign n524 = ~n509 & ~n510 ;
  assign n534 = n523 & n524 ;
  assign n535 = n533 & n534 ;
  assign n519 = \InstQueue_reg[2][6]/NET0131  & n478 ;
  assign n520 = \InstQueue_reg[9][6]/NET0131  & n469 ;
  assign n529 = ~n519 & ~n520 ;
  assign n521 = \InstQueue_reg[13][6]/NET0131  & n471 ;
  assign n522 = \InstQueue_reg[4][6]/NET0131  & n463 ;
  assign n530 = ~n521 & ~n522 ;
  assign n531 = n529 & n530 ;
  assign n515 = \InstQueue_reg[7][6]/NET0131  & n482 ;
  assign n516 = \InstQueue_reg[12][6]/NET0131  & n488 ;
  assign n527 = ~n515 & ~n516 ;
  assign n517 = \InstQueue_reg[10][6]/NET0131  & n490 ;
  assign n518 = \InstQueue_reg[15][6]/NET0131  & n476 ;
  assign n528 = ~n517 & ~n518 ;
  assign n532 = n527 & n528 ;
  assign n536 = n531 & n532 ;
  assign n537 = n535 & n536 ;
  assign n538 = ~n506 & ~n537 ;
  assign n543 = \InstQueue_reg[11][2]/NET0131  & n474 ;
  assign n544 = \InstQueue_reg[14][2]/NET0131  & n454 ;
  assign n557 = ~n543 & ~n544 ;
  assign n545 = \InstQueue_reg[7][2]/NET0131  & n482 ;
  assign n546 = \InstQueue_reg[8][2]/NET0131  & n486 ;
  assign n558 = ~n545 & ~n546 ;
  assign n565 = n557 & n558 ;
  assign n539 = \InstQueue_reg[13][2]/NET0131  & n471 ;
  assign n540 = \InstQueue_reg[2][2]/NET0131  & n478 ;
  assign n555 = ~n539 & ~n540 ;
  assign n541 = \InstQueue_reg[10][2]/NET0131  & n490 ;
  assign n542 = \InstQueue_reg[15][2]/NET0131  & n476 ;
  assign n556 = ~n541 & ~n542 ;
  assign n566 = n555 & n556 ;
  assign n567 = n565 & n566 ;
  assign n551 = \InstQueue_reg[5][2]/NET0131  & n484 ;
  assign n552 = \InstQueue_reg[0][2]/NET0131  & n461 ;
  assign n561 = ~n551 & ~n552 ;
  assign n553 = \InstQueue_reg[9][2]/NET0131  & n469 ;
  assign n554 = \InstQueue_reg[12][2]/NET0131  & n488 ;
  assign n562 = ~n553 & ~n554 ;
  assign n563 = n561 & n562 ;
  assign n547 = \InstQueue_reg[4][2]/NET0131  & n463 ;
  assign n548 = \InstQueue_reg[3][2]/NET0131  & n480 ;
  assign n559 = ~n547 & ~n548 ;
  assign n549 = \InstQueue_reg[1][2]/NET0131  & n466 ;
  assign n550 = \InstQueue_reg[6][2]/NET0131  & n457 ;
  assign n560 = ~n549 & ~n550 ;
  assign n564 = n559 & n560 ;
  assign n568 = n563 & n564 ;
  assign n569 = n567 & n568 ;
  assign n574 = \InstQueue_reg[5][1]/NET0131  & n484 ;
  assign n575 = \InstQueue_reg[14][1]/NET0131  & n454 ;
  assign n588 = ~n574 & ~n575 ;
  assign n576 = \InstQueue_reg[15][1]/NET0131  & n476 ;
  assign n577 = \InstQueue_reg[8][1]/NET0131  & n486 ;
  assign n589 = ~n576 & ~n577 ;
  assign n596 = n588 & n589 ;
  assign n570 = \InstQueue_reg[1][1]/NET0131  & n466 ;
  assign n571 = \InstQueue_reg[0][1]/NET0131  & n461 ;
  assign n586 = ~n570 & ~n571 ;
  assign n572 = \InstQueue_reg[12][1]/NET0131  & n488 ;
  assign n573 = \InstQueue_reg[7][1]/NET0131  & n482 ;
  assign n587 = ~n572 & ~n573 ;
  assign n597 = n586 & n587 ;
  assign n598 = n596 & n597 ;
  assign n582 = \InstQueue_reg[2][1]/NET0131  & n478 ;
  assign n583 = \InstQueue_reg[9][1]/NET0131  & n469 ;
  assign n592 = ~n582 & ~n583 ;
  assign n584 = \InstQueue_reg[3][1]/NET0131  & n480 ;
  assign n585 = \InstQueue_reg[11][1]/NET0131  & n474 ;
  assign n593 = ~n584 & ~n585 ;
  assign n594 = n592 & n593 ;
  assign n578 = \InstQueue_reg[6][1]/NET0131  & n457 ;
  assign n579 = \InstQueue_reg[10][1]/NET0131  & n490 ;
  assign n590 = ~n578 & ~n579 ;
  assign n580 = \InstQueue_reg[13][1]/NET0131  & n471 ;
  assign n581 = \InstQueue_reg[4][1]/NET0131  & n463 ;
  assign n591 = ~n580 & ~n581 ;
  assign n595 = n590 & n591 ;
  assign n599 = n594 & n595 ;
  assign n600 = n598 & n599 ;
  assign n601 = n569 & n600 ;
  assign n606 = \InstQueue_reg[0][3]/NET0131  & n461 ;
  assign n607 = \InstQueue_reg[14][3]/NET0131  & n454 ;
  assign n620 = ~n606 & ~n607 ;
  assign n608 = \InstQueue_reg[12][3]/NET0131  & n488 ;
  assign n609 = \InstQueue_reg[5][3]/NET0131  & n484 ;
  assign n621 = ~n608 & ~n609 ;
  assign n628 = n620 & n621 ;
  assign n602 = \InstQueue_reg[10][3]/NET0131  & n490 ;
  assign n603 = \InstQueue_reg[15][3]/NET0131  & n476 ;
  assign n618 = ~n602 & ~n603 ;
  assign n604 = \InstQueue_reg[1][3]/NET0131  & n466 ;
  assign n605 = \InstQueue_reg[4][3]/NET0131  & n463 ;
  assign n619 = ~n604 & ~n605 ;
  assign n629 = n618 & n619 ;
  assign n630 = n628 & n629 ;
  assign n614 = \InstQueue_reg[6][3]/NET0131  & n457 ;
  assign n615 = \InstQueue_reg[13][3]/NET0131  & n471 ;
  assign n624 = ~n614 & ~n615 ;
  assign n616 = \InstQueue_reg[3][3]/NET0131  & n480 ;
  assign n617 = \InstQueue_reg[7][3]/NET0131  & n482 ;
  assign n625 = ~n616 & ~n617 ;
  assign n626 = n624 & n625 ;
  assign n610 = \InstQueue_reg[2][3]/NET0131  & n478 ;
  assign n611 = \InstQueue_reg[11][3]/NET0131  & n474 ;
  assign n622 = ~n610 & ~n611 ;
  assign n612 = \InstQueue_reg[9][3]/NET0131  & n469 ;
  assign n613 = \InstQueue_reg[8][3]/NET0131  & n486 ;
  assign n623 = ~n612 & ~n613 ;
  assign n627 = n622 & n623 ;
  assign n631 = n626 & n627 ;
  assign n632 = n630 & n631 ;
  assign n637 = \InstQueue_reg[11][0]/NET0131  & n474 ;
  assign n638 = \InstQueue_reg[14][0]/NET0131  & n454 ;
  assign n651 = ~n637 & ~n638 ;
  assign n639 = \InstQueue_reg[9][0]/NET0131  & n469 ;
  assign n640 = \InstQueue_reg[6][0]/NET0131  & n457 ;
  assign n652 = ~n639 & ~n640 ;
  assign n659 = n651 & n652 ;
  assign n633 = \InstQueue_reg[10][0]/NET0131  & n490 ;
  assign n634 = \InstQueue_reg[13][0]/NET0131  & n471 ;
  assign n649 = ~n633 & ~n634 ;
  assign n635 = \InstQueue_reg[1][0]/NET0131  & n466 ;
  assign n636 = \InstQueue_reg[0][0]/NET0131  & n461 ;
  assign n650 = ~n635 & ~n636 ;
  assign n660 = n649 & n650 ;
  assign n661 = n659 & n660 ;
  assign n645 = \InstQueue_reg[8][0]/NET0131  & n486 ;
  assign n646 = \InstQueue_reg[2][0]/NET0131  & n478 ;
  assign n655 = ~n645 & ~n646 ;
  assign n647 = \InstQueue_reg[12][0]/NET0131  & n488 ;
  assign n648 = \InstQueue_reg[15][0]/NET0131  & n476 ;
  assign n656 = ~n647 & ~n648 ;
  assign n657 = n655 & n656 ;
  assign n641 = \InstQueue_reg[4][0]/NET0131  & n463 ;
  assign n642 = \InstQueue_reg[3][0]/NET0131  & n480 ;
  assign n653 = ~n641 & ~n642 ;
  assign n643 = \InstQueue_reg[5][0]/NET0131  & n484 ;
  assign n644 = \InstQueue_reg[7][0]/NET0131  & n482 ;
  assign n654 = ~n643 & ~n644 ;
  assign n658 = n653 & n654 ;
  assign n662 = n657 & n658 ;
  assign n663 = n661 & n662 ;
  assign n664 = n632 & n663 ;
  assign n665 = n601 & n664 ;
  assign n666 = n538 & n665 ;
  assign n671 = \InstQueue_reg[5][5]/NET0131  & n484 ;
  assign n672 = \InstQueue_reg[1][5]/NET0131  & n466 ;
  assign n685 = ~n671 & ~n672 ;
  assign n673 = \InstQueue_reg[15][5]/NET0131  & n476 ;
  assign n674 = \InstQueue_reg[12][5]/NET0131  & n488 ;
  assign n686 = ~n673 & ~n674 ;
  assign n693 = n685 & n686 ;
  assign n667 = \InstQueue_reg[14][5]/NET0131  & n454 ;
  assign n668 = \InstQueue_reg[4][5]/NET0131  & n463 ;
  assign n683 = ~n667 & ~n668 ;
  assign n669 = \InstQueue_reg[10][5]/NET0131  & n490 ;
  assign n670 = \InstQueue_reg[2][5]/NET0131  & n478 ;
  assign n684 = ~n669 & ~n670 ;
  assign n694 = n683 & n684 ;
  assign n695 = n693 & n694 ;
  assign n679 = \InstQueue_reg[13][5]/NET0131  & n471 ;
  assign n680 = \InstQueue_reg[0][5]/NET0131  & n461 ;
  assign n689 = ~n679 & ~n680 ;
  assign n681 = \InstQueue_reg[11][5]/NET0131  & n474 ;
  assign n682 = \InstQueue_reg[7][5]/NET0131  & n482 ;
  assign n690 = ~n681 & ~n682 ;
  assign n691 = n689 & n690 ;
  assign n675 = \InstQueue_reg[9][5]/NET0131  & n469 ;
  assign n676 = \InstQueue_reg[6][5]/NET0131  & n457 ;
  assign n687 = ~n675 & ~n676 ;
  assign n677 = \InstQueue_reg[3][5]/NET0131  & n480 ;
  assign n678 = \InstQueue_reg[8][5]/NET0131  & n486 ;
  assign n688 = ~n677 & ~n678 ;
  assign n692 = n687 & n688 ;
  assign n696 = n691 & n692 ;
  assign n697 = n695 & n696 ;
  assign n698 = n666 & n697 ;
  assign n699 = ~n632 & ~n663 ;
  assign n700 = n569 & ~n600 ;
  assign n701 = n699 & n700 ;
  assign n702 = ~n506 & n537 ;
  assign n707 = \InstQueue_reg[11][4]/NET0131  & n474 ;
  assign n708 = \InstQueue_reg[3][4]/NET0131  & n480 ;
  assign n721 = ~n707 & ~n708 ;
  assign n709 = \InstQueue_reg[15][4]/NET0131  & n476 ;
  assign n710 = \InstQueue_reg[8][4]/NET0131  & n486 ;
  assign n722 = ~n709 & ~n710 ;
  assign n729 = n721 & n722 ;
  assign n703 = \InstQueue_reg[14][4]/NET0131  & n454 ;
  assign n704 = \InstQueue_reg[12][4]/NET0131  & n488 ;
  assign n719 = ~n703 & ~n704 ;
  assign n705 = \InstQueue_reg[2][4]/NET0131  & n478 ;
  assign n706 = \InstQueue_reg[1][4]/NET0131  & n466 ;
  assign n720 = ~n705 & ~n706 ;
  assign n730 = n719 & n720 ;
  assign n731 = n729 & n730 ;
  assign n715 = \InstQueue_reg[0][4]/NET0131  & n461 ;
  assign n716 = \InstQueue_reg[5][4]/NET0131  & n484 ;
  assign n725 = ~n715 & ~n716 ;
  assign n717 = \InstQueue_reg[10][4]/NET0131  & n490 ;
  assign n718 = \InstQueue_reg[7][4]/NET0131  & n482 ;
  assign n726 = ~n717 & ~n718 ;
  assign n727 = n725 & n726 ;
  assign n711 = \InstQueue_reg[6][4]/NET0131  & n457 ;
  assign n712 = \InstQueue_reg[13][4]/NET0131  & n471 ;
  assign n723 = ~n711 & ~n712 ;
  assign n713 = \InstQueue_reg[4][4]/NET0131  & n463 ;
  assign n714 = \InstQueue_reg[9][4]/NET0131  & n469 ;
  assign n724 = ~n713 & ~n714 ;
  assign n728 = n723 & n724 ;
  assign n732 = n727 & n728 ;
  assign n733 = n731 & n732 ;
  assign n734 = n697 & n733 ;
  assign n735 = n702 & n734 ;
  assign n736 = n701 & n735 ;
  assign n737 = ~n697 & n733 ;
  assign n738 = n538 & n737 ;
  assign n739 = ~n569 & n664 ;
  assign n740 = n738 & n739 ;
  assign n741 = n601 & n699 ;
  assign n742 = n735 & n741 ;
  assign n743 = ~n740 & ~n742 ;
  assign n744 = ~n736 & n743 ;
  assign n745 = ~n698 & n744 ;
  assign n746 = n738 & n741 ;
  assign n747 = n700 & n738 ;
  assign n748 = n699 & n747 ;
  assign n749 = ~n746 & ~n748 ;
  assign n750 = n702 & ~n733 ;
  assign n751 = ~n697 & n750 ;
  assign n752 = n701 & n751 ;
  assign n753 = ~n632 & n663 ;
  assign n754 = n601 & n753 ;
  assign n755 = n751 & n754 ;
  assign n756 = ~n752 & ~n755 ;
  assign n757 = n749 & n756 ;
  assign n758 = n745 & n757 ;
  assign n759 = n506 & n537 ;
  assign n760 = n600 & n759 ;
  assign n761 = n734 & n760 ;
  assign n762 = n506 & ~n537 ;
  assign n763 = ~n600 & n737 ;
  assign n764 = n762 & n763 ;
  assign n765 = ~n761 & ~n764 ;
  assign n766 = n739 & ~n765 ;
  assign n767 = n734 & n762 ;
  assign n768 = ~n750 & ~n767 ;
  assign n769 = n665 & ~n768 ;
  assign n771 = n632 & ~n663 ;
  assign n772 = n700 & n771 ;
  assign n773 = n767 & n772 ;
  assign n776 = ~n769 & ~n773 ;
  assign n770 = n747 & n753 ;
  assign n774 = ~n569 & n771 ;
  assign n775 = n761 & n774 ;
  assign n777 = ~n770 & ~n775 ;
  assign n778 = n776 & n777 ;
  assign n779 = ~n766 & n778 ;
  assign n780 = ~n758 & n779 ;
  assign n781 = ~\InstQueueRd_Addr_reg[0]/NET0131  & \InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n782 = \InstQueueRd_Addr_reg[0]/NET0131  & ~\InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n783 = ~\InstQueueRd_Addr_reg[1]/NET0131  & \InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n784 = \InstQueueRd_Addr_reg[1]/NET0131  & ~\InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n785 = ~n783 & ~n784 ;
  assign n786 = ~n782 & n785 ;
  assign n787 = ~n781 & n786 ;
  assign n788 = ~n782 & ~n784 ;
  assign n789 = ~n783 & ~n788 ;
  assign n790 = ~\InstQueueRd_Addr_reg[2]/NET0131  & \InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n791 = \InstQueueRd_Addr_reg[2]/NET0131  & ~\InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n792 = ~n790 & ~n791 ;
  assign n793 = n789 & n792 ;
  assign n794 = ~n789 & ~n792 ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = ~n787 & ~n795 ;
  assign n797 = ~\InstQueueRd_Addr_reg[3]/NET0131  & \InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n798 = \InstQueueRd_Addr_reg[3]/NET0131  & ~\InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n799 = ~n797 & ~n798 ;
  assign n800 = ~n789 & ~n791 ;
  assign n801 = ~n790 & ~n800 ;
  assign n802 = n799 & n801 ;
  assign n803 = ~n799 & ~n801 ;
  assign n804 = ~n802 & ~n803 ;
  assign n805 = ~n796 & n804 ;
  assign n806 = ~n798 & ~n801 ;
  assign n807 = ~n797 & ~n806 ;
  assign n808 = ~n805 & ~n807 ;
  assign n809 = ~n756 & n808 ;
  assign n810 = n780 & ~n809 ;
  assign n819 = ~n453 & ~n465 ;
  assign n820 = ~n810 & ~n819 ;
  assign n821 = n795 & n804 ;
  assign n822 = n782 & ~n785 ;
  assign n823 = ~n786 & ~n822 ;
  assign n824 = n821 & ~n823 ;
  assign n825 = ~n807 & ~n824 ;
  assign n826 = ~READY_n_pad & n825 ;
  assign n827 = ~n600 & n740 ;
  assign n828 = ~n742 & ~n827 ;
  assign n829 = ~\State_reg[0]/NET0131  & \State_reg[1]/NET0131  ;
  assign n830 = ~\State_reg[2]/NET0131  & n829 ;
  assign n831 = ~\State_reg[0]/NET0131  & ~\State_reg[1]/NET0131  ;
  assign n832 = \State_reg[2]/NET0131  & n831 ;
  assign n833 = ~n830 & ~n832 ;
  assign n834 = ~n828 & ~n833 ;
  assign n835 = n600 & n740 ;
  assign n836 = ~n736 & ~n835 ;
  assign n837 = ~n834 & n836 ;
  assign n838 = n826 & ~n837 ;
  assign n839 = ~n698 & ~n838 ;
  assign n840 = ~\InstQueueRd_Addr_reg[1]/NET0131  & n839 ;
  assign n841 = ~n828 & n833 ;
  assign n842 = ~n743 & ~n826 ;
  assign n843 = ~n841 & ~n842 ;
  assign n844 = n736 & ~n826 ;
  assign n845 = n843 & ~n844 ;
  assign n812 = ~n756 & ~n808 ;
  assign n813 = n749 & ~n812 ;
  assign n846 = \InstQueueRd_Addr_reg[1]/NET0131  & n813 ;
  assign n847 = n845 & n846 ;
  assign n848 = ~n840 & ~n847 ;
  assign n849 = ~n820 & ~n848 ;
  assign n811 = ~\InstQueueRd_Addr_reg[0]/NET0131  & n810 ;
  assign n814 = \InstQueueRd_Addr_reg[0]/NET0131  & n745 ;
  assign n815 = n813 & n814 ;
  assign n816 = ~n811 & ~n815 ;
  assign n817 = \InstQueueWr_Addr_reg[0]/NET0131  & ~n816 ;
  assign n850 = ~\InstQueueWr_Addr_reg[1]/NET0131  & ~n817 ;
  assign n851 = n849 & ~n850 ;
  assign n861 = ~READY_n_pad & ~n833 ;
  assign n862 = n825 & n861 ;
  assign n872 = ~n826 & n835 ;
  assign n873 = ~n844 & ~n872 ;
  assign n874 = n828 & n873 ;
  assign n875 = ~n862 & ~n874 ;
  assign n857 = ~\InstQueueRd_Addr_reg[2]/NET0131  & ~n473 ;
  assign n858 = n808 & ~n857 ;
  assign n876 = ~n756 & ~n858 ;
  assign n877 = n749 & ~n876 ;
  assign n878 = ~n875 & n877 ;
  assign n879 = \InstQueueRd_Addr_reg[3]/NET0131  & ~n878 ;
  assign n864 = n825 & ~n836 ;
  assign n865 = ~READY_n_pad & n864 ;
  assign n863 = ~n828 & n862 ;
  assign n866 = ~n698 & ~n863 ;
  assign n867 = ~n865 & n866 ;
  assign n852 = \InstQueueRd_Addr_reg[1]/NET0131  & \InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n868 = ~\InstQueueRd_Addr_reg[3]/NET0131  & ~n852 ;
  assign n869 = \InstQueueRd_Addr_reg[3]/NET0131  & n852 ;
  assign n870 = ~n868 & ~n869 ;
  assign n871 = ~n867 & n870 ;
  assign n853 = \InstQueueRd_Addr_reg[0]/NET0131  & n852 ;
  assign n854 = \InstQueueRd_Addr_reg[3]/NET0131  & ~n853 ;
  assign n855 = ~n482 & ~n854 ;
  assign n856 = ~n780 & ~n855 ;
  assign n859 = ~\InstQueueRd_Addr_reg[3]/NET0131  & n858 ;
  assign n860 = ~n756 & n859 ;
  assign n880 = ~n856 & ~n860 ;
  assign n881 = ~n871 & n880 ;
  assign n882 = ~n879 & n881 ;
  assign n883 = \InstQueueWr_Addr_reg[3]/NET0131  & n882 ;
  assign n818 = \InstQueueWr_Addr_reg[1]/NET0131  & n817 ;
  assign n884 = ~n853 & ~n857 ;
  assign n885 = ~n780 & n884 ;
  assign n887 = ~\InstQueueRd_Addr_reg[1]/NET0131  & ~\InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n888 = ~n852 & ~n887 ;
  assign n889 = ~READY_n_pad & ~n888 ;
  assign n890 = ~\InstQueueRd_Addr_reg[2]/NET0131  & READY_n_pad ;
  assign n891 = ~n889 & ~n890 ;
  assign n895 = n825 & ~n833 ;
  assign n897 = ~n891 & n895 ;
  assign n896 = ~\InstQueueRd_Addr_reg[2]/NET0131  & ~n895 ;
  assign n898 = ~n828 & ~n896 ;
  assign n899 = ~n897 & n898 ;
  assign n886 = ~\InstQueueRd_Addr_reg[2]/NET0131  & ~n825 ;
  assign n892 = n825 & ~n891 ;
  assign n893 = ~n886 & ~n892 ;
  assign n894 = ~n836 & n893 ;
  assign n904 = n698 & n888 ;
  assign n906 = ~n894 & ~n904 ;
  assign n900 = ~\InstQueueRd_Addr_reg[2]/NET0131  & ~n808 ;
  assign n901 = n808 & n884 ;
  assign n902 = ~n900 & ~n901 ;
  assign n903 = ~n756 & n902 ;
  assign n905 = \InstQueueRd_Addr_reg[2]/NET0131  & ~n749 ;
  assign n907 = ~n903 & ~n905 ;
  assign n908 = n906 & n907 ;
  assign n909 = ~n899 & n908 ;
  assign n910 = ~n885 & n909 ;
  assign n911 = \InstQueueWr_Addr_reg[2]/NET0131  & n910 ;
  assign n912 = ~n818 & ~n911 ;
  assign n913 = ~n883 & n912 ;
  assign n914 = ~n851 & n913 ;
  assign n937 = ~\InstQueueWr_Addr_reg[2]/NET0131  & ~n910 ;
  assign n938 = ~n883 & n937 ;
  assign n927 = \InstQueueWr_Addr_reg[3]/NET0131  & n910 ;
  assign n928 = ~n882 & ~n927 ;
  assign n915 = \More_reg/NET0131  & ~n861 ;
  assign n916 = n825 & ~n915 ;
  assign n917 = ~n874 & ~n916 ;
  assign n918 = ~n781 & ~n785 ;
  assign n919 = ~n786 & ~n918 ;
  assign n920 = n821 & ~n919 ;
  assign n921 = ~n807 & ~n920 ;
  assign n922 = n748 & ~n921 ;
  assign n923 = n746 & ~n808 ;
  assign n924 = ~n812 & ~n923 ;
  assign n925 = ~n922 & n924 ;
  assign n926 = ~n917 & n925 ;
  assign n931 = READY_n_pad & ~n744 ;
  assign n932 = ~n841 & ~n931 ;
  assign n933 = \Flush_reg/NET0131  & n825 ;
  assign n934 = ~n932 & n933 ;
  assign n929 = n748 & n921 ;
  assign n930 = n746 & n808 ;
  assign n935 = ~n929 & ~n930 ;
  assign n936 = ~n934 & n935 ;
  assign n939 = n926 & n936 ;
  assign n940 = ~n928 & n939 ;
  assign n941 = ~n938 & n940 ;
  assign n942 = ~n914 & n941 ;
  assign n943 = ~\DataWidth_reg[1]/NET0131  & n742 ;
  assign n944 = n862 & n943 ;
  assign n945 = n942 & ~n944 ;
  assign n946 = \State2_reg[0]/NET0131  & ~\State2_reg[3]/NET0131  ;
  assign n947 = ~\State2_reg[1]/NET0131  & \State2_reg[2]/NET0131  ;
  assign n948 = n946 & n947 ;
  assign n949 = ~n945 & n948 ;
  assign n954 = \State2_reg[1]/NET0131  & \State2_reg[2]/NET0131  ;
  assign n955 = ~\State2_reg[3]/NET0131  & n954 ;
  assign n956 = ~\State2_reg[0]/NET0131  & n955 ;
  assign n950 = \State2_reg[1]/NET0131  & ~\State2_reg[2]/NET0131  ;
  assign n951 = ~\State2_reg[3]/NET0131  & n950 ;
  assign n957 = \State2_reg[0]/NET0131  & n951 ;
  assign n958 = ~n956 & ~n957 ;
  assign n959 = READY_n_pad & ~n958 ;
  assign n952 = ~\State2_reg[0]/NET0131  & n951 ;
  assign n953 = ~\DataWidth_reg[1]/NET0131  & n952 ;
  assign n960 = ~\State2_reg[1]/NET0131  & ~\State2_reg[2]/NET0131  ;
  assign n961 = \State2_reg[0]/NET0131  & n960 ;
  assign n962 = ~\State2_reg[3]/NET0131  & n961 ;
  assign n963 = ~READY_n_pad & n962 ;
  assign n964 = ~n953 & ~n963 ;
  assign n965 = ~n959 & n964 ;
  assign n966 = ~n949 & n965 ;
  assign n968 = ~\State2_reg[0]/NET0131  & ~\State2_reg[3]/NET0131  ;
  assign n969 = \State2_reg[2]/NET0131  & n968 ;
  assign n970 = ~\State2_reg[1]/NET0131  & n969 ;
  assign n971 = \DataWidth_reg[1]/NET0131  & n952 ;
  assign n972 = ~n970 & ~n971 ;
  assign n967 = ~READY_n_pad & n957 ;
  assign n973 = ~n948 & ~n956 ;
  assign n974 = ~n967 & n973 ;
  assign n975 = n972 & n974 ;
  assign n976 = n942 & n944 ;
  assign n977 = n948 & ~n976 ;
  assign n984 = \State2_reg[0]/NET0131  & n955 ;
  assign n985 = ~\Flush_reg/NET0131  & \InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n986 = \InstQueueRd_Addr_reg[3]/NET0131  & ~n460 ;
  assign n987 = n985 & n986 ;
  assign n988 = n984 & ~n987 ;
  assign n982 = ~\State2_reg[2]/NET0131  & n946 ;
  assign n983 = READY_n_pad & n982 ;
  assign n978 = READY_n_pad & n954 ;
  assign n979 = n968 & ~n978 ;
  assign n980 = \State2_reg[3]/NET0131  & n960 ;
  assign n981 = \State2_reg[0]/NET0131  & n980 ;
  assign n989 = ~n979 & ~n981 ;
  assign n990 = ~n983 & n989 ;
  assign n991 = ~n988 & n990 ;
  assign n992 = ~n977 & n991 ;
  assign n993 = ~\State2_reg[0]/NET0131  & n980 ;
  assign n994 = ~n984 & ~n993 ;
  assign n995 = \InstAddrPointer_reg[31]/NET0131  & ~n921 ;
  assign n996 = \InstAddrPointer_reg[1]/NET0131  & \InstAddrPointer_reg[2]/NET0131  ;
  assign n997 = \InstAddrPointer_reg[3]/NET0131  & n996 ;
  assign n998 = \InstAddrPointer_reg[4]/NET0131  & n997 ;
  assign n999 = \InstAddrPointer_reg[5]/NET0131  & \InstAddrPointer_reg[6]/NET0131  ;
  assign n1000 = n998 & n999 ;
  assign n1001 = \InstAddrPointer_reg[7]/NET0131  & n1000 ;
  assign n1002 = \InstAddrPointer_reg[8]/NET0131  & n1001 ;
  assign n1006 = \InstAddrPointer_reg[9]/NET0131  & n1002 ;
  assign n1007 = \InstAddrPointer_reg[10]/NET0131  & n1006 ;
  assign n1008 = ~\InstAddrPointer_reg[11]/NET0131  & ~n1007 ;
  assign n1009 = \InstAddrPointer_reg[10]/NET0131  & \InstAddrPointer_reg[11]/NET0131  ;
  assign n1010 = n1006 & n1009 ;
  assign n1011 = ~n1008 & ~n1010 ;
  assign n1012 = \InstAddrPointer_reg[12]/NET0131  & n1011 ;
  assign n1013 = \InstAddrPointer_reg[13]/NET0131  & n1012 ;
  assign n1003 = ~\InstAddrPointer_reg[8]/NET0131  & ~n1001 ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1005 = \InstAddrPointer_reg[9]/NET0131  & n1004 ;
  assign n1014 = \InstAddrPointer_reg[10]/NET0131  & n1005 ;
  assign n1015 = n1013 & n1014 ;
  assign n1019 = n855 & ~n884 ;
  assign n1158 = \InstQueue_reg[2][3]/NET0131  & n465 ;
  assign n1159 = \InstQueue_reg[1][3]/NET0131  & n460 ;
  assign n1160 = ~n1158 & ~n1159 ;
  assign n1161 = n1019 & ~n1160 ;
  assign n1162 = \InstQueue_reg[0][3]/NET0131  & n476 ;
  assign n1163 = \InstQueue_reg[13][3]/NET0131  & n488 ;
  assign n1176 = ~n1162 & ~n1163 ;
  assign n1164 = \InstQueue_reg[4][3]/NET0131  & n480 ;
  assign n1165 = \InstQueue_reg[9][3]/NET0131  & n486 ;
  assign n1177 = ~n1164 & ~n1165 ;
  assign n1166 = \InstQueue_reg[14][3]/NET0131  & n471 ;
  assign n1167 = \InstQueue_reg[3][3]/NET0131  & n478 ;
  assign n1178 = ~n1166 & ~n1167 ;
  assign n1185 = n1177 & n1178 ;
  assign n1186 = n1176 & n1185 ;
  assign n1172 = \InstQueue_reg[5][3]/NET0131  & n463 ;
  assign n1173 = \InstQueue_reg[8][3]/NET0131  & n482 ;
  assign n1181 = ~n1172 & ~n1173 ;
  assign n1174 = \InstQueue_reg[6][3]/NET0131  & n484 ;
  assign n1175 = \InstQueue_reg[12][3]/NET0131  & n474 ;
  assign n1182 = ~n1174 & ~n1175 ;
  assign n1183 = n1181 & n1182 ;
  assign n1168 = \InstQueue_reg[11][3]/NET0131  & n490 ;
  assign n1169 = \InstQueue_reg[7][3]/NET0131  & n457 ;
  assign n1179 = ~n1168 & ~n1169 ;
  assign n1170 = \InstQueue_reg[10][3]/NET0131  & n469 ;
  assign n1171 = \InstQueue_reg[15][3]/NET0131  & n454 ;
  assign n1180 = ~n1170 & ~n1171 ;
  assign n1184 = n1179 & n1180 ;
  assign n1187 = n1183 & n1184 ;
  assign n1188 = n1186 & n1187 ;
  assign n1189 = ~n1161 & n1188 ;
  assign n1190 = ~\InstAddrPointer_reg[3]/NET0131  & ~n996 ;
  assign n1191 = ~n997 & ~n1190 ;
  assign n1192 = n1189 & ~n1191 ;
  assign n1193 = ~\InstAddrPointer_reg[1]/NET0131  & ~\InstAddrPointer_reg[2]/NET0131  ;
  assign n1194 = ~n996 & ~n1193 ;
  assign n1199 = \InstQueue_reg[10][2]/NET0131  & n469 ;
  assign n1200 = \InstQueue_reg[6][2]/NET0131  & n484 ;
  assign n1213 = ~n1199 & ~n1200 ;
  assign n1201 = \InstQueue_reg[12][2]/NET0131  & n474 ;
  assign n1202 = \InstQueue_reg[11][2]/NET0131  & n490 ;
  assign n1214 = ~n1201 & ~n1202 ;
  assign n1221 = n1213 & n1214 ;
  assign n1195 = \InstQueue_reg[15][2]/NET0131  & n454 ;
  assign n1196 = \InstQueue_reg[14][2]/NET0131  & n471 ;
  assign n1211 = ~n1195 & ~n1196 ;
  assign n1197 = \InstQueue_reg[9][2]/NET0131  & n486 ;
  assign n1198 = \InstQueue_reg[2][2]/NET0131  & n466 ;
  assign n1212 = ~n1197 & ~n1198 ;
  assign n1222 = n1211 & n1212 ;
  assign n1223 = n1221 & n1222 ;
  assign n1207 = \InstQueue_reg[8][2]/NET0131  & n482 ;
  assign n1208 = \InstQueue_reg[3][2]/NET0131  & n478 ;
  assign n1217 = ~n1207 & ~n1208 ;
  assign n1209 = \InstQueue_reg[13][2]/NET0131  & n488 ;
  assign n1210 = \InstQueue_reg[0][2]/NET0131  & n476 ;
  assign n1218 = ~n1209 & ~n1210 ;
  assign n1219 = n1217 & n1218 ;
  assign n1203 = \InstQueue_reg[1][2]/NET0131  & n461 ;
  assign n1204 = \InstQueue_reg[5][2]/NET0131  & n463 ;
  assign n1215 = ~n1203 & ~n1204 ;
  assign n1205 = \InstQueue_reg[7][2]/NET0131  & n457 ;
  assign n1206 = \InstQueue_reg[4][2]/NET0131  & n480 ;
  assign n1216 = ~n1205 & ~n1206 ;
  assign n1220 = n1215 & n1216 ;
  assign n1224 = n1219 & n1220 ;
  assign n1225 = n1223 & n1224 ;
  assign n1226 = ~n1194 & n1225 ;
  assign n1227 = ~n1192 & ~n1226 ;
  assign n1232 = \InstQueue_reg[7][1]/NET0131  & n457 ;
  assign n1233 = \InstQueue_reg[13][1]/NET0131  & n488 ;
  assign n1250 = ~n1232 & ~n1233 ;
  assign n1234 = \InstQueue_reg[1][1]/NET0131  & n461 ;
  assign n1235 = \InstQueue_reg[6][1]/NET0131  & n484 ;
  assign n1251 = ~n1234 & ~n1235 ;
  assign n1255 = n1250 & n1251 ;
  assign n1228 = \InstQueue_reg[12][1]/NET0131  & n474 ;
  assign n1229 = \InstQueue_reg[14][1]/NET0131  & n471 ;
  assign n1248 = ~n1228 & ~n1229 ;
  assign n1230 = \InstQueue_reg[5][1]/NET0131  & n463 ;
  assign n1231 = \InstQueue_reg[11][1]/NET0131  & n490 ;
  assign n1249 = ~n1230 & ~n1231 ;
  assign n1256 = n1248 & n1249 ;
  assign n1257 = n1255 & n1256 ;
  assign n1133 = \InstQueueRd_Addr_reg[3]/NET0131  & n884 ;
  assign n1236 = \InstQueue_reg[15][1]/NET0131  & n453 ;
  assign n1237 = n1133 & n1236 ;
  assign n1238 = \InstQueue_reg[9][1]/NET0131  & n486 ;
  assign n1239 = \InstQueue_reg[4][1]/NET0131  & n480 ;
  assign n1252 = ~n1238 & ~n1239 ;
  assign n1240 = \InstQueue_reg[8][1]/NET0131  & n482 ;
  assign n1241 = \InstQueue_reg[0][1]/NET0131  & n476 ;
  assign n1253 = ~n1240 & ~n1241 ;
  assign n1254 = n1252 & n1253 ;
  assign n1258 = ~n1237 & n1254 ;
  assign n1259 = n1257 & n1258 ;
  assign n1021 = ~n855 & ~n884 ;
  assign n1242 = \InstQueue_reg[10][1]/NET0131  & n465 ;
  assign n1243 = n1021 & n1242 ;
  assign n1244 = \InstQueue_reg[2][1]/NET0131  & n465 ;
  assign n1245 = \InstQueue_reg[3][1]/NET0131  & n453 ;
  assign n1246 = ~n1244 & ~n1245 ;
  assign n1247 = n1019 & ~n1246 ;
  assign n1260 = ~n1243 & ~n1247 ;
  assign n1261 = n1259 & n1260 ;
  assign n1262 = ~\InstAddrPointer_reg[1]/NET0131  & ~n1261 ;
  assign n1263 = \InstAddrPointer_reg[1]/NET0131  & n1261 ;
  assign n1268 = \InstQueue_reg[10][0]/NET0131  & n469 ;
  assign n1269 = \InstQueue_reg[2][0]/NET0131  & n466 ;
  assign n1282 = ~n1268 & ~n1269 ;
  assign n1270 = \InstQueue_reg[3][0]/NET0131  & n478 ;
  assign n1271 = \InstQueue_reg[13][0]/NET0131  & n488 ;
  assign n1283 = ~n1270 & ~n1271 ;
  assign n1290 = n1282 & n1283 ;
  assign n1264 = \InstQueue_reg[15][0]/NET0131  & n454 ;
  assign n1265 = \InstQueue_reg[9][0]/NET0131  & n486 ;
  assign n1280 = ~n1264 & ~n1265 ;
  assign n1266 = \InstQueue_reg[7][0]/NET0131  & n457 ;
  assign n1267 = \InstQueue_reg[5][0]/NET0131  & n463 ;
  assign n1281 = ~n1266 & ~n1267 ;
  assign n1291 = n1280 & n1281 ;
  assign n1292 = n1290 & n1291 ;
  assign n1276 = \InstQueue_reg[8][0]/NET0131  & n482 ;
  assign n1277 = \InstQueue_reg[1][0]/NET0131  & n461 ;
  assign n1286 = ~n1276 & ~n1277 ;
  assign n1278 = \InstQueue_reg[6][0]/NET0131  & n484 ;
  assign n1279 = \InstQueue_reg[0][0]/NET0131  & n476 ;
  assign n1287 = ~n1278 & ~n1279 ;
  assign n1288 = n1286 & n1287 ;
  assign n1272 = \InstQueue_reg[14][0]/NET0131  & n471 ;
  assign n1273 = \InstQueue_reg[11][0]/NET0131  & n490 ;
  assign n1284 = ~n1272 & ~n1273 ;
  assign n1274 = \InstQueue_reg[12][0]/NET0131  & n474 ;
  assign n1275 = \InstQueue_reg[4][0]/NET0131  & n480 ;
  assign n1285 = ~n1274 & ~n1275 ;
  assign n1289 = n1284 & n1285 ;
  assign n1293 = n1288 & n1289 ;
  assign n1294 = n1292 & n1293 ;
  assign n1295 = \InstAddrPointer_reg[0]/NET0131  & ~n1294 ;
  assign n1296 = ~n1263 & n1295 ;
  assign n1297 = ~n1262 & ~n1296 ;
  assign n1298 = n1227 & ~n1297 ;
  assign n1299 = ~n1189 & n1191 ;
  assign n1300 = n1194 & ~n1225 ;
  assign n1301 = ~n1192 & n1300 ;
  assign n1302 = ~n1299 & ~n1301 ;
  assign n1303 = ~n1298 & n1302 ;
  assign n1053 = \InstAddrPointer_reg[5]/NET0131  & n998 ;
  assign n1088 = ~\InstAddrPointer_reg[5]/NET0131  & ~n998 ;
  assign n1089 = ~n1053 & ~n1088 ;
  assign n1094 = \InstQueue_reg[4][5]/NET0131  & n480 ;
  assign n1095 = \InstQueue_reg[15][5]/NET0131  & n454 ;
  assign n1108 = ~n1094 & ~n1095 ;
  assign n1096 = \InstQueue_reg[11][5]/NET0131  & n490 ;
  assign n1097 = \InstQueue_reg[13][5]/NET0131  & n488 ;
  assign n1109 = ~n1096 & ~n1097 ;
  assign n1116 = n1108 & n1109 ;
  assign n1090 = \InstQueue_reg[9][5]/NET0131  & n486 ;
  assign n1091 = \InstQueue_reg[12][5]/NET0131  & n474 ;
  assign n1106 = ~n1090 & ~n1091 ;
  assign n1092 = \InstQueue_reg[2][5]/NET0131  & n466 ;
  assign n1093 = \InstQueue_reg[0][5]/NET0131  & n476 ;
  assign n1107 = ~n1092 & ~n1093 ;
  assign n1117 = n1106 & n1107 ;
  assign n1118 = n1116 & n1117 ;
  assign n1102 = \InstQueue_reg[1][5]/NET0131  & n461 ;
  assign n1103 = \InstQueue_reg[6][5]/NET0131  & n484 ;
  assign n1112 = ~n1102 & ~n1103 ;
  assign n1104 = \InstQueue_reg[14][5]/NET0131  & n471 ;
  assign n1105 = \InstQueue_reg[10][5]/NET0131  & n469 ;
  assign n1113 = ~n1104 & ~n1105 ;
  assign n1114 = n1112 & n1113 ;
  assign n1098 = \InstQueue_reg[8][5]/NET0131  & n482 ;
  assign n1099 = \InstQueue_reg[3][5]/NET0131  & n478 ;
  assign n1110 = ~n1098 & ~n1099 ;
  assign n1100 = \InstQueue_reg[5][5]/NET0131  & n463 ;
  assign n1101 = \InstQueue_reg[7][5]/NET0131  & n457 ;
  assign n1111 = ~n1100 & ~n1101 ;
  assign n1115 = n1110 & n1111 ;
  assign n1119 = n1114 & n1115 ;
  assign n1120 = n1118 & n1119 ;
  assign n1121 = ~n1089 & n1120 ;
  assign n1122 = ~\InstAddrPointer_reg[4]/NET0131  & ~n997 ;
  assign n1123 = ~n998 & ~n1122 ;
  assign n1128 = \InstQueue_reg[11][4]/NET0131  & n490 ;
  assign n1129 = \InstQueue_reg[1][4]/NET0131  & n461 ;
  assign n1144 = ~n1128 & ~n1129 ;
  assign n1130 = \InstQueue_reg[4][4]/NET0131  & n480 ;
  assign n1131 = \InstQueue_reg[6][4]/NET0131  & n484 ;
  assign n1145 = ~n1130 & ~n1131 ;
  assign n1151 = n1144 & n1145 ;
  assign n1124 = \InstQueue_reg[5][4]/NET0131  & n463 ;
  assign n1125 = \InstQueue_reg[2][4]/NET0131  & n466 ;
  assign n1142 = ~n1124 & ~n1125 ;
  assign n1126 = \InstQueue_reg[10][4]/NET0131  & n469 ;
  assign n1127 = \InstQueue_reg[15][4]/NET0131  & n454 ;
  assign n1143 = ~n1126 & ~n1127 ;
  assign n1152 = n1142 & n1143 ;
  assign n1153 = n1151 & n1152 ;
  assign n1134 = \InstQueue_reg[13][4]/NET0131  & n460 ;
  assign n1135 = n1133 & n1134 ;
  assign n1141 = \InstQueue_reg[9][4]/NET0131  & n486 ;
  assign n1139 = \InstQueue_reg[7][4]/NET0131  & n457 ;
  assign n1140 = \InstQueue_reg[3][4]/NET0131  & n478 ;
  assign n1148 = ~n1139 & ~n1140 ;
  assign n1149 = ~n1141 & n1148 ;
  assign n1132 = \InstQueue_reg[12][4]/NET0131  & n474 ;
  assign n1136 = \InstQueue_reg[8][4]/NET0131  & n482 ;
  assign n1146 = ~n1132 & ~n1136 ;
  assign n1137 = \InstQueue_reg[14][4]/NET0131  & n471 ;
  assign n1138 = \InstQueue_reg[0][4]/NET0131  & n476 ;
  assign n1147 = ~n1137 & ~n1138 ;
  assign n1150 = n1146 & n1147 ;
  assign n1154 = n1149 & n1150 ;
  assign n1155 = ~n1135 & n1154 ;
  assign n1156 = n1153 & n1155 ;
  assign n1157 = ~n1123 & n1156 ;
  assign n1304 = ~n1121 & ~n1157 ;
  assign n1305 = ~n1303 & n1304 ;
  assign n1306 = n1089 & ~n1120 ;
  assign n1307 = n1123 & ~n1156 ;
  assign n1308 = ~n1121 & n1307 ;
  assign n1309 = ~n1306 & ~n1308 ;
  assign n1310 = ~n1305 & n1309 ;
  assign n1016 = ~\InstAddrPointer_reg[7]/NET0131  & ~n1000 ;
  assign n1017 = ~n1001 & ~n1016 ;
  assign n1020 = \InstQueue_reg[0][7]/NET0131  & n1019 ;
  assign n1022 = \InstQueue_reg[8][7]/NET0131  & n1021 ;
  assign n1023 = ~n1020 & ~n1022 ;
  assign n1024 = n473 & ~n1023 ;
  assign n1018 = \InstQueue_reg[6][7]/NET0131  & n484 ;
  assign n1025 = \InstQueue_reg[9][7]/NET0131  & n486 ;
  assign n1038 = ~n1018 & ~n1025 ;
  assign n1026 = \InstQueue_reg[13][7]/NET0131  & n488 ;
  assign n1027 = \InstQueue_reg[14][7]/NET0131  & n471 ;
  assign n1039 = ~n1026 & ~n1027 ;
  assign n1028 = \InstQueue_reg[15][7]/NET0131  & n454 ;
  assign n1029 = \InstQueue_reg[10][7]/NET0131  & n469 ;
  assign n1040 = ~n1028 & ~n1029 ;
  assign n1047 = n1039 & n1040 ;
  assign n1048 = n1038 & n1047 ;
  assign n1034 = \InstQueue_reg[11][7]/NET0131  & n490 ;
  assign n1035 = \InstQueue_reg[1][7]/NET0131  & n461 ;
  assign n1043 = ~n1034 & ~n1035 ;
  assign n1036 = \InstQueue_reg[3][7]/NET0131  & n478 ;
  assign n1037 = \InstQueue_reg[5][7]/NET0131  & n463 ;
  assign n1044 = ~n1036 & ~n1037 ;
  assign n1045 = n1043 & n1044 ;
  assign n1030 = \InstQueue_reg[2][7]/NET0131  & n466 ;
  assign n1031 = \InstQueue_reg[7][7]/NET0131  & n457 ;
  assign n1041 = ~n1030 & ~n1031 ;
  assign n1032 = \InstQueue_reg[4][7]/NET0131  & n480 ;
  assign n1033 = \InstQueue_reg[12][7]/NET0131  & n474 ;
  assign n1042 = ~n1032 & ~n1033 ;
  assign n1046 = n1041 & n1042 ;
  assign n1049 = n1045 & n1046 ;
  assign n1050 = n1048 & n1049 ;
  assign n1051 = ~n1024 & n1050 ;
  assign n1052 = ~n1017 & n1051 ;
  assign n1054 = ~\InstAddrPointer_reg[6]/NET0131  & ~n1053 ;
  assign n1055 = ~n1000 & ~n1054 ;
  assign n1060 = \InstQueue_reg[9][6]/NET0131  & n486 ;
  assign n1061 = \InstQueue_reg[15][6]/NET0131  & n454 ;
  assign n1074 = ~n1060 & ~n1061 ;
  assign n1062 = \InstQueue_reg[13][6]/NET0131  & n488 ;
  assign n1063 = \InstQueue_reg[10][6]/NET0131  & n469 ;
  assign n1075 = ~n1062 & ~n1063 ;
  assign n1082 = n1074 & n1075 ;
  assign n1056 = \InstQueue_reg[8][6]/NET0131  & n482 ;
  assign n1057 = \InstQueue_reg[11][6]/NET0131  & n490 ;
  assign n1072 = ~n1056 & ~n1057 ;
  assign n1058 = \InstQueue_reg[6][6]/NET0131  & n484 ;
  assign n1059 = \InstQueue_reg[3][6]/NET0131  & n478 ;
  assign n1073 = ~n1058 & ~n1059 ;
  assign n1083 = n1072 & n1073 ;
  assign n1084 = n1082 & n1083 ;
  assign n1068 = \InstQueue_reg[1][6]/NET0131  & n461 ;
  assign n1069 = \InstQueue_reg[12][6]/NET0131  & n474 ;
  assign n1078 = ~n1068 & ~n1069 ;
  assign n1070 = \InstQueue_reg[5][6]/NET0131  & n463 ;
  assign n1071 = \InstQueue_reg[0][6]/NET0131  & n476 ;
  assign n1079 = ~n1070 & ~n1071 ;
  assign n1080 = n1078 & n1079 ;
  assign n1064 = \InstQueue_reg[7][6]/NET0131  & n457 ;
  assign n1065 = \InstQueue_reg[4][6]/NET0131  & n480 ;
  assign n1076 = ~n1064 & ~n1065 ;
  assign n1066 = \InstQueue_reg[14][6]/NET0131  & n471 ;
  assign n1067 = \InstQueue_reg[2][6]/NET0131  & n466 ;
  assign n1077 = ~n1066 & ~n1067 ;
  assign n1081 = n1076 & n1077 ;
  assign n1085 = n1080 & n1081 ;
  assign n1086 = n1084 & n1085 ;
  assign n1087 = ~n1055 & n1086 ;
  assign n1311 = ~n1052 & ~n1087 ;
  assign n1312 = ~n1310 & n1311 ;
  assign n1313 = n1017 & ~n1051 ;
  assign n1314 = n1055 & ~n1086 ;
  assign n1315 = ~n1052 & n1314 ;
  assign n1316 = ~n1313 & ~n1315 ;
  assign n1317 = ~n1312 & n1316 ;
  assign n1318 = n1015 & ~n1317 ;
  assign n1319 = \InstAddrPointer_reg[12]/NET0131  & n1009 ;
  assign n1320 = \InstAddrPointer_reg[9]/NET0131  & n1319 ;
  assign n1321 = n1002 & n1320 ;
  assign n1322 = \InstAddrPointer_reg[13]/NET0131  & n1321 ;
  assign n1323 = ~\InstAddrPointer_reg[14]/NET0131  & ~n1322 ;
  assign n1324 = \InstAddrPointer_reg[14]/NET0131  & n1322 ;
  assign n1325 = ~n1323 & ~n1324 ;
  assign n1326 = n1318 & n1325 ;
  assign n1331 = \InstAddrPointer_reg[13]/NET0131  & \InstAddrPointer_reg[14]/NET0131  ;
  assign n1332 = \InstAddrPointer_reg[15]/NET0131  & n1331 ;
  assign n1333 = \InstAddrPointer_reg[16]/NET0131  & n1319 ;
  assign n1334 = n1332 & n1333 ;
  assign n1335 = \InstAddrPointer_reg[9]/NET0131  & n1334 ;
  assign n1336 = n1002 & n1335 ;
  assign n1337 = \InstAddrPointer_reg[18]/NET0131  & \InstAddrPointer_reg[19]/NET0131  ;
  assign n1338 = \InstAddrPointer_reg[17]/NET0131  & n1337 ;
  assign n1339 = n1336 & n1338 ;
  assign n1329 = \InstAddrPointer_reg[20]/NET0131  & \InstAddrPointer_reg[21]/NET0131  ;
  assign n1330 = \InstAddrPointer_reg[22]/NET0131  & n1329 ;
  assign n1347 = \InstAddrPointer_reg[23]/NET0131  & n1330 ;
  assign n1348 = \InstAddrPointer_reg[24]/NET0131  & n1347 ;
  assign n1349 = n1339 & n1348 ;
  assign n1350 = \InstAddrPointer_reg[25]/NET0131  & n1349 ;
  assign n1351 = ~\InstAddrPointer_reg[26]/NET0131  & ~n1350 ;
  assign n1352 = \InstAddrPointer_reg[26]/NET0131  & n1350 ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = ~\InstAddrPointer_reg[25]/NET0131  & ~n1349 ;
  assign n1355 = ~n1350 & ~n1354 ;
  assign n1356 = n1353 & n1355 ;
  assign n1340 = n1330 & n1339 ;
  assign n1341 = \InstAddrPointer_reg[23]/NET0131  & n1340 ;
  assign n1357 = ~\InstAddrPointer_reg[24]/NET0131  & ~n1341 ;
  assign n1358 = ~n1349 & ~n1357 ;
  assign n1359 = n1356 & n1358 ;
  assign n1360 = ~\InstAddrPointer_reg[23]/NET0131  & ~n1340 ;
  assign n1361 = ~n1341 & ~n1360 ;
  assign n1362 = n1359 & n1361 ;
  assign n1327 = \InstAddrPointer_reg[24]/NET0131  & \InstAddrPointer_reg[25]/NET0131  ;
  assign n1328 = \InstAddrPointer_reg[26]/NET0131  & n1327 ;
  assign n1342 = n1328 & n1341 ;
  assign n1343 = ~\InstAddrPointer_reg[27]/NET0131  & ~n1342 ;
  assign n1344 = \InstAddrPointer_reg[27]/NET0131  & n1342 ;
  assign n1345 = ~n1343 & ~n1344 ;
  assign n1346 = \InstAddrPointer_reg[28]/NET0131  & n1345 ;
  assign n1363 = \InstAddrPointer_reg[27]/NET0131  & \InstAddrPointer_reg[28]/NET0131  ;
  assign n1364 = n1352 & n1363 ;
  assign n1365 = ~\InstAddrPointer_reg[29]/NET0131  & ~n1364 ;
  assign n1366 = \InstAddrPointer_reg[29]/NET0131  & n1363 ;
  assign n1367 = n1352 & n1366 ;
  assign n1368 = ~n1365 & ~n1367 ;
  assign n1369 = n1346 & n1368 ;
  assign n1370 = n1362 & n1369 ;
  assign n1371 = \InstAddrPointer_reg[30]/NET0131  & n1370 ;
  assign n1372 = ~\InstAddrPointer_reg[15]/NET0131  & ~n1324 ;
  assign n1373 = \InstAddrPointer_reg[15]/NET0131  & n1324 ;
  assign n1374 = ~n1372 & ~n1373 ;
  assign n1378 = \InstAddrPointer_reg[16]/NET0131  & ~n1373 ;
  assign n1379 = ~\InstAddrPointer_reg[16]/NET0131  & n1373 ;
  assign n1380 = ~n1378 & ~n1379 ;
  assign n1381 = \InstAddrPointer_reg[17]/NET0131  & n1336 ;
  assign n1382 = ~\InstAddrPointer_reg[17]/NET0131  & ~n1336 ;
  assign n1383 = ~n1381 & ~n1382 ;
  assign n1384 = ~n1380 & n1383 ;
  assign n1385 = \InstAddrPointer_reg[18]/NET0131  & n1381 ;
  assign n1386 = ~\InstAddrPointer_reg[18]/NET0131  & ~n1381 ;
  assign n1387 = ~n1385 & ~n1386 ;
  assign n1388 = \InstAddrPointer_reg[19]/NET0131  & n1387 ;
  assign n1389 = n1384 & n1388 ;
  assign n1375 = n1329 & n1339 ;
  assign n1376 = ~\InstAddrPointer_reg[22]/NET0131  & ~n1375 ;
  assign n1377 = ~n1340 & ~n1376 ;
  assign n1390 = \InstAddrPointer_reg[20]/NET0131  & n1339 ;
  assign n1391 = ~\InstAddrPointer_reg[20]/NET0131  & ~n1339 ;
  assign n1392 = ~n1390 & ~n1391 ;
  assign n1393 = \InstAddrPointer_reg[21]/NET0131  & n1392 ;
  assign n1394 = n1377 & n1393 ;
  assign n1395 = n1389 & n1394 ;
  assign n1396 = n1374 & n1395 ;
  assign n1397 = n1371 & n1396 ;
  assign n1398 = n1326 & n1397 ;
  assign n1399 = \InstAddrPointer_reg[30]/NET0131  & n1366 ;
  assign n1400 = n1342 & n1399 ;
  assign n1401 = \InstAddrPointer_reg[31]/NET0131  & ~n1400 ;
  assign n1402 = ~\InstAddrPointer_reg[31]/NET0131  & n1400 ;
  assign n1403 = ~n1401 & ~n1402 ;
  assign n1404 = ~n1398 & n1403 ;
  assign n1405 = n1297 & ~n1300 ;
  assign n1406 = ~n1157 & n1227 ;
  assign n1407 = ~n1405 & n1406 ;
  assign n1408 = ~n1157 & n1299 ;
  assign n1409 = ~n1307 & ~n1408 ;
  assign n1410 = ~n1407 & n1409 ;
  assign n1411 = ~n1087 & ~n1121 ;
  assign n1412 = ~n1410 & n1411 ;
  assign n1413 = ~n1087 & n1306 ;
  assign n1414 = ~n1314 & ~n1413 ;
  assign n1415 = ~n1313 & n1414 ;
  assign n1416 = ~n1412 & n1415 ;
  assign n1417 = n1004 & ~n1052 ;
  assign n1418 = ~n1416 & n1417 ;
  assign n1419 = ~\InstAddrPointer_reg[9]/NET0131  & ~n1002 ;
  assign n1420 = ~n1006 & ~n1419 ;
  assign n1421 = \InstAddrPointer_reg[10]/NET0131  & n1420 ;
  assign n1422 = n1418 & n1421 ;
  assign n1423 = \InstAddrPointer_reg[15]/NET0131  & n1325 ;
  assign n1424 = n1013 & n1423 ;
  assign n1425 = n1395 & n1424 ;
  assign n1426 = n1422 & n1425 ;
  assign n1427 = n1371 & ~n1403 ;
  assign n1428 = n1426 & n1427 ;
  assign n1429 = n1051 & ~n1428 ;
  assign n1430 = ~n1404 & n1429 ;
  assign n1431 = \InstAddrPointer_reg[0]/NET0131  & \InstAddrPointer_reg[1]/NET0131  ;
  assign n1432 = \InstAddrPointer_reg[2]/NET0131  & n1431 ;
  assign n1433 = \InstAddrPointer_reg[3]/NET0131  & n1432 ;
  assign n1434 = \InstAddrPointer_reg[4]/NET0131  & n1433 ;
  assign n1435 = n999 & n1434 ;
  assign n1436 = ~\InstAddrPointer_reg[7]/NET0131  & ~n1435 ;
  assign n1437 = \InstAddrPointer_reg[7]/NET0131  & n1435 ;
  assign n1438 = ~n1436 & ~n1437 ;
  assign n1439 = n1051 & ~n1438 ;
  assign n1440 = \InstAddrPointer_reg[5]/NET0131  & n1434 ;
  assign n1441 = ~\InstAddrPointer_reg[6]/NET0131  & ~n1440 ;
  assign n1442 = ~n1435 & ~n1441 ;
  assign n1443 = n1086 & ~n1442 ;
  assign n1444 = ~\InstAddrPointer_reg[5]/NET0131  & ~n1434 ;
  assign n1445 = ~n1440 & ~n1444 ;
  assign n1446 = n1120 & ~n1445 ;
  assign n1447 = ~n1443 & ~n1446 ;
  assign n1448 = ~\InstAddrPointer_reg[2]/NET0131  & ~n1431 ;
  assign n1449 = ~n1432 & ~n1448 ;
  assign n1450 = ~n1225 & n1449 ;
  assign n1451 = \InstAddrPointer_reg[0]/NET0131  & n1294 ;
  assign n1452 = ~n1262 & n1451 ;
  assign n1453 = n1225 & ~n1449 ;
  assign n1454 = ~\InstAddrPointer_reg[0]/NET0131  & ~\InstAddrPointer_reg[1]/NET0131  ;
  assign n1455 = ~n1431 & ~n1454 ;
  assign n1456 = n1261 & ~n1455 ;
  assign n1457 = ~n1453 & ~n1456 ;
  assign n1458 = ~n1452 & n1457 ;
  assign n1459 = ~n1450 & ~n1458 ;
  assign n1460 = ~\InstAddrPointer_reg[4]/NET0131  & ~n1433 ;
  assign n1461 = ~n1434 & ~n1460 ;
  assign n1462 = n1156 & ~n1461 ;
  assign n1463 = ~\InstAddrPointer_reg[3]/NET0131  & ~n1432 ;
  assign n1464 = ~n1433 & ~n1463 ;
  assign n1465 = n1189 & ~n1464 ;
  assign n1466 = ~n1462 & ~n1465 ;
  assign n1467 = ~n1459 & n1466 ;
  assign n1468 = n1447 & n1467 ;
  assign n1469 = ~n1156 & n1461 ;
  assign n1470 = ~n1189 & n1464 ;
  assign n1471 = ~n1462 & n1470 ;
  assign n1472 = ~n1469 & ~n1471 ;
  assign n1473 = n1447 & ~n1472 ;
  assign n1474 = ~n1086 & n1442 ;
  assign n1475 = ~n1120 & n1445 ;
  assign n1476 = ~n1443 & n1475 ;
  assign n1477 = ~n1474 & ~n1476 ;
  assign n1478 = ~n1473 & n1477 ;
  assign n1479 = ~n1468 & n1478 ;
  assign n1480 = ~n1439 & ~n1479 ;
  assign n1481 = \InstAddrPointer_reg[0]/NET0131  & n1006 ;
  assign n1482 = ~\InstAddrPointer_reg[10]/NET0131  & ~n1481 ;
  assign n1483 = \InstAddrPointer_reg[10]/NET0131  & n1481 ;
  assign n1484 = ~n1482 & ~n1483 ;
  assign n1485 = \InstAddrPointer_reg[8]/NET0131  & n1437 ;
  assign n1486 = ~\InstAddrPointer_reg[9]/NET0131  & ~n1485 ;
  assign n1487 = ~n1481 & ~n1486 ;
  assign n1488 = ~n1484 & ~n1487 ;
  assign n1489 = ~n1051 & n1438 ;
  assign n1490 = ~\InstAddrPointer_reg[8]/NET0131  & ~n1437 ;
  assign n1491 = ~n1485 & ~n1490 ;
  assign n1492 = ~n1489 & ~n1491 ;
  assign n1493 = n1488 & n1492 ;
  assign n1494 = ~n1480 & n1493 ;
  assign n1495 = n1009 & n1481 ;
  assign n1496 = ~\InstAddrPointer_reg[12]/NET0131  & ~n1495 ;
  assign n1497 = n1320 & n1485 ;
  assign n1498 = ~n1496 & ~n1497 ;
  assign n1499 = ~\InstAddrPointer_reg[11]/NET0131  & ~n1483 ;
  assign n1500 = ~n1495 & ~n1499 ;
  assign n1501 = ~n1498 & ~n1500 ;
  assign n1502 = ~\InstAddrPointer_reg[13]/NET0131  & ~n1497 ;
  assign n1503 = \InstAddrPointer_reg[13]/NET0131  & n1497 ;
  assign n1504 = ~n1502 & ~n1503 ;
  assign n1505 = ~\InstAddrPointer_reg[14]/NET0131  & ~n1503 ;
  assign n1506 = \InstAddrPointer_reg[0]/NET0131  & n1324 ;
  assign n1507 = ~n1505 & ~n1506 ;
  assign n1508 = ~n1504 & ~n1507 ;
  assign n1509 = n1501 & n1508 ;
  assign n1510 = ~\InstAddrPointer_reg[15]/NET0131  & ~n1506 ;
  assign n1511 = \InstAddrPointer_reg[15]/NET0131  & n1506 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = n1509 & ~n1512 ;
  assign n1514 = ~\InstAddrPointer_reg[16]/NET0131  & ~n1511 ;
  assign n1515 = \InstAddrPointer_reg[0]/NET0131  & n1336 ;
  assign n1516 = ~n1514 & ~n1515 ;
  assign n1517 = \InstAddrPointer_reg[0]/NET0131  & n1381 ;
  assign n1518 = ~\InstAddrPointer_reg[18]/NET0131  & ~n1517 ;
  assign n1519 = \InstAddrPointer_reg[0]/NET0131  & n1385 ;
  assign n1520 = ~n1518 & ~n1519 ;
  assign n1521 = ~\InstAddrPointer_reg[17]/NET0131  & ~n1515 ;
  assign n1522 = ~n1517 & ~n1521 ;
  assign n1523 = ~n1520 & ~n1522 ;
  assign n1524 = ~n1516 & n1523 ;
  assign n1525 = n1513 & n1524 ;
  assign n1526 = n1494 & n1525 ;
  assign n1527 = ~\InstAddrPointer_reg[19]/NET0131  & ~n1519 ;
  assign n1528 = n1338 & n1515 ;
  assign n1529 = ~n1527 & ~n1528 ;
  assign n1537 = n1348 & n1528 ;
  assign n1545 = \InstAddrPointer_reg[0]/NET0131  & n1340 ;
  assign n1547 = \InstAddrPointer_reg[23]/NET0131  & n1545 ;
  assign n1551 = ~\InstAddrPointer_reg[24]/NET0131  & ~n1547 ;
  assign n1552 = ~n1537 & ~n1551 ;
  assign n1546 = ~\InstAddrPointer_reg[23]/NET0131  & ~n1545 ;
  assign n1548 = ~n1546 & ~n1547 ;
  assign n1532 = \InstAddrPointer_reg[0]/NET0131  & n1375 ;
  assign n1549 = ~\InstAddrPointer_reg[22]/NET0131  & ~n1532 ;
  assign n1550 = ~n1545 & ~n1549 ;
  assign n1553 = ~n1548 & ~n1550 ;
  assign n1554 = ~n1552 & n1553 ;
  assign n1530 = \InstAddrPointer_reg[20]/NET0131  & n1528 ;
  assign n1531 = ~\InstAddrPointer_reg[21]/NET0131  & ~n1530 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = ~\InstAddrPointer_reg[20]/NET0131  & ~n1528 ;
  assign n1535 = ~n1530 & ~n1534 ;
  assign n1536 = ~n1533 & ~n1535 ;
  assign n1538 = \InstAddrPointer_reg[25]/NET0131  & n1537 ;
  assign n1539 = ~\InstAddrPointer_reg[25]/NET0131  & ~n1537 ;
  assign n1540 = ~n1538 & ~n1539 ;
  assign n1541 = \InstAddrPointer_reg[26]/NET0131  & ~n1538 ;
  assign n1542 = ~\InstAddrPointer_reg[26]/NET0131  & n1538 ;
  assign n1543 = ~n1541 & ~n1542 ;
  assign n1544 = ~n1540 & n1543 ;
  assign n1555 = n1536 & n1544 ;
  assign n1556 = n1554 & n1555 ;
  assign n1557 = ~n1529 & n1556 ;
  assign n1558 = n1526 & n1557 ;
  assign n1559 = \InstAddrPointer_reg[0]/NET0131  & n1364 ;
  assign n1560 = \InstAddrPointer_reg[29]/NET0131  & n1559 ;
  assign n1561 = \InstAddrPointer_reg[30]/NET0131  & ~n1560 ;
  assign n1562 = ~\InstAddrPointer_reg[30]/NET0131  & n1560 ;
  assign n1563 = ~n1561 & ~n1562 ;
  assign n1564 = \InstAddrPointer_reg[0]/NET0131  & n1342 ;
  assign n1565 = ~\InstAddrPointer_reg[27]/NET0131  & ~n1564 ;
  assign n1566 = \InstAddrPointer_reg[27]/NET0131  & n1564 ;
  assign n1567 = ~n1565 & ~n1566 ;
  assign n1568 = ~\InstAddrPointer_reg[28]/NET0131  & ~n1566 ;
  assign n1569 = n1363 & n1564 ;
  assign n1570 = ~n1568 & ~n1569 ;
  assign n1571 = ~n1567 & ~n1570 ;
  assign n1572 = \InstAddrPointer_reg[29]/NET0131  & ~n1559 ;
  assign n1573 = ~\InstAddrPointer_reg[29]/NET0131  & n1559 ;
  assign n1574 = ~n1572 & ~n1573 ;
  assign n1575 = n1571 & n1574 ;
  assign n1576 = n1563 & n1575 ;
  assign n1577 = n1558 & n1576 ;
  assign n1578 = \InstAddrPointer_reg[0]/NET0131  & n1400 ;
  assign n1579 = \InstAddrPointer_reg[31]/NET0131  & ~n1578 ;
  assign n1580 = \InstAddrPointer_reg[0]/NET0131  & n1402 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1582 = ~n1051 & ~n1581 ;
  assign n1583 = ~n1577 & n1582 ;
  assign n1584 = ~n1051 & n1581 ;
  assign n1585 = n1577 & n1584 ;
  assign n1586 = ~n1583 & ~n1585 ;
  assign n1587 = ~n1430 & n1586 ;
  assign n1588 = n921 & ~n1587 ;
  assign n1589 = ~n995 & ~n1588 ;
  assign n1590 = n748 & ~n1589 ;
  assign n1591 = \InstAddrPointer_reg[3]/NET0131  & ~n1448 ;
  assign n1592 = \InstAddrPointer_reg[4]/NET0131  & n1591 ;
  assign n1608 = ~\InstAddrPointer_reg[4]/NET0131  & ~n1591 ;
  assign n1609 = ~n1592 & ~n1608 ;
  assign n1610 = n1156 & ~n1609 ;
  assign n1611 = ~\InstAddrPointer_reg[3]/NET0131  & n1448 ;
  assign n1612 = ~n1591 & ~n1611 ;
  assign n1613 = n1189 & ~n1612 ;
  assign n1614 = ~n1610 & ~n1613 ;
  assign n1615 = n1225 & n1449 ;
  assign n1616 = ~n1225 & ~n1449 ;
  assign n1617 = ~n1261 & n1455 ;
  assign n1618 = ~\InstAddrPointer_reg[0]/NET0131  & ~n1294 ;
  assign n1619 = ~n1617 & ~n1618 ;
  assign n1620 = ~n1456 & ~n1619 ;
  assign n1621 = ~n1616 & ~n1620 ;
  assign n1622 = ~n1615 & ~n1621 ;
  assign n1623 = n1614 & n1622 ;
  assign n1624 = ~n1156 & n1609 ;
  assign n1625 = ~n1189 & n1612 ;
  assign n1626 = ~n1610 & n1625 ;
  assign n1627 = ~n1624 & ~n1626 ;
  assign n1628 = ~n1623 & n1627 ;
  assign n1601 = \InstAddrPointer_reg[5]/NET0131  & n1592 ;
  assign n1602 = ~\InstAddrPointer_reg[5]/NET0131  & ~n1592 ;
  assign n1603 = ~n1601 & ~n1602 ;
  assign n1604 = n1120 & ~n1603 ;
  assign n1593 = n999 & n1592 ;
  assign n1605 = ~\InstAddrPointer_reg[6]/NET0131  & ~n1601 ;
  assign n1606 = ~n1593 & ~n1605 ;
  assign n1607 = n1086 & ~n1606 ;
  assign n1629 = ~n1604 & ~n1607 ;
  assign n1630 = ~n1628 & n1629 ;
  assign n1594 = \InstAddrPointer_reg[7]/NET0131  & n1593 ;
  assign n1631 = ~\InstAddrPointer_reg[7]/NET0131  & ~n1593 ;
  assign n1632 = ~n1594 & ~n1631 ;
  assign n1633 = ~n1051 & n1632 ;
  assign n1634 = ~n1086 & n1606 ;
  assign n1635 = ~n1120 & n1603 ;
  assign n1636 = ~n1607 & n1635 ;
  assign n1637 = ~n1634 & ~n1636 ;
  assign n1638 = ~n1633 & n1637 ;
  assign n1639 = ~n1630 & n1638 ;
  assign n1640 = n1051 & ~n1632 ;
  assign n1595 = \InstAddrPointer_reg[8]/NET0131  & n1594 ;
  assign n1641 = ~\InstAddrPointer_reg[8]/NET0131  & ~n1594 ;
  assign n1642 = ~n1595 & ~n1641 ;
  assign n1643 = ~n1640 & n1642 ;
  assign n1644 = ~n1639 & n1643 ;
  assign n1645 = n1320 & n1595 ;
  assign n1646 = \InstAddrPointer_reg[13]/NET0131  & n1645 ;
  assign n1659 = \InstAddrPointer_reg[14]/NET0131  & n1646 ;
  assign n1660 = ~\InstAddrPointer_reg[15]/NET0131  & ~n1659 ;
  assign n1661 = \InstAddrPointer_reg[15]/NET0131  & n1659 ;
  assign n1662 = ~n1660 & ~n1661 ;
  assign n1663 = \InstAddrPointer_reg[16]/NET0131  & n1662 ;
  assign n1596 = \InstAddrPointer_reg[9]/NET0131  & n1595 ;
  assign n1649 = \InstAddrPointer_reg[10]/NET0131  & n1596 ;
  assign n1650 = ~\InstAddrPointer_reg[11]/NET0131  & ~n1649 ;
  assign n1651 = \InstAddrPointer_reg[11]/NET0131  & n1649 ;
  assign n1652 = ~n1650 & ~n1651 ;
  assign n1653 = \InstAddrPointer_reg[12]/NET0131  & n1652 ;
  assign n1647 = ~\InstAddrPointer_reg[13]/NET0131  & ~n1645 ;
  assign n1648 = ~n1646 & ~n1647 ;
  assign n1654 = \InstAddrPointer_reg[14]/NET0131  & n1648 ;
  assign n1655 = n1653 & n1654 ;
  assign n1656 = ~\InstAddrPointer_reg[9]/NET0131  & ~n1595 ;
  assign n1657 = ~n1596 & ~n1656 ;
  assign n1658 = \InstAddrPointer_reg[10]/NET0131  & n1657 ;
  assign n1664 = n1655 & n1658 ;
  assign n1665 = n1663 & n1664 ;
  assign n1666 = n1644 & n1665 ;
  assign n1597 = n1334 & n1596 ;
  assign n1598 = ~\InstAddrPointer_reg[17]/NET0131  & ~n1597 ;
  assign n1599 = \InstAddrPointer_reg[17]/NET0131  & n1597 ;
  assign n1600 = ~n1598 & ~n1599 ;
  assign n1667 = n1337 & n1600 ;
  assign n1668 = n1666 & n1667 ;
  assign n1669 = n1338 & n1597 ;
  assign n1670 = \InstAddrPointer_reg[20]/NET0131  & n1669 ;
  assign n1671 = ~\InstAddrPointer_reg[20]/NET0131  & ~n1669 ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = \InstAddrPointer_reg[21]/NET0131  & n1672 ;
  assign n1674 = n1668 & n1673 ;
  assign n1675 = n1347 & n1669 ;
  assign n1676 = n1328 & n1675 ;
  assign n1677 = n1363 & n1676 ;
  assign n1678 = \InstAddrPointer_reg[29]/NET0131  & n1677 ;
  assign n1679 = ~\InstAddrPointer_reg[30]/NET0131  & ~n1678 ;
  assign n1680 = \InstAddrPointer_reg[30]/NET0131  & n1678 ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1685 = \InstAddrPointer_reg[24]/NET0131  & n1675 ;
  assign n1686 = \InstAddrPointer_reg[25]/NET0131  & n1685 ;
  assign n1687 = ~\InstAddrPointer_reg[26]/NET0131  & ~n1686 ;
  assign n1688 = ~n1676 & ~n1687 ;
  assign n1689 = n1329 & n1669 ;
  assign n1690 = ~\InstAddrPointer_reg[22]/NET0131  & ~n1689 ;
  assign n1691 = \InstAddrPointer_reg[22]/NET0131  & n1689 ;
  assign n1692 = ~n1690 & ~n1691 ;
  assign n1693 = \InstAddrPointer_reg[23]/NET0131  & n1692 ;
  assign n1694 = ~\InstAddrPointer_reg[24]/NET0131  & ~n1675 ;
  assign n1695 = ~n1685 & ~n1694 ;
  assign n1696 = n1693 & n1695 ;
  assign n1697 = \InstAddrPointer_reg[25]/NET0131  & n1696 ;
  assign n1698 = n1688 & n1697 ;
  assign n1699 = ~\InstAddrPointer_reg[29]/NET0131  & ~n1677 ;
  assign n1700 = ~n1678 & ~n1699 ;
  assign n1682 = \InstAddrPointer_reg[27]/NET0131  & n1676 ;
  assign n1683 = ~\InstAddrPointer_reg[28]/NET0131  & ~n1682 ;
  assign n1684 = ~n1677 & ~n1683 ;
  assign n1701 = \InstAddrPointer_reg[27]/NET0131  & n1684 ;
  assign n1702 = n1700 & n1701 ;
  assign n1703 = n1698 & n1702 ;
  assign n1704 = n1681 & n1703 ;
  assign n1705 = n1674 & n1704 ;
  assign n1706 = \InstAddrPointer_reg[31]/NET0131  & ~n1680 ;
  assign n1707 = ~\InstAddrPointer_reg[31]/NET0131  & n1680 ;
  assign n1708 = ~n1706 & ~n1707 ;
  assign n1710 = n1705 & ~n1708 ;
  assign n1709 = ~n1705 & n1708 ;
  assign n1711 = n930 & ~n1709 ;
  assign n1712 = ~n1710 & n1711 ;
  assign n1714 = ~n828 & ~n862 ;
  assign n1715 = n736 & ~n825 ;
  assign n1716 = n924 & ~n1715 ;
  assign n1717 = ~n872 & n1716 ;
  assign n1718 = ~n1714 & n1717 ;
  assign n1719 = n736 & n825 ;
  assign n1720 = READY_n_pad & n1719 ;
  assign n1721 = n1718 & ~n1720 ;
  assign n1722 = \InstAddrPointer_reg[31]/NET0131  & ~n1721 ;
  assign n1724 = n809 & ~n1708 ;
  assign n1713 = ~n780 & ~n1581 ;
  assign n1723 = ~n867 & ~n1403 ;
  assign n1725 = ~n1713 & ~n1723 ;
  assign n1726 = ~n1724 & n1725 ;
  assign n1727 = ~n1722 & n1726 ;
  assign n1728 = ~n1712 & n1727 ;
  assign n1729 = ~n1590 & n1728 ;
  assign n1730 = n948 & ~n1729 ;
  assign n1731 = n960 & n968 ;
  assign n1732 = \rEIP_reg[31]/NET0131  & n1731 ;
  assign n1733 = n960 & ~n968 ;
  assign n1734 = ~n951 & ~n970 ;
  assign n1735 = ~n955 & n1734 ;
  assign n1736 = ~n1733 & n1735 ;
  assign n1737 = \InstAddrPointer_reg[31]/NET0131  & ~n1736 ;
  assign n1738 = ~n1732 & ~n1737 ;
  assign n1739 = ~n1730 & n1738 ;
  assign n1740 = n1015 & n1423 ;
  assign n1741 = ~n1317 & n1740 ;
  assign n1742 = n1395 & n1741 ;
  assign n1743 = n1370 & n1742 ;
  assign n1744 = ~\InstAddrPointer_reg[30]/NET0131  & ~n1367 ;
  assign n1745 = \InstAddrPointer_reg[30]/NET0131  & n1367 ;
  assign n1746 = ~n1744 & ~n1745 ;
  assign n1747 = ~n1743 & ~n1746 ;
  assign n1748 = n1371 & n1742 ;
  assign n1749 = n1051 & ~n1748 ;
  assign n1750 = ~n1747 & n1749 ;
  assign n1751 = ~n1450 & ~n1470 ;
  assign n1752 = ~n1458 & n1751 ;
  assign n1753 = ~n1446 & n1466 ;
  assign n1754 = ~n1752 & n1753 ;
  assign n1755 = ~n1446 & n1469 ;
  assign n1756 = ~n1475 & ~n1755 ;
  assign n1757 = ~n1754 & n1756 ;
  assign n1758 = ~n1439 & ~n1443 ;
  assign n1759 = ~n1757 & n1758 ;
  assign n1760 = ~n1474 & ~n1489 ;
  assign n1761 = ~n1439 & ~n1760 ;
  assign n1762 = ~n1759 & ~n1761 ;
  assign n1763 = ~n1491 & n1762 ;
  assign n1764 = n1488 & n1501 ;
  assign n1765 = ~n1504 & n1764 ;
  assign n1766 = n1763 & n1765 ;
  assign n1767 = n1524 & ~n1529 ;
  assign n1768 = ~n1512 & n1767 ;
  assign n1769 = ~n1507 & n1536 ;
  assign n1770 = n1768 & n1769 ;
  assign n1771 = ~n1540 & n1554 ;
  assign n1772 = n1770 & n1771 ;
  assign n1773 = n1766 & n1772 ;
  assign n1774 = n1543 & n1575 ;
  assign n1775 = n1773 & n1774 ;
  assign n1776 = ~n1051 & ~n1563 ;
  assign n1777 = ~n1775 & n1776 ;
  assign n1778 = ~n1051 & n1577 ;
  assign n1779 = ~n1777 & ~n1778 ;
  assign n1780 = ~n1750 & n1779 ;
  assign n1781 = n921 & ~n1780 ;
  assign n1782 = \InstAddrPointer_reg[30]/NET0131  & ~n921 ;
  assign n1783 = ~n1781 & ~n1782 ;
  assign n1784 = n748 & ~n1783 ;
  assign n1785 = \InstAddrPointer_reg[9]/NET0131  & n1642 ;
  assign n1786 = ~n1622 & ~n1625 ;
  assign n1787 = ~n1604 & n1614 ;
  assign n1788 = ~n1786 & n1787 ;
  assign n1789 = ~n1624 & ~n1635 ;
  assign n1790 = ~n1604 & ~n1789 ;
  assign n1791 = ~n1788 & ~n1790 ;
  assign n1792 = ~n1607 & ~n1640 ;
  assign n1793 = ~n1791 & n1792 ;
  assign n1794 = n1634 & ~n1640 ;
  assign n1795 = ~n1633 & ~n1794 ;
  assign n1796 = ~n1793 & n1795 ;
  assign n1797 = n1785 & ~n1796 ;
  assign n1800 = \InstAddrPointer_reg[13]/NET0131  & n1653 ;
  assign n1801 = ~\InstAddrPointer_reg[14]/NET0131  & ~n1646 ;
  assign n1802 = ~n1659 & ~n1801 ;
  assign n1798 = ~\InstAddrPointer_reg[10]/NET0131  & ~n1596 ;
  assign n1799 = ~n1649 & ~n1798 ;
  assign n1803 = n1600 & n1799 ;
  assign n1804 = n1802 & n1803 ;
  assign n1805 = n1663 & n1804 ;
  assign n1806 = n1800 & n1805 ;
  assign n1807 = n1797 & n1806 ;
  assign n1808 = \InstAddrPointer_reg[18]/NET0131  & n1599 ;
  assign n1809 = ~\InstAddrPointer_reg[18]/NET0131  & ~n1599 ;
  assign n1810 = ~n1808 & ~n1809 ;
  assign n1811 = \InstAddrPointer_reg[19]/NET0131  & n1810 ;
  assign n1812 = n1673 & n1811 ;
  assign n1813 = n1807 & n1812 ;
  assign n1814 = n1703 & n1813 ;
  assign n1816 = n1681 & n1814 ;
  assign n1815 = ~n1681 & ~n1814 ;
  assign n1817 = n930 & ~n1815 ;
  assign n1818 = ~n1816 & n1817 ;
  assign n1819 = ~n780 & ~n1563 ;
  assign n1820 = n843 & ~n1720 ;
  assign n1821 = n1716 & n1820 ;
  assign n1822 = \InstAddrPointer_reg[30]/NET0131  & ~n1821 ;
  assign n1825 = ~n1819 & ~n1822 ;
  assign n1823 = n809 & n1681 ;
  assign n1824 = ~n839 & n1746 ;
  assign n1826 = ~n1823 & ~n1824 ;
  assign n1827 = n1825 & n1826 ;
  assign n1828 = ~n1818 & n1827 ;
  assign n1829 = ~n1784 & n1828 ;
  assign n1830 = n948 & ~n1829 ;
  assign n1831 = \rEIP_reg[30]/NET0131  & n1731 ;
  assign n1832 = \InstAddrPointer_reg[30]/NET0131  & ~n1736 ;
  assign n1833 = ~n1831 & ~n1832 ;
  assign n1834 = ~n1830 & n1833 ;
  assign n1835 = \InstAddrPointer_reg[28]/NET0131  & ~n921 ;
  assign n1846 = n1389 & n1740 ;
  assign n1847 = ~n1317 & n1846 ;
  assign n1848 = \InstAddrPointer_reg[23]/NET0131  & n1377 ;
  assign n1849 = n1393 & n1848 ;
  assign n1850 = n1847 & n1849 ;
  assign n1851 = n1345 & n1359 ;
  assign n1852 = n1850 & n1851 ;
  assign n1853 = \InstAddrPointer_reg[28]/NET0131  & ~n1344 ;
  assign n1854 = ~\InstAddrPointer_reg[28]/NET0131  & n1344 ;
  assign n1855 = ~n1853 & ~n1854 ;
  assign n1857 = n1852 & n1855 ;
  assign n1856 = ~n1852 & ~n1855 ;
  assign n1858 = n1051 & ~n1856 ;
  assign n1859 = ~n1857 & n1858 ;
  assign n1836 = n1488 & n1513 ;
  assign n1837 = ~n1491 & n1836 ;
  assign n1838 = n1762 & n1837 ;
  assign n1839 = n1767 & n1838 ;
  assign n1840 = n1556 & ~n1567 ;
  assign n1841 = n1839 & n1840 ;
  assign n1843 = n1570 & ~n1841 ;
  assign n1842 = ~n1570 & n1841 ;
  assign n1844 = ~n1051 & ~n1842 ;
  assign n1845 = ~n1843 & n1844 ;
  assign n1860 = n921 & ~n1845 ;
  assign n1861 = ~n1859 & n1860 ;
  assign n1862 = ~n1835 & ~n1861 ;
  assign n1863 = n748 & ~n1862 ;
  assign n1866 = \InstAddrPointer_reg[11]/NET0131  & n1785 ;
  assign n1867 = n1799 & n1866 ;
  assign n1868 = ~n1796 & n1867 ;
  assign n1864 = ~\InstAddrPointer_reg[12]/NET0131  & ~n1651 ;
  assign n1865 = ~n1645 & ~n1864 ;
  assign n1869 = n1332 & n1865 ;
  assign n1870 = n1868 & n1869 ;
  assign n1871 = ~\InstAddrPointer_reg[16]/NET0131  & ~n1661 ;
  assign n1872 = ~n1597 & ~n1871 ;
  assign n1873 = n1338 & n1872 ;
  assign n1874 = n1870 & n1873 ;
  assign n1875 = ~\InstAddrPointer_reg[27]/NET0131  & ~n1676 ;
  assign n1876 = ~n1682 & ~n1875 ;
  assign n1877 = n1673 & n1876 ;
  assign n1878 = n1698 & n1877 ;
  assign n1879 = n1874 & n1878 ;
  assign n1881 = ~n1684 & ~n1879 ;
  assign n1880 = n1684 & n1879 ;
  assign n1882 = n930 & ~n1880 ;
  assign n1883 = ~n1881 & n1882 ;
  assign n1888 = ~n828 & ~n895 ;
  assign n1889 = ~n825 & ~n836 ;
  assign n1890 = ~n923 & ~n1889 ;
  assign n1891 = ~n1888 & n1890 ;
  assign n1892 = ~n812 & n1891 ;
  assign n1893 = n828 & ~n864 ;
  assign n1894 = READY_n_pad & ~n1893 ;
  assign n1895 = n1892 & ~n1894 ;
  assign n1896 = \InstAddrPointer_reg[28]/NET0131  & ~n1895 ;
  assign n1885 = \InstAddrPointer_reg[28]/NET0131  & ~n828 ;
  assign n1886 = n839 & ~n1885 ;
  assign n1887 = ~n1855 & ~n1886 ;
  assign n1884 = n809 & n1684 ;
  assign n1897 = ~n780 & n1570 ;
  assign n1898 = ~n1884 & ~n1897 ;
  assign n1899 = ~n1887 & n1898 ;
  assign n1900 = ~n1896 & n1899 ;
  assign n1901 = ~n1883 & n1900 ;
  assign n1902 = ~n1863 & n1901 ;
  assign n1903 = n948 & ~n1902 ;
  assign n1904 = \rEIP_reg[28]/NET0131  & n1731 ;
  assign n1905 = \InstAddrPointer_reg[28]/NET0131  & ~n1736 ;
  assign n1906 = ~n1904 & ~n1905 ;
  assign n1907 = ~n1903 & n1906 ;
  assign n1908 = \InstAddrPointer_reg[23]/NET0131  & ~n921 ;
  assign n1909 = n1536 & ~n1550 ;
  assign n1910 = n1494 & n1509 ;
  assign n1911 = ~n1512 & n1910 ;
  assign n1912 = n1767 & n1911 ;
  assign n1913 = n1909 & n1912 ;
  assign n1914 = n1548 & ~n1913 ;
  assign n1915 = ~n1548 & n1909 ;
  assign n1916 = n1912 & n1915 ;
  assign n1917 = ~n1051 & ~n1916 ;
  assign n1918 = ~n1914 & n1917 ;
  assign n1919 = ~n1361 & ~n1426 ;
  assign n1920 = ~n1850 & ~n1919 ;
  assign n1921 = n1051 & ~n1920 ;
  assign n1922 = n921 & ~n1921 ;
  assign n1923 = ~n1918 & n1922 ;
  assign n1924 = ~n1908 & ~n1923 ;
  assign n1925 = n748 & ~n1924 ;
  assign n1930 = n1673 & n1874 ;
  assign n1931 = n1693 & n1930 ;
  assign n1926 = ~\InstAddrPointer_reg[23]/NET0131  & ~n1691 ;
  assign n1927 = ~n1675 & ~n1926 ;
  assign n1928 = n1674 & n1692 ;
  assign n1929 = ~n1927 & ~n1928 ;
  assign n1932 = n930 & ~n1929 ;
  assign n1933 = ~n1931 & n1932 ;
  assign n1935 = n873 & ~n923 ;
  assign n1936 = ~n1714 & n1935 ;
  assign n1937 = ~n812 & n1936 ;
  assign n1938 = ~n756 & ~n1691 ;
  assign n1939 = n1937 & ~n1938 ;
  assign n1940 = \InstAddrPointer_reg[23]/NET0131  & ~n1939 ;
  assign n1934 = ~n839 & n1361 ;
  assign n1941 = n809 & n1927 ;
  assign n1942 = ~n780 & n1548 ;
  assign n1943 = ~n1941 & ~n1942 ;
  assign n1944 = ~n1934 & n1943 ;
  assign n1945 = ~n1940 & n1944 ;
  assign n1946 = ~n1933 & n1945 ;
  assign n1947 = ~n1925 & n1946 ;
  assign n1948 = n948 & ~n1947 ;
  assign n1949 = \rEIP_reg[23]/NET0131  & n1731 ;
  assign n1950 = \InstAddrPointer_reg[23]/NET0131  & ~n1736 ;
  assign n1951 = ~n1949 & ~n1950 ;
  assign n1952 = ~n1948 & n1951 ;
  assign n1953 = n1362 & n1426 ;
  assign n1954 = ~n1345 & ~n1953 ;
  assign n1955 = n1051 & ~n1852 ;
  assign n1956 = ~n1954 & n1955 ;
  assign n1958 = n1558 & n1567 ;
  assign n1957 = ~n1558 & ~n1567 ;
  assign n1959 = ~n1051 & ~n1957 ;
  assign n1960 = ~n1958 & n1959 ;
  assign n1961 = ~n1956 & ~n1960 ;
  assign n1962 = n921 & ~n1961 ;
  assign n1963 = \InstAddrPointer_reg[27]/NET0131  & ~n921 ;
  assign n1964 = ~n1962 & ~n1963 ;
  assign n1965 = n748 & ~n1964 ;
  assign n1967 = n1674 & n1698 ;
  assign n1968 = ~n1876 & ~n1967 ;
  assign n1966 = n1668 & n1878 ;
  assign n1969 = n930 & ~n1966 ;
  assign n1970 = ~n1968 & n1969 ;
  assign n1972 = ~n756 & ~n1676 ;
  assign n1973 = n1718 & ~n1972 ;
  assign n1974 = \InstAddrPointer_reg[27]/NET0131  & ~n1973 ;
  assign n1975 = READY_n_pad & n736 ;
  assign n1976 = \InstAddrPointer_reg[27]/NET0131  & n1975 ;
  assign n1977 = ~READY_n_pad & n1345 ;
  assign n1978 = ~n837 & n1977 ;
  assign n1979 = ~n1976 & ~n1978 ;
  assign n1980 = n825 & ~n1979 ;
  assign n1982 = ~n780 & n1567 ;
  assign n1971 = n698 & n1345 ;
  assign n1981 = n809 & n1876 ;
  assign n1983 = ~n1971 & ~n1981 ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = ~n1980 & n1984 ;
  assign n1986 = ~n1974 & n1985 ;
  assign n1987 = ~n1970 & n1986 ;
  assign n1988 = ~n1965 & n1987 ;
  assign n1989 = n948 & ~n1988 ;
  assign n1990 = \rEIP_reg[27]/NET0131  & n1731 ;
  assign n1991 = \InstAddrPointer_reg[27]/NET0131  & ~n1736 ;
  assign n1992 = ~n1990 & ~n1991 ;
  assign n1993 = ~n1989 & n1992 ;
  assign n1994 = \PhyAddrPointer_reg[31]/NET0131  & ~n921 ;
  assign n1995 = ~n1588 & ~n1994 ;
  assign n1996 = n748 & ~n1995 ;
  assign n1997 = ~n749 & ~n923 ;
  assign n1998 = \PhyAddrPointer_reg[31]/NET0131  & ~n1997 ;
  assign n1999 = ~n1712 & ~n1998 ;
  assign n2000 = ~n1996 & n1999 ;
  assign n2001 = n948 & ~n2000 ;
  assign n2005 = \PhyAddrPointer_reg[2]/NET0131  & \PhyAddrPointer_reg[3]/NET0131  ;
  assign n2006 = \PhyAddrPointer_reg[4]/NET0131  & n2005 ;
  assign n2007 = \PhyAddrPointer_reg[5]/NET0131  & n2006 ;
  assign n2008 = \PhyAddrPointer_reg[6]/NET0131  & n2007 ;
  assign n2009 = \PhyAddrPointer_reg[7]/NET0131  & n2008 ;
  assign n2010 = \PhyAddrPointer_reg[8]/NET0131  & n2009 ;
  assign n2011 = \PhyAddrPointer_reg[9]/NET0131  & n2010 ;
  assign n2012 = \PhyAddrPointer_reg[10]/NET0131  & n2011 ;
  assign n2013 = \PhyAddrPointer_reg[11]/NET0131  & n2012 ;
  assign n2014 = \PhyAddrPointer_reg[12]/NET0131  & n2013 ;
  assign n2015 = \PhyAddrPointer_reg[13]/NET0131  & n2014 ;
  assign n2018 = \PhyAddrPointer_reg[14]/NET0131  & \PhyAddrPointer_reg[15]/NET0131  ;
  assign n2019 = \PhyAddrPointer_reg[16]/NET0131  & n2018 ;
  assign n2020 = \PhyAddrPointer_reg[17]/NET0131  & n2019 ;
  assign n2016 = \PhyAddrPointer_reg[18]/NET0131  & \PhyAddrPointer_reg[19]/NET0131  ;
  assign n2017 = \PhyAddrPointer_reg[20]/NET0131  & n2016 ;
  assign n2021 = \PhyAddrPointer_reg[21]/NET0131  & n2017 ;
  assign n2022 = n2020 & n2021 ;
  assign n2023 = n2015 & n2022 ;
  assign n2024 = \PhyAddrPointer_reg[22]/NET0131  & \PhyAddrPointer_reg[23]/NET0131  ;
  assign n2025 = n2023 & n2024 ;
  assign n2026 = \PhyAddrPointer_reg[24]/NET0131  & n2025 ;
  assign n2027 = \PhyAddrPointer_reg[25]/NET0131  & \PhyAddrPointer_reg[26]/NET0131  ;
  assign n2028 = n2026 & n2027 ;
  assign n2029 = \PhyAddrPointer_reg[27]/NET0131  & n2028 ;
  assign n2030 = \PhyAddrPointer_reg[28]/NET0131  & n2029 ;
  assign n2031 = \PhyAddrPointer_reg[29]/NET0131  & n2030 ;
  assign n2032 = \PhyAddrPointer_reg[30]/NET0131  & n2031 ;
  assign n2033 = \PhyAddrPointer_reg[1]/NET0131  & n2032 ;
  assign n2034 = ~\PhyAddrPointer_reg[31]/NET0131  & ~n2033 ;
  assign n2035 = \PhyAddrPointer_reg[31]/NET0131  & n2033 ;
  assign n2036 = ~n2034 & ~n2035 ;
  assign n2037 = ~n952 & ~n970 ;
  assign n2038 = \DataWidth_reg[1]/NET0131  & ~n970 ;
  assign n2039 = ~n2037 & ~n2038 ;
  assign n2040 = n2036 & n2039 ;
  assign n2042 = ~\PhyAddrPointer_reg[31]/NET0131  & ~n2032 ;
  assign n2041 = \PhyAddrPointer_reg[31]/NET0131  & n2032 ;
  assign n2043 = n971 & ~n2041 ;
  assign n2044 = ~n2042 & n2043 ;
  assign n2002 = ~n955 & ~n982 ;
  assign n2003 = ~n980 & n2002 ;
  assign n2004 = \PhyAddrPointer_reg[31]/NET0131  & ~n2003 ;
  assign n2045 = ~n1732 & ~n2004 ;
  assign n2046 = ~n2044 & n2045 ;
  assign n2047 = ~n2040 & n2046 ;
  assign n2048 = ~n2001 & n2047 ;
  assign n2049 = \InstAddrPointer_reg[19]/NET0131  & ~n921 ;
  assign n2050 = ~\InstAddrPointer_reg[19]/NET0131  & ~n1385 ;
  assign n2051 = ~n1339 & ~n2050 ;
  assign n2052 = n1384 & n1741 ;
  assign n2053 = n1387 & n2052 ;
  assign n2054 = ~n2051 & ~n2053 ;
  assign n2055 = n1051 & ~n1847 ;
  assign n2056 = ~n2054 & n2055 ;
  assign n2057 = ~n1526 & n1529 ;
  assign n2058 = ~n1912 & ~n2057 ;
  assign n2059 = ~n1051 & ~n2058 ;
  assign n2060 = ~n2056 & ~n2059 ;
  assign n2061 = n921 & ~n2060 ;
  assign n2062 = ~n2049 & ~n2061 ;
  assign n2063 = n748 & ~n2062 ;
  assign n2065 = ~\InstAddrPointer_reg[19]/NET0131  & ~n1808 ;
  assign n2066 = ~n1669 & ~n2065 ;
  assign n2067 = n1600 & n1666 ;
  assign n2068 = \InstAddrPointer_reg[18]/NET0131  & n2067 ;
  assign n2069 = ~n2066 & ~n2068 ;
  assign n2070 = n930 & ~n1668 ;
  assign n2071 = ~n2069 & n2070 ;
  assign n2073 = n845 & n924 ;
  assign n2074 = \InstAddrPointer_reg[19]/NET0131  & ~n2073 ;
  assign n2072 = ~n839 & n2051 ;
  assign n2064 = ~n780 & n1529 ;
  assign n2075 = n809 & n2066 ;
  assign n2076 = ~n2064 & ~n2075 ;
  assign n2077 = ~n2072 & n2076 ;
  assign n2078 = ~n2074 & n2077 ;
  assign n2079 = ~n2071 & n2078 ;
  assign n2080 = ~n2063 & n2079 ;
  assign n2081 = n948 & ~n2080 ;
  assign n2082 = \rEIP_reg[19]/NET0131  & n1731 ;
  assign n2083 = \InstAddrPointer_reg[19]/NET0131  & ~n1736 ;
  assign n2084 = ~n2082 & ~n2083 ;
  assign n2085 = ~n2081 & n2084 ;
  assign n2087 = \InstAddrPointer_reg[20]/NET0131  & ~n921 ;
  assign n2093 = ~n1535 & n1839 ;
  assign n2092 = n1535 & ~n1839 ;
  assign n2094 = ~n1051 & ~n2092 ;
  assign n2095 = ~n2093 & n2094 ;
  assign n2088 = n1392 & n1847 ;
  assign n2089 = ~n1392 & ~n1847 ;
  assign n2090 = ~n2088 & ~n2089 ;
  assign n2091 = n1051 & ~n2090 ;
  assign n2096 = n921 & ~n2091 ;
  assign n2097 = ~n2095 & n2096 ;
  assign n2098 = ~n2087 & ~n2097 ;
  assign n2099 = n748 & ~n2098 ;
  assign n2101 = n1672 & n1874 ;
  assign n2100 = ~n1672 & ~n1874 ;
  assign n2102 = n930 & ~n2100 ;
  assign n2103 = ~n2101 & n2102 ;
  assign n2106 = \InstAddrPointer_reg[20]/NET0131  & ~n836 ;
  assign n2107 = n867 & ~n2106 ;
  assign n2108 = n1392 & ~n2107 ;
  assign n2105 = \InstAddrPointer_reg[20]/NET0131  & ~n1937 ;
  assign n2086 = n809 & n1672 ;
  assign n2104 = ~n780 & n1535 ;
  assign n2109 = ~n2086 & ~n2104 ;
  assign n2110 = ~n2105 & n2109 ;
  assign n2111 = ~n2108 & n2110 ;
  assign n2112 = ~n2103 & n2111 ;
  assign n2113 = ~n2099 & n2112 ;
  assign n2114 = n948 & ~n2113 ;
  assign n2115 = \rEIP_reg[20]/NET0131  & n1731 ;
  assign n2116 = \InstAddrPointer_reg[20]/NET0131  & ~n1736 ;
  assign n2117 = ~n2115 & ~n2116 ;
  assign n2118 = ~n2114 & n2117 ;
  assign n2119 = \InstAddrPointer_reg[22]/NET0131  & ~n921 ;
  assign n2125 = n1393 & n1847 ;
  assign n2126 = ~n1377 & ~n2125 ;
  assign n2127 = ~n1742 & ~n2126 ;
  assign n2128 = n1051 & ~n2127 ;
  assign n2120 = n1766 & n1770 ;
  assign n2122 = n1550 & ~n2120 ;
  assign n2121 = ~n1550 & n2120 ;
  assign n2123 = ~n1051 & ~n2121 ;
  assign n2124 = ~n2122 & n2123 ;
  assign n2129 = n921 & ~n2124 ;
  assign n2130 = ~n2128 & n2129 ;
  assign n2131 = ~n2119 & ~n2130 ;
  assign n2132 = n748 & ~n2131 ;
  assign n2135 = n1692 & n1813 ;
  assign n2134 = ~n1692 & ~n1813 ;
  assign n2136 = n930 & ~n2134 ;
  assign n2137 = ~n2135 & n2136 ;
  assign n2138 = ~n736 & ~n834 ;
  assign n2139 = n825 & ~n2138 ;
  assign n2140 = READY_n_pad & n2139 ;
  assign n2141 = n1717 & ~n1888 ;
  assign n2142 = ~n2140 & n2141 ;
  assign n2143 = \InstAddrPointer_reg[22]/NET0131  & ~n2142 ;
  assign n2144 = ~n839 & n1377 ;
  assign n2133 = ~n780 & n1550 ;
  assign n2145 = n809 & n1692 ;
  assign n2146 = ~n2133 & ~n2145 ;
  assign n2147 = ~n2144 & n2146 ;
  assign n2148 = ~n2143 & n2147 ;
  assign n2149 = ~n2137 & n2148 ;
  assign n2150 = ~n2132 & n2149 ;
  assign n2151 = n948 & ~n2150 ;
  assign n2152 = \rEIP_reg[22]/NET0131  & n1731 ;
  assign n2153 = \InstAddrPointer_reg[22]/NET0131  & ~n1736 ;
  assign n2154 = ~n2152 & ~n2153 ;
  assign n2155 = ~n2151 & n2154 ;
  assign n2181 = ~n1695 & ~n1931 ;
  assign n2182 = n1696 & n1930 ;
  assign n2183 = n930 & ~n2182 ;
  assign n2184 = ~n2181 & n2183 ;
  assign n2156 = \InstAddrPointer_reg[24]/NET0131  & ~n921 ;
  assign n2173 = ~n1358 & ~n1850 ;
  assign n2174 = n1358 & n1850 ;
  assign n2175 = ~n2173 & ~n2174 ;
  assign n2176 = n1051 & ~n2175 ;
  assign n2157 = n1839 & n1915 ;
  assign n2158 = n1552 & ~n2157 ;
  assign n2160 = ~n1467 & n1472 ;
  assign n2161 = ~n1439 & n1447 ;
  assign n2162 = ~n2160 & n2161 ;
  assign n2159 = ~n1439 & ~n1477 ;
  assign n2163 = n1492 & ~n2159 ;
  assign n2164 = ~n2162 & n2163 ;
  assign n2165 = n1764 & n2164 ;
  assign n2166 = n1508 & ~n1535 ;
  assign n2167 = n1768 & n2166 ;
  assign n2168 = n2165 & n2167 ;
  assign n2169 = ~n1533 & n1554 ;
  assign n2170 = n2168 & n2169 ;
  assign n2171 = ~n1051 & ~n2170 ;
  assign n2172 = ~n2158 & n2171 ;
  assign n2177 = n921 & ~n2172 ;
  assign n2178 = ~n2176 & n2177 ;
  assign n2179 = ~n2156 & ~n2178 ;
  assign n2180 = n748 & ~n2179 ;
  assign n2188 = \InstAddrPointer_reg[24]/NET0131  & ~n1937 ;
  assign n2187 = ~n867 & n1358 ;
  assign n2185 = ~n780 & n1552 ;
  assign n2186 = n809 & n1695 ;
  assign n2189 = ~n2185 & ~n2186 ;
  assign n2190 = ~n2187 & n2189 ;
  assign n2191 = ~n2188 & n2190 ;
  assign n2192 = ~n2180 & n2191 ;
  assign n2193 = ~n2184 & n2192 ;
  assign n2194 = n948 & ~n2193 ;
  assign n2195 = \rEIP_reg[24]/NET0131  & n1731 ;
  assign n2196 = \InstAddrPointer_reg[24]/NET0131  & ~n1736 ;
  assign n2197 = ~n2195 & ~n2196 ;
  assign n2198 = ~n2194 & n2197 ;
  assign n2199 = \PhyAddrPointer_reg[30]/NET0131  & ~n921 ;
  assign n2200 = ~n1781 & ~n2199 ;
  assign n2201 = n748 & ~n2200 ;
  assign n2202 = \PhyAddrPointer_reg[30]/NET0131  & ~n1997 ;
  assign n2203 = ~n1818 & ~n2202 ;
  assign n2204 = ~n2201 & n2203 ;
  assign n2205 = n948 & ~n2204 ;
  assign n2209 = \PhyAddrPointer_reg[1]/NET0131  & n2031 ;
  assign n2210 = ~\PhyAddrPointer_reg[30]/NET0131  & ~n2209 ;
  assign n2211 = ~n2033 & ~n2210 ;
  assign n2212 = n2039 & n2211 ;
  assign n2206 = ~\PhyAddrPointer_reg[30]/NET0131  & ~n2031 ;
  assign n2207 = n971 & ~n2032 ;
  assign n2208 = ~n2206 & n2207 ;
  assign n2213 = \PhyAddrPointer_reg[30]/NET0131  & ~n2003 ;
  assign n2214 = ~n1831 & ~n2213 ;
  assign n2215 = ~n2208 & n2214 ;
  assign n2216 = ~n2212 & n2215 ;
  assign n2217 = ~n2205 & n2216 ;
  assign n2221 = \InstAddrPointer_reg[11]/NET0131  & ~n921 ;
  assign n2226 = ~n1011 & ~n1422 ;
  assign n2227 = n1011 & n1422 ;
  assign n2228 = ~n2226 & ~n2227 ;
  assign n2229 = n1051 & ~n2228 ;
  assign n2223 = ~n1494 & n1500 ;
  assign n2222 = n1494 & ~n1500 ;
  assign n2224 = ~n1051 & ~n2222 ;
  assign n2225 = ~n2223 & n2224 ;
  assign n2230 = n921 & ~n2225 ;
  assign n2231 = ~n2229 & n2230 ;
  assign n2232 = ~n2221 & ~n2231 ;
  assign n2233 = n748 & ~n2232 ;
  assign n2243 = n1644 & n1658 ;
  assign n2245 = n1652 & n2243 ;
  assign n2244 = ~n1652 & ~n2243 ;
  assign n2246 = n930 & ~n2244 ;
  assign n2247 = ~n2245 & n2246 ;
  assign n2234 = n833 & n836 ;
  assign n2235 = n826 & ~n2234 ;
  assign n2236 = n1011 & n2235 ;
  assign n2237 = n862 & n1007 ;
  assign n2238 = \InstAddrPointer_reg[11]/NET0131  & ~n2237 ;
  assign n2239 = ~n2236 & ~n2238 ;
  assign n2240 = ~n836 & n1011 ;
  assign n2241 = n874 & ~n2240 ;
  assign n2242 = ~n2239 & ~n2241 ;
  assign n2220 = ~n780 & n1500 ;
  assign n2249 = n808 & ~n1652 ;
  assign n2248 = ~\InstAddrPointer_reg[11]/NET0131  & ~n808 ;
  assign n2250 = ~n756 & ~n2248 ;
  assign n2251 = ~n2249 & n2250 ;
  assign n2252 = \InstAddrPointer_reg[11]/NET0131  & n923 ;
  assign n2253 = n698 & n1011 ;
  assign n2254 = ~n2252 & ~n2253 ;
  assign n2255 = ~n2251 & n2254 ;
  assign n2256 = ~n2220 & n2255 ;
  assign n2257 = ~n2242 & n2256 ;
  assign n2258 = ~n2247 & n2257 ;
  assign n2259 = ~n2233 & n2258 ;
  assign n2260 = n948 & ~n2259 ;
  assign n2218 = \rEIP_reg[11]/NET0131  & n1731 ;
  assign n2219 = \InstAddrPointer_reg[11]/NET0131  & ~n1736 ;
  assign n2261 = ~n2218 & ~n2219 ;
  assign n2262 = ~n2260 & n2261 ;
  assign n2264 = \InstAddrPointer_reg[14]/NET0131  & ~n921 ;
  assign n2265 = n1507 & ~n1766 ;
  assign n2266 = ~n1910 & ~n2265 ;
  assign n2267 = ~n1051 & ~n2266 ;
  assign n2268 = ~n1318 & ~n1325 ;
  assign n2269 = n1051 & ~n1326 ;
  assign n2270 = ~n2268 & n2269 ;
  assign n2271 = ~n2267 & ~n2270 ;
  assign n2272 = n921 & ~n2271 ;
  assign n2273 = ~n2264 & ~n2272 ;
  assign n2274 = n748 & ~n2273 ;
  assign n2275 = n1642 & ~n1796 ;
  assign n2276 = n1658 & n2275 ;
  assign n2277 = n1800 & n2276 ;
  assign n2279 = n1802 & n2277 ;
  assign n2278 = ~n1802 & ~n2277 ;
  assign n2280 = n930 & ~n2278 ;
  assign n2281 = ~n2279 & n2280 ;
  assign n2284 = \InstAddrPointer_reg[14]/NET0131  & ~n1937 ;
  assign n2283 = ~n867 & n1325 ;
  assign n2263 = ~n780 & n1507 ;
  assign n2282 = n809 & n1802 ;
  assign n2285 = ~n2263 & ~n2282 ;
  assign n2286 = ~n2283 & n2285 ;
  assign n2287 = ~n2284 & n2286 ;
  assign n2288 = ~n2281 & n2287 ;
  assign n2289 = ~n2274 & n2288 ;
  assign n2290 = n948 & ~n2289 ;
  assign n2291 = \rEIP_reg[14]/NET0131  & n1731 ;
  assign n2292 = \InstAddrPointer_reg[14]/NET0131  & ~n1736 ;
  assign n2293 = ~n2291 & ~n2292 ;
  assign n2294 = ~n2290 & n2293 ;
  assign n2295 = \InstAddrPointer_reg[25]/NET0131  & ~n921 ;
  assign n2296 = n1358 & n1848 ;
  assign n2297 = ~\InstAddrPointer_reg[21]/NET0131  & ~n1390 ;
  assign n2298 = ~n1375 & ~n2297 ;
  assign n2299 = n2296 & n2298 ;
  assign n2300 = ~n1380 & n1421 ;
  assign n2301 = n1424 & n2300 ;
  assign n2302 = n1418 & n2301 ;
  assign n2303 = \InstAddrPointer_reg[20]/NET0131  & n1383 ;
  assign n2304 = n1388 & n2303 ;
  assign n2305 = n2302 & n2304 ;
  assign n2306 = n2299 & n2305 ;
  assign n2307 = ~n1355 & ~n2306 ;
  assign n2308 = \InstAddrPointer_reg[25]/NET0131  & n2296 ;
  assign n2309 = n2125 & n2308 ;
  assign n2310 = ~n2307 & ~n2309 ;
  assign n2311 = n1051 & ~n2310 ;
  assign n2313 = n1540 & ~n2170 ;
  assign n2312 = ~n1540 & n2170 ;
  assign n2314 = ~n1051 & ~n2312 ;
  assign n2315 = ~n2313 & n2314 ;
  assign n2316 = n921 & ~n2315 ;
  assign n2317 = ~n2311 & n2316 ;
  assign n2318 = ~n2295 & ~n2317 ;
  assign n2319 = n748 & ~n2318 ;
  assign n2320 = n1674 & n1696 ;
  assign n2321 = ~\InstAddrPointer_reg[25]/NET0131  & ~n1685 ;
  assign n2322 = ~n1686 & ~n2321 ;
  assign n2324 = n2320 & n2322 ;
  assign n2323 = ~n2320 & ~n2322 ;
  assign n2325 = n930 & ~n2323 ;
  assign n2326 = ~n2324 & n2325 ;
  assign n2334 = \InstAddrPointer_reg[25]/NET0131  & ~n2142 ;
  assign n2328 = ~READY_n_pad & n2139 ;
  assign n2327 = n826 & n835 ;
  assign n2329 = ~n698 & ~n2327 ;
  assign n2330 = ~n2328 & n2329 ;
  assign n2331 = n1355 & ~n2330 ;
  assign n2332 = ~n780 & n1540 ;
  assign n2333 = n809 & n2322 ;
  assign n2335 = ~n2332 & ~n2333 ;
  assign n2336 = ~n2331 & n2335 ;
  assign n2337 = ~n2334 & n2336 ;
  assign n2338 = ~n2326 & n2337 ;
  assign n2339 = ~n2319 & n2338 ;
  assign n2340 = n948 & ~n2339 ;
  assign n2341 = \rEIP_reg[25]/NET0131  & n1731 ;
  assign n2342 = \InstAddrPointer_reg[25]/NET0131  & ~n1736 ;
  assign n2343 = ~n2341 & ~n2342 ;
  assign n2344 = ~n2340 & n2343 ;
  assign n2345 = \PhyAddrPointer_reg[15]/NET0131  & ~n921 ;
  assign n2349 = ~n1326 & ~n1374 ;
  assign n2350 = ~n1741 & ~n2349 ;
  assign n2351 = n1051 & ~n2350 ;
  assign n2346 = n1512 & ~n1910 ;
  assign n2347 = ~n1051 & ~n1911 ;
  assign n2348 = ~n2346 & n2347 ;
  assign n2352 = n921 & ~n2348 ;
  assign n2353 = ~n2351 & n2352 ;
  assign n2354 = ~n2345 & ~n2353 ;
  assign n2355 = n748 & ~n2354 ;
  assign n2356 = \PhyAddrPointer_reg[15]/NET0131  & ~n1997 ;
  assign n2357 = n1655 & n2243 ;
  assign n2359 = n1662 & n2357 ;
  assign n2358 = ~n1662 & ~n2357 ;
  assign n2360 = n930 & ~n2358 ;
  assign n2361 = ~n2359 & n2360 ;
  assign n2362 = ~n2356 & ~n2361 ;
  assign n2363 = ~n2355 & n2362 ;
  assign n2364 = n948 & ~n2363 ;
  assign n2372 = \PhyAddrPointer_reg[1]/NET0131  & n2013 ;
  assign n2373 = \PhyAddrPointer_reg[12]/NET0131  & n2372 ;
  assign n2374 = \PhyAddrPointer_reg[13]/NET0131  & n2373 ;
  assign n2375 = \PhyAddrPointer_reg[14]/NET0131  & n2374 ;
  assign n2376 = ~\PhyAddrPointer_reg[15]/NET0131  & ~n2375 ;
  assign n2377 = n2018 & n2374 ;
  assign n2378 = ~n2376 & ~n2377 ;
  assign n2379 = n970 & n2378 ;
  assign n2365 = \PhyAddrPointer_reg[14]/NET0131  & n2015 ;
  assign n2366 = ~\DataWidth_reg[1]/NET0131  & ~\PhyAddrPointer_reg[1]/NET0131  ;
  assign n2367 = n2365 & ~n2366 ;
  assign n2369 = \PhyAddrPointer_reg[15]/NET0131  & n2367 ;
  assign n2368 = ~\PhyAddrPointer_reg[15]/NET0131  & ~n2367 ;
  assign n2370 = n952 & ~n2368 ;
  assign n2371 = ~n2369 & n2370 ;
  assign n2380 = \rEIP_reg[15]/NET0131  & n1731 ;
  assign n2381 = \PhyAddrPointer_reg[15]/NET0131  & ~n2003 ;
  assign n2382 = ~n2380 & ~n2381 ;
  assign n2383 = ~n2371 & n2382 ;
  assign n2384 = ~n2379 & n2383 ;
  assign n2385 = ~n2364 & n2384 ;
  assign n2386 = \PhyAddrPointer_reg[23]/NET0131  & ~n921 ;
  assign n2387 = ~n1923 & ~n2386 ;
  assign n2388 = n748 & ~n2387 ;
  assign n2389 = \PhyAddrPointer_reg[23]/NET0131  & ~n1997 ;
  assign n2390 = ~n1933 & ~n2389 ;
  assign n2391 = ~n2388 & n2390 ;
  assign n2392 = n948 & ~n2391 ;
  assign n2393 = \PhyAddrPointer_reg[1]/NET0131  & n2023 ;
  assign n2394 = \PhyAddrPointer_reg[22]/NET0131  & n2393 ;
  assign n2395 = ~\PhyAddrPointer_reg[23]/NET0131  & ~n2394 ;
  assign n2396 = \PhyAddrPointer_reg[1]/NET0131  & n2025 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = n2039 & n2397 ;
  assign n2399 = n971 & ~n2025 ;
  assign n2400 = n2003 & ~n2399 ;
  assign n2401 = \PhyAddrPointer_reg[23]/NET0131  & ~n2400 ;
  assign n2402 = \PhyAddrPointer_reg[22]/NET0131  & n2023 ;
  assign n2403 = n2399 & n2402 ;
  assign n2404 = ~n1949 & ~n2403 ;
  assign n2405 = ~n2401 & n2404 ;
  assign n2406 = ~n2398 & n2405 ;
  assign n2407 = ~n2392 & n2406 ;
  assign n2408 = \PhyAddrPointer_reg[27]/NET0131  & ~n921 ;
  assign n2409 = ~n1962 & ~n2408 ;
  assign n2410 = n748 & ~n2409 ;
  assign n2411 = \PhyAddrPointer_reg[27]/NET0131  & ~n1997 ;
  assign n2412 = ~n1970 & ~n2411 ;
  assign n2413 = ~n2410 & n2412 ;
  assign n2414 = n948 & ~n2413 ;
  assign n2418 = \PhyAddrPointer_reg[1]/NET0131  & n2029 ;
  assign n2419 = \PhyAddrPointer_reg[1]/NET0131  & n2026 ;
  assign n2420 = n2027 & n2419 ;
  assign n2421 = ~\PhyAddrPointer_reg[27]/NET0131  & ~n2420 ;
  assign n2422 = ~n2418 & ~n2421 ;
  assign n2423 = n2039 & n2422 ;
  assign n2415 = ~\PhyAddrPointer_reg[27]/NET0131  & ~n2028 ;
  assign n2416 = n971 & ~n2029 ;
  assign n2417 = ~n2415 & n2416 ;
  assign n2424 = \PhyAddrPointer_reg[27]/NET0131  & ~n2003 ;
  assign n2425 = ~n1990 & ~n2424 ;
  assign n2426 = ~n2417 & n2425 ;
  assign n2427 = ~n2423 & n2426 ;
  assign n2428 = ~n2414 & n2427 ;
  assign n2429 = \PhyAddrPointer_reg[28]/NET0131  & ~n921 ;
  assign n2430 = ~n1861 & ~n2429 ;
  assign n2431 = n748 & ~n2430 ;
  assign n2432 = \PhyAddrPointer_reg[28]/NET0131  & ~n1997 ;
  assign n2433 = ~n1883 & ~n2432 ;
  assign n2434 = ~n2431 & n2433 ;
  assign n2435 = n948 & ~n2434 ;
  assign n2439 = ~\PhyAddrPointer_reg[28]/NET0131  & ~n2418 ;
  assign n2440 = \PhyAddrPointer_reg[1]/NET0131  & n2030 ;
  assign n2441 = ~n2439 & ~n2440 ;
  assign n2442 = n2039 & n2441 ;
  assign n2436 = ~\PhyAddrPointer_reg[28]/NET0131  & ~n2029 ;
  assign n2437 = n971 & ~n2030 ;
  assign n2438 = ~n2436 & n2437 ;
  assign n2443 = \PhyAddrPointer_reg[28]/NET0131  & ~n2003 ;
  assign n2444 = ~n1904 & ~n2443 ;
  assign n2445 = ~n2438 & n2444 ;
  assign n2446 = ~n2442 & n2445 ;
  assign n2447 = ~n2435 & n2446 ;
  assign n2448 = \PhyAddrPointer_reg[29]/NET0131  & ~n921 ;
  assign n2449 = n1346 & n1356 ;
  assign n2450 = n2299 & n2449 ;
  assign n2451 = n2088 & n2450 ;
  assign n2452 = ~n1368 & ~n2451 ;
  assign n2453 = n1368 & n2450 ;
  assign n2454 = n2088 & n2453 ;
  assign n2455 = n1051 & ~n2454 ;
  assign n2456 = ~n2452 & n2455 ;
  assign n2457 = n1544 & n1571 ;
  assign n2458 = n2170 & n2457 ;
  assign n2459 = ~n1051 & ~n1574 ;
  assign n2460 = ~n2458 & n2459 ;
  assign n2461 = ~n1051 & n1574 ;
  assign n2462 = n2458 & n2461 ;
  assign n2463 = ~n2460 & ~n2462 ;
  assign n2464 = ~n2456 & n2463 ;
  assign n2465 = n921 & ~n2464 ;
  assign n2466 = ~n2448 & ~n2465 ;
  assign n2467 = n748 & ~n2466 ;
  assign n2468 = \PhyAddrPointer_reg[29]/NET0131  & ~n1997 ;
  assign n2469 = n1684 & n1966 ;
  assign n2471 = ~n1700 & ~n2469 ;
  assign n2470 = \InstAddrPointer_reg[29]/NET0131  & n2469 ;
  assign n2472 = n930 & ~n2470 ;
  assign n2473 = ~n2471 & n2472 ;
  assign n2474 = ~n2468 & ~n2473 ;
  assign n2475 = ~n2467 & n2474 ;
  assign n2476 = n948 & ~n2475 ;
  assign n2482 = ~\PhyAddrPointer_reg[29]/NET0131  & ~n2440 ;
  assign n2483 = ~n2209 & ~n2482 ;
  assign n2484 = n970 & n2483 ;
  assign n2477 = n2030 & ~n2366 ;
  assign n2479 = \PhyAddrPointer_reg[29]/NET0131  & n2477 ;
  assign n2478 = ~\PhyAddrPointer_reg[29]/NET0131  & ~n2477 ;
  assign n2480 = n952 & ~n2478 ;
  assign n2481 = ~n2479 & n2480 ;
  assign n2485 = \rEIP_reg[29]/NET0131  & n1731 ;
  assign n2486 = \PhyAddrPointer_reg[29]/NET0131  & ~n2003 ;
  assign n2487 = ~n2485 & ~n2486 ;
  assign n2488 = ~n2481 & n2487 ;
  assign n2489 = ~n2484 & n2488 ;
  assign n2490 = ~n2476 & n2489 ;
  assign n2494 = \InstAddrPointer_reg[8]/NET0131  & ~n921 ;
  assign n2499 = n1004 & n1317 ;
  assign n2498 = ~n1004 & ~n1317 ;
  assign n2500 = n1051 & ~n2498 ;
  assign n2501 = ~n2499 & n2500 ;
  assign n2495 = n1491 & ~n1762 ;
  assign n2496 = ~n1051 & ~n1763 ;
  assign n2497 = ~n2495 & n2496 ;
  assign n2502 = n921 & ~n2497 ;
  assign n2503 = ~n2501 & n2502 ;
  assign n2504 = ~n2494 & ~n2503 ;
  assign n2505 = n748 & ~n2504 ;
  assign n2510 = ~n1642 & n1796 ;
  assign n2511 = n930 & ~n2275 ;
  assign n2512 = ~n2510 & n2511 ;
  assign n2506 = n825 & ~n837 ;
  assign n2507 = READY_n_pad & n2506 ;
  assign n2508 = n1892 & ~n2507 ;
  assign n2509 = \InstAddrPointer_reg[8]/NET0131  & ~n2508 ;
  assign n2513 = ~n839 & n1004 ;
  assign n2493 = ~n780 & n1491 ;
  assign n2514 = n809 & n1642 ;
  assign n2515 = ~n2493 & ~n2514 ;
  assign n2516 = ~n2513 & n2515 ;
  assign n2517 = ~n2509 & n2516 ;
  assign n2518 = ~n2512 & n2517 ;
  assign n2519 = ~n2505 & n2518 ;
  assign n2520 = n948 & ~n2519 ;
  assign n2491 = \InstAddrPointer_reg[8]/NET0131  & ~n1736 ;
  assign n2492 = \rEIP_reg[8]/NET0131  & n1731 ;
  assign n2521 = ~n2491 & ~n2492 ;
  assign n2522 = ~n2520 & n2521 ;
  assign n2523 = \InstAddrPointer_reg[12]/NET0131  & ~n921 ;
  assign n2531 = ~\InstAddrPointer_reg[12]/NET0131  & ~n1010 ;
  assign n2532 = ~n1321 & ~n2531 ;
  assign n2533 = n1005 & ~n1317 ;
  assign n2534 = ~\InstAddrPointer_reg[10]/NET0131  & ~n1006 ;
  assign n2535 = ~n1007 & ~n2534 ;
  assign n2536 = n2533 & n2535 ;
  assign n2537 = \InstAddrPointer_reg[11]/NET0131  & n2536 ;
  assign n2539 = ~n2532 & n2537 ;
  assign n2538 = n2532 & ~n2537 ;
  assign n2540 = n1051 & ~n2538 ;
  assign n2541 = ~n2539 & n2540 ;
  assign n2525 = ~n1487 & n1763 ;
  assign n2526 = ~n1484 & ~n1500 ;
  assign n2527 = n2525 & n2526 ;
  assign n2528 = n1498 & ~n2527 ;
  assign n2524 = n1763 & n1764 ;
  assign n2529 = ~n1051 & ~n2524 ;
  assign n2530 = ~n2528 & n2529 ;
  assign n2542 = n921 & ~n2530 ;
  assign n2543 = ~n2541 & n2542 ;
  assign n2544 = ~n2523 & ~n2543 ;
  assign n2545 = n748 & ~n2544 ;
  assign n2548 = n1865 & n1868 ;
  assign n2547 = ~n1865 & ~n1868 ;
  assign n2549 = n930 & ~n2547 ;
  assign n2550 = ~n2548 & n2549 ;
  assign n2552 = \InstAddrPointer_reg[12]/NET0131  & ~n836 ;
  assign n2553 = n867 & ~n2552 ;
  assign n2554 = n2532 & ~n2553 ;
  assign n2551 = ~n780 & n1498 ;
  assign n2546 = \InstAddrPointer_reg[12]/NET0131  & ~n1936 ;
  assign n2556 = n808 & ~n1865 ;
  assign n2555 = ~\InstAddrPointer_reg[12]/NET0131  & ~n808 ;
  assign n2557 = ~n756 & ~n2555 ;
  assign n2558 = ~n2556 & n2557 ;
  assign n2559 = ~n2546 & ~n2558 ;
  assign n2560 = ~n2551 & n2559 ;
  assign n2561 = ~n2554 & n2560 ;
  assign n2562 = ~n2550 & n2561 ;
  assign n2563 = ~n2545 & n2562 ;
  assign n2564 = n948 & ~n2563 ;
  assign n2565 = \rEIP_reg[12]/NET0131  & n1731 ;
  assign n2566 = \InstAddrPointer_reg[12]/NET0131  & ~n1736 ;
  assign n2567 = ~n2565 & ~n2566 ;
  assign n2568 = ~n2564 & n2567 ;
  assign n2569 = \PhyAddrPointer_reg[11]/NET0131  & ~n921 ;
  assign n2570 = ~n2231 & ~n2569 ;
  assign n2571 = n748 & ~n2570 ;
  assign n2572 = \PhyAddrPointer_reg[11]/NET0131  & ~n1997 ;
  assign n2573 = ~n2247 & ~n2572 ;
  assign n2574 = ~n2571 & n2573 ;
  assign n2575 = n948 & ~n2574 ;
  assign n2579 = \PhyAddrPointer_reg[1]/NET0131  & n2012 ;
  assign n2580 = ~\PhyAddrPointer_reg[11]/NET0131  & ~n2579 ;
  assign n2581 = ~n2372 & ~n2580 ;
  assign n2582 = n2039 & n2581 ;
  assign n2576 = ~\PhyAddrPointer_reg[11]/NET0131  & ~n2012 ;
  assign n2577 = n971 & ~n2013 ;
  assign n2578 = ~n2576 & n2577 ;
  assign n2583 = \PhyAddrPointer_reg[11]/NET0131  & ~n2003 ;
  assign n2584 = ~n2218 & ~n2583 ;
  assign n2585 = ~n2578 & n2584 ;
  assign n2586 = ~n2582 & n2585 ;
  assign n2587 = ~n2575 & n2586 ;
  assign n2588 = \PhyAddrPointer_reg[14]/NET0131  & ~n921 ;
  assign n2589 = ~n2272 & ~n2588 ;
  assign n2590 = n748 & ~n2589 ;
  assign n2591 = \PhyAddrPointer_reg[14]/NET0131  & ~n1997 ;
  assign n2592 = ~n2281 & ~n2591 ;
  assign n2593 = ~n2590 & n2592 ;
  assign n2594 = n948 & ~n2593 ;
  assign n2598 = ~\PhyAddrPointer_reg[14]/NET0131  & ~n2374 ;
  assign n2599 = ~n2375 & ~n2598 ;
  assign n2600 = n2039 & n2599 ;
  assign n2595 = ~\PhyAddrPointer_reg[14]/NET0131  & ~n2015 ;
  assign n2596 = n971 & ~n2365 ;
  assign n2597 = ~n2595 & n2596 ;
  assign n2601 = \PhyAddrPointer_reg[14]/NET0131  & ~n2003 ;
  assign n2602 = ~n2291 & ~n2601 ;
  assign n2603 = ~n2597 & n2602 ;
  assign n2604 = ~n2600 & n2603 ;
  assign n2605 = ~n2594 & n2604 ;
  assign n2606 = \PhyAddrPointer_reg[19]/NET0131  & ~n921 ;
  assign n2607 = ~n2061 & ~n2606 ;
  assign n2608 = n748 & ~n2607 ;
  assign n2609 = \PhyAddrPointer_reg[19]/NET0131  & ~n1997 ;
  assign n2610 = ~n2071 & ~n2609 ;
  assign n2611 = ~n2608 & n2610 ;
  assign n2612 = n948 & ~n2611 ;
  assign n2613 = n2015 & n2020 ;
  assign n2614 = \PhyAddrPointer_reg[18]/NET0131  & n2613 ;
  assign n2620 = \PhyAddrPointer_reg[1]/NET0131  & n2614 ;
  assign n2621 = ~\PhyAddrPointer_reg[19]/NET0131  & ~n2620 ;
  assign n2622 = \PhyAddrPointer_reg[19]/NET0131  & n2620 ;
  assign n2623 = ~n2621 & ~n2622 ;
  assign n2624 = n2039 & n2623 ;
  assign n2615 = n971 & ~n2614 ;
  assign n2616 = n2003 & ~n2615 ;
  assign n2617 = \PhyAddrPointer_reg[19]/NET0131  & ~n2616 ;
  assign n2618 = ~\PhyAddrPointer_reg[19]/NET0131  & n971 ;
  assign n2619 = n2614 & n2618 ;
  assign n2625 = ~n2082 & ~n2619 ;
  assign n2626 = ~n2617 & n2625 ;
  assign n2627 = ~n2624 & n2626 ;
  assign n2628 = ~n2612 & n2627 ;
  assign n2629 = \PhyAddrPointer_reg[20]/NET0131  & ~n921 ;
  assign n2630 = ~n2097 & ~n2629 ;
  assign n2631 = n748 & ~n2630 ;
  assign n2632 = \PhyAddrPointer_reg[20]/NET0131  & ~n1997 ;
  assign n2633 = ~n2103 & ~n2632 ;
  assign n2634 = ~n2631 & n2633 ;
  assign n2635 = n948 & ~n2634 ;
  assign n2637 = ~\PhyAddrPointer_reg[20]/NET0131  & ~n2622 ;
  assign n2638 = n2017 & n2613 ;
  assign n2639 = \PhyAddrPointer_reg[1]/NET0131  & n2638 ;
  assign n2640 = ~n2637 & ~n2639 ;
  assign n2641 = n970 & n2640 ;
  assign n2643 = \PhyAddrPointer_reg[19]/NET0131  & ~n2366 ;
  assign n2644 = n2614 & n2643 ;
  assign n2645 = ~\PhyAddrPointer_reg[20]/NET0131  & ~n2644 ;
  assign n2642 = ~n2366 & n2638 ;
  assign n2646 = n952 & ~n2642 ;
  assign n2647 = ~n2645 & n2646 ;
  assign n2636 = \PhyAddrPointer_reg[20]/NET0131  & ~n2003 ;
  assign n2648 = ~n2115 & ~n2636 ;
  assign n2649 = ~n2647 & n2648 ;
  assign n2650 = ~n2641 & n2649 ;
  assign n2651 = ~n2635 & n2650 ;
  assign n2652 = \PhyAddrPointer_reg[22]/NET0131  & ~n921 ;
  assign n2653 = ~n2130 & ~n2652 ;
  assign n2654 = n748 & ~n2653 ;
  assign n2655 = \PhyAddrPointer_reg[22]/NET0131  & ~n1997 ;
  assign n2656 = ~n2137 & ~n2655 ;
  assign n2657 = ~n2654 & n2656 ;
  assign n2658 = n948 & ~n2657 ;
  assign n2664 = ~\PhyAddrPointer_reg[22]/NET0131  & ~n2393 ;
  assign n2665 = ~n2394 & ~n2664 ;
  assign n2666 = n970 & n2665 ;
  assign n2659 = n2023 & ~n2366 ;
  assign n2661 = \PhyAddrPointer_reg[22]/NET0131  & n2659 ;
  assign n2660 = ~\PhyAddrPointer_reg[22]/NET0131  & ~n2659 ;
  assign n2662 = n952 & ~n2660 ;
  assign n2663 = ~n2661 & n2662 ;
  assign n2667 = \PhyAddrPointer_reg[22]/NET0131  & ~n2003 ;
  assign n2668 = ~n2152 & ~n2667 ;
  assign n2669 = ~n2663 & n2668 ;
  assign n2670 = ~n2666 & n2669 ;
  assign n2671 = ~n2658 & n2670 ;
  assign n2672 = \PhyAddrPointer_reg[24]/NET0131  & ~n921 ;
  assign n2673 = ~n2178 & ~n2672 ;
  assign n2674 = n748 & ~n2673 ;
  assign n2675 = \PhyAddrPointer_reg[24]/NET0131  & ~n1997 ;
  assign n2676 = ~n2184 & ~n2675 ;
  assign n2677 = ~n2674 & n2676 ;
  assign n2678 = n948 & ~n2677 ;
  assign n2682 = ~\PhyAddrPointer_reg[24]/NET0131  & ~n2396 ;
  assign n2683 = ~n2419 & ~n2682 ;
  assign n2684 = n2039 & n2683 ;
  assign n2681 = \PhyAddrPointer_reg[24]/NET0131  & ~n2400 ;
  assign n2679 = ~\PhyAddrPointer_reg[24]/NET0131  & n971 ;
  assign n2680 = n2025 & n2679 ;
  assign n2685 = ~n2195 & ~n2680 ;
  assign n2686 = ~n2681 & n2685 ;
  assign n2687 = ~n2684 & n2686 ;
  assign n2688 = ~n2678 & n2687 ;
  assign n2689 = \PhyAddrPointer_reg[26]/NET0131  & ~n921 ;
  assign n2690 = ~n1353 & ~n2309 ;
  assign n2691 = n1051 & ~n1953 ;
  assign n2692 = ~n2690 & n2691 ;
  assign n2694 = ~n1543 & n1773 ;
  assign n2693 = n1543 & ~n1773 ;
  assign n2695 = ~n1051 & ~n2693 ;
  assign n2696 = ~n2694 & n2695 ;
  assign n2697 = ~n2692 & ~n2696 ;
  assign n2698 = n921 & ~n2697 ;
  assign n2699 = ~n2689 & ~n2698 ;
  assign n2700 = n748 & ~n2699 ;
  assign n2701 = \PhyAddrPointer_reg[26]/NET0131  & ~n1997 ;
  assign n2702 = n1697 & n1813 ;
  assign n2703 = ~n1688 & ~n2702 ;
  assign n2704 = n1698 & n1813 ;
  assign n2705 = n930 & ~n2704 ;
  assign n2706 = ~n2703 & n2705 ;
  assign n2707 = ~n2701 & ~n2706 ;
  assign n2708 = ~n2700 & n2707 ;
  assign n2709 = n948 & ~n2708 ;
  assign n2710 = n2026 & ~n2366 ;
  assign n2711 = \PhyAddrPointer_reg[25]/NET0131  & n2710 ;
  assign n2718 = n952 & ~n2711 ;
  assign n2719 = n2003 & ~n2718 ;
  assign n2720 = \PhyAddrPointer_reg[26]/NET0131  & ~n2719 ;
  assign n2714 = \PhyAddrPointer_reg[25]/NET0131  & n2419 ;
  assign n2715 = ~\PhyAddrPointer_reg[26]/NET0131  & ~n2714 ;
  assign n2716 = ~n2420 & ~n2715 ;
  assign n2717 = n970 & n2716 ;
  assign n2712 = ~\PhyAddrPointer_reg[26]/NET0131  & n952 ;
  assign n2713 = n2711 & n2712 ;
  assign n2721 = \rEIP_reg[26]/NET0131  & n1731 ;
  assign n2722 = ~n2713 & ~n2721 ;
  assign n2723 = ~n2717 & n2722 ;
  assign n2724 = ~n2720 & n2723 ;
  assign n2725 = ~n2709 & n2724 ;
  assign n2729 = \InstAddrPointer_reg[9]/NET0131  & ~n921 ;
  assign n2734 = ~n1418 & ~n1420 ;
  assign n2735 = n1418 & n1420 ;
  assign n2736 = ~n2734 & ~n2735 ;
  assign n2737 = n1051 & ~n2736 ;
  assign n2730 = ~n1487 & ~n2164 ;
  assign n2731 = n1487 & n2164 ;
  assign n2732 = ~n2730 & ~n2731 ;
  assign n2733 = ~n1051 & ~n2732 ;
  assign n2738 = n921 & ~n2733 ;
  assign n2739 = ~n2737 & n2738 ;
  assign n2740 = ~n2729 & ~n2739 ;
  assign n2741 = n748 & ~n2740 ;
  assign n2744 = ~n1644 & ~n1657 ;
  assign n2743 = n1644 & n1657 ;
  assign n2745 = n930 & ~n2743 ;
  assign n2746 = ~n2744 & n2745 ;
  assign n2747 = ~n839 & n1420 ;
  assign n2742 = \InstAddrPointer_reg[9]/NET0131  & ~n2073 ;
  assign n2728 = ~n780 & n1487 ;
  assign n2748 = n809 & n1657 ;
  assign n2749 = ~n2728 & ~n2748 ;
  assign n2750 = ~n2742 & n2749 ;
  assign n2751 = ~n2747 & n2750 ;
  assign n2752 = ~n2746 & n2751 ;
  assign n2753 = ~n2741 & n2752 ;
  assign n2754 = n948 & ~n2753 ;
  assign n2726 = \rEIP_reg[9]/NET0131  & n1731 ;
  assign n2727 = \InstAddrPointer_reg[9]/NET0131  & ~n1736 ;
  assign n2755 = ~n2726 & ~n2727 ;
  assign n2756 = ~n2754 & n2755 ;
  assign n2765 = \PhyAddrPointer_reg[16]/NET0131  & ~n921 ;
  assign n2771 = n1380 & n1741 ;
  assign n2770 = ~n1380 & ~n1741 ;
  assign n2772 = n1051 & ~n2770 ;
  assign n2773 = ~n2771 & n2772 ;
  assign n2767 = n1516 & ~n1838 ;
  assign n2766 = ~n1516 & n1838 ;
  assign n2768 = ~n1051 & ~n2766 ;
  assign n2769 = ~n2767 & n2768 ;
  assign n2774 = n921 & ~n2769 ;
  assign n2775 = ~n2773 & n2774 ;
  assign n2776 = ~n2765 & ~n2775 ;
  assign n2777 = n748 & ~n2776 ;
  assign n2762 = n1870 & n1872 ;
  assign n2761 = ~n1870 & ~n1872 ;
  assign n2763 = n930 & ~n2761 ;
  assign n2764 = ~n2762 & n2763 ;
  assign n2778 = \PhyAddrPointer_reg[16]/NET0131  & ~n1997 ;
  assign n2779 = ~n2764 & ~n2778 ;
  assign n2780 = ~n2777 & n2779 ;
  assign n2781 = n948 & ~n2780 ;
  assign n2785 = ~\PhyAddrPointer_reg[16]/NET0131  & ~n2377 ;
  assign n2757 = n2015 & n2019 ;
  assign n2786 = \PhyAddrPointer_reg[1]/NET0131  & n2757 ;
  assign n2787 = ~n2785 & ~n2786 ;
  assign n2788 = n2039 & n2787 ;
  assign n2758 = n971 & ~n2757 ;
  assign n2782 = n2003 & ~n2758 ;
  assign n2783 = \PhyAddrPointer_reg[16]/NET0131  & ~n2782 ;
  assign n2759 = \PhyAddrPointer_reg[15]/NET0131  & n2365 ;
  assign n2760 = n2758 & n2759 ;
  assign n2784 = \rEIP_reg[16]/NET0131  & n1731 ;
  assign n2789 = ~n2760 & ~n2784 ;
  assign n2790 = ~n2783 & n2789 ;
  assign n2791 = ~n2788 & n2790 ;
  assign n2792 = ~n2781 & n2791 ;
  assign n2807 = \PhyAddrPointer_reg[17]/NET0131  & ~n921 ;
  assign n2815 = ~n1383 & n2302 ;
  assign n2814 = n1383 & ~n2302 ;
  assign n2816 = n1051 & ~n2814 ;
  assign n2817 = ~n2815 & n2816 ;
  assign n2808 = ~n1516 & n1836 ;
  assign n2809 = n2164 & n2808 ;
  assign n2811 = ~n1522 & n2809 ;
  assign n2810 = n1522 & ~n2809 ;
  assign n2812 = ~n1051 & ~n2810 ;
  assign n2813 = ~n2811 & n2812 ;
  assign n2818 = n921 & ~n2813 ;
  assign n2819 = ~n2817 & n2818 ;
  assign n2820 = ~n2807 & ~n2819 ;
  assign n2821 = n748 & ~n2820 ;
  assign n2804 = ~n1600 & ~n1666 ;
  assign n2805 = n930 & ~n2067 ;
  assign n2806 = ~n2804 & n2805 ;
  assign n2822 = \PhyAddrPointer_reg[17]/NET0131  & ~n1997 ;
  assign n2823 = ~n2806 & ~n2822 ;
  assign n2824 = ~n2821 & n2823 ;
  assign n2825 = n948 & ~n2824 ;
  assign n2800 = ~\PhyAddrPointer_reg[17]/NET0131  & ~n2786 ;
  assign n2801 = \PhyAddrPointer_reg[1]/NET0131  & n2613 ;
  assign n2802 = ~n2800 & ~n2801 ;
  assign n2803 = n2039 & n2802 ;
  assign n2793 = ~n955 & ~n957 ;
  assign n2794 = ~n1733 & n2793 ;
  assign n2795 = ~n2758 & n2794 ;
  assign n2796 = \PhyAddrPointer_reg[17]/NET0131  & ~n2795 ;
  assign n2797 = ~\PhyAddrPointer_reg[17]/NET0131  & n971 ;
  assign n2798 = n2757 & n2797 ;
  assign n2799 = \rEIP_reg[17]/NET0131  & n1731 ;
  assign n2826 = ~n2798 & ~n2799 ;
  assign n2827 = ~n2796 & n2826 ;
  assign n2828 = ~n2803 & n2827 ;
  assign n2829 = ~n2825 & n2828 ;
  assign n2830 = \PhyAddrPointer_reg[18]/NET0131  & ~n921 ;
  assign n2835 = ~n1387 & ~n2052 ;
  assign n2836 = ~n2053 & ~n2835 ;
  assign n2837 = n1051 & ~n2836 ;
  assign n2831 = n1520 & ~n2811 ;
  assign n2832 = n1523 & n2809 ;
  assign n2833 = ~n1051 & ~n2832 ;
  assign n2834 = ~n2831 & n2833 ;
  assign n2838 = n921 & ~n2834 ;
  assign n2839 = ~n2837 & n2838 ;
  assign n2840 = ~n2830 & ~n2839 ;
  assign n2841 = n748 & ~n2840 ;
  assign n2842 = \PhyAddrPointer_reg[18]/NET0131  & ~n1997 ;
  assign n2844 = n1807 & n1810 ;
  assign n2843 = ~n1807 & ~n1810 ;
  assign n2845 = n930 & ~n2843 ;
  assign n2846 = ~n2844 & n2845 ;
  assign n2847 = ~n2842 & ~n2846 ;
  assign n2848 = ~n2841 & n2847 ;
  assign n2849 = n948 & ~n2848 ;
  assign n2851 = ~\PhyAddrPointer_reg[18]/NET0131  & ~n2801 ;
  assign n2852 = ~n2620 & ~n2851 ;
  assign n2853 = n2039 & n2852 ;
  assign n2854 = ~\PhyAddrPointer_reg[18]/NET0131  & ~n2613 ;
  assign n2855 = n2615 & ~n2854 ;
  assign n2850 = \rEIP_reg[18]/NET0131  & n1731 ;
  assign n2856 = \PhyAddrPointer_reg[18]/NET0131  & ~n2003 ;
  assign n2857 = ~n2850 & ~n2856 ;
  assign n2858 = ~n2855 & n2857 ;
  assign n2859 = ~n2853 & n2858 ;
  assign n2860 = ~n2849 & n2859 ;
  assign n2861 = \PhyAddrPointer_reg[25]/NET0131  & ~n921 ;
  assign n2862 = ~n2317 & ~n2861 ;
  assign n2863 = n748 & ~n2862 ;
  assign n2864 = \PhyAddrPointer_reg[25]/NET0131  & ~n1997 ;
  assign n2865 = ~n2326 & ~n2864 ;
  assign n2866 = ~n2863 & n2865 ;
  assign n2867 = n948 & ~n2866 ;
  assign n2871 = ~\PhyAddrPointer_reg[25]/NET0131  & ~n2710 ;
  assign n2872 = n2718 & ~n2871 ;
  assign n2868 = ~\PhyAddrPointer_reg[25]/NET0131  & ~n2419 ;
  assign n2869 = ~n2714 & ~n2868 ;
  assign n2870 = n970 & n2869 ;
  assign n2873 = \PhyAddrPointer_reg[25]/NET0131  & ~n2003 ;
  assign n2874 = ~n2341 & ~n2873 ;
  assign n2875 = ~n2870 & n2874 ;
  assign n2876 = ~n2872 & n2875 ;
  assign n2877 = ~n2867 & n2876 ;
  assign n2883 = \PhyAddrPointer_reg[8]/NET0131  & ~n921 ;
  assign n2884 = ~n2503 & ~n2883 ;
  assign n2885 = n748 & ~n2884 ;
  assign n2886 = \PhyAddrPointer_reg[8]/NET0131  & ~n1997 ;
  assign n2887 = ~n2512 & ~n2886 ;
  assign n2888 = ~n2885 & n2887 ;
  assign n2889 = n948 & ~n2888 ;
  assign n2878 = \PhyAddrPointer_reg[1]/NET0131  & n2009 ;
  assign n2879 = ~\PhyAddrPointer_reg[8]/NET0131  & ~n2878 ;
  assign n2880 = \PhyAddrPointer_reg[1]/NET0131  & n2010 ;
  assign n2881 = ~n2879 & ~n2880 ;
  assign n2890 = ~\DataWidth_reg[1]/NET0131  & ~n2881 ;
  assign n2891 = ~\PhyAddrPointer_reg[8]/NET0131  & ~n2009 ;
  assign n2892 = ~n2010 & ~n2891 ;
  assign n2893 = \DataWidth_reg[1]/NET0131  & ~n2892 ;
  assign n2894 = n952 & ~n2893 ;
  assign n2895 = ~n2890 & n2894 ;
  assign n2882 = n970 & n2881 ;
  assign n2896 = \PhyAddrPointer_reg[8]/NET0131  & ~n2003 ;
  assign n2897 = ~n2492 & ~n2896 ;
  assign n2898 = ~n2882 & n2897 ;
  assign n2899 = ~n2895 & n2898 ;
  assign n2900 = ~n2889 & n2899 ;
  assign n2908 = ~n875 & n924 ;
  assign n2909 = ~n836 & ~n997 ;
  assign n2910 = n2908 & ~n2909 ;
  assign n2911 = \InstAddrPointer_reg[4]/NET0131  & ~n2910 ;
  assign n2907 = ~n780 & n1461 ;
  assign n2903 = ~n808 & n1591 ;
  assign n2904 = n1609 & ~n2903 ;
  assign n2905 = ~n756 & n2904 ;
  assign n2906 = ~n867 & n1123 ;
  assign n2926 = ~n2905 & ~n2906 ;
  assign n2927 = ~n2907 & n2926 ;
  assign n2928 = ~n2911 & n2927 ;
  assign n2912 = \InstAddrPointer_reg[4]/NET0131  & ~n921 ;
  assign n2913 = ~n1157 & ~n1307 ;
  assign n2914 = ~n1303 & ~n2913 ;
  assign n2915 = n1303 & n2913 ;
  assign n2916 = ~n2914 & ~n2915 ;
  assign n2917 = n921 & ~n2916 ;
  assign n2918 = ~n2912 & ~n2917 ;
  assign n2919 = n748 & ~n2918 ;
  assign n2920 = ~n1610 & ~n1624 ;
  assign n2921 = ~n1613 & ~n1786 ;
  assign n2923 = n2920 & n2921 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2924 = n930 & ~n2922 ;
  assign n2925 = ~n2923 & n2924 ;
  assign n2929 = ~n2919 & ~n2925 ;
  assign n2930 = n2928 & n2929 ;
  assign n2931 = n948 & ~n2930 ;
  assign n2901 = \rEIP_reg[4]/NET0131  & n1731 ;
  assign n2902 = \InstAddrPointer_reg[4]/NET0131  & ~n1736 ;
  assign n2932 = ~n2901 & ~n2902 ;
  assign n2933 = ~n2931 & n2932 ;
  assign n2941 = \InstAddrPointer_reg[6]/NET0131  & ~n921 ;
  assign n2947 = ~n1087 & ~n1314 ;
  assign n2948 = n1310 & ~n2947 ;
  assign n2949 = ~n1310 & n2947 ;
  assign n2950 = ~n2948 & ~n2949 ;
  assign n2951 = n1051 & ~n2950 ;
  assign n2942 = ~n1443 & ~n1474 ;
  assign n2944 = n1757 & n2942 ;
  assign n2943 = ~n1757 & ~n2942 ;
  assign n2945 = ~n1051 & ~n2943 ;
  assign n2946 = ~n2944 & n2945 ;
  assign n2952 = n921 & ~n2946 ;
  assign n2953 = ~n2951 & n2952 ;
  assign n2954 = ~n2941 & ~n2953 ;
  assign n2955 = n748 & ~n2954 ;
  assign n2957 = ~n1607 & ~n1634 ;
  assign n2959 = ~n1791 & n2957 ;
  assign n2958 = n1791 & ~n2957 ;
  assign n2960 = n930 & ~n2958 ;
  assign n2961 = ~n2959 & n2960 ;
  assign n2938 = ~n1053 & n2506 ;
  assign n2939 = n839 & ~n2938 ;
  assign n2940 = n1055 & ~n2939 ;
  assign n2937 = \InstAddrPointer_reg[6]/NET0131  & ~n2508 ;
  assign n2936 = n809 & n1606 ;
  assign n2956 = ~n780 & n1442 ;
  assign n2962 = ~n2936 & ~n2956 ;
  assign n2963 = ~n2937 & n2962 ;
  assign n2964 = ~n2940 & n2963 ;
  assign n2965 = ~n2961 & n2964 ;
  assign n2966 = ~n2955 & n2965 ;
  assign n2967 = n948 & ~n2966 ;
  assign n2934 = \rEIP_reg[6]/NET0131  & n1731 ;
  assign n2935 = \InstAddrPointer_reg[6]/NET0131  & ~n1736 ;
  assign n2968 = ~n2934 & ~n2935 ;
  assign n2969 = ~n2967 & n2968 ;
  assign n2973 = \PhyAddrPointer_reg[10]/NET0131  & ~n921 ;
  assign n2977 = ~n2533 & ~n2535 ;
  assign n2978 = ~n2536 & ~n2977 ;
  assign n2979 = n1051 & ~n2978 ;
  assign n2974 = n1484 & ~n2525 ;
  assign n2975 = ~n1051 & ~n1494 ;
  assign n2976 = ~n2974 & n2975 ;
  assign n2980 = n921 & ~n2976 ;
  assign n2981 = ~n2979 & n2980 ;
  assign n2982 = ~n2973 & ~n2981 ;
  assign n2983 = n748 & ~n2982 ;
  assign n2970 = ~n1797 & ~n1799 ;
  assign n2971 = n930 & ~n2276 ;
  assign n2972 = ~n2970 & n2971 ;
  assign n2984 = \PhyAddrPointer_reg[10]/NET0131  & ~n1997 ;
  assign n2985 = ~n2972 & ~n2984 ;
  assign n2986 = ~n2983 & n2985 ;
  assign n2987 = n948 & ~n2986 ;
  assign n2988 = \PhyAddrPointer_reg[1]/NET0131  & n2011 ;
  assign n2989 = ~\PhyAddrPointer_reg[10]/NET0131  & ~n2988 ;
  assign n2990 = ~n2579 & ~n2989 ;
  assign n2992 = ~\DataWidth_reg[1]/NET0131  & ~n2990 ;
  assign n2993 = ~\PhyAddrPointer_reg[10]/NET0131  & ~n2011 ;
  assign n2994 = ~n2012 & ~n2993 ;
  assign n2995 = \DataWidth_reg[1]/NET0131  & ~n2994 ;
  assign n2996 = n952 & ~n2995 ;
  assign n2997 = ~n2992 & n2996 ;
  assign n2991 = n970 & n2990 ;
  assign n2998 = \rEIP_reg[10]/NET0131  & n1731 ;
  assign n2999 = \PhyAddrPointer_reg[10]/NET0131  & ~n2003 ;
  assign n3000 = ~n2998 & ~n2999 ;
  assign n3001 = ~n2991 & n3000 ;
  assign n3002 = ~n2997 & n3001 ;
  assign n3003 = ~n2987 & n3002 ;
  assign n3015 = \PhyAddrPointer_reg[7]/NET0131  & ~n921 ;
  assign n3020 = ~n1412 & n1414 ;
  assign n3022 = n1017 & n3020 ;
  assign n3021 = ~n1017 & ~n3020 ;
  assign n3023 = n1051 & ~n3021 ;
  assign n3024 = ~n3022 & n3023 ;
  assign n3017 = ~n1438 & n1479 ;
  assign n3016 = n1438 & ~n1479 ;
  assign n3018 = ~n1051 & ~n3016 ;
  assign n3019 = ~n3017 & n3018 ;
  assign n3025 = n921 & ~n3019 ;
  assign n3026 = ~n3024 & n3025 ;
  assign n3027 = ~n3015 & ~n3026 ;
  assign n3028 = n748 & ~n3027 ;
  assign n3009 = ~n1633 & ~n1640 ;
  assign n3010 = ~n1630 & n1637 ;
  assign n3012 = n3009 & ~n3010 ;
  assign n3011 = ~n3009 & n3010 ;
  assign n3013 = n930 & ~n3011 ;
  assign n3014 = ~n3012 & n3013 ;
  assign n3029 = \PhyAddrPointer_reg[7]/NET0131  & ~n1997 ;
  assign n3030 = ~n3014 & ~n3029 ;
  assign n3031 = ~n3028 & n3030 ;
  assign n3032 = n948 & ~n3031 ;
  assign n3004 = \PhyAddrPointer_reg[1]/NET0131  & n2007 ;
  assign n3005 = \PhyAddrPointer_reg[6]/NET0131  & n3004 ;
  assign n3006 = ~\PhyAddrPointer_reg[7]/NET0131  & ~n3005 ;
  assign n3007 = ~n2878 & ~n3006 ;
  assign n3033 = ~\DataWidth_reg[1]/NET0131  & ~n3007 ;
  assign n3034 = ~\PhyAddrPointer_reg[7]/NET0131  & ~n2008 ;
  assign n3035 = ~n2009 & ~n3034 ;
  assign n3036 = \DataWidth_reg[1]/NET0131  & ~n3035 ;
  assign n3037 = n952 & ~n3036 ;
  assign n3038 = ~n3033 & n3037 ;
  assign n3008 = n970 & n3007 ;
  assign n3039 = \rEIP_reg[7]/NET0131  & n1731 ;
  assign n3040 = \PhyAddrPointer_reg[7]/NET0131  & ~n2003 ;
  assign n3041 = ~n3039 & ~n3040 ;
  assign n3042 = ~n3008 & n3041 ;
  assign n3043 = ~n3038 & n3042 ;
  assign n3044 = ~n3032 & n3043 ;
  assign n3062 = \InstAddrPointer_reg[3]/NET0131  & ~n921 ;
  assign n3068 = ~n1192 & ~n1299 ;
  assign n3069 = ~n1226 & ~n1405 ;
  assign n3070 = ~n3068 & ~n3069 ;
  assign n3071 = n3068 & n3069 ;
  assign n3072 = ~n3070 & ~n3071 ;
  assign n3073 = n1051 & ~n3072 ;
  assign n3065 = ~n1465 & n1752 ;
  assign n3063 = ~n1465 & ~n1470 ;
  assign n3064 = ~n1459 & ~n3063 ;
  assign n3066 = ~n1051 & ~n3064 ;
  assign n3067 = ~n3065 & n3066 ;
  assign n3074 = n921 & ~n3067 ;
  assign n3075 = ~n3073 & n3074 ;
  assign n3076 = ~n3062 & ~n3075 ;
  assign n3077 = n748 & ~n3076 ;
  assign n3061 = ~n780 & n1464 ;
  assign n3049 = ~n1613 & ~n1625 ;
  assign n3051 = ~n1622 & ~n3049 ;
  assign n3050 = n1622 & n3049 ;
  assign n3052 = n930 & ~n3050 ;
  assign n3053 = ~n3051 & n3052 ;
  assign n3047 = n809 & n1612 ;
  assign n3048 = n698 & n1191 ;
  assign n3078 = ~n3047 & ~n3048 ;
  assign n3079 = ~n3053 & n3078 ;
  assign n3080 = ~n3061 & n3079 ;
  assign n3055 = \InstAddrPointer_reg[3]/NET0131  & n835 ;
  assign n3056 = ~n2506 & ~n3055 ;
  assign n3054 = ~\InstAddrPointer_reg[3]/NET0131  & READY_n_pad ;
  assign n3057 = ~READY_n_pad & ~n1191 ;
  assign n3058 = ~n3054 & ~n3057 ;
  assign n3059 = ~n3056 & n3058 ;
  assign n3060 = \InstAddrPointer_reg[3]/NET0131  & ~n1892 ;
  assign n3081 = ~n3059 & ~n3060 ;
  assign n3082 = n3080 & n3081 ;
  assign n3083 = ~n3077 & n3082 ;
  assign n3084 = n948 & ~n3083 ;
  assign n3045 = \rEIP_reg[3]/NET0131  & n1731 ;
  assign n3046 = \InstAddrPointer_reg[3]/NET0131  & ~n1736 ;
  assign n3085 = ~n3045 & ~n3046 ;
  assign n3086 = ~n3084 & n3085 ;
  assign n3089 = \InstAddrPointer_reg[5]/NET0131  & ~n921 ;
  assign n3090 = ~n1121 & ~n1306 ;
  assign n3091 = ~n1410 & ~n3090 ;
  assign n3092 = n1410 & n3090 ;
  assign n3093 = ~n3091 & ~n3092 ;
  assign n3094 = n921 & ~n3093 ;
  assign n3095 = ~n3089 & ~n3094 ;
  assign n3096 = n748 & ~n3095 ;
  assign n3101 = ~n1604 & ~n1635 ;
  assign n3103 = ~n1628 & n3101 ;
  assign n3102 = n1628 & ~n3101 ;
  assign n3104 = n930 & ~n3102 ;
  assign n3105 = ~n3103 & n3104 ;
  assign n3098 = \InstAddrPointer_reg[5]/NET0131  & ~n2908 ;
  assign n3100 = ~n867 & n1089 ;
  assign n3097 = ~n780 & n1445 ;
  assign n3099 = n809 & n1603 ;
  assign n3106 = ~n3097 & ~n3099 ;
  assign n3107 = ~n3100 & n3106 ;
  assign n3108 = ~n3098 & n3107 ;
  assign n3109 = ~n3105 & n3108 ;
  assign n3110 = ~n3096 & n3109 ;
  assign n3111 = n948 & ~n3110 ;
  assign n3087 = \rEIP_reg[5]/NET0131  & n1731 ;
  assign n3088 = \InstAddrPointer_reg[5]/NET0131  & ~n1736 ;
  assign n3112 = ~n3087 & ~n3088 ;
  assign n3113 = ~n3111 & n3112 ;
  assign n3114 = ~n980 & ~n984 ;
  assign n3115 = ~n968 & ~n982 ;
  assign n3116 = n3114 & n3115 ;
  assign n3117 = \EAX_reg[31]/NET0131  & ~n3116 ;
  assign n3119 = \EAX_reg[0]/NET0131  & \EAX_reg[1]/NET0131  ;
  assign n3120 = \EAX_reg[2]/NET0131  & n3119 ;
  assign n3121 = \EAX_reg[3]/NET0131  & n3120 ;
  assign n3122 = \EAX_reg[4]/NET0131  & n3121 ;
  assign n3123 = \EAX_reg[5]/NET0131  & n3122 ;
  assign n3124 = \EAX_reg[6]/NET0131  & n3123 ;
  assign n3125 = \EAX_reg[7]/NET0131  & n3124 ;
  assign n3126 = \EAX_reg[8]/NET0131  & n3125 ;
  assign n3127 = \EAX_reg[9]/NET0131  & n3126 ;
  assign n3128 = \EAX_reg[10]/NET0131  & n3127 ;
  assign n3129 = \EAX_reg[11]/NET0131  & n3128 ;
  assign n3130 = \EAX_reg[12]/NET0131  & n3129 ;
  assign n3131 = \EAX_reg[13]/NET0131  & n3130 ;
  assign n3132 = \EAX_reg[14]/NET0131  & n3131 ;
  assign n3133 = \EAX_reg[15]/NET0131  & n3132 ;
  assign n3134 = \EAX_reg[16]/NET0131  & n3133 ;
  assign n3135 = \EAX_reg[17]/NET0131  & n3134 ;
  assign n3136 = \EAX_reg[18]/NET0131  & n3135 ;
  assign n3137 = \EAX_reg[19]/NET0131  & n3136 ;
  assign n3138 = \EAX_reg[20]/NET0131  & \EAX_reg[21]/NET0131  ;
  assign n3139 = \EAX_reg[22]/NET0131  & n3138 ;
  assign n3140 = n3137 & n3139 ;
  assign n3141 = \EAX_reg[23]/NET0131  & \EAX_reg[24]/NET0131  ;
  assign n3142 = \EAX_reg[25]/NET0131  & n3141 ;
  assign n3143 = \EAX_reg[26]/NET0131  & \EAX_reg[27]/NET0131  ;
  assign n3144 = n3142 & n3143 ;
  assign n3145 = n3140 & n3144 ;
  assign n3146 = \EAX_reg[28]/NET0131  & \EAX_reg[29]/NET0131  ;
  assign n3147 = n3145 & n3146 ;
  assign n3148 = \EAX_reg[30]/NET0131  & n3147 ;
  assign n3150 = \EAX_reg[31]/NET0131  & n3148 ;
  assign n3118 = n665 & n767 ;
  assign n3149 = ~\EAX_reg[31]/NET0131  & ~n3148 ;
  assign n3151 = n3118 & ~n3149 ;
  assign n3152 = ~n3150 & n3151 ;
  assign n3153 = n755 & n808 ;
  assign n3443 = n836 & ~n3118 ;
  assign n3444 = ~n755 & ~n3443 ;
  assign n3445 = ~n3153 & ~n3444 ;
  assign n3446 = ~n844 & ~n3445 ;
  assign n3447 = ~n872 & n3446 ;
  assign n3448 = \EAX_reg[31]/NET0131  & ~n3447 ;
  assign n3158 = \InstQueue_reg[14][7]/NET0131  & n474 ;
  assign n3159 = \InstQueue_reg[0][7]/NET0131  & n471 ;
  assign n3172 = ~n3158 & ~n3159 ;
  assign n3160 = \InstQueue_reg[2][7]/NET0131  & n476 ;
  assign n3161 = \InstQueue_reg[9][7]/NET0131  & n457 ;
  assign n3173 = ~n3160 & ~n3161 ;
  assign n3180 = n3172 & n3173 ;
  assign n3154 = \InstQueue_reg[5][7]/NET0131  & n478 ;
  assign n3155 = \InstQueue_reg[11][7]/NET0131  & n486 ;
  assign n3170 = ~n3154 & ~n3155 ;
  assign n3156 = \InstQueue_reg[8][7]/NET0131  & n484 ;
  assign n3157 = \InstQueue_reg[4][7]/NET0131  & n466 ;
  assign n3171 = ~n3156 & ~n3157 ;
  assign n3181 = n3170 & n3171 ;
  assign n3182 = n3180 & n3181 ;
  assign n3166 = \InstQueue_reg[15][7]/NET0131  & n488 ;
  assign n3167 = \InstQueue_reg[10][7]/NET0131  & n482 ;
  assign n3176 = ~n3166 & ~n3167 ;
  assign n3168 = \InstQueue_reg[13][7]/NET0131  & n490 ;
  assign n3169 = \InstQueue_reg[6][7]/NET0131  & n480 ;
  assign n3177 = ~n3168 & ~n3169 ;
  assign n3178 = n3176 & n3177 ;
  assign n3162 = \InstQueue_reg[3][7]/NET0131  & n461 ;
  assign n3163 = \InstQueue_reg[1][7]/NET0131  & n454 ;
  assign n3174 = ~n3162 & ~n3163 ;
  assign n3164 = \InstQueue_reg[7][7]/NET0131  & n463 ;
  assign n3165 = \InstQueue_reg[12][7]/NET0131  & n469 ;
  assign n3175 = ~n3164 & ~n3165 ;
  assign n3179 = n3174 & n3175 ;
  assign n3183 = n3178 & n3179 ;
  assign n3184 = n3182 & n3183 ;
  assign n3189 = \InstQueue_reg[7][0]/NET0131  & n480 ;
  assign n3190 = \InstQueue_reg[15][0]/NET0131  & n474 ;
  assign n3203 = ~n3189 & ~n3190 ;
  assign n3191 = \InstQueue_reg[3][0]/NET0131  & n476 ;
  assign n3192 = \InstQueue_reg[4][0]/NET0131  & n461 ;
  assign n3204 = ~n3191 & ~n3192 ;
  assign n3211 = n3203 & n3204 ;
  assign n3185 = \InstQueue_reg[10][0]/NET0131  & n457 ;
  assign n3186 = \InstQueue_reg[0][0]/NET0131  & n488 ;
  assign n3201 = ~n3185 & ~n3186 ;
  assign n3187 = \InstQueue_reg[8][0]/NET0131  & n463 ;
  assign n3188 = \InstQueue_reg[9][0]/NET0131  & n484 ;
  assign n3202 = ~n3187 & ~n3188 ;
  assign n3212 = n3201 & n3202 ;
  assign n3213 = n3211 & n3212 ;
  assign n3197 = \InstQueue_reg[5][0]/NET0131  & n466 ;
  assign n3198 = \InstQueue_reg[11][0]/NET0131  & n482 ;
  assign n3207 = ~n3197 & ~n3198 ;
  assign n3199 = \InstQueue_reg[6][0]/NET0131  & n478 ;
  assign n3200 = \InstQueue_reg[13][0]/NET0131  & n469 ;
  assign n3208 = ~n3199 & ~n3200 ;
  assign n3209 = n3207 & n3208 ;
  assign n3193 = \InstQueue_reg[12][0]/NET0131  & n486 ;
  assign n3194 = \InstQueue_reg[2][0]/NET0131  & n454 ;
  assign n3205 = ~n3193 & ~n3194 ;
  assign n3195 = \InstQueue_reg[1][0]/NET0131  & n471 ;
  assign n3196 = \InstQueue_reg[14][0]/NET0131  & n490 ;
  assign n3206 = ~n3195 & ~n3196 ;
  assign n3210 = n3205 & n3206 ;
  assign n3214 = n3209 & n3210 ;
  assign n3215 = n3213 & n3214 ;
  assign n3216 = ~n3184 & ~n3215 ;
  assign n3221 = \InstQueue_reg[11][1]/NET0131  & n482 ;
  assign n3222 = \InstQueue_reg[9][1]/NET0131  & n484 ;
  assign n3235 = ~n3221 & ~n3222 ;
  assign n3223 = \InstQueue_reg[15][1]/NET0131  & n474 ;
  assign n3224 = \InstQueue_reg[4][1]/NET0131  & n461 ;
  assign n3236 = ~n3223 & ~n3224 ;
  assign n3243 = n3235 & n3236 ;
  assign n3217 = \InstQueue_reg[8][1]/NET0131  & n463 ;
  assign n3218 = \InstQueue_reg[1][1]/NET0131  & n471 ;
  assign n3233 = ~n3217 & ~n3218 ;
  assign n3219 = \InstQueue_reg[0][1]/NET0131  & n488 ;
  assign n3220 = \InstQueue_reg[6][1]/NET0131  & n478 ;
  assign n3234 = ~n3219 & ~n3220 ;
  assign n3244 = n3233 & n3234 ;
  assign n3245 = n3243 & n3244 ;
  assign n3229 = \InstQueue_reg[7][1]/NET0131  & n480 ;
  assign n3230 = \InstQueue_reg[3][1]/NET0131  & n476 ;
  assign n3239 = ~n3229 & ~n3230 ;
  assign n3231 = \InstQueue_reg[13][1]/NET0131  & n469 ;
  assign n3232 = \InstQueue_reg[14][1]/NET0131  & n490 ;
  assign n3240 = ~n3231 & ~n3232 ;
  assign n3241 = n3239 & n3240 ;
  assign n3225 = \InstQueue_reg[12][1]/NET0131  & n486 ;
  assign n3226 = \InstQueue_reg[2][1]/NET0131  & n454 ;
  assign n3237 = ~n3225 & ~n3226 ;
  assign n3227 = \InstQueue_reg[5][1]/NET0131  & n466 ;
  assign n3228 = \InstQueue_reg[10][1]/NET0131  & n457 ;
  assign n3238 = ~n3227 & ~n3228 ;
  assign n3242 = n3237 & n3238 ;
  assign n3246 = n3241 & n3242 ;
  assign n3247 = n3245 & n3246 ;
  assign n3248 = n3216 & ~n3247 ;
  assign n3253 = \InstQueue_reg[3][2]/NET0131  & n476 ;
  assign n3254 = \InstQueue_reg[5][2]/NET0131  & n466 ;
  assign n3267 = ~n3253 & ~n3254 ;
  assign n3255 = \InstQueue_reg[8][2]/NET0131  & n463 ;
  assign n3256 = \InstQueue_reg[14][2]/NET0131  & n490 ;
  assign n3268 = ~n3255 & ~n3256 ;
  assign n3275 = n3267 & n3268 ;
  assign n3249 = \InstQueue_reg[15][2]/NET0131  & n474 ;
  assign n3250 = \InstQueue_reg[1][2]/NET0131  & n471 ;
  assign n3265 = ~n3249 & ~n3250 ;
  assign n3251 = \InstQueue_reg[4][2]/NET0131  & n461 ;
  assign n3252 = \InstQueue_reg[13][2]/NET0131  & n469 ;
  assign n3266 = ~n3251 & ~n3252 ;
  assign n3276 = n3265 & n3266 ;
  assign n3277 = n3275 & n3276 ;
  assign n3261 = \InstQueue_reg[9][2]/NET0131  & n484 ;
  assign n3262 = \InstQueue_reg[11][2]/NET0131  & n482 ;
  assign n3271 = ~n3261 & ~n3262 ;
  assign n3263 = \InstQueue_reg[7][2]/NET0131  & n480 ;
  assign n3264 = \InstQueue_reg[10][2]/NET0131  & n457 ;
  assign n3272 = ~n3263 & ~n3264 ;
  assign n3273 = n3271 & n3272 ;
  assign n3257 = \InstQueue_reg[6][2]/NET0131  & n478 ;
  assign n3258 = \InstQueue_reg[2][2]/NET0131  & n454 ;
  assign n3269 = ~n3257 & ~n3258 ;
  assign n3259 = \InstQueue_reg[0][2]/NET0131  & n488 ;
  assign n3260 = \InstQueue_reg[12][2]/NET0131  & n486 ;
  assign n3270 = ~n3259 & ~n3260 ;
  assign n3274 = n3269 & n3270 ;
  assign n3278 = n3273 & n3274 ;
  assign n3279 = n3277 & n3278 ;
  assign n3280 = n3248 & ~n3279 ;
  assign n3285 = \InstQueue_reg[3][3]/NET0131  & n476 ;
  assign n3286 = \InstQueue_reg[5][3]/NET0131  & n466 ;
  assign n3299 = ~n3285 & ~n3286 ;
  assign n3287 = \InstQueue_reg[8][3]/NET0131  & n463 ;
  assign n3288 = \InstQueue_reg[14][3]/NET0131  & n490 ;
  assign n3300 = ~n3287 & ~n3288 ;
  assign n3307 = n3299 & n3300 ;
  assign n3281 = \InstQueue_reg[15][3]/NET0131  & n474 ;
  assign n3282 = \InstQueue_reg[1][3]/NET0131  & n471 ;
  assign n3297 = ~n3281 & ~n3282 ;
  assign n3283 = \InstQueue_reg[4][3]/NET0131  & n461 ;
  assign n3284 = \InstQueue_reg[13][3]/NET0131  & n469 ;
  assign n3298 = ~n3283 & ~n3284 ;
  assign n3308 = n3297 & n3298 ;
  assign n3309 = n3307 & n3308 ;
  assign n3293 = \InstQueue_reg[9][3]/NET0131  & n484 ;
  assign n3294 = \InstQueue_reg[11][3]/NET0131  & n482 ;
  assign n3303 = ~n3293 & ~n3294 ;
  assign n3295 = \InstQueue_reg[7][3]/NET0131  & n480 ;
  assign n3296 = \InstQueue_reg[10][3]/NET0131  & n457 ;
  assign n3304 = ~n3295 & ~n3296 ;
  assign n3305 = n3303 & n3304 ;
  assign n3289 = \InstQueue_reg[6][3]/NET0131  & n478 ;
  assign n3290 = \InstQueue_reg[2][3]/NET0131  & n454 ;
  assign n3301 = ~n3289 & ~n3290 ;
  assign n3291 = \InstQueue_reg[0][3]/NET0131  & n488 ;
  assign n3292 = \InstQueue_reg[12][3]/NET0131  & n486 ;
  assign n3302 = ~n3291 & ~n3292 ;
  assign n3306 = n3301 & n3302 ;
  assign n3310 = n3305 & n3306 ;
  assign n3311 = n3309 & n3310 ;
  assign n3312 = n3280 & ~n3311 ;
  assign n3317 = \InstQueue_reg[11][4]/NET0131  & n482 ;
  assign n3318 = \InstQueue_reg[9][4]/NET0131  & n484 ;
  assign n3331 = ~n3317 & ~n3318 ;
  assign n3319 = \InstQueue_reg[15][4]/NET0131  & n474 ;
  assign n3320 = \InstQueue_reg[4][4]/NET0131  & n461 ;
  assign n3332 = ~n3319 & ~n3320 ;
  assign n3339 = n3331 & n3332 ;
  assign n3313 = \InstQueue_reg[8][4]/NET0131  & n463 ;
  assign n3314 = \InstQueue_reg[1][4]/NET0131  & n471 ;
  assign n3329 = ~n3313 & ~n3314 ;
  assign n3315 = \InstQueue_reg[0][4]/NET0131  & n488 ;
  assign n3316 = \InstQueue_reg[6][4]/NET0131  & n478 ;
  assign n3330 = ~n3315 & ~n3316 ;
  assign n3340 = n3329 & n3330 ;
  assign n3341 = n3339 & n3340 ;
  assign n3325 = \InstQueue_reg[7][4]/NET0131  & n480 ;
  assign n3326 = \InstQueue_reg[3][4]/NET0131  & n476 ;
  assign n3335 = ~n3325 & ~n3326 ;
  assign n3327 = \InstQueue_reg[13][4]/NET0131  & n469 ;
  assign n3328 = \InstQueue_reg[14][4]/NET0131  & n490 ;
  assign n3336 = ~n3327 & ~n3328 ;
  assign n3337 = n3335 & n3336 ;
  assign n3321 = \InstQueue_reg[12][4]/NET0131  & n486 ;
  assign n3322 = \InstQueue_reg[2][4]/NET0131  & n454 ;
  assign n3333 = ~n3321 & ~n3322 ;
  assign n3323 = \InstQueue_reg[5][4]/NET0131  & n466 ;
  assign n3324 = \InstQueue_reg[10][4]/NET0131  & n457 ;
  assign n3334 = ~n3323 & ~n3324 ;
  assign n3338 = n3333 & n3334 ;
  assign n3342 = n3337 & n3338 ;
  assign n3343 = n3341 & n3342 ;
  assign n3344 = n3312 & ~n3343 ;
  assign n3349 = \InstQueue_reg[3][5]/NET0131  & n476 ;
  assign n3350 = \InstQueue_reg[9][5]/NET0131  & n484 ;
  assign n3363 = ~n3349 & ~n3350 ;
  assign n3351 = \InstQueue_reg[14][5]/NET0131  & n490 ;
  assign n3352 = \InstQueue_reg[6][5]/NET0131  & n478 ;
  assign n3364 = ~n3351 & ~n3352 ;
  assign n3371 = n3363 & n3364 ;
  assign n3345 = \InstQueue_reg[10][5]/NET0131  & n457 ;
  assign n3346 = \InstQueue_reg[12][5]/NET0131  & n486 ;
  assign n3361 = ~n3345 & ~n3346 ;
  assign n3347 = \InstQueue_reg[4][5]/NET0131  & n461 ;
  assign n3348 = \InstQueue_reg[13][5]/NET0131  & n469 ;
  assign n3362 = ~n3347 & ~n3348 ;
  assign n3372 = n3361 & n3362 ;
  assign n3373 = n3371 & n3372 ;
  assign n3357 = \InstQueue_reg[5][5]/NET0131  & n466 ;
  assign n3358 = \InstQueue_reg[11][5]/NET0131  & n482 ;
  assign n3367 = ~n3357 & ~n3358 ;
  assign n3359 = \InstQueue_reg[1][5]/NET0131  & n471 ;
  assign n3360 = \InstQueue_reg[8][5]/NET0131  & n463 ;
  assign n3368 = ~n3359 & ~n3360 ;
  assign n3369 = n3367 & n3368 ;
  assign n3353 = \InstQueue_reg[0][5]/NET0131  & n488 ;
  assign n3354 = \InstQueue_reg[2][5]/NET0131  & n454 ;
  assign n3365 = ~n3353 & ~n3354 ;
  assign n3355 = \InstQueue_reg[7][5]/NET0131  & n480 ;
  assign n3356 = \InstQueue_reg[15][5]/NET0131  & n474 ;
  assign n3366 = ~n3355 & ~n3356 ;
  assign n3370 = n3365 & n3366 ;
  assign n3374 = n3369 & n3370 ;
  assign n3375 = n3373 & n3374 ;
  assign n3376 = n3344 & ~n3375 ;
  assign n3381 = \InstQueue_reg[3][6]/NET0131  & n476 ;
  assign n3382 = \InstQueue_reg[15][6]/NET0131  & n474 ;
  assign n3395 = ~n3381 & ~n3382 ;
  assign n3383 = \InstQueue_reg[10][6]/NET0131  & n457 ;
  assign n3384 = \InstQueue_reg[9][6]/NET0131  & n484 ;
  assign n3396 = ~n3383 & ~n3384 ;
  assign n3403 = n3395 & n3396 ;
  assign n3377 = \InstQueue_reg[14][6]/NET0131  & n490 ;
  assign n3378 = \InstQueue_reg[1][6]/NET0131  & n471 ;
  assign n3393 = ~n3377 & ~n3378 ;
  assign n3379 = \InstQueue_reg[8][6]/NET0131  & n463 ;
  assign n3380 = \InstQueue_reg[0][6]/NET0131  & n488 ;
  assign n3394 = ~n3379 & ~n3380 ;
  assign n3404 = n3393 & n3394 ;
  assign n3405 = n3403 & n3404 ;
  assign n3389 = \InstQueue_reg[5][6]/NET0131  & n466 ;
  assign n3390 = \InstQueue_reg[11][6]/NET0131  & n482 ;
  assign n3399 = ~n3389 & ~n3390 ;
  assign n3391 = \InstQueue_reg[6][6]/NET0131  & n478 ;
  assign n3392 = \InstQueue_reg[4][6]/NET0131  & n461 ;
  assign n3400 = ~n3391 & ~n3392 ;
  assign n3401 = n3399 & n3400 ;
  assign n3385 = \InstQueue_reg[12][6]/NET0131  & n486 ;
  assign n3386 = \InstQueue_reg[2][6]/NET0131  & n454 ;
  assign n3397 = ~n3385 & ~n3386 ;
  assign n3387 = \InstQueue_reg[13][6]/NET0131  & n469 ;
  assign n3388 = \InstQueue_reg[7][6]/NET0131  & n480 ;
  assign n3398 = ~n3387 & ~n3388 ;
  assign n3402 = n3397 & n3398 ;
  assign n3406 = n3401 & n3402 ;
  assign n3407 = n3405 & n3406 ;
  assign n3408 = n3376 & ~n3407 ;
  assign n3413 = \InstQueue_reg[3][7]/NET0131  & n476 ;
  assign n3414 = \InstQueue_reg[5][7]/NET0131  & n466 ;
  assign n3427 = ~n3413 & ~n3414 ;
  assign n3415 = \InstQueue_reg[8][7]/NET0131  & n463 ;
  assign n3416 = \InstQueue_reg[14][7]/NET0131  & n490 ;
  assign n3428 = ~n3415 & ~n3416 ;
  assign n3435 = n3427 & n3428 ;
  assign n3409 = \InstQueue_reg[15][7]/NET0131  & n474 ;
  assign n3410 = \InstQueue_reg[1][7]/NET0131  & n471 ;
  assign n3425 = ~n3409 & ~n3410 ;
  assign n3411 = \InstQueue_reg[4][7]/NET0131  & n461 ;
  assign n3412 = \InstQueue_reg[13][7]/NET0131  & n469 ;
  assign n3426 = ~n3411 & ~n3412 ;
  assign n3436 = n3425 & n3426 ;
  assign n3437 = n3435 & n3436 ;
  assign n3421 = \InstQueue_reg[9][7]/NET0131  & n484 ;
  assign n3422 = \InstQueue_reg[11][7]/NET0131  & n482 ;
  assign n3431 = ~n3421 & ~n3422 ;
  assign n3423 = \InstQueue_reg[7][7]/NET0131  & n480 ;
  assign n3424 = \InstQueue_reg[10][7]/NET0131  & n457 ;
  assign n3432 = ~n3423 & ~n3424 ;
  assign n3433 = n3431 & n3432 ;
  assign n3417 = \InstQueue_reg[6][7]/NET0131  & n478 ;
  assign n3418 = \InstQueue_reg[2][7]/NET0131  & n454 ;
  assign n3429 = ~n3417 & ~n3418 ;
  assign n3419 = \InstQueue_reg[0][7]/NET0131  & n488 ;
  assign n3420 = \InstQueue_reg[12][7]/NET0131  & n486 ;
  assign n3430 = ~n3419 & ~n3420 ;
  assign n3434 = n3429 & n3430 ;
  assign n3438 = n3433 & n3434 ;
  assign n3439 = n3437 & n3438 ;
  assign n3440 = n3408 & ~n3439 ;
  assign n3441 = n3153 & n3440 ;
  assign n3442 = \Datai[31]_pad  & n2327 ;
  assign n3449 = ~n3441 & ~n3442 ;
  assign n3450 = ~n3448 & n3449 ;
  assign n3451 = ~n3152 & n3450 ;
  assign n3452 = n948 & ~n3451 ;
  assign n3453 = ~n3117 & ~n3452 ;
  assign n3458 = \EBX_reg[25]/NET0131  & \EBX_reg[26]/NET0131  ;
  assign n3459 = \EBX_reg[21]/NET0131  & \EBX_reg[22]/NET0131  ;
  assign n3460 = \EBX_reg[0]/NET0131  & \EBX_reg[1]/NET0131  ;
  assign n3461 = \EBX_reg[2]/NET0131  & n3460 ;
  assign n3462 = \EBX_reg[3]/NET0131  & n3461 ;
  assign n3463 = \EBX_reg[4]/NET0131  & n3462 ;
  assign n3464 = \EBX_reg[5]/NET0131  & n3463 ;
  assign n3465 = \EBX_reg[6]/NET0131  & n3464 ;
  assign n3466 = \EBX_reg[7]/NET0131  & n3465 ;
  assign n3467 = \EBX_reg[8]/NET0131  & n3466 ;
  assign n3468 = \EBX_reg[9]/NET0131  & n3467 ;
  assign n3469 = \EBX_reg[10]/NET0131  & n3468 ;
  assign n3470 = \EBX_reg[11]/NET0131  & n3469 ;
  assign n3471 = \EBX_reg[12]/NET0131  & n3470 ;
  assign n3472 = \EBX_reg[13]/NET0131  & n3471 ;
  assign n3473 = \EBX_reg[14]/NET0131  & n3472 ;
  assign n3474 = \EBX_reg[15]/NET0131  & n3473 ;
  assign n3475 = \EBX_reg[16]/NET0131  & n3474 ;
  assign n3476 = \EBX_reg[17]/NET0131  & n3475 ;
  assign n3477 = \EBX_reg[18]/NET0131  & \EBX_reg[19]/NET0131  ;
  assign n3478 = \EBX_reg[20]/NET0131  & n3477 ;
  assign n3479 = n3476 & n3478 ;
  assign n3480 = n3459 & n3479 ;
  assign n3481 = \EBX_reg[23]/NET0131  & n3480 ;
  assign n3482 = \EBX_reg[24]/NET0131  & n3481 ;
  assign n3483 = n3458 & n3482 ;
  assign n3484 = n773 & ~n3483 ;
  assign n3454 = n752 & n808 ;
  assign n3485 = ~n752 & n773 ;
  assign n3486 = ~n3454 & ~n3485 ;
  assign n3487 = ~n3484 & ~n3486 ;
  assign n3488 = \EBX_reg[27]/NET0131  & ~n3487 ;
  assign n3455 = ~n3312 & n3343 ;
  assign n3456 = ~n3344 & ~n3455 ;
  assign n3457 = n3454 & n3456 ;
  assign n3489 = ~\EBX_reg[27]/NET0131  & n773 ;
  assign n3490 = n3483 & n3489 ;
  assign n3491 = ~n3457 & ~n3490 ;
  assign n3492 = ~n3488 & n3491 ;
  assign n3493 = n948 & ~n3492 ;
  assign n3494 = \EBX_reg[27]/NET0131  & ~n3116 ;
  assign n3495 = ~n3493 & ~n3494 ;
  assign n3496 = ~n922 & n1997 ;
  assign n3497 = \PhyAddrPointer_reg[4]/NET0131  & ~n3496 ;
  assign n3498 = n748 & n2917 ;
  assign n3499 = ~n3497 & ~n3498 ;
  assign n3500 = ~n2925 & n3499 ;
  assign n3501 = n948 & ~n3500 ;
  assign n3506 = \PhyAddrPointer_reg[1]/NET0131  & \PhyAddrPointer_reg[2]/NET0131  ;
  assign n3507 = \PhyAddrPointer_reg[3]/NET0131  & n3506 ;
  assign n3508 = ~\PhyAddrPointer_reg[4]/NET0131  & ~n3507 ;
  assign n3509 = \PhyAddrPointer_reg[4]/NET0131  & n3507 ;
  assign n3510 = ~n3508 & ~n3509 ;
  assign n3511 = n2039 & n3510 ;
  assign n3505 = \PhyAddrPointer_reg[4]/NET0131  & ~n2003 ;
  assign n3502 = ~\PhyAddrPointer_reg[4]/NET0131  & ~n2005 ;
  assign n3503 = ~n2006 & ~n3502 ;
  assign n3504 = n971 & n3503 ;
  assign n3512 = ~n2901 & ~n3504 ;
  assign n3513 = ~n3505 & n3512 ;
  assign n3514 = ~n3511 & n3513 ;
  assign n3515 = ~n3501 & n3514 ;
  assign n3518 = ~READY_n_pad & ~n1194 ;
  assign n3519 = n864 & ~n3518 ;
  assign n3520 = ~n922 & ~n1714 ;
  assign n3521 = n1890 & n3520 ;
  assign n3522 = ~n3519 & n3521 ;
  assign n3523 = \InstAddrPointer_reg[2]/NET0131  & ~n3522 ;
  assign n3529 = ~n780 & n1449 ;
  assign n3528 = ~n867 & n1194 ;
  assign n3524 = ~\InstAddrPointer_reg[2]/NET0131  & ~n808 ;
  assign n3525 = n808 & n1449 ;
  assign n3526 = ~n3524 & ~n3525 ;
  assign n3527 = ~n756 & n3526 ;
  assign n3530 = ~n1450 & ~n1453 ;
  assign n3532 = n1620 & ~n3530 ;
  assign n3531 = ~n1620 & n3530 ;
  assign n3533 = n930 & ~n3531 ;
  assign n3534 = ~n3532 & n3533 ;
  assign n3535 = ~n1226 & ~n1300 ;
  assign n3537 = n1297 & ~n3535 ;
  assign n3536 = ~n1297 & n3535 ;
  assign n3538 = n929 & ~n3536 ;
  assign n3539 = ~n3537 & n3538 ;
  assign n3540 = ~n3534 & ~n3539 ;
  assign n3541 = ~n3527 & n3540 ;
  assign n3542 = ~n3528 & n3541 ;
  assign n3543 = ~n3529 & n3542 ;
  assign n3544 = ~n3523 & n3543 ;
  assign n3545 = n948 & ~n3544 ;
  assign n3516 = \rEIP_reg[2]/NET0131  & n1731 ;
  assign n3517 = \InstAddrPointer_reg[2]/NET0131  & ~n1736 ;
  assign n3546 = ~n3516 & ~n3517 ;
  assign n3547 = ~n3545 & n3546 ;
  assign n3549 = ~n1451 & ~n1618 ;
  assign n3550 = n929 & ~n3549 ;
  assign n3551 = n930 & n3549 ;
  assign n3552 = ~n3550 & ~n3551 ;
  assign n3553 = ~\InstAddrPointer_reg[0]/NET0131  & n810 ;
  assign n3554 = \InstAddrPointer_reg[0]/NET0131  & n745 ;
  assign n3555 = n925 & n3554 ;
  assign n3556 = ~n3553 & ~n3555 ;
  assign n3557 = n3552 & ~n3556 ;
  assign n3558 = n948 & ~n3557 ;
  assign n3548 = \InstAddrPointer_reg[0]/NET0131  & ~n1736 ;
  assign n3559 = \rEIP_reg[0]/NET0131  & n1731 ;
  assign n3560 = ~n3548 & ~n3559 ;
  assign n3561 = ~n3558 & n3560 ;
  assign n3562 = \EAX_reg[26]/NET0131  & ~n3116 ;
  assign n3565 = n3140 & n3142 ;
  assign n3566 = ~\EAX_reg[26]/NET0131  & ~n3565 ;
  assign n3567 = \EAX_reg[26]/NET0131  & n3565 ;
  assign n3568 = n3118 & ~n3567 ;
  assign n3569 = ~n3566 & n3568 ;
  assign n3570 = \EAX_reg[26]/NET0131  & ~n3447 ;
  assign n3574 = \Datai[26]_pad  & n2327 ;
  assign n3563 = \Datai[10]_pad  & ~READY_n_pad ;
  assign n3564 = n1719 & n3563 ;
  assign n3571 = ~n3280 & n3311 ;
  assign n3572 = ~n3312 & ~n3571 ;
  assign n3573 = n3153 & n3572 ;
  assign n3575 = ~n3564 & ~n3573 ;
  assign n3576 = ~n3574 & n3575 ;
  assign n3577 = ~n3570 & n3576 ;
  assign n3578 = ~n3569 & n3577 ;
  assign n3579 = n948 & ~n3578 ;
  assign n3580 = ~n3562 & ~n3579 ;
  assign n3581 = ~n962 & ~n1731 ;
  assign n3582 = ~n980 & n2037 ;
  assign n3583 = n2793 & n3582 ;
  assign n3584 = n3581 & n3583 ;
  assign n3585 = \uWord_reg[12]/NET0131  & ~n3584 ;
  assign n3588 = ~\EAX_reg[13]/NET0131  & ~\EAX_reg[14]/NET0131  ;
  assign n3589 = ~\EAX_reg[15]/NET0131  & ~\EAX_reg[1]/NET0131  ;
  assign n3596 = n3588 & n3589 ;
  assign n3586 = ~\EAX_reg[0]/NET0131  & ~\EAX_reg[10]/NET0131  ;
  assign n3587 = ~\EAX_reg[11]/NET0131  & ~\EAX_reg[12]/NET0131  ;
  assign n3597 = n3586 & n3587 ;
  assign n3598 = n3596 & n3597 ;
  assign n3592 = ~\EAX_reg[6]/NET0131  & ~\EAX_reg[7]/NET0131  ;
  assign n3593 = ~\EAX_reg[8]/NET0131  & ~\EAX_reg[9]/NET0131  ;
  assign n3594 = n3592 & n3593 ;
  assign n3590 = ~\EAX_reg[2]/NET0131  & ~\EAX_reg[3]/NET0131  ;
  assign n3591 = ~\EAX_reg[4]/NET0131  & ~\EAX_reg[5]/NET0131  ;
  assign n3595 = n3590 & n3591 ;
  assign n3599 = n3594 & n3595 ;
  assign n3600 = n3598 & n3599 ;
  assign n3601 = \EAX_reg[31]/NET0131  & ~n3600 ;
  assign n3602 = \EAX_reg[16]/NET0131  & n3601 ;
  assign n3603 = \EAX_reg[17]/NET0131  & n3602 ;
  assign n3604 = \EAX_reg[18]/NET0131  & n3603 ;
  assign n3605 = \EAX_reg[19]/NET0131  & n3604 ;
  assign n3606 = n3139 & n3605 ;
  assign n3607 = n3141 & n3606 ;
  assign n3608 = \EAX_reg[25]/NET0131  & n3607 ;
  assign n3609 = \EAX_reg[26]/NET0131  & n3608 ;
  assign n3610 = \EAX_reg[27]/NET0131  & n3609 ;
  assign n3611 = ~\EAX_reg[28]/NET0131  & ~n3610 ;
  assign n3612 = \EAX_reg[28]/NET0131  & n3610 ;
  assign n3613 = ~n3611 & ~n3612 ;
  assign n3614 = n742 & n3613 ;
  assign n3615 = \Datai[12]_pad  & n736 ;
  assign n3616 = ~READY_n_pad & n3615 ;
  assign n3617 = ~n3614 & ~n3616 ;
  assign n3618 = n825 & ~n3617 ;
  assign n3619 = ~n736 & ~n742 ;
  assign n3620 = n825 & ~n3619 ;
  assign n3621 = ~n1975 & n3620 ;
  assign n3622 = \uWord_reg[12]/NET0131  & ~n3621 ;
  assign n3623 = ~n3618 & ~n3622 ;
  assign n3624 = n948 & ~n3623 ;
  assign n3625 = ~n3585 & ~n3624 ;
  assign n3627 = n816 & n948 ;
  assign n3628 = ~n956 & ~n981 ;
  assign n3629 = n1734 & n3628 ;
  assign n3630 = n3581 & n3629 ;
  assign n3631 = \InstQueueRd_Addr_reg[0]/NET0131  & ~n3630 ;
  assign n3626 = ~\InstQueueRd_Addr_reg[0]/NET0131  & n993 ;
  assign n3632 = \Flush_reg/NET0131  & \InstAddrPointer_reg[0]/NET0131  ;
  assign n3633 = ~\Flush_reg/NET0131  & ~\InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n3634 = ~n3632 & ~n3633 ;
  assign n3635 = n984 & n3634 ;
  assign n3636 = ~n3626 & ~n3635 ;
  assign n3637 = ~n3631 & n3636 ;
  assign n3638 = ~n3627 & n3637 ;
  assign n3643 = ~n910 & n948 ;
  assign n3644 = \InstAddrPointer_reg[31]/NET0131  & ~n1455 ;
  assign n3645 = ~\InstAddrPointer_reg[1]/NET0131  & ~\InstAddrPointer_reg[31]/NET0131  ;
  assign n3646 = ~n3644 & ~n3645 ;
  assign n3647 = n3632 & n3646 ;
  assign n3648 = ~n985 & ~n3647 ;
  assign n3649 = n984 & ~n3648 ;
  assign n3639 = ~n969 & ~n981 ;
  assign n3640 = ~n951 & n3581 ;
  assign n3641 = n3639 & n3640 ;
  assign n3642 = \InstQueueRd_Addr_reg[2]/NET0131  & ~n3641 ;
  assign n3650 = n884 & n993 ;
  assign n3651 = ~n3642 & ~n3650 ;
  assign n3652 = ~n3649 & n3651 ;
  assign n3653 = ~n3643 & n3652 ;
  assign n3654 = \PhyAddrPointer_reg[3]/NET0131  & ~n921 ;
  assign n3655 = ~n3075 & ~n3654 ;
  assign n3656 = n748 & ~n3655 ;
  assign n3657 = \PhyAddrPointer_reg[3]/NET0131  & ~n1997 ;
  assign n3658 = ~n3053 & ~n3657 ;
  assign n3659 = ~n3656 & n3658 ;
  assign n3660 = n948 & ~n3659 ;
  assign n3661 = \PhyAddrPointer_reg[2]/NET0131  & ~n2366 ;
  assign n3662 = n952 & n3661 ;
  assign n3663 = ~\PhyAddrPointer_reg[3]/NET0131  & ~n3662 ;
  assign n3665 = n952 & ~n3661 ;
  assign n3664 = ~n993 & n2002 ;
  assign n3666 = \PhyAddrPointer_reg[3]/NET0131  & n3664 ;
  assign n3667 = ~n3665 & n3666 ;
  assign n3668 = ~n3663 & ~n3667 ;
  assign n3670 = ~\PhyAddrPointer_reg[3]/NET0131  & ~n3506 ;
  assign n3671 = ~n3507 & ~n3670 ;
  assign n3672 = n970 & n3671 ;
  assign n3669 = \PhyAddrPointer_reg[3]/NET0131  & n981 ;
  assign n3673 = ~n3045 & ~n3669 ;
  assign n3674 = ~n3672 & n3673 ;
  assign n3675 = ~n3668 & n3674 ;
  assign n3676 = ~n3660 & n3675 ;
  assign n3680 = \PhyAddrPointer_reg[5]/NET0131  & ~n921 ;
  assign n3681 = ~n3094 & ~n3680 ;
  assign n3682 = n748 & ~n3681 ;
  assign n3683 = \PhyAddrPointer_reg[5]/NET0131  & ~n1997 ;
  assign n3684 = ~n3105 & ~n3683 ;
  assign n3685 = ~n3682 & n3684 ;
  assign n3686 = n948 & ~n3685 ;
  assign n3677 = ~\PhyAddrPointer_reg[5]/NET0131  & ~n3509 ;
  assign n3678 = ~n3004 & ~n3677 ;
  assign n3687 = ~\DataWidth_reg[1]/NET0131  & ~n3678 ;
  assign n3688 = ~\PhyAddrPointer_reg[5]/NET0131  & ~n2006 ;
  assign n3689 = ~n2007 & ~n3688 ;
  assign n3690 = \DataWidth_reg[1]/NET0131  & ~n3689 ;
  assign n3691 = n952 & ~n3690 ;
  assign n3692 = ~n3687 & n3691 ;
  assign n3679 = n970 & n3678 ;
  assign n3693 = \PhyAddrPointer_reg[5]/NET0131  & ~n2003 ;
  assign n3694 = ~n3087 & ~n3693 ;
  assign n3695 = ~n3679 & n3694 ;
  assign n3696 = ~n3692 & n3695 ;
  assign n3697 = ~n3686 & n3696 ;
  assign n3701 = \PhyAddrPointer_reg[6]/NET0131  & ~n921 ;
  assign n3702 = ~n2953 & ~n3701 ;
  assign n3703 = n748 & ~n3702 ;
  assign n3704 = \PhyAddrPointer_reg[6]/NET0131  & ~n1997 ;
  assign n3705 = ~n2961 & ~n3704 ;
  assign n3706 = ~n3703 & n3705 ;
  assign n3707 = n948 & ~n3706 ;
  assign n3709 = n2007 & ~n2366 ;
  assign n3710 = ~\PhyAddrPointer_reg[6]/NET0131  & ~n3709 ;
  assign n3708 = n2008 & ~n2366 ;
  assign n3711 = n952 & ~n3708 ;
  assign n3712 = ~n3710 & n3711 ;
  assign n3698 = ~\PhyAddrPointer_reg[6]/NET0131  & ~n3004 ;
  assign n3699 = ~n3005 & ~n3698 ;
  assign n3700 = n970 & n3699 ;
  assign n3713 = \PhyAddrPointer_reg[6]/NET0131  & ~n2003 ;
  assign n3714 = ~n2934 & ~n3713 ;
  assign n3715 = ~n3700 & n3714 ;
  assign n3716 = ~n3712 & n3715 ;
  assign n3717 = ~n3707 & n3716 ;
  assign n3720 = ~n922 & n1937 ;
  assign n3721 = \InstAddrPointer_reg[1]/NET0131  & ~n3720 ;
  assign n3719 = ~n810 & n1455 ;
  assign n3724 = ~n1456 & ~n1617 ;
  assign n3725 = ~n1451 & n3724 ;
  assign n3722 = ~n1262 & ~n1263 ;
  assign n3723 = n1451 & ~n3722 ;
  assign n3726 = ~n1051 & ~n3723 ;
  assign n3727 = ~n3725 & n3726 ;
  assign n3729 = n1295 & n3722 ;
  assign n3728 = ~n1295 & ~n3722 ;
  assign n3730 = n1051 & ~n3728 ;
  assign n3731 = ~n3729 & n3730 ;
  assign n3732 = ~n3727 & ~n3731 ;
  assign n3733 = n929 & ~n3732 ;
  assign n3735 = n1618 & ~n3722 ;
  assign n3734 = ~n1618 & ~n3724 ;
  assign n3736 = n930 & ~n3734 ;
  assign n3737 = ~n3735 & n3736 ;
  assign n3738 = ~n3733 & ~n3737 ;
  assign n3739 = ~\InstAddrPointer_reg[1]/NET0131  & ~n867 ;
  assign n3740 = n3738 & ~n3739 ;
  assign n3741 = ~n3719 & n3740 ;
  assign n3742 = ~n3721 & n3741 ;
  assign n3743 = n948 & ~n3742 ;
  assign n3718 = \rEIP_reg[1]/NET0131  & n1731 ;
  assign n3744 = \InstAddrPointer_reg[1]/NET0131  & ~n1736 ;
  assign n3745 = ~n3718 & ~n3744 ;
  assign n3746 = ~n3743 & n3745 ;
  assign n3748 = ~n849 & n948 ;
  assign n3749 = ~\Flush_reg/NET0131  & \InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n3750 = n3632 & ~n3646 ;
  assign n3751 = ~n3749 & ~n3750 ;
  assign n3752 = n984 & ~n3751 ;
  assign n3747 = \InstQueueRd_Addr_reg[1]/NET0131  & ~n3641 ;
  assign n3753 = ~n819 & n993 ;
  assign n3754 = ~n3747 & ~n3753 ;
  assign n3755 = ~n3752 & n3754 ;
  assign n3756 = ~n3748 & n3755 ;
  assign n3757 = \EAX_reg[29]/NET0131  & ~n3116 ;
  assign n3758 = \EAX_reg[28]/NET0131  & n3145 ;
  assign n3759 = n3118 & ~n3758 ;
  assign n3760 = n3446 & ~n3759 ;
  assign n3761 = \EAX_reg[29]/NET0131  & ~n3760 ;
  assign n3762 = ~\EAX_reg[29]/NET0131  & n3118 ;
  assign n3763 = n3758 & n3762 ;
  assign n3764 = ~n3376 & n3407 ;
  assign n3765 = ~n3408 & ~n3764 ;
  assign n3766 = n3153 & n3765 ;
  assign n3767 = \Datai[13]_pad  & n826 ;
  assign n3768 = n736 & n3767 ;
  assign n3770 = ~\Datai[29]_pad  & n826 ;
  assign n3769 = ~\EAX_reg[29]/NET0131  & ~n826 ;
  assign n3771 = n835 & ~n3769 ;
  assign n3772 = ~n3770 & n3771 ;
  assign n3773 = ~n3768 & ~n3772 ;
  assign n3774 = ~n3766 & n3773 ;
  assign n3775 = ~n3763 & n3774 ;
  assign n3776 = ~n3761 & n3775 ;
  assign n3777 = n948 & ~n3776 ;
  assign n3778 = ~n3757 & ~n3777 ;
  assign n3781 = \EBX_reg[18]/NET0131  & n3476 ;
  assign n3782 = \EBX_reg[19]/NET0131  & n3781 ;
  assign n3783 = \EBX_reg[20]/NET0131  & \EBX_reg[23]/NET0131  ;
  assign n3784 = n3459 & n3783 ;
  assign n3785 = n3782 & n3784 ;
  assign n3786 = \EBX_reg[24]/NET0131  & n3785 ;
  assign n3788 = \EBX_reg[25]/NET0131  & n3786 ;
  assign n3789 = ~\EBX_reg[26]/NET0131  & ~n3788 ;
  assign n3787 = n3458 & n3786 ;
  assign n3790 = n773 & ~n3787 ;
  assign n3791 = ~n3789 & n3790 ;
  assign n3779 = n3454 & n3572 ;
  assign n3780 = \EBX_reg[26]/NET0131  & n3486 ;
  assign n3792 = ~n3779 & ~n3780 ;
  assign n3793 = ~n3791 & n3792 ;
  assign n3794 = n948 & ~n3793 ;
  assign n3795 = \EBX_reg[26]/NET0131  & ~n3116 ;
  assign n3796 = ~n3794 & ~n3795 ;
  assign n3798 = n742 & n825 ;
  assign n3799 = \EAX_reg[23]/NET0131  & n3606 ;
  assign n3800 = ~\EAX_reg[24]/NET0131  & ~n3799 ;
  assign n3801 = ~n3607 & ~n3800 ;
  assign n3802 = ~n833 & ~n3801 ;
  assign n3803 = n3798 & ~n3802 ;
  assign n3804 = n825 & ~n828 ;
  assign n3805 = n827 & n833 ;
  assign n3806 = n3804 & ~n3805 ;
  assign n3807 = ~n3803 & n3806 ;
  assign n3808 = \Datao[24]_pad  & ~n3807 ;
  assign n3809 = n742 & n3801 ;
  assign n3810 = n895 & n3809 ;
  assign n3811 = ~n3808 & ~n3810 ;
  assign n3812 = n948 & ~n3811 ;
  assign n3797 = \uWord_reg[8]/NET0131  & n956 ;
  assign n3813 = \State2_reg[1]/NET0131  & \State2_reg[3]/NET0131  ;
  assign n3814 = \State2_reg[2]/NET0131  & ~n970 ;
  assign n3815 = ~n3813 & ~n3814 ;
  assign n3816 = ~n984 & ~n3815 ;
  assign n3817 = \Datao[24]_pad  & ~n3816 ;
  assign n3818 = ~n3797 & ~n3817 ;
  assign n3819 = ~n3812 & n3818 ;
  assign n3821 = ~n833 & ~n3613 ;
  assign n3822 = n3798 & ~n3821 ;
  assign n3823 = n3806 & ~n3822 ;
  assign n3824 = \Datao[28]_pad  & ~n3823 ;
  assign n3825 = n895 & n3614 ;
  assign n3826 = ~n3824 & ~n3825 ;
  assign n3827 = n948 & ~n3826 ;
  assign n3820 = \uWord_reg[12]/NET0131  & n956 ;
  assign n3828 = \Datao[28]_pad  & ~n3816 ;
  assign n3829 = ~n3820 & ~n3828 ;
  assign n3830 = ~n3827 & n3829 ;
  assign n3832 = ~n882 & n948 ;
  assign n3833 = ~\Flush_reg/NET0131  & \InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n3834 = ~n3647 & ~n3833 ;
  assign n3835 = n984 & ~n3834 ;
  assign n3831 = \InstQueueRd_Addr_reg[3]/NET0131  & ~n3641 ;
  assign n3836 = ~n855 & n993 ;
  assign n3837 = ~n3831 & ~n3836 ;
  assign n3838 = ~n3835 & n3837 ;
  assign n3839 = ~n3832 & n3838 ;
  assign n3840 = n948 & ~n3621 ;
  assign n3841 = n3584 & ~n3840 ;
  assign n3842 = \uWord_reg[8]/NET0131  & ~n3841 ;
  assign n3843 = n825 & n948 ;
  assign n3844 = \Datai[8]_pad  & n736 ;
  assign n3845 = ~READY_n_pad & n3844 ;
  assign n3846 = ~n3809 & ~n3845 ;
  assign n3847 = n3843 & ~n3846 ;
  assign n3848 = ~n3842 & ~n3847 ;
  assign n3851 = \EBX_reg[27]/NET0131  & \EBX_reg[28]/NET0131  ;
  assign n3852 = n3483 & n3851 ;
  assign n3854 = \EBX_reg[29]/NET0131  & n3852 ;
  assign n3853 = ~\EBX_reg[29]/NET0131  & ~n3852 ;
  assign n3855 = n773 & ~n3853 ;
  assign n3856 = ~n3854 & n3855 ;
  assign n3849 = \EBX_reg[29]/NET0131  & n3486 ;
  assign n3850 = n3454 & n3765 ;
  assign n3857 = ~n3849 & ~n3850 ;
  assign n3858 = ~n3856 & n3857 ;
  assign n3859 = n948 & ~n3858 ;
  assign n3860 = \EBX_reg[29]/NET0131  & ~n3116 ;
  assign n3861 = ~n3859 & ~n3860 ;
  assign n3874 = \InstQueueWr_Addr_reg[0]/NET0131  & ~\InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3875 = \InstQueueWr_Addr_reg[2]/NET0131  & n3874 ;
  assign n3876 = \InstQueueWr_Addr_reg[3]/NET0131  & n3875 ;
  assign n3879 = ~\Datai[13]_pad  & ~\Datai[14]_pad  ;
  assign n3880 = ~\Datai[15]_pad  & ~\Datai[1]_pad  ;
  assign n3887 = n3879 & n3880 ;
  assign n3877 = ~\Datai[0]_pad  & ~\Datai[10]_pad  ;
  assign n3878 = ~\Datai[11]_pad  & ~\Datai[12]_pad  ;
  assign n3888 = n3877 & n3878 ;
  assign n3889 = n3887 & n3888 ;
  assign n3883 = ~\Datai[6]_pad  & ~\Datai[7]_pad  ;
  assign n3884 = ~\Datai[8]_pad  & ~\Datai[9]_pad  ;
  assign n3885 = n3883 & n3884 ;
  assign n3881 = ~\Datai[2]_pad  & ~\Datai[3]_pad  ;
  assign n3882 = ~\Datai[4]_pad  & ~\Datai[5]_pad  ;
  assign n3886 = n3881 & n3882 ;
  assign n3890 = n3885 & n3886 ;
  assign n3891 = n3889 & n3890 ;
  assign n3894 = ~\Datai[20]_pad  & ~\Datai[21]_pad  ;
  assign n3895 = ~\Datai[22]_pad  & ~\Datai[23]_pad  ;
  assign n3896 = n3894 & n3895 ;
  assign n3892 = ~\Datai[16]_pad  & ~\Datai[17]_pad  ;
  assign n3893 = ~\Datai[18]_pad  & ~\Datai[19]_pad  ;
  assign n3897 = n3892 & n3893 ;
  assign n3898 = n3896 & n3897 ;
  assign n3899 = n3891 & n3898 ;
  assign n3900 = \Datai[31]_pad  & ~n3899 ;
  assign n3901 = \Datai[24]_pad  & n3900 ;
  assign n3902 = \Datai[25]_pad  & n3901 ;
  assign n3903 = \Datai[26]_pad  & n3902 ;
  assign n3904 = \Datai[27]_pad  & n3903 ;
  assign n3905 = \Datai[28]_pad  & n3904 ;
  assign n3906 = ~\Datai[28]_pad  & ~n3904 ;
  assign n3907 = ~n3905 & ~n3906 ;
  assign n3908 = n3876 & n3907 ;
  assign n3909 = \Datai[31]_pad  & ~n3891 ;
  assign n3910 = \Datai[16]_pad  & n3909 ;
  assign n3911 = \Datai[17]_pad  & n3910 ;
  assign n3912 = \Datai[18]_pad  & n3911 ;
  assign n3913 = \Datai[19]_pad  & n3912 ;
  assign n3914 = ~\Datai[20]_pad  & ~n3913 ;
  assign n3915 = \Datai[20]_pad  & n3913 ;
  assign n3916 = ~n3914 & ~n3915 ;
  assign n3917 = ~\InstQueueWr_Addr_reg[0]/NET0131  & \InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3918 = \InstQueueWr_Addr_reg[2]/NET0131  & n3917 ;
  assign n3919 = \InstQueueWr_Addr_reg[3]/NET0131  & n3918 ;
  assign n3920 = n3916 & n3919 ;
  assign n3921 = ~n3908 & ~n3920 ;
  assign n3922 = \DataWidth_reg[1]/NET0131  & ~n3921 ;
  assign n3862 = ~\InstQueueWr_Addr_reg[0]/NET0131  & ~\InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3863 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3862 ;
  assign n3864 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3863 ;
  assign n3865 = \InstQueueWr_Addr_reg[0]/NET0131  & \InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3866 = \InstQueueWr_Addr_reg[2]/NET0131  & n3865 ;
  assign n3867 = \InstQueueWr_Addr_reg[3]/NET0131  & n3866 ;
  assign n3868 = ~n3864 & ~n3867 ;
  assign n3869 = \Datai[4]_pad  & ~n3868 ;
  assign n3870 = \InstQueue_reg[0][4]/NET0131  & ~n3864 ;
  assign n3871 = ~n3867 & n3870 ;
  assign n3872 = ~n3869 & ~n3871 ;
  assign n3923 = ~n3876 & ~n3919 ;
  assign n3924 = \DataWidth_reg[1]/NET0131  & ~n3923 ;
  assign n3925 = ~n3872 & ~n3924 ;
  assign n3926 = ~n3922 & ~n3925 ;
  assign n3927 = n952 & ~n3926 ;
  assign n3928 = ~n733 & n3864 ;
  assign n3929 = ~n3870 & ~n3928 ;
  assign n3930 = n993 & ~n3929 ;
  assign n3873 = n970 & ~n3872 ;
  assign n3931 = ~n948 & ~n961 ;
  assign n3932 = ~n1731 & n3931 ;
  assign n3933 = n2793 & n3932 ;
  assign n3934 = \InstQueue_reg[0][4]/NET0131  & ~n3933 ;
  assign n3935 = ~n3873 & ~n3934 ;
  assign n3936 = ~n3930 & n3935 ;
  assign n3937 = ~n3927 & n3936 ;
  assign n3948 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3866 ;
  assign n3949 = n3907 & n3948 ;
  assign n3950 = \InstQueueWr_Addr_reg[3]/NET0131  & n3863 ;
  assign n3951 = n3916 & n3950 ;
  assign n3952 = ~n3949 & ~n3951 ;
  assign n3953 = \DataWidth_reg[1]/NET0131  & ~n3952 ;
  assign n3938 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3917 ;
  assign n3939 = \InstQueueWr_Addr_reg[3]/NET0131  & n3938 ;
  assign n3940 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3874 ;
  assign n3941 = \InstQueueWr_Addr_reg[3]/NET0131  & n3940 ;
  assign n3942 = ~n3939 & ~n3941 ;
  assign n3943 = \Datai[4]_pad  & ~n3942 ;
  assign n3944 = \InstQueue_reg[10][4]/NET0131  & ~n3939 ;
  assign n3945 = ~n3941 & n3944 ;
  assign n3946 = ~n3943 & ~n3945 ;
  assign n3954 = ~n3948 & ~n3950 ;
  assign n3955 = \DataWidth_reg[1]/NET0131  & ~n3954 ;
  assign n3956 = ~n3946 & ~n3955 ;
  assign n3957 = ~n3953 & ~n3956 ;
  assign n3958 = n952 & ~n3957 ;
  assign n3959 = ~n733 & n3939 ;
  assign n3960 = ~n3944 & ~n3959 ;
  assign n3961 = n993 & ~n3960 ;
  assign n3947 = n970 & ~n3946 ;
  assign n3962 = \InstQueue_reg[10][4]/NET0131  & ~n3933 ;
  assign n3963 = ~n3947 & ~n3962 ;
  assign n3964 = ~n3961 & n3963 ;
  assign n3965 = ~n3958 & n3964 ;
  assign n3974 = n3907 & n3950 ;
  assign n3975 = n3916 & n3941 ;
  assign n3976 = ~n3974 & ~n3975 ;
  assign n3977 = \DataWidth_reg[1]/NET0131  & ~n3976 ;
  assign n3966 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3865 ;
  assign n3967 = \InstQueueWr_Addr_reg[3]/NET0131  & n3966 ;
  assign n3968 = ~n3939 & ~n3967 ;
  assign n3969 = \Datai[4]_pad  & ~n3968 ;
  assign n3970 = \InstQueue_reg[11][4]/NET0131  & ~n3967 ;
  assign n3971 = ~n3939 & n3970 ;
  assign n3972 = ~n3969 & ~n3971 ;
  assign n3978 = ~n3941 & ~n3950 ;
  assign n3979 = \DataWidth_reg[1]/NET0131  & ~n3978 ;
  assign n3980 = ~n3972 & ~n3979 ;
  assign n3981 = ~n3977 & ~n3980 ;
  assign n3982 = n952 & ~n3981 ;
  assign n3983 = ~n733 & n3967 ;
  assign n3984 = ~n3970 & ~n3983 ;
  assign n3985 = n993 & ~n3984 ;
  assign n3973 = n970 & ~n3972 ;
  assign n3986 = \InstQueue_reg[11][4]/NET0131  & ~n3933 ;
  assign n3987 = ~n3973 & ~n3986 ;
  assign n3988 = ~n3985 & n3987 ;
  assign n3989 = ~n3982 & n3988 ;
  assign n3998 = n3907 & n3941 ;
  assign n3999 = n3916 & n3939 ;
  assign n4000 = ~n3998 & ~n3999 ;
  assign n4001 = \DataWidth_reg[1]/NET0131  & ~n4000 ;
  assign n3990 = \InstQueueWr_Addr_reg[2]/NET0131  & n3862 ;
  assign n3991 = \InstQueueWr_Addr_reg[3]/NET0131  & n3990 ;
  assign n3992 = ~n3967 & ~n3991 ;
  assign n3993 = \Datai[4]_pad  & ~n3992 ;
  assign n3994 = \InstQueue_reg[12][4]/NET0131  & ~n3991 ;
  assign n3995 = ~n3967 & n3994 ;
  assign n3996 = ~n3993 & ~n3995 ;
  assign n4002 = \DataWidth_reg[1]/NET0131  & ~n3942 ;
  assign n4003 = ~n3996 & ~n4002 ;
  assign n4004 = ~n4001 & ~n4003 ;
  assign n4005 = n952 & ~n4004 ;
  assign n4006 = ~n733 & n3991 ;
  assign n4007 = ~n3994 & ~n4006 ;
  assign n4008 = n993 & ~n4007 ;
  assign n3997 = n970 & ~n3996 ;
  assign n4009 = \InstQueue_reg[12][4]/NET0131  & ~n3933 ;
  assign n4010 = ~n3997 & ~n4009 ;
  assign n4011 = ~n4008 & n4010 ;
  assign n4012 = ~n4005 & n4011 ;
  assign n4019 = n3907 & n3939 ;
  assign n4020 = n3916 & n3967 ;
  assign n4021 = ~n4019 & ~n4020 ;
  assign n4022 = \DataWidth_reg[1]/NET0131  & ~n4021 ;
  assign n4013 = ~n3876 & ~n3991 ;
  assign n4014 = \Datai[4]_pad  & ~n4013 ;
  assign n4015 = \InstQueue_reg[13][4]/NET0131  & ~n3876 ;
  assign n4016 = ~n3991 & n4015 ;
  assign n4017 = ~n4014 & ~n4016 ;
  assign n4023 = \DataWidth_reg[1]/NET0131  & ~n3968 ;
  assign n4024 = ~n4017 & ~n4023 ;
  assign n4025 = ~n4022 & ~n4024 ;
  assign n4026 = n952 & ~n4025 ;
  assign n4027 = ~n733 & n3876 ;
  assign n4028 = ~n4015 & ~n4027 ;
  assign n4029 = n993 & ~n4028 ;
  assign n4018 = n970 & ~n4017 ;
  assign n4030 = \InstQueue_reg[13][4]/NET0131  & ~n3933 ;
  assign n4031 = ~n4018 & ~n4030 ;
  assign n4032 = ~n4029 & n4031 ;
  assign n4033 = ~n4026 & n4032 ;
  assign n4039 = n3907 & n3967 ;
  assign n4040 = n3916 & n3991 ;
  assign n4041 = ~n4039 & ~n4040 ;
  assign n4042 = \DataWidth_reg[1]/NET0131  & ~n4041 ;
  assign n4034 = \Datai[4]_pad  & ~n3923 ;
  assign n4035 = \InstQueue_reg[14][4]/NET0131  & ~n3919 ;
  assign n4036 = ~n3876 & n4035 ;
  assign n4037 = ~n4034 & ~n4036 ;
  assign n4043 = \DataWidth_reg[1]/NET0131  & ~n3992 ;
  assign n4044 = ~n4037 & ~n4043 ;
  assign n4045 = ~n4042 & ~n4044 ;
  assign n4046 = n952 & ~n4045 ;
  assign n4047 = ~n733 & n3919 ;
  assign n4048 = ~n4035 & ~n4047 ;
  assign n4049 = n993 & ~n4048 ;
  assign n4038 = n970 & ~n4037 ;
  assign n4050 = \InstQueue_reg[14][4]/NET0131  & ~n3933 ;
  assign n4051 = ~n4038 & ~n4050 ;
  assign n4052 = ~n4049 & n4051 ;
  assign n4053 = ~n4046 & n4052 ;
  assign n4060 = n3907 & n3991 ;
  assign n4061 = n3876 & n3916 ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = \DataWidth_reg[1]/NET0131  & ~n4062 ;
  assign n4054 = ~n3867 & ~n3919 ;
  assign n4055 = \Datai[4]_pad  & ~n4054 ;
  assign n4056 = \InstQueue_reg[15][4]/NET0131  & ~n3867 ;
  assign n4057 = ~n3919 & n4056 ;
  assign n4058 = ~n4055 & ~n4057 ;
  assign n4064 = \DataWidth_reg[1]/NET0131  & ~n4013 ;
  assign n4065 = ~n4058 & ~n4064 ;
  assign n4066 = ~n4063 & ~n4065 ;
  assign n4067 = n952 & ~n4066 ;
  assign n4068 = ~n733 & n3867 ;
  assign n4069 = ~n4056 & ~n4068 ;
  assign n4070 = n993 & ~n4069 ;
  assign n4059 = n970 & ~n4058 ;
  assign n4071 = \InstQueue_reg[15][4]/NET0131  & ~n3933 ;
  assign n4072 = ~n4059 & ~n4071 ;
  assign n4073 = ~n4070 & n4072 ;
  assign n4074 = ~n4067 & n4073 ;
  assign n4082 = n3907 & n3919 ;
  assign n4083 = n3867 & n3916 ;
  assign n4084 = ~n4082 & ~n4083 ;
  assign n4085 = \DataWidth_reg[1]/NET0131  & ~n4084 ;
  assign n4075 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3940 ;
  assign n4076 = ~n3864 & ~n4075 ;
  assign n4077 = \Datai[4]_pad  & ~n4076 ;
  assign n4078 = \InstQueue_reg[1][4]/NET0131  & ~n4075 ;
  assign n4079 = ~n3864 & n4078 ;
  assign n4080 = ~n4077 & ~n4079 ;
  assign n4086 = \DataWidth_reg[1]/NET0131  & ~n4054 ;
  assign n4087 = ~n4080 & ~n4086 ;
  assign n4088 = ~n4085 & ~n4087 ;
  assign n4089 = n952 & ~n4088 ;
  assign n4090 = ~n733 & n4075 ;
  assign n4091 = ~n4078 & ~n4090 ;
  assign n4092 = n993 & ~n4091 ;
  assign n4081 = n970 & ~n4080 ;
  assign n4093 = \InstQueue_reg[1][4]/NET0131  & ~n3933 ;
  assign n4094 = ~n4081 & ~n4093 ;
  assign n4095 = ~n4092 & n4094 ;
  assign n4096 = ~n4089 & n4095 ;
  assign n4104 = n3864 & n3916 ;
  assign n4105 = n3867 & n3907 ;
  assign n4106 = ~n4104 & ~n4105 ;
  assign n4107 = \DataWidth_reg[1]/NET0131  & ~n4106 ;
  assign n4097 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3938 ;
  assign n4098 = ~n4075 & ~n4097 ;
  assign n4099 = \Datai[4]_pad  & ~n4098 ;
  assign n4100 = \InstQueue_reg[2][4]/NET0131  & ~n4097 ;
  assign n4101 = ~n4075 & n4100 ;
  assign n4102 = ~n4099 & ~n4101 ;
  assign n4108 = \DataWidth_reg[1]/NET0131  & ~n3868 ;
  assign n4109 = ~n4102 & ~n4108 ;
  assign n4110 = ~n4107 & ~n4109 ;
  assign n4111 = n952 & ~n4110 ;
  assign n4112 = ~n733 & n4097 ;
  assign n4113 = ~n4100 & ~n4112 ;
  assign n4114 = n993 & ~n4113 ;
  assign n4103 = n970 & ~n4102 ;
  assign n4115 = \InstQueue_reg[2][4]/NET0131  & ~n3933 ;
  assign n4116 = ~n4103 & ~n4115 ;
  assign n4117 = ~n4114 & n4116 ;
  assign n4118 = ~n4111 & n4117 ;
  assign n4126 = n3864 & n3907 ;
  assign n4127 = n3916 & n4075 ;
  assign n4128 = ~n4126 & ~n4127 ;
  assign n4129 = \DataWidth_reg[1]/NET0131  & ~n4128 ;
  assign n4119 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3966 ;
  assign n4120 = ~n4097 & ~n4119 ;
  assign n4121 = \Datai[4]_pad  & ~n4120 ;
  assign n4122 = \InstQueue_reg[3][4]/NET0131  & ~n4119 ;
  assign n4123 = ~n4097 & n4122 ;
  assign n4124 = ~n4121 & ~n4123 ;
  assign n4130 = \DataWidth_reg[1]/NET0131  & ~n4076 ;
  assign n4131 = ~n4124 & ~n4130 ;
  assign n4132 = ~n4129 & ~n4131 ;
  assign n4133 = n952 & ~n4132 ;
  assign n4134 = ~n733 & n4119 ;
  assign n4135 = ~n4122 & ~n4134 ;
  assign n4136 = n993 & ~n4135 ;
  assign n4125 = n970 & ~n4124 ;
  assign n4137 = \InstQueue_reg[3][4]/NET0131  & ~n3933 ;
  assign n4138 = ~n4125 & ~n4137 ;
  assign n4139 = ~n4136 & n4138 ;
  assign n4140 = ~n4133 & n4139 ;
  assign n4148 = n3907 & n4075 ;
  assign n4149 = n3916 & n4097 ;
  assign n4150 = ~n4148 & ~n4149 ;
  assign n4151 = \DataWidth_reg[1]/NET0131  & ~n4150 ;
  assign n4141 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3990 ;
  assign n4142 = ~n4119 & ~n4141 ;
  assign n4143 = \Datai[4]_pad  & ~n4142 ;
  assign n4144 = \InstQueue_reg[4][4]/NET0131  & ~n4141 ;
  assign n4145 = ~n4119 & n4144 ;
  assign n4146 = ~n4143 & ~n4145 ;
  assign n4152 = \DataWidth_reg[1]/NET0131  & ~n4098 ;
  assign n4153 = ~n4146 & ~n4152 ;
  assign n4154 = ~n4151 & ~n4153 ;
  assign n4155 = n952 & ~n4154 ;
  assign n4156 = ~n733 & n4141 ;
  assign n4157 = ~n4144 & ~n4156 ;
  assign n4158 = n993 & ~n4157 ;
  assign n4147 = n970 & ~n4146 ;
  assign n4159 = \InstQueue_reg[4][4]/NET0131  & ~n3933 ;
  assign n4160 = ~n4147 & ~n4159 ;
  assign n4161 = ~n4158 & n4160 ;
  assign n4162 = ~n4155 & n4161 ;
  assign n4170 = n3907 & n4097 ;
  assign n4171 = n3916 & n4119 ;
  assign n4172 = ~n4170 & ~n4171 ;
  assign n4173 = \DataWidth_reg[1]/NET0131  & ~n4172 ;
  assign n4163 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3875 ;
  assign n4164 = ~n4141 & ~n4163 ;
  assign n4165 = \Datai[4]_pad  & ~n4164 ;
  assign n4166 = \InstQueue_reg[5][4]/NET0131  & ~n4163 ;
  assign n4167 = ~n4141 & n4166 ;
  assign n4168 = ~n4165 & ~n4167 ;
  assign n4174 = \DataWidth_reg[1]/NET0131  & ~n4120 ;
  assign n4175 = ~n4168 & ~n4174 ;
  assign n4176 = ~n4173 & ~n4175 ;
  assign n4177 = n952 & ~n4176 ;
  assign n4178 = ~n733 & n4163 ;
  assign n4179 = ~n4166 & ~n4178 ;
  assign n4180 = n993 & ~n4179 ;
  assign n4169 = n970 & ~n4168 ;
  assign n4181 = \InstQueue_reg[5][4]/NET0131  & ~n3933 ;
  assign n4182 = ~n4169 & ~n4181 ;
  assign n4183 = ~n4180 & n4182 ;
  assign n4184 = ~n4177 & n4183 ;
  assign n4192 = n3907 & n4119 ;
  assign n4193 = n3916 & n4141 ;
  assign n4194 = ~n4192 & ~n4193 ;
  assign n4195 = \DataWidth_reg[1]/NET0131  & ~n4194 ;
  assign n4185 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3918 ;
  assign n4186 = ~n4163 & ~n4185 ;
  assign n4187 = \Datai[4]_pad  & ~n4186 ;
  assign n4188 = \InstQueue_reg[6][4]/NET0131  & ~n4185 ;
  assign n4189 = ~n4163 & n4188 ;
  assign n4190 = ~n4187 & ~n4189 ;
  assign n4196 = \DataWidth_reg[1]/NET0131  & ~n4142 ;
  assign n4197 = ~n4190 & ~n4196 ;
  assign n4198 = ~n4195 & ~n4197 ;
  assign n4199 = n952 & ~n4198 ;
  assign n4200 = ~n733 & n4185 ;
  assign n4201 = ~n4188 & ~n4200 ;
  assign n4202 = n993 & ~n4201 ;
  assign n4191 = n970 & ~n4190 ;
  assign n4203 = \InstQueue_reg[6][4]/NET0131  & ~n3933 ;
  assign n4204 = ~n4191 & ~n4203 ;
  assign n4205 = ~n4202 & n4204 ;
  assign n4206 = ~n4199 & n4205 ;
  assign n4213 = n3907 & n4141 ;
  assign n4214 = n3916 & n4163 ;
  assign n4215 = ~n4213 & ~n4214 ;
  assign n4216 = \DataWidth_reg[1]/NET0131  & ~n4215 ;
  assign n4207 = ~n3948 & ~n4185 ;
  assign n4208 = \Datai[4]_pad  & ~n4207 ;
  assign n4209 = \InstQueue_reg[7][4]/NET0131  & ~n3948 ;
  assign n4210 = ~n4185 & n4209 ;
  assign n4211 = ~n4208 & ~n4210 ;
  assign n4217 = \DataWidth_reg[1]/NET0131  & ~n4164 ;
  assign n4218 = ~n4211 & ~n4217 ;
  assign n4219 = ~n4216 & ~n4218 ;
  assign n4220 = n952 & ~n4219 ;
  assign n4221 = ~n733 & n3948 ;
  assign n4222 = ~n4209 & ~n4221 ;
  assign n4223 = n993 & ~n4222 ;
  assign n4212 = n970 & ~n4211 ;
  assign n4224 = \InstQueue_reg[7][4]/NET0131  & ~n3933 ;
  assign n4225 = ~n4212 & ~n4224 ;
  assign n4226 = ~n4223 & n4225 ;
  assign n4227 = ~n4220 & n4226 ;
  assign n4233 = n3907 & n4163 ;
  assign n4234 = n3916 & n4185 ;
  assign n4235 = ~n4233 & ~n4234 ;
  assign n4236 = \DataWidth_reg[1]/NET0131  & ~n4235 ;
  assign n4228 = \Datai[4]_pad  & ~n3954 ;
  assign n4229 = \InstQueue_reg[8][4]/NET0131  & ~n3950 ;
  assign n4230 = ~n3948 & n4229 ;
  assign n4231 = ~n4228 & ~n4230 ;
  assign n4237 = \DataWidth_reg[1]/NET0131  & ~n4186 ;
  assign n4238 = ~n4231 & ~n4237 ;
  assign n4239 = ~n4236 & ~n4238 ;
  assign n4240 = n952 & ~n4239 ;
  assign n4241 = ~n733 & n3950 ;
  assign n4242 = ~n4229 & ~n4241 ;
  assign n4243 = n993 & ~n4242 ;
  assign n4232 = n970 & ~n4231 ;
  assign n4244 = \InstQueue_reg[8][4]/NET0131  & ~n3933 ;
  assign n4245 = ~n4232 & ~n4244 ;
  assign n4246 = ~n4243 & n4245 ;
  assign n4247 = ~n4240 & n4246 ;
  assign n4253 = n3907 & n4185 ;
  assign n4254 = n3916 & n3948 ;
  assign n4255 = ~n4253 & ~n4254 ;
  assign n4256 = \DataWidth_reg[1]/NET0131  & ~n4255 ;
  assign n4248 = \Datai[4]_pad  & ~n3978 ;
  assign n4249 = \InstQueue_reg[9][4]/NET0131  & ~n3941 ;
  assign n4250 = ~n3950 & n4249 ;
  assign n4251 = ~n4248 & ~n4250 ;
  assign n4257 = \DataWidth_reg[1]/NET0131  & ~n4207 ;
  assign n4258 = ~n4251 & ~n4257 ;
  assign n4259 = ~n4256 & ~n4258 ;
  assign n4260 = n952 & ~n4259 ;
  assign n4261 = ~n733 & n3941 ;
  assign n4262 = ~n4249 & ~n4261 ;
  assign n4263 = n993 & ~n4262 ;
  assign n4252 = n970 & ~n4251 ;
  assign n4264 = \InstQueue_reg[9][4]/NET0131  & ~n3933 ;
  assign n4265 = ~n4252 & ~n4264 ;
  assign n4266 = ~n4263 & n4265 ;
  assign n4267 = ~n4260 & n4266 ;
  assign n4271 = \PhyAddrPointer_reg[2]/NET0131  & ~n3496 ;
  assign n4272 = n3540 & ~n4271 ;
  assign n4273 = n948 & ~n4272 ;
  assign n4274 = \PhyAddrPointer_reg[2]/NET0131  & ~n2794 ;
  assign n4268 = ~\PhyAddrPointer_reg[1]/NET0131  & ~\PhyAddrPointer_reg[2]/NET0131  ;
  assign n4269 = ~n3506 & ~n4268 ;
  assign n4270 = n2039 & n4269 ;
  assign n4275 = ~\PhyAddrPointer_reg[2]/NET0131  & n971 ;
  assign n4276 = ~n3516 & ~n4275 ;
  assign n4277 = ~n4270 & n4276 ;
  assign n4278 = ~n4274 & n4277 ;
  assign n4279 = ~n4273 & n4278 ;
  assign n4281 = ~\EAX_reg[20]/NET0131  & ~n3605 ;
  assign n4282 = \EAX_reg[20]/NET0131  & n3605 ;
  assign n4283 = ~n4281 & ~n4282 ;
  assign n4284 = n3798 & n4283 ;
  assign n4285 = ~n833 & n4284 ;
  assign n4286 = ~n828 & n895 ;
  assign n4287 = \Datao[20]_pad  & ~n4286 ;
  assign n4288 = ~n4285 & ~n4287 ;
  assign n4289 = n948 & ~n4288 ;
  assign n4280 = \uWord_reg[4]/NET0131  & n956 ;
  assign n4290 = \Datao[20]_pad  & ~n3816 ;
  assign n4291 = ~n4280 & ~n4290 ;
  assign n4292 = ~n4289 & n4291 ;
  assign n4293 = \uWord_reg[4]/NET0131  & ~n3841 ;
  assign n4294 = \Datai[4]_pad  & n736 ;
  assign n4295 = n826 & n4294 ;
  assign n4296 = ~n4284 & ~n4295 ;
  assign n4297 = n948 & ~n4296 ;
  assign n4298 = ~n4293 & ~n4297 ;
  assign n4299 = \EAX_reg[25]/NET0131  & ~n3116 ;
  assign n4304 = \EAX_reg[23]/NET0131  & n3140 ;
  assign n4305 = \EAX_reg[24]/NET0131  & n4304 ;
  assign n4306 = ~\EAX_reg[25]/NET0131  & ~n4305 ;
  assign n4307 = n3118 & ~n3565 ;
  assign n4308 = ~n4306 & n4307 ;
  assign n4309 = \EAX_reg[25]/NET0131  & ~n3447 ;
  assign n4300 = ~n3248 & n3279 ;
  assign n4301 = n808 & ~n3280 ;
  assign n4302 = ~n4300 & n4301 ;
  assign n4303 = n755 & n4302 ;
  assign n4310 = \Datai[25]_pad  & n835 ;
  assign n4311 = \Datai[9]_pad  & n736 ;
  assign n4312 = ~n4310 & ~n4311 ;
  assign n4313 = n826 & ~n4312 ;
  assign n4314 = ~n4303 & ~n4313 ;
  assign n4315 = ~n4309 & n4314 ;
  assign n4316 = ~n4308 & n4315 ;
  assign n4317 = n948 & ~n4316 ;
  assign n4318 = ~n4299 & ~n4317 ;
  assign n4324 = \Datai[29]_pad  & n3905 ;
  assign n4325 = \Datai[30]_pad  & n4324 ;
  assign n4326 = \Datai[31]_pad  & ~n4325 ;
  assign n4327 = n3876 & n4326 ;
  assign n4328 = \Datai[21]_pad  & n3915 ;
  assign n4329 = \Datai[22]_pad  & n4328 ;
  assign n4330 = ~\Datai[23]_pad  & ~n4329 ;
  assign n4331 = \Datai[23]_pad  & n4329 ;
  assign n4332 = ~n4330 & ~n4331 ;
  assign n4333 = n3919 & n4332 ;
  assign n4334 = ~n4327 & ~n4333 ;
  assign n4335 = \DataWidth_reg[1]/NET0131  & ~n4334 ;
  assign n4319 = \Datai[7]_pad  & ~n3868 ;
  assign n4320 = \InstQueue_reg[0][7]/NET0131  & ~n3864 ;
  assign n4321 = ~n3867 & n4320 ;
  assign n4322 = ~n4319 & ~n4321 ;
  assign n4336 = ~n3924 & ~n4322 ;
  assign n4337 = ~n4335 & ~n4336 ;
  assign n4338 = n952 & ~n4337 ;
  assign n4339 = ~n506 & n3864 ;
  assign n4340 = ~n4320 & ~n4339 ;
  assign n4341 = n993 & ~n4340 ;
  assign n4323 = n970 & ~n4322 ;
  assign n4342 = \InstQueue_reg[0][7]/NET0131  & ~n3933 ;
  assign n4343 = ~n4323 & ~n4342 ;
  assign n4344 = ~n4341 & n4343 ;
  assign n4345 = ~n4338 & n4344 ;
  assign n4351 = n3948 & n4326 ;
  assign n4352 = n3950 & n4332 ;
  assign n4353 = ~n4351 & ~n4352 ;
  assign n4354 = \DataWidth_reg[1]/NET0131  & ~n4353 ;
  assign n4346 = \Datai[7]_pad  & ~n3942 ;
  assign n4347 = \InstQueue_reg[10][7]/NET0131  & ~n3939 ;
  assign n4348 = ~n3941 & n4347 ;
  assign n4349 = ~n4346 & ~n4348 ;
  assign n4355 = ~n3955 & ~n4349 ;
  assign n4356 = ~n4354 & ~n4355 ;
  assign n4357 = n952 & ~n4356 ;
  assign n4358 = ~n506 & n3939 ;
  assign n4359 = ~n4347 & ~n4358 ;
  assign n4360 = n993 & ~n4359 ;
  assign n4350 = n970 & ~n4349 ;
  assign n4361 = \InstQueue_reg[10][7]/NET0131  & ~n3933 ;
  assign n4362 = ~n4350 & ~n4361 ;
  assign n4363 = ~n4360 & n4362 ;
  assign n4364 = ~n4357 & n4363 ;
  assign n4370 = n3950 & n4326 ;
  assign n4371 = n3941 & n4332 ;
  assign n4372 = ~n4370 & ~n4371 ;
  assign n4373 = \DataWidth_reg[1]/NET0131  & ~n4372 ;
  assign n4365 = \Datai[7]_pad  & ~n3968 ;
  assign n4366 = \InstQueue_reg[11][7]/NET0131  & ~n3967 ;
  assign n4367 = ~n3939 & n4366 ;
  assign n4368 = ~n4365 & ~n4367 ;
  assign n4374 = ~n3979 & ~n4368 ;
  assign n4375 = ~n4373 & ~n4374 ;
  assign n4376 = n952 & ~n4375 ;
  assign n4377 = ~n506 & n3967 ;
  assign n4378 = ~n4366 & ~n4377 ;
  assign n4379 = n993 & ~n4378 ;
  assign n4369 = n970 & ~n4368 ;
  assign n4380 = \InstQueue_reg[11][7]/NET0131  & ~n3933 ;
  assign n4381 = ~n4369 & ~n4380 ;
  assign n4382 = ~n4379 & n4381 ;
  assign n4383 = ~n4376 & n4382 ;
  assign n4389 = n3941 & n4326 ;
  assign n4390 = n3939 & n4332 ;
  assign n4391 = ~n4389 & ~n4390 ;
  assign n4392 = \DataWidth_reg[1]/NET0131  & ~n4391 ;
  assign n4384 = \Datai[7]_pad  & ~n3992 ;
  assign n4385 = \InstQueue_reg[12][7]/NET0131  & ~n3991 ;
  assign n4386 = ~n3967 & n4385 ;
  assign n4387 = ~n4384 & ~n4386 ;
  assign n4393 = ~n4002 & ~n4387 ;
  assign n4394 = ~n4392 & ~n4393 ;
  assign n4395 = n952 & ~n4394 ;
  assign n4396 = ~n506 & n3991 ;
  assign n4397 = ~n4385 & ~n4396 ;
  assign n4398 = n993 & ~n4397 ;
  assign n4388 = n970 & ~n4387 ;
  assign n4399 = \InstQueue_reg[12][7]/NET0131  & ~n3933 ;
  assign n4400 = ~n4388 & ~n4399 ;
  assign n4401 = ~n4398 & n4400 ;
  assign n4402 = ~n4395 & n4401 ;
  assign n4408 = n3939 & n4326 ;
  assign n4409 = n3967 & n4332 ;
  assign n4410 = ~n4408 & ~n4409 ;
  assign n4411 = \DataWidth_reg[1]/NET0131  & ~n4410 ;
  assign n4403 = \Datai[7]_pad  & ~n4013 ;
  assign n4404 = \InstQueue_reg[13][7]/NET0131  & ~n3876 ;
  assign n4405 = ~n3991 & n4404 ;
  assign n4406 = ~n4403 & ~n4405 ;
  assign n4412 = ~n4023 & ~n4406 ;
  assign n4413 = ~n4411 & ~n4412 ;
  assign n4414 = n952 & ~n4413 ;
  assign n4415 = ~n506 & n3876 ;
  assign n4416 = ~n4404 & ~n4415 ;
  assign n4417 = n993 & ~n4416 ;
  assign n4407 = n970 & ~n4406 ;
  assign n4418 = \InstQueue_reg[13][7]/NET0131  & ~n3933 ;
  assign n4419 = ~n4407 & ~n4418 ;
  assign n4420 = ~n4417 & n4419 ;
  assign n4421 = ~n4414 & n4420 ;
  assign n4427 = n3967 & n4326 ;
  assign n4428 = n3991 & n4332 ;
  assign n4429 = ~n4427 & ~n4428 ;
  assign n4430 = \DataWidth_reg[1]/NET0131  & ~n4429 ;
  assign n4422 = \Datai[7]_pad  & ~n3923 ;
  assign n4423 = \InstQueue_reg[14][7]/NET0131  & ~n3919 ;
  assign n4424 = ~n3876 & n4423 ;
  assign n4425 = ~n4422 & ~n4424 ;
  assign n4431 = ~n4043 & ~n4425 ;
  assign n4432 = ~n4430 & ~n4431 ;
  assign n4433 = n952 & ~n4432 ;
  assign n4434 = ~n506 & n3919 ;
  assign n4435 = ~n4423 & ~n4434 ;
  assign n4436 = n993 & ~n4435 ;
  assign n4426 = n970 & ~n4425 ;
  assign n4437 = \InstQueue_reg[14][7]/NET0131  & ~n3933 ;
  assign n4438 = ~n4426 & ~n4437 ;
  assign n4439 = ~n4436 & n4438 ;
  assign n4440 = ~n4433 & n4439 ;
  assign n4446 = n3991 & n4326 ;
  assign n4447 = n3876 & n4332 ;
  assign n4448 = ~n4446 & ~n4447 ;
  assign n4449 = \DataWidth_reg[1]/NET0131  & ~n4448 ;
  assign n4441 = \Datai[7]_pad  & ~n4054 ;
  assign n4442 = \InstQueue_reg[15][7]/NET0131  & ~n3867 ;
  assign n4443 = ~n3919 & n4442 ;
  assign n4444 = ~n4441 & ~n4443 ;
  assign n4450 = ~n4064 & ~n4444 ;
  assign n4451 = ~n4449 & ~n4450 ;
  assign n4452 = n952 & ~n4451 ;
  assign n4453 = ~n506 & n3867 ;
  assign n4454 = ~n4442 & ~n4453 ;
  assign n4455 = n993 & ~n4454 ;
  assign n4445 = n970 & ~n4444 ;
  assign n4456 = \InstQueue_reg[15][7]/NET0131  & ~n3933 ;
  assign n4457 = ~n4445 & ~n4456 ;
  assign n4458 = ~n4455 & n4457 ;
  assign n4459 = ~n4452 & n4458 ;
  assign n4465 = n3919 & n4326 ;
  assign n4466 = n3867 & n4332 ;
  assign n4467 = ~n4465 & ~n4466 ;
  assign n4468 = \DataWidth_reg[1]/NET0131  & ~n4467 ;
  assign n4460 = \Datai[7]_pad  & ~n4076 ;
  assign n4461 = \InstQueue_reg[1][7]/NET0131  & ~n4075 ;
  assign n4462 = ~n3864 & n4461 ;
  assign n4463 = ~n4460 & ~n4462 ;
  assign n4469 = ~n4086 & ~n4463 ;
  assign n4470 = ~n4468 & ~n4469 ;
  assign n4471 = n952 & ~n4470 ;
  assign n4472 = ~n506 & n4075 ;
  assign n4473 = ~n4461 & ~n4472 ;
  assign n4474 = n993 & ~n4473 ;
  assign n4464 = n970 & ~n4463 ;
  assign n4475 = \InstQueue_reg[1][7]/NET0131  & ~n3933 ;
  assign n4476 = ~n4464 & ~n4475 ;
  assign n4477 = ~n4474 & n4476 ;
  assign n4478 = ~n4471 & n4477 ;
  assign n4484 = n3864 & n4332 ;
  assign n4485 = n3867 & n4326 ;
  assign n4486 = ~n4484 & ~n4485 ;
  assign n4487 = \DataWidth_reg[1]/NET0131  & ~n4486 ;
  assign n4479 = \Datai[7]_pad  & ~n4098 ;
  assign n4480 = \InstQueue_reg[2][7]/NET0131  & ~n4097 ;
  assign n4481 = ~n4075 & n4480 ;
  assign n4482 = ~n4479 & ~n4481 ;
  assign n4488 = ~n4108 & ~n4482 ;
  assign n4489 = ~n4487 & ~n4488 ;
  assign n4490 = n952 & ~n4489 ;
  assign n4491 = ~n506 & n4097 ;
  assign n4492 = ~n4480 & ~n4491 ;
  assign n4493 = n993 & ~n4492 ;
  assign n4483 = n970 & ~n4482 ;
  assign n4494 = \InstQueue_reg[2][7]/NET0131  & ~n3933 ;
  assign n4495 = ~n4483 & ~n4494 ;
  assign n4496 = ~n4493 & n4495 ;
  assign n4497 = ~n4490 & n4496 ;
  assign n4503 = n3864 & n4326 ;
  assign n4504 = n4075 & n4332 ;
  assign n4505 = ~n4503 & ~n4504 ;
  assign n4506 = \DataWidth_reg[1]/NET0131  & ~n4505 ;
  assign n4498 = \Datai[7]_pad  & ~n4120 ;
  assign n4499 = \InstQueue_reg[3][7]/NET0131  & ~n4119 ;
  assign n4500 = ~n4097 & n4499 ;
  assign n4501 = ~n4498 & ~n4500 ;
  assign n4507 = ~n4130 & ~n4501 ;
  assign n4508 = ~n4506 & ~n4507 ;
  assign n4509 = n952 & ~n4508 ;
  assign n4510 = ~n506 & n4119 ;
  assign n4511 = ~n4499 & ~n4510 ;
  assign n4512 = n993 & ~n4511 ;
  assign n4502 = n970 & ~n4501 ;
  assign n4513 = \InstQueue_reg[3][7]/NET0131  & ~n3933 ;
  assign n4514 = ~n4502 & ~n4513 ;
  assign n4515 = ~n4512 & n4514 ;
  assign n4516 = ~n4509 & n4515 ;
  assign n4522 = n4075 & n4326 ;
  assign n4523 = n4097 & n4332 ;
  assign n4524 = ~n4522 & ~n4523 ;
  assign n4525 = \DataWidth_reg[1]/NET0131  & ~n4524 ;
  assign n4517 = \Datai[7]_pad  & ~n4142 ;
  assign n4518 = \InstQueue_reg[4][7]/NET0131  & ~n4141 ;
  assign n4519 = ~n4119 & n4518 ;
  assign n4520 = ~n4517 & ~n4519 ;
  assign n4526 = ~n4152 & ~n4520 ;
  assign n4527 = ~n4525 & ~n4526 ;
  assign n4528 = n952 & ~n4527 ;
  assign n4529 = ~n506 & n4141 ;
  assign n4530 = ~n4518 & ~n4529 ;
  assign n4531 = n993 & ~n4530 ;
  assign n4521 = n970 & ~n4520 ;
  assign n4532 = \InstQueue_reg[4][7]/NET0131  & ~n3933 ;
  assign n4533 = ~n4521 & ~n4532 ;
  assign n4534 = ~n4531 & n4533 ;
  assign n4535 = ~n4528 & n4534 ;
  assign n4541 = n4097 & n4326 ;
  assign n4542 = n4119 & n4332 ;
  assign n4543 = ~n4541 & ~n4542 ;
  assign n4544 = \DataWidth_reg[1]/NET0131  & ~n4543 ;
  assign n4536 = \Datai[7]_pad  & ~n4164 ;
  assign n4537 = \InstQueue_reg[5][7]/NET0131  & ~n4163 ;
  assign n4538 = ~n4141 & n4537 ;
  assign n4539 = ~n4536 & ~n4538 ;
  assign n4545 = ~n4174 & ~n4539 ;
  assign n4546 = ~n4544 & ~n4545 ;
  assign n4547 = n952 & ~n4546 ;
  assign n4548 = ~n506 & n4163 ;
  assign n4549 = ~n4537 & ~n4548 ;
  assign n4550 = n993 & ~n4549 ;
  assign n4540 = n970 & ~n4539 ;
  assign n4551 = \InstQueue_reg[5][7]/NET0131  & ~n3933 ;
  assign n4552 = ~n4540 & ~n4551 ;
  assign n4553 = ~n4550 & n4552 ;
  assign n4554 = ~n4547 & n4553 ;
  assign n4560 = n4119 & n4326 ;
  assign n4561 = n4141 & n4332 ;
  assign n4562 = ~n4560 & ~n4561 ;
  assign n4563 = \DataWidth_reg[1]/NET0131  & ~n4562 ;
  assign n4555 = \Datai[7]_pad  & ~n4186 ;
  assign n4556 = \InstQueue_reg[6][7]/NET0131  & ~n4185 ;
  assign n4557 = ~n4163 & n4556 ;
  assign n4558 = ~n4555 & ~n4557 ;
  assign n4564 = ~n4196 & ~n4558 ;
  assign n4565 = ~n4563 & ~n4564 ;
  assign n4566 = n952 & ~n4565 ;
  assign n4567 = ~n506 & n4185 ;
  assign n4568 = ~n4556 & ~n4567 ;
  assign n4569 = n993 & ~n4568 ;
  assign n4559 = n970 & ~n4558 ;
  assign n4570 = \InstQueue_reg[6][7]/NET0131  & ~n3933 ;
  assign n4571 = ~n4559 & ~n4570 ;
  assign n4572 = ~n4569 & n4571 ;
  assign n4573 = ~n4566 & n4572 ;
  assign n4579 = n4141 & n4326 ;
  assign n4580 = n4163 & n4332 ;
  assign n4581 = ~n4579 & ~n4580 ;
  assign n4582 = \DataWidth_reg[1]/NET0131  & ~n4581 ;
  assign n4574 = \Datai[7]_pad  & ~n4207 ;
  assign n4575 = \InstQueue_reg[7][7]/NET0131  & ~n3948 ;
  assign n4576 = ~n4185 & n4575 ;
  assign n4577 = ~n4574 & ~n4576 ;
  assign n4583 = ~n4217 & ~n4577 ;
  assign n4584 = ~n4582 & ~n4583 ;
  assign n4585 = n952 & ~n4584 ;
  assign n4586 = ~n506 & n3948 ;
  assign n4587 = ~n4575 & ~n4586 ;
  assign n4588 = n993 & ~n4587 ;
  assign n4578 = n970 & ~n4577 ;
  assign n4589 = \InstQueue_reg[7][7]/NET0131  & ~n3933 ;
  assign n4590 = ~n4578 & ~n4589 ;
  assign n4591 = ~n4588 & n4590 ;
  assign n4592 = ~n4585 & n4591 ;
  assign n4598 = n4163 & n4326 ;
  assign n4599 = n4185 & n4332 ;
  assign n4600 = ~n4598 & ~n4599 ;
  assign n4601 = \DataWidth_reg[1]/NET0131  & ~n4600 ;
  assign n4593 = \Datai[7]_pad  & ~n3954 ;
  assign n4594 = \InstQueue_reg[8][7]/NET0131  & ~n3950 ;
  assign n4595 = ~n3948 & n4594 ;
  assign n4596 = ~n4593 & ~n4595 ;
  assign n4602 = ~n4237 & ~n4596 ;
  assign n4603 = ~n4601 & ~n4602 ;
  assign n4604 = n952 & ~n4603 ;
  assign n4605 = ~n506 & n3950 ;
  assign n4606 = ~n4594 & ~n4605 ;
  assign n4607 = n993 & ~n4606 ;
  assign n4597 = n970 & ~n4596 ;
  assign n4608 = \InstQueue_reg[8][7]/NET0131  & ~n3933 ;
  assign n4609 = ~n4597 & ~n4608 ;
  assign n4610 = ~n4607 & n4609 ;
  assign n4611 = ~n4604 & n4610 ;
  assign n4617 = n4185 & n4326 ;
  assign n4618 = n3948 & n4332 ;
  assign n4619 = ~n4617 & ~n4618 ;
  assign n4620 = \DataWidth_reg[1]/NET0131  & ~n4619 ;
  assign n4612 = \Datai[7]_pad  & ~n3978 ;
  assign n4613 = \InstQueue_reg[9][7]/NET0131  & ~n3941 ;
  assign n4614 = ~n3950 & n4613 ;
  assign n4615 = ~n4612 & ~n4614 ;
  assign n4621 = ~n4257 & ~n4615 ;
  assign n4622 = ~n4620 & ~n4621 ;
  assign n4623 = n952 & ~n4622 ;
  assign n4624 = ~n506 & n3941 ;
  assign n4625 = ~n4613 & ~n4624 ;
  assign n4626 = n993 & ~n4625 ;
  assign n4616 = n970 & ~n4615 ;
  assign n4627 = \InstQueue_reg[9][7]/NET0131  & ~n3933 ;
  assign n4628 = ~n4616 & ~n4627 ;
  assign n4629 = ~n4626 & n4628 ;
  assign n4630 = ~n4623 & n4629 ;
  assign n4652 = \rEIP_reg[22]/NET0131  & \rEIP_reg[23]/NET0131  ;
  assign n4653 = \rEIP_reg[1]/NET0131  & \rEIP_reg[2]/NET0131  ;
  assign n4654 = \rEIP_reg[3]/NET0131  & n4653 ;
  assign n4655 = \rEIP_reg[4]/NET0131  & n4654 ;
  assign n4656 = \rEIP_reg[5]/NET0131  & n4655 ;
  assign n4657 = \rEIP_reg[6]/NET0131  & n4656 ;
  assign n4658 = \rEIP_reg[7]/NET0131  & n4657 ;
  assign n4659 = \rEIP_reg[8]/NET0131  & n4658 ;
  assign n4660 = \rEIP_reg[9]/NET0131  & n4659 ;
  assign n4661 = \rEIP_reg[10]/NET0131  & n4660 ;
  assign n4662 = \rEIP_reg[11]/NET0131  & n4661 ;
  assign n4663 = \rEIP_reg[12]/NET0131  & n4662 ;
  assign n4664 = \rEIP_reg[13]/NET0131  & n4663 ;
  assign n4665 = \rEIP_reg[14]/NET0131  & n4664 ;
  assign n4666 = \rEIP_reg[15]/NET0131  & n4665 ;
  assign n4667 = \rEIP_reg[16]/NET0131  & n4666 ;
  assign n4668 = \rEIP_reg[17]/NET0131  & \rEIP_reg[18]/NET0131  ;
  assign n4669 = \rEIP_reg[19]/NET0131  & n4668 ;
  assign n4670 = \rEIP_reg[20]/NET0131  & \rEIP_reg[21]/NET0131  ;
  assign n4671 = n4669 & n4670 ;
  assign n4672 = n4667 & n4671 ;
  assign n4673 = n4652 & n4672 ;
  assign n4674 = \rEIP_reg[24]/NET0131  & \rEIP_reg[25]/NET0131  ;
  assign n4675 = \rEIP_reg[26]/NET0131  & n4674 ;
  assign n4676 = n4673 & n4675 ;
  assign n4677 = \rEIP_reg[27]/NET0131  & \rEIP_reg[28]/NET0131  ;
  assign n4678 = \rEIP_reg[29]/NET0131  & n4677 ;
  assign n4679 = \rEIP_reg[30]/NET0131  & n4678 ;
  assign n4680 = n4676 & n4679 ;
  assign n4681 = \rEIP_reg[31]/NET0131  & n4680 ;
  assign n4682 = ~\rEIP_reg[31]/NET0131  & ~n4680 ;
  assign n4683 = ~n4681 & ~n4682 ;
  assign n4684 = ~\DataWidth_reg[1]/NET0131  & ~READY_n_pad ;
  assign n4685 = n4683 & n4684 ;
  assign n4689 = ~\EBX_reg[0]/NET0131  & ~\EBX_reg[1]/NET0131  ;
  assign n4690 = ~\EBX_reg[2]/NET0131  & n4689 ;
  assign n4691 = ~\EBX_reg[3]/NET0131  & n4690 ;
  assign n4692 = ~\EBX_reg[4]/NET0131  & n4691 ;
  assign n4693 = ~\EBX_reg[5]/NET0131  & n4692 ;
  assign n4694 = ~\EBX_reg[6]/NET0131  & n4693 ;
  assign n4695 = ~\EBX_reg[7]/NET0131  & n4694 ;
  assign n4696 = ~\EBX_reg[8]/NET0131  & n4695 ;
  assign n4697 = ~\EBX_reg[9]/NET0131  & n4696 ;
  assign n4698 = ~\EBX_reg[10]/NET0131  & ~\EBX_reg[11]/NET0131  ;
  assign n4699 = ~\EBX_reg[12]/NET0131  & n4698 ;
  assign n4700 = n4697 & n4699 ;
  assign n4701 = ~\EBX_reg[13]/NET0131  & n4700 ;
  assign n4702 = ~\EBX_reg[14]/NET0131  & n4701 ;
  assign n4703 = ~\EBX_reg[15]/NET0131  & n4702 ;
  assign n4704 = ~\EBX_reg[16]/NET0131  & n4703 ;
  assign n4705 = ~\EBX_reg[17]/NET0131  & n4704 ;
  assign n4706 = ~\EBX_reg[18]/NET0131  & n4705 ;
  assign n4707 = ~\EBX_reg[19]/NET0131  & n4706 ;
  assign n4708 = ~\EBX_reg[20]/NET0131  & ~\EBX_reg[21]/NET0131  ;
  assign n4709 = ~\EBX_reg[22]/NET0131  & ~\EBX_reg[23]/NET0131  ;
  assign n4710 = n4708 & n4709 ;
  assign n4711 = n4707 & n4710 ;
  assign n4688 = ~\EBX_reg[24]/NET0131  & ~\EBX_reg[25]/NET0131  ;
  assign n4712 = ~\EBX_reg[26]/NET0131  & n4688 ;
  assign n4713 = n4711 & n4712 ;
  assign n4687 = ~\EBX_reg[29]/NET0131  & ~n4684 ;
  assign n4686 = ~\EBX_reg[27]/NET0131  & ~\EBX_reg[28]/NET0131  ;
  assign n4714 = ~\EBX_reg[30]/NET0131  & \EBX_reg[31]/NET0131  ;
  assign n4715 = n4686 & n4714 ;
  assign n4716 = n4687 & n4715 ;
  assign n4717 = n4713 & n4716 ;
  assign n4718 = ~n4685 & ~n4717 ;
  assign n4719 = n1719 & ~n4718 ;
  assign n4650 = ~n744 & n825 ;
  assign n4651 = \rEIP_reg[31]/NET0131  & ~n4650 ;
  assign n4720 = ~\DataWidth_reg[1]/NET0131  & n861 ;
  assign n4722 = ~n4683 & n4720 ;
  assign n4721 = ~\EBX_reg[31]/NET0131  & ~n4720 ;
  assign n4723 = n3798 & ~n4721 ;
  assign n4724 = ~n4722 & n4723 ;
  assign n4725 = ~n4651 & ~n4724 ;
  assign n4726 = ~n4719 & n4725 ;
  assign n4727 = n948 & ~n4726 ;
  assign n4631 = \DataWidth_reg[1]/NET0131  & \rEIP_reg[31]/NET0131  ;
  assign n4639 = ~n2422 & ~n2441 ;
  assign n4635 = ~n2397 & ~n2683 ;
  assign n4632 = ~\PhyAddrPointer_reg[0]/NET0131  & n2801 ;
  assign n4633 = n2022 & n4632 ;
  assign n4634 = \PhyAddrPointer_reg[22]/NET0131  & n4633 ;
  assign n4636 = ~n2869 & n4634 ;
  assign n4637 = n4635 & n4636 ;
  assign n4638 = ~n2716 & n4637 ;
  assign n4640 = ~n2483 & n4638 ;
  assign n4641 = n4639 & n4640 ;
  assign n4642 = ~\DataWidth_reg[1]/NET0131  & ~n2211 ;
  assign n4643 = n2036 & n4642 ;
  assign n4644 = n4641 & n4643 ;
  assign n4645 = ~n4631 & ~n4644 ;
  assign n4646 = n952 & ~n4645 ;
  assign n4647 = ~n970 & n3664 ;
  assign n4648 = \rEIP_reg[31]/NET0131  & ~n4647 ;
  assign n4649 = \PhyAddrPointer_reg[31]/NET0131  & n981 ;
  assign n4728 = ~n4648 & ~n4649 ;
  assign n4729 = ~n4646 & n4728 ;
  assign n4730 = ~n4727 & n4729 ;
  assign n4732 = ~\EAX_reg[27]/NET0131  & ~n3609 ;
  assign n4733 = ~n3610 & n3798 ;
  assign n4734 = ~n4732 & n4733 ;
  assign n4735 = ~n833 & n4734 ;
  assign n4736 = \Datao[27]_pad  & ~n4286 ;
  assign n4737 = ~n4735 & ~n4736 ;
  assign n4738 = n948 & ~n4737 ;
  assign n4731 = \uWord_reg[11]/NET0131  & n956 ;
  assign n4739 = \Datao[27]_pad  & ~n3816 ;
  assign n4740 = ~n4731 & ~n4739 ;
  assign n4741 = ~n4738 & n4740 ;
  assign n4742 = n948 & ~n3447 ;
  assign n4743 = n3116 & ~n4742 ;
  assign n4744 = \EAX_reg[2]/NET0131  & ~n4743 ;
  assign n4746 = \Datai[2]_pad  & n826 ;
  assign n4747 = ~n836 & n4746 ;
  assign n4745 = ~n1225 & n3153 ;
  assign n4748 = ~\EAX_reg[2]/NET0131  & ~n3119 ;
  assign n4749 = ~n3120 & ~n4748 ;
  assign n4750 = n3118 & n4749 ;
  assign n4751 = ~n4745 & ~n4750 ;
  assign n4752 = ~n4747 & n4751 ;
  assign n4753 = n948 & ~n4752 ;
  assign n4754 = ~n4744 & ~n4753 ;
  assign n4755 = \uWord_reg[11]/NET0131  & ~n3584 ;
  assign n4756 = \uWord_reg[11]/NET0131  & ~n3621 ;
  assign n4757 = \Datai[11]_pad  & n826 ;
  assign n4758 = n736 & n4757 ;
  assign n4759 = ~n4756 & ~n4758 ;
  assign n4760 = ~n4734 & n4759 ;
  assign n4761 = n948 & ~n4760 ;
  assign n4762 = ~n4755 & ~n4761 ;
  assign n4763 = \EAX_reg[3]/NET0131  & ~n4743 ;
  assign n4765 = \Datai[3]_pad  & n826 ;
  assign n4766 = ~n836 & n4765 ;
  assign n4764 = ~n1189 & n3153 ;
  assign n4767 = ~\EAX_reg[3]/NET0131  & ~n3120 ;
  assign n4768 = ~n3121 & ~n4767 ;
  assign n4769 = n3118 & n4768 ;
  assign n4770 = ~n4764 & ~n4769 ;
  assign n4771 = ~n4766 & n4770 ;
  assign n4772 = n948 & ~n4771 ;
  assign n4773 = ~n4763 & ~n4772 ;
  assign n4774 = \EAX_reg[4]/NET0131  & ~n4743 ;
  assign n4776 = \Datai[4]_pad  & n865 ;
  assign n4775 = ~n1156 & n3153 ;
  assign n4777 = ~\EAX_reg[4]/NET0131  & ~n3121 ;
  assign n4778 = ~n3122 & ~n4777 ;
  assign n4779 = n3118 & n4778 ;
  assign n4780 = ~n4775 & ~n4779 ;
  assign n4781 = ~n4776 & n4780 ;
  assign n4782 = n948 & ~n4781 ;
  assign n4783 = ~n4774 & ~n4782 ;
  assign n4784 = \EAX_reg[5]/NET0131  & ~n4743 ;
  assign n4786 = \Datai[5]_pad  & n865 ;
  assign n4785 = ~n1120 & n3153 ;
  assign n4787 = ~\EAX_reg[5]/NET0131  & ~n3122 ;
  assign n4788 = ~n3123 & ~n4787 ;
  assign n4789 = n3118 & n4788 ;
  assign n4790 = ~n4785 & ~n4789 ;
  assign n4791 = ~n4786 & n4790 ;
  assign n4792 = n948 & ~n4791 ;
  assign n4793 = ~n4784 & ~n4792 ;
  assign n4794 = \EAX_reg[6]/NET0131  & ~n4743 ;
  assign n4796 = \Datai[6]_pad  & n865 ;
  assign n4795 = ~n1086 & n3153 ;
  assign n4797 = ~\EAX_reg[6]/NET0131  & ~n3123 ;
  assign n4798 = ~n3124 & ~n4797 ;
  assign n4799 = n3118 & n4798 ;
  assign n4800 = ~n4795 & ~n4799 ;
  assign n4801 = ~n4796 & n4800 ;
  assign n4802 = n948 & ~n4801 ;
  assign n4803 = ~n4794 & ~n4802 ;
  assign n4804 = \EAX_reg[7]/NET0131  & ~n4743 ;
  assign n4806 = \Datai[7]_pad  & n865 ;
  assign n4805 = ~n1051 & n3153 ;
  assign n4807 = ~\EAX_reg[7]/NET0131  & ~n3124 ;
  assign n4808 = ~n3125 & ~n4807 ;
  assign n4809 = n3118 & n4808 ;
  assign n4810 = ~n4805 & ~n4809 ;
  assign n4811 = ~n4806 & n4810 ;
  assign n4812 = n948 & ~n4811 ;
  assign n4813 = ~n4804 & ~n4812 ;
  assign n4814 = \EAX_reg[9]/NET0131  & ~n4743 ;
  assign n4815 = \Datai[9]_pad  & n865 ;
  assign n4820 = \InstQueue_reg[4][1]/NET0131  & n478 ;
  assign n4821 = \InstQueue_reg[7][1]/NET0131  & n484 ;
  assign n4834 = ~n4820 & ~n4821 ;
  assign n4822 = \InstQueue_reg[8][1]/NET0131  & n457 ;
  assign n4823 = \InstQueue_reg[12][1]/NET0131  & n490 ;
  assign n4835 = ~n4822 & ~n4823 ;
  assign n4842 = n4834 & n4835 ;
  assign n4816 = \InstQueue_reg[13][1]/NET0131  & n474 ;
  assign n4817 = \InstQueue_reg[10][1]/NET0131  & n486 ;
  assign n4832 = ~n4816 & ~n4817 ;
  assign n4818 = \InstQueue_reg[9][1]/NET0131  & n482 ;
  assign n4819 = \InstQueue_reg[1][1]/NET0131  & n476 ;
  assign n4833 = ~n4818 & ~n4819 ;
  assign n4843 = n4832 & n4833 ;
  assign n4844 = n4842 & n4843 ;
  assign n4828 = \InstQueue_reg[14][1]/NET0131  & n488 ;
  assign n4829 = \InstQueue_reg[15][1]/NET0131  & n471 ;
  assign n4838 = ~n4828 & ~n4829 ;
  assign n4830 = \InstQueue_reg[5][1]/NET0131  & n480 ;
  assign n4831 = \InstQueue_reg[3][1]/NET0131  & n466 ;
  assign n4839 = ~n4830 & ~n4831 ;
  assign n4840 = n4838 & n4839 ;
  assign n4824 = \InstQueue_reg[11][1]/NET0131  & n469 ;
  assign n4825 = \InstQueue_reg[0][1]/NET0131  & n454 ;
  assign n4836 = ~n4824 & ~n4825 ;
  assign n4826 = \InstQueue_reg[6][1]/NET0131  & n463 ;
  assign n4827 = \InstQueue_reg[2][1]/NET0131  & n461 ;
  assign n4837 = ~n4826 & ~n4827 ;
  assign n4841 = n4836 & n4837 ;
  assign n4845 = n4840 & n4841 ;
  assign n4846 = n4844 & n4845 ;
  assign n4847 = n3153 & ~n4846 ;
  assign n4848 = ~\EAX_reg[9]/NET0131  & ~n3126 ;
  assign n4849 = ~n3127 & ~n4848 ;
  assign n4850 = n3118 & n4849 ;
  assign n4851 = ~n4847 & ~n4850 ;
  assign n4852 = ~n4815 & n4851 ;
  assign n4853 = n948 & ~n4852 ;
  assign n4854 = ~n4814 & ~n4853 ;
  assign n4855 = \EAX_reg[8]/NET0131  & ~n4743 ;
  assign n4856 = \Datai[8]_pad  & n865 ;
  assign n4861 = \InstQueue_reg[14][0]/NET0131  & n488 ;
  assign n4862 = \InstQueue_reg[6][0]/NET0131  & n463 ;
  assign n4875 = ~n4861 & ~n4862 ;
  assign n4863 = \InstQueue_reg[13][0]/NET0131  & n474 ;
  assign n4864 = \InstQueue_reg[2][0]/NET0131  & n461 ;
  assign n4876 = ~n4863 & ~n4864 ;
  assign n4883 = n4875 & n4876 ;
  assign n4857 = \InstQueue_reg[8][0]/NET0131  & n457 ;
  assign n4858 = \InstQueue_reg[10][0]/NET0131  & n486 ;
  assign n4873 = ~n4857 & ~n4858 ;
  assign n4859 = \InstQueue_reg[9][0]/NET0131  & n482 ;
  assign n4860 = \InstQueue_reg[1][0]/NET0131  & n476 ;
  assign n4874 = ~n4859 & ~n4860 ;
  assign n4884 = n4873 & n4874 ;
  assign n4885 = n4883 & n4884 ;
  assign n4869 = \InstQueue_reg[11][0]/NET0131  & n469 ;
  assign n4870 = \InstQueue_reg[15][0]/NET0131  & n471 ;
  assign n4879 = ~n4869 & ~n4870 ;
  assign n4871 = \InstQueue_reg[4][0]/NET0131  & n478 ;
  assign n4872 = \InstQueue_reg[7][0]/NET0131  & n484 ;
  assign n4880 = ~n4871 & ~n4872 ;
  assign n4881 = n4879 & n4880 ;
  assign n4865 = \InstQueue_reg[5][0]/NET0131  & n480 ;
  assign n4866 = \InstQueue_reg[0][0]/NET0131  & n454 ;
  assign n4877 = ~n4865 & ~n4866 ;
  assign n4867 = \InstQueue_reg[3][0]/NET0131  & n466 ;
  assign n4868 = \InstQueue_reg[12][0]/NET0131  & n490 ;
  assign n4878 = ~n4867 & ~n4868 ;
  assign n4882 = n4877 & n4878 ;
  assign n4886 = n4881 & n4882 ;
  assign n4887 = n4885 & n4886 ;
  assign n4888 = n3153 & ~n4887 ;
  assign n4889 = ~\EAX_reg[8]/NET0131  & ~n3125 ;
  assign n4890 = ~n3126 & ~n4889 ;
  assign n4891 = n3118 & n4890 ;
  assign n4892 = ~n4888 & ~n4891 ;
  assign n4893 = ~n4856 & n4892 ;
  assign n4894 = n948 & ~n4893 ;
  assign n4895 = ~n4855 & ~n4894 ;
  assign n4896 = \EAX_reg[11]/NET0131  & ~n4743 ;
  assign n4932 = ~n836 & n4757 ;
  assign n4897 = ~\EAX_reg[11]/NET0131  & ~n3128 ;
  assign n4898 = n3118 & ~n3129 ;
  assign n4899 = ~n4897 & n4898 ;
  assign n4904 = \InstQueue_reg[13][3]/NET0131  & n474 ;
  assign n4905 = \InstQueue_reg[7][3]/NET0131  & n484 ;
  assign n4918 = ~n4904 & ~n4905 ;
  assign n4906 = \InstQueue_reg[10][3]/NET0131  & n486 ;
  assign n4907 = \InstQueue_reg[12][3]/NET0131  & n490 ;
  assign n4919 = ~n4906 & ~n4907 ;
  assign n4926 = n4918 & n4919 ;
  assign n4900 = \InstQueue_reg[3][3]/NET0131  & n466 ;
  assign n4901 = \InstQueue_reg[2][3]/NET0131  & n461 ;
  assign n4916 = ~n4900 & ~n4901 ;
  assign n4902 = \InstQueue_reg[1][3]/NET0131  & n476 ;
  assign n4903 = \InstQueue_reg[9][3]/NET0131  & n482 ;
  assign n4917 = ~n4902 & ~n4903 ;
  assign n4927 = n4916 & n4917 ;
  assign n4928 = n4926 & n4927 ;
  assign n4912 = \InstQueue_reg[4][3]/NET0131  & n478 ;
  assign n4913 = \InstQueue_reg[11][3]/NET0131  & n469 ;
  assign n4922 = ~n4912 & ~n4913 ;
  assign n4914 = \InstQueue_reg[8][3]/NET0131  & n457 ;
  assign n4915 = \InstQueue_reg[6][3]/NET0131  & n463 ;
  assign n4923 = ~n4914 & ~n4915 ;
  assign n4924 = n4922 & n4923 ;
  assign n4908 = \InstQueue_reg[15][3]/NET0131  & n471 ;
  assign n4909 = \InstQueue_reg[0][3]/NET0131  & n454 ;
  assign n4920 = ~n4908 & ~n4909 ;
  assign n4910 = \InstQueue_reg[14][3]/NET0131  & n488 ;
  assign n4911 = \InstQueue_reg[5][3]/NET0131  & n480 ;
  assign n4921 = ~n4910 & ~n4911 ;
  assign n4925 = n4920 & n4921 ;
  assign n4929 = n4924 & n4925 ;
  assign n4930 = n4928 & n4929 ;
  assign n4931 = n3153 & ~n4930 ;
  assign n4933 = ~n4899 & ~n4931 ;
  assign n4934 = ~n4932 & n4933 ;
  assign n4935 = n948 & ~n4934 ;
  assign n4936 = ~n4896 & ~n4935 ;
  assign n4940 = \EBX_reg[25]/NET0131  & n3482 ;
  assign n4939 = ~\EBX_reg[25]/NET0131  & ~n3482 ;
  assign n4941 = n773 & ~n4939 ;
  assign n4942 = ~n4940 & n4941 ;
  assign n4937 = n752 & n4302 ;
  assign n4938 = \EBX_reg[25]/NET0131  & n3486 ;
  assign n4943 = ~n4937 & ~n4938 ;
  assign n4944 = ~n4942 & n4943 ;
  assign n4945 = n948 & ~n4944 ;
  assign n4946 = \EBX_reg[25]/NET0131  & ~n3116 ;
  assign n4947 = ~n4945 & ~n4946 ;
  assign n4948 = \EAX_reg[10]/NET0131  & ~n4743 ;
  assign n4981 = n864 & n3563 ;
  assign n4953 = \InstQueue_reg[4][2]/NET0131  & n478 ;
  assign n4954 = \InstQueue_reg[7][2]/NET0131  & n484 ;
  assign n4967 = ~n4953 & ~n4954 ;
  assign n4955 = \InstQueue_reg[8][2]/NET0131  & n457 ;
  assign n4956 = \InstQueue_reg[12][2]/NET0131  & n490 ;
  assign n4968 = ~n4955 & ~n4956 ;
  assign n4975 = n4967 & n4968 ;
  assign n4949 = \InstQueue_reg[13][2]/NET0131  & n474 ;
  assign n4950 = \InstQueue_reg[10][2]/NET0131  & n486 ;
  assign n4965 = ~n4949 & ~n4950 ;
  assign n4951 = \InstQueue_reg[9][2]/NET0131  & n482 ;
  assign n4952 = \InstQueue_reg[1][2]/NET0131  & n476 ;
  assign n4966 = ~n4951 & ~n4952 ;
  assign n4976 = n4965 & n4966 ;
  assign n4977 = n4975 & n4976 ;
  assign n4961 = \InstQueue_reg[14][2]/NET0131  & n488 ;
  assign n4962 = \InstQueue_reg[15][2]/NET0131  & n471 ;
  assign n4971 = ~n4961 & ~n4962 ;
  assign n4963 = \InstQueue_reg[5][2]/NET0131  & n480 ;
  assign n4964 = \InstQueue_reg[3][2]/NET0131  & n466 ;
  assign n4972 = ~n4963 & ~n4964 ;
  assign n4973 = n4971 & n4972 ;
  assign n4957 = \InstQueue_reg[11][2]/NET0131  & n469 ;
  assign n4958 = \InstQueue_reg[0][2]/NET0131  & n454 ;
  assign n4969 = ~n4957 & ~n4958 ;
  assign n4959 = \InstQueue_reg[6][2]/NET0131  & n463 ;
  assign n4960 = \InstQueue_reg[2][2]/NET0131  & n461 ;
  assign n4970 = ~n4959 & ~n4960 ;
  assign n4974 = n4969 & n4970 ;
  assign n4978 = n4973 & n4974 ;
  assign n4979 = n4977 & n4978 ;
  assign n4980 = n3153 & ~n4979 ;
  assign n4982 = ~\EAX_reg[10]/NET0131  & ~n3127 ;
  assign n4983 = n3118 & ~n3128 ;
  assign n4984 = ~n4982 & n4983 ;
  assign n4985 = ~n4980 & ~n4984 ;
  assign n4986 = ~n4981 & n4985 ;
  assign n4987 = n948 & ~n4986 ;
  assign n4988 = ~n4948 & ~n4987 ;
  assign n4989 = \EAX_reg[12]/NET0131  & ~n3116 ;
  assign n4991 = n3447 & ~n4898 ;
  assign n4992 = \EAX_reg[12]/NET0131  & ~n4991 ;
  assign n4990 = \Datai[12]_pad  & n865 ;
  assign n4993 = n3118 & ~n3130 ;
  assign n4994 = n3129 & n4993 ;
  assign n4999 = \InstQueue_reg[4][4]/NET0131  & n478 ;
  assign n5000 = \InstQueue_reg[7][4]/NET0131  & n484 ;
  assign n5013 = ~n4999 & ~n5000 ;
  assign n5001 = \InstQueue_reg[12][4]/NET0131  & n490 ;
  assign n5002 = \InstQueue_reg[6][4]/NET0131  & n463 ;
  assign n5014 = ~n5001 & ~n5002 ;
  assign n5021 = n5013 & n5014 ;
  assign n4995 = \InstQueue_reg[2][4]/NET0131  & n461 ;
  assign n4996 = \InstQueue_reg[3][4]/NET0131  & n466 ;
  assign n5011 = ~n4995 & ~n4996 ;
  assign n4997 = \InstQueue_reg[10][4]/NET0131  & n486 ;
  assign n4998 = \InstQueue_reg[1][4]/NET0131  & n476 ;
  assign n5012 = ~n4997 & ~n4998 ;
  assign n5022 = n5011 & n5012 ;
  assign n5023 = n5021 & n5022 ;
  assign n5007 = \InstQueue_reg[14][4]/NET0131  & n488 ;
  assign n5008 = \InstQueue_reg[9][4]/NET0131  & n482 ;
  assign n5017 = ~n5007 & ~n5008 ;
  assign n5009 = \InstQueue_reg[15][4]/NET0131  & n471 ;
  assign n5010 = \InstQueue_reg[13][4]/NET0131  & n474 ;
  assign n5018 = ~n5009 & ~n5010 ;
  assign n5019 = n5017 & n5018 ;
  assign n5003 = \InstQueue_reg[11][4]/NET0131  & n469 ;
  assign n5004 = \InstQueue_reg[0][4]/NET0131  & n454 ;
  assign n5015 = ~n5003 & ~n5004 ;
  assign n5005 = \InstQueue_reg[5][4]/NET0131  & n480 ;
  assign n5006 = \InstQueue_reg[8][4]/NET0131  & n457 ;
  assign n5016 = ~n5005 & ~n5006 ;
  assign n5020 = n5015 & n5016 ;
  assign n5024 = n5019 & n5020 ;
  assign n5025 = n5023 & n5024 ;
  assign n5026 = n3153 & ~n5025 ;
  assign n5027 = ~n4994 & ~n5026 ;
  assign n5028 = ~n4990 & n5027 ;
  assign n5029 = ~n4992 & n5028 ;
  assign n5030 = n948 & ~n5029 ;
  assign n5031 = ~n4989 & ~n5030 ;
  assign n5032 = \EAX_reg[13]/NET0131  & ~n3116 ;
  assign n5033 = ~n3445 & ~n4993 ;
  assign n5034 = \EAX_reg[13]/NET0131  & ~n5033 ;
  assign n5069 = \EAX_reg[13]/NET0131  & ~n826 ;
  assign n5070 = ~n3767 & ~n5069 ;
  assign n5071 = ~n836 & ~n5070 ;
  assign n5035 = ~\EAX_reg[13]/NET0131  & n3118 ;
  assign n5036 = n3130 & n5035 ;
  assign n5041 = \InstQueue_reg[4][5]/NET0131  & n478 ;
  assign n5042 = \InstQueue_reg[7][5]/NET0131  & n484 ;
  assign n5055 = ~n5041 & ~n5042 ;
  assign n5043 = \InstQueue_reg[8][5]/NET0131  & n457 ;
  assign n5044 = \InstQueue_reg[12][5]/NET0131  & n490 ;
  assign n5056 = ~n5043 & ~n5044 ;
  assign n5063 = n5055 & n5056 ;
  assign n5037 = \InstQueue_reg[13][5]/NET0131  & n474 ;
  assign n5038 = \InstQueue_reg[10][5]/NET0131  & n486 ;
  assign n5053 = ~n5037 & ~n5038 ;
  assign n5039 = \InstQueue_reg[9][5]/NET0131  & n482 ;
  assign n5040 = \InstQueue_reg[1][5]/NET0131  & n476 ;
  assign n5054 = ~n5039 & ~n5040 ;
  assign n5064 = n5053 & n5054 ;
  assign n5065 = n5063 & n5064 ;
  assign n5049 = \InstQueue_reg[14][5]/NET0131  & n488 ;
  assign n5050 = \InstQueue_reg[15][5]/NET0131  & n471 ;
  assign n5059 = ~n5049 & ~n5050 ;
  assign n5051 = \InstQueue_reg[5][5]/NET0131  & n480 ;
  assign n5052 = \InstQueue_reg[3][5]/NET0131  & n466 ;
  assign n5060 = ~n5051 & ~n5052 ;
  assign n5061 = n5059 & n5060 ;
  assign n5045 = \InstQueue_reg[11][5]/NET0131  & n469 ;
  assign n5046 = \InstQueue_reg[0][5]/NET0131  & n454 ;
  assign n5057 = ~n5045 & ~n5046 ;
  assign n5047 = \InstQueue_reg[6][5]/NET0131  & n463 ;
  assign n5048 = \InstQueue_reg[2][5]/NET0131  & n461 ;
  assign n5058 = ~n5047 & ~n5048 ;
  assign n5062 = n5057 & n5058 ;
  assign n5066 = n5061 & n5062 ;
  assign n5067 = n5065 & n5066 ;
  assign n5068 = n3153 & ~n5067 ;
  assign n5072 = ~n5036 & ~n5068 ;
  assign n5073 = ~n5071 & n5072 ;
  assign n5074 = ~n5034 & n5073 ;
  assign n5075 = n948 & ~n5074 ;
  assign n5076 = ~n5032 & ~n5075 ;
  assign n5077 = \EAX_reg[14]/NET0131  & ~n3116 ;
  assign n5079 = n3118 & ~n3131 ;
  assign n5080 = n3447 & ~n5079 ;
  assign n5081 = \EAX_reg[14]/NET0131  & ~n5080 ;
  assign n5078 = \Datai[14]_pad  & n865 ;
  assign n5086 = \InstQueue_reg[7][6]/NET0131  & n484 ;
  assign n5087 = \InstQueue_reg[6][6]/NET0131  & n463 ;
  assign n5100 = ~n5086 & ~n5087 ;
  assign n5088 = \InstQueue_reg[15][6]/NET0131  & n471 ;
  assign n5089 = \InstQueue_reg[12][6]/NET0131  & n490 ;
  assign n5101 = ~n5088 & ~n5089 ;
  assign n5108 = n5100 & n5101 ;
  assign n5082 = \InstQueue_reg[3][6]/NET0131  & n466 ;
  assign n5083 = \InstQueue_reg[2][6]/NET0131  & n461 ;
  assign n5098 = ~n5082 & ~n5083 ;
  assign n5084 = \InstQueue_reg[1][6]/NET0131  & n476 ;
  assign n5085 = \InstQueue_reg[9][6]/NET0131  & n482 ;
  assign n5099 = ~n5084 & ~n5085 ;
  assign n5109 = n5098 & n5099 ;
  assign n5110 = n5108 & n5109 ;
  assign n5094 = \InstQueue_reg[4][6]/NET0131  & n478 ;
  assign n5095 = \InstQueue_reg[11][6]/NET0131  & n469 ;
  assign n5104 = ~n5094 & ~n5095 ;
  assign n5096 = \InstQueue_reg[8][6]/NET0131  & n457 ;
  assign n5097 = \InstQueue_reg[13][6]/NET0131  & n474 ;
  assign n5105 = ~n5096 & ~n5097 ;
  assign n5106 = n5104 & n5105 ;
  assign n5090 = \InstQueue_reg[10][6]/NET0131  & n486 ;
  assign n5091 = \InstQueue_reg[0][6]/NET0131  & n454 ;
  assign n5102 = ~n5090 & ~n5091 ;
  assign n5092 = \InstQueue_reg[14][6]/NET0131  & n488 ;
  assign n5093 = \InstQueue_reg[5][6]/NET0131  & n480 ;
  assign n5103 = ~n5092 & ~n5093 ;
  assign n5107 = n5102 & n5103 ;
  assign n5111 = n5106 & n5107 ;
  assign n5112 = n5110 & n5111 ;
  assign n5113 = n3153 & ~n5112 ;
  assign n5114 = ~\EAX_reg[14]/NET0131  & n3118 ;
  assign n5115 = n3131 & n5114 ;
  assign n5116 = ~n5113 & ~n5115 ;
  assign n5117 = ~n5078 & n5116 ;
  assign n5118 = ~n5081 & n5117 ;
  assign n5119 = n948 & ~n5118 ;
  assign n5120 = ~n5077 & ~n5119 ;
  assign n5121 = \EAX_reg[15]/NET0131  & ~n3116 ;
  assign n5123 = n3118 & ~n3132 ;
  assign n5124 = n3447 & ~n5123 ;
  assign n5125 = \EAX_reg[15]/NET0131  & ~n5124 ;
  assign n5158 = ~\EAX_reg[15]/NET0131  & n3118 ;
  assign n5159 = n3132 & n5158 ;
  assign n5122 = \Datai[15]_pad  & n865 ;
  assign n5130 = \InstQueue_reg[7][7]/NET0131  & n484 ;
  assign n5131 = \InstQueue_reg[6][7]/NET0131  & n463 ;
  assign n5144 = ~n5130 & ~n5131 ;
  assign n5132 = \InstQueue_reg[15][7]/NET0131  & n471 ;
  assign n5133 = \InstQueue_reg[3][7]/NET0131  & n466 ;
  assign n5145 = ~n5132 & ~n5133 ;
  assign n5152 = n5144 & n5145 ;
  assign n5126 = \InstQueue_reg[8][7]/NET0131  & n457 ;
  assign n5127 = \InstQueue_reg[2][7]/NET0131  & n461 ;
  assign n5142 = ~n5126 & ~n5127 ;
  assign n5128 = \InstQueue_reg[1][7]/NET0131  & n476 ;
  assign n5129 = \InstQueue_reg[9][7]/NET0131  & n482 ;
  assign n5143 = ~n5128 & ~n5129 ;
  assign n5153 = n5142 & n5143 ;
  assign n5154 = n5152 & n5153 ;
  assign n5138 = \InstQueue_reg[4][7]/NET0131  & n478 ;
  assign n5139 = \InstQueue_reg[14][7]/NET0131  & n488 ;
  assign n5148 = ~n5138 & ~n5139 ;
  assign n5140 = \InstQueue_reg[12][7]/NET0131  & n490 ;
  assign n5141 = \InstQueue_reg[13][7]/NET0131  & n474 ;
  assign n5149 = ~n5140 & ~n5141 ;
  assign n5150 = n5148 & n5149 ;
  assign n5134 = \InstQueue_reg[10][7]/NET0131  & n486 ;
  assign n5135 = \InstQueue_reg[0][7]/NET0131  & n454 ;
  assign n5146 = ~n5134 & ~n5135 ;
  assign n5136 = \InstQueue_reg[5][7]/NET0131  & n480 ;
  assign n5137 = \InstQueue_reg[11][7]/NET0131  & n469 ;
  assign n5147 = ~n5136 & ~n5137 ;
  assign n5151 = n5146 & n5147 ;
  assign n5155 = n5150 & n5151 ;
  assign n5156 = n5154 & n5155 ;
  assign n5157 = n3153 & ~n5156 ;
  assign n5160 = ~n5122 & ~n5157 ;
  assign n5161 = ~n5159 & n5160 ;
  assign n5162 = ~n5125 & n5161 ;
  assign n5163 = n948 & ~n5162 ;
  assign n5164 = ~n5121 & ~n5163 ;
  assign n5165 = \EAX_reg[1]/NET0131  & ~n4743 ;
  assign n5167 = \Datai[1]_pad  & n826 ;
  assign n5168 = ~n836 & n5167 ;
  assign n5166 = ~n1261 & n3153 ;
  assign n5169 = ~\EAX_reg[0]/NET0131  & ~\EAX_reg[1]/NET0131  ;
  assign n5170 = ~n3119 & ~n5169 ;
  assign n5171 = n3118 & n5170 ;
  assign n5172 = ~n5166 & ~n5171 ;
  assign n5173 = ~n5168 & n5172 ;
  assign n5174 = n948 & ~n5173 ;
  assign n5175 = ~n5165 & ~n5174 ;
  assign n5181 = ~\Datai[27]_pad  & ~n3903 ;
  assign n5182 = ~n3904 & ~n5181 ;
  assign n5183 = n3876 & n5182 ;
  assign n5184 = ~\Datai[19]_pad  & ~n3912 ;
  assign n5185 = ~n3913 & ~n5184 ;
  assign n5186 = n3919 & n5185 ;
  assign n5187 = ~n5183 & ~n5186 ;
  assign n5188 = \DataWidth_reg[1]/NET0131  & ~n5187 ;
  assign n5176 = \Datai[3]_pad  & ~n3868 ;
  assign n5177 = \InstQueue_reg[0][3]/NET0131  & ~n3864 ;
  assign n5178 = ~n3867 & n5177 ;
  assign n5179 = ~n5176 & ~n5178 ;
  assign n5189 = ~n3924 & ~n5179 ;
  assign n5190 = ~n5188 & ~n5189 ;
  assign n5191 = n952 & ~n5190 ;
  assign n5192 = ~n632 & n3864 ;
  assign n5193 = ~n5177 & ~n5192 ;
  assign n5194 = n993 & ~n5193 ;
  assign n5180 = n970 & ~n5179 ;
  assign n5195 = \InstQueue_reg[0][3]/NET0131  & ~n3933 ;
  assign n5196 = ~n5180 & ~n5195 ;
  assign n5197 = ~n5194 & n5196 ;
  assign n5198 = ~n5191 & n5197 ;
  assign n5204 = ~\Datai[30]_pad  & ~n4324 ;
  assign n5205 = ~n4325 & ~n5204 ;
  assign n5206 = n3876 & n5205 ;
  assign n5207 = ~\Datai[22]_pad  & ~n4328 ;
  assign n5208 = ~n4329 & ~n5207 ;
  assign n5209 = n3919 & n5208 ;
  assign n5210 = ~n5206 & ~n5209 ;
  assign n5211 = \DataWidth_reg[1]/NET0131  & ~n5210 ;
  assign n5199 = \Datai[6]_pad  & ~n3868 ;
  assign n5200 = \InstQueue_reg[0][6]/NET0131  & ~n3864 ;
  assign n5201 = ~n3867 & n5200 ;
  assign n5202 = ~n5199 & ~n5201 ;
  assign n5212 = ~n3924 & ~n5202 ;
  assign n5213 = ~n5211 & ~n5212 ;
  assign n5214 = n952 & ~n5213 ;
  assign n5215 = ~n537 & n3864 ;
  assign n5216 = ~n5200 & ~n5215 ;
  assign n5217 = n993 & ~n5216 ;
  assign n5203 = n970 & ~n5202 ;
  assign n5218 = \InstQueue_reg[0][6]/NET0131  & ~n3933 ;
  assign n5219 = ~n5203 & ~n5218 ;
  assign n5220 = ~n5217 & n5219 ;
  assign n5221 = ~n5214 & n5220 ;
  assign n5227 = n3948 & n5182 ;
  assign n5228 = n3950 & n5185 ;
  assign n5229 = ~n5227 & ~n5228 ;
  assign n5230 = \DataWidth_reg[1]/NET0131  & ~n5229 ;
  assign n5222 = \Datai[3]_pad  & ~n3942 ;
  assign n5223 = \InstQueue_reg[10][3]/NET0131  & ~n3939 ;
  assign n5224 = ~n3941 & n5223 ;
  assign n5225 = ~n5222 & ~n5224 ;
  assign n5231 = ~n3955 & ~n5225 ;
  assign n5232 = ~n5230 & ~n5231 ;
  assign n5233 = n952 & ~n5232 ;
  assign n5234 = ~n632 & n3939 ;
  assign n5235 = ~n5223 & ~n5234 ;
  assign n5236 = n993 & ~n5235 ;
  assign n5226 = n970 & ~n5225 ;
  assign n5237 = \InstQueue_reg[10][3]/NET0131  & ~n3933 ;
  assign n5238 = ~n5226 & ~n5237 ;
  assign n5239 = ~n5236 & n5238 ;
  assign n5240 = ~n5233 & n5239 ;
  assign n5246 = n3948 & n5205 ;
  assign n5247 = n3950 & n5208 ;
  assign n5248 = ~n5246 & ~n5247 ;
  assign n5249 = \DataWidth_reg[1]/NET0131  & ~n5248 ;
  assign n5241 = \Datai[6]_pad  & ~n3942 ;
  assign n5242 = \InstQueue_reg[10][6]/NET0131  & ~n3939 ;
  assign n5243 = ~n3941 & n5242 ;
  assign n5244 = ~n5241 & ~n5243 ;
  assign n5250 = ~n3955 & ~n5244 ;
  assign n5251 = ~n5249 & ~n5250 ;
  assign n5252 = n952 & ~n5251 ;
  assign n5253 = ~n537 & n3939 ;
  assign n5254 = ~n5242 & ~n5253 ;
  assign n5255 = n993 & ~n5254 ;
  assign n5245 = n970 & ~n5244 ;
  assign n5256 = \InstQueue_reg[10][6]/NET0131  & ~n3933 ;
  assign n5257 = ~n5245 & ~n5256 ;
  assign n5258 = ~n5255 & n5257 ;
  assign n5259 = ~n5252 & n5258 ;
  assign n5265 = n3950 & n5182 ;
  assign n5266 = n3941 & n5185 ;
  assign n5267 = ~n5265 & ~n5266 ;
  assign n5268 = \DataWidth_reg[1]/NET0131  & ~n5267 ;
  assign n5260 = \Datai[3]_pad  & ~n3968 ;
  assign n5261 = \InstQueue_reg[11][3]/NET0131  & ~n3967 ;
  assign n5262 = ~n3939 & n5261 ;
  assign n5263 = ~n5260 & ~n5262 ;
  assign n5269 = ~n3979 & ~n5263 ;
  assign n5270 = ~n5268 & ~n5269 ;
  assign n5271 = n952 & ~n5270 ;
  assign n5272 = ~n632 & n3967 ;
  assign n5273 = ~n5261 & ~n5272 ;
  assign n5274 = n993 & ~n5273 ;
  assign n5264 = n970 & ~n5263 ;
  assign n5275 = \InstQueue_reg[11][3]/NET0131  & ~n3933 ;
  assign n5276 = ~n5264 & ~n5275 ;
  assign n5277 = ~n5274 & n5276 ;
  assign n5278 = ~n5271 & n5277 ;
  assign n5284 = n3950 & n5205 ;
  assign n5285 = n3941 & n5208 ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = \DataWidth_reg[1]/NET0131  & ~n5286 ;
  assign n5279 = \Datai[6]_pad  & ~n3968 ;
  assign n5280 = \InstQueue_reg[11][6]/NET0131  & ~n3967 ;
  assign n5281 = ~n3939 & n5280 ;
  assign n5282 = ~n5279 & ~n5281 ;
  assign n5288 = ~n3979 & ~n5282 ;
  assign n5289 = ~n5287 & ~n5288 ;
  assign n5290 = n952 & ~n5289 ;
  assign n5291 = ~n537 & n3967 ;
  assign n5292 = ~n5280 & ~n5291 ;
  assign n5293 = n993 & ~n5292 ;
  assign n5283 = n970 & ~n5282 ;
  assign n5294 = \InstQueue_reg[11][6]/NET0131  & ~n3933 ;
  assign n5295 = ~n5283 & ~n5294 ;
  assign n5296 = ~n5293 & n5295 ;
  assign n5297 = ~n5290 & n5296 ;
  assign n5303 = n3941 & n5182 ;
  assign n5304 = n3939 & n5185 ;
  assign n5305 = ~n5303 & ~n5304 ;
  assign n5306 = \DataWidth_reg[1]/NET0131  & ~n5305 ;
  assign n5298 = \Datai[3]_pad  & ~n3992 ;
  assign n5299 = \InstQueue_reg[12][3]/NET0131  & ~n3991 ;
  assign n5300 = ~n3967 & n5299 ;
  assign n5301 = ~n5298 & ~n5300 ;
  assign n5307 = ~n4002 & ~n5301 ;
  assign n5308 = ~n5306 & ~n5307 ;
  assign n5309 = n952 & ~n5308 ;
  assign n5310 = ~n632 & n3991 ;
  assign n5311 = ~n5299 & ~n5310 ;
  assign n5312 = n993 & ~n5311 ;
  assign n5302 = n970 & ~n5301 ;
  assign n5313 = \InstQueue_reg[12][3]/NET0131  & ~n3933 ;
  assign n5314 = ~n5302 & ~n5313 ;
  assign n5315 = ~n5312 & n5314 ;
  assign n5316 = ~n5309 & n5315 ;
  assign n5322 = n3941 & n5205 ;
  assign n5323 = n3939 & n5208 ;
  assign n5324 = ~n5322 & ~n5323 ;
  assign n5325 = \DataWidth_reg[1]/NET0131  & ~n5324 ;
  assign n5317 = \Datai[6]_pad  & ~n3992 ;
  assign n5318 = \InstQueue_reg[12][6]/NET0131  & ~n3991 ;
  assign n5319 = ~n3967 & n5318 ;
  assign n5320 = ~n5317 & ~n5319 ;
  assign n5326 = ~n4002 & ~n5320 ;
  assign n5327 = ~n5325 & ~n5326 ;
  assign n5328 = n952 & ~n5327 ;
  assign n5329 = ~n537 & n3991 ;
  assign n5330 = ~n5318 & ~n5329 ;
  assign n5331 = n993 & ~n5330 ;
  assign n5321 = n970 & ~n5320 ;
  assign n5332 = \InstQueue_reg[12][6]/NET0131  & ~n3933 ;
  assign n5333 = ~n5321 & ~n5332 ;
  assign n5334 = ~n5331 & n5333 ;
  assign n5335 = ~n5328 & n5334 ;
  assign n5341 = n3939 & n5182 ;
  assign n5342 = n3967 & n5185 ;
  assign n5343 = ~n5341 & ~n5342 ;
  assign n5344 = \DataWidth_reg[1]/NET0131  & ~n5343 ;
  assign n5336 = \Datai[3]_pad  & ~n4013 ;
  assign n5337 = \InstQueue_reg[13][3]/NET0131  & ~n3876 ;
  assign n5338 = ~n3991 & n5337 ;
  assign n5339 = ~n5336 & ~n5338 ;
  assign n5345 = ~n4023 & ~n5339 ;
  assign n5346 = ~n5344 & ~n5345 ;
  assign n5347 = n952 & ~n5346 ;
  assign n5348 = ~n632 & n3876 ;
  assign n5349 = ~n5337 & ~n5348 ;
  assign n5350 = n993 & ~n5349 ;
  assign n5340 = n970 & ~n5339 ;
  assign n5351 = \InstQueue_reg[13][3]/NET0131  & ~n3933 ;
  assign n5352 = ~n5340 & ~n5351 ;
  assign n5353 = ~n5350 & n5352 ;
  assign n5354 = ~n5347 & n5353 ;
  assign n5360 = n3939 & n5205 ;
  assign n5361 = n3967 & n5208 ;
  assign n5362 = ~n5360 & ~n5361 ;
  assign n5363 = \DataWidth_reg[1]/NET0131  & ~n5362 ;
  assign n5355 = \Datai[6]_pad  & ~n4013 ;
  assign n5356 = \InstQueue_reg[13][6]/NET0131  & ~n3876 ;
  assign n5357 = ~n3991 & n5356 ;
  assign n5358 = ~n5355 & ~n5357 ;
  assign n5364 = ~n4023 & ~n5358 ;
  assign n5365 = ~n5363 & ~n5364 ;
  assign n5366 = n952 & ~n5365 ;
  assign n5367 = ~n537 & n3876 ;
  assign n5368 = ~n5356 & ~n5367 ;
  assign n5369 = n993 & ~n5368 ;
  assign n5359 = n970 & ~n5358 ;
  assign n5370 = \InstQueue_reg[13][6]/NET0131  & ~n3933 ;
  assign n5371 = ~n5359 & ~n5370 ;
  assign n5372 = ~n5369 & n5371 ;
  assign n5373 = ~n5366 & n5372 ;
  assign n5379 = n3967 & n5182 ;
  assign n5380 = n3991 & n5185 ;
  assign n5381 = ~n5379 & ~n5380 ;
  assign n5382 = \DataWidth_reg[1]/NET0131  & ~n5381 ;
  assign n5374 = \Datai[3]_pad  & ~n3923 ;
  assign n5375 = \InstQueue_reg[14][3]/NET0131  & ~n3919 ;
  assign n5376 = ~n3876 & n5375 ;
  assign n5377 = ~n5374 & ~n5376 ;
  assign n5383 = ~n4043 & ~n5377 ;
  assign n5384 = ~n5382 & ~n5383 ;
  assign n5385 = n952 & ~n5384 ;
  assign n5386 = ~n632 & n3919 ;
  assign n5387 = ~n5375 & ~n5386 ;
  assign n5388 = n993 & ~n5387 ;
  assign n5378 = n970 & ~n5377 ;
  assign n5389 = \InstQueue_reg[14][3]/NET0131  & ~n3933 ;
  assign n5390 = ~n5378 & ~n5389 ;
  assign n5391 = ~n5388 & n5390 ;
  assign n5392 = ~n5385 & n5391 ;
  assign n5398 = n3967 & n5205 ;
  assign n5399 = n3991 & n5208 ;
  assign n5400 = ~n5398 & ~n5399 ;
  assign n5401 = \DataWidth_reg[1]/NET0131  & ~n5400 ;
  assign n5393 = \Datai[6]_pad  & ~n3923 ;
  assign n5394 = \InstQueue_reg[14][6]/NET0131  & ~n3919 ;
  assign n5395 = ~n3876 & n5394 ;
  assign n5396 = ~n5393 & ~n5395 ;
  assign n5402 = ~n4043 & ~n5396 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = n952 & ~n5403 ;
  assign n5405 = ~n537 & n3919 ;
  assign n5406 = ~n5394 & ~n5405 ;
  assign n5407 = n993 & ~n5406 ;
  assign n5397 = n970 & ~n5396 ;
  assign n5408 = \InstQueue_reg[14][6]/NET0131  & ~n3933 ;
  assign n5409 = ~n5397 & ~n5408 ;
  assign n5410 = ~n5407 & n5409 ;
  assign n5411 = ~n5404 & n5410 ;
  assign n5417 = n3991 & n5182 ;
  assign n5418 = n3876 & n5185 ;
  assign n5419 = ~n5417 & ~n5418 ;
  assign n5420 = \DataWidth_reg[1]/NET0131  & ~n5419 ;
  assign n5412 = \Datai[3]_pad  & ~n4054 ;
  assign n5413 = \InstQueue_reg[15][3]/NET0131  & ~n3867 ;
  assign n5414 = ~n3919 & n5413 ;
  assign n5415 = ~n5412 & ~n5414 ;
  assign n5421 = ~n4064 & ~n5415 ;
  assign n5422 = ~n5420 & ~n5421 ;
  assign n5423 = n952 & ~n5422 ;
  assign n5424 = ~n632 & n3867 ;
  assign n5425 = ~n5413 & ~n5424 ;
  assign n5426 = n993 & ~n5425 ;
  assign n5416 = n970 & ~n5415 ;
  assign n5427 = \InstQueue_reg[15][3]/NET0131  & ~n3933 ;
  assign n5428 = ~n5416 & ~n5427 ;
  assign n5429 = ~n5426 & n5428 ;
  assign n5430 = ~n5423 & n5429 ;
  assign n5436 = n3991 & n5205 ;
  assign n5437 = n3876 & n5208 ;
  assign n5438 = ~n5436 & ~n5437 ;
  assign n5439 = \DataWidth_reg[1]/NET0131  & ~n5438 ;
  assign n5431 = \Datai[6]_pad  & ~n4054 ;
  assign n5432 = \InstQueue_reg[15][6]/NET0131  & ~n3867 ;
  assign n5433 = ~n3919 & n5432 ;
  assign n5434 = ~n5431 & ~n5433 ;
  assign n5440 = ~n4064 & ~n5434 ;
  assign n5441 = ~n5439 & ~n5440 ;
  assign n5442 = n952 & ~n5441 ;
  assign n5443 = ~n537 & n3867 ;
  assign n5444 = ~n5432 & ~n5443 ;
  assign n5445 = n993 & ~n5444 ;
  assign n5435 = n970 & ~n5434 ;
  assign n5446 = \InstQueue_reg[15][6]/NET0131  & ~n3933 ;
  assign n5447 = ~n5435 & ~n5446 ;
  assign n5448 = ~n5445 & n5447 ;
  assign n5449 = ~n5442 & n5448 ;
  assign n5455 = n3919 & n5182 ;
  assign n5456 = n3867 & n5185 ;
  assign n5457 = ~n5455 & ~n5456 ;
  assign n5458 = \DataWidth_reg[1]/NET0131  & ~n5457 ;
  assign n5450 = \Datai[3]_pad  & ~n4076 ;
  assign n5451 = \InstQueue_reg[1][3]/NET0131  & ~n4075 ;
  assign n5452 = ~n3864 & n5451 ;
  assign n5453 = ~n5450 & ~n5452 ;
  assign n5459 = ~n4086 & ~n5453 ;
  assign n5460 = ~n5458 & ~n5459 ;
  assign n5461 = n952 & ~n5460 ;
  assign n5462 = ~n632 & n4075 ;
  assign n5463 = ~n5451 & ~n5462 ;
  assign n5464 = n993 & ~n5463 ;
  assign n5454 = n970 & ~n5453 ;
  assign n5465 = \InstQueue_reg[1][3]/NET0131  & ~n3933 ;
  assign n5466 = ~n5454 & ~n5465 ;
  assign n5467 = ~n5464 & n5466 ;
  assign n5468 = ~n5461 & n5467 ;
  assign n5474 = n3919 & n5205 ;
  assign n5475 = n3867 & n5208 ;
  assign n5476 = ~n5474 & ~n5475 ;
  assign n5477 = \DataWidth_reg[1]/NET0131  & ~n5476 ;
  assign n5469 = \Datai[6]_pad  & ~n4076 ;
  assign n5470 = \InstQueue_reg[1][6]/NET0131  & ~n4075 ;
  assign n5471 = ~n3864 & n5470 ;
  assign n5472 = ~n5469 & ~n5471 ;
  assign n5478 = ~n4086 & ~n5472 ;
  assign n5479 = ~n5477 & ~n5478 ;
  assign n5480 = n952 & ~n5479 ;
  assign n5481 = ~n537 & n4075 ;
  assign n5482 = ~n5470 & ~n5481 ;
  assign n5483 = n993 & ~n5482 ;
  assign n5473 = n970 & ~n5472 ;
  assign n5484 = \InstQueue_reg[1][6]/NET0131  & ~n3933 ;
  assign n5485 = ~n5473 & ~n5484 ;
  assign n5486 = ~n5483 & n5485 ;
  assign n5487 = ~n5480 & n5486 ;
  assign n5493 = n3864 & n5185 ;
  assign n5494 = n3867 & n5182 ;
  assign n5495 = ~n5493 & ~n5494 ;
  assign n5496 = \DataWidth_reg[1]/NET0131  & ~n5495 ;
  assign n5488 = \Datai[3]_pad  & ~n4098 ;
  assign n5489 = \InstQueue_reg[2][3]/NET0131  & ~n4097 ;
  assign n5490 = ~n4075 & n5489 ;
  assign n5491 = ~n5488 & ~n5490 ;
  assign n5497 = ~n4108 & ~n5491 ;
  assign n5498 = ~n5496 & ~n5497 ;
  assign n5499 = n952 & ~n5498 ;
  assign n5500 = ~n632 & n4097 ;
  assign n5501 = ~n5489 & ~n5500 ;
  assign n5502 = n993 & ~n5501 ;
  assign n5492 = n970 & ~n5491 ;
  assign n5503 = \InstQueue_reg[2][3]/NET0131  & ~n3933 ;
  assign n5504 = ~n5492 & ~n5503 ;
  assign n5505 = ~n5502 & n5504 ;
  assign n5506 = ~n5499 & n5505 ;
  assign n5512 = n3864 & n5208 ;
  assign n5513 = n3867 & n5205 ;
  assign n5514 = ~n5512 & ~n5513 ;
  assign n5515 = \DataWidth_reg[1]/NET0131  & ~n5514 ;
  assign n5507 = \Datai[6]_pad  & ~n4098 ;
  assign n5508 = \InstQueue_reg[2][6]/NET0131  & ~n4097 ;
  assign n5509 = ~n4075 & n5508 ;
  assign n5510 = ~n5507 & ~n5509 ;
  assign n5516 = ~n4108 & ~n5510 ;
  assign n5517 = ~n5515 & ~n5516 ;
  assign n5518 = n952 & ~n5517 ;
  assign n5519 = ~n537 & n4097 ;
  assign n5520 = ~n5508 & ~n5519 ;
  assign n5521 = n993 & ~n5520 ;
  assign n5511 = n970 & ~n5510 ;
  assign n5522 = \InstQueue_reg[2][6]/NET0131  & ~n3933 ;
  assign n5523 = ~n5511 & ~n5522 ;
  assign n5524 = ~n5521 & n5523 ;
  assign n5525 = ~n5518 & n5524 ;
  assign n5531 = n3864 & n5182 ;
  assign n5532 = n4075 & n5185 ;
  assign n5533 = ~n5531 & ~n5532 ;
  assign n5534 = \DataWidth_reg[1]/NET0131  & ~n5533 ;
  assign n5526 = \Datai[3]_pad  & ~n4120 ;
  assign n5527 = \InstQueue_reg[3][3]/NET0131  & ~n4119 ;
  assign n5528 = ~n4097 & n5527 ;
  assign n5529 = ~n5526 & ~n5528 ;
  assign n5535 = ~n4130 & ~n5529 ;
  assign n5536 = ~n5534 & ~n5535 ;
  assign n5537 = n952 & ~n5536 ;
  assign n5538 = ~n632 & n4119 ;
  assign n5539 = ~n5527 & ~n5538 ;
  assign n5540 = n993 & ~n5539 ;
  assign n5530 = n970 & ~n5529 ;
  assign n5541 = \InstQueue_reg[3][3]/NET0131  & ~n3933 ;
  assign n5542 = ~n5530 & ~n5541 ;
  assign n5543 = ~n5540 & n5542 ;
  assign n5544 = ~n5537 & n5543 ;
  assign n5550 = n3864 & n5205 ;
  assign n5551 = n4075 & n5208 ;
  assign n5552 = ~n5550 & ~n5551 ;
  assign n5553 = \DataWidth_reg[1]/NET0131  & ~n5552 ;
  assign n5545 = \Datai[6]_pad  & ~n4120 ;
  assign n5546 = \InstQueue_reg[3][6]/NET0131  & ~n4119 ;
  assign n5547 = ~n4097 & n5546 ;
  assign n5548 = ~n5545 & ~n5547 ;
  assign n5554 = ~n4130 & ~n5548 ;
  assign n5555 = ~n5553 & ~n5554 ;
  assign n5556 = n952 & ~n5555 ;
  assign n5557 = ~n537 & n4119 ;
  assign n5558 = ~n5546 & ~n5557 ;
  assign n5559 = n993 & ~n5558 ;
  assign n5549 = n970 & ~n5548 ;
  assign n5560 = \InstQueue_reg[3][6]/NET0131  & ~n3933 ;
  assign n5561 = ~n5549 & ~n5560 ;
  assign n5562 = ~n5559 & n5561 ;
  assign n5563 = ~n5556 & n5562 ;
  assign n5569 = n4075 & n5182 ;
  assign n5570 = n4097 & n5185 ;
  assign n5571 = ~n5569 & ~n5570 ;
  assign n5572 = \DataWidth_reg[1]/NET0131  & ~n5571 ;
  assign n5564 = \Datai[3]_pad  & ~n4142 ;
  assign n5565 = \InstQueue_reg[4][3]/NET0131  & ~n4141 ;
  assign n5566 = ~n4119 & n5565 ;
  assign n5567 = ~n5564 & ~n5566 ;
  assign n5573 = ~n4152 & ~n5567 ;
  assign n5574 = ~n5572 & ~n5573 ;
  assign n5575 = n952 & ~n5574 ;
  assign n5576 = ~n632 & n4141 ;
  assign n5577 = ~n5565 & ~n5576 ;
  assign n5578 = n993 & ~n5577 ;
  assign n5568 = n970 & ~n5567 ;
  assign n5579 = \InstQueue_reg[4][3]/NET0131  & ~n3933 ;
  assign n5580 = ~n5568 & ~n5579 ;
  assign n5581 = ~n5578 & n5580 ;
  assign n5582 = ~n5575 & n5581 ;
  assign n5588 = n4075 & n5205 ;
  assign n5589 = n4097 & n5208 ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5591 = \DataWidth_reg[1]/NET0131  & ~n5590 ;
  assign n5583 = \Datai[6]_pad  & ~n4142 ;
  assign n5584 = \InstQueue_reg[4][6]/NET0131  & ~n4141 ;
  assign n5585 = ~n4119 & n5584 ;
  assign n5586 = ~n5583 & ~n5585 ;
  assign n5592 = ~n4152 & ~n5586 ;
  assign n5593 = ~n5591 & ~n5592 ;
  assign n5594 = n952 & ~n5593 ;
  assign n5595 = ~n537 & n4141 ;
  assign n5596 = ~n5584 & ~n5595 ;
  assign n5597 = n993 & ~n5596 ;
  assign n5587 = n970 & ~n5586 ;
  assign n5598 = \InstQueue_reg[4][6]/NET0131  & ~n3933 ;
  assign n5599 = ~n5587 & ~n5598 ;
  assign n5600 = ~n5597 & n5599 ;
  assign n5601 = ~n5594 & n5600 ;
  assign n5607 = n4097 & n5182 ;
  assign n5608 = n4119 & n5185 ;
  assign n5609 = ~n5607 & ~n5608 ;
  assign n5610 = \DataWidth_reg[1]/NET0131  & ~n5609 ;
  assign n5602 = \Datai[3]_pad  & ~n4164 ;
  assign n5603 = \InstQueue_reg[5][3]/NET0131  & ~n4163 ;
  assign n5604 = ~n4141 & n5603 ;
  assign n5605 = ~n5602 & ~n5604 ;
  assign n5611 = ~n4174 & ~n5605 ;
  assign n5612 = ~n5610 & ~n5611 ;
  assign n5613 = n952 & ~n5612 ;
  assign n5614 = ~n632 & n4163 ;
  assign n5615 = ~n5603 & ~n5614 ;
  assign n5616 = n993 & ~n5615 ;
  assign n5606 = n970 & ~n5605 ;
  assign n5617 = \InstQueue_reg[5][3]/NET0131  & ~n3933 ;
  assign n5618 = ~n5606 & ~n5617 ;
  assign n5619 = ~n5616 & n5618 ;
  assign n5620 = ~n5613 & n5619 ;
  assign n5626 = n4097 & n5205 ;
  assign n5627 = n4119 & n5208 ;
  assign n5628 = ~n5626 & ~n5627 ;
  assign n5629 = \DataWidth_reg[1]/NET0131  & ~n5628 ;
  assign n5621 = \Datai[6]_pad  & ~n4164 ;
  assign n5622 = \InstQueue_reg[5][6]/NET0131  & ~n4163 ;
  assign n5623 = ~n4141 & n5622 ;
  assign n5624 = ~n5621 & ~n5623 ;
  assign n5630 = ~n4174 & ~n5624 ;
  assign n5631 = ~n5629 & ~n5630 ;
  assign n5632 = n952 & ~n5631 ;
  assign n5633 = ~n537 & n4163 ;
  assign n5634 = ~n5622 & ~n5633 ;
  assign n5635 = n993 & ~n5634 ;
  assign n5625 = n970 & ~n5624 ;
  assign n5636 = \InstQueue_reg[5][6]/NET0131  & ~n3933 ;
  assign n5637 = ~n5625 & ~n5636 ;
  assign n5638 = ~n5635 & n5637 ;
  assign n5639 = ~n5632 & n5638 ;
  assign n5645 = n4119 & n5182 ;
  assign n5646 = n4141 & n5185 ;
  assign n5647 = ~n5645 & ~n5646 ;
  assign n5648 = \DataWidth_reg[1]/NET0131  & ~n5647 ;
  assign n5640 = \Datai[3]_pad  & ~n4186 ;
  assign n5641 = \InstQueue_reg[6][3]/NET0131  & ~n4185 ;
  assign n5642 = ~n4163 & n5641 ;
  assign n5643 = ~n5640 & ~n5642 ;
  assign n5649 = ~n4196 & ~n5643 ;
  assign n5650 = ~n5648 & ~n5649 ;
  assign n5651 = n952 & ~n5650 ;
  assign n5652 = ~n632 & n4185 ;
  assign n5653 = ~n5641 & ~n5652 ;
  assign n5654 = n993 & ~n5653 ;
  assign n5644 = n970 & ~n5643 ;
  assign n5655 = \InstQueue_reg[6][3]/NET0131  & ~n3933 ;
  assign n5656 = ~n5644 & ~n5655 ;
  assign n5657 = ~n5654 & n5656 ;
  assign n5658 = ~n5651 & n5657 ;
  assign n5664 = n4119 & n5205 ;
  assign n5665 = n4141 & n5208 ;
  assign n5666 = ~n5664 & ~n5665 ;
  assign n5667 = \DataWidth_reg[1]/NET0131  & ~n5666 ;
  assign n5659 = \Datai[6]_pad  & ~n4186 ;
  assign n5660 = \InstQueue_reg[6][6]/NET0131  & ~n4185 ;
  assign n5661 = ~n4163 & n5660 ;
  assign n5662 = ~n5659 & ~n5661 ;
  assign n5668 = ~n4196 & ~n5662 ;
  assign n5669 = ~n5667 & ~n5668 ;
  assign n5670 = n952 & ~n5669 ;
  assign n5671 = ~n537 & n4185 ;
  assign n5672 = ~n5660 & ~n5671 ;
  assign n5673 = n993 & ~n5672 ;
  assign n5663 = n970 & ~n5662 ;
  assign n5674 = \InstQueue_reg[6][6]/NET0131  & ~n3933 ;
  assign n5675 = ~n5663 & ~n5674 ;
  assign n5676 = ~n5673 & n5675 ;
  assign n5677 = ~n5670 & n5676 ;
  assign n5683 = n4141 & n5182 ;
  assign n5684 = n4163 & n5185 ;
  assign n5685 = ~n5683 & ~n5684 ;
  assign n5686 = \DataWidth_reg[1]/NET0131  & ~n5685 ;
  assign n5678 = \Datai[3]_pad  & ~n4207 ;
  assign n5679 = \InstQueue_reg[7][3]/NET0131  & ~n3948 ;
  assign n5680 = ~n4185 & n5679 ;
  assign n5681 = ~n5678 & ~n5680 ;
  assign n5687 = ~n4217 & ~n5681 ;
  assign n5688 = ~n5686 & ~n5687 ;
  assign n5689 = n952 & ~n5688 ;
  assign n5690 = ~n632 & n3948 ;
  assign n5691 = ~n5679 & ~n5690 ;
  assign n5692 = n993 & ~n5691 ;
  assign n5682 = n970 & ~n5681 ;
  assign n5693 = \InstQueue_reg[7][3]/NET0131  & ~n3933 ;
  assign n5694 = ~n5682 & ~n5693 ;
  assign n5695 = ~n5692 & n5694 ;
  assign n5696 = ~n5689 & n5695 ;
  assign n5702 = n4141 & n5205 ;
  assign n5703 = n4163 & n5208 ;
  assign n5704 = ~n5702 & ~n5703 ;
  assign n5705 = \DataWidth_reg[1]/NET0131  & ~n5704 ;
  assign n5697 = \Datai[6]_pad  & ~n4207 ;
  assign n5698 = \InstQueue_reg[7][6]/NET0131  & ~n3948 ;
  assign n5699 = ~n4185 & n5698 ;
  assign n5700 = ~n5697 & ~n5699 ;
  assign n5706 = ~n4217 & ~n5700 ;
  assign n5707 = ~n5705 & ~n5706 ;
  assign n5708 = n952 & ~n5707 ;
  assign n5709 = ~n537 & n3948 ;
  assign n5710 = ~n5698 & ~n5709 ;
  assign n5711 = n993 & ~n5710 ;
  assign n5701 = n970 & ~n5700 ;
  assign n5712 = \InstQueue_reg[7][6]/NET0131  & ~n3933 ;
  assign n5713 = ~n5701 & ~n5712 ;
  assign n5714 = ~n5711 & n5713 ;
  assign n5715 = ~n5708 & n5714 ;
  assign n5721 = n4163 & n5182 ;
  assign n5722 = n4185 & n5185 ;
  assign n5723 = ~n5721 & ~n5722 ;
  assign n5724 = \DataWidth_reg[1]/NET0131  & ~n5723 ;
  assign n5716 = \Datai[3]_pad  & ~n3954 ;
  assign n5717 = \InstQueue_reg[8][3]/NET0131  & ~n3950 ;
  assign n5718 = ~n3948 & n5717 ;
  assign n5719 = ~n5716 & ~n5718 ;
  assign n5725 = ~n4237 & ~n5719 ;
  assign n5726 = ~n5724 & ~n5725 ;
  assign n5727 = n952 & ~n5726 ;
  assign n5728 = ~n632 & n3950 ;
  assign n5729 = ~n5717 & ~n5728 ;
  assign n5730 = n993 & ~n5729 ;
  assign n5720 = n970 & ~n5719 ;
  assign n5731 = \InstQueue_reg[8][3]/NET0131  & ~n3933 ;
  assign n5732 = ~n5720 & ~n5731 ;
  assign n5733 = ~n5730 & n5732 ;
  assign n5734 = ~n5727 & n5733 ;
  assign n5740 = n4163 & n5205 ;
  assign n5741 = n4185 & n5208 ;
  assign n5742 = ~n5740 & ~n5741 ;
  assign n5743 = \DataWidth_reg[1]/NET0131  & ~n5742 ;
  assign n5735 = \Datai[6]_pad  & ~n3954 ;
  assign n5736 = \InstQueue_reg[8][6]/NET0131  & ~n3950 ;
  assign n5737 = ~n3948 & n5736 ;
  assign n5738 = ~n5735 & ~n5737 ;
  assign n5744 = ~n4237 & ~n5738 ;
  assign n5745 = ~n5743 & ~n5744 ;
  assign n5746 = n952 & ~n5745 ;
  assign n5747 = ~n537 & n3950 ;
  assign n5748 = ~n5736 & ~n5747 ;
  assign n5749 = n993 & ~n5748 ;
  assign n5739 = n970 & ~n5738 ;
  assign n5750 = \InstQueue_reg[8][6]/NET0131  & ~n3933 ;
  assign n5751 = ~n5739 & ~n5750 ;
  assign n5752 = ~n5749 & n5751 ;
  assign n5753 = ~n5746 & n5752 ;
  assign n5759 = n4185 & n5182 ;
  assign n5760 = n3948 & n5185 ;
  assign n5761 = ~n5759 & ~n5760 ;
  assign n5762 = \DataWidth_reg[1]/NET0131  & ~n5761 ;
  assign n5754 = \Datai[3]_pad  & ~n3978 ;
  assign n5755 = \InstQueue_reg[9][3]/NET0131  & ~n3941 ;
  assign n5756 = ~n3950 & n5755 ;
  assign n5757 = ~n5754 & ~n5756 ;
  assign n5763 = ~n4257 & ~n5757 ;
  assign n5764 = ~n5762 & ~n5763 ;
  assign n5765 = n952 & ~n5764 ;
  assign n5766 = ~n632 & n3941 ;
  assign n5767 = ~n5755 & ~n5766 ;
  assign n5768 = n993 & ~n5767 ;
  assign n5758 = n970 & ~n5757 ;
  assign n5769 = \InstQueue_reg[9][3]/NET0131  & ~n3933 ;
  assign n5770 = ~n5758 & ~n5769 ;
  assign n5771 = ~n5768 & n5770 ;
  assign n5772 = ~n5765 & n5771 ;
  assign n5778 = n4185 & n5205 ;
  assign n5779 = n3948 & n5208 ;
  assign n5780 = ~n5778 & ~n5779 ;
  assign n5781 = \DataWidth_reg[1]/NET0131  & ~n5780 ;
  assign n5773 = \Datai[6]_pad  & ~n3978 ;
  assign n5774 = \InstQueue_reg[9][6]/NET0131  & ~n3941 ;
  assign n5775 = ~n3950 & n5774 ;
  assign n5776 = ~n5773 & ~n5775 ;
  assign n5782 = ~n4257 & ~n5776 ;
  assign n5783 = ~n5781 & ~n5782 ;
  assign n5784 = n952 & ~n5783 ;
  assign n5785 = ~n537 & n3941 ;
  assign n5786 = ~n5774 & ~n5785 ;
  assign n5787 = n993 & ~n5786 ;
  assign n5777 = n970 & ~n5776 ;
  assign n5788 = \InstQueue_reg[9][6]/NET0131  & ~n3933 ;
  assign n5789 = ~n5777 & ~n5788 ;
  assign n5790 = ~n5787 & n5789 ;
  assign n5791 = ~n5784 & n5790 ;
  assign n5794 = n948 & ~n3496 ;
  assign n5793 = ~n982 & n994 ;
  assign n5795 = ~n952 & n3639 ;
  assign n5796 = n5793 & n5795 ;
  assign n5797 = ~n5794 & n5796 ;
  assign n5798 = \PhyAddrPointer_reg[0]/NET0131  & ~n5797 ;
  assign n5792 = n948 & ~n3552 ;
  assign n5799 = ~n3559 & ~n5792 ;
  assign n5800 = ~n5798 & n5799 ;
  assign n5823 = \PhyAddrPointer_reg[0]/NET0131  & n2036 ;
  assign n5825 = \PhyAddrPointer_reg[1]/NET0131  & n5823 ;
  assign n5824 = ~\PhyAddrPointer_reg[1]/NET0131  & ~n5823 ;
  assign n5826 = ~\DataWidth_reg[1]/NET0131  & ~n5824 ;
  assign n5827 = ~n5825 & n5826 ;
  assign n5822 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[1]/NET0131  ;
  assign n5828 = n952 & ~n5822 ;
  assign n5829 = ~n5827 & n5828 ;
  assign n5802 = \rEIP_reg[1]/NET0131  & ~n4650 ;
  assign n5803 = ~\EBX_reg[1]/NET0131  & ~n4720 ;
  assign n5804 = n742 & ~n5803 ;
  assign n5807 = ~n3460 & ~n4689 ;
  assign n5808 = \EBX_reg[31]/NET0131  & n5807 ;
  assign n5809 = \EBX_reg[1]/NET0131  & ~\EBX_reg[31]/NET0131  ;
  assign n5810 = ~n4684 & ~n5809 ;
  assign n5811 = ~n5808 & n5810 ;
  assign n5812 = n736 & ~n5811 ;
  assign n5813 = ~n5804 & ~n5812 ;
  assign n5814 = \rEIP_reg[1]/NET0131  & n4684 ;
  assign n5815 = ~n5813 & ~n5814 ;
  assign n5805 = n833 & n5804 ;
  assign n5806 = n740 & ~n819 ;
  assign n5816 = ~n5805 & ~n5806 ;
  assign n5817 = ~n5815 & n5816 ;
  assign n5818 = n825 & ~n5817 ;
  assign n5819 = ~n5802 & ~n5818 ;
  assign n5820 = n948 & ~n5819 ;
  assign n5801 = \PhyAddrPointer_reg[1]/NET0131  & n981 ;
  assign n5821 = \rEIP_reg[1]/NET0131  & ~n4647 ;
  assign n5830 = ~n5801 & ~n5821 ;
  assign n5831 = ~n5820 & n5830 ;
  assign n5832 = ~n5829 & n5831 ;
  assign n5857 = n2016 & n4632 ;
  assign n5858 = n2036 & ~n5857 ;
  assign n5860 = ~n2640 & n5858 ;
  assign n5859 = n2640 & ~n5858 ;
  assign n5861 = ~\DataWidth_reg[1]/NET0131  & ~n5859 ;
  assign n5862 = ~n5860 & n5861 ;
  assign n5856 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[20]/NET0131  ;
  assign n5863 = n952 & ~n5856 ;
  assign n5864 = ~n5862 & n5863 ;
  assign n5835 = \rEIP_reg[20]/NET0131  & ~n4650 ;
  assign n5840 = ~\EBX_reg[20]/NET0131  & ~n4720 ;
  assign n5841 = n742 & ~n5840 ;
  assign n5845 = \EBX_reg[31]/NET0131  & ~n4707 ;
  assign n5847 = ~\EBX_reg[20]/NET0131  & n5845 ;
  assign n5846 = \EBX_reg[20]/NET0131  & ~n5845 ;
  assign n5848 = ~n4684 & ~n5846 ;
  assign n5849 = ~n5847 & n5848 ;
  assign n5850 = n736 & ~n5849 ;
  assign n5851 = ~n5841 & ~n5850 ;
  assign n5836 = n4667 & n4669 ;
  assign n5837 = ~\rEIP_reg[20]/NET0131  & ~n5836 ;
  assign n5838 = \rEIP_reg[20]/NET0131  & n5836 ;
  assign n5839 = ~n5837 & ~n5838 ;
  assign n5842 = n833 & n5841 ;
  assign n5843 = n4684 & ~n5842 ;
  assign n5844 = ~n5839 & n5843 ;
  assign n5852 = n825 & ~n5844 ;
  assign n5853 = ~n5851 & n5852 ;
  assign n5854 = ~n5835 & ~n5853 ;
  assign n5855 = n948 & ~n5854 ;
  assign n5833 = \rEIP_reg[20]/NET0131  & ~n4647 ;
  assign n5834 = \PhyAddrPointer_reg[20]/NET0131  & n981 ;
  assign n5865 = ~n5833 & ~n5834 ;
  assign n5866 = ~n5855 & n5865 ;
  assign n5867 = ~n5864 & n5866 ;
  assign n5888 = ~\PhyAddrPointer_reg[21]/NET0131  & ~n2639 ;
  assign n5889 = ~n2393 & ~n5888 ;
  assign n5890 = ~\PhyAddrPointer_reg[0]/NET0131  & \PhyAddrPointer_reg[1]/NET0131  ;
  assign n5891 = n2005 & n5890 ;
  assign n5892 = \PhyAddrPointer_reg[4]/NET0131  & n5891 ;
  assign n5893 = n2010 & n5892 ;
  assign n5894 = n2639 & n5893 ;
  assign n5895 = n2036 & ~n5894 ;
  assign n5897 = ~n5889 & n5895 ;
  assign n5896 = n5889 & ~n5895 ;
  assign n5898 = ~\DataWidth_reg[1]/NET0131  & ~n5896 ;
  assign n5899 = ~n5897 & n5898 ;
  assign n5887 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[21]/NET0131  ;
  assign n5900 = n952 & ~n5887 ;
  assign n5901 = ~n5899 & n5900 ;
  assign n5871 = ~\EBX_reg[20]/NET0131  & n4707 ;
  assign n5872 = \EBX_reg[31]/NET0131  & ~n5871 ;
  assign n5874 = ~\EBX_reg[21]/NET0131  & n5872 ;
  assign n5873 = \EBX_reg[21]/NET0131  & ~n5872 ;
  assign n5875 = ~n4684 & ~n5873 ;
  assign n5876 = ~n5874 & n5875 ;
  assign n5868 = ~\rEIP_reg[21]/NET0131  & ~n5838 ;
  assign n5869 = ~n4672 & ~n5868 ;
  assign n5870 = n4684 & ~n5869 ;
  assign n5877 = n1719 & ~n5870 ;
  assign n5878 = ~n5876 & n5877 ;
  assign n5879 = \rEIP_reg[21]/NET0131  & ~n4650 ;
  assign n5881 = ~n833 & n5870 ;
  assign n5880 = ~\EBX_reg[21]/NET0131  & ~n4720 ;
  assign n5882 = n3798 & ~n5880 ;
  assign n5883 = ~n5881 & n5882 ;
  assign n5884 = ~n5879 & ~n5883 ;
  assign n5885 = ~n5878 & n5884 ;
  assign n5886 = n948 & ~n5885 ;
  assign n5902 = \rEIP_reg[21]/NET0131  & ~n4647 ;
  assign n5903 = \PhyAddrPointer_reg[21]/NET0131  & n981 ;
  assign n5904 = ~n5902 & ~n5903 ;
  assign n5905 = ~n5886 & n5904 ;
  assign n5906 = ~n5901 & n5905 ;
  assign n5930 = n2036 & ~n4633 ;
  assign n5932 = ~n2665 & n5930 ;
  assign n5931 = n2665 & ~n5930 ;
  assign n5933 = ~\DataWidth_reg[1]/NET0131  & ~n5931 ;
  assign n5934 = ~n5932 & n5933 ;
  assign n5929 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[22]/NET0131  ;
  assign n5935 = n952 & ~n5929 ;
  assign n5936 = ~n5934 & n5935 ;
  assign n5916 = ~\EBX_reg[21]/NET0131  & n5871 ;
  assign n5917 = \EBX_reg[31]/NET0131  & ~n5916 ;
  assign n5919 = ~\EBX_reg[22]/NET0131  & n5917 ;
  assign n5918 = \EBX_reg[22]/NET0131  & ~n5917 ;
  assign n5920 = ~n4684 & ~n5918 ;
  assign n5921 = ~n5919 & n5920 ;
  assign n5909 = ~\rEIP_reg[22]/NET0131  & ~n4672 ;
  assign n5910 = \rEIP_reg[22]/NET0131  & n4672 ;
  assign n5911 = ~n5909 & ~n5910 ;
  assign n5915 = n4684 & ~n5911 ;
  assign n5922 = n1719 & ~n5915 ;
  assign n5923 = ~n5921 & n5922 ;
  assign n5907 = \rEIP_reg[22]/NET0131  & ~n4650 ;
  assign n5912 = n4720 & ~n5911 ;
  assign n5908 = ~\EBX_reg[22]/NET0131  & ~n4720 ;
  assign n5913 = n3798 & ~n5908 ;
  assign n5914 = ~n5912 & n5913 ;
  assign n5924 = ~n5907 & ~n5914 ;
  assign n5925 = ~n5923 & n5924 ;
  assign n5926 = n948 & ~n5925 ;
  assign n5927 = \PhyAddrPointer_reg[22]/NET0131  & n981 ;
  assign n5928 = \rEIP_reg[22]/NET0131  & ~n4647 ;
  assign n5937 = ~n5927 & ~n5928 ;
  assign n5938 = ~n5926 & n5937 ;
  assign n5939 = ~n5936 & n5938 ;
  assign n5960 = n2036 & ~n4634 ;
  assign n5962 = ~n2397 & n5960 ;
  assign n5961 = n2397 & ~n5960 ;
  assign n5963 = ~\DataWidth_reg[1]/NET0131  & ~n5961 ;
  assign n5964 = ~n5962 & n5963 ;
  assign n5959 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[23]/NET0131  ;
  assign n5965 = n952 & ~n5959 ;
  assign n5966 = ~n5964 & n5965 ;
  assign n5948 = ~\EBX_reg[22]/NET0131  & n5916 ;
  assign n5949 = \EBX_reg[31]/NET0131  & ~n5948 ;
  assign n5951 = ~\EBX_reg[23]/NET0131  & n5949 ;
  assign n5950 = \EBX_reg[23]/NET0131  & ~n5949 ;
  assign n5952 = ~n4684 & ~n5950 ;
  assign n5953 = ~n5951 & n5952 ;
  assign n5942 = ~\rEIP_reg[23]/NET0131  & ~n5910 ;
  assign n5943 = ~n4673 & ~n5942 ;
  assign n5947 = n4684 & ~n5943 ;
  assign n5954 = n1719 & ~n5947 ;
  assign n5955 = ~n5953 & n5954 ;
  assign n5940 = \rEIP_reg[23]/NET0131  & ~n4650 ;
  assign n5944 = n4720 & ~n5943 ;
  assign n5941 = ~\EBX_reg[23]/NET0131  & ~n4720 ;
  assign n5945 = n3798 & ~n5941 ;
  assign n5946 = ~n5944 & n5945 ;
  assign n5956 = ~n5940 & ~n5946 ;
  assign n5957 = ~n5955 & n5956 ;
  assign n5958 = n948 & ~n5957 ;
  assign n5967 = \PhyAddrPointer_reg[23]/NET0131  & n981 ;
  assign n5968 = \rEIP_reg[23]/NET0131  & ~n4647 ;
  assign n5969 = ~n5967 & ~n5968 ;
  assign n5970 = ~n5958 & n5969 ;
  assign n5971 = ~n5966 & n5970 ;
  assign n6001 = ~n2397 & n4634 ;
  assign n6002 = n2036 & ~n6001 ;
  assign n6004 = ~n2683 & n6002 ;
  assign n6003 = n2683 & ~n6002 ;
  assign n6005 = ~\DataWidth_reg[1]/NET0131  & ~n6003 ;
  assign n6006 = ~n6004 & n6005 ;
  assign n6000 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[24]/NET0131  ;
  assign n6007 = n952 & ~n6000 ;
  assign n6008 = ~n6006 & n6007 ;
  assign n5990 = \EBX_reg[31]/NET0131  & ~n4711 ;
  assign n5992 = ~\EBX_reg[24]/NET0131  & n5990 ;
  assign n5991 = \EBX_reg[24]/NET0131  & ~n5990 ;
  assign n5993 = ~n4684 & ~n5991 ;
  assign n5994 = ~n5992 & n5993 ;
  assign n5977 = \rEIP_reg[24]/NET0131  & n4673 ;
  assign n5978 = ~\rEIP_reg[24]/NET0131  & ~n4673 ;
  assign n5979 = ~n5977 & ~n5978 ;
  assign n5980 = n4684 & ~n5979 ;
  assign n5995 = n1719 & ~n5980 ;
  assign n5996 = ~n5994 & n5995 ;
  assign n5981 = ~\EBX_reg[24]/NET0131  & ~n4684 ;
  assign n5982 = n895 & ~n5981 ;
  assign n5983 = ~n5980 & n5982 ;
  assign n5974 = \rEIP_reg[24]/NET0131  & ~n825 ;
  assign n5975 = n825 & n833 ;
  assign n5976 = \EBX_reg[24]/NET0131  & n5975 ;
  assign n5984 = ~n5974 & ~n5976 ;
  assign n5985 = ~n5983 & n5984 ;
  assign n5986 = n742 & ~n5985 ;
  assign n5987 = ~n740 & n742 ;
  assign n5988 = ~n4650 & ~n5987 ;
  assign n5989 = \rEIP_reg[24]/NET0131  & n5988 ;
  assign n5997 = ~n5986 & ~n5989 ;
  assign n5998 = ~n5996 & n5997 ;
  assign n5999 = n948 & ~n5998 ;
  assign n5972 = \PhyAddrPointer_reg[24]/NET0131  & n981 ;
  assign n5973 = \rEIP_reg[24]/NET0131  & ~n4647 ;
  assign n6009 = ~n5972 & ~n5973 ;
  assign n6010 = ~n5999 & n6009 ;
  assign n6011 = ~n6008 & n6010 ;
  assign n6035 = n2402 & n5894 ;
  assign n6036 = n4635 & n6035 ;
  assign n6037 = n2036 & ~n6036 ;
  assign n6039 = ~n2869 & n6037 ;
  assign n6038 = n2869 & ~n6037 ;
  assign n6040 = ~\DataWidth_reg[1]/NET0131  & ~n6038 ;
  assign n6041 = ~n6039 & n6040 ;
  assign n6034 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[25]/NET0131  ;
  assign n6042 = n952 & ~n6034 ;
  assign n6043 = ~n6041 & n6042 ;
  assign n6019 = ~\EBX_reg[24]/NET0131  & n4711 ;
  assign n6020 = \EBX_reg[31]/NET0131  & ~n6019 ;
  assign n6022 = ~\EBX_reg[25]/NET0131  & n6020 ;
  assign n6021 = \EBX_reg[25]/NET0131  & ~n6020 ;
  assign n6023 = ~n4684 & ~n6021 ;
  assign n6024 = ~n6022 & n6023 ;
  assign n6015 = ~\rEIP_reg[25]/NET0131  & ~n5977 ;
  assign n6016 = \rEIP_reg[25]/NET0131  & n5977 ;
  assign n6017 = ~n6015 & ~n6016 ;
  assign n6018 = n4684 & ~n6017 ;
  assign n6025 = n1719 & ~n6018 ;
  assign n6026 = ~n6024 & n6025 ;
  assign n6014 = \rEIP_reg[25]/NET0131  & ~n4650 ;
  assign n6028 = n4720 & ~n6017 ;
  assign n6027 = ~\EBX_reg[25]/NET0131  & ~n4720 ;
  assign n6029 = n3798 & ~n6027 ;
  assign n6030 = ~n6028 & n6029 ;
  assign n6031 = ~n6014 & ~n6030 ;
  assign n6032 = ~n6026 & n6031 ;
  assign n6033 = n948 & ~n6032 ;
  assign n6012 = \PhyAddrPointer_reg[25]/NET0131  & n981 ;
  assign n6013 = \rEIP_reg[25]/NET0131  & ~n4647 ;
  assign n6044 = ~n6012 & ~n6013 ;
  assign n6045 = ~n6033 & n6044 ;
  assign n6046 = ~n6043 & n6045 ;
  assign n6069 = n2036 & ~n4637 ;
  assign n6071 = ~n2716 & n6069 ;
  assign n6070 = n2716 & ~n6069 ;
  assign n6072 = ~\DataWidth_reg[1]/NET0131  & ~n6070 ;
  assign n6073 = ~n6071 & n6072 ;
  assign n6068 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[26]/NET0131  ;
  assign n6074 = n952 & ~n6068 ;
  assign n6075 = ~n6073 & n6074 ;
  assign n6053 = n4688 & n4711 ;
  assign n6054 = \EBX_reg[31]/NET0131  & ~n6053 ;
  assign n6056 = ~\EBX_reg[26]/NET0131  & n6054 ;
  assign n6055 = \EBX_reg[26]/NET0131  & ~n6054 ;
  assign n6057 = ~n4684 & ~n6055 ;
  assign n6058 = ~n6056 & n6057 ;
  assign n6050 = ~\rEIP_reg[26]/NET0131  & ~n6016 ;
  assign n6051 = ~n4676 & ~n6050 ;
  assign n6052 = n4684 & ~n6051 ;
  assign n6059 = n1719 & ~n6052 ;
  assign n6060 = ~n6058 & n6059 ;
  assign n6049 = \rEIP_reg[26]/NET0131  & ~n4650 ;
  assign n6062 = n4720 & ~n6051 ;
  assign n6061 = ~\EBX_reg[26]/NET0131  & ~n4720 ;
  assign n6063 = n3798 & ~n6061 ;
  assign n6064 = ~n6062 & n6063 ;
  assign n6065 = ~n6049 & ~n6064 ;
  assign n6066 = ~n6060 & n6065 ;
  assign n6067 = n948 & ~n6066 ;
  assign n6047 = \PhyAddrPointer_reg[26]/NET0131  & n981 ;
  assign n6048 = \rEIP_reg[26]/NET0131  & ~n4647 ;
  assign n6076 = ~n6047 & ~n6048 ;
  assign n6077 = ~n6067 & n6076 ;
  assign n6078 = ~n6075 & n6077 ;
  assign n6101 = n2036 & ~n4638 ;
  assign n6103 = ~n2422 & n6101 ;
  assign n6102 = n2422 & ~n6101 ;
  assign n6104 = ~\DataWidth_reg[1]/NET0131  & ~n6102 ;
  assign n6105 = ~n6103 & n6104 ;
  assign n6100 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[27]/NET0131  ;
  assign n6106 = n952 & ~n6100 ;
  assign n6107 = ~n6105 & n6106 ;
  assign n6086 = \EBX_reg[31]/NET0131  & ~n4713 ;
  assign n6088 = ~\EBX_reg[27]/NET0131  & n6086 ;
  assign n6087 = \EBX_reg[27]/NET0131  & ~n6086 ;
  assign n6089 = ~n4684 & ~n6087 ;
  assign n6090 = ~n6088 & n6089 ;
  assign n6082 = ~\rEIP_reg[27]/NET0131  & ~n4676 ;
  assign n6083 = \rEIP_reg[27]/NET0131  & n4676 ;
  assign n6084 = ~n6082 & ~n6083 ;
  assign n6085 = n4684 & ~n6084 ;
  assign n6091 = n1719 & ~n6085 ;
  assign n6092 = ~n6090 & n6091 ;
  assign n6081 = \rEIP_reg[27]/NET0131  & ~n4650 ;
  assign n6094 = ~n833 & n6085 ;
  assign n6093 = ~\EBX_reg[27]/NET0131  & ~n4720 ;
  assign n6095 = n3798 & ~n6093 ;
  assign n6096 = ~n6094 & n6095 ;
  assign n6097 = ~n6081 & ~n6096 ;
  assign n6098 = ~n6092 & n6097 ;
  assign n6099 = n948 & ~n6098 ;
  assign n6079 = \rEIP_reg[27]/NET0131  & ~n4647 ;
  assign n6080 = \PhyAddrPointer_reg[27]/NET0131  & n981 ;
  assign n6108 = ~n6079 & ~n6080 ;
  assign n6109 = ~n6099 & n6108 ;
  assign n6110 = ~n6107 & n6109 ;
  assign n6134 = ~n2422 & n4638 ;
  assign n6135 = n2036 & ~n6134 ;
  assign n6137 = n2441 & ~n6135 ;
  assign n6136 = ~n2441 & n6135 ;
  assign n6138 = ~\DataWidth_reg[1]/NET0131  & ~n6136 ;
  assign n6139 = ~n6137 & n6138 ;
  assign n6133 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[28]/NET0131  ;
  assign n6140 = n952 & ~n6133 ;
  assign n6141 = ~n6139 & n6140 ;
  assign n6115 = ~\EBX_reg[27]/NET0131  & n4713 ;
  assign n6116 = \EBX_reg[31]/NET0131  & ~n6115 ;
  assign n6118 = ~\EBX_reg[28]/NET0131  & n6116 ;
  assign n6117 = \EBX_reg[28]/NET0131  & ~n6116 ;
  assign n6119 = ~n4684 & ~n6117 ;
  assign n6120 = ~n6118 & n6119 ;
  assign n6111 = ~\rEIP_reg[28]/NET0131  & ~n6083 ;
  assign n6112 = n4676 & n4677 ;
  assign n6113 = ~n6111 & ~n6112 ;
  assign n6114 = n4684 & ~n6113 ;
  assign n6121 = n1719 & ~n6114 ;
  assign n6122 = ~n6120 & n6121 ;
  assign n6123 = \rEIP_reg[28]/NET0131  & ~n4650 ;
  assign n6125 = n4720 & ~n6113 ;
  assign n6124 = ~\EBX_reg[28]/NET0131  & ~n4720 ;
  assign n6126 = n3798 & ~n6124 ;
  assign n6127 = ~n6125 & n6126 ;
  assign n6128 = ~n6123 & ~n6127 ;
  assign n6129 = ~n6122 & n6128 ;
  assign n6130 = n948 & ~n6129 ;
  assign n6131 = \PhyAddrPointer_reg[28]/NET0131  & n981 ;
  assign n6132 = \rEIP_reg[28]/NET0131  & ~n4647 ;
  assign n6142 = ~n6131 & ~n6132 ;
  assign n6143 = ~n6130 & n6142 ;
  assign n6144 = ~n6141 & n6143 ;
  assign n6157 = ~\EBX_reg[28]/NET0131  & n6115 ;
  assign n6158 = \EBX_reg[31]/NET0131  & ~n6157 ;
  assign n6160 = ~\EBX_reg[29]/NET0131  & n6158 ;
  assign n6159 = \EBX_reg[29]/NET0131  & ~n6158 ;
  assign n6161 = ~n4684 & ~n6159 ;
  assign n6162 = ~n6160 & n6161 ;
  assign n6146 = ~\rEIP_reg[29]/NET0131  & ~n6112 ;
  assign n6147 = n4676 & n4678 ;
  assign n6148 = ~n6146 & ~n6147 ;
  assign n6149 = n4684 & ~n6148 ;
  assign n6163 = n1719 & ~n6149 ;
  assign n6164 = ~n6162 & n6163 ;
  assign n6145 = \rEIP_reg[29]/NET0131  & n5988 ;
  assign n6150 = n895 & ~n4687 ;
  assign n6151 = ~n6149 & n6150 ;
  assign n6152 = \EBX_reg[29]/NET0131  & n5975 ;
  assign n6153 = \rEIP_reg[29]/NET0131  & ~n825 ;
  assign n6154 = ~n6152 & ~n6153 ;
  assign n6155 = ~n6151 & n6154 ;
  assign n6156 = n742 & ~n6155 ;
  assign n6165 = ~n6145 & ~n6156 ;
  assign n6166 = ~n6164 & n6165 ;
  assign n6167 = n948 & ~n6166 ;
  assign n6169 = ~n2716 & ~n2869 ;
  assign n6170 = n6036 & n6169 ;
  assign n6171 = n4639 & n6170 ;
  assign n6172 = n2036 & ~n6171 ;
  assign n6174 = n2483 & ~n6172 ;
  assign n6173 = ~n2483 & n6172 ;
  assign n6175 = ~\DataWidth_reg[1]/NET0131  & ~n6173 ;
  assign n6176 = ~n6174 & n6175 ;
  assign n6168 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[29]/NET0131  ;
  assign n6177 = n952 & ~n6168 ;
  assign n6178 = ~n6176 & n6177 ;
  assign n6179 = \PhyAddrPointer_reg[29]/NET0131  & n981 ;
  assign n6180 = \rEIP_reg[29]/NET0131  & ~n4647 ;
  assign n6181 = ~n6179 & ~n6180 ;
  assign n6182 = ~n6178 & n6181 ;
  assign n6183 = ~n6167 & n6182 ;
  assign n6185 = n2036 & ~n5890 ;
  assign n6187 = ~n4269 & n6185 ;
  assign n6186 = n4269 & ~n6185 ;
  assign n6188 = ~\DataWidth_reg[1]/NET0131  & ~n6186 ;
  assign n6189 = ~n6187 & n6188 ;
  assign n6184 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[2]/NET0131  ;
  assign n6190 = n952 & ~n6184 ;
  assign n6191 = ~n6189 & n6190 ;
  assign n6194 = \rEIP_reg[2]/NET0131  & ~n4650 ;
  assign n6207 = \EBX_reg[2]/NET0131  & ~n4720 ;
  assign n6196 = ~\rEIP_reg[1]/NET0131  & ~\rEIP_reg[2]/NET0131  ;
  assign n6197 = ~\DataWidth_reg[1]/NET0131  & ~n4653 ;
  assign n6198 = ~n6196 & n6197 ;
  assign n6208 = n861 & n6198 ;
  assign n6209 = ~n6207 & ~n6208 ;
  assign n6210 = n742 & ~n6209 ;
  assign n6195 = n740 & n884 ;
  assign n6199 = ~READY_n_pad & n6198 ;
  assign n6200 = \EBX_reg[31]/NET0131  & ~n4689 ;
  assign n6202 = \EBX_reg[2]/NET0131  & n6200 ;
  assign n6201 = ~\EBX_reg[2]/NET0131  & ~n6200 ;
  assign n6203 = ~n4684 & ~n6201 ;
  assign n6204 = ~n6202 & n6203 ;
  assign n6205 = ~n6199 & ~n6204 ;
  assign n6206 = n736 & ~n6205 ;
  assign n6211 = ~n6195 & ~n6206 ;
  assign n6212 = ~n6210 & n6211 ;
  assign n6213 = n825 & ~n6212 ;
  assign n6214 = ~n6194 & ~n6213 ;
  assign n6215 = n948 & ~n6214 ;
  assign n6192 = \PhyAddrPointer_reg[2]/NET0131  & n981 ;
  assign n6193 = \rEIP_reg[2]/NET0131  & ~n4647 ;
  assign n6216 = ~n6192 & ~n6193 ;
  assign n6217 = ~n6215 & n6216 ;
  assign n6218 = ~n6191 & n6217 ;
  assign n6219 = ~\rEIP_reg[30]/NET0131  & ~n6147 ;
  assign n6220 = ~n4680 & n4684 ;
  assign n6221 = ~n6219 & n6220 ;
  assign n6222 = ~\EBX_reg[26]/NET0131  & ~\EBX_reg[29]/NET0131  ;
  assign n6223 = n4686 & n6222 ;
  assign n6224 = n6053 & n6223 ;
  assign n6225 = \EBX_reg[31]/NET0131  & ~n6224 ;
  assign n6227 = \EBX_reg[30]/NET0131  & n6225 ;
  assign n6226 = ~\EBX_reg[30]/NET0131  & ~n6225 ;
  assign n6228 = ~n4684 & ~n6226 ;
  assign n6229 = ~n6227 & n6228 ;
  assign n6230 = ~n6221 & ~n6229 ;
  assign n6231 = n1719 & ~n6230 ;
  assign n6232 = \rEIP_reg[30]/NET0131  & n5988 ;
  assign n6233 = \EBX_reg[30]/NET0131  & ~n4684 ;
  assign n6234 = ~n6221 & ~n6233 ;
  assign n6235 = n895 & ~n6234 ;
  assign n6236 = \EBX_reg[30]/NET0131  & n5975 ;
  assign n6237 = \rEIP_reg[30]/NET0131  & ~n825 ;
  assign n6238 = ~n6236 & ~n6237 ;
  assign n6239 = ~n6235 & n6238 ;
  assign n6240 = n742 & ~n6239 ;
  assign n6241 = ~n6232 & ~n6240 ;
  assign n6242 = ~n6231 & n6241 ;
  assign n6243 = n948 & ~n6242 ;
  assign n6245 = n2036 & ~n4641 ;
  assign n6247 = n2211 & ~n6245 ;
  assign n6246 = ~n2211 & n6245 ;
  assign n6248 = ~\DataWidth_reg[1]/NET0131  & ~n6246 ;
  assign n6249 = ~n6247 & n6248 ;
  assign n6244 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[30]/NET0131  ;
  assign n6250 = n952 & ~n6244 ;
  assign n6251 = ~n6249 & n6250 ;
  assign n6252 = \PhyAddrPointer_reg[30]/NET0131  & n981 ;
  assign n6253 = \rEIP_reg[30]/NET0131  & ~n4647 ;
  assign n6254 = ~n6252 & ~n6253 ;
  assign n6255 = ~n6251 & n6254 ;
  assign n6256 = ~n6243 & n6255 ;
  assign n6258 = ~\PhyAddrPointer_reg[0]/NET0131  & n3506 ;
  assign n6259 = n2036 & ~n6258 ;
  assign n6261 = n3671 & ~n6259 ;
  assign n6260 = ~n3671 & n6259 ;
  assign n6262 = ~\DataWidth_reg[1]/NET0131  & ~n6260 ;
  assign n6263 = ~n6261 & n6262 ;
  assign n6257 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[3]/NET0131  ;
  assign n6264 = n952 & ~n6257 ;
  assign n6265 = ~n6263 & n6264 ;
  assign n6267 = \rEIP_reg[3]/NET0131  & ~n4650 ;
  assign n6276 = \EBX_reg[31]/NET0131  & ~n4690 ;
  assign n6278 = \EBX_reg[3]/NET0131  & n6276 ;
  assign n6277 = ~\EBX_reg[3]/NET0131  & ~n6276 ;
  assign n6279 = ~n4684 & ~n6277 ;
  assign n6280 = ~n6278 & n6279 ;
  assign n6270 = ~\rEIP_reg[3]/NET0131  & ~n4653 ;
  assign n6271 = ~\DataWidth_reg[1]/NET0131  & ~n4654 ;
  assign n6272 = ~n6270 & n6271 ;
  assign n6281 = ~READY_n_pad & n6272 ;
  assign n6282 = ~n6280 & ~n6281 ;
  assign n6283 = n736 & ~n6282 ;
  assign n6268 = n740 & ~n855 ;
  assign n6269 = \EBX_reg[3]/NET0131  & ~n4720 ;
  assign n6273 = n861 & n6272 ;
  assign n6274 = ~n6269 & ~n6273 ;
  assign n6275 = n742 & ~n6274 ;
  assign n6284 = ~n6268 & ~n6275 ;
  assign n6285 = ~n6283 & n6284 ;
  assign n6286 = n825 & ~n6285 ;
  assign n6287 = ~n6267 & ~n6286 ;
  assign n6288 = n948 & ~n6287 ;
  assign n6266 = \rEIP_reg[3]/NET0131  & ~n4647 ;
  assign n6289 = ~n3669 & ~n6266 ;
  assign n6290 = ~n6288 & n6289 ;
  assign n6291 = ~n6265 & n6290 ;
  assign n6293 = n2036 & ~n5891 ;
  assign n6295 = ~n3510 & n6293 ;
  assign n6294 = n3510 & ~n6293 ;
  assign n6296 = ~\DataWidth_reg[1]/NET0131  & ~n6294 ;
  assign n6297 = ~n6295 & n6296 ;
  assign n6292 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[4]/NET0131  ;
  assign n6298 = n952 & ~n6292 ;
  assign n6299 = ~n6297 & n6298 ;
  assign n6302 = \rEIP_reg[4]/NET0131  & ~n4650 ;
  assign n6303 = \EBX_reg[31]/NET0131  & ~n4691 ;
  assign n6305 = ~\EBX_reg[4]/NET0131  & n6303 ;
  assign n6304 = \EBX_reg[4]/NET0131  & ~n6303 ;
  assign n6306 = ~n4684 & ~n6304 ;
  assign n6307 = ~n6305 & n6306 ;
  assign n6308 = ~\rEIP_reg[4]/NET0131  & ~n4654 ;
  assign n6309 = ~n4655 & ~n6308 ;
  assign n6310 = n4684 & ~n6309 ;
  assign n6311 = ~n6307 & ~n6310 ;
  assign n6312 = n1719 & n6311 ;
  assign n6313 = ~\EBX_reg[4]/NET0131  & ~n4720 ;
  assign n6314 = n4720 & ~n6309 ;
  assign n6315 = ~n6313 & ~n6314 ;
  assign n6316 = n3798 & n6315 ;
  assign n6317 = ~n6312 & ~n6316 ;
  assign n6318 = ~n6302 & n6317 ;
  assign n6319 = n948 & ~n6318 ;
  assign n6300 = ~n969 & n5793 ;
  assign n6301 = \rEIP_reg[4]/NET0131  & ~n6300 ;
  assign n6320 = \PhyAddrPointer_reg[4]/NET0131  & n981 ;
  assign n6321 = ~n1731 & ~n6320 ;
  assign n6322 = ~n6301 & n6321 ;
  assign n6323 = ~n6319 & n6322 ;
  assign n6324 = ~n6299 & n6323 ;
  assign n6326 = n2036 & ~n5892 ;
  assign n6328 = ~n3678 & n6326 ;
  assign n6327 = n3678 & ~n6326 ;
  assign n6329 = ~\DataWidth_reg[1]/NET0131  & ~n6327 ;
  assign n6330 = ~n6328 & n6329 ;
  assign n6325 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[5]/NET0131  ;
  assign n6331 = n952 & ~n6325 ;
  assign n6332 = ~n6330 & n6331 ;
  assign n6334 = \rEIP_reg[5]/NET0131  & ~n4650 ;
  assign n6335 = \EBX_reg[31]/NET0131  & ~n4692 ;
  assign n6337 = ~\EBX_reg[5]/NET0131  & n6335 ;
  assign n6336 = \EBX_reg[5]/NET0131  & ~n6335 ;
  assign n6338 = ~n4684 & ~n6336 ;
  assign n6339 = ~n6337 & n6338 ;
  assign n6340 = ~\rEIP_reg[5]/NET0131  & ~n4655 ;
  assign n6341 = ~n4656 & ~n6340 ;
  assign n6342 = n4684 & ~n6341 ;
  assign n6343 = ~n6339 & ~n6342 ;
  assign n6344 = n1719 & n6343 ;
  assign n6345 = ~\EBX_reg[5]/NET0131  & ~n4720 ;
  assign n6346 = n4720 & ~n6341 ;
  assign n6347 = ~n6345 & ~n6346 ;
  assign n6348 = n3798 & n6347 ;
  assign n6349 = ~n6344 & ~n6348 ;
  assign n6350 = ~n6334 & n6349 ;
  assign n6351 = n948 & ~n6350 ;
  assign n6333 = \rEIP_reg[5]/NET0131  & ~n6300 ;
  assign n6352 = \PhyAddrPointer_reg[5]/NET0131  & n981 ;
  assign n6353 = ~n1731 & ~n6352 ;
  assign n6354 = ~n6333 & n6353 ;
  assign n6355 = ~n6351 & n6354 ;
  assign n6356 = ~n6332 & n6355 ;
  assign n6358 = ~\PhyAddrPointer_reg[0]/NET0131  & n3004 ;
  assign n6359 = n2036 & ~n6358 ;
  assign n6361 = n3699 & ~n6359 ;
  assign n6360 = ~n3699 & n6359 ;
  assign n6362 = ~\DataWidth_reg[1]/NET0131  & ~n6360 ;
  assign n6363 = ~n6361 & n6362 ;
  assign n6357 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[6]/NET0131  ;
  assign n6364 = n952 & ~n6357 ;
  assign n6365 = ~n6363 & n6364 ;
  assign n6367 = ~\EBX_reg[6]/NET0131  & ~n4720 ;
  assign n6368 = ~\rEIP_reg[6]/NET0131  & ~n4656 ;
  assign n6369 = ~n4657 & ~n6368 ;
  assign n6370 = n4720 & ~n6369 ;
  assign n6371 = ~n6367 & ~n6370 ;
  assign n6372 = n742 & n6371 ;
  assign n6373 = n4684 & ~n6369 ;
  assign n6374 = \EBX_reg[31]/NET0131  & ~n4693 ;
  assign n6376 = ~\EBX_reg[6]/NET0131  & n6374 ;
  assign n6375 = \EBX_reg[6]/NET0131  & ~n6374 ;
  assign n6377 = ~n4684 & ~n6375 ;
  assign n6378 = ~n6376 & n6377 ;
  assign n6379 = ~n6373 & ~n6378 ;
  assign n6380 = n736 & n6379 ;
  assign n6381 = ~n6372 & ~n6380 ;
  assign n6382 = n825 & ~n6381 ;
  assign n6383 = \rEIP_reg[6]/NET0131  & ~n4650 ;
  assign n6384 = ~n6382 & ~n6383 ;
  assign n6385 = n948 & ~n6384 ;
  assign n6366 = \rEIP_reg[6]/NET0131  & ~n6300 ;
  assign n6386 = \PhyAddrPointer_reg[6]/NET0131  & n981 ;
  assign n6387 = ~n1731 & ~n6386 ;
  assign n6388 = ~n6366 & n6387 ;
  assign n6389 = ~n6385 & n6388 ;
  assign n6390 = ~n6365 & n6389 ;
  assign n6392 = ~\PhyAddrPointer_reg[0]/NET0131  & n3005 ;
  assign n6393 = n2036 & ~n6392 ;
  assign n6395 = n3007 & ~n6393 ;
  assign n6394 = ~n3007 & n6393 ;
  assign n6396 = ~\DataWidth_reg[1]/NET0131  & ~n6394 ;
  assign n6397 = ~n6395 & n6396 ;
  assign n6391 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[7]/NET0131  ;
  assign n6398 = n952 & ~n6391 ;
  assign n6399 = ~n6397 & n6398 ;
  assign n6401 = \rEIP_reg[7]/NET0131  & ~n4650 ;
  assign n6402 = ~\EBX_reg[7]/NET0131  & ~n4720 ;
  assign n6403 = ~\rEIP_reg[7]/NET0131  & ~n4657 ;
  assign n6404 = ~n4658 & ~n6403 ;
  assign n6405 = n4720 & ~n6404 ;
  assign n6406 = ~n6402 & ~n6405 ;
  assign n6407 = n3798 & n6406 ;
  assign n6408 = n4684 & ~n6404 ;
  assign n6409 = \EBX_reg[31]/NET0131  & ~n4694 ;
  assign n6411 = ~\EBX_reg[7]/NET0131  & n6409 ;
  assign n6410 = \EBX_reg[7]/NET0131  & ~n6409 ;
  assign n6412 = ~n4684 & ~n6410 ;
  assign n6413 = ~n6411 & n6412 ;
  assign n6414 = ~n6408 & ~n6413 ;
  assign n6415 = n1719 & n6414 ;
  assign n6416 = ~n6407 & ~n6415 ;
  assign n6417 = ~n6401 & n6416 ;
  assign n6418 = n948 & ~n6417 ;
  assign n6400 = \rEIP_reg[7]/NET0131  & ~n6300 ;
  assign n6419 = \PhyAddrPointer_reg[7]/NET0131  & n981 ;
  assign n6420 = ~n1731 & ~n6419 ;
  assign n6421 = ~n6400 & n6420 ;
  assign n6422 = ~n6418 & n6421 ;
  assign n6423 = ~n6399 & n6422 ;
  assign n6425 = \PhyAddrPointer_reg[7]/NET0131  & n6392 ;
  assign n6426 = n2036 & ~n6425 ;
  assign n6428 = n2881 & ~n6426 ;
  assign n6427 = ~n2881 & n6426 ;
  assign n6429 = ~\DataWidth_reg[1]/NET0131  & ~n6427 ;
  assign n6430 = ~n6428 & n6429 ;
  assign n6424 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[8]/NET0131  ;
  assign n6431 = n952 & ~n6424 ;
  assign n6432 = ~n6430 & n6431 ;
  assign n6434 = \rEIP_reg[8]/NET0131  & ~n4650 ;
  assign n6435 = ~\EBX_reg[8]/NET0131  & ~n4720 ;
  assign n6436 = ~\rEIP_reg[8]/NET0131  & ~n4658 ;
  assign n6437 = ~n4659 & ~n6436 ;
  assign n6438 = n4720 & ~n6437 ;
  assign n6439 = ~n6435 & ~n6438 ;
  assign n6440 = n742 & n6439 ;
  assign n6442 = \EBX_reg[31]/NET0131  & ~n4695 ;
  assign n6444 = ~\EBX_reg[8]/NET0131  & n6442 ;
  assign n6443 = \EBX_reg[8]/NET0131  & ~n6442 ;
  assign n6445 = ~n4684 & ~n6443 ;
  assign n6446 = ~n6444 & n6445 ;
  assign n6441 = n4684 & ~n6437 ;
  assign n6447 = n736 & ~n6441 ;
  assign n6448 = ~n6446 & n6447 ;
  assign n6449 = ~n6440 & ~n6448 ;
  assign n6450 = n825 & ~n6449 ;
  assign n6451 = ~n6434 & ~n6450 ;
  assign n6452 = n948 & ~n6451 ;
  assign n6433 = \rEIP_reg[8]/NET0131  & ~n6300 ;
  assign n6453 = \PhyAddrPointer_reg[8]/NET0131  & n981 ;
  assign n6454 = ~n1731 & ~n6453 ;
  assign n6455 = ~n6433 & n6454 ;
  assign n6456 = ~n6452 & n6455 ;
  assign n6457 = ~n6432 & n6456 ;
  assign n6459 = ~\PhyAddrPointer_reg[9]/NET0131  & ~n2880 ;
  assign n6460 = ~n2988 & ~n6459 ;
  assign n6461 = n2036 & ~n5893 ;
  assign n6463 = ~n6460 & n6461 ;
  assign n6462 = n6460 & ~n6461 ;
  assign n6464 = ~\DataWidth_reg[1]/NET0131  & ~n6462 ;
  assign n6465 = ~n6463 & n6464 ;
  assign n6458 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[9]/NET0131  ;
  assign n6466 = n952 & ~n6458 ;
  assign n6467 = ~n6465 & n6466 ;
  assign n6469 = \rEIP_reg[9]/NET0131  & ~n4650 ;
  assign n6471 = ~\rEIP_reg[9]/NET0131  & ~n4659 ;
  assign n6472 = ~n4660 & ~n6471 ;
  assign n6473 = n4720 & ~n6472 ;
  assign n6470 = ~\EBX_reg[9]/NET0131  & ~n4720 ;
  assign n6474 = n742 & ~n6470 ;
  assign n6475 = ~n6473 & n6474 ;
  assign n6477 = \EBX_reg[31]/NET0131  & ~n4696 ;
  assign n6479 = ~\EBX_reg[9]/NET0131  & n6477 ;
  assign n6478 = \EBX_reg[9]/NET0131  & ~n6477 ;
  assign n6480 = ~n4684 & ~n6478 ;
  assign n6481 = ~n6479 & n6480 ;
  assign n6476 = n4684 & ~n6472 ;
  assign n6482 = n736 & ~n6476 ;
  assign n6483 = ~n6481 & n6482 ;
  assign n6484 = ~n6475 & ~n6483 ;
  assign n6485 = n825 & ~n6484 ;
  assign n6486 = ~n6469 & ~n6485 ;
  assign n6487 = n948 & ~n6486 ;
  assign n6468 = \rEIP_reg[9]/NET0131  & ~n6300 ;
  assign n6488 = \PhyAddrPointer_reg[9]/NET0131  & n981 ;
  assign n6489 = ~n1731 & ~n6488 ;
  assign n6490 = ~n6468 & n6489 ;
  assign n6491 = ~n6487 & n6490 ;
  assign n6492 = ~n6467 & n6491 ;
  assign n6494 = \PhyAddrPointer_reg[1]/NET0131  & ~n3496 ;
  assign n6495 = n3738 & ~n6494 ;
  assign n6496 = n948 & ~n6495 ;
  assign n6497 = ~n971 & n2003 ;
  assign n6498 = \PhyAddrPointer_reg[1]/NET0131  & ~n6497 ;
  assign n6493 = ~\PhyAddrPointer_reg[1]/NET0131  & n2039 ;
  assign n6499 = ~n3718 & ~n6493 ;
  assign n6500 = ~n6498 & n6499 ;
  assign n6501 = ~n6496 & n6500 ;
  assign n6503 = n2011 & n5890 ;
  assign n6504 = n2036 & ~n6503 ;
  assign n6506 = ~n2990 & n6504 ;
  assign n6505 = n2990 & ~n6504 ;
  assign n6507 = ~\DataWidth_reg[1]/NET0131  & ~n6505 ;
  assign n6508 = ~n6506 & n6507 ;
  assign n6502 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[10]/NET0131  ;
  assign n6509 = n952 & ~n6502 ;
  assign n6510 = ~n6508 & n6509 ;
  assign n6512 = \rEIP_reg[10]/NET0131  & ~n4650 ;
  assign n6513 = ~\rEIP_reg[10]/NET0131  & ~n4660 ;
  assign n6514 = ~n4661 & ~n6513 ;
  assign n6515 = n4684 & ~n6514 ;
  assign n6516 = ~\EBX_reg[10]/NET0131  & ~n4720 ;
  assign n6517 = n742 & ~n6516 ;
  assign n6518 = \EBX_reg[31]/NET0131  & ~n4697 ;
  assign n6520 = ~\EBX_reg[10]/NET0131  & n6518 ;
  assign n6519 = \EBX_reg[10]/NET0131  & ~n6518 ;
  assign n6521 = ~n4684 & ~n6519 ;
  assign n6522 = ~n6520 & n6521 ;
  assign n6523 = n736 & ~n6522 ;
  assign n6524 = ~n6517 & ~n6523 ;
  assign n6525 = ~n6515 & ~n6524 ;
  assign n6526 = n833 & n6517 ;
  assign n6527 = ~n6525 & ~n6526 ;
  assign n6528 = n825 & ~n6527 ;
  assign n6529 = ~n6512 & ~n6528 ;
  assign n6530 = n948 & ~n6529 ;
  assign n6511 = \rEIP_reg[10]/NET0131  & ~n6300 ;
  assign n6531 = \PhyAddrPointer_reg[10]/NET0131  & n981 ;
  assign n6532 = ~n1731 & ~n6531 ;
  assign n6533 = ~n6511 & n6532 ;
  assign n6534 = ~n6530 & n6533 ;
  assign n6535 = ~n6510 & n6534 ;
  assign n6537 = ~\PhyAddrPointer_reg[0]/NET0131  & n2579 ;
  assign n6538 = n2036 & ~n6537 ;
  assign n6540 = ~n2581 & n6538 ;
  assign n6539 = n2581 & ~n6538 ;
  assign n6541 = ~\DataWidth_reg[1]/NET0131  & ~n6539 ;
  assign n6542 = ~n6540 & n6541 ;
  assign n6536 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[11]/NET0131  ;
  assign n6543 = n952 & ~n6536 ;
  assign n6544 = ~n6542 & n6543 ;
  assign n6546 = \rEIP_reg[11]/NET0131  & ~n4650 ;
  assign n6547 = ~\rEIP_reg[11]/NET0131  & ~n4661 ;
  assign n6548 = ~n4662 & ~n6547 ;
  assign n6549 = n4684 & ~n6548 ;
  assign n6550 = ~\EBX_reg[11]/NET0131  & ~n4720 ;
  assign n6551 = n742 & ~n6550 ;
  assign n6552 = ~\EBX_reg[10]/NET0131  & n4697 ;
  assign n6553 = \EBX_reg[31]/NET0131  & ~n6552 ;
  assign n6555 = \EBX_reg[11]/NET0131  & ~n6553 ;
  assign n6554 = ~\EBX_reg[11]/NET0131  & n6553 ;
  assign n6556 = ~n4684 & ~n6554 ;
  assign n6557 = ~n6555 & n6556 ;
  assign n6558 = n736 & ~n6557 ;
  assign n6559 = ~n6551 & ~n6558 ;
  assign n6560 = ~n6549 & ~n6559 ;
  assign n6561 = n833 & n6551 ;
  assign n6562 = ~n6560 & ~n6561 ;
  assign n6563 = n825 & ~n6562 ;
  assign n6564 = ~n6546 & ~n6563 ;
  assign n6565 = n948 & ~n6564 ;
  assign n6545 = \rEIP_reg[11]/NET0131  & ~n6300 ;
  assign n6566 = \PhyAddrPointer_reg[11]/NET0131  & n981 ;
  assign n6567 = ~n1731 & ~n6566 ;
  assign n6568 = ~n6545 & n6567 ;
  assign n6569 = ~n6565 & n6568 ;
  assign n6570 = ~n6544 & n6569 ;
  assign n6572 = ~\PhyAddrPointer_reg[12]/NET0131  & ~n2372 ;
  assign n6573 = ~n2373 & ~n6572 ;
  assign n6574 = n2013 & n5890 ;
  assign n6575 = n2036 & ~n6574 ;
  assign n6577 = n6573 & ~n6575 ;
  assign n6576 = ~n6573 & n6575 ;
  assign n6578 = ~\DataWidth_reg[1]/NET0131  & ~n6576 ;
  assign n6579 = ~n6577 & n6578 ;
  assign n6571 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[12]/NET0131  ;
  assign n6580 = n952 & ~n6571 ;
  assign n6581 = ~n6579 & n6580 ;
  assign n6583 = \rEIP_reg[12]/NET0131  & ~n4650 ;
  assign n6584 = ~\rEIP_reg[12]/NET0131  & ~n4662 ;
  assign n6585 = ~n4663 & ~n6584 ;
  assign n6586 = n4684 & ~n6585 ;
  assign n6587 = ~\EBX_reg[12]/NET0131  & ~n4720 ;
  assign n6588 = n742 & ~n6587 ;
  assign n6589 = ~\EBX_reg[11]/NET0131  & n6552 ;
  assign n6590 = \EBX_reg[31]/NET0131  & ~n6589 ;
  assign n6592 = ~\EBX_reg[12]/NET0131  & n6590 ;
  assign n6591 = \EBX_reg[12]/NET0131  & ~n6590 ;
  assign n6593 = ~n4684 & ~n6591 ;
  assign n6594 = ~n6592 & n6593 ;
  assign n6595 = n736 & ~n6594 ;
  assign n6596 = ~n6588 & ~n6595 ;
  assign n6597 = ~n6586 & ~n6596 ;
  assign n6598 = n833 & n6588 ;
  assign n6599 = ~n6597 & ~n6598 ;
  assign n6600 = n825 & ~n6599 ;
  assign n6601 = ~n6583 & ~n6600 ;
  assign n6602 = n948 & ~n6601 ;
  assign n6582 = \rEIP_reg[12]/NET0131  & ~n6300 ;
  assign n6603 = \PhyAddrPointer_reg[12]/NET0131  & n981 ;
  assign n6604 = ~n1731 & ~n6603 ;
  assign n6605 = ~n6582 & n6604 ;
  assign n6606 = ~n6602 & n6605 ;
  assign n6607 = ~n6581 & n6606 ;
  assign n6609 = ~\PhyAddrPointer_reg[13]/NET0131  & ~n2373 ;
  assign n6610 = ~n2374 & ~n6609 ;
  assign n6611 = n2373 & n5893 ;
  assign n6612 = n2036 & ~n6611 ;
  assign n6614 = ~n6610 & n6612 ;
  assign n6613 = n6610 & ~n6612 ;
  assign n6615 = ~\DataWidth_reg[1]/NET0131  & ~n6613 ;
  assign n6616 = ~n6614 & n6615 ;
  assign n6608 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[13]/NET0131  ;
  assign n6617 = n952 & ~n6608 ;
  assign n6618 = ~n6616 & n6617 ;
  assign n6620 = \rEIP_reg[13]/NET0131  & ~n4650 ;
  assign n6622 = ~\rEIP_reg[13]/NET0131  & ~n4663 ;
  assign n6623 = ~n4664 & ~n6622 ;
  assign n6624 = n4720 & ~n6623 ;
  assign n6621 = ~\EBX_reg[13]/NET0131  & ~n4720 ;
  assign n6625 = n742 & ~n6621 ;
  assign n6626 = ~n6624 & n6625 ;
  assign n6628 = \EBX_reg[31]/NET0131  & ~n4700 ;
  assign n6630 = \EBX_reg[13]/NET0131  & ~n6628 ;
  assign n6629 = ~\EBX_reg[13]/NET0131  & n6628 ;
  assign n6631 = ~n4684 & ~n6629 ;
  assign n6632 = ~n6630 & n6631 ;
  assign n6627 = n4684 & ~n6623 ;
  assign n6633 = n736 & ~n6627 ;
  assign n6634 = ~n6632 & n6633 ;
  assign n6635 = ~n6626 & ~n6634 ;
  assign n6636 = n825 & ~n6635 ;
  assign n6637 = ~n6620 & ~n6636 ;
  assign n6638 = n948 & ~n6637 ;
  assign n6619 = \rEIP_reg[13]/NET0131  & ~n6300 ;
  assign n6639 = \PhyAddrPointer_reg[13]/NET0131  & n981 ;
  assign n6640 = ~n1731 & ~n6639 ;
  assign n6641 = ~n6619 & n6640 ;
  assign n6642 = ~n6638 & n6641 ;
  assign n6643 = ~n6618 & n6642 ;
  assign n6645 = ~\PhyAddrPointer_reg[0]/NET0131  & n2374 ;
  assign n6646 = n2036 & ~n6645 ;
  assign n6648 = ~n2599 & n6646 ;
  assign n6647 = n2599 & ~n6646 ;
  assign n6649 = ~\DataWidth_reg[1]/NET0131  & ~n6647 ;
  assign n6650 = ~n6648 & n6649 ;
  assign n6644 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[14]/NET0131  ;
  assign n6651 = n952 & ~n6644 ;
  assign n6652 = ~n6650 & n6651 ;
  assign n6654 = \rEIP_reg[14]/NET0131  & ~n4650 ;
  assign n6656 = ~\rEIP_reg[14]/NET0131  & ~n4664 ;
  assign n6657 = ~n4665 & ~n6656 ;
  assign n6658 = n4720 & ~n6657 ;
  assign n6655 = ~\EBX_reg[14]/NET0131  & ~n4720 ;
  assign n6659 = n742 & ~n6655 ;
  assign n6660 = ~n6658 & n6659 ;
  assign n6662 = \EBX_reg[31]/NET0131  & ~n4701 ;
  assign n6664 = \EBX_reg[14]/NET0131  & ~n6662 ;
  assign n6663 = ~\EBX_reg[14]/NET0131  & n6662 ;
  assign n6665 = ~n4684 & ~n6663 ;
  assign n6666 = ~n6664 & n6665 ;
  assign n6661 = n4684 & ~n6657 ;
  assign n6667 = n736 & ~n6661 ;
  assign n6668 = ~n6666 & n6667 ;
  assign n6669 = ~n6660 & ~n6668 ;
  assign n6670 = n825 & ~n6669 ;
  assign n6671 = ~n6654 & ~n6670 ;
  assign n6672 = n948 & ~n6671 ;
  assign n6653 = \rEIP_reg[14]/NET0131  & ~n6300 ;
  assign n6673 = \PhyAddrPointer_reg[14]/NET0131  & n981 ;
  assign n6674 = ~n1731 & ~n6673 ;
  assign n6675 = ~n6653 & n6674 ;
  assign n6676 = ~n6672 & n6675 ;
  assign n6677 = ~n6652 & n6676 ;
  assign n6679 = \PhyAddrPointer_reg[14]/NET0131  & n6645 ;
  assign n6680 = n2036 & ~n6679 ;
  assign n6682 = ~n2378 & n6680 ;
  assign n6681 = n2378 & ~n6680 ;
  assign n6683 = ~\DataWidth_reg[1]/NET0131  & ~n6681 ;
  assign n6684 = ~n6682 & n6683 ;
  assign n6678 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[15]/NET0131  ;
  assign n6685 = n952 & ~n6678 ;
  assign n6686 = ~n6684 & n6685 ;
  assign n6688 = \rEIP_reg[15]/NET0131  & ~n4650 ;
  assign n6691 = ~\EBX_reg[15]/NET0131  & ~n4720 ;
  assign n6692 = n742 & ~n6691 ;
  assign n6696 = \EBX_reg[31]/NET0131  & ~n4702 ;
  assign n6698 = \EBX_reg[15]/NET0131  & ~n6696 ;
  assign n6697 = ~\EBX_reg[15]/NET0131  & n6696 ;
  assign n6699 = ~n4684 & ~n6697 ;
  assign n6700 = ~n6698 & n6699 ;
  assign n6701 = n736 & ~n6700 ;
  assign n6702 = ~n6692 & ~n6701 ;
  assign n6689 = ~\rEIP_reg[15]/NET0131  & ~n4665 ;
  assign n6690 = ~n4666 & ~n6689 ;
  assign n6693 = n833 & n6692 ;
  assign n6694 = n4684 & ~n6693 ;
  assign n6695 = ~n6690 & n6694 ;
  assign n6703 = n825 & ~n6695 ;
  assign n6704 = ~n6702 & n6703 ;
  assign n6705 = ~n6688 & ~n6704 ;
  assign n6706 = n948 & ~n6705 ;
  assign n6687 = \rEIP_reg[15]/NET0131  & ~n6300 ;
  assign n6707 = \PhyAddrPointer_reg[15]/NET0131  & n981 ;
  assign n6708 = ~n1731 & ~n6707 ;
  assign n6709 = ~n6687 & n6708 ;
  assign n6710 = ~n6706 & n6709 ;
  assign n6711 = ~n6686 & n6710 ;
  assign n6713 = n2759 & n5890 ;
  assign n6714 = n2036 & ~n6713 ;
  assign n6716 = n2787 & ~n6714 ;
  assign n6715 = ~n2787 & n6714 ;
  assign n6717 = ~\DataWidth_reg[1]/NET0131  & ~n6715 ;
  assign n6718 = ~n6716 & n6717 ;
  assign n6712 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[16]/NET0131  ;
  assign n6719 = n952 & ~n6712 ;
  assign n6720 = ~n6718 & n6719 ;
  assign n6722 = ~\rEIP_reg[16]/NET0131  & ~n4666 ;
  assign n6723 = ~n4667 & ~n6722 ;
  assign n6724 = n4684 & ~n6723 ;
  assign n6734 = ~n833 & n6724 ;
  assign n6733 = ~\EBX_reg[16]/NET0131  & ~n4720 ;
  assign n6735 = n3798 & ~n6733 ;
  assign n6736 = ~n6734 & n6735 ;
  assign n6725 = \EBX_reg[31]/NET0131  & ~n4703 ;
  assign n6727 = ~\EBX_reg[16]/NET0131  & n6725 ;
  assign n6726 = \EBX_reg[16]/NET0131  & ~n6725 ;
  assign n6728 = ~n4684 & ~n6726 ;
  assign n6729 = ~n6727 & n6728 ;
  assign n6730 = n1719 & ~n6724 ;
  assign n6731 = ~n6729 & n6730 ;
  assign n6732 = \rEIP_reg[16]/NET0131  & ~n4650 ;
  assign n6737 = ~n6731 & ~n6732 ;
  assign n6738 = ~n6736 & n6737 ;
  assign n6739 = n948 & ~n6738 ;
  assign n6721 = \rEIP_reg[16]/NET0131  & ~n6300 ;
  assign n6740 = \PhyAddrPointer_reg[16]/NET0131  & n981 ;
  assign n6741 = ~n1731 & ~n6740 ;
  assign n6742 = ~n6721 & n6741 ;
  assign n6743 = ~n6739 & n6742 ;
  assign n6744 = ~n6720 & n6743 ;
  assign n6746 = n2786 & n5893 ;
  assign n6747 = n2036 & ~n6746 ;
  assign n6749 = ~n2802 & n6747 ;
  assign n6748 = n2802 & ~n6747 ;
  assign n6750 = ~\DataWidth_reg[1]/NET0131  & ~n6748 ;
  assign n6751 = ~n6749 & n6750 ;
  assign n6745 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[17]/NET0131  ;
  assign n6752 = n952 & ~n6745 ;
  assign n6753 = ~n6751 & n6752 ;
  assign n6757 = ~\rEIP_reg[17]/NET0131  & ~n4667 ;
  assign n6756 = \rEIP_reg[17]/NET0131  & n4667 ;
  assign n6758 = n4684 & ~n6756 ;
  assign n6759 = ~n6757 & n6758 ;
  assign n6768 = \EBX_reg[17]/NET0131  & ~n4684 ;
  assign n6769 = ~n6759 & ~n6768 ;
  assign n6770 = n895 & ~n6769 ;
  assign n6767 = \rEIP_reg[17]/NET0131  & ~n825 ;
  assign n6771 = \EBX_reg[17]/NET0131  & n5975 ;
  assign n6772 = ~n6767 & ~n6771 ;
  assign n6773 = ~n6770 & n6772 ;
  assign n6774 = n742 & ~n6773 ;
  assign n6755 = \rEIP_reg[17]/NET0131  & n5988 ;
  assign n6760 = \EBX_reg[31]/NET0131  & ~n4704 ;
  assign n6762 = \EBX_reg[17]/NET0131  & n6760 ;
  assign n6761 = ~\EBX_reg[17]/NET0131  & ~n6760 ;
  assign n6763 = ~n4684 & ~n6761 ;
  assign n6764 = ~n6762 & n6763 ;
  assign n6765 = ~n6759 & ~n6764 ;
  assign n6766 = n1719 & ~n6765 ;
  assign n6775 = ~n6755 & ~n6766 ;
  assign n6776 = ~n6774 & n6775 ;
  assign n6777 = n948 & ~n6776 ;
  assign n6754 = \rEIP_reg[17]/NET0131  & ~n6300 ;
  assign n6778 = \PhyAddrPointer_reg[17]/NET0131  & n981 ;
  assign n6779 = ~n1731 & ~n6778 ;
  assign n6780 = ~n6754 & n6779 ;
  assign n6781 = ~n6777 & n6780 ;
  assign n6782 = ~n6753 & n6781 ;
  assign n6784 = n2036 & ~n4632 ;
  assign n6786 = ~n2852 & n6784 ;
  assign n6785 = n2852 & ~n6784 ;
  assign n6787 = ~\DataWidth_reg[1]/NET0131  & ~n6785 ;
  assign n6788 = ~n6786 & n6787 ;
  assign n6783 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[18]/NET0131  ;
  assign n6789 = n952 & ~n6783 ;
  assign n6790 = ~n6788 & n6789 ;
  assign n6801 = \EBX_reg[31]/NET0131  & ~n4705 ;
  assign n6803 = ~\EBX_reg[18]/NET0131  & n6801 ;
  assign n6802 = \EBX_reg[18]/NET0131  & ~n6801 ;
  assign n6804 = ~n4684 & ~n6802 ;
  assign n6805 = ~n6803 & n6804 ;
  assign n6794 = ~\rEIP_reg[18]/NET0131  & ~n6756 ;
  assign n6795 = \rEIP_reg[18]/NET0131  & n6756 ;
  assign n6796 = ~n6794 & ~n6795 ;
  assign n6800 = n4684 & ~n6796 ;
  assign n6806 = n1719 & ~n6800 ;
  assign n6807 = ~n6805 & n6806 ;
  assign n6792 = \rEIP_reg[18]/NET0131  & ~n4650 ;
  assign n6797 = n4720 & ~n6796 ;
  assign n6793 = ~\EBX_reg[18]/NET0131  & ~n4720 ;
  assign n6798 = n3798 & ~n6793 ;
  assign n6799 = ~n6797 & n6798 ;
  assign n6808 = ~n6792 & ~n6799 ;
  assign n6809 = ~n6807 & n6808 ;
  assign n6810 = n948 & ~n6809 ;
  assign n6791 = \rEIP_reg[18]/NET0131  & ~n6300 ;
  assign n6811 = \PhyAddrPointer_reg[18]/NET0131  & n981 ;
  assign n6812 = ~n1731 & ~n6811 ;
  assign n6813 = ~n6791 & n6812 ;
  assign n6814 = ~n6810 & n6813 ;
  assign n6815 = ~n6790 & n6814 ;
  assign n6817 = ~\PhyAddrPointer_reg[0]/NET0131  & n2620 ;
  assign n6818 = n2036 & ~n6817 ;
  assign n6820 = ~n2623 & n6818 ;
  assign n6819 = n2623 & ~n6818 ;
  assign n6821 = ~\DataWidth_reg[1]/NET0131  & ~n6819 ;
  assign n6822 = ~n6820 & n6821 ;
  assign n6816 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[19]/NET0131  ;
  assign n6823 = n952 & ~n6816 ;
  assign n6824 = ~n6822 & n6823 ;
  assign n6826 = ~\rEIP_reg[19]/NET0131  & ~n6795 ;
  assign n6827 = ~n5836 & ~n6826 ;
  assign n6828 = n4684 & ~n6827 ;
  assign n6838 = ~n833 & n6828 ;
  assign n6837 = ~\EBX_reg[19]/NET0131  & ~n4720 ;
  assign n6839 = n3798 & ~n6837 ;
  assign n6840 = ~n6838 & n6839 ;
  assign n6829 = \EBX_reg[31]/NET0131  & ~n4706 ;
  assign n6831 = ~\EBX_reg[19]/NET0131  & n6829 ;
  assign n6830 = \EBX_reg[19]/NET0131  & ~n6829 ;
  assign n6832 = ~n4684 & ~n6830 ;
  assign n6833 = ~n6831 & n6832 ;
  assign n6834 = n1719 & ~n6828 ;
  assign n6835 = ~n6833 & n6834 ;
  assign n6836 = \rEIP_reg[19]/NET0131  & ~n4650 ;
  assign n6841 = ~n6835 & ~n6836 ;
  assign n6842 = ~n6840 & n6841 ;
  assign n6843 = n948 & ~n6842 ;
  assign n6825 = \rEIP_reg[19]/NET0131  & ~n6300 ;
  assign n6844 = \PhyAddrPointer_reg[19]/NET0131  & n981 ;
  assign n6845 = ~n1731 & ~n6844 ;
  assign n6846 = ~n6825 & n6845 ;
  assign n6847 = ~n6843 & n6846 ;
  assign n6848 = ~n6824 & n6847 ;
  assign n6854 = ~READY_n_pad & ~n943 ;
  assign n6855 = ~n841 & n6854 ;
  assign n6856 = n4650 & n6855 ;
  assign n6853 = ~\RequestPending_reg/NET0131  & ~n4650 ;
  assign n6857 = n948 & ~n6853 ;
  assign n6858 = ~n6856 & n6857 ;
  assign n6849 = ~n982 & ~n1731 ;
  assign n6850 = n968 & n978 ;
  assign n6851 = n3114 & ~n6850 ;
  assign n6852 = \RequestPending_reg/NET0131  & ~n6851 ;
  assign n6859 = n6849 & ~n6852 ;
  assign n6860 = ~n6858 & n6859 ;
  assign n6862 = ~\EAX_reg[23]/NET0131  & ~n3606 ;
  assign n6863 = ~n3799 & ~n6862 ;
  assign n6864 = ~n833 & ~n6863 ;
  assign n6865 = n3798 & ~n6864 ;
  assign n6866 = n3806 & ~n6865 ;
  assign n6867 = \Datao[23]_pad  & ~n6866 ;
  assign n6868 = n742 & n6863 ;
  assign n6869 = n895 & n6868 ;
  assign n6870 = ~n6867 & ~n6869 ;
  assign n6871 = n948 & ~n6870 ;
  assign n6861 = \uWord_reg[7]/NET0131  & n956 ;
  assign n6872 = \Datao[23]_pad  & ~n3816 ;
  assign n6873 = ~n6861 & ~n6872 ;
  assign n6874 = ~n6871 & n6873 ;
  assign n6876 = ~\EAX_reg[19]/NET0131  & ~n3604 ;
  assign n6877 = ~n3605 & ~n6876 ;
  assign n6878 = ~n833 & ~n6877 ;
  assign n6879 = n3798 & ~n6878 ;
  assign n6880 = n3806 & ~n6879 ;
  assign n6881 = \Datao[19]_pad  & ~n6880 ;
  assign n6882 = n3798 & n6877 ;
  assign n6883 = ~n833 & n6882 ;
  assign n6884 = ~n6881 & ~n6883 ;
  assign n6885 = n948 & ~n6884 ;
  assign n6875 = \uWord_reg[3]/NET0131  & n956 ;
  assign n6886 = \Datao[19]_pad  & ~n3816 ;
  assign n6887 = ~n6875 & ~n6886 ;
  assign n6888 = ~n6885 & n6887 ;
  assign n6889 = \uWord_reg[3]/NET0131  & ~n3584 ;
  assign n6890 = READY_n_pad & \uWord_reg[3]/NET0131  ;
  assign n6891 = ~n4765 & ~n6890 ;
  assign n6892 = n736 & ~n6891 ;
  assign n6893 = \uWord_reg[3]/NET0131  & ~n3620 ;
  assign n6894 = ~n6882 & ~n6893 ;
  assign n6895 = ~n6892 & n6894 ;
  assign n6896 = n948 & ~n6895 ;
  assign n6897 = ~n6889 & ~n6896 ;
  assign n6898 = \uWord_reg[7]/NET0131  & ~n3841 ;
  assign n6899 = \Datai[7]_pad  & n736 ;
  assign n6900 = ~READY_n_pad & n6899 ;
  assign n6901 = ~n6868 & ~n6900 ;
  assign n6902 = n3843 & ~n6901 ;
  assign n6903 = ~n6898 & ~n6902 ;
  assign n6905 = n740 & n825 ;
  assign n6906 = \MemoryFetch_reg/NET0131  & ~n6905 ;
  assign n6907 = ~n3620 & ~n6906 ;
  assign n6908 = n948 & ~n6907 ;
  assign n6904 = \MemoryFetch_reg/NET0131  & ~n3583 ;
  assign n6909 = n3581 & ~n6904 ;
  assign n6910 = ~n6908 & n6909 ;
  assign n6912 = \ReadRequest_reg/NET0131  & ~n3804 ;
  assign n6913 = ~n864 & ~n6912 ;
  assign n6914 = n948 & ~n6913 ;
  assign n6911 = \ReadRequest_reg/NET0131  & ~n3583 ;
  assign n6915 = n3581 & ~n6911 ;
  assign n6916 = ~n6914 & n6915 ;
  assign n6917 = ~\EBX_reg[0]/NET0131  & n833 ;
  assign n6918 = n3798 & ~n6917 ;
  assign n6919 = ~n1719 & ~n6918 ;
  assign n6920 = ~\EBX_reg[0]/NET0131  & ~n4684 ;
  assign n6921 = ~n6919 & ~n6920 ;
  assign n6922 = n4650 & ~n6921 ;
  assign n6923 = \rEIP_reg[0]/NET0131  & ~n6922 ;
  assign n6924 = ~\InstQueueRd_Addr_reg[0]/NET0131  & n740 ;
  assign n6925 = n742 & n833 ;
  assign n6926 = ~n3619 & ~n4684 ;
  assign n6927 = ~n6925 & ~n6926 ;
  assign n6928 = \EBX_reg[0]/NET0131  & ~n6927 ;
  assign n6929 = ~n6924 & ~n6928 ;
  assign n6930 = n825 & ~n6929 ;
  assign n6931 = ~n6923 & ~n6930 ;
  assign n6932 = n948 & ~n6931 ;
  assign n6933 = ~n953 & ~n981 ;
  assign n6934 = \PhyAddrPointer_reg[0]/NET0131  & ~n6933 ;
  assign n6935 = n972 & n3664 ;
  assign n6936 = \rEIP_reg[0]/NET0131  & ~n6935 ;
  assign n6937 = ~n6934 & ~n6936 ;
  assign n6938 = ~n6932 & n6937 ;
  assign n6940 = \EAX_reg[29]/NET0131  & n3612 ;
  assign n6941 = \EAX_reg[30]/NET0131  & ~n6940 ;
  assign n6942 = ~\EAX_reg[30]/NET0131  & n6940 ;
  assign n6943 = ~n6941 & ~n6942 ;
  assign n6944 = ~n833 & n6943 ;
  assign n6945 = n3798 & ~n6944 ;
  assign n6946 = n3806 & ~n6945 ;
  assign n6947 = \Datao[30]_pad  & ~n6946 ;
  assign n6948 = n742 & ~n6943 ;
  assign n6949 = n895 & n6948 ;
  assign n6950 = ~n6947 & ~n6949 ;
  assign n6951 = n948 & ~n6950 ;
  assign n6939 = \uWord_reg[14]/NET0131  & n956 ;
  assign n6952 = \Datao[30]_pad  & ~n3816 ;
  assign n6953 = ~n6939 & ~n6952 ;
  assign n6954 = ~n6951 & n6953 ;
  assign n6959 = ~\EAX_reg[28]/NET0131  & ~n3145 ;
  assign n6960 = n3759 & ~n6959 ;
  assign n6961 = \EAX_reg[28]/NET0131  & ~n3447 ;
  assign n6955 = ~n3344 & n3375 ;
  assign n6956 = n808 & ~n3376 ;
  assign n6957 = ~n6955 & n6956 ;
  assign n6958 = n755 & n6957 ;
  assign n6962 = \Datai[28]_pad  & n835 ;
  assign n6963 = ~n3615 & ~n6962 ;
  assign n6964 = n826 & ~n6963 ;
  assign n6965 = ~n6958 & ~n6964 ;
  assign n6966 = ~n6961 & n6965 ;
  assign n6967 = ~n6960 & n6966 ;
  assign n6968 = n948 & ~n6967 ;
  assign n6969 = \EAX_reg[28]/NET0131  & ~n3116 ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = \uWord_reg[14]/NET0131  & ~n3584 ;
  assign n6972 = \Datai[14]_pad  & n736 ;
  assign n6973 = ~READY_n_pad & n6972 ;
  assign n6974 = ~n6948 & ~n6973 ;
  assign n6975 = n825 & ~n6974 ;
  assign n6976 = \uWord_reg[14]/NET0131  & ~n3621 ;
  assign n6977 = ~n6975 & ~n6976 ;
  assign n6978 = n948 & ~n6977 ;
  assign n6979 = ~n6971 & ~n6978 ;
  assign n6980 = \EAX_reg[0]/NET0131  & ~n4743 ;
  assign n6981 = \Datai[0]_pad  & n865 ;
  assign n6982 = ~n1294 & n3153 ;
  assign n6983 = ~\EAX_reg[0]/NET0131  & n3118 ;
  assign n6984 = ~n6982 & ~n6983 ;
  assign n6985 = ~n6981 & n6984 ;
  assign n6986 = n948 & ~n6985 ;
  assign n6987 = ~n6980 & ~n6986 ;
  assign n6991 = \EBX_reg[27]/NET0131  & n3787 ;
  assign n6992 = ~\EBX_reg[28]/NET0131  & ~n6991 ;
  assign n6990 = n3787 & n3851 ;
  assign n6993 = n773 & ~n6990 ;
  assign n6994 = ~n6992 & n6993 ;
  assign n6988 = \EBX_reg[28]/NET0131  & n3486 ;
  assign n6989 = n752 & n6957 ;
  assign n6995 = ~n6988 & ~n6989 ;
  assign n6996 = ~n6994 & n6995 ;
  assign n6997 = n948 & ~n6996 ;
  assign n6998 = \EBX_reg[28]/NET0131  & ~n3116 ;
  assign n6999 = ~n6997 & ~n6998 ;
  assign n7039 = \EAX_reg[16]/NET0131  & ~n3447 ;
  assign n7032 = ~\EAX_reg[16]/NET0131  & ~n3133 ;
  assign n7033 = n3118 & ~n3134 ;
  assign n7034 = ~n7032 & n7033 ;
  assign n7004 = \InstQueue_reg[12][0]/NET0131  & n469 ;
  assign n7005 = \InstQueue_reg[1][0]/NET0131  & n454 ;
  assign n7018 = ~n7004 & ~n7005 ;
  assign n7006 = \InstQueue_reg[15][0]/NET0131  & n488 ;
  assign n7007 = \InstQueue_reg[13][0]/NET0131  & n490 ;
  assign n7019 = ~n7006 & ~n7007 ;
  assign n7026 = n7018 & n7019 ;
  assign n7000 = \InstQueue_reg[6][0]/NET0131  & n480 ;
  assign n7001 = \InstQueue_reg[2][0]/NET0131  & n476 ;
  assign n7016 = ~n7000 & ~n7001 ;
  assign n7002 = \InstQueue_reg[5][0]/NET0131  & n478 ;
  assign n7003 = \InstQueue_reg[7][0]/NET0131  & n463 ;
  assign n7017 = ~n7002 & ~n7003 ;
  assign n7027 = n7016 & n7017 ;
  assign n7028 = n7026 & n7027 ;
  assign n7012 = \InstQueue_reg[9][0]/NET0131  & n457 ;
  assign n7013 = \InstQueue_reg[11][0]/NET0131  & n486 ;
  assign n7022 = ~n7012 & ~n7013 ;
  assign n7014 = \InstQueue_reg[3][0]/NET0131  & n461 ;
  assign n7015 = \InstQueue_reg[10][0]/NET0131  & n482 ;
  assign n7023 = ~n7014 & ~n7015 ;
  assign n7024 = n7022 & n7023 ;
  assign n7008 = \InstQueue_reg[0][0]/NET0131  & n471 ;
  assign n7009 = \InstQueue_reg[8][0]/NET0131  & n484 ;
  assign n7020 = ~n7008 & ~n7009 ;
  assign n7010 = \InstQueue_reg[14][0]/NET0131  & n474 ;
  assign n7011 = \InstQueue_reg[4][0]/NET0131  & n466 ;
  assign n7021 = ~n7010 & ~n7011 ;
  assign n7025 = n7020 & n7021 ;
  assign n7029 = n7024 & n7025 ;
  assign n7030 = n7028 & n7029 ;
  assign n7031 = n3153 & ~n7030 ;
  assign n7035 = \Datai[16]_pad  & n835 ;
  assign n7036 = \Datai[0]_pad  & n736 ;
  assign n7037 = ~n7035 & ~n7036 ;
  assign n7038 = n826 & ~n7037 ;
  assign n7040 = ~n7031 & ~n7038 ;
  assign n7041 = ~n7034 & n7040 ;
  assign n7042 = ~n7039 & n7041 ;
  assign n7043 = n948 & ~n7042 ;
  assign n7044 = \EAX_reg[16]/NET0131  & ~n3116 ;
  assign n7045 = ~n7043 & ~n7044 ;
  assign n7078 = ~\EAX_reg[17]/NET0131  & ~n3134 ;
  assign n7079 = n3118 & ~n3135 ;
  assign n7080 = ~n7078 & n7079 ;
  assign n7085 = \EAX_reg[17]/NET0131  & ~n3447 ;
  assign n7050 = \InstQueue_reg[12][1]/NET0131  & n469 ;
  assign n7051 = \InstQueue_reg[1][1]/NET0131  & n454 ;
  assign n7064 = ~n7050 & ~n7051 ;
  assign n7052 = \InstQueue_reg[15][1]/NET0131  & n488 ;
  assign n7053 = \InstQueue_reg[8][1]/NET0131  & n484 ;
  assign n7065 = ~n7052 & ~n7053 ;
  assign n7072 = n7064 & n7065 ;
  assign n7046 = \InstQueue_reg[6][1]/NET0131  & n480 ;
  assign n7047 = \InstQueue_reg[2][1]/NET0131  & n476 ;
  assign n7062 = ~n7046 & ~n7047 ;
  assign n7048 = \InstQueue_reg[5][1]/NET0131  & n478 ;
  assign n7049 = \InstQueue_reg[7][1]/NET0131  & n463 ;
  assign n7063 = ~n7048 & ~n7049 ;
  assign n7073 = n7062 & n7063 ;
  assign n7074 = n7072 & n7073 ;
  assign n7058 = \InstQueue_reg[9][1]/NET0131  & n457 ;
  assign n7059 = \InstQueue_reg[11][1]/NET0131  & n486 ;
  assign n7068 = ~n7058 & ~n7059 ;
  assign n7060 = \InstQueue_reg[13][1]/NET0131  & n490 ;
  assign n7061 = \InstQueue_reg[10][1]/NET0131  & n482 ;
  assign n7069 = ~n7060 & ~n7061 ;
  assign n7070 = n7068 & n7069 ;
  assign n7054 = \InstQueue_reg[0][1]/NET0131  & n471 ;
  assign n7055 = \InstQueue_reg[3][1]/NET0131  & n461 ;
  assign n7066 = ~n7054 & ~n7055 ;
  assign n7056 = \InstQueue_reg[14][1]/NET0131  & n474 ;
  assign n7057 = \InstQueue_reg[4][1]/NET0131  & n466 ;
  assign n7067 = ~n7056 & ~n7057 ;
  assign n7071 = n7066 & n7067 ;
  assign n7075 = n7070 & n7071 ;
  assign n7076 = n7074 & n7075 ;
  assign n7077 = n3153 & ~n7076 ;
  assign n7081 = \Datai[17]_pad  & n835 ;
  assign n7082 = \Datai[1]_pad  & n736 ;
  assign n7083 = ~n7081 & ~n7082 ;
  assign n7084 = n826 & ~n7083 ;
  assign n7086 = ~n7077 & ~n7084 ;
  assign n7087 = ~n7085 & n7086 ;
  assign n7088 = ~n7080 & n7087 ;
  assign n7089 = n948 & ~n7088 ;
  assign n7090 = \EAX_reg[17]/NET0131  & ~n3116 ;
  assign n7091 = ~n7089 & ~n7090 ;
  assign n7092 = \EAX_reg[18]/NET0131  & ~n3116 ;
  assign n7125 = ~n3445 & ~n7079 ;
  assign n7126 = \EAX_reg[18]/NET0131  & ~n7125 ;
  assign n7133 = ~\EAX_reg[18]/NET0131  & n3118 ;
  assign n7134 = n3135 & n7133 ;
  assign n7127 = \EAX_reg[18]/NET0131  & ~n826 ;
  assign n7130 = \Datai[18]_pad  & n826 ;
  assign n7131 = ~n7127 & ~n7130 ;
  assign n7132 = n835 & ~n7131 ;
  assign n7097 = \InstQueue_reg[9][2]/NET0131  & n457 ;
  assign n7098 = \InstQueue_reg[0][2]/NET0131  & n471 ;
  assign n7111 = ~n7097 & ~n7098 ;
  assign n7099 = \InstQueue_reg[11][2]/NET0131  & n486 ;
  assign n7100 = \InstQueue_reg[13][2]/NET0131  & n490 ;
  assign n7112 = ~n7099 & ~n7100 ;
  assign n7119 = n7111 & n7112 ;
  assign n7093 = \InstQueue_reg[3][2]/NET0131  & n461 ;
  assign n7094 = \InstQueue_reg[15][2]/NET0131  & n488 ;
  assign n7109 = ~n7093 & ~n7094 ;
  assign n7095 = \InstQueue_reg[10][2]/NET0131  & n482 ;
  assign n7096 = \InstQueue_reg[2][2]/NET0131  & n476 ;
  assign n7110 = ~n7095 & ~n7096 ;
  assign n7120 = n7109 & n7110 ;
  assign n7121 = n7119 & n7120 ;
  assign n7105 = \InstQueue_reg[12][2]/NET0131  & n469 ;
  assign n7106 = \InstQueue_reg[5][2]/NET0131  & n478 ;
  assign n7115 = ~n7105 & ~n7106 ;
  assign n7107 = \InstQueue_reg[4][2]/NET0131  & n466 ;
  assign n7108 = \InstQueue_reg[8][2]/NET0131  & n484 ;
  assign n7116 = ~n7107 & ~n7108 ;
  assign n7117 = n7115 & n7116 ;
  assign n7101 = \InstQueue_reg[6][2]/NET0131  & n480 ;
  assign n7102 = \InstQueue_reg[1][2]/NET0131  & n454 ;
  assign n7113 = ~n7101 & ~n7102 ;
  assign n7103 = \InstQueue_reg[7][2]/NET0131  & n463 ;
  assign n7104 = \InstQueue_reg[14][2]/NET0131  & n474 ;
  assign n7114 = ~n7103 & ~n7104 ;
  assign n7118 = n7113 & n7114 ;
  assign n7122 = n7117 & n7118 ;
  assign n7123 = n7121 & n7122 ;
  assign n7124 = n3153 & ~n7123 ;
  assign n7128 = ~n4746 & ~n7127 ;
  assign n7129 = n736 & ~n7128 ;
  assign n7135 = ~n7124 & ~n7129 ;
  assign n7136 = ~n7132 & n7135 ;
  assign n7137 = ~n7134 & n7136 ;
  assign n7138 = ~n7126 & n7137 ;
  assign n7139 = n948 & ~n7138 ;
  assign n7140 = ~n7092 & ~n7139 ;
  assign n7173 = ~\EAX_reg[19]/NET0131  & ~n3136 ;
  assign n7174 = n3118 & ~n3137 ;
  assign n7175 = ~n7173 & n7174 ;
  assign n7180 = \EAX_reg[19]/NET0131  & ~n3447 ;
  assign n7145 = \InstQueue_reg[6][3]/NET0131  & n480 ;
  assign n7146 = \InstQueue_reg[1][3]/NET0131  & n454 ;
  assign n7159 = ~n7145 & ~n7146 ;
  assign n7147 = \InstQueue_reg[0][3]/NET0131  & n471 ;
  assign n7148 = \InstQueue_reg[3][3]/NET0131  & n461 ;
  assign n7160 = ~n7147 & ~n7148 ;
  assign n7167 = n7159 & n7160 ;
  assign n7141 = \InstQueue_reg[8][3]/NET0131  & n484 ;
  assign n7142 = \InstQueue_reg[2][3]/NET0131  & n476 ;
  assign n7157 = ~n7141 & ~n7142 ;
  assign n7143 = \InstQueue_reg[11][3]/NET0131  & n486 ;
  assign n7144 = \InstQueue_reg[4][3]/NET0131  & n466 ;
  assign n7158 = ~n7143 & ~n7144 ;
  assign n7168 = n7157 & n7158 ;
  assign n7169 = n7167 & n7168 ;
  assign n7153 = \InstQueue_reg[15][3]/NET0131  & n488 ;
  assign n7154 = \InstQueue_reg[12][3]/NET0131  & n469 ;
  assign n7163 = ~n7153 & ~n7154 ;
  assign n7155 = \InstQueue_reg[5][3]/NET0131  & n478 ;
  assign n7156 = \InstQueue_reg[10][3]/NET0131  & n482 ;
  assign n7164 = ~n7155 & ~n7156 ;
  assign n7165 = n7163 & n7164 ;
  assign n7149 = \InstQueue_reg[9][3]/NET0131  & n457 ;
  assign n7150 = \InstQueue_reg[14][3]/NET0131  & n474 ;
  assign n7161 = ~n7149 & ~n7150 ;
  assign n7151 = \InstQueue_reg[7][3]/NET0131  & n463 ;
  assign n7152 = \InstQueue_reg[13][3]/NET0131  & n490 ;
  assign n7162 = ~n7151 & ~n7152 ;
  assign n7166 = n7161 & n7162 ;
  assign n7170 = n7165 & n7166 ;
  assign n7171 = n7169 & n7170 ;
  assign n7172 = n3153 & ~n7171 ;
  assign n7176 = \Datai[19]_pad  & n835 ;
  assign n7177 = \Datai[3]_pad  & n736 ;
  assign n7178 = ~n7176 & ~n7177 ;
  assign n7179 = n826 & ~n7178 ;
  assign n7181 = ~n7172 & ~n7179 ;
  assign n7182 = ~n7180 & n7181 ;
  assign n7183 = ~n7175 & n7182 ;
  assign n7184 = n948 & ~n7183 ;
  assign n7185 = \EAX_reg[19]/NET0131  & ~n3116 ;
  assign n7186 = ~n7184 & ~n7185 ;
  assign n7187 = ~n926 & n948 ;
  assign n7188 = \More_reg/NET0131  & ~n3116 ;
  assign n7189 = ~n7187 & ~n7188 ;
  assign n7223 = ~\EAX_reg[20]/NET0131  & ~n3137 ;
  assign n7222 = \EAX_reg[20]/NET0131  & n3137 ;
  assign n7224 = n3118 & ~n7222 ;
  assign n7225 = ~n7223 & n7224 ;
  assign n7229 = \EAX_reg[20]/NET0131  & ~n3447 ;
  assign n7194 = \InstQueue_reg[6][4]/NET0131  & n480 ;
  assign n7195 = \InstQueue_reg[1][4]/NET0131  & n454 ;
  assign n7208 = ~n7194 & ~n7195 ;
  assign n7196 = \InstQueue_reg[15][4]/NET0131  & n488 ;
  assign n7197 = \InstQueue_reg[3][4]/NET0131  & n461 ;
  assign n7209 = ~n7196 & ~n7197 ;
  assign n7216 = n7208 & n7209 ;
  assign n7190 = \InstQueue_reg[8][4]/NET0131  & n484 ;
  assign n7191 = \InstQueue_reg[2][4]/NET0131  & n476 ;
  assign n7206 = ~n7190 & ~n7191 ;
  assign n7192 = \InstQueue_reg[11][4]/NET0131  & n486 ;
  assign n7193 = \InstQueue_reg[7][4]/NET0131  & n463 ;
  assign n7207 = ~n7192 & ~n7193 ;
  assign n7217 = n7206 & n7207 ;
  assign n7218 = n7216 & n7217 ;
  assign n7202 = \InstQueue_reg[9][4]/NET0131  & n457 ;
  assign n7203 = \InstQueue_reg[12][4]/NET0131  & n469 ;
  assign n7212 = ~n7202 & ~n7203 ;
  assign n7204 = \InstQueue_reg[5][4]/NET0131  & n478 ;
  assign n7205 = \InstQueue_reg[10][4]/NET0131  & n482 ;
  assign n7213 = ~n7204 & ~n7205 ;
  assign n7214 = n7212 & n7213 ;
  assign n7198 = \InstQueue_reg[0][4]/NET0131  & n471 ;
  assign n7199 = \InstQueue_reg[14][4]/NET0131  & n474 ;
  assign n7210 = ~n7198 & ~n7199 ;
  assign n7200 = \InstQueue_reg[4][4]/NET0131  & n466 ;
  assign n7201 = \InstQueue_reg[13][4]/NET0131  & n490 ;
  assign n7211 = ~n7200 & ~n7201 ;
  assign n7215 = n7210 & n7211 ;
  assign n7219 = n7214 & n7215 ;
  assign n7220 = n7218 & n7219 ;
  assign n7221 = n3153 & ~n7220 ;
  assign n7226 = \Datai[20]_pad  & n835 ;
  assign n7227 = ~n4294 & ~n7226 ;
  assign n7228 = n826 & ~n7227 ;
  assign n7230 = ~n7221 & ~n7228 ;
  assign n7231 = ~n7229 & n7230 ;
  assign n7232 = ~n7225 & n7231 ;
  assign n7233 = n948 & ~n7232 ;
  assign n7234 = \EAX_reg[20]/NET0131  & ~n3116 ;
  assign n7235 = ~n7233 & ~n7234 ;
  assign n7268 = ~\EAX_reg[21]/NET0131  & ~n7222 ;
  assign n7269 = \EAX_reg[21]/NET0131  & n7222 ;
  assign n7270 = n3118 & ~n7269 ;
  assign n7271 = ~n7268 & n7270 ;
  assign n7272 = \EAX_reg[21]/NET0131  & ~n3447 ;
  assign n7240 = \InstQueue_reg[0][5]/NET0131  & n471 ;
  assign n7241 = \InstQueue_reg[1][5]/NET0131  & n454 ;
  assign n7254 = ~n7240 & ~n7241 ;
  assign n7242 = \InstQueue_reg[6][5]/NET0131  & n480 ;
  assign n7243 = \InstQueue_reg[3][5]/NET0131  & n461 ;
  assign n7255 = ~n7242 & ~n7243 ;
  assign n7262 = n7254 & n7255 ;
  assign n7236 = \InstQueue_reg[8][5]/NET0131  & n484 ;
  assign n7237 = \InstQueue_reg[2][5]/NET0131  & n476 ;
  assign n7252 = ~n7236 & ~n7237 ;
  assign n7238 = \InstQueue_reg[10][5]/NET0131  & n482 ;
  assign n7239 = \InstQueue_reg[7][5]/NET0131  & n463 ;
  assign n7253 = ~n7238 & ~n7239 ;
  assign n7263 = n7252 & n7253 ;
  assign n7264 = n7262 & n7263 ;
  assign n7248 = \InstQueue_reg[13][5]/NET0131  & n490 ;
  assign n7249 = \InstQueue_reg[5][5]/NET0131  & n478 ;
  assign n7258 = ~n7248 & ~n7249 ;
  assign n7250 = \InstQueue_reg[11][5]/NET0131  & n486 ;
  assign n7251 = \InstQueue_reg[15][5]/NET0131  & n488 ;
  assign n7259 = ~n7250 & ~n7251 ;
  assign n7260 = n7258 & n7259 ;
  assign n7244 = \InstQueue_reg[4][5]/NET0131  & n466 ;
  assign n7245 = \InstQueue_reg[14][5]/NET0131  & n474 ;
  assign n7256 = ~n7244 & ~n7245 ;
  assign n7246 = \InstQueue_reg[9][5]/NET0131  & n457 ;
  assign n7247 = \InstQueue_reg[12][5]/NET0131  & n469 ;
  assign n7257 = ~n7246 & ~n7247 ;
  assign n7261 = n7256 & n7257 ;
  assign n7265 = n7260 & n7261 ;
  assign n7266 = n7264 & n7265 ;
  assign n7267 = n3153 & ~n7266 ;
  assign n7273 = \Datai[5]_pad  & n736 ;
  assign n7274 = \Datai[21]_pad  & n835 ;
  assign n7275 = ~n7273 & ~n7274 ;
  assign n7276 = n826 & ~n7275 ;
  assign n7277 = ~n7267 & ~n7276 ;
  assign n7278 = ~n7272 & n7277 ;
  assign n7279 = ~n7271 & n7278 ;
  assign n7280 = n948 & ~n7279 ;
  assign n7281 = \EAX_reg[21]/NET0131  & ~n3116 ;
  assign n7282 = ~n7280 & ~n7281 ;
  assign n7283 = \EAX_reg[22]/NET0131  & ~n3116 ;
  assign n7316 = n3447 & ~n7270 ;
  assign n7317 = \EAX_reg[22]/NET0131  & ~n7316 ;
  assign n7322 = ~\EAX_reg[22]/NET0131  & n3118 ;
  assign n7323 = n7269 & n7322 ;
  assign n7288 = \InstQueue_reg[5][6]/NET0131  & n478 ;
  assign n7289 = \InstQueue_reg[6][6]/NET0131  & n480 ;
  assign n7302 = ~n7288 & ~n7289 ;
  assign n7290 = \InstQueue_reg[12][6]/NET0131  & n469 ;
  assign n7291 = \InstQueue_reg[13][6]/NET0131  & n490 ;
  assign n7303 = ~n7290 & ~n7291 ;
  assign n7310 = n7302 & n7303 ;
  assign n7284 = \InstQueue_reg[14][6]/NET0131  & n474 ;
  assign n7285 = \InstQueue_reg[15][6]/NET0131  & n488 ;
  assign n7300 = ~n7284 & ~n7285 ;
  assign n7286 = \InstQueue_reg[10][6]/NET0131  & n482 ;
  assign n7287 = \InstQueue_reg[2][6]/NET0131  & n476 ;
  assign n7301 = ~n7286 & ~n7287 ;
  assign n7311 = n7300 & n7301 ;
  assign n7312 = n7310 & n7311 ;
  assign n7296 = \InstQueue_reg[0][6]/NET0131  & n471 ;
  assign n7297 = \InstQueue_reg[11][6]/NET0131  & n486 ;
  assign n7306 = ~n7296 & ~n7297 ;
  assign n7298 = \InstQueue_reg[8][6]/NET0131  & n484 ;
  assign n7299 = \InstQueue_reg[3][6]/NET0131  & n461 ;
  assign n7307 = ~n7298 & ~n7299 ;
  assign n7308 = n7306 & n7307 ;
  assign n7292 = \InstQueue_reg[9][6]/NET0131  & n457 ;
  assign n7293 = \InstQueue_reg[1][6]/NET0131  & n454 ;
  assign n7304 = ~n7292 & ~n7293 ;
  assign n7294 = \InstQueue_reg[4][6]/NET0131  & n466 ;
  assign n7295 = \InstQueue_reg[7][6]/NET0131  & n463 ;
  assign n7305 = ~n7294 & ~n7295 ;
  assign n7309 = n7304 & n7305 ;
  assign n7313 = n7308 & n7309 ;
  assign n7314 = n7312 & n7313 ;
  assign n7315 = n3153 & ~n7314 ;
  assign n7318 = \Datai[6]_pad  & n736 ;
  assign n7319 = \Datai[22]_pad  & n835 ;
  assign n7320 = ~n7318 & ~n7319 ;
  assign n7321 = n826 & ~n7320 ;
  assign n7324 = ~n7315 & ~n7321 ;
  assign n7325 = ~n7323 & n7324 ;
  assign n7326 = ~n7317 & n7325 ;
  assign n7327 = n948 & ~n7326 ;
  assign n7328 = ~n7283 & ~n7327 ;
  assign n7332 = ~\EAX_reg[23]/NET0131  & ~n3140 ;
  assign n7333 = n3118 & ~n4304 ;
  assign n7334 = ~n7332 & n7333 ;
  assign n7335 = \EAX_reg[23]/NET0131  & ~n3447 ;
  assign n7329 = n3184 & n3215 ;
  assign n7330 = ~n3216 & ~n7329 ;
  assign n7331 = n3153 & n7330 ;
  assign n7336 = \Datai[23]_pad  & n835 ;
  assign n7337 = ~n6899 & ~n7336 ;
  assign n7338 = n826 & ~n7337 ;
  assign n7339 = ~n7331 & ~n7338 ;
  assign n7340 = ~n7335 & n7339 ;
  assign n7341 = ~n7334 & n7340 ;
  assign n7342 = n948 & ~n7341 ;
  assign n7343 = \EAX_reg[23]/NET0131  & ~n3116 ;
  assign n7344 = ~n7342 & ~n7343 ;
  assign n7345 = \EAX_reg[24]/NET0131  & ~n3116 ;
  assign n7346 = n3447 & ~n7333 ;
  assign n7347 = \EAX_reg[24]/NET0131  & ~n7346 ;
  assign n7348 = ~\EAX_reg[24]/NET0131  & n3118 ;
  assign n7349 = n4304 & n7348 ;
  assign n7350 = ~n3216 & n3247 ;
  assign n7351 = ~n3248 & ~n7350 ;
  assign n7352 = n3153 & n7351 ;
  assign n7353 = \Datai[24]_pad  & n835 ;
  assign n7354 = ~n3844 & ~n7353 ;
  assign n7355 = n826 & ~n7354 ;
  assign n7356 = ~n7352 & ~n7355 ;
  assign n7357 = ~n7349 & n7356 ;
  assign n7358 = ~n7347 & n7357 ;
  assign n7359 = n948 & ~n7358 ;
  assign n7360 = ~n7345 & ~n7359 ;
  assign n7362 = \Datao[26]_pad  & ~n4286 ;
  assign n7363 = ~\EAX_reg[26]/NET0131  & ~n3608 ;
  assign n7364 = n742 & ~n3609 ;
  assign n7365 = ~n7363 & n7364 ;
  assign n7366 = n895 & n7365 ;
  assign n7367 = ~n7362 & ~n7366 ;
  assign n7368 = n948 & ~n7367 ;
  assign n7361 = \uWord_reg[10]/NET0131  & n956 ;
  assign n7369 = \Datao[26]_pad  & ~n3816 ;
  assign n7370 = ~n7361 & ~n7369 ;
  assign n7371 = ~n7368 & n7370 ;
  assign n7372 = \uWord_reg[0]/NET0131  & ~n3841 ;
  assign n7373 = ~\EAX_reg[16]/NET0131  & ~n3601 ;
  assign n7374 = ~n3602 & ~n7373 ;
  assign n7375 = n3798 & n7374 ;
  assign n7376 = n826 & n7036 ;
  assign n7377 = ~n7375 & ~n7376 ;
  assign n7378 = n948 & ~n7377 ;
  assign n7379 = ~n7372 & ~n7378 ;
  assign n7380 = \uWord_reg[10]/NET0131  & ~n3841 ;
  assign n7381 = n736 & n3563 ;
  assign n7382 = ~n7365 & ~n7381 ;
  assign n7383 = n3843 & ~n7382 ;
  assign n7384 = ~n7380 & ~n7383 ;
  assign n7385 = \uWord_reg[13]/NET0131  & ~n3584 ;
  assign n7386 = ~\EAX_reg[29]/NET0131  & ~n3612 ;
  assign n7387 = n3798 & ~n6940 ;
  assign n7388 = ~n7386 & n7387 ;
  assign n7389 = \uWord_reg[13]/NET0131  & ~n3621 ;
  assign n7390 = ~n3768 & ~n7389 ;
  assign n7391 = ~n7388 & n7390 ;
  assign n7392 = n948 & ~n7391 ;
  assign n7393 = ~n7385 & ~n7392 ;
  assign n7394 = \uWord_reg[1]/NET0131  & ~n3584 ;
  assign n7396 = READY_n_pad & \uWord_reg[1]/NET0131  ;
  assign n7397 = ~n5167 & ~n7396 ;
  assign n7398 = n736 & ~n7397 ;
  assign n7395 = \uWord_reg[1]/NET0131  & ~n3620 ;
  assign n7399 = ~\EAX_reg[17]/NET0131  & ~n3602 ;
  assign n7400 = ~n3603 & ~n7399 ;
  assign n7401 = n3798 & n7400 ;
  assign n7402 = ~n7395 & ~n7401 ;
  assign n7403 = ~n7398 & n7402 ;
  assign n7404 = n948 & ~n7403 ;
  assign n7405 = ~n7394 & ~n7404 ;
  assign n7406 = \uWord_reg[2]/NET0131  & ~n3841 ;
  assign n7407 = n736 & n4746 ;
  assign n7408 = ~\EAX_reg[18]/NET0131  & ~n3603 ;
  assign n7409 = ~n3604 & ~n7408 ;
  assign n7410 = n3798 & n7409 ;
  assign n7411 = ~n7407 & ~n7410 ;
  assign n7412 = n948 & ~n7411 ;
  assign n7413 = ~n7406 & ~n7412 ;
  assign n7414 = \uWord_reg[5]/NET0131  & ~n3841 ;
  assign n7415 = ~READY_n_pad & n7273 ;
  assign n7417 = ~\EAX_reg[21]/NET0131  & ~n4282 ;
  assign n7416 = n3138 & n3605 ;
  assign n7418 = n742 & ~n7416 ;
  assign n7419 = ~n7417 & n7418 ;
  assign n7420 = ~n7415 & ~n7419 ;
  assign n7421 = n3843 & ~n7420 ;
  assign n7422 = ~n7414 & ~n7421 ;
  assign n7423 = \uWord_reg[6]/NET0131  & ~n3841 ;
  assign n7424 = ~READY_n_pad & n7318 ;
  assign n7425 = ~\EAX_reg[22]/NET0131  & ~n7416 ;
  assign n7426 = n742 & ~n3606 ;
  assign n7427 = ~n7425 & n7426 ;
  assign n7428 = ~n7424 & ~n7427 ;
  assign n7429 = n3843 & ~n7428 ;
  assign n7430 = ~n7423 & ~n7429 ;
  assign n7431 = \uWord_reg[9]/NET0131  & ~n3841 ;
  assign n7432 = n826 & n4311 ;
  assign n7433 = ~\EAX_reg[25]/NET0131  & ~n3607 ;
  assign n7434 = ~n3608 & n3798 ;
  assign n7435 = ~n7433 & n7434 ;
  assign n7436 = ~n7432 & ~n7435 ;
  assign n7437 = n948 & ~n7436 ;
  assign n7438 = ~n7431 & ~n7437 ;
  assign n7439 = n948 & n3486 ;
  assign n7440 = n3116 & ~n7439 ;
  assign n7441 = \EBX_reg[0]/NET0131  & ~n7440 ;
  assign n7442 = ~\EBX_reg[0]/NET0131  & n773 ;
  assign n7443 = ~n1294 & n3454 ;
  assign n7444 = ~n7442 & ~n7443 ;
  assign n7445 = n948 & ~n7444 ;
  assign n7446 = ~n7441 & ~n7445 ;
  assign n7448 = \EBX_reg[10]/NET0131  & n3486 ;
  assign n7447 = n3454 & ~n4979 ;
  assign n7449 = ~\EBX_reg[10]/NET0131  & ~n3468 ;
  assign n7450 = n773 & ~n3469 ;
  assign n7451 = ~n7449 & n7450 ;
  assign n7452 = ~n7447 & ~n7451 ;
  assign n7453 = ~n7448 & n7452 ;
  assign n7454 = n948 & ~n7453 ;
  assign n7455 = \EBX_reg[10]/NET0131  & ~n3116 ;
  assign n7456 = ~n7454 & ~n7455 ;
  assign n7458 = ~n3486 & ~n7450 ;
  assign n7459 = \EBX_reg[11]/NET0131  & ~n7458 ;
  assign n7457 = n3454 & ~n4930 ;
  assign n7460 = ~\EBX_reg[11]/NET0131  & n773 ;
  assign n7461 = n3469 & n7460 ;
  assign n7462 = ~n7457 & ~n7461 ;
  assign n7463 = ~n7459 & n7462 ;
  assign n7464 = n948 & ~n7463 ;
  assign n7465 = \EBX_reg[11]/NET0131  & ~n3116 ;
  assign n7466 = ~n7464 & ~n7465 ;
  assign n7469 = ~\EBX_reg[12]/NET0131  & ~n3470 ;
  assign n7470 = n773 & ~n3471 ;
  assign n7471 = ~n7469 & n7470 ;
  assign n7467 = n3454 & ~n5025 ;
  assign n7468 = \EBX_reg[12]/NET0131  & n3486 ;
  assign n7472 = ~n7467 & ~n7468 ;
  assign n7473 = ~n7471 & n7472 ;
  assign n7474 = n948 & ~n7473 ;
  assign n7475 = \EBX_reg[12]/NET0131  & ~n3116 ;
  assign n7476 = ~n7474 & ~n7475 ;
  assign n7477 = \EBX_reg[14]/NET0131  & ~n3116 ;
  assign n7479 = n773 & ~n3472 ;
  assign n7480 = ~n3486 & ~n7479 ;
  assign n7481 = \EBX_reg[14]/NET0131  & ~n7480 ;
  assign n7478 = n3454 & ~n5112 ;
  assign n7482 = ~\EBX_reg[14]/NET0131  & n773 ;
  assign n7483 = n3472 & n7482 ;
  assign n7484 = ~n7478 & ~n7483 ;
  assign n7485 = ~n7481 & n7484 ;
  assign n7486 = n948 & ~n7485 ;
  assign n7487 = ~n7477 & ~n7486 ;
  assign n7489 = ~\EBX_reg[13]/NET0131  & ~n3471 ;
  assign n7490 = n7479 & ~n7489 ;
  assign n7488 = \EBX_reg[13]/NET0131  & n3486 ;
  assign n7491 = n3454 & ~n5067 ;
  assign n7492 = ~n7488 & ~n7491 ;
  assign n7493 = ~n7490 & n7492 ;
  assign n7494 = n948 & ~n7493 ;
  assign n7495 = \EBX_reg[13]/NET0131  & ~n3116 ;
  assign n7496 = ~n7494 & ~n7495 ;
  assign n7499 = ~\EBX_reg[15]/NET0131  & ~n3473 ;
  assign n7500 = n773 & ~n3474 ;
  assign n7501 = ~n7499 & n7500 ;
  assign n7497 = \EBX_reg[15]/NET0131  & n3486 ;
  assign n7498 = n3454 & ~n5156 ;
  assign n7502 = ~n7497 & ~n7498 ;
  assign n7503 = ~n7501 & n7502 ;
  assign n7504 = n948 & ~n7503 ;
  assign n7505 = \EBX_reg[15]/NET0131  & ~n3116 ;
  assign n7506 = ~n7504 & ~n7505 ;
  assign n7509 = ~\EBX_reg[16]/NET0131  & ~n3474 ;
  assign n7510 = n773 & ~n3475 ;
  assign n7511 = ~n7509 & n7510 ;
  assign n7507 = \EBX_reg[16]/NET0131  & n3486 ;
  assign n7508 = n3454 & ~n7030 ;
  assign n7512 = ~n7507 & ~n7508 ;
  assign n7513 = ~n7511 & n7512 ;
  assign n7514 = n948 & ~n7513 ;
  assign n7515 = \EBX_reg[16]/NET0131  & ~n3116 ;
  assign n7516 = ~n7514 & ~n7515 ;
  assign n7519 = ~\EBX_reg[17]/NET0131  & ~n3475 ;
  assign n7520 = n773 & ~n3476 ;
  assign n7521 = ~n7519 & n7520 ;
  assign n7517 = \EBX_reg[17]/NET0131  & n3486 ;
  assign n7518 = n3454 & ~n7076 ;
  assign n7522 = ~n7517 & ~n7518 ;
  assign n7523 = ~n7521 & n7522 ;
  assign n7524 = n948 & ~n7523 ;
  assign n7525 = \EBX_reg[17]/NET0131  & ~n3116 ;
  assign n7526 = ~n7524 & ~n7525 ;
  assign n7529 = ~\EBX_reg[18]/NET0131  & ~n3476 ;
  assign n7530 = n773 & ~n3781 ;
  assign n7531 = ~n7529 & n7530 ;
  assign n7527 = \EBX_reg[18]/NET0131  & n3486 ;
  assign n7528 = n3454 & ~n7123 ;
  assign n7532 = ~n7527 & ~n7528 ;
  assign n7533 = ~n7531 & n7532 ;
  assign n7534 = n948 & ~n7533 ;
  assign n7535 = \EBX_reg[18]/NET0131  & ~n3116 ;
  assign n7536 = ~n7534 & ~n7535 ;
  assign n7539 = ~\EBX_reg[19]/NET0131  & ~n3781 ;
  assign n7540 = n773 & ~n3782 ;
  assign n7541 = ~n7539 & n7540 ;
  assign n7537 = \EBX_reg[19]/NET0131  & n3486 ;
  assign n7538 = n3454 & ~n7171 ;
  assign n7542 = ~n7537 & ~n7538 ;
  assign n7543 = ~n7541 & n7542 ;
  assign n7544 = n948 & ~n7543 ;
  assign n7545 = \EBX_reg[19]/NET0131  & ~n3116 ;
  assign n7546 = ~n7544 & ~n7545 ;
  assign n7548 = \EBX_reg[1]/NET0131  & n3486 ;
  assign n7547 = ~n1261 & n3454 ;
  assign n7549 = n773 & n5807 ;
  assign n7550 = ~n7547 & ~n7549 ;
  assign n7551 = ~n7548 & n7550 ;
  assign n7552 = n948 & ~n7551 ;
  assign n7553 = \EBX_reg[1]/NET0131  & ~n3116 ;
  assign n7554 = ~n7552 & ~n7553 ;
  assign n7557 = ~\EBX_reg[20]/NET0131  & ~n3782 ;
  assign n7558 = n773 & ~n3479 ;
  assign n7559 = ~n7557 & n7558 ;
  assign n7555 = \EBX_reg[20]/NET0131  & n3486 ;
  assign n7556 = n3454 & ~n7220 ;
  assign n7560 = ~n7555 & ~n7556 ;
  assign n7561 = ~n7559 & n7560 ;
  assign n7562 = n948 & ~n7561 ;
  assign n7563 = \EBX_reg[20]/NET0131  & ~n3116 ;
  assign n7564 = ~n7562 & ~n7563 ;
  assign n7568 = \EBX_reg[21]/NET0131  & n3479 ;
  assign n7567 = ~\EBX_reg[21]/NET0131  & ~n3479 ;
  assign n7569 = n773 & ~n7567 ;
  assign n7570 = ~n7568 & n7569 ;
  assign n7565 = \EBX_reg[21]/NET0131  & n3486 ;
  assign n7566 = n3454 & ~n7266 ;
  assign n7571 = ~n7565 & ~n7566 ;
  assign n7572 = ~n7570 & n7571 ;
  assign n7573 = n948 & ~n7572 ;
  assign n7574 = \EBX_reg[21]/NET0131  & ~n3116 ;
  assign n7575 = ~n7573 & ~n7574 ;
  assign n7578 = ~\EBX_reg[22]/NET0131  & ~n7568 ;
  assign n7579 = n773 & ~n3480 ;
  assign n7580 = ~n7578 & n7579 ;
  assign n7576 = \EBX_reg[22]/NET0131  & n3486 ;
  assign n7577 = n3454 & ~n7314 ;
  assign n7581 = ~n7576 & ~n7577 ;
  assign n7582 = ~n7580 & n7581 ;
  assign n7583 = n948 & ~n7582 ;
  assign n7584 = \EBX_reg[22]/NET0131  & ~n3116 ;
  assign n7585 = ~n7583 & ~n7584 ;
  assign n7588 = ~\EBX_reg[23]/NET0131  & ~n3480 ;
  assign n7589 = n773 & ~n3481 ;
  assign n7590 = ~n7588 & n7589 ;
  assign n7586 = n3454 & n7330 ;
  assign n7587 = \EBX_reg[23]/NET0131  & n3486 ;
  assign n7591 = ~n7586 & ~n7587 ;
  assign n7592 = ~n7590 & n7591 ;
  assign n7593 = n948 & ~n7592 ;
  assign n7594 = \EBX_reg[23]/NET0131  & ~n3116 ;
  assign n7595 = ~n7593 & ~n7594 ;
  assign n7598 = ~\EBX_reg[24]/NET0131  & ~n3785 ;
  assign n7599 = n773 & ~n3786 ;
  assign n7600 = ~n7598 & n7599 ;
  assign n7596 = \EBX_reg[24]/NET0131  & n3486 ;
  assign n7597 = n3454 & n7351 ;
  assign n7601 = ~n7596 & ~n7597 ;
  assign n7602 = ~n7600 & n7601 ;
  assign n7603 = n948 & ~n7602 ;
  assign n7604 = \EBX_reg[24]/NET0131  & ~n3116 ;
  assign n7605 = ~n7603 & ~n7604 ;
  assign n7607 = \EBX_reg[2]/NET0131  & n3486 ;
  assign n7606 = ~n1225 & n3454 ;
  assign n7608 = ~\EBX_reg[2]/NET0131  & ~n3460 ;
  assign n7609 = ~n3461 & ~n7608 ;
  assign n7610 = n773 & n7609 ;
  assign n7611 = ~n7606 & ~n7610 ;
  assign n7612 = ~n7607 & n7611 ;
  assign n7613 = n948 & ~n7612 ;
  assign n7614 = \EBX_reg[2]/NET0131  & ~n3116 ;
  assign n7615 = ~n7613 & ~n7614 ;
  assign n7617 = \EBX_reg[3]/NET0131  & n3486 ;
  assign n7616 = ~n1189 & n3454 ;
  assign n7618 = ~\EBX_reg[3]/NET0131  & ~n3461 ;
  assign n7619 = ~n3462 & ~n7618 ;
  assign n7620 = n773 & n7619 ;
  assign n7621 = ~n7616 & ~n7620 ;
  assign n7622 = ~n7617 & n7621 ;
  assign n7623 = n948 & ~n7622 ;
  assign n7624 = \EBX_reg[3]/NET0131  & ~n3116 ;
  assign n7625 = ~n7623 & ~n7624 ;
  assign n7627 = \EBX_reg[4]/NET0131  & n3486 ;
  assign n7626 = ~n1156 & n3454 ;
  assign n7628 = ~\EBX_reg[4]/NET0131  & ~n3462 ;
  assign n7629 = ~n3463 & ~n7628 ;
  assign n7630 = n773 & n7629 ;
  assign n7631 = ~n7626 & ~n7630 ;
  assign n7632 = ~n7627 & n7631 ;
  assign n7633 = n948 & ~n7632 ;
  assign n7634 = \EBX_reg[4]/NET0131  & ~n3116 ;
  assign n7635 = ~n7633 & ~n7634 ;
  assign n7637 = \EBX_reg[5]/NET0131  & n3486 ;
  assign n7636 = ~n1120 & n3454 ;
  assign n7638 = ~\EBX_reg[5]/NET0131  & ~n3463 ;
  assign n7639 = ~n3464 & ~n7638 ;
  assign n7640 = n773 & n7639 ;
  assign n7641 = ~n7636 & ~n7640 ;
  assign n7642 = ~n7637 & n7641 ;
  assign n7643 = n948 & ~n7642 ;
  assign n7644 = \EBX_reg[5]/NET0131  & ~n3116 ;
  assign n7645 = ~n7643 & ~n7644 ;
  assign n7647 = \EBX_reg[6]/NET0131  & n3486 ;
  assign n7646 = ~n1086 & n3454 ;
  assign n7648 = ~\EBX_reg[6]/NET0131  & ~n3464 ;
  assign n7649 = ~n3465 & ~n7648 ;
  assign n7650 = n773 & n7649 ;
  assign n7651 = ~n7646 & ~n7650 ;
  assign n7652 = ~n7647 & n7651 ;
  assign n7653 = n948 & ~n7652 ;
  assign n7654 = \EBX_reg[6]/NET0131  & ~n3116 ;
  assign n7655 = ~n7653 & ~n7654 ;
  assign n7657 = \EBX_reg[7]/NET0131  & n3486 ;
  assign n7656 = ~n1051 & n3454 ;
  assign n7658 = ~\EBX_reg[7]/NET0131  & ~n3465 ;
  assign n7659 = ~n3466 & ~n7658 ;
  assign n7660 = n773 & n7659 ;
  assign n7661 = ~n7656 & ~n7660 ;
  assign n7662 = ~n7657 & n7661 ;
  assign n7663 = n948 & ~n7662 ;
  assign n7664 = \EBX_reg[7]/NET0131  & ~n3116 ;
  assign n7665 = ~n7663 & ~n7664 ;
  assign n7667 = \EBX_reg[8]/NET0131  & n3486 ;
  assign n7666 = n3454 & ~n4887 ;
  assign n7668 = ~\EBX_reg[8]/NET0131  & ~n3466 ;
  assign n7669 = ~n3467 & ~n7668 ;
  assign n7670 = n773 & n7669 ;
  assign n7671 = ~n7666 & ~n7670 ;
  assign n7672 = ~n7667 & n7671 ;
  assign n7673 = n948 & ~n7672 ;
  assign n7674 = \EBX_reg[8]/NET0131  & ~n3116 ;
  assign n7675 = ~n7673 & ~n7674 ;
  assign n7677 = \EBX_reg[9]/NET0131  & n3486 ;
  assign n7676 = n3454 & ~n4846 ;
  assign n7678 = ~\EBX_reg[9]/NET0131  & ~n3467 ;
  assign n7679 = ~n3468 & ~n7678 ;
  assign n7680 = n773 & n7679 ;
  assign n7681 = ~n7676 & ~n7680 ;
  assign n7682 = ~n7677 & n7681 ;
  assign n7683 = n948 & ~n7682 ;
  assign n7684 = \EBX_reg[9]/NET0131  & ~n3116 ;
  assign n7685 = ~n7683 & ~n7684 ;
  assign n7686 = ~n936 & n948 ;
  assign n7687 = \Flush_reg/NET0131  & ~n3116 ;
  assign n7688 = ~n7686 & ~n7687 ;
  assign n7694 = ~\Datai[26]_pad  & ~n3902 ;
  assign n7695 = ~n3903 & ~n7694 ;
  assign n7696 = n3876 & n7695 ;
  assign n7697 = ~\Datai[18]_pad  & ~n3911 ;
  assign n7698 = ~n3912 & ~n7697 ;
  assign n7699 = n3919 & n7698 ;
  assign n7700 = ~n7696 & ~n7699 ;
  assign n7701 = \DataWidth_reg[1]/NET0131  & ~n7700 ;
  assign n7689 = \Datai[2]_pad  & ~n3868 ;
  assign n7690 = \InstQueue_reg[0][2]/NET0131  & ~n3864 ;
  assign n7691 = ~n3867 & n7690 ;
  assign n7692 = ~n7689 & ~n7691 ;
  assign n7702 = ~n3924 & ~n7692 ;
  assign n7703 = ~n7701 & ~n7702 ;
  assign n7704 = n952 & ~n7703 ;
  assign n7705 = ~n569 & n3864 ;
  assign n7706 = ~n7690 & ~n7705 ;
  assign n7707 = n993 & ~n7706 ;
  assign n7693 = n970 & ~n7692 ;
  assign n7708 = \InstQueue_reg[0][2]/NET0131  & ~n3933 ;
  assign n7709 = ~n7693 & ~n7708 ;
  assign n7710 = ~n7707 & n7709 ;
  assign n7711 = ~n7704 & n7710 ;
  assign n7717 = n3948 & n7695 ;
  assign n7718 = n3950 & n7698 ;
  assign n7719 = ~n7717 & ~n7718 ;
  assign n7720 = \DataWidth_reg[1]/NET0131  & ~n7719 ;
  assign n7712 = \Datai[2]_pad  & ~n3942 ;
  assign n7713 = \InstQueue_reg[10][2]/NET0131  & ~n3939 ;
  assign n7714 = ~n3941 & n7713 ;
  assign n7715 = ~n7712 & ~n7714 ;
  assign n7721 = ~n3955 & ~n7715 ;
  assign n7722 = ~n7720 & ~n7721 ;
  assign n7723 = n952 & ~n7722 ;
  assign n7724 = ~n569 & n3939 ;
  assign n7725 = ~n7713 & ~n7724 ;
  assign n7726 = n993 & ~n7725 ;
  assign n7716 = n970 & ~n7715 ;
  assign n7727 = \InstQueue_reg[10][2]/NET0131  & ~n3933 ;
  assign n7728 = ~n7716 & ~n7727 ;
  assign n7729 = ~n7726 & n7728 ;
  assign n7730 = ~n7723 & n7729 ;
  assign n7736 = n3950 & n7695 ;
  assign n7737 = n3941 & n7698 ;
  assign n7738 = ~n7736 & ~n7737 ;
  assign n7739 = \DataWidth_reg[1]/NET0131  & ~n7738 ;
  assign n7731 = \Datai[2]_pad  & ~n3968 ;
  assign n7732 = \InstQueue_reg[11][2]/NET0131  & ~n3967 ;
  assign n7733 = ~n3939 & n7732 ;
  assign n7734 = ~n7731 & ~n7733 ;
  assign n7740 = ~n3979 & ~n7734 ;
  assign n7741 = ~n7739 & ~n7740 ;
  assign n7742 = n952 & ~n7741 ;
  assign n7743 = ~n569 & n3967 ;
  assign n7744 = ~n7732 & ~n7743 ;
  assign n7745 = n993 & ~n7744 ;
  assign n7735 = n970 & ~n7734 ;
  assign n7746 = \InstQueue_reg[11][2]/NET0131  & ~n3933 ;
  assign n7747 = ~n7735 & ~n7746 ;
  assign n7748 = ~n7745 & n7747 ;
  assign n7749 = ~n7742 & n7748 ;
  assign n7755 = n3941 & n7695 ;
  assign n7756 = n3939 & n7698 ;
  assign n7757 = ~n7755 & ~n7756 ;
  assign n7758 = \DataWidth_reg[1]/NET0131  & ~n7757 ;
  assign n7750 = \Datai[2]_pad  & ~n3992 ;
  assign n7751 = \InstQueue_reg[12][2]/NET0131  & ~n3991 ;
  assign n7752 = ~n3967 & n7751 ;
  assign n7753 = ~n7750 & ~n7752 ;
  assign n7759 = ~n4002 & ~n7753 ;
  assign n7760 = ~n7758 & ~n7759 ;
  assign n7761 = n952 & ~n7760 ;
  assign n7762 = ~n569 & n3991 ;
  assign n7763 = ~n7751 & ~n7762 ;
  assign n7764 = n993 & ~n7763 ;
  assign n7754 = n970 & ~n7753 ;
  assign n7765 = \InstQueue_reg[12][2]/NET0131  & ~n3933 ;
  assign n7766 = ~n7754 & ~n7765 ;
  assign n7767 = ~n7764 & n7766 ;
  assign n7768 = ~n7761 & n7767 ;
  assign n7774 = n3939 & n7695 ;
  assign n7775 = n3967 & n7698 ;
  assign n7776 = ~n7774 & ~n7775 ;
  assign n7777 = \DataWidth_reg[1]/NET0131  & ~n7776 ;
  assign n7769 = \Datai[2]_pad  & ~n4013 ;
  assign n7770 = \InstQueue_reg[13][2]/NET0131  & ~n3876 ;
  assign n7771 = ~n3991 & n7770 ;
  assign n7772 = ~n7769 & ~n7771 ;
  assign n7778 = ~n4023 & ~n7772 ;
  assign n7779 = ~n7777 & ~n7778 ;
  assign n7780 = n952 & ~n7779 ;
  assign n7781 = ~n569 & n3876 ;
  assign n7782 = ~n7770 & ~n7781 ;
  assign n7783 = n993 & ~n7782 ;
  assign n7773 = n970 & ~n7772 ;
  assign n7784 = \InstQueue_reg[13][2]/NET0131  & ~n3933 ;
  assign n7785 = ~n7773 & ~n7784 ;
  assign n7786 = ~n7783 & n7785 ;
  assign n7787 = ~n7780 & n7786 ;
  assign n7793 = n3967 & n7695 ;
  assign n7794 = n3991 & n7698 ;
  assign n7795 = ~n7793 & ~n7794 ;
  assign n7796 = \DataWidth_reg[1]/NET0131  & ~n7795 ;
  assign n7788 = \Datai[2]_pad  & ~n3923 ;
  assign n7789 = \InstQueue_reg[14][2]/NET0131  & ~n3919 ;
  assign n7790 = ~n3876 & n7789 ;
  assign n7791 = ~n7788 & ~n7790 ;
  assign n7797 = ~n4043 & ~n7791 ;
  assign n7798 = ~n7796 & ~n7797 ;
  assign n7799 = n952 & ~n7798 ;
  assign n7800 = ~n569 & n3919 ;
  assign n7801 = ~n7789 & ~n7800 ;
  assign n7802 = n993 & ~n7801 ;
  assign n7792 = n970 & ~n7791 ;
  assign n7803 = \InstQueue_reg[14][2]/NET0131  & ~n3933 ;
  assign n7804 = ~n7792 & ~n7803 ;
  assign n7805 = ~n7802 & n7804 ;
  assign n7806 = ~n7799 & n7805 ;
  assign n7812 = n3991 & n7695 ;
  assign n7813 = n3876 & n7698 ;
  assign n7814 = ~n7812 & ~n7813 ;
  assign n7815 = \DataWidth_reg[1]/NET0131  & ~n7814 ;
  assign n7807 = \Datai[2]_pad  & ~n4054 ;
  assign n7808 = \InstQueue_reg[15][2]/NET0131  & ~n3867 ;
  assign n7809 = ~n3919 & n7808 ;
  assign n7810 = ~n7807 & ~n7809 ;
  assign n7816 = ~n4064 & ~n7810 ;
  assign n7817 = ~n7815 & ~n7816 ;
  assign n7818 = n952 & ~n7817 ;
  assign n7819 = ~n569 & n3867 ;
  assign n7820 = ~n7808 & ~n7819 ;
  assign n7821 = n993 & ~n7820 ;
  assign n7811 = n970 & ~n7810 ;
  assign n7822 = \InstQueue_reg[15][2]/NET0131  & ~n3933 ;
  assign n7823 = ~n7811 & ~n7822 ;
  assign n7824 = ~n7821 & n7823 ;
  assign n7825 = ~n7818 & n7824 ;
  assign n7831 = n3919 & n7695 ;
  assign n7832 = n3867 & n7698 ;
  assign n7833 = ~n7831 & ~n7832 ;
  assign n7834 = \DataWidth_reg[1]/NET0131  & ~n7833 ;
  assign n7826 = \Datai[2]_pad  & ~n4076 ;
  assign n7827 = \InstQueue_reg[1][2]/NET0131  & ~n4075 ;
  assign n7828 = ~n3864 & n7827 ;
  assign n7829 = ~n7826 & ~n7828 ;
  assign n7835 = ~n4086 & ~n7829 ;
  assign n7836 = ~n7834 & ~n7835 ;
  assign n7837 = n952 & ~n7836 ;
  assign n7838 = ~n569 & n4075 ;
  assign n7839 = ~n7827 & ~n7838 ;
  assign n7840 = n993 & ~n7839 ;
  assign n7830 = n970 & ~n7829 ;
  assign n7841 = \InstQueue_reg[1][2]/NET0131  & ~n3933 ;
  assign n7842 = ~n7830 & ~n7841 ;
  assign n7843 = ~n7840 & n7842 ;
  assign n7844 = ~n7837 & n7843 ;
  assign n7850 = n3864 & n7698 ;
  assign n7851 = n3867 & n7695 ;
  assign n7852 = ~n7850 & ~n7851 ;
  assign n7853 = \DataWidth_reg[1]/NET0131  & ~n7852 ;
  assign n7845 = \Datai[2]_pad  & ~n4098 ;
  assign n7846 = \InstQueue_reg[2][2]/NET0131  & ~n4097 ;
  assign n7847 = ~n4075 & n7846 ;
  assign n7848 = ~n7845 & ~n7847 ;
  assign n7854 = ~n4108 & ~n7848 ;
  assign n7855 = ~n7853 & ~n7854 ;
  assign n7856 = n952 & ~n7855 ;
  assign n7857 = ~n569 & n4097 ;
  assign n7858 = ~n7846 & ~n7857 ;
  assign n7859 = n993 & ~n7858 ;
  assign n7849 = n970 & ~n7848 ;
  assign n7860 = \InstQueue_reg[2][2]/NET0131  & ~n3933 ;
  assign n7861 = ~n7849 & ~n7860 ;
  assign n7862 = ~n7859 & n7861 ;
  assign n7863 = ~n7856 & n7862 ;
  assign n7869 = n3864 & n7695 ;
  assign n7870 = n4075 & n7698 ;
  assign n7871 = ~n7869 & ~n7870 ;
  assign n7872 = \DataWidth_reg[1]/NET0131  & ~n7871 ;
  assign n7864 = \Datai[2]_pad  & ~n4120 ;
  assign n7865 = \InstQueue_reg[3][2]/NET0131  & ~n4119 ;
  assign n7866 = ~n4097 & n7865 ;
  assign n7867 = ~n7864 & ~n7866 ;
  assign n7873 = ~n4130 & ~n7867 ;
  assign n7874 = ~n7872 & ~n7873 ;
  assign n7875 = n952 & ~n7874 ;
  assign n7876 = ~n569 & n4119 ;
  assign n7877 = ~n7865 & ~n7876 ;
  assign n7878 = n993 & ~n7877 ;
  assign n7868 = n970 & ~n7867 ;
  assign n7879 = \InstQueue_reg[3][2]/NET0131  & ~n3933 ;
  assign n7880 = ~n7868 & ~n7879 ;
  assign n7881 = ~n7878 & n7880 ;
  assign n7882 = ~n7875 & n7881 ;
  assign n7888 = n4075 & n7695 ;
  assign n7889 = n4097 & n7698 ;
  assign n7890 = ~n7888 & ~n7889 ;
  assign n7891 = \DataWidth_reg[1]/NET0131  & ~n7890 ;
  assign n7883 = \Datai[2]_pad  & ~n4142 ;
  assign n7884 = \InstQueue_reg[4][2]/NET0131  & ~n4141 ;
  assign n7885 = ~n4119 & n7884 ;
  assign n7886 = ~n7883 & ~n7885 ;
  assign n7892 = ~n4152 & ~n7886 ;
  assign n7893 = ~n7891 & ~n7892 ;
  assign n7894 = n952 & ~n7893 ;
  assign n7895 = ~n569 & n4141 ;
  assign n7896 = ~n7884 & ~n7895 ;
  assign n7897 = n993 & ~n7896 ;
  assign n7887 = n970 & ~n7886 ;
  assign n7898 = \InstQueue_reg[4][2]/NET0131  & ~n3933 ;
  assign n7899 = ~n7887 & ~n7898 ;
  assign n7900 = ~n7897 & n7899 ;
  assign n7901 = ~n7894 & n7900 ;
  assign n7907 = n4097 & n7695 ;
  assign n7908 = n4119 & n7698 ;
  assign n7909 = ~n7907 & ~n7908 ;
  assign n7910 = \DataWidth_reg[1]/NET0131  & ~n7909 ;
  assign n7902 = \Datai[2]_pad  & ~n4164 ;
  assign n7903 = \InstQueue_reg[5][2]/NET0131  & ~n4163 ;
  assign n7904 = ~n4141 & n7903 ;
  assign n7905 = ~n7902 & ~n7904 ;
  assign n7911 = ~n4174 & ~n7905 ;
  assign n7912 = ~n7910 & ~n7911 ;
  assign n7913 = n952 & ~n7912 ;
  assign n7914 = ~n569 & n4163 ;
  assign n7915 = ~n7903 & ~n7914 ;
  assign n7916 = n993 & ~n7915 ;
  assign n7906 = n970 & ~n7905 ;
  assign n7917 = \InstQueue_reg[5][2]/NET0131  & ~n3933 ;
  assign n7918 = ~n7906 & ~n7917 ;
  assign n7919 = ~n7916 & n7918 ;
  assign n7920 = ~n7913 & n7919 ;
  assign n7926 = n4119 & n7695 ;
  assign n7927 = n4141 & n7698 ;
  assign n7928 = ~n7926 & ~n7927 ;
  assign n7929 = \DataWidth_reg[1]/NET0131  & ~n7928 ;
  assign n7921 = \Datai[2]_pad  & ~n4186 ;
  assign n7922 = \InstQueue_reg[6][2]/NET0131  & ~n4185 ;
  assign n7923 = ~n4163 & n7922 ;
  assign n7924 = ~n7921 & ~n7923 ;
  assign n7930 = ~n4196 & ~n7924 ;
  assign n7931 = ~n7929 & ~n7930 ;
  assign n7932 = n952 & ~n7931 ;
  assign n7933 = ~n569 & n4185 ;
  assign n7934 = ~n7922 & ~n7933 ;
  assign n7935 = n993 & ~n7934 ;
  assign n7925 = n970 & ~n7924 ;
  assign n7936 = \InstQueue_reg[6][2]/NET0131  & ~n3933 ;
  assign n7937 = ~n7925 & ~n7936 ;
  assign n7938 = ~n7935 & n7937 ;
  assign n7939 = ~n7932 & n7938 ;
  assign n7945 = n4141 & n7695 ;
  assign n7946 = n4163 & n7698 ;
  assign n7947 = ~n7945 & ~n7946 ;
  assign n7948 = \DataWidth_reg[1]/NET0131  & ~n7947 ;
  assign n7940 = \Datai[2]_pad  & ~n4207 ;
  assign n7941 = \InstQueue_reg[7][2]/NET0131  & ~n3948 ;
  assign n7942 = ~n4185 & n7941 ;
  assign n7943 = ~n7940 & ~n7942 ;
  assign n7949 = ~n4217 & ~n7943 ;
  assign n7950 = ~n7948 & ~n7949 ;
  assign n7951 = n952 & ~n7950 ;
  assign n7952 = ~n569 & n3948 ;
  assign n7953 = ~n7941 & ~n7952 ;
  assign n7954 = n993 & ~n7953 ;
  assign n7944 = n970 & ~n7943 ;
  assign n7955 = \InstQueue_reg[7][2]/NET0131  & ~n3933 ;
  assign n7956 = ~n7944 & ~n7955 ;
  assign n7957 = ~n7954 & n7956 ;
  assign n7958 = ~n7951 & n7957 ;
  assign n7964 = n4163 & n7695 ;
  assign n7965 = n4185 & n7698 ;
  assign n7966 = ~n7964 & ~n7965 ;
  assign n7967 = \DataWidth_reg[1]/NET0131  & ~n7966 ;
  assign n7959 = \Datai[2]_pad  & ~n3954 ;
  assign n7960 = \InstQueue_reg[8][2]/NET0131  & ~n3950 ;
  assign n7961 = ~n3948 & n7960 ;
  assign n7962 = ~n7959 & ~n7961 ;
  assign n7968 = ~n4237 & ~n7962 ;
  assign n7969 = ~n7967 & ~n7968 ;
  assign n7970 = n952 & ~n7969 ;
  assign n7971 = ~n569 & n3950 ;
  assign n7972 = ~n7960 & ~n7971 ;
  assign n7973 = n993 & ~n7972 ;
  assign n7963 = n970 & ~n7962 ;
  assign n7974 = \InstQueue_reg[8][2]/NET0131  & ~n3933 ;
  assign n7975 = ~n7963 & ~n7974 ;
  assign n7976 = ~n7973 & n7975 ;
  assign n7977 = ~n7970 & n7976 ;
  assign n7983 = n4185 & n7695 ;
  assign n7984 = n3948 & n7698 ;
  assign n7985 = ~n7983 & ~n7984 ;
  assign n7986 = \DataWidth_reg[1]/NET0131  & ~n7985 ;
  assign n7978 = \Datai[2]_pad  & ~n3978 ;
  assign n7979 = \InstQueue_reg[9][2]/NET0131  & ~n3941 ;
  assign n7980 = ~n3950 & n7979 ;
  assign n7981 = ~n7978 & ~n7980 ;
  assign n7987 = ~n4257 & ~n7981 ;
  assign n7988 = ~n7986 & ~n7987 ;
  assign n7989 = n952 & ~n7988 ;
  assign n7990 = ~n569 & n3941 ;
  assign n7991 = ~n7979 & ~n7990 ;
  assign n7992 = n993 & ~n7991 ;
  assign n7982 = n970 & ~n7981 ;
  assign n7993 = \InstQueue_reg[9][2]/NET0131  & ~n3933 ;
  assign n7994 = ~n7982 & ~n7993 ;
  assign n7995 = ~n7992 & n7994 ;
  assign n7996 = ~n7989 & n7995 ;
  assign n7998 = \Datao[29]_pad  & ~n4286 ;
  assign n7999 = ~n833 & n7388 ;
  assign n8000 = ~n7998 & ~n7999 ;
  assign n8001 = n948 & ~n8000 ;
  assign n7997 = \uWord_reg[13]/NET0131  & n956 ;
  assign n8002 = \Datao[29]_pad  & ~n3816 ;
  assign n8003 = ~n7997 & ~n8002 ;
  assign n8004 = ~n8001 & n8003 ;
  assign n8007 = \CodeFetch_reg/NET0131  & n948 ;
  assign n8008 = ~n4650 & n8007 ;
  assign n8005 = ~n960 & n1735 ;
  assign n8006 = \CodeFetch_reg/NET0131  & ~n8005 ;
  assign n8009 = ~n962 & ~n8006 ;
  assign n8010 = ~n8008 & n8009 ;
  assign n8012 = \Datao[18]_pad  & ~n4286 ;
  assign n8013 = ~n833 & n7410 ;
  assign n8014 = ~n8012 & ~n8013 ;
  assign n8015 = n948 & ~n8014 ;
  assign n8011 = \uWord_reg[2]/NET0131  & n956 ;
  assign n8016 = \Datao[18]_pad  & ~n3816 ;
  assign n8017 = ~n8011 & ~n8016 ;
  assign n8018 = ~n8015 & n8017 ;
  assign n8019 = \lWord_reg[0]/NET0131  & ~n3841 ;
  assign n8020 = \EAX_reg[0]/NET0131  & n3798 ;
  assign n8021 = ~n7376 & ~n8020 ;
  assign n8022 = n948 & ~n8021 ;
  assign n8023 = ~n8019 & ~n8022 ;
  assign n8024 = \lWord_reg[10]/NET0131  & ~n3841 ;
  assign n8025 = \EAX_reg[10]/NET0131  & n742 ;
  assign n8026 = ~n7381 & ~n8025 ;
  assign n8027 = n3843 & ~n8026 ;
  assign n8028 = ~n8024 & ~n8027 ;
  assign n8029 = \lWord_reg[11]/NET0131  & ~n3841 ;
  assign n8030 = \EAX_reg[11]/NET0131  & n3798 ;
  assign n8031 = ~n4758 & ~n8030 ;
  assign n8032 = n948 & ~n8031 ;
  assign n8033 = ~n8029 & ~n8032 ;
  assign n8034 = \lWord_reg[12]/NET0131  & ~n3841 ;
  assign n8035 = \EAX_reg[12]/NET0131  & n3798 ;
  assign n8036 = n826 & n3615 ;
  assign n8037 = ~n8035 & ~n8036 ;
  assign n8038 = n948 & ~n8037 ;
  assign n8039 = ~n8034 & ~n8038 ;
  assign n8040 = \lWord_reg[13]/NET0131  & ~n3841 ;
  assign n8041 = \EAX_reg[13]/NET0131  & n3798 ;
  assign n8042 = ~n3768 & ~n8041 ;
  assign n8043 = n948 & ~n8042 ;
  assign n8044 = ~n8040 & ~n8043 ;
  assign n8045 = \lWord_reg[14]/NET0131  & ~n3841 ;
  assign n8046 = \EAX_reg[14]/NET0131  & n3798 ;
  assign n8047 = n826 & n6972 ;
  assign n8048 = ~n8046 & ~n8047 ;
  assign n8049 = n948 & ~n8048 ;
  assign n8050 = ~n8045 & ~n8049 ;
  assign n8052 = \Datai[15]_pad  & n826 ;
  assign n8053 = READY_n_pad & \lWord_reg[15]/NET0131  ;
  assign n8054 = ~n8052 & ~n8053 ;
  assign n8055 = n736 & ~n8054 ;
  assign n8051 = \lWord_reg[15]/NET0131  & ~n3620 ;
  assign n8056 = \EAX_reg[15]/NET0131  & n3798 ;
  assign n8057 = ~n8051 & ~n8056 ;
  assign n8058 = ~n8055 & n8057 ;
  assign n8059 = n948 & ~n8058 ;
  assign n8060 = \lWord_reg[15]/NET0131  & ~n3584 ;
  assign n8061 = ~n8059 & ~n8060 ;
  assign n8062 = \lWord_reg[1]/NET0131  & ~n3841 ;
  assign n8063 = \EAX_reg[1]/NET0131  & n3798 ;
  assign n8064 = n736 & n5167 ;
  assign n8065 = ~n8063 & ~n8064 ;
  assign n8066 = n948 & ~n8065 ;
  assign n8067 = ~n8062 & ~n8066 ;
  assign n8068 = \lWord_reg[2]/NET0131  & ~n3841 ;
  assign n8069 = \EAX_reg[2]/NET0131  & n3798 ;
  assign n8070 = ~n7407 & ~n8069 ;
  assign n8071 = n948 & ~n8070 ;
  assign n8072 = ~n8068 & ~n8071 ;
  assign n8073 = \lWord_reg[3]/NET0131  & ~n3841 ;
  assign n8074 = \EAX_reg[3]/NET0131  & n3798 ;
  assign n8075 = n736 & n4765 ;
  assign n8076 = ~n8074 & ~n8075 ;
  assign n8077 = n948 & ~n8076 ;
  assign n8078 = ~n8073 & ~n8077 ;
  assign n8079 = \lWord_reg[4]/NET0131  & ~n3841 ;
  assign n8080 = \EAX_reg[4]/NET0131  & n3798 ;
  assign n8081 = ~n4295 & ~n8080 ;
  assign n8082 = n948 & ~n8081 ;
  assign n8083 = ~n8079 & ~n8082 ;
  assign n8084 = \lWord_reg[5]/NET0131  & ~n3841 ;
  assign n8085 = \EAX_reg[5]/NET0131  & n3798 ;
  assign n8086 = n826 & n7273 ;
  assign n8087 = ~n8085 & ~n8086 ;
  assign n8088 = n948 & ~n8087 ;
  assign n8089 = ~n8084 & ~n8088 ;
  assign n8090 = \lWord_reg[6]/NET0131  & ~n3841 ;
  assign n8091 = \EAX_reg[6]/NET0131  & n3798 ;
  assign n8092 = n826 & n7318 ;
  assign n8093 = ~n8091 & ~n8092 ;
  assign n8094 = n948 & ~n8093 ;
  assign n8095 = ~n8090 & ~n8094 ;
  assign n8096 = \lWord_reg[7]/NET0131  & ~n3841 ;
  assign n8097 = \EAX_reg[7]/NET0131  & n3798 ;
  assign n8098 = n826 & n6899 ;
  assign n8099 = ~n8097 & ~n8098 ;
  assign n8100 = n948 & ~n8099 ;
  assign n8101 = ~n8096 & ~n8100 ;
  assign n8102 = \lWord_reg[8]/NET0131  & ~n3841 ;
  assign n8103 = \EAX_reg[8]/NET0131  & n3798 ;
  assign n8104 = n826 & n3844 ;
  assign n8105 = ~n8103 & ~n8104 ;
  assign n8106 = n948 & ~n8105 ;
  assign n8107 = ~n8102 & ~n8106 ;
  assign n8108 = \lWord_reg[9]/NET0131  & ~n3841 ;
  assign n8109 = \EAX_reg[9]/NET0131  & n3798 ;
  assign n8110 = ~n7432 & ~n8109 ;
  assign n8111 = n948 & ~n8110 ;
  assign n8112 = ~n8108 & ~n8111 ;
  assign n8113 = \InstAddrPointer_reg[29]/NET0131  & ~n921 ;
  assign n8114 = ~n2465 & ~n8113 ;
  assign n8115 = n748 & ~n8114 ;
  assign n8119 = \InstAddrPointer_reg[29]/NET0131  & ~n2073 ;
  assign n8116 = ~n839 & n1368 ;
  assign n8117 = n809 & n1700 ;
  assign n8118 = ~n780 & ~n1574 ;
  assign n8120 = ~n8117 & ~n8118 ;
  assign n8121 = ~n8116 & n8120 ;
  assign n8122 = ~n8119 & n8121 ;
  assign n8123 = ~n2473 & n8122 ;
  assign n8124 = ~n8115 & n8123 ;
  assign n8125 = n948 & ~n8124 ;
  assign n8126 = \InstAddrPointer_reg[29]/NET0131  & ~n1736 ;
  assign n8127 = ~n2485 & ~n8126 ;
  assign n8128 = ~n8125 & n8127 ;
  assign n8134 = ~\Datai[29]_pad  & ~n3905 ;
  assign n8135 = ~n4324 & ~n8134 ;
  assign n8136 = n3876 & n8135 ;
  assign n8137 = ~\Datai[21]_pad  & ~n3915 ;
  assign n8138 = ~n4328 & ~n8137 ;
  assign n8139 = n3919 & n8138 ;
  assign n8140 = ~n8136 & ~n8139 ;
  assign n8141 = \DataWidth_reg[1]/NET0131  & ~n8140 ;
  assign n8129 = \Datai[5]_pad  & ~n3868 ;
  assign n8130 = \InstQueue_reg[0][5]/NET0131  & ~n3864 ;
  assign n8131 = ~n3867 & n8130 ;
  assign n8132 = ~n8129 & ~n8131 ;
  assign n8142 = ~n3924 & ~n8132 ;
  assign n8143 = ~n8141 & ~n8142 ;
  assign n8144 = n952 & ~n8143 ;
  assign n8145 = ~n697 & n3864 ;
  assign n8146 = ~n8130 & ~n8145 ;
  assign n8147 = n993 & ~n8146 ;
  assign n8133 = n970 & ~n8132 ;
  assign n8148 = \InstQueue_reg[0][5]/NET0131  & ~n3933 ;
  assign n8149 = ~n8133 & ~n8148 ;
  assign n8150 = ~n8147 & n8149 ;
  assign n8151 = ~n8144 & n8150 ;
  assign n8157 = n3948 & n8135 ;
  assign n8158 = n3950 & n8138 ;
  assign n8159 = ~n8157 & ~n8158 ;
  assign n8160 = \DataWidth_reg[1]/NET0131  & ~n8159 ;
  assign n8152 = \Datai[5]_pad  & ~n3942 ;
  assign n8153 = \InstQueue_reg[10][5]/NET0131  & ~n3939 ;
  assign n8154 = ~n3941 & n8153 ;
  assign n8155 = ~n8152 & ~n8154 ;
  assign n8161 = ~n3955 & ~n8155 ;
  assign n8162 = ~n8160 & ~n8161 ;
  assign n8163 = n952 & ~n8162 ;
  assign n8164 = ~n697 & n3939 ;
  assign n8165 = ~n8153 & ~n8164 ;
  assign n8166 = n993 & ~n8165 ;
  assign n8156 = n970 & ~n8155 ;
  assign n8167 = \InstQueue_reg[10][5]/NET0131  & ~n3933 ;
  assign n8168 = ~n8156 & ~n8167 ;
  assign n8169 = ~n8166 & n8168 ;
  assign n8170 = ~n8163 & n8169 ;
  assign n8176 = n3950 & n8135 ;
  assign n8177 = n3941 & n8138 ;
  assign n8178 = ~n8176 & ~n8177 ;
  assign n8179 = \DataWidth_reg[1]/NET0131  & ~n8178 ;
  assign n8171 = \Datai[5]_pad  & ~n3968 ;
  assign n8172 = \InstQueue_reg[11][5]/NET0131  & ~n3967 ;
  assign n8173 = ~n3939 & n8172 ;
  assign n8174 = ~n8171 & ~n8173 ;
  assign n8180 = ~n3979 & ~n8174 ;
  assign n8181 = ~n8179 & ~n8180 ;
  assign n8182 = n952 & ~n8181 ;
  assign n8183 = ~n697 & n3967 ;
  assign n8184 = ~n8172 & ~n8183 ;
  assign n8185 = n993 & ~n8184 ;
  assign n8175 = n970 & ~n8174 ;
  assign n8186 = \InstQueue_reg[11][5]/NET0131  & ~n3933 ;
  assign n8187 = ~n8175 & ~n8186 ;
  assign n8188 = ~n8185 & n8187 ;
  assign n8189 = ~n8182 & n8188 ;
  assign n8195 = n3941 & n8135 ;
  assign n8196 = n3939 & n8138 ;
  assign n8197 = ~n8195 & ~n8196 ;
  assign n8198 = \DataWidth_reg[1]/NET0131  & ~n8197 ;
  assign n8190 = \Datai[5]_pad  & ~n3992 ;
  assign n8191 = \InstQueue_reg[12][5]/NET0131  & ~n3991 ;
  assign n8192 = ~n3967 & n8191 ;
  assign n8193 = ~n8190 & ~n8192 ;
  assign n8199 = ~n4002 & ~n8193 ;
  assign n8200 = ~n8198 & ~n8199 ;
  assign n8201 = n952 & ~n8200 ;
  assign n8202 = ~n697 & n3991 ;
  assign n8203 = ~n8191 & ~n8202 ;
  assign n8204 = n993 & ~n8203 ;
  assign n8194 = n970 & ~n8193 ;
  assign n8205 = \InstQueue_reg[12][5]/NET0131  & ~n3933 ;
  assign n8206 = ~n8194 & ~n8205 ;
  assign n8207 = ~n8204 & n8206 ;
  assign n8208 = ~n8201 & n8207 ;
  assign n8214 = n3939 & n8135 ;
  assign n8215 = n3967 & n8138 ;
  assign n8216 = ~n8214 & ~n8215 ;
  assign n8217 = \DataWidth_reg[1]/NET0131  & ~n8216 ;
  assign n8209 = \Datai[5]_pad  & ~n4013 ;
  assign n8210 = \InstQueue_reg[13][5]/NET0131  & ~n3876 ;
  assign n8211 = ~n3991 & n8210 ;
  assign n8212 = ~n8209 & ~n8211 ;
  assign n8218 = ~n4023 & ~n8212 ;
  assign n8219 = ~n8217 & ~n8218 ;
  assign n8220 = n952 & ~n8219 ;
  assign n8221 = ~n697 & n3876 ;
  assign n8222 = ~n8210 & ~n8221 ;
  assign n8223 = n993 & ~n8222 ;
  assign n8213 = n970 & ~n8212 ;
  assign n8224 = \InstQueue_reg[13][5]/NET0131  & ~n3933 ;
  assign n8225 = ~n8213 & ~n8224 ;
  assign n8226 = ~n8223 & n8225 ;
  assign n8227 = ~n8220 & n8226 ;
  assign n8233 = n3967 & n8135 ;
  assign n8234 = n3991 & n8138 ;
  assign n8235 = ~n8233 & ~n8234 ;
  assign n8236 = \DataWidth_reg[1]/NET0131  & ~n8235 ;
  assign n8228 = \Datai[5]_pad  & ~n3923 ;
  assign n8229 = \InstQueue_reg[14][5]/NET0131  & ~n3919 ;
  assign n8230 = ~n3876 & n8229 ;
  assign n8231 = ~n8228 & ~n8230 ;
  assign n8237 = ~n4043 & ~n8231 ;
  assign n8238 = ~n8236 & ~n8237 ;
  assign n8239 = n952 & ~n8238 ;
  assign n8240 = ~n697 & n3919 ;
  assign n8241 = ~n8229 & ~n8240 ;
  assign n8242 = n993 & ~n8241 ;
  assign n8232 = n970 & ~n8231 ;
  assign n8243 = \InstQueue_reg[14][5]/NET0131  & ~n3933 ;
  assign n8244 = ~n8232 & ~n8243 ;
  assign n8245 = ~n8242 & n8244 ;
  assign n8246 = ~n8239 & n8245 ;
  assign n8252 = n3991 & n8135 ;
  assign n8253 = n3876 & n8138 ;
  assign n8254 = ~n8252 & ~n8253 ;
  assign n8255 = \DataWidth_reg[1]/NET0131  & ~n8254 ;
  assign n8247 = \Datai[5]_pad  & ~n4054 ;
  assign n8248 = \InstQueue_reg[15][5]/NET0131  & ~n3867 ;
  assign n8249 = ~n3919 & n8248 ;
  assign n8250 = ~n8247 & ~n8249 ;
  assign n8256 = ~n4064 & ~n8250 ;
  assign n8257 = ~n8255 & ~n8256 ;
  assign n8258 = n952 & ~n8257 ;
  assign n8259 = ~n697 & n3867 ;
  assign n8260 = ~n8248 & ~n8259 ;
  assign n8261 = n993 & ~n8260 ;
  assign n8251 = n970 & ~n8250 ;
  assign n8262 = \InstQueue_reg[15][5]/NET0131  & ~n3933 ;
  assign n8263 = ~n8251 & ~n8262 ;
  assign n8264 = ~n8261 & n8263 ;
  assign n8265 = ~n8258 & n8264 ;
  assign n8271 = n3919 & n8135 ;
  assign n8272 = n3867 & n8138 ;
  assign n8273 = ~n8271 & ~n8272 ;
  assign n8274 = \DataWidth_reg[1]/NET0131  & ~n8273 ;
  assign n8266 = \Datai[5]_pad  & ~n4076 ;
  assign n8267 = \InstQueue_reg[1][5]/NET0131  & ~n4075 ;
  assign n8268 = ~n3864 & n8267 ;
  assign n8269 = ~n8266 & ~n8268 ;
  assign n8275 = ~n4086 & ~n8269 ;
  assign n8276 = ~n8274 & ~n8275 ;
  assign n8277 = n952 & ~n8276 ;
  assign n8278 = ~n697 & n4075 ;
  assign n8279 = ~n8267 & ~n8278 ;
  assign n8280 = n993 & ~n8279 ;
  assign n8270 = n970 & ~n8269 ;
  assign n8281 = \InstQueue_reg[1][5]/NET0131  & ~n3933 ;
  assign n8282 = ~n8270 & ~n8281 ;
  assign n8283 = ~n8280 & n8282 ;
  assign n8284 = ~n8277 & n8283 ;
  assign n8290 = n3864 & n8138 ;
  assign n8291 = n3867 & n8135 ;
  assign n8292 = ~n8290 & ~n8291 ;
  assign n8293 = \DataWidth_reg[1]/NET0131  & ~n8292 ;
  assign n8285 = \Datai[5]_pad  & ~n4098 ;
  assign n8286 = \InstQueue_reg[2][5]/NET0131  & ~n4097 ;
  assign n8287 = ~n4075 & n8286 ;
  assign n8288 = ~n8285 & ~n8287 ;
  assign n8294 = ~n4108 & ~n8288 ;
  assign n8295 = ~n8293 & ~n8294 ;
  assign n8296 = n952 & ~n8295 ;
  assign n8297 = ~n697 & n4097 ;
  assign n8298 = ~n8286 & ~n8297 ;
  assign n8299 = n993 & ~n8298 ;
  assign n8289 = n970 & ~n8288 ;
  assign n8300 = \InstQueue_reg[2][5]/NET0131  & ~n3933 ;
  assign n8301 = ~n8289 & ~n8300 ;
  assign n8302 = ~n8299 & n8301 ;
  assign n8303 = ~n8296 & n8302 ;
  assign n8309 = n3864 & n8135 ;
  assign n8310 = n4075 & n8138 ;
  assign n8311 = ~n8309 & ~n8310 ;
  assign n8312 = \DataWidth_reg[1]/NET0131  & ~n8311 ;
  assign n8304 = \Datai[5]_pad  & ~n4120 ;
  assign n8305 = \InstQueue_reg[3][5]/NET0131  & ~n4119 ;
  assign n8306 = ~n4097 & n8305 ;
  assign n8307 = ~n8304 & ~n8306 ;
  assign n8313 = ~n4130 & ~n8307 ;
  assign n8314 = ~n8312 & ~n8313 ;
  assign n8315 = n952 & ~n8314 ;
  assign n8316 = ~n697 & n4119 ;
  assign n8317 = ~n8305 & ~n8316 ;
  assign n8318 = n993 & ~n8317 ;
  assign n8308 = n970 & ~n8307 ;
  assign n8319 = \InstQueue_reg[3][5]/NET0131  & ~n3933 ;
  assign n8320 = ~n8308 & ~n8319 ;
  assign n8321 = ~n8318 & n8320 ;
  assign n8322 = ~n8315 & n8321 ;
  assign n8328 = n4075 & n8135 ;
  assign n8329 = n4097 & n8138 ;
  assign n8330 = ~n8328 & ~n8329 ;
  assign n8331 = \DataWidth_reg[1]/NET0131  & ~n8330 ;
  assign n8323 = \Datai[5]_pad  & ~n4142 ;
  assign n8324 = \InstQueue_reg[4][5]/NET0131  & ~n4141 ;
  assign n8325 = ~n4119 & n8324 ;
  assign n8326 = ~n8323 & ~n8325 ;
  assign n8332 = ~n4152 & ~n8326 ;
  assign n8333 = ~n8331 & ~n8332 ;
  assign n8334 = n952 & ~n8333 ;
  assign n8335 = ~n697 & n4141 ;
  assign n8336 = ~n8324 & ~n8335 ;
  assign n8337 = n993 & ~n8336 ;
  assign n8327 = n970 & ~n8326 ;
  assign n8338 = \InstQueue_reg[4][5]/NET0131  & ~n3933 ;
  assign n8339 = ~n8327 & ~n8338 ;
  assign n8340 = ~n8337 & n8339 ;
  assign n8341 = ~n8334 & n8340 ;
  assign n8347 = n4097 & n8135 ;
  assign n8348 = n4119 & n8138 ;
  assign n8349 = ~n8347 & ~n8348 ;
  assign n8350 = \DataWidth_reg[1]/NET0131  & ~n8349 ;
  assign n8342 = \Datai[5]_pad  & ~n4164 ;
  assign n8343 = \InstQueue_reg[5][5]/NET0131  & ~n4163 ;
  assign n8344 = ~n4141 & n8343 ;
  assign n8345 = ~n8342 & ~n8344 ;
  assign n8351 = ~n4174 & ~n8345 ;
  assign n8352 = ~n8350 & ~n8351 ;
  assign n8353 = n952 & ~n8352 ;
  assign n8354 = ~n697 & n4163 ;
  assign n8355 = ~n8343 & ~n8354 ;
  assign n8356 = n993 & ~n8355 ;
  assign n8346 = n970 & ~n8345 ;
  assign n8357 = \InstQueue_reg[5][5]/NET0131  & ~n3933 ;
  assign n8358 = ~n8346 & ~n8357 ;
  assign n8359 = ~n8356 & n8358 ;
  assign n8360 = ~n8353 & n8359 ;
  assign n8366 = n4119 & n8135 ;
  assign n8367 = n4141 & n8138 ;
  assign n8368 = ~n8366 & ~n8367 ;
  assign n8369 = \DataWidth_reg[1]/NET0131  & ~n8368 ;
  assign n8361 = \Datai[5]_pad  & ~n4186 ;
  assign n8362 = \InstQueue_reg[6][5]/NET0131  & ~n4185 ;
  assign n8363 = ~n4163 & n8362 ;
  assign n8364 = ~n8361 & ~n8363 ;
  assign n8370 = ~n4196 & ~n8364 ;
  assign n8371 = ~n8369 & ~n8370 ;
  assign n8372 = n952 & ~n8371 ;
  assign n8373 = ~n697 & n4185 ;
  assign n8374 = ~n8362 & ~n8373 ;
  assign n8375 = n993 & ~n8374 ;
  assign n8365 = n970 & ~n8364 ;
  assign n8376 = \InstQueue_reg[6][5]/NET0131  & ~n3933 ;
  assign n8377 = ~n8365 & ~n8376 ;
  assign n8378 = ~n8375 & n8377 ;
  assign n8379 = ~n8372 & n8378 ;
  assign n8385 = n4141 & n8135 ;
  assign n8386 = n4163 & n8138 ;
  assign n8387 = ~n8385 & ~n8386 ;
  assign n8388 = \DataWidth_reg[1]/NET0131  & ~n8387 ;
  assign n8380 = \Datai[5]_pad  & ~n4207 ;
  assign n8381 = \InstQueue_reg[7][5]/NET0131  & ~n3948 ;
  assign n8382 = ~n4185 & n8381 ;
  assign n8383 = ~n8380 & ~n8382 ;
  assign n8389 = ~n4217 & ~n8383 ;
  assign n8390 = ~n8388 & ~n8389 ;
  assign n8391 = n952 & ~n8390 ;
  assign n8392 = ~n697 & n3948 ;
  assign n8393 = ~n8381 & ~n8392 ;
  assign n8394 = n993 & ~n8393 ;
  assign n8384 = n970 & ~n8383 ;
  assign n8395 = \InstQueue_reg[7][5]/NET0131  & ~n3933 ;
  assign n8396 = ~n8384 & ~n8395 ;
  assign n8397 = ~n8394 & n8396 ;
  assign n8398 = ~n8391 & n8397 ;
  assign n8404 = n4163 & n8135 ;
  assign n8405 = n4185 & n8138 ;
  assign n8406 = ~n8404 & ~n8405 ;
  assign n8407 = \DataWidth_reg[1]/NET0131  & ~n8406 ;
  assign n8399 = \Datai[5]_pad  & ~n3954 ;
  assign n8400 = \InstQueue_reg[8][5]/NET0131  & ~n3950 ;
  assign n8401 = ~n3948 & n8400 ;
  assign n8402 = ~n8399 & ~n8401 ;
  assign n8408 = ~n4237 & ~n8402 ;
  assign n8409 = ~n8407 & ~n8408 ;
  assign n8410 = n952 & ~n8409 ;
  assign n8411 = ~n697 & n3950 ;
  assign n8412 = ~n8400 & ~n8411 ;
  assign n8413 = n993 & ~n8412 ;
  assign n8403 = n970 & ~n8402 ;
  assign n8414 = \InstQueue_reg[8][5]/NET0131  & ~n3933 ;
  assign n8415 = ~n8403 & ~n8414 ;
  assign n8416 = ~n8413 & n8415 ;
  assign n8417 = ~n8410 & n8416 ;
  assign n8423 = n4185 & n8135 ;
  assign n8424 = n3948 & n8138 ;
  assign n8425 = ~n8423 & ~n8424 ;
  assign n8426 = \DataWidth_reg[1]/NET0131  & ~n8425 ;
  assign n8418 = \Datai[5]_pad  & ~n3978 ;
  assign n8419 = \InstQueue_reg[9][5]/NET0131  & ~n3941 ;
  assign n8420 = ~n3950 & n8419 ;
  assign n8421 = ~n8418 & ~n8420 ;
  assign n8427 = ~n4257 & ~n8421 ;
  assign n8428 = ~n8426 & ~n8427 ;
  assign n8429 = n952 & ~n8428 ;
  assign n8430 = ~n697 & n3941 ;
  assign n8431 = ~n8419 & ~n8430 ;
  assign n8432 = n993 & ~n8431 ;
  assign n8422 = n970 & ~n8421 ;
  assign n8433 = \InstQueue_reg[9][5]/NET0131  & ~n3933 ;
  assign n8434 = ~n8422 & ~n8433 ;
  assign n8435 = ~n8432 & n8434 ;
  assign n8436 = ~n8429 & n8435 ;
  assign n8447 = ~\rEIP_reg[0]/NET0131  & ~\rEIP_reg[1]/NET0131  ;
  assign n8448 = \rEIP_reg[31]/NET0131  & ~n8447 ;
  assign n8449 = \rEIP_reg[2]/NET0131  & n8448 ;
  assign n8450 = \rEIP_reg[3]/NET0131  & n8449 ;
  assign n8451 = \rEIP_reg[4]/NET0131  & n8450 ;
  assign n8452 = \rEIP_reg[5]/NET0131  & n8451 ;
  assign n8453 = \rEIP_reg[6]/NET0131  & n8452 ;
  assign n8454 = \rEIP_reg[7]/NET0131  & n8453 ;
  assign n8455 = \rEIP_reg[8]/NET0131  & n8454 ;
  assign n8456 = \rEIP_reg[9]/NET0131  & n8455 ;
  assign n8457 = \rEIP_reg[10]/NET0131  & n8456 ;
  assign n8458 = \rEIP_reg[11]/NET0131  & n8457 ;
  assign n8459 = \rEIP_reg[12]/NET0131  & n8458 ;
  assign n8460 = \rEIP_reg[13]/NET0131  & n8459 ;
  assign n8461 = \rEIP_reg[14]/NET0131  & n8460 ;
  assign n8462 = \rEIP_reg[15]/NET0131  & n8461 ;
  assign n8463 = \rEIP_reg[16]/NET0131  & n8462 ;
  assign n8464 = n4671 & n8463 ;
  assign n8465 = n4652 & n8464 ;
  assign n8466 = n4674 & n8465 ;
  assign n8467 = \rEIP_reg[26]/NET0131  & n8466 ;
  assign n8468 = n4678 & n8467 ;
  assign n8469 = ~\rEIP_reg[30]/NET0131  & ~n8468 ;
  assign n8470 = n4679 & n8467 ;
  assign n8471 = n830 & ~n8470 ;
  assign n8472 = ~n8469 & n8471 ;
  assign n8437 = \Address[28]_pad  & ~n829 ;
  assign n8439 = \rEIP_reg[0]/NET0131  & \rEIP_reg[31]/NET0131  ;
  assign n8440 = n4673 & n8439 ;
  assign n8441 = n4675 & n8440 ;
  assign n8442 = n4677 & n8441 ;
  assign n8443 = ~\rEIP_reg[29]/NET0131  & ~n8442 ;
  assign n8438 = \State_reg[2]/NET0131  & n829 ;
  assign n8444 = n4678 & n8441 ;
  assign n8445 = n8438 & ~n8444 ;
  assign n8446 = ~n8443 & n8445 ;
  assign n8473 = ~n8437 & ~n8446 ;
  assign n8474 = ~n8472 & n8473 ;
  assign n8476 = \Datao[25]_pad  & ~n4286 ;
  assign n8477 = ~n833 & n7435 ;
  assign n8478 = ~n8476 & ~n8477 ;
  assign n8479 = n948 & ~n8478 ;
  assign n8475 = \uWord_reg[9]/NET0131  & n956 ;
  assign n8480 = \Datao[25]_pad  & ~n3816 ;
  assign n8481 = ~n8475 & ~n8480 ;
  assign n8482 = ~n8479 & n8481 ;
  assign n8484 = ~n833 & ~n7400 ;
  assign n8485 = n3798 & ~n8484 ;
  assign n8486 = n3806 & ~n8485 ;
  assign n8487 = \Datao[17]_pad  & ~n8486 ;
  assign n8488 = ~n833 & n7401 ;
  assign n8489 = ~n8487 & ~n8488 ;
  assign n8490 = n948 & ~n8489 ;
  assign n8483 = \uWord_reg[1]/NET0131  & n956 ;
  assign n8491 = \Datao[17]_pad  & ~n3816 ;
  assign n8492 = ~n8483 & ~n8491 ;
  assign n8493 = ~n8490 & n8492 ;
  assign n8495 = ~n833 & ~n7374 ;
  assign n8496 = n3798 & ~n8495 ;
  assign n8497 = n3806 & ~n8496 ;
  assign n8498 = \Datao[16]_pad  & ~n8497 ;
  assign n8499 = ~n833 & n7375 ;
  assign n8500 = ~n8498 & ~n8499 ;
  assign n8501 = n948 & ~n8500 ;
  assign n8494 = \uWord_reg[0]/NET0131  & n956 ;
  assign n8502 = \Datao[16]_pad  & ~n3816 ;
  assign n8503 = ~n8494 & ~n8502 ;
  assign n8504 = ~n8501 & n8503 ;
  assign n8506 = \Datao[21]_pad  & ~n4286 ;
  assign n8507 = n895 & n7419 ;
  assign n8508 = ~n8506 & ~n8507 ;
  assign n8509 = n948 & ~n8508 ;
  assign n8505 = \uWord_reg[5]/NET0131  & n956 ;
  assign n8510 = \Datao[21]_pad  & ~n3816 ;
  assign n8511 = ~n8505 & ~n8510 ;
  assign n8512 = ~n8509 & n8511 ;
  assign n8513 = ~\Flush_reg/NET0131  & n988 ;
  assign n8514 = n973 & ~n981 ;
  assign n8515 = ~n8513 & n8514 ;
  assign n8516 = n6849 & n8515 ;
  assign n8517 = \InstQueueWr_Addr_reg[2]/NET0131  & ~n8516 ;
  assign n8518 = ~n2038 & ~n3917 ;
  assign n8519 = \InstQueueWr_Addr_reg[2]/NET0131  & ~n8518 ;
  assign n8520 = ~n2037 & ~n8519 ;
  assign n8521 = ~n993 & ~n8520 ;
  assign n8522 = ~n2037 & n3917 ;
  assign n8523 = ~\InstQueueWr_Addr_reg[2]/NET0131  & ~n3865 ;
  assign n8524 = ~n971 & n8523 ;
  assign n8525 = ~n8522 & n8524 ;
  assign n8526 = ~n3866 & ~n8525 ;
  assign n8527 = ~n8521 & n8526 ;
  assign n8528 = ~n8517 & ~n8527 ;
  assign n8537 = \rEIP_reg[17]/NET0131  & n8463 ;
  assign n8538 = ~\rEIP_reg[18]/NET0131  & ~n8537 ;
  assign n8539 = n4668 & n8463 ;
  assign n8540 = n830 & ~n8539 ;
  assign n8541 = ~n8538 & n8540 ;
  assign n8529 = \Address[16]_pad  & ~n829 ;
  assign n8530 = n4665 & n8439 ;
  assign n8531 = \rEIP_reg[15]/NET0131  & n8530 ;
  assign n8532 = \rEIP_reg[16]/NET0131  & n8531 ;
  assign n8534 = ~\rEIP_reg[17]/NET0131  & ~n8532 ;
  assign n8533 = \rEIP_reg[17]/NET0131  & n8532 ;
  assign n8535 = n8438 & ~n8533 ;
  assign n8536 = ~n8534 & n8535 ;
  assign n8542 = ~n8529 & ~n8536 ;
  assign n8543 = ~n8541 & n8542 ;
  assign n8547 = ~\EAX_reg[2]/NET0131  & n4286 ;
  assign n8546 = ~\Datao[2]_pad  & ~n4286 ;
  assign n8548 = n948 & ~n8546 ;
  assign n8549 = ~n8547 & n8548 ;
  assign n8544 = \lWord_reg[2]/NET0131  & n956 ;
  assign n8545 = \Datao[2]_pad  & ~n3816 ;
  assign n8550 = ~n8544 & ~n8545 ;
  assign n8551 = ~n8549 & n8550 ;
  assign n8555 = ~\EAX_reg[3]/NET0131  & n4286 ;
  assign n8554 = ~\Datao[3]_pad  & ~n4286 ;
  assign n8556 = n948 & ~n8554 ;
  assign n8557 = ~n8555 & n8556 ;
  assign n8552 = \lWord_reg[3]/NET0131  & n956 ;
  assign n8553 = \Datao[3]_pad  & ~n3816 ;
  assign n8558 = ~n8552 & ~n8553 ;
  assign n8559 = ~n8557 & n8558 ;
  assign n8563 = ~\EAX_reg[4]/NET0131  & n4286 ;
  assign n8562 = ~\Datao[4]_pad  & ~n4286 ;
  assign n8564 = n948 & ~n8562 ;
  assign n8565 = ~n8563 & n8564 ;
  assign n8560 = \lWord_reg[4]/NET0131  & n956 ;
  assign n8561 = \Datao[4]_pad  & ~n3816 ;
  assign n8566 = ~n8560 & ~n8561 ;
  assign n8567 = ~n8565 & n8566 ;
  assign n8571 = ~\EAX_reg[5]/NET0131  & n4286 ;
  assign n8570 = ~\Datao[5]_pad  & ~n4286 ;
  assign n8572 = n948 & ~n8570 ;
  assign n8573 = ~n8571 & n8572 ;
  assign n8568 = \lWord_reg[5]/NET0131  & n956 ;
  assign n8569 = \Datao[5]_pad  & ~n3816 ;
  assign n8574 = ~n8568 & ~n8569 ;
  assign n8575 = ~n8573 & n8574 ;
  assign n8579 = ~\EAX_reg[6]/NET0131  & n4286 ;
  assign n8578 = ~\Datao[6]_pad  & ~n4286 ;
  assign n8580 = n948 & ~n8578 ;
  assign n8581 = ~n8579 & n8580 ;
  assign n8576 = \lWord_reg[6]/NET0131  & n956 ;
  assign n8577 = \Datao[6]_pad  & ~n3816 ;
  assign n8582 = ~n8576 & ~n8577 ;
  assign n8583 = ~n8581 & n8582 ;
  assign n8587 = ~\EAX_reg[7]/NET0131  & n4286 ;
  assign n8586 = ~\Datao[7]_pad  & ~n4286 ;
  assign n8588 = n948 & ~n8586 ;
  assign n8589 = ~n8587 & n8588 ;
  assign n8584 = \lWord_reg[7]/NET0131  & n956 ;
  assign n8585 = \Datao[7]_pad  & ~n3816 ;
  assign n8590 = ~n8584 & ~n8585 ;
  assign n8591 = ~n8589 & n8590 ;
  assign n8595 = ~\EAX_reg[8]/NET0131  & n4286 ;
  assign n8594 = ~\Datao[8]_pad  & ~n4286 ;
  assign n8596 = n948 & ~n8594 ;
  assign n8597 = ~n8595 & n8596 ;
  assign n8592 = \lWord_reg[8]/NET0131  & n956 ;
  assign n8593 = \Datao[8]_pad  & ~n3816 ;
  assign n8598 = ~n8592 & ~n8593 ;
  assign n8599 = ~n8597 & n8598 ;
  assign n8603 = ~\EAX_reg[9]/NET0131  & n4286 ;
  assign n8602 = ~\Datao[9]_pad  & ~n4286 ;
  assign n8604 = n948 & ~n8602 ;
  assign n8605 = ~n8603 & n8604 ;
  assign n8600 = \lWord_reg[9]/NET0131  & n956 ;
  assign n8601 = \Datao[9]_pad  & ~n3816 ;
  assign n8606 = ~n8600 & ~n8601 ;
  assign n8607 = ~n8605 & n8606 ;
  assign n8611 = ~\EAX_reg[0]/NET0131  & n4286 ;
  assign n8610 = ~\Datao[0]_pad  & ~n4286 ;
  assign n8612 = n948 & ~n8610 ;
  assign n8613 = ~n8611 & n8612 ;
  assign n8608 = \lWord_reg[0]/NET0131  & n956 ;
  assign n8609 = \Datao[0]_pad  & ~n3816 ;
  assign n8614 = ~n8608 & ~n8609 ;
  assign n8615 = ~n8613 & n8614 ;
  assign n8619 = ~\EAX_reg[10]/NET0131  & n4286 ;
  assign n8618 = ~\Datao[10]_pad  & ~n4286 ;
  assign n8620 = n948 & ~n8618 ;
  assign n8621 = ~n8619 & n8620 ;
  assign n8616 = \lWord_reg[10]/NET0131  & n956 ;
  assign n8617 = \Datao[10]_pad  & ~n3816 ;
  assign n8622 = ~n8616 & ~n8617 ;
  assign n8623 = ~n8621 & n8622 ;
  assign n8627 = ~\EAX_reg[12]/NET0131  & n4286 ;
  assign n8626 = ~\Datao[12]_pad  & ~n4286 ;
  assign n8628 = n948 & ~n8626 ;
  assign n8629 = ~n8627 & n8628 ;
  assign n8624 = \lWord_reg[12]/NET0131  & n956 ;
  assign n8625 = \Datao[12]_pad  & ~n3816 ;
  assign n8630 = ~n8624 & ~n8625 ;
  assign n8631 = ~n8629 & n8630 ;
  assign n8635 = ~\EAX_reg[11]/NET0131  & n4286 ;
  assign n8634 = ~\Datao[11]_pad  & ~n4286 ;
  assign n8636 = n948 & ~n8634 ;
  assign n8637 = ~n8635 & n8636 ;
  assign n8632 = \lWord_reg[11]/NET0131  & n956 ;
  assign n8633 = \Datao[11]_pad  & ~n3816 ;
  assign n8638 = ~n8632 & ~n8633 ;
  assign n8639 = ~n8637 & n8638 ;
  assign n8643 = ~\EAX_reg[13]/NET0131  & n4286 ;
  assign n8642 = ~\Datao[13]_pad  & ~n4286 ;
  assign n8644 = n948 & ~n8642 ;
  assign n8645 = ~n8643 & n8644 ;
  assign n8640 = \lWord_reg[13]/NET0131  & n956 ;
  assign n8641 = \Datao[13]_pad  & ~n3816 ;
  assign n8646 = ~n8640 & ~n8641 ;
  assign n8647 = ~n8645 & n8646 ;
  assign n8651 = ~\EAX_reg[14]/NET0131  & n4286 ;
  assign n8650 = ~\Datao[14]_pad  & ~n4286 ;
  assign n8652 = n948 & ~n8650 ;
  assign n8653 = ~n8651 & n8652 ;
  assign n8648 = \lWord_reg[14]/NET0131  & n956 ;
  assign n8649 = \Datao[14]_pad  & ~n3816 ;
  assign n8654 = ~n8648 & ~n8649 ;
  assign n8655 = ~n8653 & n8654 ;
  assign n8659 = ~\EAX_reg[15]/NET0131  & n4286 ;
  assign n8658 = ~\Datao[15]_pad  & ~n4286 ;
  assign n8660 = n948 & ~n8658 ;
  assign n8661 = ~n8659 & n8660 ;
  assign n8656 = \lWord_reg[15]/NET0131  & n956 ;
  assign n8657 = \Datao[15]_pad  & ~n3816 ;
  assign n8662 = ~n8656 & ~n8657 ;
  assign n8663 = ~n8661 & n8662 ;
  assign n8667 = ~\EAX_reg[1]/NET0131  & n4286 ;
  assign n8666 = ~\Datao[1]_pad  & ~n4286 ;
  assign n8668 = n948 & ~n8666 ;
  assign n8669 = ~n8667 & n8668 ;
  assign n8664 = \lWord_reg[1]/NET0131  & n956 ;
  assign n8665 = \Datao[1]_pad  & ~n3816 ;
  assign n8670 = ~n8664 & ~n8665 ;
  assign n8671 = ~n8669 & n8670 ;
  assign n8676 = n971 & ~n3991 ;
  assign n8679 = ~n3875 & n8676 ;
  assign n8680 = ~n2039 & ~n8679 ;
  assign n8672 = \InstQueueWr_Addr_reg[3]/NET0131  & ~n3866 ;
  assign n8673 = ~n3948 & ~n8672 ;
  assign n8681 = ~n3918 & n8673 ;
  assign n8682 = ~n3919 & ~n8681 ;
  assign n8683 = ~n8680 & n8682 ;
  assign n8675 = \InstQueueWr_Addr_reg[3]/NET0131  & ~n8516 ;
  assign n8674 = n993 & ~n8673 ;
  assign n8677 = ~n3990 & ~n4163 ;
  assign n8678 = n8676 & ~n8677 ;
  assign n8684 = ~n8674 & ~n8678 ;
  assign n8685 = ~n8675 & n8684 ;
  assign n8686 = ~n8683 & n8685 ;
  assign n8687 = \InstQueueWr_Addr_reg[1]/NET0131  & ~n8515 ;
  assign n8688 = ~\InstQueueWr_Addr_reg[0]/NET0131  & n993 ;
  assign n8689 = \InstQueueWr_Addr_reg[1]/NET0131  & n6849 ;
  assign n8690 = ~n971 & n8689 ;
  assign n8691 = ~n8688 & n8690 ;
  assign n8692 = \InstQueueWr_Addr_reg[0]/NET0131  & n993 ;
  assign n8693 = ~\InstQueueWr_Addr_reg[1]/NET0131  & ~n8692 ;
  assign n8694 = ~n2039 & n8693 ;
  assign n8695 = ~n8691 & ~n8694 ;
  assign n8696 = ~n8687 & ~n8695 ;
  assign n8699 = ~n948 & n3630 ;
  assign n8700 = \InstQueueWr_Addr_reg[0]/NET0131  & ~n8699 ;
  assign n8697 = ~\Flush_reg/NET0131  & ~\InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n8698 = n988 & ~n8697 ;
  assign n8701 = ~n8688 & ~n8698 ;
  assign n8702 = ~n8700 & n8701 ;
  assign n8708 = ~\Datai[25]_pad  & ~n3901 ;
  assign n8709 = ~n3902 & ~n8708 ;
  assign n8710 = n3876 & n8709 ;
  assign n8711 = ~\Datai[17]_pad  & ~n3910 ;
  assign n8712 = ~n3911 & ~n8711 ;
  assign n8713 = n3919 & n8712 ;
  assign n8714 = ~n8710 & ~n8713 ;
  assign n8715 = \DataWidth_reg[1]/NET0131  & ~n8714 ;
  assign n8703 = \Datai[1]_pad  & ~n3868 ;
  assign n8704 = \InstQueue_reg[0][1]/NET0131  & ~n3864 ;
  assign n8705 = ~n3867 & n8704 ;
  assign n8706 = ~n8703 & ~n8705 ;
  assign n8716 = ~n3924 & ~n8706 ;
  assign n8717 = ~n8715 & ~n8716 ;
  assign n8718 = n952 & ~n8717 ;
  assign n8719 = ~n600 & n3864 ;
  assign n8720 = ~n8704 & ~n8719 ;
  assign n8721 = n993 & ~n8720 ;
  assign n8707 = n970 & ~n8706 ;
  assign n8722 = \InstQueue_reg[0][1]/NET0131  & ~n3933 ;
  assign n8723 = ~n8707 & ~n8722 ;
  assign n8724 = ~n8721 & n8723 ;
  assign n8725 = ~n8718 & n8724 ;
  assign n8731 = n3948 & n8709 ;
  assign n8732 = n3950 & n8712 ;
  assign n8733 = ~n8731 & ~n8732 ;
  assign n8734 = \DataWidth_reg[1]/NET0131  & ~n8733 ;
  assign n8726 = \Datai[1]_pad  & ~n3942 ;
  assign n8727 = \InstQueue_reg[10][1]/NET0131  & ~n3939 ;
  assign n8728 = ~n3941 & n8727 ;
  assign n8729 = ~n8726 & ~n8728 ;
  assign n8735 = ~n3955 & ~n8729 ;
  assign n8736 = ~n8734 & ~n8735 ;
  assign n8737 = n952 & ~n8736 ;
  assign n8738 = ~n600 & n3939 ;
  assign n8739 = ~n8727 & ~n8738 ;
  assign n8740 = n993 & ~n8739 ;
  assign n8730 = n970 & ~n8729 ;
  assign n8741 = \InstQueue_reg[10][1]/NET0131  & ~n3933 ;
  assign n8742 = ~n8730 & ~n8741 ;
  assign n8743 = ~n8740 & n8742 ;
  assign n8744 = ~n8737 & n8743 ;
  assign n8750 = ~\Datai[24]_pad  & ~n3900 ;
  assign n8751 = ~n3901 & ~n8750 ;
  assign n8752 = n3950 & n8751 ;
  assign n8753 = ~\Datai[16]_pad  & ~n3909 ;
  assign n8754 = ~n3910 & ~n8753 ;
  assign n8755 = n3941 & n8754 ;
  assign n8756 = ~n8752 & ~n8755 ;
  assign n8757 = \DataWidth_reg[1]/NET0131  & ~n8756 ;
  assign n8745 = \Datai[0]_pad  & ~n3968 ;
  assign n8746 = \InstQueue_reg[11][0]/NET0131  & ~n3967 ;
  assign n8747 = ~n3939 & n8746 ;
  assign n8748 = ~n8745 & ~n8747 ;
  assign n8758 = ~n3979 & ~n8748 ;
  assign n8759 = ~n8757 & ~n8758 ;
  assign n8760 = n952 & ~n8759 ;
  assign n8761 = ~n663 & n3967 ;
  assign n8762 = ~n8746 & ~n8761 ;
  assign n8763 = n993 & ~n8762 ;
  assign n8749 = n970 & ~n8748 ;
  assign n8764 = \InstQueue_reg[11][0]/NET0131  & ~n3933 ;
  assign n8765 = ~n8749 & ~n8764 ;
  assign n8766 = ~n8763 & n8765 ;
  assign n8767 = ~n8760 & n8766 ;
  assign n8773 = n3950 & n8709 ;
  assign n8774 = n3941 & n8712 ;
  assign n8775 = ~n8773 & ~n8774 ;
  assign n8776 = \DataWidth_reg[1]/NET0131  & ~n8775 ;
  assign n8768 = \Datai[1]_pad  & ~n3968 ;
  assign n8769 = \InstQueue_reg[11][1]/NET0131  & ~n3967 ;
  assign n8770 = ~n3939 & n8769 ;
  assign n8771 = ~n8768 & ~n8770 ;
  assign n8777 = ~n3979 & ~n8771 ;
  assign n8778 = ~n8776 & ~n8777 ;
  assign n8779 = n952 & ~n8778 ;
  assign n8780 = ~n600 & n3967 ;
  assign n8781 = ~n8769 & ~n8780 ;
  assign n8782 = n993 & ~n8781 ;
  assign n8772 = n970 & ~n8771 ;
  assign n8783 = \InstQueue_reg[11][1]/NET0131  & ~n3933 ;
  assign n8784 = ~n8772 & ~n8783 ;
  assign n8785 = ~n8782 & n8784 ;
  assign n8786 = ~n8779 & n8785 ;
  assign n8792 = n3941 & n8709 ;
  assign n8793 = n3939 & n8712 ;
  assign n8794 = ~n8792 & ~n8793 ;
  assign n8795 = \DataWidth_reg[1]/NET0131  & ~n8794 ;
  assign n8787 = \Datai[1]_pad  & ~n3992 ;
  assign n8788 = \InstQueue_reg[12][1]/NET0131  & ~n3991 ;
  assign n8789 = ~n3967 & n8788 ;
  assign n8790 = ~n8787 & ~n8789 ;
  assign n8796 = ~n4002 & ~n8790 ;
  assign n8797 = ~n8795 & ~n8796 ;
  assign n8798 = n952 & ~n8797 ;
  assign n8799 = ~n600 & n3991 ;
  assign n8800 = ~n8788 & ~n8799 ;
  assign n8801 = n993 & ~n8800 ;
  assign n8791 = n970 & ~n8790 ;
  assign n8802 = \InstQueue_reg[12][1]/NET0131  & ~n3933 ;
  assign n8803 = ~n8791 & ~n8802 ;
  assign n8804 = ~n8801 & n8803 ;
  assign n8805 = ~n8798 & n8804 ;
  assign n8811 = n3939 & n8709 ;
  assign n8812 = n3967 & n8712 ;
  assign n8813 = ~n8811 & ~n8812 ;
  assign n8814 = \DataWidth_reg[1]/NET0131  & ~n8813 ;
  assign n8806 = \Datai[1]_pad  & ~n4013 ;
  assign n8807 = \InstQueue_reg[13][1]/NET0131  & ~n3876 ;
  assign n8808 = ~n3991 & n8807 ;
  assign n8809 = ~n8806 & ~n8808 ;
  assign n8815 = ~n4023 & ~n8809 ;
  assign n8816 = ~n8814 & ~n8815 ;
  assign n8817 = n952 & ~n8816 ;
  assign n8818 = ~n600 & n3876 ;
  assign n8819 = ~n8807 & ~n8818 ;
  assign n8820 = n993 & ~n8819 ;
  assign n8810 = n970 & ~n8809 ;
  assign n8821 = \InstQueue_reg[13][1]/NET0131  & ~n3933 ;
  assign n8822 = ~n8810 & ~n8821 ;
  assign n8823 = ~n8820 & n8822 ;
  assign n8824 = ~n8817 & n8823 ;
  assign n8830 = n3967 & n8709 ;
  assign n8831 = n3991 & n8712 ;
  assign n8832 = ~n8830 & ~n8831 ;
  assign n8833 = \DataWidth_reg[1]/NET0131  & ~n8832 ;
  assign n8825 = \Datai[1]_pad  & ~n3923 ;
  assign n8826 = \InstQueue_reg[14][1]/NET0131  & ~n3919 ;
  assign n8827 = ~n3876 & n8826 ;
  assign n8828 = ~n8825 & ~n8827 ;
  assign n8834 = ~n4043 & ~n8828 ;
  assign n8835 = ~n8833 & ~n8834 ;
  assign n8836 = n952 & ~n8835 ;
  assign n8837 = ~n600 & n3919 ;
  assign n8838 = ~n8826 & ~n8837 ;
  assign n8839 = n993 & ~n8838 ;
  assign n8829 = n970 & ~n8828 ;
  assign n8840 = \InstQueue_reg[14][1]/NET0131  & ~n3933 ;
  assign n8841 = ~n8829 & ~n8840 ;
  assign n8842 = ~n8839 & n8841 ;
  assign n8843 = ~n8836 & n8842 ;
  assign n8849 = n3991 & n8709 ;
  assign n8850 = n3876 & n8712 ;
  assign n8851 = ~n8849 & ~n8850 ;
  assign n8852 = \DataWidth_reg[1]/NET0131  & ~n8851 ;
  assign n8844 = \Datai[1]_pad  & ~n4054 ;
  assign n8845 = \InstQueue_reg[15][1]/NET0131  & ~n3867 ;
  assign n8846 = ~n3919 & n8845 ;
  assign n8847 = ~n8844 & ~n8846 ;
  assign n8853 = ~n4064 & ~n8847 ;
  assign n8854 = ~n8852 & ~n8853 ;
  assign n8855 = n952 & ~n8854 ;
  assign n8856 = ~n600 & n3867 ;
  assign n8857 = ~n8845 & ~n8856 ;
  assign n8858 = n993 & ~n8857 ;
  assign n8848 = n970 & ~n8847 ;
  assign n8859 = \InstQueue_reg[15][1]/NET0131  & ~n3933 ;
  assign n8860 = ~n8848 & ~n8859 ;
  assign n8861 = ~n8858 & n8860 ;
  assign n8862 = ~n8855 & n8861 ;
  assign n8868 = n3919 & n8709 ;
  assign n8869 = n3867 & n8712 ;
  assign n8870 = ~n8868 & ~n8869 ;
  assign n8871 = \DataWidth_reg[1]/NET0131  & ~n8870 ;
  assign n8863 = \Datai[1]_pad  & ~n4076 ;
  assign n8864 = \InstQueue_reg[1][1]/NET0131  & ~n4075 ;
  assign n8865 = ~n3864 & n8864 ;
  assign n8866 = ~n8863 & ~n8865 ;
  assign n8872 = ~n4086 & ~n8866 ;
  assign n8873 = ~n8871 & ~n8872 ;
  assign n8874 = n952 & ~n8873 ;
  assign n8875 = ~n600 & n4075 ;
  assign n8876 = ~n8864 & ~n8875 ;
  assign n8877 = n993 & ~n8876 ;
  assign n8867 = n970 & ~n8866 ;
  assign n8878 = \InstQueue_reg[1][1]/NET0131  & ~n3933 ;
  assign n8879 = ~n8867 & ~n8878 ;
  assign n8880 = ~n8877 & n8879 ;
  assign n8881 = ~n8874 & n8880 ;
  assign n8887 = n3864 & n8712 ;
  assign n8888 = n3867 & n8709 ;
  assign n8889 = ~n8887 & ~n8888 ;
  assign n8890 = \DataWidth_reg[1]/NET0131  & ~n8889 ;
  assign n8882 = \Datai[1]_pad  & ~n4098 ;
  assign n8883 = \InstQueue_reg[2][1]/NET0131  & ~n4097 ;
  assign n8884 = ~n4075 & n8883 ;
  assign n8885 = ~n8882 & ~n8884 ;
  assign n8891 = ~n4108 & ~n8885 ;
  assign n8892 = ~n8890 & ~n8891 ;
  assign n8893 = n952 & ~n8892 ;
  assign n8894 = ~n600 & n4097 ;
  assign n8895 = ~n8883 & ~n8894 ;
  assign n8896 = n993 & ~n8895 ;
  assign n8886 = n970 & ~n8885 ;
  assign n8897 = \InstQueue_reg[2][1]/NET0131  & ~n3933 ;
  assign n8898 = ~n8886 & ~n8897 ;
  assign n8899 = ~n8896 & n8898 ;
  assign n8900 = ~n8893 & n8899 ;
  assign n8906 = n3864 & n8751 ;
  assign n8907 = n4075 & n8754 ;
  assign n8908 = ~n8906 & ~n8907 ;
  assign n8909 = \DataWidth_reg[1]/NET0131  & ~n8908 ;
  assign n8901 = \Datai[0]_pad  & ~n4120 ;
  assign n8902 = \InstQueue_reg[3][0]/NET0131  & ~n4119 ;
  assign n8903 = ~n4097 & n8902 ;
  assign n8904 = ~n8901 & ~n8903 ;
  assign n8910 = ~n4130 & ~n8904 ;
  assign n8911 = ~n8909 & ~n8910 ;
  assign n8912 = n952 & ~n8911 ;
  assign n8913 = ~n663 & n4119 ;
  assign n8914 = ~n8902 & ~n8913 ;
  assign n8915 = n993 & ~n8914 ;
  assign n8905 = n970 & ~n8904 ;
  assign n8916 = \InstQueue_reg[3][0]/NET0131  & ~n3933 ;
  assign n8917 = ~n8905 & ~n8916 ;
  assign n8918 = ~n8915 & n8917 ;
  assign n8919 = ~n8912 & n8918 ;
  assign n8925 = n3864 & n8709 ;
  assign n8926 = n4075 & n8712 ;
  assign n8927 = ~n8925 & ~n8926 ;
  assign n8928 = \DataWidth_reg[1]/NET0131  & ~n8927 ;
  assign n8920 = \Datai[1]_pad  & ~n4120 ;
  assign n8921 = \InstQueue_reg[3][1]/NET0131  & ~n4119 ;
  assign n8922 = ~n4097 & n8921 ;
  assign n8923 = ~n8920 & ~n8922 ;
  assign n8929 = ~n4130 & ~n8923 ;
  assign n8930 = ~n8928 & ~n8929 ;
  assign n8931 = n952 & ~n8930 ;
  assign n8932 = ~n600 & n4119 ;
  assign n8933 = ~n8921 & ~n8932 ;
  assign n8934 = n993 & ~n8933 ;
  assign n8924 = n970 & ~n8923 ;
  assign n8935 = \InstQueue_reg[3][1]/NET0131  & ~n3933 ;
  assign n8936 = ~n8924 & ~n8935 ;
  assign n8937 = ~n8934 & n8936 ;
  assign n8938 = ~n8931 & n8937 ;
  assign n8944 = n4075 & n8709 ;
  assign n8945 = n4097 & n8712 ;
  assign n8946 = ~n8944 & ~n8945 ;
  assign n8947 = \DataWidth_reg[1]/NET0131  & ~n8946 ;
  assign n8939 = \Datai[1]_pad  & ~n4142 ;
  assign n8940 = \InstQueue_reg[4][1]/NET0131  & ~n4141 ;
  assign n8941 = ~n4119 & n8940 ;
  assign n8942 = ~n8939 & ~n8941 ;
  assign n8948 = ~n4152 & ~n8942 ;
  assign n8949 = ~n8947 & ~n8948 ;
  assign n8950 = n952 & ~n8949 ;
  assign n8951 = ~n600 & n4141 ;
  assign n8952 = ~n8940 & ~n8951 ;
  assign n8953 = n993 & ~n8952 ;
  assign n8943 = n970 & ~n8942 ;
  assign n8954 = \InstQueue_reg[4][1]/NET0131  & ~n3933 ;
  assign n8955 = ~n8943 & ~n8954 ;
  assign n8956 = ~n8953 & n8955 ;
  assign n8957 = ~n8950 & n8956 ;
  assign n8963 = n4097 & n8709 ;
  assign n8964 = n4119 & n8712 ;
  assign n8965 = ~n8963 & ~n8964 ;
  assign n8966 = \DataWidth_reg[1]/NET0131  & ~n8965 ;
  assign n8958 = \Datai[1]_pad  & ~n4164 ;
  assign n8959 = \InstQueue_reg[5][1]/NET0131  & ~n4163 ;
  assign n8960 = ~n4141 & n8959 ;
  assign n8961 = ~n8958 & ~n8960 ;
  assign n8967 = ~n4174 & ~n8961 ;
  assign n8968 = ~n8966 & ~n8967 ;
  assign n8969 = n952 & ~n8968 ;
  assign n8970 = ~n600 & n4163 ;
  assign n8971 = ~n8959 & ~n8970 ;
  assign n8972 = n993 & ~n8971 ;
  assign n8962 = n970 & ~n8961 ;
  assign n8973 = \InstQueue_reg[5][1]/NET0131  & ~n3933 ;
  assign n8974 = ~n8962 & ~n8973 ;
  assign n8975 = ~n8972 & n8974 ;
  assign n8976 = ~n8969 & n8975 ;
  assign n8982 = n4119 & n8709 ;
  assign n8983 = n4141 & n8712 ;
  assign n8984 = ~n8982 & ~n8983 ;
  assign n8985 = \DataWidth_reg[1]/NET0131  & ~n8984 ;
  assign n8977 = \Datai[1]_pad  & ~n4186 ;
  assign n8978 = \InstQueue_reg[6][1]/NET0131  & ~n4185 ;
  assign n8979 = ~n4163 & n8978 ;
  assign n8980 = ~n8977 & ~n8979 ;
  assign n8986 = ~n4196 & ~n8980 ;
  assign n8987 = ~n8985 & ~n8986 ;
  assign n8988 = n952 & ~n8987 ;
  assign n8989 = ~n600 & n4185 ;
  assign n8990 = ~n8978 & ~n8989 ;
  assign n8991 = n993 & ~n8990 ;
  assign n8981 = n970 & ~n8980 ;
  assign n8992 = \InstQueue_reg[6][1]/NET0131  & ~n3933 ;
  assign n8993 = ~n8981 & ~n8992 ;
  assign n8994 = ~n8991 & n8993 ;
  assign n8995 = ~n8988 & n8994 ;
  assign n9001 = n4141 & n8751 ;
  assign n9002 = n4163 & n8754 ;
  assign n9003 = ~n9001 & ~n9002 ;
  assign n9004 = \DataWidth_reg[1]/NET0131  & ~n9003 ;
  assign n8996 = \Datai[0]_pad  & ~n4207 ;
  assign n8997 = \InstQueue_reg[7][0]/NET0131  & ~n3948 ;
  assign n8998 = ~n4185 & n8997 ;
  assign n8999 = ~n8996 & ~n8998 ;
  assign n9005 = ~n4217 & ~n8999 ;
  assign n9006 = ~n9004 & ~n9005 ;
  assign n9007 = n952 & ~n9006 ;
  assign n9008 = ~n663 & n3948 ;
  assign n9009 = ~n8997 & ~n9008 ;
  assign n9010 = n993 & ~n9009 ;
  assign n9000 = n970 & ~n8999 ;
  assign n9011 = \InstQueue_reg[7][0]/NET0131  & ~n3933 ;
  assign n9012 = ~n9000 & ~n9011 ;
  assign n9013 = ~n9010 & n9012 ;
  assign n9014 = ~n9007 & n9013 ;
  assign n9020 = n4141 & n8709 ;
  assign n9021 = n4163 & n8712 ;
  assign n9022 = ~n9020 & ~n9021 ;
  assign n9023 = \DataWidth_reg[1]/NET0131  & ~n9022 ;
  assign n9015 = \Datai[1]_pad  & ~n4207 ;
  assign n9016 = \InstQueue_reg[7][1]/NET0131  & ~n3948 ;
  assign n9017 = ~n4185 & n9016 ;
  assign n9018 = ~n9015 & ~n9017 ;
  assign n9024 = ~n4217 & ~n9018 ;
  assign n9025 = ~n9023 & ~n9024 ;
  assign n9026 = n952 & ~n9025 ;
  assign n9027 = ~n600 & n3948 ;
  assign n9028 = ~n9016 & ~n9027 ;
  assign n9029 = n993 & ~n9028 ;
  assign n9019 = n970 & ~n9018 ;
  assign n9030 = \InstQueue_reg[7][1]/NET0131  & ~n3933 ;
  assign n9031 = ~n9019 & ~n9030 ;
  assign n9032 = ~n9029 & n9031 ;
  assign n9033 = ~n9026 & n9032 ;
  assign n9039 = n4163 & n8709 ;
  assign n9040 = n4185 & n8712 ;
  assign n9041 = ~n9039 & ~n9040 ;
  assign n9042 = \DataWidth_reg[1]/NET0131  & ~n9041 ;
  assign n9034 = \Datai[1]_pad  & ~n3954 ;
  assign n9035 = \InstQueue_reg[8][1]/NET0131  & ~n3950 ;
  assign n9036 = ~n3948 & n9035 ;
  assign n9037 = ~n9034 & ~n9036 ;
  assign n9043 = ~n4237 & ~n9037 ;
  assign n9044 = ~n9042 & ~n9043 ;
  assign n9045 = n952 & ~n9044 ;
  assign n9046 = ~n600 & n3950 ;
  assign n9047 = ~n9035 & ~n9046 ;
  assign n9048 = n993 & ~n9047 ;
  assign n9038 = n970 & ~n9037 ;
  assign n9049 = \InstQueue_reg[8][1]/NET0131  & ~n3933 ;
  assign n9050 = ~n9038 & ~n9049 ;
  assign n9051 = ~n9048 & n9050 ;
  assign n9052 = ~n9045 & n9051 ;
  assign n9058 = n4185 & n8709 ;
  assign n9059 = n3948 & n8712 ;
  assign n9060 = ~n9058 & ~n9059 ;
  assign n9061 = \DataWidth_reg[1]/NET0131  & ~n9060 ;
  assign n9053 = \Datai[1]_pad  & ~n3978 ;
  assign n9054 = \InstQueue_reg[9][1]/NET0131  & ~n3941 ;
  assign n9055 = ~n3950 & n9054 ;
  assign n9056 = ~n9053 & ~n9055 ;
  assign n9062 = ~n4257 & ~n9056 ;
  assign n9063 = ~n9061 & ~n9062 ;
  assign n9064 = n952 & ~n9063 ;
  assign n9065 = ~n600 & n3941 ;
  assign n9066 = ~n9054 & ~n9065 ;
  assign n9067 = n993 & ~n9066 ;
  assign n9057 = n970 & ~n9056 ;
  assign n9068 = \InstQueue_reg[9][1]/NET0131  & ~n3933 ;
  assign n9069 = ~n9057 & ~n9068 ;
  assign n9070 = ~n9067 & n9069 ;
  assign n9071 = ~n9064 & n9070 ;
  assign n9078 = ~\rEIP_reg[26]/NET0131  & ~n8466 ;
  assign n9079 = n830 & ~n8467 ;
  assign n9080 = ~n9078 & n9079 ;
  assign n9072 = \Address[24]_pad  & ~n829 ;
  assign n9075 = n6016 & n8439 ;
  assign n9073 = n5977 & n8439 ;
  assign n9074 = ~\rEIP_reg[25]/NET0131  & ~n9073 ;
  assign n9076 = n8438 & ~n9074 ;
  assign n9077 = ~n9075 & n9076 ;
  assign n9081 = ~n9072 & ~n9077 ;
  assign n9082 = ~n9080 & n9081 ;
  assign n9089 = ~\rEIP_reg[14]/NET0131  & ~n8460 ;
  assign n9090 = n830 & ~n8461 ;
  assign n9091 = ~n9089 & n9090 ;
  assign n9083 = \Address[12]_pad  & ~n829 ;
  assign n9086 = n4664 & n8439 ;
  assign n9084 = n4663 & n8439 ;
  assign n9085 = ~\rEIP_reg[13]/NET0131  & ~n9084 ;
  assign n9087 = n8438 & ~n9085 ;
  assign n9088 = ~n9086 & n9087 ;
  assign n9092 = ~n9083 & ~n9088 ;
  assign n9093 = ~n9091 & n9092 ;
  assign n9102 = ~\rEIP_reg[22]/NET0131  & ~n8464 ;
  assign n9101 = \rEIP_reg[22]/NET0131  & n8464 ;
  assign n9103 = n830 & ~n9101 ;
  assign n9104 = ~n9102 & n9103 ;
  assign n9094 = \Address[20]_pad  & ~n829 ;
  assign n9095 = n5836 & n8439 ;
  assign n9096 = \rEIP_reg[20]/NET0131  & n9095 ;
  assign n9097 = ~\rEIP_reg[21]/NET0131  & ~n9096 ;
  assign n9098 = n4672 & n8439 ;
  assign n9099 = n8438 & ~n9098 ;
  assign n9100 = ~n9097 & n9099 ;
  assign n9105 = ~n9094 & ~n9100 ;
  assign n9106 = ~n9104 & n9105 ;
  assign n9115 = ~\rEIP_reg[10]/NET0131  & ~n8456 ;
  assign n9116 = n830 & ~n8457 ;
  assign n9117 = ~n9115 & n9116 ;
  assign n9107 = \Address[8]_pad  & ~n829 ;
  assign n9108 = n4657 & n8439 ;
  assign n9109 = \rEIP_reg[7]/NET0131  & n9108 ;
  assign n9110 = \rEIP_reg[8]/NET0131  & n9109 ;
  assign n9112 = ~\rEIP_reg[9]/NET0131  & ~n9110 ;
  assign n9111 = \rEIP_reg[9]/NET0131  & n9110 ;
  assign n9113 = n8438 & ~n9111 ;
  assign n9114 = ~n9112 & n9113 ;
  assign n9118 = ~n9107 & ~n9114 ;
  assign n9119 = ~n9117 & n9118 ;
  assign n9125 = n3876 & n8751 ;
  assign n9126 = n3919 & n8754 ;
  assign n9127 = ~n9125 & ~n9126 ;
  assign n9128 = \DataWidth_reg[1]/NET0131  & ~n9127 ;
  assign n9120 = \Datai[0]_pad  & ~n3868 ;
  assign n9121 = \InstQueue_reg[0][0]/NET0131  & ~n3864 ;
  assign n9122 = ~n3867 & n9121 ;
  assign n9123 = ~n9120 & ~n9122 ;
  assign n9129 = ~n3924 & ~n9123 ;
  assign n9130 = ~n9128 & ~n9129 ;
  assign n9131 = n952 & ~n9130 ;
  assign n9132 = ~n663 & n3864 ;
  assign n9133 = ~n9121 & ~n9132 ;
  assign n9134 = n993 & ~n9133 ;
  assign n9124 = n970 & ~n9123 ;
  assign n9135 = \InstQueue_reg[0][0]/NET0131  & ~n3933 ;
  assign n9136 = ~n9124 & ~n9135 ;
  assign n9137 = ~n9134 & n9136 ;
  assign n9138 = ~n9131 & n9137 ;
  assign n9144 = n3950 & n8754 ;
  assign n9145 = n3948 & n8751 ;
  assign n9146 = ~n9144 & ~n9145 ;
  assign n9147 = \DataWidth_reg[1]/NET0131  & ~n9146 ;
  assign n9139 = \Datai[0]_pad  & ~n3942 ;
  assign n9140 = \InstQueue_reg[10][0]/NET0131  & ~n3939 ;
  assign n9141 = ~n3941 & n9140 ;
  assign n9142 = ~n9139 & ~n9141 ;
  assign n9148 = ~n3955 & ~n9142 ;
  assign n9149 = ~n9147 & ~n9148 ;
  assign n9150 = n952 & ~n9149 ;
  assign n9151 = ~n663 & n3939 ;
  assign n9152 = ~n9140 & ~n9151 ;
  assign n9153 = n993 & ~n9152 ;
  assign n9143 = n970 & ~n9142 ;
  assign n9154 = \InstQueue_reg[10][0]/NET0131  & ~n3933 ;
  assign n9155 = ~n9143 & ~n9154 ;
  assign n9156 = ~n9153 & n9155 ;
  assign n9157 = ~n9150 & n9156 ;
  assign n9163 = n3941 & n8751 ;
  assign n9164 = n3939 & n8754 ;
  assign n9165 = ~n9163 & ~n9164 ;
  assign n9166 = \DataWidth_reg[1]/NET0131  & ~n9165 ;
  assign n9158 = \Datai[0]_pad  & ~n3992 ;
  assign n9159 = \InstQueue_reg[12][0]/NET0131  & ~n3991 ;
  assign n9160 = ~n3967 & n9159 ;
  assign n9161 = ~n9158 & ~n9160 ;
  assign n9167 = ~n4002 & ~n9161 ;
  assign n9168 = ~n9166 & ~n9167 ;
  assign n9169 = n952 & ~n9168 ;
  assign n9170 = ~n663 & n3991 ;
  assign n9171 = ~n9159 & ~n9170 ;
  assign n9172 = n993 & ~n9171 ;
  assign n9162 = n970 & ~n9161 ;
  assign n9173 = \InstQueue_reg[12][0]/NET0131  & ~n3933 ;
  assign n9174 = ~n9162 & ~n9173 ;
  assign n9175 = ~n9172 & n9174 ;
  assign n9176 = ~n9169 & n9175 ;
  assign n9182 = n3939 & n8751 ;
  assign n9183 = n3967 & n8754 ;
  assign n9184 = ~n9182 & ~n9183 ;
  assign n9185 = \DataWidth_reg[1]/NET0131  & ~n9184 ;
  assign n9177 = \Datai[0]_pad  & ~n4013 ;
  assign n9178 = \InstQueue_reg[13][0]/NET0131  & ~n3876 ;
  assign n9179 = ~n3991 & n9178 ;
  assign n9180 = ~n9177 & ~n9179 ;
  assign n9186 = ~n4023 & ~n9180 ;
  assign n9187 = ~n9185 & ~n9186 ;
  assign n9188 = n952 & ~n9187 ;
  assign n9189 = ~n663 & n3876 ;
  assign n9190 = ~n9178 & ~n9189 ;
  assign n9191 = n993 & ~n9190 ;
  assign n9181 = n970 & ~n9180 ;
  assign n9192 = \InstQueue_reg[13][0]/NET0131  & ~n3933 ;
  assign n9193 = ~n9181 & ~n9192 ;
  assign n9194 = ~n9191 & n9193 ;
  assign n9195 = ~n9188 & n9194 ;
  assign n9201 = n3967 & n8751 ;
  assign n9202 = n3991 & n8754 ;
  assign n9203 = ~n9201 & ~n9202 ;
  assign n9204 = \DataWidth_reg[1]/NET0131  & ~n9203 ;
  assign n9196 = \Datai[0]_pad  & ~n3923 ;
  assign n9197 = \InstQueue_reg[14][0]/NET0131  & ~n3919 ;
  assign n9198 = ~n3876 & n9197 ;
  assign n9199 = ~n9196 & ~n9198 ;
  assign n9205 = ~n4043 & ~n9199 ;
  assign n9206 = ~n9204 & ~n9205 ;
  assign n9207 = n952 & ~n9206 ;
  assign n9208 = ~n663 & n3919 ;
  assign n9209 = ~n9197 & ~n9208 ;
  assign n9210 = n993 & ~n9209 ;
  assign n9200 = n970 & ~n9199 ;
  assign n9211 = \InstQueue_reg[14][0]/NET0131  & ~n3933 ;
  assign n9212 = ~n9200 & ~n9211 ;
  assign n9213 = ~n9210 & n9212 ;
  assign n9214 = ~n9207 & n9213 ;
  assign n9220 = n3991 & n8751 ;
  assign n9221 = n3876 & n8754 ;
  assign n9222 = ~n9220 & ~n9221 ;
  assign n9223 = \DataWidth_reg[1]/NET0131  & ~n9222 ;
  assign n9215 = \Datai[0]_pad  & ~n4054 ;
  assign n9216 = \InstQueue_reg[15][0]/NET0131  & ~n3867 ;
  assign n9217 = ~n3919 & n9216 ;
  assign n9218 = ~n9215 & ~n9217 ;
  assign n9224 = ~n4064 & ~n9218 ;
  assign n9225 = ~n9223 & ~n9224 ;
  assign n9226 = n952 & ~n9225 ;
  assign n9227 = ~n663 & n3867 ;
  assign n9228 = ~n9216 & ~n9227 ;
  assign n9229 = n993 & ~n9228 ;
  assign n9219 = n970 & ~n9218 ;
  assign n9230 = \InstQueue_reg[15][0]/NET0131  & ~n3933 ;
  assign n9231 = ~n9219 & ~n9230 ;
  assign n9232 = ~n9229 & n9231 ;
  assign n9233 = ~n9226 & n9232 ;
  assign n9239 = n3919 & n8751 ;
  assign n9240 = n3867 & n8754 ;
  assign n9241 = ~n9239 & ~n9240 ;
  assign n9242 = \DataWidth_reg[1]/NET0131  & ~n9241 ;
  assign n9234 = \Datai[0]_pad  & ~n4076 ;
  assign n9235 = \InstQueue_reg[1][0]/NET0131  & ~n4075 ;
  assign n9236 = ~n3864 & n9235 ;
  assign n9237 = ~n9234 & ~n9236 ;
  assign n9243 = ~n4086 & ~n9237 ;
  assign n9244 = ~n9242 & ~n9243 ;
  assign n9245 = n952 & ~n9244 ;
  assign n9246 = ~n663 & n4075 ;
  assign n9247 = ~n9235 & ~n9246 ;
  assign n9248 = n993 & ~n9247 ;
  assign n9238 = n970 & ~n9237 ;
  assign n9249 = \InstQueue_reg[1][0]/NET0131  & ~n3933 ;
  assign n9250 = ~n9238 & ~n9249 ;
  assign n9251 = ~n9248 & n9250 ;
  assign n9252 = ~n9245 & n9251 ;
  assign n9258 = n3864 & n8754 ;
  assign n9259 = n3867 & n8751 ;
  assign n9260 = ~n9258 & ~n9259 ;
  assign n9261 = \DataWidth_reg[1]/NET0131  & ~n9260 ;
  assign n9253 = \Datai[0]_pad  & ~n4098 ;
  assign n9254 = \InstQueue_reg[2][0]/NET0131  & ~n4097 ;
  assign n9255 = ~n4075 & n9254 ;
  assign n9256 = ~n9253 & ~n9255 ;
  assign n9262 = ~n4108 & ~n9256 ;
  assign n9263 = ~n9261 & ~n9262 ;
  assign n9264 = n952 & ~n9263 ;
  assign n9265 = ~n663 & n4097 ;
  assign n9266 = ~n9254 & ~n9265 ;
  assign n9267 = n993 & ~n9266 ;
  assign n9257 = n970 & ~n9256 ;
  assign n9268 = \InstQueue_reg[2][0]/NET0131  & ~n3933 ;
  assign n9269 = ~n9257 & ~n9268 ;
  assign n9270 = ~n9267 & n9269 ;
  assign n9271 = ~n9264 & n9270 ;
  assign n9277 = n4075 & n8751 ;
  assign n9278 = n4097 & n8754 ;
  assign n9279 = ~n9277 & ~n9278 ;
  assign n9280 = \DataWidth_reg[1]/NET0131  & ~n9279 ;
  assign n9272 = \Datai[0]_pad  & ~n4142 ;
  assign n9273 = \InstQueue_reg[4][0]/NET0131  & ~n4141 ;
  assign n9274 = ~n4119 & n9273 ;
  assign n9275 = ~n9272 & ~n9274 ;
  assign n9281 = ~n4152 & ~n9275 ;
  assign n9282 = ~n9280 & ~n9281 ;
  assign n9283 = n952 & ~n9282 ;
  assign n9284 = ~n663 & n4141 ;
  assign n9285 = ~n9273 & ~n9284 ;
  assign n9286 = n993 & ~n9285 ;
  assign n9276 = n970 & ~n9275 ;
  assign n9287 = \InstQueue_reg[4][0]/NET0131  & ~n3933 ;
  assign n9288 = ~n9276 & ~n9287 ;
  assign n9289 = ~n9286 & n9288 ;
  assign n9290 = ~n9283 & n9289 ;
  assign n9296 = n4097 & n8751 ;
  assign n9297 = n4119 & n8754 ;
  assign n9298 = ~n9296 & ~n9297 ;
  assign n9299 = \DataWidth_reg[1]/NET0131  & ~n9298 ;
  assign n9291 = \Datai[0]_pad  & ~n4164 ;
  assign n9292 = \InstQueue_reg[5][0]/NET0131  & ~n4163 ;
  assign n9293 = ~n4141 & n9292 ;
  assign n9294 = ~n9291 & ~n9293 ;
  assign n9300 = ~n4174 & ~n9294 ;
  assign n9301 = ~n9299 & ~n9300 ;
  assign n9302 = n952 & ~n9301 ;
  assign n9303 = ~n663 & n4163 ;
  assign n9304 = ~n9292 & ~n9303 ;
  assign n9305 = n993 & ~n9304 ;
  assign n9295 = n970 & ~n9294 ;
  assign n9306 = \InstQueue_reg[5][0]/NET0131  & ~n3933 ;
  assign n9307 = ~n9295 & ~n9306 ;
  assign n9308 = ~n9305 & n9307 ;
  assign n9309 = ~n9302 & n9308 ;
  assign n9315 = n4119 & n8751 ;
  assign n9316 = n4141 & n8754 ;
  assign n9317 = ~n9315 & ~n9316 ;
  assign n9318 = \DataWidth_reg[1]/NET0131  & ~n9317 ;
  assign n9310 = \Datai[0]_pad  & ~n4186 ;
  assign n9311 = \InstQueue_reg[6][0]/NET0131  & ~n4185 ;
  assign n9312 = ~n4163 & n9311 ;
  assign n9313 = ~n9310 & ~n9312 ;
  assign n9319 = ~n4196 & ~n9313 ;
  assign n9320 = ~n9318 & ~n9319 ;
  assign n9321 = n952 & ~n9320 ;
  assign n9322 = ~n663 & n4185 ;
  assign n9323 = ~n9311 & ~n9322 ;
  assign n9324 = n993 & ~n9323 ;
  assign n9314 = n970 & ~n9313 ;
  assign n9325 = \InstQueue_reg[6][0]/NET0131  & ~n3933 ;
  assign n9326 = ~n9314 & ~n9325 ;
  assign n9327 = ~n9324 & n9326 ;
  assign n9328 = ~n9321 & n9327 ;
  assign n9334 = n4163 & n8751 ;
  assign n9335 = n4185 & n8754 ;
  assign n9336 = ~n9334 & ~n9335 ;
  assign n9337 = \DataWidth_reg[1]/NET0131  & ~n9336 ;
  assign n9329 = \Datai[0]_pad  & ~n3954 ;
  assign n9330 = \InstQueue_reg[8][0]/NET0131  & ~n3950 ;
  assign n9331 = ~n3948 & n9330 ;
  assign n9332 = ~n9329 & ~n9331 ;
  assign n9338 = ~n4237 & ~n9332 ;
  assign n9339 = ~n9337 & ~n9338 ;
  assign n9340 = n952 & ~n9339 ;
  assign n9341 = ~n663 & n3950 ;
  assign n9342 = ~n9330 & ~n9341 ;
  assign n9343 = n993 & ~n9342 ;
  assign n9333 = n970 & ~n9332 ;
  assign n9344 = \InstQueue_reg[8][0]/NET0131  & ~n3933 ;
  assign n9345 = ~n9333 & ~n9344 ;
  assign n9346 = ~n9343 & n9345 ;
  assign n9347 = ~n9340 & n9346 ;
  assign n9353 = n4185 & n8751 ;
  assign n9354 = n3948 & n8754 ;
  assign n9355 = ~n9353 & ~n9354 ;
  assign n9356 = \DataWidth_reg[1]/NET0131  & ~n9355 ;
  assign n9348 = \Datai[0]_pad  & ~n3978 ;
  assign n9349 = \InstQueue_reg[9][0]/NET0131  & ~n3941 ;
  assign n9350 = ~n3950 & n9349 ;
  assign n9351 = ~n9348 & ~n9350 ;
  assign n9357 = ~n4257 & ~n9351 ;
  assign n9358 = ~n9356 & ~n9357 ;
  assign n9359 = n952 & ~n9358 ;
  assign n9360 = ~n663 & n3941 ;
  assign n9361 = ~n9349 & ~n9360 ;
  assign n9362 = n993 & ~n9361 ;
  assign n9352 = n970 & ~n9351 ;
  assign n9363 = \InstQueue_reg[9][0]/NET0131  & ~n3933 ;
  assign n9364 = ~n9352 & ~n9363 ;
  assign n9365 = ~n9362 & n9364 ;
  assign n9366 = ~n9359 & n9365 ;
  assign n9376 = ~\rEIP_reg[6]/NET0131  & ~n8452 ;
  assign n9377 = n830 & ~n8453 ;
  assign n9378 = ~n9376 & n9377 ;
  assign n9367 = \Address[4]_pad  & ~n829 ;
  assign n9368 = \rEIP_reg[1]/NET0131  & n8439 ;
  assign n9369 = \rEIP_reg[2]/NET0131  & n9368 ;
  assign n9370 = \rEIP_reg[3]/NET0131  & n9369 ;
  assign n9371 = \rEIP_reg[4]/NET0131  & n9370 ;
  assign n9373 = ~\rEIP_reg[5]/NET0131  & ~n9371 ;
  assign n9372 = \rEIP_reg[5]/NET0131  & n9371 ;
  assign n9374 = n8438 & ~n9372 ;
  assign n9375 = ~n9373 & n9374 ;
  assign n9379 = ~n9367 & ~n9375 ;
  assign n9380 = ~n9378 & n9379 ;
  assign n9386 = n4677 & n8467 ;
  assign n9387 = ~\rEIP_reg[29]/NET0131  & ~n9386 ;
  assign n9388 = n830 & ~n8468 ;
  assign n9389 = ~n9387 & n9388 ;
  assign n9381 = \Address[27]_pad  & ~n829 ;
  assign n9382 = \rEIP_reg[27]/NET0131  & n8441 ;
  assign n9383 = ~\rEIP_reg[28]/NET0131  & ~n9382 ;
  assign n9384 = n8438 & ~n8442 ;
  assign n9385 = ~n9383 & n9384 ;
  assign n9390 = ~n9381 & ~n9385 ;
  assign n9391 = ~n9389 & n9390 ;
  assign n9392 = ~\Address[15]_pad  & ~n829 ;
  assign n9396 = ~\rEIP_reg[17]/NET0131  & ~n8463 ;
  assign n9397 = ~\State_reg[2]/NET0131  & ~n8537 ;
  assign n9398 = ~n9396 & n9397 ;
  assign n9393 = ~\rEIP_reg[16]/NET0131  & ~n8531 ;
  assign n9394 = \State_reg[2]/NET0131  & ~n8532 ;
  assign n9395 = ~n9393 & n9394 ;
  assign n9399 = n829 & ~n9395 ;
  assign n9400 = ~n9398 & n9399 ;
  assign n9401 = ~n9392 & ~n9400 ;
  assign n9406 = \rEIP_reg[24]/NET0131  & n8465 ;
  assign n9407 = ~\rEIP_reg[25]/NET0131  & ~n9406 ;
  assign n9408 = n830 & ~n8466 ;
  assign n9409 = ~n9407 & n9408 ;
  assign n9402 = \Address[23]_pad  & ~n829 ;
  assign n9403 = ~\rEIP_reg[24]/NET0131  & ~n8440 ;
  assign n9404 = n8438 & ~n9073 ;
  assign n9405 = ~n9403 & n9404 ;
  assign n9410 = ~n9402 & ~n9405 ;
  assign n9411 = ~n9409 & n9410 ;
  assign n9417 = ~\rEIP_reg[13]/NET0131  & ~n8459 ;
  assign n9418 = n830 & ~n8460 ;
  assign n9419 = ~n9417 & n9418 ;
  assign n9412 = \Address[11]_pad  & ~n829 ;
  assign n9414 = ~n6585 & n8439 ;
  assign n9413 = ~\rEIP_reg[12]/NET0131  & ~n8439 ;
  assign n9415 = n8438 & ~n9413 ;
  assign n9416 = ~n9414 & n9415 ;
  assign n9420 = ~n9412 & ~n9416 ;
  assign n9421 = ~n9419 & n9420 ;
  assign n9426 = ~\rEIP_reg[5]/NET0131  & ~n8451 ;
  assign n9427 = n830 & ~n8452 ;
  assign n9428 = ~n9426 & n9427 ;
  assign n9422 = \Address[3]_pad  & ~n829 ;
  assign n9423 = ~\rEIP_reg[4]/NET0131  & ~n9370 ;
  assign n9424 = n8438 & ~n9371 ;
  assign n9425 = ~n9423 & n9424 ;
  assign n9429 = ~n9422 & ~n9425 ;
  assign n9430 = ~n9428 & n9429 ;
  assign n9435 = \rEIP_reg[19]/NET0131  & n8539 ;
  assign n9436 = \rEIP_reg[20]/NET0131  & n9435 ;
  assign n9437 = ~\rEIP_reg[21]/NET0131  & ~n9436 ;
  assign n9438 = n830 & ~n8464 ;
  assign n9439 = ~n9437 & n9438 ;
  assign n9431 = \Address[19]_pad  & ~n829 ;
  assign n9432 = ~\rEIP_reg[20]/NET0131  & ~n9095 ;
  assign n9433 = n8438 & ~n9096 ;
  assign n9434 = ~n9432 & n9433 ;
  assign n9440 = ~n9431 & ~n9434 ;
  assign n9441 = ~n9439 & n9440 ;
  assign n9446 = ~\rEIP_reg[9]/NET0131  & ~n8455 ;
  assign n9447 = n830 & ~n8456 ;
  assign n9448 = ~n9446 & n9447 ;
  assign n9442 = \Address[7]_pad  & ~n829 ;
  assign n9443 = ~\rEIP_reg[8]/NET0131  & ~n9109 ;
  assign n9444 = n8438 & ~n9110 ;
  assign n9445 = ~n9443 & n9444 ;
  assign n9449 = ~n9442 & ~n9445 ;
  assign n9450 = ~n9448 & n9449 ;
  assign n9455 = ~\rEIP_reg[16]/NET0131  & ~n8462 ;
  assign n9456 = n830 & ~n8463 ;
  assign n9457 = ~n9455 & n9456 ;
  assign n9451 = \Address[14]_pad  & ~n829 ;
  assign n9452 = ~\rEIP_reg[15]/NET0131  & ~n8530 ;
  assign n9453 = n8438 & ~n8531 ;
  assign n9454 = ~n9452 & n9453 ;
  assign n9458 = ~n9451 & ~n9454 ;
  assign n9459 = ~n9457 & n9458 ;
  assign n9464 = \rEIP_reg[27]/NET0131  & n8467 ;
  assign n9465 = ~\rEIP_reg[28]/NET0131  & ~n9464 ;
  assign n9466 = n830 & ~n9386 ;
  assign n9467 = ~n9465 & n9466 ;
  assign n9460 = \Address[26]_pad  & ~n829 ;
  assign n9461 = ~\rEIP_reg[27]/NET0131  & ~n8441 ;
  assign n9462 = n8438 & ~n9382 ;
  assign n9463 = ~n9461 & n9462 ;
  assign n9468 = ~n9460 & ~n9463 ;
  assign n9469 = ~n9467 & n9468 ;
  assign n9475 = ~\rEIP_reg[24]/NET0131  & ~n8465 ;
  assign n9476 = n830 & ~n9406 ;
  assign n9477 = ~n9475 & n9476 ;
  assign n9470 = \Address[22]_pad  & ~n829 ;
  assign n9471 = n5910 & n8439 ;
  assign n9472 = ~\rEIP_reg[23]/NET0131  & ~n9471 ;
  assign n9473 = n8438 & ~n8440 ;
  assign n9474 = ~n9472 & n9473 ;
  assign n9478 = ~n9470 & ~n9474 ;
  assign n9479 = ~n9477 & n9478 ;
  assign n9485 = ~\rEIP_reg[12]/NET0131  & ~n8458 ;
  assign n9486 = n830 & ~n8459 ;
  assign n9487 = ~n9485 & n9486 ;
  assign n9480 = \Address[10]_pad  & ~n829 ;
  assign n9482 = ~n6548 & n8439 ;
  assign n9481 = ~\rEIP_reg[11]/NET0131  & ~n8439 ;
  assign n9483 = n8438 & ~n9481 ;
  assign n9484 = ~n9482 & n9483 ;
  assign n9488 = ~n9480 & ~n9484 ;
  assign n9489 = ~n9487 & n9488 ;
  assign n9494 = ~\rEIP_reg[4]/NET0131  & ~n8450 ;
  assign n9495 = n830 & ~n8451 ;
  assign n9496 = ~n9494 & n9495 ;
  assign n9490 = \Address[2]_pad  & ~n829 ;
  assign n9491 = ~\rEIP_reg[3]/NET0131  & ~n9369 ;
  assign n9492 = n8438 & ~n9370 ;
  assign n9493 = ~n9491 & n9492 ;
  assign n9497 = ~n9490 & ~n9493 ;
  assign n9498 = ~n9496 & n9497 ;
  assign n9504 = ~\rEIP_reg[20]/NET0131  & ~n9435 ;
  assign n9505 = n830 & ~n9436 ;
  assign n9506 = ~n9504 & n9505 ;
  assign n9499 = \Address[18]_pad  & ~n829 ;
  assign n9500 = \rEIP_reg[18]/NET0131  & n8533 ;
  assign n9501 = ~\rEIP_reg[19]/NET0131  & ~n9500 ;
  assign n9502 = n8438 & ~n9095 ;
  assign n9503 = ~n9501 & n9502 ;
  assign n9507 = ~n9499 & ~n9503 ;
  assign n9508 = ~n9506 & n9507 ;
  assign n9513 = ~\rEIP_reg[8]/NET0131  & ~n8454 ;
  assign n9514 = n830 & ~n8455 ;
  assign n9515 = ~n9513 & n9514 ;
  assign n9509 = \Address[6]_pad  & ~n829 ;
  assign n9510 = ~\rEIP_reg[7]/NET0131  & ~n9108 ;
  assign n9511 = n8438 & ~n9109 ;
  assign n9512 = ~n9510 & n9511 ;
  assign n9516 = ~n9509 & ~n9512 ;
  assign n9517 = ~n9515 & n9516 ;
  assign n9522 = ~\rEIP_reg[27]/NET0131  & ~n8467 ;
  assign n9523 = n830 & ~n9464 ;
  assign n9524 = ~n9522 & n9523 ;
  assign n9518 = \Address[25]_pad  & ~n829 ;
  assign n9519 = ~\rEIP_reg[26]/NET0131  & ~n9075 ;
  assign n9520 = n8438 & ~n8441 ;
  assign n9521 = ~n9519 & n9520 ;
  assign n9525 = ~n9518 & ~n9521 ;
  assign n9526 = ~n9524 & n9525 ;
  assign n9533 = \rEIP_reg[31]/NET0131  & n8470 ;
  assign n9532 = ~\rEIP_reg[31]/NET0131  & ~n8470 ;
  assign n9534 = n830 & ~n9532 ;
  assign n9535 = ~n9533 & n9534 ;
  assign n9527 = \Address[29]_pad  & ~n829 ;
  assign n9529 = \rEIP_reg[0]/NET0131  & n4681 ;
  assign n9528 = ~\rEIP_reg[30]/NET0131  & ~n8444 ;
  assign n9530 = n8438 & ~n9528 ;
  assign n9531 = ~n9529 & n9530 ;
  assign n9536 = ~n9527 & ~n9531 ;
  assign n9537 = ~n9535 & n9536 ;
  assign n9542 = ~\rEIP_reg[15]/NET0131  & ~n8461 ;
  assign n9543 = n830 & ~n8462 ;
  assign n9544 = ~n9542 & n9543 ;
  assign n9538 = \Address[13]_pad  & ~n829 ;
  assign n9539 = ~\rEIP_reg[14]/NET0131  & ~n9086 ;
  assign n9540 = n8438 & ~n8530 ;
  assign n9541 = ~n9539 & n9540 ;
  assign n9545 = ~n9538 & ~n9541 ;
  assign n9546 = ~n9544 & n9545 ;
  assign n9552 = ~\rEIP_reg[11]/NET0131  & ~n8457 ;
  assign n9553 = n830 & ~n8458 ;
  assign n9554 = ~n9552 & n9553 ;
  assign n9547 = \Address[9]_pad  & ~n829 ;
  assign n9549 = \rEIP_reg[10]/NET0131  & n9111 ;
  assign n9548 = ~\rEIP_reg[10]/NET0131  & ~n9111 ;
  assign n9550 = n8438 & ~n9548 ;
  assign n9551 = ~n9549 & n9550 ;
  assign n9555 = ~n9547 & ~n9551 ;
  assign n9556 = ~n9554 & n9555 ;
  assign n9561 = ~\rEIP_reg[23]/NET0131  & ~n9101 ;
  assign n9562 = n830 & ~n8465 ;
  assign n9563 = ~n9561 & n9562 ;
  assign n9557 = \Address[21]_pad  & ~n829 ;
  assign n9558 = ~\rEIP_reg[22]/NET0131  & ~n9098 ;
  assign n9559 = n8438 & ~n9471 ;
  assign n9560 = ~n9558 & n9559 ;
  assign n9564 = ~n9557 & ~n9560 ;
  assign n9565 = ~n9563 & n9564 ;
  assign n9566 = \DataWidth_reg[0]/NET0131  & \DataWidth_reg[1]/NET0131  ;
  assign n9567 = \ByteEnable_reg[2]/NET0131  & n9566 ;
  assign n9568 = ~\DataWidth_reg[1]/NET0131  & \rEIP_reg[1]/NET0131  ;
  assign n9569 = \DataWidth_reg[0]/NET0131  & ~n9568 ;
  assign n9570 = \rEIP_reg[0]/NET0131  & ~n9569 ;
  assign n9571 = ~n8447 & ~n9570 ;
  assign n9572 = ~n5822 & ~n9571 ;
  assign n9573 = ~n9567 & ~n9572 ;
  assign n9577 = ~HOLD_pad & \State_reg[0]/NET0131  ;
  assign n9578 = ~\State_reg[2]/NET0131  & ~n9577 ;
  assign n9579 = ~READY_n_pad & ~n9578 ;
  assign n9580 = \State_reg[1]/NET0131  & ~n9579 ;
  assign n9574 = HOLD_pad & \State_reg[2]/NET0131  ;
  assign n9575 = \RequestPending_reg/NET0131  & \State_reg[0]/NET0131  ;
  assign n9576 = ~n9574 & n9575 ;
  assign n9581 = ~n832 & ~n9576 ;
  assign n9582 = ~n9580 & n9581 ;
  assign n9585 = ~\DataWidth_reg[0]/NET0131  & ~\DataWidth_reg[1]/NET0131  ;
  assign n9586 = ~\rEIP_reg[0]/NET0131  & n9585 ;
  assign n9583 = \ByteEnable_reg[1]/NET0131  & n9566 ;
  assign n9584 = \rEIP_reg[1]/NET0131  & ~n9566 ;
  assign n9587 = ~n9583 & ~n9584 ;
  assign n9588 = ~n9586 & n9587 ;
  assign n9589 = ~READY_n_pad & \State_reg[0]/NET0131  ;
  assign n9590 = NA_n_pad & ~\State_reg[0]/NET0131  ;
  assign n9591 = \State_reg[2]/NET0131  & ~n9590 ;
  assign n9592 = ~n9589 & ~n9591 ;
  assign n9593 = ~HOLD_pad & ~n9592 ;
  assign n9594 = \State_reg[0]/NET0131  & ~\State_reg[1]/NET0131  ;
  assign n9595 = ~\State_reg[2]/NET0131  & n9594 ;
  assign n9596 = ~n9593 & ~n9595 ;
  assign n9597 = \RequestPending_reg/NET0131  & ~n9596 ;
  assign n9598 = ~n8438 & ~n9597 ;
  assign n9603 = ~\rEIP_reg[3]/NET0131  & ~n8449 ;
  assign n9604 = n830 & ~n8450 ;
  assign n9605 = ~n9603 & n9604 ;
  assign n9599 = \Address[1]_pad  & ~n829 ;
  assign n9600 = ~\rEIP_reg[2]/NET0131  & ~n9368 ;
  assign n9601 = n8438 & ~n9369 ;
  assign n9602 = ~n9600 & n9601 ;
  assign n9606 = ~n9599 & ~n9602 ;
  assign n9607 = ~n9605 & n9606 ;
  assign n9612 = ~\rEIP_reg[19]/NET0131  & ~n8539 ;
  assign n9613 = n830 & ~n9435 ;
  assign n9614 = ~n9612 & n9613 ;
  assign n9608 = \Address[17]_pad  & ~n829 ;
  assign n9609 = ~\rEIP_reg[18]/NET0131  & ~n8533 ;
  assign n9610 = n8438 & ~n9500 ;
  assign n9611 = ~n9609 & n9610 ;
  assign n9615 = ~n9608 & ~n9611 ;
  assign n9616 = ~n9614 & n9615 ;
  assign n9621 = ~\rEIP_reg[7]/NET0131  & ~n8453 ;
  assign n9622 = n830 & ~n8454 ;
  assign n9623 = ~n9621 & n9622 ;
  assign n9617 = \Address[5]_pad  & ~n829 ;
  assign n9618 = ~\rEIP_reg[6]/NET0131  & ~n9372 ;
  assign n9619 = n8438 & ~n9108 ;
  assign n9620 = ~n9618 & n9619 ;
  assign n9624 = ~n9617 & ~n9620 ;
  assign n9625 = ~n9623 & n9624 ;
  assign n9626 = \State_reg[0]/NET0131  & \State_reg[1]/NET0131  ;
  assign n9627 = ~\State_reg[2]/NET0131  & n9626 ;
  assign n9628 = ~HOLD_pad & ~\RequestPending_reg/NET0131  ;
  assign n9629 = READY_n_pad & ~n9628 ;
  assign n9630 = n9627 & n9629 ;
  assign n9631 = ~n832 & ~n9630 ;
  assign n9632 = ~NA_n_pad & ~n9631 ;
  assign n9633 = ~\RequestPending_reg/NET0131  & ~\State_reg[1]/NET0131  ;
  assign n9634 = ~\State_reg[2]/NET0131  & ~n9633 ;
  assign n9635 = HOLD_pad & \State_reg[0]/NET0131  ;
  assign n9636 = ~n9634 & n9635 ;
  assign n9637 = \State_reg[1]/NET0131  & \State_reg[2]/NET0131  ;
  assign n9638 = ~n9589 & n9637 ;
  assign n9639 = ~n9636 & ~n9638 ;
  assign n9640 = ~n9632 & n9639 ;
  assign n9641 = \ByteEnable_reg[3]/NET0131  & n9566 ;
  assign n9642 = \rEIP_reg[1]/NET0131  & ~n9586 ;
  assign n9643 = ~\DataWidth_reg[1]/NET0131  & ~n9642 ;
  assign n9644 = ~n9641 & ~n9643 ;
  assign n9649 = ~\rEIP_reg[2]/NET0131  & ~n8448 ;
  assign n9650 = n830 & ~n8449 ;
  assign n9651 = ~n9649 & n9650 ;
  assign n9645 = \Address[0]_pad  & ~n829 ;
  assign n9646 = ~\rEIP_reg[1]/NET0131  & ~n8439 ;
  assign n9647 = n8438 & ~n9368 ;
  assign n9648 = ~n9646 & n9647 ;
  assign n9652 = ~n9645 & ~n9648 ;
  assign n9653 = ~n9651 & n9652 ;
  assign n9654 = ~n831 & ~n9627 ;
  assign n9655 = ~\DataWidth_reg[1]/NET0131  & n9654 ;
  assign n9656 = ~n832 & ~n9627 ;
  assign n9657 = ~\BS16_n_pad  & ~n9656 ;
  assign n9658 = ~n9655 & ~n9657 ;
  assign n9659 = ADS_n_pad & \State_reg[0]/NET0131  ;
  assign n9660 = n9654 & ~n9659 ;
  assign n9661 = \BE_n[2]_pad  & ~n829 ;
  assign n9662 = \ByteEnable_reg[2]/NET0131  & n829 ;
  assign n9663 = ~n9661 & ~n9662 ;
  assign n9664 = \BE_n[0]_pad  & ~n829 ;
  assign n9665 = \ByteEnable_reg[0]/NET0131  & n829 ;
  assign n9666 = ~n9664 & ~n9665 ;
  assign n9667 = \BE_n[1]_pad  & ~n829 ;
  assign n9668 = \ByteEnable_reg[1]/NET0131  & n829 ;
  assign n9669 = ~n9667 & ~n9668 ;
  assign n9670 = \BE_n[3]_pad  & ~n829 ;
  assign n9671 = \ByteEnable_reg[3]/NET0131  & n829 ;
  assign n9672 = ~n9670 & ~n9671 ;
  assign n9673 = W_R_n_pad & ~n829 ;
  assign n9674 = ~\ReadRequest_reg/NET0131  & n829 ;
  assign n9675 = ~n9673 & ~n9674 ;
  assign n9676 = M_IO_n_pad & ~n829 ;
  assign n9677 = \MemoryFetch_reg/NET0131  & n829 ;
  assign n9678 = ~n9676 & ~n9677 ;
  assign n9679 = ~\State_reg[1]/NET0131  & \State_reg[2]/NET0131  ;
  assign n9680 = ~\State_reg[0]/NET0131  & ~n9679 ;
  assign n9681 = ~D_C_n_pad & ~n9680 ;
  assign n9682 = \CodeFetch_reg/NET0131  & n829 ;
  assign n9683 = ~n9681 & ~n9682 ;
  assign n9684 = \DataWidth_reg[0]/NET0131  & n9654 ;
  assign n9685 = ~n9657 & ~n9684 ;
  assign n9686 = \InstAddrPointer_reg[13]/NET0131  & ~n921 ;
  assign n9690 = n1012 & n1422 ;
  assign n9692 = ~\InstAddrPointer_reg[13]/NET0131  & ~n1321 ;
  assign n9693 = ~n1322 & ~n9692 ;
  assign n9694 = ~n9690 & n9693 ;
  assign n9691 = ~\InstAddrPointer_reg[13]/NET0131  & n9690 ;
  assign n9695 = n1051 & ~n9691 ;
  assign n9696 = ~n9694 & n9695 ;
  assign n9687 = n1504 & ~n2165 ;
  assign n9688 = ~n1051 & ~n1766 ;
  assign n9689 = ~n9687 & n9688 ;
  assign n9697 = n921 & ~n9689 ;
  assign n9698 = ~n9696 & n9697 ;
  assign n9699 = ~n9686 & ~n9698 ;
  assign n9700 = n748 & ~n9699 ;
  assign n9702 = n1653 & n2243 ;
  assign n9704 = n1648 & n9702 ;
  assign n9703 = ~n1648 & ~n9702 ;
  assign n9705 = n930 & ~n9703 ;
  assign n9706 = ~n9704 & n9705 ;
  assign n9707 = \InstAddrPointer_reg[13]/NET0131  & ~n1937 ;
  assign n9708 = ~n867 & n9693 ;
  assign n9701 = ~n780 & n1504 ;
  assign n9709 = n809 & n1648 ;
  assign n9710 = ~n9701 & ~n9709 ;
  assign n9711 = ~n9708 & n9710 ;
  assign n9712 = ~n9707 & n9711 ;
  assign n9713 = ~n9706 & n9712 ;
  assign n9714 = ~n9700 & n9713 ;
  assign n9715 = n948 & ~n9714 ;
  assign n9716 = \rEIP_reg[13]/NET0131  & n1731 ;
  assign n9717 = \InstAddrPointer_reg[13]/NET0131  & ~n1736 ;
  assign n9718 = ~n9716 & ~n9717 ;
  assign n9719 = ~n9715 & n9718 ;
  assign n9722 = \InstAddrPointer_reg[16]/NET0131  & ~n921 ;
  assign n9723 = ~n2775 & ~n9722 ;
  assign n9724 = n748 & ~n9723 ;
  assign n9730 = ~n836 & ~n1380 ;
  assign n9731 = n874 & ~n9730 ;
  assign n9732 = n862 & n1373 ;
  assign n9733 = \InstAddrPointer_reg[16]/NET0131  & ~n9732 ;
  assign n9734 = n1379 & n2235 ;
  assign n9735 = ~n9733 & ~n9734 ;
  assign n9736 = ~n9731 & ~n9735 ;
  assign n9729 = ~n780 & n1516 ;
  assign n9721 = n698 & ~n1380 ;
  assign n9725 = ~\InstAddrPointer_reg[16]/NET0131  & ~n808 ;
  assign n9726 = ~n756 & n1872 ;
  assign n9727 = n924 & ~n9726 ;
  assign n9728 = ~n9725 & ~n9727 ;
  assign n9737 = ~n9721 & ~n9728 ;
  assign n9738 = ~n9729 & n9737 ;
  assign n9739 = ~n9736 & n9738 ;
  assign n9740 = ~n2764 & n9739 ;
  assign n9741 = ~n9724 & n9740 ;
  assign n9742 = n948 & ~n9741 ;
  assign n9720 = \InstAddrPointer_reg[16]/NET0131  & ~n1736 ;
  assign n9743 = ~n2784 & ~n9720 ;
  assign n9744 = ~n9742 & n9743 ;
  assign n9747 = \InstAddrPointer_reg[17]/NET0131  & ~n921 ;
  assign n9748 = ~n2819 & ~n9747 ;
  assign n9749 = n748 & ~n9748 ;
  assign n9751 = ~READY_n_pad & ~n1383 ;
  assign n9754 = ~n828 & ~n9751 ;
  assign n9755 = n1891 & ~n9754 ;
  assign n9756 = \InstAddrPointer_reg[17]/NET0131  & ~n9755 ;
  assign n9757 = ~n780 & n1522 ;
  assign n9750 = ~\InstAddrPointer_reg[17]/NET0131  & READY_n_pad ;
  assign n9752 = ~n9750 & ~n9751 ;
  assign n9753 = n2506 & n9752 ;
  assign n9746 = n698 & n1383 ;
  assign n9759 = n808 & ~n1600 ;
  assign n9758 = ~\InstAddrPointer_reg[17]/NET0131  & ~n808 ;
  assign n9760 = ~n756 & ~n9758 ;
  assign n9761 = ~n9759 & n9760 ;
  assign n9762 = ~n9746 & ~n9761 ;
  assign n9763 = ~n9753 & n9762 ;
  assign n9764 = ~n9757 & n9763 ;
  assign n9765 = ~n9756 & n9764 ;
  assign n9766 = ~n2806 & n9765 ;
  assign n9767 = ~n9749 & n9766 ;
  assign n9768 = n948 & ~n9767 ;
  assign n9745 = \InstAddrPointer_reg[17]/NET0131  & ~n1736 ;
  assign n9769 = ~n2799 & ~n9745 ;
  assign n9770 = ~n9768 & n9769 ;
  assign n9773 = \InstAddrPointer_reg[10]/NET0131  & ~n921 ;
  assign n9774 = ~n2981 & ~n9773 ;
  assign n9775 = n748 & ~n9774 ;
  assign n9777 = \InstAddrPointer_reg[10]/NET0131  & n2506 ;
  assign n9778 = n839 & ~n9777 ;
  assign n9779 = n2535 & ~n9778 ;
  assign n9772 = \InstAddrPointer_reg[10]/NET0131  & ~n2508 ;
  assign n9776 = n809 & n1799 ;
  assign n9780 = ~n780 & n1484 ;
  assign n9781 = ~n9776 & ~n9780 ;
  assign n9782 = ~n9772 & n9781 ;
  assign n9783 = ~n9779 & n9782 ;
  assign n9784 = ~n2972 & n9783 ;
  assign n9785 = ~n9775 & n9784 ;
  assign n9786 = n948 & ~n9785 ;
  assign n9771 = \InstAddrPointer_reg[10]/NET0131  & ~n1736 ;
  assign n9787 = ~n2998 & ~n9771 ;
  assign n9788 = ~n9786 & n9787 ;
  assign n9789 = \EBX_reg[29]/NET0131  & n6990 ;
  assign n9790 = ~\EBX_reg[30]/NET0131  & ~n9789 ;
  assign n9791 = \EBX_reg[29]/NET0131  & \EBX_reg[30]/NET0131  ;
  assign n9792 = n6990 & n9791 ;
  assign n9793 = n773 & ~n9792 ;
  assign n9794 = ~n9790 & n9793 ;
  assign n9795 = \EBX_reg[30]/NET0131  & n3486 ;
  assign n9796 = ~n3408 & n3439 ;
  assign n9797 = ~n3440 & ~n9796 ;
  assign n9798 = n3454 & n9797 ;
  assign n9799 = ~n9795 & ~n9798 ;
  assign n9800 = ~n9794 & n9799 ;
  assign n9801 = n948 & ~n9800 ;
  assign n9802 = \EBX_reg[30]/NET0131  & ~n3116 ;
  assign n9803 = ~n9801 & ~n9802 ;
  assign n9805 = \InstAddrPointer_reg[26]/NET0131  & ~n921 ;
  assign n9806 = ~n2698 & ~n9805 ;
  assign n9807 = n748 & ~n9806 ;
  assign n9808 = ~n756 & ~n1686 ;
  assign n9809 = n2073 & ~n9808 ;
  assign n9810 = \InstAddrPointer_reg[26]/NET0131  & ~n9809 ;
  assign n9811 = ~n839 & n1353 ;
  assign n9812 = n809 & n1688 ;
  assign n9813 = ~n780 & ~n1543 ;
  assign n9814 = ~n9812 & ~n9813 ;
  assign n9815 = ~n9811 & n9814 ;
  assign n9816 = ~n9810 & n9815 ;
  assign n9817 = ~n2706 & n9816 ;
  assign n9818 = ~n9807 & n9817 ;
  assign n9819 = n948 & ~n9818 ;
  assign n9804 = \InstAddrPointer_reg[26]/NET0131  & ~n1736 ;
  assign n9820 = ~n2721 & ~n9804 ;
  assign n9821 = ~n9819 & n9820 ;
  assign n9823 = ~\EAX_reg[30]/NET0131  & ~n3147 ;
  assign n9824 = n3118 & ~n3148 ;
  assign n9825 = ~n9823 & n9824 ;
  assign n9826 = \EAX_reg[30]/NET0131  & ~n3447 ;
  assign n9822 = n3153 & n9797 ;
  assign n9827 = \Datai[30]_pad  & n835 ;
  assign n9828 = ~n6972 & ~n9827 ;
  assign n9829 = n826 & ~n9828 ;
  assign n9830 = ~n9822 & ~n9829 ;
  assign n9831 = ~n9826 & n9830 ;
  assign n9832 = ~n9825 & n9831 ;
  assign n9833 = n948 & ~n9832 ;
  assign n9834 = \EAX_reg[30]/NET0131  & ~n3116 ;
  assign n9835 = ~n9833 & ~n9834 ;
  assign n9838 = n3851 & n9791 ;
  assign n9839 = n3483 & n9838 ;
  assign n9841 = \EBX_reg[31]/NET0131  & n9839 ;
  assign n9840 = ~\EBX_reg[31]/NET0131  & ~n9839 ;
  assign n9842 = n773 & ~n9840 ;
  assign n9843 = ~n9841 & n9842 ;
  assign n9836 = \EBX_reg[31]/NET0131  & n3486 ;
  assign n9837 = n3440 & n3454 ;
  assign n9844 = ~n9836 & ~n9837 ;
  assign n9845 = ~n9843 & n9844 ;
  assign n9846 = n948 & ~n9845 ;
  assign n9847 = \EBX_reg[31]/NET0131  & ~n3116 ;
  assign n9848 = ~n9846 & ~n9847 ;
  assign n9850 = n948 & ~n4286 ;
  assign n9851 = n3816 & ~n9850 ;
  assign n9852 = \Datao_reg[22]/NET0131  & ~n9851 ;
  assign n9849 = \uWord_reg[6]/NET0131  & n956 ;
  assign n9853 = n895 & n948 ;
  assign n9854 = n7427 & n9853 ;
  assign n9855 = ~n9849 & ~n9854 ;
  assign n9856 = ~n9852 & n9855 ;
  assign n9859 = \InstAddrPointer_reg[7]/NET0131  & ~n921 ;
  assign n9860 = ~n3026 & ~n9859 ;
  assign n9861 = n748 & ~n9860 ;
  assign n9864 = \InstAddrPointer_reg[7]/NET0131  & ~n1937 ;
  assign n9863 = ~n867 & n1017 ;
  assign n9858 = ~n780 & n1438 ;
  assign n9862 = n809 & n1632 ;
  assign n9865 = ~n9858 & ~n9862 ;
  assign n9866 = ~n9863 & n9865 ;
  assign n9867 = ~n9864 & n9866 ;
  assign n9868 = ~n3014 & n9867 ;
  assign n9869 = ~n9861 & n9868 ;
  assign n9870 = n948 & ~n9869 ;
  assign n9857 = \InstAddrPointer_reg[7]/NET0131  & ~n1736 ;
  assign n9871 = ~n3039 & ~n9857 ;
  assign n9872 = ~n9870 & n9871 ;
  assign n9886 = \PhyAddrPointer_reg[21]/NET0131  & ~n921 ;
  assign n9891 = ~n2298 & ~n2305 ;
  assign n9892 = n2298 & n2305 ;
  assign n9893 = ~n9891 & ~n9892 ;
  assign n9894 = n1051 & ~n9893 ;
  assign n9887 = ~n1533 & ~n2168 ;
  assign n9888 = n1533 & n2168 ;
  assign n9889 = ~n9887 & ~n9888 ;
  assign n9890 = ~n1051 & ~n9889 ;
  assign n9895 = n921 & ~n9890 ;
  assign n9896 = ~n9894 & n9895 ;
  assign n9897 = ~n9886 & ~n9896 ;
  assign n9898 = n748 & ~n9897 ;
  assign n9880 = ~\InstAddrPointer_reg[21]/NET0131  & ~n1670 ;
  assign n9881 = ~n1689 & ~n9880 ;
  assign n9882 = n1668 & n1672 ;
  assign n9883 = ~n9881 & ~n9882 ;
  assign n9884 = n930 & ~n1674 ;
  assign n9885 = ~n9883 & n9884 ;
  assign n9899 = \PhyAddrPointer_reg[21]/NET0131  & ~n1997 ;
  assign n9900 = ~n9885 & ~n9899 ;
  assign n9901 = ~n9898 & n9900 ;
  assign n9902 = n948 & ~n9901 ;
  assign n9879 = n2039 & n5889 ;
  assign n9873 = n971 & ~n2638 ;
  assign n9874 = n2003 & ~n9873 ;
  assign n9875 = \PhyAddrPointer_reg[21]/NET0131  & ~n9874 ;
  assign n9876 = ~\PhyAddrPointer_reg[21]/NET0131  & n971 ;
  assign n9877 = n2638 & n9876 ;
  assign n9878 = \rEIP_reg[21]/NET0131  & n1731 ;
  assign n9903 = ~n9877 & ~n9878 ;
  assign n9904 = ~n9875 & n9903 ;
  assign n9905 = ~n9879 & n9904 ;
  assign n9906 = ~n9902 & n9905 ;
  assign n9908 = \InstAddrPointer_reg[15]/NET0131  & ~n921 ;
  assign n9909 = ~n2353 & ~n9908 ;
  assign n9910 = n748 & ~n9909 ;
  assign n9919 = ~\InstAddrPointer_reg[15]/NET0131  & ~n838 ;
  assign n9920 = ~n744 & ~n9919 ;
  assign n9921 = n666 & n734 ;
  assign n9922 = ~n9920 & ~n9921 ;
  assign n9923 = ~n875 & n1373 ;
  assign n9924 = ~n1372 & ~n9923 ;
  assign n9925 = ~n9922 & n9924 ;
  assign n9913 = ~n780 & n1512 ;
  assign n9911 = \InstAddrPointer_reg[15]/NET0131  & ~n808 ;
  assign n9914 = n808 & n1662 ;
  assign n9915 = ~n9911 & ~n9914 ;
  assign n9916 = ~n756 & ~n9915 ;
  assign n9912 = n746 & n9911 ;
  assign n9917 = n698 & ~n733 ;
  assign n9918 = n1374 & n9917 ;
  assign n9926 = ~n9912 & ~n9918 ;
  assign n9927 = ~n9916 & n9926 ;
  assign n9928 = ~n9913 & n9927 ;
  assign n9929 = ~n9925 & n9928 ;
  assign n9930 = ~n2361 & n9929 ;
  assign n9931 = ~n9910 & n9930 ;
  assign n9932 = n948 & ~n9931 ;
  assign n9907 = \InstAddrPointer_reg[15]/NET0131  & ~n1736 ;
  assign n9933 = ~n2380 & ~n9907 ;
  assign n9934 = ~n9932 & n9933 ;
  assign n9935 = \PhyAddrPointer_reg[13]/NET0131  & ~n921 ;
  assign n9936 = ~n9698 & ~n9935 ;
  assign n9937 = n748 & ~n9936 ;
  assign n9938 = \PhyAddrPointer_reg[13]/NET0131  & ~n1997 ;
  assign n9939 = ~n9706 & ~n9938 ;
  assign n9940 = ~n9937 & n9939 ;
  assign n9941 = n948 & ~n9940 ;
  assign n9947 = n2039 & n6610 ;
  assign n9942 = n971 & ~n2014 ;
  assign n9943 = n2003 & ~n9942 ;
  assign n9944 = \PhyAddrPointer_reg[13]/NET0131  & ~n9943 ;
  assign n9945 = ~\PhyAddrPointer_reg[13]/NET0131  & n971 ;
  assign n9946 = n2014 & n9945 ;
  assign n9948 = ~n9716 & ~n9946 ;
  assign n9949 = ~n9944 & n9948 ;
  assign n9950 = ~n9947 & n9949 ;
  assign n9951 = ~n9941 & n9950 ;
  assign n9952 = \EAX_reg[27]/NET0131  & ~n3116 ;
  assign n9954 = ~n3445 & ~n3568 ;
  assign n9955 = \EAX_reg[27]/NET0131  & ~n9954 ;
  assign n9962 = ~\EAX_reg[27]/NET0131  & n3118 ;
  assign n9963 = n3567 & n9962 ;
  assign n9956 = \EAX_reg[27]/NET0131  & ~n826 ;
  assign n9959 = \Datai[27]_pad  & n826 ;
  assign n9960 = ~n9956 & ~n9959 ;
  assign n9961 = n835 & ~n9960 ;
  assign n9953 = n3153 & n3456 ;
  assign n9957 = ~n4757 & ~n9956 ;
  assign n9958 = n736 & ~n9957 ;
  assign n9964 = ~n9953 & ~n9958 ;
  assign n9965 = ~n9961 & n9964 ;
  assign n9966 = ~n9963 & n9965 ;
  assign n9967 = ~n9955 & n9966 ;
  assign n9968 = n948 & ~n9967 ;
  assign n9969 = ~n9952 & ~n9968 ;
  assign n9970 = \PhyAddrPointer_reg[9]/NET0131  & ~n921 ;
  assign n9971 = ~n2739 & ~n9970 ;
  assign n9972 = n748 & ~n9971 ;
  assign n9973 = \PhyAddrPointer_reg[9]/NET0131  & ~n1997 ;
  assign n9974 = ~n2746 & ~n9973 ;
  assign n9975 = ~n9972 & n9974 ;
  assign n9976 = n948 & ~n9975 ;
  assign n9980 = n2039 & n6460 ;
  assign n9977 = ~\PhyAddrPointer_reg[9]/NET0131  & ~n2010 ;
  assign n9978 = n971 & ~n2011 ;
  assign n9979 = ~n9977 & n9978 ;
  assign n9981 = \PhyAddrPointer_reg[9]/NET0131  & ~n2003 ;
  assign n9982 = ~n2726 & ~n9981 ;
  assign n9983 = ~n9979 & n9982 ;
  assign n9984 = ~n9980 & n9983 ;
  assign n9985 = ~n9976 & n9984 ;
  assign n9986 = \PhyAddrPointer_reg[12]/NET0131  & ~n921 ;
  assign n9987 = ~n2543 & ~n9986 ;
  assign n9988 = n748 & ~n9987 ;
  assign n9989 = \PhyAddrPointer_reg[12]/NET0131  & ~n1997 ;
  assign n9990 = ~n2550 & ~n9989 ;
  assign n9991 = ~n9988 & n9990 ;
  assign n9992 = n948 & ~n9991 ;
  assign n9994 = ~\DataWidth_reg[1]/NET0131  & ~n6573 ;
  assign n9995 = ~\PhyAddrPointer_reg[12]/NET0131  & ~n2013 ;
  assign n9996 = ~n2014 & ~n9995 ;
  assign n9997 = \DataWidth_reg[1]/NET0131  & ~n9996 ;
  assign n9998 = n952 & ~n9997 ;
  assign n9999 = ~n9994 & n9998 ;
  assign n9993 = n970 & n6573 ;
  assign n10000 = \PhyAddrPointer_reg[12]/NET0131  & ~n2003 ;
  assign n10001 = ~n2565 & ~n10000 ;
  assign n10002 = ~n9993 & n10001 ;
  assign n10003 = ~n9999 & n10002 ;
  assign n10004 = ~n9992 & n10003 ;
  assign n10006 = \InstAddrPointer_reg[18]/NET0131  & ~n921 ;
  assign n10007 = ~n2839 & ~n10006 ;
  assign n10008 = n748 & ~n10007 ;
  assign n10009 = \InstAddrPointer_reg[18]/NET0131  & ~n2908 ;
  assign n10011 = ~n867 & n1387 ;
  assign n10010 = ~n780 & n1520 ;
  assign n10012 = n809 & n1810 ;
  assign n10013 = ~n10010 & ~n10012 ;
  assign n10014 = ~n10011 & n10013 ;
  assign n10015 = ~n10009 & n10014 ;
  assign n10016 = ~n2846 & n10015 ;
  assign n10017 = ~n10008 & n10016 ;
  assign n10018 = n948 & ~n10017 ;
  assign n10005 = \InstAddrPointer_reg[18]/NET0131  & ~n1736 ;
  assign n10019 = ~n2850 & ~n10005 ;
  assign n10020 = ~n10018 & n10019 ;
  assign n10022 = \InstAddrPointer_reg[21]/NET0131  & ~n921 ;
  assign n10023 = ~n9896 & ~n10022 ;
  assign n10024 = n748 & ~n10023 ;
  assign n10025 = ~n756 & ~n1670 ;
  assign n10026 = n2908 & ~n10025 ;
  assign n10027 = \InstAddrPointer_reg[21]/NET0131  & ~n10026 ;
  assign n10029 = ~n780 & n1533 ;
  assign n10021 = ~n867 & n2298 ;
  assign n10028 = n809 & n9881 ;
  assign n10030 = ~n10021 & ~n10028 ;
  assign n10031 = ~n10029 & n10030 ;
  assign n10032 = ~n10027 & n10031 ;
  assign n10033 = ~n9885 & n10032 ;
  assign n10034 = ~n10024 & n10033 ;
  assign n10035 = n948 & ~n10034 ;
  assign n10036 = \InstAddrPointer_reg[21]/NET0131  & ~n1736 ;
  assign n10037 = ~n9878 & ~n10036 ;
  assign n10038 = ~n10035 & n10037 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g47521/_2_  = ~n966 ;
  assign \g47523/_0_  = ~n975 ;
  assign \g47526/_0_  = ~n992 ;
  assign \g47529/_0_  = ~n994 ;
  assign \g47533/_0_  = ~n1739 ;
  assign \g47540/_0_  = ~n1834 ;
  assign \g47551/_0_  = ~n1907 ;
  assign \g47552/_0_  = ~n1952 ;
  assign \g47553/_0_  = ~n1993 ;
  assign \g47563/_2_  = ~n2048 ;
  assign \g47566/_0_  = ~n2085 ;
  assign \g47567/_0_  = ~n2118 ;
  assign \g47568/_0_  = ~n2155 ;
  assign \g47569/_0_  = ~n2198 ;
  assign \g47583/_2_  = ~n2217 ;
  assign \g47584/_0_  = ~n2262 ;
  assign \g47585/_0_  = ~n2294 ;
  assign \g47589/_0_  = ~n2344 ;
  assign \g47602/_0_  = ~n2385 ;
  assign \g47603/_0_  = ~n2407 ;
  assign \g47604/_2_  = ~n2428 ;
  assign \g47605/_0_  = ~n2447 ;
  assign \g47606/_2_  = ~n2490 ;
  assign \g47609/_0_  = ~n2522 ;
  assign \g47611/_0_  = ~n2568 ;
  assign \g47631/_0_  = ~n2587 ;
  assign \g47632/_0_  = ~n2605 ;
  assign \g47633/_0_  = ~n2628 ;
  assign \g47635/_0_  = ~n2651 ;
  assign \g47636/_0_  = ~n2671 ;
  assign \g47637/_0_  = ~n2688 ;
  assign \g47638/_2_  = ~n2725 ;
  assign \g47643/_0_  = ~n2756 ;
  assign \g47665/_2_  = ~n2792 ;
  assign \g47666/_0_  = ~n2829 ;
  assign \g47667/_0_  = ~n2860 ;
  assign \g47670/_0_  = ~n2877 ;
  assign \g47672/_0_  = ~n2900 ;
  assign \g47677/_0_  = ~n2933 ;
  assign \g47678/_0_  = ~n2969 ;
  assign \g47706/_0_  = ~n3003 ;
  assign \g47711/_0_  = ~n3044 ;
  assign \g47717/_0_  = ~n3086 ;
  assign \g47718/_0_  = ~n3113 ;
  assign \g47721/_0_  = ~n3453 ;
  assign \g47722/_0_  = ~n3495 ;
  assign \g47751/_0_  = ~n3515 ;
  assign \g47755/_0_  = ~n3547 ;
  assign \g47756/_0_  = ~n3561 ;
  assign \g47757/_0_  = ~n3580 ;
  assign \g47759/_0_  = ~n3625 ;
  assign \g47789/_0_  = ~n3638 ;
  assign \g47793/_0_  = ~n3653 ;
  assign \g47797/_0_  = ~n3676 ;
  assign \g47798/_0_  = ~n3697 ;
  assign \g47799/_0_  = ~n3717 ;
  assign \g47802/_0_  = ~n3746 ;
  assign \g47804/_0_  = ~n3756 ;
  assign \g47807/_0_  = ~n3778 ;
  assign \g47809/_0_  = ~n3796 ;
  assign \g47862/_0_  = ~n3819 ;
  assign \g47863/_0_  = ~n3830 ;
  assign \g47864/_0_  = ~n3839 ;
  assign \g47869/_0_  = ~n3848 ;
  assign \g47870/_0_  = ~n3861 ;
  assign \g47924/_0_  = ~n3937 ;
  assign \g47925/_0_  = ~n3965 ;
  assign \g47926/_0_  = ~n3989 ;
  assign \g47927/_0_  = ~n4012 ;
  assign \g47928/_0_  = ~n4033 ;
  assign \g47930/_0_  = ~n4053 ;
  assign \g47932/_0_  = ~n4074 ;
  assign \g47933/_0_  = ~n4096 ;
  assign \g47934/_0_  = ~n4118 ;
  assign \g47935/_0_  = ~n4140 ;
  assign \g47936/_0_  = ~n4162 ;
  assign \g47937/_0_  = ~n4184 ;
  assign \g47938/_0_  = ~n4206 ;
  assign \g47939/_0_  = ~n4227 ;
  assign \g47940/_0_  = ~n4247 ;
  assign \g47941/_0_  = ~n4267 ;
  assign \g47957/_0_  = ~n4279 ;
  assign \g47970/_0_  = ~n4292 ;
  assign \g47973/_0_  = ~n4298 ;
  assign \g47975/_0_  = ~n4318 ;
  assign \g48058/_0_  = ~n4345 ;
  assign \g48059/_0_  = ~n4364 ;
  assign \g48060/_0_  = ~n4383 ;
  assign \g48061/_0_  = ~n4402 ;
  assign \g48062/_0_  = ~n4421 ;
  assign \g48064/_0_  = ~n4440 ;
  assign \g48065/_0_  = ~n4459 ;
  assign \g48066/_0_  = ~n4478 ;
  assign \g48067/_0_  = ~n4497 ;
  assign \g48068/_0_  = ~n4516 ;
  assign \g48069/_0_  = ~n4535 ;
  assign \g48070/_0_  = ~n4554 ;
  assign \g48071/_0_  = ~n4573 ;
  assign \g48072/_0_  = ~n4592 ;
  assign \g48073/_0_  = ~n4611 ;
  assign \g48074/_0_  = ~n4630 ;
  assign \g48087/_0_  = ~n4730 ;
  assign \g48110/_0_  = ~n4741 ;
  assign \g48117/_0_  = ~n4754 ;
  assign \g48118/_0_  = ~n4762 ;
  assign \g48119/_0_  = ~n4773 ;
  assign \g48120/_0_  = ~n4783 ;
  assign \g48121/_0_  = ~n4793 ;
  assign \g48122/_0_  = ~n4803 ;
  assign \g48124/_0_  = ~n4813 ;
  assign \g48125/_0_  = ~n4854 ;
  assign \g48126/_0_  = ~n4895 ;
  assign \g48127/_0_  = ~n4936 ;
  assign \g48128/_0_  = ~n4947 ;
  assign \g48129/_0_  = ~n4988 ;
  assign \g48130/_0_  = ~n5031 ;
  assign \g48131/_0_  = ~n5076 ;
  assign \g48132/_0_  = ~n5120 ;
  assign \g48133/_0_  = ~n5164 ;
  assign \g48134/_0_  = ~n5175 ;
  assign \g48168/_0_  = ~n5198 ;
  assign \g48169/_0_  = ~n5221 ;
  assign \g48170/_0_  = ~n5240 ;
  assign \g48171/_0_  = ~n5259 ;
  assign \g48172/_0_  = ~n5278 ;
  assign \g48173/_0_  = ~n5297 ;
  assign \g48174/_0_  = ~n5316 ;
  assign \g48175/_0_  = ~n5335 ;
  assign \g48177/_0_  = ~n5354 ;
  assign \g48178/_0_  = ~n5373 ;
  assign \g48179/_0_  = ~n5392 ;
  assign \g48180/_0_  = ~n5411 ;
  assign \g48181/_0_  = ~n5430 ;
  assign \g48182/_0_  = ~n5449 ;
  assign \g48183/_0_  = ~n5468 ;
  assign \g48184/_0_  = ~n5487 ;
  assign \g48185/_0_  = ~n5506 ;
  assign \g48186/_0_  = ~n5525 ;
  assign \g48187/_0_  = ~n5544 ;
  assign \g48188/_0_  = ~n5563 ;
  assign \g48189/_0_  = ~n5582 ;
  assign \g48192/_0_  = ~n5601 ;
  assign \g48193/_0_  = ~n5620 ;
  assign \g48194/_0_  = ~n5639 ;
  assign \g48195/_0_  = ~n5658 ;
  assign \g48196/_0_  = ~n5677 ;
  assign \g48197/_0_  = ~n5696 ;
  assign \g48198/_0_  = ~n5715 ;
  assign \g48199/_0_  = ~n5734 ;
  assign \g48200/_0_  = ~n5753 ;
  assign \g48201/_0_  = ~n5772 ;
  assign \g48202/_0_  = ~n5791 ;
  assign \g48203/_0_  = ~n5800 ;
  assign \g48213/_0_  = ~n5832 ;
  assign \g48214/_0_  = ~n5867 ;
  assign \g48215/_0_  = ~n5906 ;
  assign \g48216/_0_  = ~n5939 ;
  assign \g48217/_0_  = ~n5971 ;
  assign \g48218/_0_  = ~n6011 ;
  assign \g48219/_0_  = ~n6046 ;
  assign \g48220/_0_  = ~n6078 ;
  assign \g48221/_0_  = ~n6110 ;
  assign \g48222/_0_  = ~n6144 ;
  assign \g48223/_0_  = ~n6183 ;
  assign \g48224/_0_  = ~n6218 ;
  assign \g48225/_0_  = ~n6256 ;
  assign \g48226/_0_  = ~n6291 ;
  assign \g48227/_0_  = ~n6324 ;
  assign \g48228/_0_  = ~n6356 ;
  assign \g48229/_0_  = ~n6390 ;
  assign \g48230/_0_  = ~n6423 ;
  assign \g48231/_0_  = ~n6457 ;
  assign \g48232/_0_  = ~n6492 ;
  assign \g48234/_0_  = ~n6501 ;
  assign \g48236/_0_  = ~n6535 ;
  assign \g48237/_0_  = ~n6570 ;
  assign \g48238/_0_  = ~n6607 ;
  assign \g48239/_0_  = ~n6643 ;
  assign \g48240/_0_  = ~n6677 ;
  assign \g48241/_0_  = ~n6711 ;
  assign \g48243/_0_  = ~n6744 ;
  assign \g48244/_0_  = ~n6782 ;
  assign \g48245/_0_  = ~n6815 ;
  assign \g48246/_0_  = ~n6848 ;
  assign \g48263/_0_  = ~n6860 ;
  assign \g48270/_0_  = ~n6874 ;
  assign \g48273/_0_  = ~n6888 ;
  assign \g48276/_0_  = ~n6897 ;
  assign \g48277/_0_  = ~n6903 ;
  assign \g48370/_0_  = ~n6910 ;
  assign \g48377/_0_  = ~n6916 ;
  assign \g48391/_0_  = ~n6938 ;
  assign \g48423/_0_  = ~n6954 ;
  assign \g48428/_0_  = ~n6970 ;
  assign \g48429/_0_  = ~n6979 ;
  assign \g48431/_0_  = ~n6987 ;
  assign \g48433/_0_  = ~n6999 ;
  assign \g48434/_0_  = ~n7045 ;
  assign \g48435/_0_  = ~n7091 ;
  assign \g48436/_0_  = ~n7140 ;
  assign \g48437/_0_  = ~n7186 ;
  assign \g48438/_0_  = ~n7189 ;
  assign \g48439/_0_  = ~n7235 ;
  assign \g48440/_0_  = ~n7282 ;
  assign \g48441/_0_  = ~n7328 ;
  assign \g48442/_0_  = ~n7344 ;
  assign \g48443/_0_  = ~n7360 ;
  assign \g48610/_0_  = ~n7371 ;
  assign \g48634/_0_  = ~n7379 ;
  assign \g48635/_0_  = ~n7384 ;
  assign \g48636/_0_  = ~n7393 ;
  assign \g48637/_0_  = ~n7405 ;
  assign \g48638/_0_  = ~n7413 ;
  assign \g48639/_0_  = ~n7422 ;
  assign \g48640/_0_  = ~n7430 ;
  assign \g48642/_0_  = ~n7438 ;
  assign \g48643/_0_  = ~n7446 ;
  assign \g48644/_0_  = ~n7456 ;
  assign \g48645/_0_  = ~n7466 ;
  assign \g48646/_0_  = ~n7476 ;
  assign \g48647/_0_  = ~n7487 ;
  assign \g48648/_0_  = ~n7496 ;
  assign \g48649/_0_  = ~n7506 ;
  assign \g48650/_0_  = ~n7516 ;
  assign \g48651/_0_  = ~n7526 ;
  assign \g48652/_0_  = ~n7536 ;
  assign \g48653/_0_  = ~n7546 ;
  assign \g48654/_0_  = ~n7554 ;
  assign \g48655/_0_  = ~n7564 ;
  assign \g48656/_0_  = ~n7575 ;
  assign \g48657/_0_  = ~n7585 ;
  assign \g48658/_0_  = ~n7595 ;
  assign \g48659/_0_  = ~n7605 ;
  assign \g48660/_0_  = ~n7615 ;
  assign \g48662/_0_  = ~n7625 ;
  assign \g48663/_0_  = ~n7635 ;
  assign \g48664/_0_  = ~n7645 ;
  assign \g48665/_0_  = ~n7655 ;
  assign \g48666/_0_  = ~n7665 ;
  assign \g48667/_0_  = ~n7675 ;
  assign \g48668/_0_  = ~n7685 ;
  assign \g48669/_0_  = ~n7688 ;
  assign \g48750/_0_  = ~n7711 ;
  assign \g48753/_0_  = ~n7730 ;
  assign \g48756/_0_  = ~n7749 ;
  assign \g48759/_0_  = ~n7768 ;
  assign \g48763/_0_  = ~n7787 ;
  assign \g48766/_0_  = ~n7806 ;
  assign \g48769/_0_  = ~n7825 ;
  assign \g48772/_0_  = ~n7844 ;
  assign \g48775/_0_  = ~n7863 ;
  assign \g48778/_0_  = ~n7882 ;
  assign \g48781/_0_  = ~n7901 ;
  assign \g48785/_0_  = ~n7920 ;
  assign \g48789/_0_  = ~n7939 ;
  assign \g48792/_0_  = ~n7958 ;
  assign \g48796/_0_  = ~n7977 ;
  assign \g48799/_0_  = ~n7996 ;
  assign \g48937/_0_  = ~n8004 ;
  assign \g48958/_0_  = ~n8010 ;
  assign \g48959/_0_  = ~n8018 ;
  assign \g48964/_0_  = ~n8023 ;
  assign \g48965/_0_  = ~n8028 ;
  assign \g48966/_0_  = ~n8033 ;
  assign \g48967/_0_  = ~n8039 ;
  assign \g48968/_0_  = ~n8044 ;
  assign \g48969/_0_  = ~n8050 ;
  assign \g48970/_0_  = ~n8061 ;
  assign \g48971/_0_  = ~n8067 ;
  assign \g48972/_0_  = ~n8072 ;
  assign \g48973/_0_  = ~n8078 ;
  assign \g48974/_0_  = ~n8083 ;
  assign \g48975/_0_  = ~n8089 ;
  assign \g48976/_0_  = ~n8095 ;
  assign \g48977/_0_  = ~n8101 ;
  assign \g48978/_0_  = ~n8107 ;
  assign \g48979/_0_  = ~n8112 ;
  assign \g49/_0_  = ~n8128 ;
  assign \g49069/_0_  = ~n8151 ;
  assign \g49070/_0_  = ~n8170 ;
  assign \g49071/_0_  = ~n8189 ;
  assign \g49073/_0_  = ~n8208 ;
  assign \g49074/_0_  = ~n8227 ;
  assign \g49076/_0_  = ~n8246 ;
  assign \g49078/_0_  = ~n8265 ;
  assign \g49081/_0_  = ~n8284 ;
  assign \g49083/_0_  = ~n8303 ;
  assign \g49085/_0_  = ~n8322 ;
  assign \g49087/_0_  = ~n8341 ;
  assign \g49088/_0_  = ~n8360 ;
  assign \g49090/_0_  = ~n8379 ;
  assign \g49092/_0_  = ~n8398 ;
  assign \g49095/_0_  = ~n8417 ;
  assign \g49098/_0_  = ~n8436 ;
  assign \g49125/_0_  = ~n8474 ;
  assign \g49162/_0_  = ~n8482 ;
  assign \g49202/_0_  = ~n8493 ;
  assign \g49203/_0_  = ~n8504 ;
  assign \g49206/_0_  = ~n8512 ;
  assign \g49340/_0_  = ~n8528 ;
  assign \g49457/_0_  = ~n8543 ;
  assign \g49512/_0_  = ~n8551 ;
  assign \g49513/_0_  = ~n8559 ;
  assign \g49514/_0_  = ~n8567 ;
  assign \g49515/_0_  = ~n8575 ;
  assign \g49516/_0_  = ~n8583 ;
  assign \g49517/_0_  = ~n8591 ;
  assign \g49518/_0_  = ~n8599 ;
  assign \g49519/_0_  = ~n8607 ;
  assign \g49520/_0_  = ~n8615 ;
  assign \g49521/_0_  = ~n8623 ;
  assign \g49522/_0_  = ~n8631 ;
  assign \g49523/_0_  = ~n8639 ;
  assign \g49524/_0_  = ~n8647 ;
  assign \g49525/_0_  = ~n8655 ;
  assign \g49526/_0_  = ~n8663 ;
  assign \g49527/_0_  = ~n8671 ;
  assign \g49534/_0_  = ~n8686 ;
  assign \g49551/_0_  = ~n8696 ;
  assign \g49573/_0_  = ~n8702 ;
  assign \g49574/_0_  = ~n8725 ;
  assign \g49578/_0_  = ~n8744 ;
  assign \g49582/_0_  = ~n8767 ;
  assign \g49584/_0_  = ~n8786 ;
  assign \g49592/_0_  = ~n8805 ;
  assign \g49600/_0_  = ~n8824 ;
  assign \g49604/_0_  = ~n8843 ;
  assign \g49608/_0_  = ~n8862 ;
  assign \g49612/_0_  = ~n8881 ;
  assign \g49616/_0_  = ~n8900 ;
  assign \g49619/_0_  = ~n8919 ;
  assign \g49620/_0_  = ~n8938 ;
  assign \g49623/_0_  = ~n8957 ;
  assign \g49627/_0_  = ~n8976 ;
  assign \g49630/_0_  = ~n8995 ;
  assign \g49634/_0_  = ~n9014 ;
  assign \g49635/_0_  = ~n9033 ;
  assign \g49639/_0_  = ~n9052 ;
  assign \g49645/_0_  = ~n9071 ;
  assign \g49744/_0_  = ~n9082 ;
  assign \g49766/_0_  = ~n9093 ;
  assign \g50098/_0_  = ~n9106 ;
  assign \g50124/_0_  = ~n9119 ;
  assign \g50195/_0_  = ~n9138 ;
  assign \g50198/_0_  = ~n9157 ;
  assign \g50201/_0_  = ~n9176 ;
  assign \g50203/_0_  = ~n9195 ;
  assign \g50205/_0_  = ~n9214 ;
  assign \g50207/_0_  = ~n9233 ;
  assign \g50209/_0_  = ~n9252 ;
  assign \g50213/_0_  = ~n9271 ;
  assign \g50222/_0_  = ~n9290 ;
  assign \g50228/_0_  = ~n9309 ;
  assign \g50231/_0_  = ~n9328 ;
  assign \g50237/_0_  = ~n9347 ;
  assign \g50240/_0_  = ~n9366 ;
  assign \g50335/_0_  = ~n9380 ;
  assign \g50477/_0_  = ~n9391 ;
  assign \g50478/_0_  = n9401 ;
  assign \g50671/_0_  = ~n9411 ;
  assign \g50757/_0_  = ~n9421 ;
  assign \g50938/_0_  = ~n9430 ;
  assign \g50998/_0_  = ~n9441 ;
  assign \g51008/_0_  = ~n9450 ;
  assign \g51579/_0_  = ~n9459 ;
  assign \g51637/_0_  = ~n9469 ;
  assign \g51662/_0_  = ~n9479 ;
  assign \g52424/_0_  = ~n9489 ;
  assign \g53184/_0_  = ~n9498 ;
  assign \g53206/_0_  = ~n9508 ;
  assign \g53270/_0_  = ~n9517 ;
  assign \g53730/_0_  = ~n9526 ;
  assign \g53754/_0_  = ~n9537 ;
  assign \g54176/_0_  = ~n9546 ;
  assign \g54214/_0_  = ~n9556 ;
  assign \g54229/_0_  = ~n9565 ;
  assign \g54392/_0_  = ~n9573 ;
  assign \g54400/_0_  = ~n9582 ;
  assign \g54415/_0_  = ~n9588 ;
  assign \g54421/_0_  = n9598 ;
  assign \g54604/_0_  = ~n9607 ;
  assign \g54607/_0_  = ~n9616 ;
  assign \g54638/_0_  = ~n9625 ;
  assign \g54694/_0_  = ~n9640 ;
  assign \g54759/_0_  = ~n9644 ;
  assign \g55607/_0_  = ~n9653 ;
  assign \g55863/_1_  = ~n9566 ;
  assign \g56073/_0_  = n9658 ;
  assign \g56292/_0_  = ~n9660 ;
  assign \g56320/_0_  = ~n9663 ;
  assign \g56527/_0_  = ~n9666 ;
  assign \g56531/_0_  = ~n9669 ;
  assign \g56533/_0_  = ~n9672 ;
  assign \g56562/_0_  = ~n9675 ;
  assign \g56615/_0_  = ~n9678 ;
  assign \g56720/_0_  = n9683 ;
  assign \g57044/_0_  = ~n9685 ;
  assign \g60635/_1_  = ~n8447 ;
  assign \g62873/_0_  = ~n9719 ;
  assign \g62886/_0_  = ~n9744 ;
  assign \g63001/_0_  = ~n9770 ;
  assign \g63101/_0_  = ~n9788 ;
  assign \g63129/_0_  = ~n9803 ;
  assign \g63198/_0_  = ~n9821 ;
  assign \g63449/_0_  = ~n9835 ;
  assign \g63471/_0_  = ~n9848 ;
  assign \g63493/_0_  = ~n9856 ;
  assign \g63626/_0_  = ~n9872 ;
  assign \g63688/_0_  = ~n9906 ;
  assign \g63800/_0_  = ~n9934 ;
  assign \g63934/_0_  = ~n9951 ;
  assign \g63954/_0_  = ~n9969 ;
  assign \g64060/_0_  = ~n9985 ;
  assign \g64375/_0_  = ~n10004 ;
  assign \g65/_0_  = ~n10020 ;
  assign \g67/_0_  = ~n10038 ;
endmodule
