module top( \data_i[0]_pad  , \data_i[10]_pad  , \data_i[11]_pad  , \data_i[12]_pad  , \data_i[13]_pad  , \data_i[14]_pad  , \data_i[15]_pad  , \data_i[16]_pad  , \data_i[17]_pad  , \data_i[18]_pad  , \data_i[19]_pad  , \data_i[1]_pad  , \data_i[20]_pad  , \data_i[21]_pad  , \data_i[22]_pad  , \data_i[23]_pad  , \data_i[24]_pad  , \data_i[25]_pad  , \data_i[26]_pad  , \data_i[27]_pad  , \data_i[28]_pad  , \data_i[29]_pad  , \data_i[2]_pad  , \data_i[30]_pad  , \data_i[31]_pad  , \data_i[32]_pad  , \data_i[33]_pad  , \data_i[34]_pad  , \data_i[35]_pad  , \data_i[36]_pad  , \data_i[37]_pad  , \data_i[38]_pad  , \data_i[39]_pad  , \data_i[3]_pad  , \data_i[40]_pad  , \data_i[41]_pad  , \data_i[42]_pad  , \data_i[43]_pad  , \data_i[44]_pad  , \data_i[45]_pad  , \data_i[46]_pad  , \data_i[47]_pad  , \data_i[48]_pad  , \data_i[49]_pad  , \data_i[4]_pad  , \data_i[50]_pad  , \data_i[51]_pad  , \data_i[52]_pad  , \data_i[53]_pad  , \data_i[54]_pad  , \data_i[55]_pad  , \data_i[56]_pad  , \data_i[57]_pad  , \data_i[58]_pad  , \data_i[59]_pad  , \data_i[5]_pad  , \data_i[60]_pad  , \data_i[61]_pad  , \data_i[62]_pad  , \data_i[63]_pad  , \data_i[6]_pad  , \data_i[7]_pad  , \data_i[8]_pad  , \data_i[9]_pad  , \data_ready_reg/NET0131  , decrypt_i_pad , \key_i[10]_pad  , \key_i[11]_pad  , \key_i[12]_pad  , \key_i[13]_pad  , \key_i[14]_pad  , \key_i[15]_pad  , \key_i[17]_pad  , \key_i[18]_pad  , \key_i[19]_pad  , \key_i[1]_pad  , \key_i[20]_pad  , \key_i[21]_pad  , \key_i[22]_pad  , \key_i[23]_pad  , \key_i[25]_pad  , \key_i[26]_pad  , \key_i[27]_pad  , \key_i[28]_pad  , \key_i[29]_pad  , \key_i[2]_pad  , \key_i[30]_pad  , \key_i[31]_pad  , \key_i[33]_pad  , \key_i[34]_pad  , \key_i[35]_pad  , \key_i[36]_pad  , \key_i[37]_pad  , \key_i[38]_pad  , \key_i[39]_pad  , \key_i[3]_pad  , \key_i[41]_pad  , \key_i[42]_pad  , \key_i[43]_pad  , \key_i[44]_pad  , \key_i[45]_pad  , \key_i[46]_pad  , \key_i[47]_pad  , \key_i[49]_pad  , \key_i[4]_pad  , \key_i[50]_pad  , \key_i[51]_pad  , \key_i[52]_pad  , \key_i[53]_pad  , \key_i[54]_pad  , \key_i[55]_pad  , \key_i[57]_pad  , \key_i[58]_pad  , \key_i[59]_pad  , \key_i[5]_pad  , \key_i[60]_pad  , \key_i[61]_pad  , \key_i[62]_pad  , \key_i[63]_pad  , \key_i[6]_pad  , \key_i[7]_pad  , \key_i[9]_pad  , load_i_pad , \rd1_Key_o_reg[0]/NET0131  , \rd1_Key_o_reg[10]/NET0131  , \rd1_Key_o_reg[11]/NET0131  , \rd1_Key_o_reg[12]/NET0131  , \rd1_Key_o_reg[13]/NET0131  , \rd1_Key_o_reg[14]/NET0131  , \rd1_Key_o_reg[15]/NET0131  , \rd1_Key_o_reg[16]/NET0131  , \rd1_Key_o_reg[17]/NET0131  , \rd1_Key_o_reg[18]/NET0131  , \rd1_Key_o_reg[19]/NET0131  , \rd1_Key_o_reg[1]/NET0131  , \rd1_Key_o_reg[20]/NET0131  , \rd1_Key_o_reg[21]/NET0131  , \rd1_Key_o_reg[22]/NET0131  , \rd1_Key_o_reg[23]/NET0131  , \rd1_Key_o_reg[24]/NET0131  , \rd1_Key_o_reg[25]/NET0131  , \rd1_Key_o_reg[26]/NET0131  , \rd1_Key_o_reg[27]/NET0131  , \rd1_Key_o_reg[28]/NET0131  , \rd1_Key_o_reg[29]/NET0131  , \rd1_Key_o_reg[2]/NET0131  , \rd1_Key_o_reg[30]/NET0131  , \rd1_Key_o_reg[31]/NET0131  , \rd1_Key_o_reg[32]/NET0131  , \rd1_Key_o_reg[33]/NET0131  , \rd1_Key_o_reg[34]/NET0131  , \rd1_Key_o_reg[35]/NET0131  , \rd1_Key_o_reg[36]/NET0131  , \rd1_Key_o_reg[37]/NET0131  , \rd1_Key_o_reg[38]/NET0131  , \rd1_Key_o_reg[39]/NET0131  , \rd1_Key_o_reg[3]/NET0131  , \rd1_Key_o_reg[40]/NET0131  , \rd1_Key_o_reg[41]/NET0131  , \rd1_Key_o_reg[42]/NET0131  , \rd1_Key_o_reg[43]/NET0131  , \rd1_Key_o_reg[44]/NET0131  , \rd1_Key_o_reg[45]/NET0131  , \rd1_Key_o_reg[46]/NET0131  , \rd1_Key_o_reg[47]/NET0131  , \rd1_Key_o_reg[48]/NET0131  , \rd1_Key_o_reg[49]/NET0131  , \rd1_Key_o_reg[4]/NET0131  , \rd1_Key_o_reg[50]/NET0131  , \rd1_Key_o_reg[51]/NET0131  , \rd1_Key_o_reg[52]/NET0131  , \rd1_Key_o_reg[53]/NET0131  , \rd1_Key_o_reg[54]/NET0131  , \rd1_Key_o_reg[55]/NET0131  , \rd1_Key_o_reg[5]/NET0131  , \rd1_Key_o_reg[6]/NET0131  , \rd1_Key_o_reg[7]/NET0131  , \rd1_Key_o_reg[8]/NET0131  , \rd1_Key_o_reg[9]/NET0131  , \rd1_L_o_reg[0]/NET0131  , \rd1_L_o_reg[10]/NET0131  , \rd1_L_o_reg[11]/NET0131  , \rd1_L_o_reg[12]/NET0131  , \rd1_L_o_reg[13]/NET0131  , \rd1_L_o_reg[14]/NET0131  , \rd1_L_o_reg[15]/NET0131  , \rd1_L_o_reg[16]/NET0131  , \rd1_L_o_reg[17]/NET0131  , \rd1_L_o_reg[18]/NET0131  , \rd1_L_o_reg[19]/NET0131  , \rd1_L_o_reg[1]/NET0131  , \rd1_L_o_reg[20]/NET0131  , \rd1_L_o_reg[21]/NET0131  , \rd1_L_o_reg[22]/NET0131  , \rd1_L_o_reg[23]/NET0131  , \rd1_L_o_reg[24]/NET0131  , \rd1_L_o_reg[25]/NET0131  , \rd1_L_o_reg[26]/NET0131  , \rd1_L_o_reg[27]/NET0131  , \rd1_L_o_reg[28]/NET0131  , \rd1_L_o_reg[29]/NET0131  , \rd1_L_o_reg[2]/NET0131  , \rd1_L_o_reg[30]/NET0131  , \rd1_L_o_reg[31]/NET0131  , \rd1_L_o_reg[3]/NET0131  , \rd1_L_o_reg[4]/NET0131  , \rd1_L_o_reg[5]/NET0131  , \rd1_L_o_reg[6]/NET0131  , \rd1_L_o_reg[7]/NET0131  , \rd1_L_o_reg[8]/NET0131  , \rd1_L_o_reg[9]/NET0131  , \rd1_R_o_reg[0]/NET0131  , \rd1_R_o_reg[10]/NET0131  , \rd1_R_o_reg[11]/NET0131  , \rd1_R_o_reg[12]/NET0131  , \rd1_R_o_reg[13]/NET0131  , \rd1_R_o_reg[14]/NET0131  , \rd1_R_o_reg[15]/NET0131  , \rd1_R_o_reg[16]/NET0131  , \rd1_R_o_reg[17]/NET0131  , \rd1_R_o_reg[18]/NET0131  , \rd1_R_o_reg[19]/NET0131  , \rd1_R_o_reg[1]/NET0131  , \rd1_R_o_reg[20]/NET0131  , \rd1_R_o_reg[21]/NET0131  , \rd1_R_o_reg[22]/NET0131  , \rd1_R_o_reg[23]/NET0131  , \rd1_R_o_reg[24]/NET0131  , \rd1_R_o_reg[25]/NET0131  , \rd1_R_o_reg[26]/NET0131  , \rd1_R_o_reg[27]/NET0131  , \rd1_R_o_reg[28]/NET0131  , \rd1_R_o_reg[29]/NET0131  , \rd1_R_o_reg[2]/NET0131  , \rd1_R_o_reg[30]/NET0131  , \rd1_R_o_reg[31]/NET0131  , \rd1_R_o_reg[3]/NET0131  , \rd1_R_o_reg[4]/NET0131  , \rd1_R_o_reg[5]/NET0131  , \rd1_R_o_reg[6]/NET0131  , \rd1_R_o_reg[7]/NET0131  , \rd1_R_o_reg[8]/NET0131  , \rd1_R_o_reg[9]/NET0131  , \stage1_iter_reg[0]/NET0131  , \stage1_iter_reg[1]/NET0131  , \stage1_iter_reg[2]/NET0131  , \stage1_iter_reg[3]/NET0131  , \_al_n0  , \_al_n1  , \g10087/_0_  , \g10220/_1_  , \g11117/_0_  , \g11124/_0_  , \g11125/_0_  , \g11170/_0_  , \g11182/_0_  , \g11184/_0_  , \g11378/_0_  , \g11393/_0_  , \g11415/_0_  , \g11432/_0_  , \g11433/_0_  , \g11453/_0_  , \g11500/_0_  , \g11588/_0_  , \g11607/_0_  , \g11616/_0_  , \g11625/_0_  , \g11641_dup/_0_  , \g11648/_0_  , \g11655/_0_  , \g11683/_0_  , \g11689/_2_  , \g11694/_0_  , \g11748/_0_  , \g11880/_0_  , \g11962/_1_  , \g12016/_0_  , \g12038/_0_  , \g12039/_0_  , \g12094/_0_  , \g12100/_0_  , \g12132/_0_  , \g12151/_0_  , \g12251/_0_  , \g12279/_0_  , \g12288/_0_  , \g12290/_0_  , \g12311/_0_  , \g12313/_0_  , \g12356/_0_  , \g12357/_0_  , \g12427/_0_  , \g12441/_0_  , \g12442/_0_  , \g12480/_0_  , \g12485/_0_  , \g12506/_0_  , \g12544/_0_  , \g12549/_2_  , \g12614/_0_  , \g12678/_0_  , \g12680/_0_  , \g12748/_0_  , \g15/_0_  , \g25/_0_  , \g31/_0_  , \g6843/_0_  , \g6861/_0_  , \g6863/_0_  , \g6865/_0_  , \g6887/_0_  , \g6888/_0_  , \g6889/_0_  , \g6890/_0_  , \g6891/_0_  , \g6892/_0_  , \g6893/_0_  , \g6894/_0_  , \g6922/_0_  , \g6923/_0_  , \g6924/_3_  , \g6926/_0_  , \g6927/_0_  , \g6928/_0_  , \g6931/_0_  , \g6933/_0_  , \g6967/_0_  , \g6968/_0_  , \g6969/_0_  , \g6974/_0_  , \g6975/_0_  , \g6976/_3_  , \g7006/_3_  , \g8882/_0_  , \g8883/_0_  , \g8884/_0_  , \g8895/_0_  , \g8896/_0_  , \g8898/_0_  , \g8900/_2_  , \g8902/_0_  , \g8907/_0_  , \g8911/_0_  , \g8924/_0_  , \g8927/_0_  , \g8929/_2_  , \g8967/_0_  , \g8969/_0_  , \g8973/_2_  , \g8987/_0_  , \g8989/_0_  , \g8991/_0_  , \g8996/_0_  , \g9099/_0_  , \g9543/_1_  , \g9751/_1_  , \g9755/_0_  , \g9786/_0_  , \g9794/_0_  , \g9817/_0_  , \g9836/_0_  , \g9859/_0_  , \g9862/_0_  , \g9867/_0_  , \g9869/_0_  , \g9876/_0_  , \g9887/_0_  , \g9895/_0_  , \g9897/_0_  , \g9908/_0_  , \g9910/_0_  , \g9915/_0_  , \g9938/_0_  , \g9970/_0_  );
  input \data_i[0]_pad  ;
  input \data_i[10]_pad  ;
  input \data_i[11]_pad  ;
  input \data_i[12]_pad  ;
  input \data_i[13]_pad  ;
  input \data_i[14]_pad  ;
  input \data_i[15]_pad  ;
  input \data_i[16]_pad  ;
  input \data_i[17]_pad  ;
  input \data_i[18]_pad  ;
  input \data_i[19]_pad  ;
  input \data_i[1]_pad  ;
  input \data_i[20]_pad  ;
  input \data_i[21]_pad  ;
  input \data_i[22]_pad  ;
  input \data_i[23]_pad  ;
  input \data_i[24]_pad  ;
  input \data_i[25]_pad  ;
  input \data_i[26]_pad  ;
  input \data_i[27]_pad  ;
  input \data_i[28]_pad  ;
  input \data_i[29]_pad  ;
  input \data_i[2]_pad  ;
  input \data_i[30]_pad  ;
  input \data_i[31]_pad  ;
  input \data_i[32]_pad  ;
  input \data_i[33]_pad  ;
  input \data_i[34]_pad  ;
  input \data_i[35]_pad  ;
  input \data_i[36]_pad  ;
  input \data_i[37]_pad  ;
  input \data_i[38]_pad  ;
  input \data_i[39]_pad  ;
  input \data_i[3]_pad  ;
  input \data_i[40]_pad  ;
  input \data_i[41]_pad  ;
  input \data_i[42]_pad  ;
  input \data_i[43]_pad  ;
  input \data_i[44]_pad  ;
  input \data_i[45]_pad  ;
  input \data_i[46]_pad  ;
  input \data_i[47]_pad  ;
  input \data_i[48]_pad  ;
  input \data_i[49]_pad  ;
  input \data_i[4]_pad  ;
  input \data_i[50]_pad  ;
  input \data_i[51]_pad  ;
  input \data_i[52]_pad  ;
  input \data_i[53]_pad  ;
  input \data_i[54]_pad  ;
  input \data_i[55]_pad  ;
  input \data_i[56]_pad  ;
  input \data_i[57]_pad  ;
  input \data_i[58]_pad  ;
  input \data_i[59]_pad  ;
  input \data_i[5]_pad  ;
  input \data_i[60]_pad  ;
  input \data_i[61]_pad  ;
  input \data_i[62]_pad  ;
  input \data_i[63]_pad  ;
  input \data_i[6]_pad  ;
  input \data_i[7]_pad  ;
  input \data_i[8]_pad  ;
  input \data_i[9]_pad  ;
  input \data_ready_reg/NET0131  ;
  input decrypt_i_pad ;
  input \key_i[10]_pad  ;
  input \key_i[11]_pad  ;
  input \key_i[12]_pad  ;
  input \key_i[13]_pad  ;
  input \key_i[14]_pad  ;
  input \key_i[15]_pad  ;
  input \key_i[17]_pad  ;
  input \key_i[18]_pad  ;
  input \key_i[19]_pad  ;
  input \key_i[1]_pad  ;
  input \key_i[20]_pad  ;
  input \key_i[21]_pad  ;
  input \key_i[22]_pad  ;
  input \key_i[23]_pad  ;
  input \key_i[25]_pad  ;
  input \key_i[26]_pad  ;
  input \key_i[27]_pad  ;
  input \key_i[28]_pad  ;
  input \key_i[29]_pad  ;
  input \key_i[2]_pad  ;
  input \key_i[30]_pad  ;
  input \key_i[31]_pad  ;
  input \key_i[33]_pad  ;
  input \key_i[34]_pad  ;
  input \key_i[35]_pad  ;
  input \key_i[36]_pad  ;
  input \key_i[37]_pad  ;
  input \key_i[38]_pad  ;
  input \key_i[39]_pad  ;
  input \key_i[3]_pad  ;
  input \key_i[41]_pad  ;
  input \key_i[42]_pad  ;
  input \key_i[43]_pad  ;
  input \key_i[44]_pad  ;
  input \key_i[45]_pad  ;
  input \key_i[46]_pad  ;
  input \key_i[47]_pad  ;
  input \key_i[49]_pad  ;
  input \key_i[4]_pad  ;
  input \key_i[50]_pad  ;
  input \key_i[51]_pad  ;
  input \key_i[52]_pad  ;
  input \key_i[53]_pad  ;
  input \key_i[54]_pad  ;
  input \key_i[55]_pad  ;
  input \key_i[57]_pad  ;
  input \key_i[58]_pad  ;
  input \key_i[59]_pad  ;
  input \key_i[5]_pad  ;
  input \key_i[60]_pad  ;
  input \key_i[61]_pad  ;
  input \key_i[62]_pad  ;
  input \key_i[63]_pad  ;
  input \key_i[6]_pad  ;
  input \key_i[7]_pad  ;
  input \key_i[9]_pad  ;
  input load_i_pad ;
  input \rd1_Key_o_reg[0]/NET0131  ;
  input \rd1_Key_o_reg[10]/NET0131  ;
  input \rd1_Key_o_reg[11]/NET0131  ;
  input \rd1_Key_o_reg[12]/NET0131  ;
  input \rd1_Key_o_reg[13]/NET0131  ;
  input \rd1_Key_o_reg[14]/NET0131  ;
  input \rd1_Key_o_reg[15]/NET0131  ;
  input \rd1_Key_o_reg[16]/NET0131  ;
  input \rd1_Key_o_reg[17]/NET0131  ;
  input \rd1_Key_o_reg[18]/NET0131  ;
  input \rd1_Key_o_reg[19]/NET0131  ;
  input \rd1_Key_o_reg[1]/NET0131  ;
  input \rd1_Key_o_reg[20]/NET0131  ;
  input \rd1_Key_o_reg[21]/NET0131  ;
  input \rd1_Key_o_reg[22]/NET0131  ;
  input \rd1_Key_o_reg[23]/NET0131  ;
  input \rd1_Key_o_reg[24]/NET0131  ;
  input \rd1_Key_o_reg[25]/NET0131  ;
  input \rd1_Key_o_reg[26]/NET0131  ;
  input \rd1_Key_o_reg[27]/NET0131  ;
  input \rd1_Key_o_reg[28]/NET0131  ;
  input \rd1_Key_o_reg[29]/NET0131  ;
  input \rd1_Key_o_reg[2]/NET0131  ;
  input \rd1_Key_o_reg[30]/NET0131  ;
  input \rd1_Key_o_reg[31]/NET0131  ;
  input \rd1_Key_o_reg[32]/NET0131  ;
  input \rd1_Key_o_reg[33]/NET0131  ;
  input \rd1_Key_o_reg[34]/NET0131  ;
  input \rd1_Key_o_reg[35]/NET0131  ;
  input \rd1_Key_o_reg[36]/NET0131  ;
  input \rd1_Key_o_reg[37]/NET0131  ;
  input \rd1_Key_o_reg[38]/NET0131  ;
  input \rd1_Key_o_reg[39]/NET0131  ;
  input \rd1_Key_o_reg[3]/NET0131  ;
  input \rd1_Key_o_reg[40]/NET0131  ;
  input \rd1_Key_o_reg[41]/NET0131  ;
  input \rd1_Key_o_reg[42]/NET0131  ;
  input \rd1_Key_o_reg[43]/NET0131  ;
  input \rd1_Key_o_reg[44]/NET0131  ;
  input \rd1_Key_o_reg[45]/NET0131  ;
  input \rd1_Key_o_reg[46]/NET0131  ;
  input \rd1_Key_o_reg[47]/NET0131  ;
  input \rd1_Key_o_reg[48]/NET0131  ;
  input \rd1_Key_o_reg[49]/NET0131  ;
  input \rd1_Key_o_reg[4]/NET0131  ;
  input \rd1_Key_o_reg[50]/NET0131  ;
  input \rd1_Key_o_reg[51]/NET0131  ;
  input \rd1_Key_o_reg[52]/NET0131  ;
  input \rd1_Key_o_reg[53]/NET0131  ;
  input \rd1_Key_o_reg[54]/NET0131  ;
  input \rd1_Key_o_reg[55]/NET0131  ;
  input \rd1_Key_o_reg[5]/NET0131  ;
  input \rd1_Key_o_reg[6]/NET0131  ;
  input \rd1_Key_o_reg[7]/NET0131  ;
  input \rd1_Key_o_reg[8]/NET0131  ;
  input \rd1_Key_o_reg[9]/NET0131  ;
  input \rd1_L_o_reg[0]/NET0131  ;
  input \rd1_L_o_reg[10]/NET0131  ;
  input \rd1_L_o_reg[11]/NET0131  ;
  input \rd1_L_o_reg[12]/NET0131  ;
  input \rd1_L_o_reg[13]/NET0131  ;
  input \rd1_L_o_reg[14]/NET0131  ;
  input \rd1_L_o_reg[15]/NET0131  ;
  input \rd1_L_o_reg[16]/NET0131  ;
  input \rd1_L_o_reg[17]/NET0131  ;
  input \rd1_L_o_reg[18]/NET0131  ;
  input \rd1_L_o_reg[19]/NET0131  ;
  input \rd1_L_o_reg[1]/NET0131  ;
  input \rd1_L_o_reg[20]/NET0131  ;
  input \rd1_L_o_reg[21]/NET0131  ;
  input \rd1_L_o_reg[22]/NET0131  ;
  input \rd1_L_o_reg[23]/NET0131  ;
  input \rd1_L_o_reg[24]/NET0131  ;
  input \rd1_L_o_reg[25]/NET0131  ;
  input \rd1_L_o_reg[26]/NET0131  ;
  input \rd1_L_o_reg[27]/NET0131  ;
  input \rd1_L_o_reg[28]/NET0131  ;
  input \rd1_L_o_reg[29]/NET0131  ;
  input \rd1_L_o_reg[2]/NET0131  ;
  input \rd1_L_o_reg[30]/NET0131  ;
  input \rd1_L_o_reg[31]/NET0131  ;
  input \rd1_L_o_reg[3]/NET0131  ;
  input \rd1_L_o_reg[4]/NET0131  ;
  input \rd1_L_o_reg[5]/NET0131  ;
  input \rd1_L_o_reg[6]/NET0131  ;
  input \rd1_L_o_reg[7]/NET0131  ;
  input \rd1_L_o_reg[8]/NET0131  ;
  input \rd1_L_o_reg[9]/NET0131  ;
  input \rd1_R_o_reg[0]/NET0131  ;
  input \rd1_R_o_reg[10]/NET0131  ;
  input \rd1_R_o_reg[11]/NET0131  ;
  input \rd1_R_o_reg[12]/NET0131  ;
  input \rd1_R_o_reg[13]/NET0131  ;
  input \rd1_R_o_reg[14]/NET0131  ;
  input \rd1_R_o_reg[15]/NET0131  ;
  input \rd1_R_o_reg[16]/NET0131  ;
  input \rd1_R_o_reg[17]/NET0131  ;
  input \rd1_R_o_reg[18]/NET0131  ;
  input \rd1_R_o_reg[19]/NET0131  ;
  input \rd1_R_o_reg[1]/NET0131  ;
  input \rd1_R_o_reg[20]/NET0131  ;
  input \rd1_R_o_reg[21]/NET0131  ;
  input \rd1_R_o_reg[22]/NET0131  ;
  input \rd1_R_o_reg[23]/NET0131  ;
  input \rd1_R_o_reg[24]/NET0131  ;
  input \rd1_R_o_reg[25]/NET0131  ;
  input \rd1_R_o_reg[26]/NET0131  ;
  input \rd1_R_o_reg[27]/NET0131  ;
  input \rd1_R_o_reg[28]/NET0131  ;
  input \rd1_R_o_reg[29]/NET0131  ;
  input \rd1_R_o_reg[2]/NET0131  ;
  input \rd1_R_o_reg[30]/NET0131  ;
  input \rd1_R_o_reg[31]/NET0131  ;
  input \rd1_R_o_reg[3]/NET0131  ;
  input \rd1_R_o_reg[4]/NET0131  ;
  input \rd1_R_o_reg[5]/NET0131  ;
  input \rd1_R_o_reg[6]/NET0131  ;
  input \rd1_R_o_reg[7]/NET0131  ;
  input \rd1_R_o_reg[8]/NET0131  ;
  input \rd1_R_o_reg[9]/NET0131  ;
  input \stage1_iter_reg[0]/NET0131  ;
  input \stage1_iter_reg[1]/NET0131  ;
  input \stage1_iter_reg[2]/NET0131  ;
  input \stage1_iter_reg[3]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g10087/_0_  ;
  output \g10220/_1_  ;
  output \g11117/_0_  ;
  output \g11124/_0_  ;
  output \g11125/_0_  ;
  output \g11170/_0_  ;
  output \g11182/_0_  ;
  output \g11184/_0_  ;
  output \g11378/_0_  ;
  output \g11393/_0_  ;
  output \g11415/_0_  ;
  output \g11432/_0_  ;
  output \g11433/_0_  ;
  output \g11453/_0_  ;
  output \g11500/_0_  ;
  output \g11588/_0_  ;
  output \g11607/_0_  ;
  output \g11616/_0_  ;
  output \g11625/_0_  ;
  output \g11641_dup/_0_  ;
  output \g11648/_0_  ;
  output \g11655/_0_  ;
  output \g11683/_0_  ;
  output \g11689/_2_  ;
  output \g11694/_0_  ;
  output \g11748/_0_  ;
  output \g11880/_0_  ;
  output \g11962/_1_  ;
  output \g12016/_0_  ;
  output \g12038/_0_  ;
  output \g12039/_0_  ;
  output \g12094/_0_  ;
  output \g12100/_0_  ;
  output \g12132/_0_  ;
  output \g12151/_0_  ;
  output \g12251/_0_  ;
  output \g12279/_0_  ;
  output \g12288/_0_  ;
  output \g12290/_0_  ;
  output \g12311/_0_  ;
  output \g12313/_0_  ;
  output \g12356/_0_  ;
  output \g12357/_0_  ;
  output \g12427/_0_  ;
  output \g12441/_0_  ;
  output \g12442/_0_  ;
  output \g12480/_0_  ;
  output \g12485/_0_  ;
  output \g12506/_0_  ;
  output \g12544/_0_  ;
  output \g12549/_2_  ;
  output \g12614/_0_  ;
  output \g12678/_0_  ;
  output \g12680/_0_  ;
  output \g12748/_0_  ;
  output \g15/_0_  ;
  output \g25/_0_  ;
  output \g31/_0_  ;
  output \g6843/_0_  ;
  output \g6861/_0_  ;
  output \g6863/_0_  ;
  output \g6865/_0_  ;
  output \g6887/_0_  ;
  output \g6888/_0_  ;
  output \g6889/_0_  ;
  output \g6890/_0_  ;
  output \g6891/_0_  ;
  output \g6892/_0_  ;
  output \g6893/_0_  ;
  output \g6894/_0_  ;
  output \g6922/_0_  ;
  output \g6923/_0_  ;
  output \g6924/_3_  ;
  output \g6926/_0_  ;
  output \g6927/_0_  ;
  output \g6928/_0_  ;
  output \g6931/_0_  ;
  output \g6933/_0_  ;
  output \g6967/_0_  ;
  output \g6968/_0_  ;
  output \g6969/_0_  ;
  output \g6974/_0_  ;
  output \g6975/_0_  ;
  output \g6976/_3_  ;
  output \g7006/_3_  ;
  output \g8882/_0_  ;
  output \g8883/_0_  ;
  output \g8884/_0_  ;
  output \g8895/_0_  ;
  output \g8896/_0_  ;
  output \g8898/_0_  ;
  output \g8900/_2_  ;
  output \g8902/_0_  ;
  output \g8907/_0_  ;
  output \g8911/_0_  ;
  output \g8924/_0_  ;
  output \g8927/_0_  ;
  output \g8929/_2_  ;
  output \g8967/_0_  ;
  output \g8969/_0_  ;
  output \g8973/_2_  ;
  output \g8987/_0_  ;
  output \g8989/_0_  ;
  output \g8991/_0_  ;
  output \g8996/_0_  ;
  output \g9099/_0_  ;
  output \g9543/_1_  ;
  output \g9751/_1_  ;
  output \g9755/_0_  ;
  output \g9786/_0_  ;
  output \g9794/_0_  ;
  output \g9817/_0_  ;
  output \g9836/_0_  ;
  output \g9859/_0_  ;
  output \g9862/_0_  ;
  output \g9867/_0_  ;
  output \g9869/_0_  ;
  output \g9876/_0_  ;
  output \g9887/_0_  ;
  output \g9895/_0_  ;
  output \g9897/_0_  ;
  output \g9908/_0_  ;
  output \g9910/_0_  ;
  output \g9915/_0_  ;
  output \g9938/_0_  ;
  output \g9970/_0_  ;
  wire n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 ;
  assign n248 = ~\stage1_iter_reg[1]/NET0131  & ~\stage1_iter_reg[2]/NET0131  ;
  assign n249 = ~\stage1_iter_reg[0]/NET0131  & ~\stage1_iter_reg[3]/NET0131  ;
  assign n250 = n248 & n249 ;
  assign n251 = ~\data_ready_reg/NET0131  & ~load_i_pad ;
  assign n252 = n250 & n251 ;
  assign n253 = ~\stage1_iter_reg[0]/NET0131  & ~\stage1_iter_reg[1]/NET0131  ;
  assign n254 = \stage1_iter_reg[0]/NET0131  & \stage1_iter_reg[1]/NET0131  ;
  assign n255 = ~n253 & ~n254 ;
  assign n256 = \rd1_Key_o_reg[26]/NET0131  & ~n250 ;
  assign n257 = ~load_i_pad & ~\rd1_Key_o_reg[26]/NET0131  ;
  assign n258 = ~\key_i[9]_pad  & load_i_pad ;
  assign n259 = ~n257 & ~n258 ;
  assign n260 = n250 & n259 ;
  assign n261 = ~n256 & ~n260 ;
  assign n262 = \stage1_iter_reg[2]/NET0131  & n254 ;
  assign n263 = \stage1_iter_reg[3]/NET0131  & n262 ;
  assign n264 = \stage1_iter_reg[0]/NET0131  & \stage1_iter_reg[3]/NET0131  ;
  assign n265 = n248 & ~n264 ;
  assign n266 = ~n263 & ~n265 ;
  assign n267 = ~n261 & ~n266 ;
  assign n268 = \rd1_Key_o_reg[25]/NET0131  & ~n250 ;
  assign n269 = ~load_i_pad & ~\rd1_Key_o_reg[25]/NET0131  ;
  assign n270 = ~\key_i[17]_pad  & load_i_pad ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = n250 & n271 ;
  assign n273 = ~n268 & ~n272 ;
  assign n274 = n266 & ~n273 ;
  assign n275 = ~n267 & ~n274 ;
  assign n276 = ~decrypt_i_pad & ~n275 ;
  assign n286 = \rd1_Key_o_reg[0]/NET0131  & ~n250 ;
  assign n287 = ~load_i_pad & ~\rd1_Key_o_reg[0]/NET0131  ;
  assign n288 = ~\key_i[60]_pad  & load_i_pad ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = n250 & n289 ;
  assign n291 = ~n286 & ~n290 ;
  assign n292 = ~n249 & ~n266 ;
  assign n293 = ~n291 & n292 ;
  assign n277 = ~load_i_pad & ~\rd1_Key_o_reg[27]/NET0131  ;
  assign n278 = ~\key_i[1]_pad  & load_i_pad ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = n250 & n279 ;
  assign n281 = load_i_pad & n250 ;
  assign n282 = \rd1_Key_o_reg[1]/NET0131  & ~n281 ;
  assign n283 = \key_i[52]_pad  & n281 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n266 & ~n284 ;
  assign n294 = ~n280 & ~n285 ;
  assign n295 = ~n293 & n294 ;
  assign n296 = decrypt_i_pad & ~n295 ;
  assign n297 = ~n276 & ~n296 ;
  assign n298 = \rd1_R_o_reg[10]/NET0131  & ~n281 ;
  assign n299 = \data_i[43]_pad  & n281 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = \rd1_Key_o_reg[3]/NET0131  & ~n281 ;
  assign n302 = \key_i[36]_pad  & n281 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = n266 & ~n303 ;
  assign n305 = \rd1_Key_o_reg[4]/NET0131  & ~n250 ;
  assign n306 = ~load_i_pad & ~\rd1_Key_o_reg[4]/NET0131  ;
  assign n307 = ~\key_i[59]_pad  & load_i_pad ;
  assign n308 = ~n306 & ~n307 ;
  assign n309 = n250 & n308 ;
  assign n310 = ~n305 & ~n309 ;
  assign n311 = ~n266 & ~n310 ;
  assign n312 = ~n304 & ~n311 ;
  assign n313 = ~decrypt_i_pad & ~n312 ;
  assign n325 = \rd1_Key_o_reg[6]/NET0131  & ~n250 ;
  assign n326 = ~load_i_pad & ~\rd1_Key_o_reg[6]/NET0131  ;
  assign n327 = ~\key_i[43]_pad  & load_i_pad ;
  assign n328 = ~n326 & ~n327 ;
  assign n329 = n250 & n328 ;
  assign n330 = ~n325 & ~n329 ;
  assign n331 = n292 & ~n330 ;
  assign n314 = \rd1_Key_o_reg[5]/NET0131  & ~n281 ;
  assign n315 = \key_i[51]_pad  & n281 ;
  assign n316 = ~n314 & ~n315 ;
  assign n317 = n250 & ~n316 ;
  assign n318 = \rd1_Key_o_reg[7]/NET0131  & ~n250 ;
  assign n319 = ~load_i_pad & ~\rd1_Key_o_reg[7]/NET0131  ;
  assign n320 = ~\key_i[35]_pad  & load_i_pad ;
  assign n321 = ~n319 & ~n320 ;
  assign n322 = n250 & n321 ;
  assign n323 = ~n318 & ~n322 ;
  assign n324 = n266 & ~n323 ;
  assign n332 = ~n317 & ~n324 ;
  assign n333 = ~n331 & n332 ;
  assign n334 = decrypt_i_pad & ~n333 ;
  assign n335 = ~n313 & ~n334 ;
  assign n336 = \rd1_Key_o_reg[28]/NET0131  & ~n250 ;
  assign n337 = ~load_i_pad & ~\rd1_Key_o_reg[28]/NET0131  ;
  assign n338 = ~\key_i[28]_pad  & load_i_pad ;
  assign n339 = ~n337 & ~n338 ;
  assign n340 = n250 & n339 ;
  assign n341 = ~n336 & ~n340 ;
  assign n342 = ~n266 & ~n341 ;
  assign n343 = \rd1_Key_o_reg[55]/NET0131  & ~n250 ;
  assign n344 = ~\key_i[7]_pad  & load_i_pad ;
  assign n345 = ~load_i_pad & ~\rd1_Key_o_reg[55]/NET0131  ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = n250 & n346 ;
  assign n348 = ~n343 & ~n347 ;
  assign n349 = n266 & ~n348 ;
  assign n350 = ~n342 & ~n349 ;
  assign n351 = ~decrypt_i_pad & ~n350 ;
  assign n363 = \rd1_Key_o_reg[30]/NET0131  & ~n250 ;
  assign n364 = ~\key_i[12]_pad  & load_i_pad ;
  assign n365 = ~load_i_pad & ~\rd1_Key_o_reg[30]/NET0131  ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = n250 & n366 ;
  assign n368 = ~n363 & ~n367 ;
  assign n369 = n292 & ~n368 ;
  assign n352 = ~load_i_pad & ~\rd1_Key_o_reg[29]/NET0131  ;
  assign n353 = ~\key_i[20]_pad  & load_i_pad ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = n250 & n354 ;
  assign n356 = \rd1_Key_o_reg[31]/NET0131  & ~n250 ;
  assign n357 = ~load_i_pad & ~\rd1_Key_o_reg[31]/NET0131  ;
  assign n358 = ~\key_i[4]_pad  & load_i_pad ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = n250 & n359 ;
  assign n361 = ~n356 & ~n360 ;
  assign n362 = n266 & ~n361 ;
  assign n370 = ~n355 & ~n362 ;
  assign n371 = ~n369 & n370 ;
  assign n372 = decrypt_i_pad & ~n371 ;
  assign n373 = ~n351 & ~n372 ;
  assign n374 = \rd1_R_o_reg[4]/NET0131  & ~n281 ;
  assign n375 = \data_i[25]_pad  & n281 ;
  assign n376 = ~n374 & ~n375 ;
  assign n377 = \rd1_Key_o_reg[21]/NET0131  & ~n250 ;
  assign n378 = ~load_i_pad & ~\rd1_Key_o_reg[21]/NET0131  ;
  assign n379 = ~\key_i[49]_pad  & load_i_pad ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = n250 & n380 ;
  assign n382 = ~n377 & ~n381 ;
  assign n383 = ~n266 & ~n382 ;
  assign n384 = \rd1_Key_o_reg[20]/NET0131  & ~n250 ;
  assign n385 = ~load_i_pad & ~\rd1_Key_o_reg[20]/NET0131  ;
  assign n386 = ~\key_i[57]_pad  & load_i_pad ;
  assign n387 = ~n385 & ~n386 ;
  assign n388 = n250 & n387 ;
  assign n389 = ~n384 & ~n388 ;
  assign n390 = n266 & ~n389 ;
  assign n391 = ~n383 & ~n390 ;
  assign n392 = ~decrypt_i_pad & ~n391 ;
  assign n400 = \rd1_Key_o_reg[23]/NET0131  & ~n281 ;
  assign n401 = \key_i[33]_pad  & n281 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = n292 & ~n402 ;
  assign n393 = \rd1_Key_o_reg[24]/NET0131  & ~n250 ;
  assign n394 = ~load_i_pad & ~\rd1_Key_o_reg[24]/NET0131  ;
  assign n395 = ~\key_i[25]_pad  & load_i_pad ;
  assign n396 = ~n394 & ~n395 ;
  assign n397 = n250 & n396 ;
  assign n398 = ~n393 & ~n397 ;
  assign n399 = n266 & ~n398 ;
  assign n404 = ~load_i_pad & ~\rd1_Key_o_reg[22]/NET0131  ;
  assign n405 = ~\key_i[41]_pad  & load_i_pad ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = n250 & n406 ;
  assign n408 = ~n399 & ~n407 ;
  assign n409 = ~n403 & n408 ;
  assign n410 = decrypt_i_pad & ~n409 ;
  assign n411 = ~n392 & ~n410 ;
  assign n412 = ~n266 & ~n330 ;
  assign n413 = n266 & ~n316 ;
  assign n414 = ~n412 & ~n413 ;
  assign n415 = ~decrypt_i_pad & ~n414 ;
  assign n420 = \rd1_Key_o_reg[8]/NET0131  & ~n281 ;
  assign n421 = \key_i[27]_pad  & n281 ;
  assign n422 = ~n420 & ~n421 ;
  assign n423 = n292 & ~n422 ;
  assign n416 = \rd1_Key_o_reg[9]/NET0131  & ~n281 ;
  assign n417 = \key_i[19]_pad  & n281 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = n266 & ~n418 ;
  assign n424 = ~n322 & ~n419 ;
  assign n425 = ~n423 & n424 ;
  assign n426 = decrypt_i_pad & ~n425 ;
  assign n427 = ~n415 & ~n426 ;
  assign n428 = \rd1_Key_o_reg[10]/NET0131  & ~n250 ;
  assign n429 = ~load_i_pad & ~\rd1_Key_o_reg[10]/NET0131  ;
  assign n430 = ~\key_i[11]_pad  & load_i_pad ;
  assign n431 = ~n429 & ~n430 ;
  assign n432 = n250 & n431 ;
  assign n433 = ~n428 & ~n432 ;
  assign n434 = ~n266 & ~n433 ;
  assign n435 = ~n419 & ~n434 ;
  assign n436 = ~decrypt_i_pad & ~n435 ;
  assign n441 = \rd1_Key_o_reg[13]/NET0131  & ~n281 ;
  assign n442 = \key_i[50]_pad  & n281 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = n266 & ~n443 ;
  assign n437 = \rd1_Key_o_reg[12]/NET0131  & ~n281 ;
  assign n438 = \key_i[58]_pad  & n281 ;
  assign n439 = ~n437 & ~n438 ;
  assign n440 = n292 & ~n439 ;
  assign n445 = ~load_i_pad & ~\rd1_Key_o_reg[11]/NET0131  ;
  assign n446 = ~\key_i[3]_pad  & load_i_pad ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = n250 & n447 ;
  assign n449 = ~n440 & ~n448 ;
  assign n450 = ~n444 & n449 ;
  assign n451 = decrypt_i_pad & ~n450 ;
  assign n452 = ~n436 & ~n451 ;
  assign n453 = \rd1_Key_o_reg[29]/NET0131  & ~n250 ;
  assign n454 = ~n355 & ~n453 ;
  assign n455 = ~n266 & ~n454 ;
  assign n456 = n266 & ~n341 ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = ~decrypt_i_pad & ~n457 ;
  assign n466 = n292 & ~n361 ;
  assign n459 = \rd1_Key_o_reg[32]/NET0131  & ~n250 ;
  assign n460 = ~load_i_pad & ~\rd1_Key_o_reg[32]/NET0131  ;
  assign n461 = ~\key_i[61]_pad  & load_i_pad ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = n250 & n462 ;
  assign n464 = ~n459 & ~n463 ;
  assign n465 = n266 & ~n464 ;
  assign n467 = ~n367 & ~n465 ;
  assign n468 = ~n466 & n467 ;
  assign n469 = decrypt_i_pad & ~n468 ;
  assign n470 = ~n458 & ~n469 ;
  assign n471 = ~n266 & ~n361 ;
  assign n472 = n266 & ~n368 ;
  assign n473 = ~n471 & ~n472 ;
  assign n474 = ~decrypt_i_pad & ~n473 ;
  assign n482 = \rd1_Key_o_reg[33]/NET0131  & ~n281 ;
  assign n483 = \key_i[53]_pad  & n281 ;
  assign n484 = ~n482 & ~n483 ;
  assign n485 = n292 & ~n484 ;
  assign n475 = \rd1_Key_o_reg[34]/NET0131  & ~n250 ;
  assign n476 = ~load_i_pad & ~\rd1_Key_o_reg[34]/NET0131  ;
  assign n477 = ~\key_i[45]_pad  & load_i_pad ;
  assign n478 = ~n476 & ~n477 ;
  assign n479 = n250 & n478 ;
  assign n480 = ~n475 & ~n479 ;
  assign n481 = n266 & ~n480 ;
  assign n486 = ~n463 & ~n481 ;
  assign n487 = ~n485 & n486 ;
  assign n488 = decrypt_i_pad & ~n487 ;
  assign n489 = ~n474 & ~n488 ;
  assign n490 = \rd1_R_o_reg[29]/NET0131  & ~n281 ;
  assign n491 = \data_i[23]_pad  & n281 ;
  assign n492 = ~n490 & ~n491 ;
  assign n495 = n250 & ~n418 ;
  assign n493 = n292 & ~n418 ;
  assign n494 = n266 & ~n422 ;
  assign n496 = ~n493 & ~n494 ;
  assign n497 = ~n495 & n496 ;
  assign n498 = ~decrypt_i_pad & ~n497 ;
  assign n500 = \rd1_Key_o_reg[11]/NET0131  & ~n250 ;
  assign n501 = ~n448 & ~n500 ;
  assign n502 = n292 & ~n501 ;
  assign n499 = n266 & ~n439 ;
  assign n503 = ~n432 & ~n499 ;
  assign n504 = ~n502 & n503 ;
  assign n505 = decrypt_i_pad & ~n504 ;
  assign n506 = ~n498 & ~n505 ;
  assign n507 = ~n266 & ~n464 ;
  assign n508 = ~n362 & ~n507 ;
  assign n509 = ~decrypt_i_pad & ~n508 ;
  assign n518 = n292 & ~n480 ;
  assign n510 = n250 & ~n484 ;
  assign n511 = \rd1_Key_o_reg[35]/NET0131  & ~n250 ;
  assign n512 = ~load_i_pad & ~\rd1_Key_o_reg[35]/NET0131  ;
  assign n513 = ~\key_i[37]_pad  & load_i_pad ;
  assign n514 = ~n512 & ~n513 ;
  assign n515 = n250 & n514 ;
  assign n516 = ~n511 & ~n515 ;
  assign n517 = n266 & ~n516 ;
  assign n519 = ~n510 & ~n517 ;
  assign n520 = ~n518 & n519 ;
  assign n521 = decrypt_i_pad & ~n520 ;
  assign n522 = ~n509 & ~n521 ;
  assign n523 = \rd1_Key_o_reg[22]/NET0131  & ~n250 ;
  assign n524 = ~n407 & ~n523 ;
  assign n525 = ~n266 & ~n524 ;
  assign n526 = n266 & ~n382 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = ~decrypt_i_pad & ~n527 ;
  assign n530 = n292 & ~n398 ;
  assign n529 = n250 & ~n402 ;
  assign n531 = ~n274 & ~n529 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = decrypt_i_pad & ~n532 ;
  assign n534 = ~n528 & ~n533 ;
  assign n535 = ~n266 & ~n291 ;
  assign n536 = \rd1_Key_o_reg[27]/NET0131  & ~n250 ;
  assign n537 = n266 & n536 ;
  assign n538 = ~n535 & ~n537 ;
  assign n539 = ~decrypt_i_pad & ~n538 ;
  assign n541 = \rd1_Key_o_reg[2]/NET0131  & ~n250 ;
  assign n542 = ~load_i_pad & ~\rd1_Key_o_reg[2]/NET0131  ;
  assign n543 = ~\key_i[44]_pad  & load_i_pad ;
  assign n544 = ~n542 & ~n543 ;
  assign n545 = n250 & n544 ;
  assign n546 = ~n541 & ~n545 ;
  assign n547 = n292 & ~n546 ;
  assign n540 = n250 & ~n284 ;
  assign n548 = ~n304 & ~n540 ;
  assign n549 = ~n547 & n548 ;
  assign n550 = decrypt_i_pad & ~n549 ;
  assign n551 = ~n539 & ~n550 ;
  assign n563 = \rd1_Key_o_reg[49]/NET0131  & ~n250 ;
  assign n564 = ~load_i_pad & ~\rd1_Key_o_reg[49]/NET0131  ;
  assign n565 = ~\key_i[55]_pad  & load_i_pad ;
  assign n566 = ~n564 & ~n565 ;
  assign n567 = n250 & n566 ;
  assign n568 = ~n563 & ~n567 ;
  assign n569 = n292 & ~n568 ;
  assign n552 = ~load_i_pad & ~\rd1_Key_o_reg[48]/NET0131  ;
  assign n553 = ~\key_i[63]_pad  & load_i_pad ;
  assign n554 = ~n552 & ~n553 ;
  assign n555 = n250 & n554 ;
  assign n556 = \rd1_Key_o_reg[50]/NET0131  & ~n250 ;
  assign n557 = ~load_i_pad & ~\rd1_Key_o_reg[50]/NET0131  ;
  assign n558 = ~\key_i[47]_pad  & load_i_pad ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = n250 & n559 ;
  assign n561 = ~n556 & ~n560 ;
  assign n562 = n266 & ~n561 ;
  assign n570 = ~n555 & ~n562 ;
  assign n571 = ~n569 & n570 ;
  assign n572 = decrypt_i_pad & ~n571 ;
  assign n573 = \rd1_Key_o_reg[47]/NET0131  & ~n281 ;
  assign n574 = \key_i[6]_pad  & n281 ;
  assign n575 = ~n573 & ~n574 ;
  assign n581 = n292 & ~n575 ;
  assign n576 = n250 & ~n575 ;
  assign n577 = \rd1_Key_o_reg[46]/NET0131  & ~n281 ;
  assign n578 = \key_i[14]_pad  & n281 ;
  assign n579 = ~n577 & ~n578 ;
  assign n580 = n266 & ~n579 ;
  assign n582 = ~n576 & ~n580 ;
  assign n583 = ~n581 & n582 ;
  assign n584 = ~decrypt_i_pad & ~n583 ;
  assign n585 = ~n572 & ~n584 ;
  assign n586 = \rd1_R_o_reg[13]/NET0131  & ~n281 ;
  assign n587 = \data_i[19]_pad  & n281 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = ~n266 & ~n516 ;
  assign n590 = ~n481 & ~n589 ;
  assign n591 = ~decrypt_i_pad & ~n590 ;
  assign n600 = \rd1_Key_o_reg[37]/NET0131  & ~n250 ;
  assign n601 = ~load_i_pad & ~\rd1_Key_o_reg[37]/NET0131  ;
  assign n602 = ~\key_i[21]_pad  & load_i_pad ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = n250 & n603 ;
  assign n605 = ~n600 & ~n604 ;
  assign n606 = n292 & ~n605 ;
  assign n592 = ~load_i_pad & ~\rd1_Key_o_reg[36]/NET0131  ;
  assign n593 = ~\key_i[29]_pad  & load_i_pad ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = n250 & n594 ;
  assign n596 = \rd1_Key_o_reg[38]/NET0131  & ~n281 ;
  assign n597 = \key_i[13]_pad  & n281 ;
  assign n598 = ~n596 & ~n597 ;
  assign n599 = n266 & ~n598 ;
  assign n607 = ~n595 & ~n599 ;
  assign n608 = ~n606 & n607 ;
  assign n609 = decrypt_i_pad & ~n608 ;
  assign n610 = ~n591 & ~n609 ;
  assign n611 = \rd1_Key_o_reg[48]/NET0131  & ~n250 ;
  assign n612 = ~n555 & ~n611 ;
  assign n613 = ~n266 & ~n612 ;
  assign n614 = n266 & ~n575 ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = ~decrypt_i_pad & ~n615 ;
  assign n624 = n292 & ~n561 ;
  assign n617 = \rd1_Key_o_reg[51]/NET0131  & ~n250 ;
  assign n618 = ~load_i_pad & ~\rd1_Key_o_reg[51]/NET0131  ;
  assign n619 = ~\key_i[39]_pad  & load_i_pad ;
  assign n620 = ~n618 & ~n619 ;
  assign n621 = n250 & n620 ;
  assign n622 = ~n617 & ~n621 ;
  assign n623 = n266 & ~n622 ;
  assign n625 = ~n567 & ~n623 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = decrypt_i_pad & ~n626 ;
  assign n628 = ~n616 & ~n627 ;
  assign n629 = \rd1_Key_o_reg[15]/NET0131  & ~n250 ;
  assign n630 = ~load_i_pad & ~\rd1_Key_o_reg[15]/NET0131  ;
  assign n631 = ~\key_i[34]_pad  & load_i_pad ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = n250 & n632 ;
  assign n634 = ~n629 & ~n633 ;
  assign n635 = n266 & ~n634 ;
  assign n636 = \rd1_Key_o_reg[16]/NET0131  & ~n250 ;
  assign n637 = ~load_i_pad & ~\rd1_Key_o_reg[16]/NET0131  ;
  assign n638 = ~\key_i[26]_pad  & load_i_pad ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = n250 & n639 ;
  assign n641 = ~n636 & ~n640 ;
  assign n642 = ~n266 & ~n641 ;
  assign n643 = ~n635 & ~n642 ;
  assign n644 = ~decrypt_i_pad & ~n643 ;
  assign n653 = \rd1_Key_o_reg[18]/NET0131  & ~n250 ;
  assign n654 = ~load_i_pad & ~\rd1_Key_o_reg[18]/NET0131  ;
  assign n655 = ~\key_i[10]_pad  & load_i_pad ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = n250 & n656 ;
  assign n658 = ~n653 & ~n657 ;
  assign n659 = n292 & ~n658 ;
  assign n645 = ~load_i_pad & ~\rd1_Key_o_reg[17]/NET0131  ;
  assign n646 = ~\key_i[18]_pad  & load_i_pad ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = n250 & n647 ;
  assign n649 = \rd1_Key_o_reg[19]/NET0131  & ~n281 ;
  assign n650 = \key_i[2]_pad  & n281 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = n266 & ~n651 ;
  assign n660 = ~n648 & ~n652 ;
  assign n661 = ~n659 & n660 ;
  assign n662 = decrypt_i_pad & ~n661 ;
  assign n663 = ~n644 & ~n662 ;
  assign n664 = \rd1_R_o_reg[0]/NET0131  & ~n281 ;
  assign n665 = \data_i[57]_pad  & n281 ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = \rd1_R_o_reg[16]/NET0131  & ~n281 ;
  assign n668 = \data_i[61]_pad  & n281 ;
  assign n669 = ~n667 & ~n668 ;
  assign n670 = \rd1_Key_o_reg[14]/NET0131  & ~n250 ;
  assign n671 = ~load_i_pad & ~\rd1_Key_o_reg[14]/NET0131  ;
  assign n672 = ~\key_i[42]_pad  & load_i_pad ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = n250 & n673 ;
  assign n675 = ~n670 & ~n674 ;
  assign n676 = ~n266 & ~n675 ;
  assign n677 = ~n444 & ~n676 ;
  assign n678 = ~decrypt_i_pad & ~n677 ;
  assign n681 = n292 & ~n641 ;
  assign n679 = \rd1_Key_o_reg[17]/NET0131  & ~n250 ;
  assign n680 = n266 & n679 ;
  assign n682 = ~n633 & ~n680 ;
  assign n683 = ~n681 & n682 ;
  assign n684 = decrypt_i_pad & ~n683 ;
  assign n685 = ~n678 & ~n684 ;
  assign n686 = \rd1_R_o_reg[7]/NET0131  & ~n281 ;
  assign n687 = \data_i[1]_pad  & n281 ;
  assign n688 = ~n686 & ~n687 ;
  assign n690 = n292 & ~n341 ;
  assign n689 = n266 & ~n454 ;
  assign n691 = ~n347 & ~n689 ;
  assign n692 = ~n690 & n691 ;
  assign n693 = decrypt_i_pad & ~n692 ;
  assign n694 = \rd1_Key_o_reg[54]/NET0131  & ~n281 ;
  assign n695 = \key_i[15]_pad  & n281 ;
  assign n696 = ~n694 & ~n695 ;
  assign n698 = n292 & ~n696 ;
  assign n697 = n250 & ~n696 ;
  assign n699 = \rd1_Key_o_reg[53]/NET0131  & ~n250 ;
  assign n700 = ~load_i_pad & ~\rd1_Key_o_reg[53]/NET0131  ;
  assign n701 = ~\key_i[23]_pad  & load_i_pad ;
  assign n702 = ~n700 & ~n701 ;
  assign n703 = n250 & n702 ;
  assign n704 = ~n699 & ~n703 ;
  assign n705 = n266 & ~n704 ;
  assign n706 = ~n697 & ~n705 ;
  assign n707 = ~n698 & n706 ;
  assign n708 = ~decrypt_i_pad & ~n707 ;
  assign n709 = ~n693 & ~n708 ;
  assign n717 = \rd1_Key_o_reg[45]/NET0131  & ~n250 ;
  assign n718 = ~load_i_pad & ~\rd1_Key_o_reg[45]/NET0131  ;
  assign n719 = ~\key_i[22]_pad  & load_i_pad ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = n250 & n720 ;
  assign n722 = ~n717 & ~n721 ;
  assign n723 = ~n266 & ~n722 ;
  assign n710 = \rd1_Key_o_reg[44]/NET0131  & ~n250 ;
  assign n711 = ~load_i_pad & ~\rd1_Key_o_reg[44]/NET0131  ;
  assign n712 = ~\key_i[30]_pad  & load_i_pad ;
  assign n713 = ~n711 & ~n712 ;
  assign n714 = n250 & n713 ;
  assign n715 = ~n710 & ~n714 ;
  assign n716 = n266 & ~n715 ;
  assign n724 = ~decrypt_i_pad & ~n716 ;
  assign n725 = ~n723 & n724 ;
  assign n726 = n250 & ~n579 ;
  assign n727 = n266 & ~n612 ;
  assign n728 = decrypt_i_pad & ~n727 ;
  assign n729 = ~n581 & n728 ;
  assign n730 = ~n726 & n729 ;
  assign n731 = ~n725 & ~n730 ;
  assign n732 = \rd1_Key_o_reg[36]/NET0131  & ~n250 ;
  assign n733 = ~n595 & ~n732 ;
  assign n734 = ~n266 & ~n733 ;
  assign n735 = ~n517 & ~n734 ;
  assign n736 = ~decrypt_i_pad & ~n735 ;
  assign n744 = n292 & ~n598 ;
  assign n737 = \rd1_Key_o_reg[39]/NET0131  & ~n250 ;
  assign n738 = ~load_i_pad & ~\rd1_Key_o_reg[39]/NET0131  ;
  assign n739 = ~\key_i[5]_pad  & load_i_pad ;
  assign n740 = ~n738 & ~n739 ;
  assign n741 = n250 & n740 ;
  assign n742 = ~n737 & ~n741 ;
  assign n743 = n266 & ~n742 ;
  assign n745 = ~n604 & ~n743 ;
  assign n746 = ~n744 & n745 ;
  assign n747 = decrypt_i_pad & ~n746 ;
  assign n748 = ~n736 & ~n747 ;
  assign n749 = \rd1_R_o_reg[30]/NET0131  & ~n281 ;
  assign n750 = \data_i[15]_pad  & n281 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = ~n266 & ~n715 ;
  assign n753 = \rd1_Key_o_reg[43]/NET0131  & ~n250 ;
  assign n754 = ~\key_i[38]_pad  & load_i_pad ;
  assign n755 = ~load_i_pad & ~\rd1_Key_o_reg[43]/NET0131  ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = n250 & n756 ;
  assign n758 = ~n753 & ~n757 ;
  assign n759 = n266 & ~n758 ;
  assign n760 = ~n752 & ~n759 ;
  assign n761 = ~decrypt_i_pad & ~n760 ;
  assign n762 = n292 & ~n579 ;
  assign n763 = ~n614 & ~n721 ;
  assign n764 = ~n762 & n763 ;
  assign n765 = decrypt_i_pad & ~n764 ;
  assign n766 = ~n761 & ~n765 ;
  assign n768 = n292 & ~n634 ;
  assign n767 = n266 & ~n641 ;
  assign n769 = ~n674 & ~n767 ;
  assign n770 = ~n768 & n769 ;
  assign n771 = decrypt_i_pad & ~n770 ;
  assign n773 = n250 & ~n443 ;
  assign n772 = n292 & ~n443 ;
  assign n774 = ~n499 & ~n772 ;
  assign n775 = ~n773 & n774 ;
  assign n776 = ~decrypt_i_pad & ~n775 ;
  assign n777 = ~n771 & ~n776 ;
  assign n778 = \rd1_R_o_reg[3]/NET0131  & ~n281 ;
  assign n779 = \data_i[33]_pad  & n281 ;
  assign n780 = ~n778 & ~n779 ;
  assign n781 = ~n777 & n780 ;
  assign n782 = n777 & ~n780 ;
  assign n783 = ~n781 & ~n782 ;
  assign n784 = n292 & ~n323 ;
  assign n785 = ~n329 & ~n494 ;
  assign n786 = ~n784 & n785 ;
  assign n787 = decrypt_i_pad & ~n786 ;
  assign n788 = n292 & ~n316 ;
  assign n789 = n266 & ~n310 ;
  assign n790 = ~n317 & ~n789 ;
  assign n791 = ~n788 & n790 ;
  assign n792 = ~decrypt_i_pad & ~n791 ;
  assign n793 = ~n787 & ~n792 ;
  assign n794 = \rd1_R_o_reg[2]/NET0131  & ~n281 ;
  assign n795 = \data_i[41]_pad  & n281 ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = ~n793 & n796 ;
  assign n798 = n793 & ~n796 ;
  assign n799 = ~n797 & ~n798 ;
  assign n800 = ~n783 & ~n799 ;
  assign n801 = n376 & ~n506 ;
  assign n802 = ~n376 & n506 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = n800 & ~n803 ;
  assign n806 = n292 & ~n382 ;
  assign n805 = n266 & ~n524 ;
  assign n807 = ~n388 & ~n805 ;
  assign n808 = ~n806 & n807 ;
  assign n809 = decrypt_i_pad & ~n808 ;
  assign n811 = n292 & ~n651 ;
  assign n810 = n250 & ~n651 ;
  assign n812 = n266 & ~n658 ;
  assign n813 = ~n810 & ~n812 ;
  assign n814 = ~n811 & n813 ;
  assign n815 = ~decrypt_i_pad & ~n814 ;
  assign n816 = ~n809 & ~n815 ;
  assign n817 = \rd1_R_o_reg[1]/NET0131  & ~n281 ;
  assign n818 = \data_i[49]_pad  & n281 ;
  assign n819 = ~n817 & ~n818 ;
  assign n820 = ~n816 & n819 ;
  assign n821 = n816 & ~n819 ;
  assign n822 = ~n820 & ~n821 ;
  assign n823 = n804 & ~n822 ;
  assign n824 = n783 & ~n803 ;
  assign n825 = n799 & n824 ;
  assign n826 = ~n822 & n825 ;
  assign n827 = ~n823 & ~n826 ;
  assign n828 = ~n799 & n803 ;
  assign n829 = n783 & n822 ;
  assign n830 = ~n799 & n829 ;
  assign n831 = ~n783 & n803 ;
  assign n832 = ~n830 & ~n831 ;
  assign n833 = ~n828 & ~n832 ;
  assign n834 = n827 & ~n833 ;
  assign n835 = ~n297 & n666 ;
  assign n836 = n297 & ~n666 ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = ~n834 & n837 ;
  assign n839 = n799 & n803 ;
  assign n840 = ~n837 & n839 ;
  assign n841 = n783 & ~n840 ;
  assign n845 = ~n799 & n837 ;
  assign n846 = n822 & ~n845 ;
  assign n847 = ~n841 & n846 ;
  assign n842 = ~n803 & n837 ;
  assign n843 = ~n822 & ~n842 ;
  assign n844 = n841 & n843 ;
  assign n848 = ~n403 & ~n805 ;
  assign n849 = ~n529 & n848 ;
  assign n850 = ~decrypt_i_pad & ~n849 ;
  assign n852 = ~n273 & n292 ;
  assign n851 = ~n261 & n266 ;
  assign n853 = ~n397 & ~n851 ;
  assign n854 = ~n852 & n853 ;
  assign n855 = decrypt_i_pad & ~n854 ;
  assign n856 = ~n850 & ~n855 ;
  assign n857 = \rd1_R_o_reg[31]/NET0131  & ~n281 ;
  assign n858 = \data_i[7]_pad  & n281 ;
  assign n859 = ~n857 & ~n858 ;
  assign n860 = ~n856 & n859 ;
  assign n861 = n856 & ~n859 ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = ~n844 & ~n862 ;
  assign n864 = ~n847 & n863 ;
  assign n865 = ~n838 & n864 ;
  assign n869 = ~n825 & n837 ;
  assign n870 = n803 & n829 ;
  assign n868 = ~n822 & n824 ;
  assign n871 = ~n800 & ~n868 ;
  assign n872 = ~n870 & n871 ;
  assign n873 = n869 & n872 ;
  assign n874 = n827 & n873 ;
  assign n875 = n803 & n822 ;
  assign n876 = n799 & ~n824 ;
  assign n877 = ~n875 & n876 ;
  assign n878 = ~n830 & ~n837 ;
  assign n879 = ~n877 & n878 ;
  assign n880 = ~n874 & ~n879 ;
  assign n866 = ~n822 & n828 ;
  assign n867 = ~n783 & n866 ;
  assign n881 = n862 & ~n867 ;
  assign n882 = ~n880 & n881 ;
  assign n883 = ~n865 & ~n882 ;
  assign n884 = ~\data_i[16]_pad  & n281 ;
  assign n885 = ~\rd1_L_o_reg[5]/NET0131  & ~n281 ;
  assign n886 = ~n884 & ~n885 ;
  assign n887 = n883 & ~n886 ;
  assign n888 = ~n883 & n886 ;
  assign n889 = ~n887 & ~n888 ;
  assign n916 = \rd1_Key_o_reg[42]/NET0131  & ~n281 ;
  assign n917 = \key_i[46]_pad  & n281 ;
  assign n918 = ~n916 & ~n917 ;
  assign n945 = n250 & ~n918 ;
  assign n944 = n292 & ~n918 ;
  assign n920 = \rd1_Key_o_reg[41]/NET0131  & ~n250 ;
  assign n921 = ~load_i_pad & ~\rd1_Key_o_reg[41]/NET0131  ;
  assign n922 = ~\key_i[54]_pad  & load_i_pad ;
  assign n923 = ~n921 & ~n922 ;
  assign n924 = n250 & n923 ;
  assign n925 = ~n920 & ~n924 ;
  assign n946 = n266 & ~n925 ;
  assign n947 = ~n944 & ~n946 ;
  assign n948 = ~n945 & n947 ;
  assign n949 = ~decrypt_i_pad & ~n948 ;
  assign n951 = n292 & ~n715 ;
  assign n950 = n266 & ~n722 ;
  assign n952 = ~n757 & ~n950 ;
  assign n953 = ~n951 & n952 ;
  assign n954 = decrypt_i_pad & ~n953 ;
  assign n955 = ~n949 & ~n954 ;
  assign n956 = n669 & ~n955 ;
  assign n957 = ~n669 & n955 ;
  assign n958 = ~n956 & ~n957 ;
  assign n896 = \rd1_R_o_reg[17]/NET0131  & ~n281 ;
  assign n897 = \data_i[53]_pad  & n281 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = ~n610 & n898 ;
  assign n900 = n610 & ~n898 ;
  assign n901 = ~n899 & ~n900 ;
  assign n903 = \rd1_R_o_reg[19]/NET0131  & ~n281 ;
  assign n904 = \data_i[37]_pad  & n281 ;
  assign n905 = ~n903 & ~n904 ;
  assign n906 = ~n628 & n905 ;
  assign n907 = n628 & ~n905 ;
  assign n908 = ~n906 & ~n907 ;
  assign n909 = ~n266 & ~n742 ;
  assign n910 = ~n599 & ~n909 ;
  assign n911 = ~decrypt_i_pad & ~n910 ;
  assign n926 = n292 & ~n925 ;
  assign n912 = ~load_i_pad & ~\rd1_Key_o_reg[40]/NET0131  ;
  assign n913 = ~\key_i[62]_pad  & load_i_pad ;
  assign n914 = ~n912 & ~n913 ;
  assign n915 = n250 & n914 ;
  assign n919 = n266 & ~n918 ;
  assign n927 = ~n915 & ~n919 ;
  assign n928 = ~n926 & n927 ;
  assign n929 = decrypt_i_pad & ~n928 ;
  assign n930 = ~n911 & ~n929 ;
  assign n931 = \rd1_R_o_reg[20]/NET0131  & ~n281 ;
  assign n932 = \data_i[29]_pad  & n281 ;
  assign n933 = ~n931 & ~n932 ;
  assign n934 = ~n930 & n933 ;
  assign n935 = n930 & ~n933 ;
  assign n936 = ~n934 & ~n935 ;
  assign n938 = n908 & n936 ;
  assign n960 = n901 & n938 ;
  assign n937 = ~n908 & ~n936 ;
  assign n939 = ~n937 & ~n938 ;
  assign n890 = \rd1_R_o_reg[18]/NET0131  & ~n281 ;
  assign n891 = \data_i[45]_pad  & n281 ;
  assign n892 = ~n890 & ~n891 ;
  assign n893 = ~n373 & n892 ;
  assign n894 = n373 & ~n892 ;
  assign n895 = ~n893 & ~n894 ;
  assign n961 = ~n895 & ~n901 ;
  assign n962 = n939 & n961 ;
  assign n963 = ~n960 & ~n962 ;
  assign n964 = n958 & ~n963 ;
  assign n902 = ~n895 & n901 ;
  assign n940 = n902 & ~n939 ;
  assign n941 = n895 & n939 ;
  assign n942 = ~n895 & n937 ;
  assign n943 = ~n941 & ~n942 ;
  assign n959 = ~n943 & ~n958 ;
  assign n965 = ~n940 & ~n959 ;
  assign n966 = ~n964 & n965 ;
  assign n967 = ~n266 & ~n704 ;
  assign n968 = \rd1_Key_o_reg[52]/NET0131  & ~n250 ;
  assign n969 = ~\key_i[31]_pad  & load_i_pad ;
  assign n970 = ~load_i_pad & ~\rd1_Key_o_reg[52]/NET0131  ;
  assign n971 = ~n969 & ~n970 ;
  assign n972 = n250 & n971 ;
  assign n973 = ~n968 & ~n972 ;
  assign n974 = n266 & ~n973 ;
  assign n975 = ~n967 & ~n974 ;
  assign n976 = ~decrypt_i_pad & ~n975 ;
  assign n977 = n292 & ~n348 ;
  assign n978 = ~n456 & ~n697 ;
  assign n979 = ~n977 & n978 ;
  assign n980 = decrypt_i_pad & ~n979 ;
  assign n981 = ~n976 & ~n980 ;
  assign n982 = \rd1_R_o_reg[15]/NET0131  & ~n281 ;
  assign n983 = \data_i[3]_pad  & n281 ;
  assign n984 = ~n982 & ~n983 ;
  assign n985 = ~n981 & n984 ;
  assign n986 = n981 & ~n984 ;
  assign n987 = ~n985 & ~n986 ;
  assign n988 = ~n966 & n987 ;
  assign n991 = ~n908 & n936 ;
  assign n992 = n901 & n991 ;
  assign n993 = ~n901 & ~n936 ;
  assign n994 = ~n908 & n993 ;
  assign n995 = ~n992 & ~n994 ;
  assign n996 = ~n941 & n995 ;
  assign n997 = n958 & ~n996 ;
  assign n989 = n902 & ~n936 ;
  assign n990 = ~n958 & n989 ;
  assign n998 = n938 & n961 ;
  assign n999 = ~n990 & ~n998 ;
  assign n1000 = ~n997 & n999 ;
  assign n1001 = ~n987 & ~n1000 ;
  assign n1004 = ~n895 & n938 ;
  assign n1005 = ~n994 & ~n1004 ;
  assign n1006 = n958 & ~n1005 ;
  assign n1007 = ~n961 & n1006 ;
  assign n1002 = n895 & n991 ;
  assign n1003 = n901 & n1002 ;
  assign n1008 = n895 & ~n901 ;
  assign n1009 = n908 & n1008 ;
  assign n1010 = n901 & n937 ;
  assign n1011 = ~n1009 & ~n1010 ;
  assign n1012 = ~n958 & ~n1011 ;
  assign n1013 = ~n1003 & ~n1012 ;
  assign n1014 = ~n1007 & n1013 ;
  assign n1015 = ~n1001 & n1014 ;
  assign n1016 = ~n988 & n1015 ;
  assign n1017 = ~\data_i[8]_pad  & n281 ;
  assign n1018 = ~\rd1_L_o_reg[6]/NET0131  & ~n281 ;
  assign n1019 = ~n1017 & ~n1018 ;
  assign n1020 = n1016 & ~n1019 ;
  assign n1021 = ~n1016 & n1019 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1023 = ~n266 & ~n273 ;
  assign n1024 = ~n399 & ~n1023 ;
  assign n1025 = ~decrypt_i_pad & ~n1024 ;
  assign n1027 = ~n280 & ~n536 ;
  assign n1028 = n292 & ~n1027 ;
  assign n1026 = n266 & ~n291 ;
  assign n1029 = ~n260 & ~n1026 ;
  assign n1030 = ~n1028 & n1029 ;
  assign n1031 = decrypt_i_pad & ~n1030 ;
  assign n1032 = ~n1025 & ~n1031 ;
  assign n1033 = ~n266 & ~n561 ;
  assign n1034 = n266 & ~n568 ;
  assign n1035 = ~n1033 & ~n1034 ;
  assign n1036 = ~decrypt_i_pad & ~n1035 ;
  assign n1037 = n292 & ~n973 ;
  assign n1038 = ~n621 & ~n705 ;
  assign n1039 = ~n1037 & n1038 ;
  assign n1040 = decrypt_i_pad & ~n1039 ;
  assign n1041 = ~n1036 & ~n1040 ;
  assign n1042 = ~n266 & ~n658 ;
  assign n1043 = ~n680 & ~n1042 ;
  assign n1044 = ~decrypt_i_pad & ~n1043 ;
  assign n1045 = n292 & ~n389 ;
  assign n1046 = ~n526 & ~n810 ;
  assign n1047 = ~n1045 & n1046 ;
  assign n1048 = decrypt_i_pad & ~n1047 ;
  assign n1049 = ~n1044 & ~n1048 ;
  assign n1050 = n266 & ~n330 ;
  assign n1051 = ~n309 & ~n1050 ;
  assign n1052 = ~n788 & n1051 ;
  assign n1053 = decrypt_i_pad & ~n1052 ;
  assign n1055 = n292 & ~n303 ;
  assign n1054 = n250 & ~n303 ;
  assign n1056 = n266 & ~n546 ;
  assign n1057 = ~n1054 & ~n1056 ;
  assign n1058 = ~n1055 & n1057 ;
  assign n1059 = ~decrypt_i_pad & ~n1058 ;
  assign n1060 = ~n1053 & ~n1059 ;
  assign n1061 = \rd1_R_o_reg[28]/NET0131  & ~n281 ;
  assign n1062 = \data_i[31]_pad  & n281 ;
  assign n1063 = ~n1061 & ~n1062 ;
  assign n1064 = ~n266 & ~n973 ;
  assign n1065 = ~n623 & ~n1064 ;
  assign n1066 = ~decrypt_i_pad & ~n1065 ;
  assign n1067 = ~n349 & ~n703 ;
  assign n1068 = ~n698 & n1067 ;
  assign n1069 = decrypt_i_pad & ~n1068 ;
  assign n1070 = ~n1066 & ~n1069 ;
  assign n1071 = \rd1_Key_o_reg[40]/NET0131  & ~n250 ;
  assign n1072 = ~n915 & ~n1071 ;
  assign n1073 = ~n266 & ~n1072 ;
  assign n1074 = ~n743 & ~n1073 ;
  assign n1075 = ~decrypt_i_pad & ~n1074 ;
  assign n1076 = ~n759 & ~n924 ;
  assign n1077 = ~n944 & n1076 ;
  assign n1078 = decrypt_i_pad & ~n1077 ;
  assign n1079 = ~n1075 & ~n1078 ;
  assign n1080 = \rd1_R_o_reg[26]/NET0131  & ~n281 ;
  assign n1081 = \data_i[47]_pad  & n281 ;
  assign n1082 = ~n1080 & ~n1081 ;
  assign n1099 = n669 & ~n685 ;
  assign n1100 = ~n669 & n685 ;
  assign n1101 = ~n1099 & ~n1100 ;
  assign n1102 = n984 & ~n1060 ;
  assign n1103 = ~n984 & n1060 ;
  assign n1104 = ~n1102 & ~n1103 ;
  assign n1105 = ~n1101 & n1104 ;
  assign n1106 = n1101 & ~n1104 ;
  assign n1107 = n588 & ~n1049 ;
  assign n1108 = ~n588 & n1049 ;
  assign n1109 = ~n1107 & ~n1108 ;
  assign n1110 = n1106 & ~n1109 ;
  assign n1111 = ~n1105 & ~n1110 ;
  assign n1112 = n266 & ~n402 ;
  assign n1113 = ~n266 & ~n398 ;
  assign n1114 = ~n1112 & ~n1113 ;
  assign n1115 = ~decrypt_i_pad & ~n1114 ;
  assign n1116 = ~n261 & n292 ;
  assign n1117 = ~n272 & ~n537 ;
  assign n1118 = ~n1116 & n1117 ;
  assign n1119 = decrypt_i_pad & ~n1118 ;
  assign n1120 = ~n1115 & ~n1119 ;
  assign n1121 = \rd1_R_o_reg[14]/NET0131  & ~n281 ;
  assign n1122 = \data_i[11]_pad  & n281 ;
  assign n1123 = ~n1121 & ~n1122 ;
  assign n1124 = ~n1120 & n1123 ;
  assign n1125 = n1120 & ~n1123 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = ~n1111 & ~n1126 ;
  assign n1130 = n1104 & ~n1109 ;
  assign n1131 = n1126 & n1130 ;
  assign n1083 = n250 & ~n422 ;
  assign n1084 = ~n324 & ~n423 ;
  assign n1085 = ~n1083 & n1084 ;
  assign n1086 = ~decrypt_i_pad & ~n1085 ;
  assign n1088 = n292 & ~n433 ;
  assign n1087 = n266 & ~n501 ;
  assign n1089 = ~n495 & ~n1087 ;
  assign n1090 = ~n1088 & n1089 ;
  assign n1091 = decrypt_i_pad & ~n1090 ;
  assign n1092 = ~n1086 & ~n1091 ;
  assign n1093 = \rd1_R_o_reg[12]/NET0131  & ~n281 ;
  assign n1094 = \data_i[27]_pad  & n281 ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = ~n1092 & n1095 ;
  assign n1097 = n1092 & ~n1095 ;
  assign n1098 = ~n1096 & ~n1097 ;
  assign n1128 = ~n1101 & ~n1104 ;
  assign n1129 = n1109 & n1128 ;
  assign n1132 = ~n1098 & ~n1129 ;
  assign n1133 = ~n1131 & n1132 ;
  assign n1134 = ~n1127 & n1133 ;
  assign n1138 = n1104 & n1109 ;
  assign n1139 = ~n1104 & n1126 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1141 = n1101 & ~n1140 ;
  assign n1135 = n1104 & ~n1126 ;
  assign n1136 = n1101 & n1135 ;
  assign n1137 = n1098 & ~n1136 ;
  assign n1142 = ~n1109 & ~n1126 ;
  assign n1143 = n1128 & n1142 ;
  assign n1144 = n1137 & ~n1143 ;
  assign n1145 = ~n1141 & n1144 ;
  assign n1146 = ~n1134 & ~n1145 ;
  assign n1147 = n1105 & n1126 ;
  assign n1148 = ~n1109 & n1147 ;
  assign n1149 = ~n1126 & n1138 ;
  assign n1150 = n1101 & n1149 ;
  assign n1151 = ~n1148 & ~n1150 ;
  assign n1152 = ~n1146 & n1151 ;
  assign n1153 = \rd1_R_o_reg[11]/NET0131  & ~n281 ;
  assign n1154 = \data_i[35]_pad  & n281 ;
  assign n1155 = ~n1153 & ~n1154 ;
  assign n1156 = ~n551 & n1155 ;
  assign n1157 = n551 & ~n1155 ;
  assign n1158 = ~n1156 & ~n1157 ;
  assign n1159 = ~n1152 & ~n1158 ;
  assign n1160 = n1101 & n1126 ;
  assign n1161 = ~n1101 & ~n1109 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = ~n1130 & ~n1162 ;
  assign n1164 = n1101 & n1142 ;
  assign n1165 = n1104 & n1164 ;
  assign n1166 = ~n1163 & ~n1165 ;
  assign n1167 = n1158 & ~n1166 ;
  assign n1168 = ~n1101 & n1138 ;
  assign n1169 = ~n1126 & n1168 ;
  assign n1170 = ~n1167 & ~n1169 ;
  assign n1171 = ~n1098 & ~n1170 ;
  assign n1172 = n1098 & n1109 ;
  assign n1173 = ~n1135 & n1172 ;
  assign n1174 = ~n1101 & n1173 ;
  assign n1175 = ~n1101 & ~n1135 ;
  assign n1176 = n1140 & ~n1175 ;
  assign n1177 = n1137 & n1176 ;
  assign n1178 = ~n1174 & ~n1177 ;
  assign n1179 = n1158 & ~n1178 ;
  assign n1180 = n1101 & n1138 ;
  assign n1181 = n1098 & ~n1126 ;
  assign n1182 = n1180 & n1181 ;
  assign n1183 = ~n1109 & n1158 ;
  assign n1184 = ~n1172 & ~n1183 ;
  assign n1185 = n1126 & n1128 ;
  assign n1186 = ~n1184 & n1185 ;
  assign n1187 = ~n1182 & ~n1186 ;
  assign n1188 = ~n1179 & n1187 ;
  assign n1189 = ~n1171 & n1188 ;
  assign n1190 = ~n1159 & n1189 ;
  assign n1191 = ~\data_i[44]_pad  & n281 ;
  assign n1192 = ~\rd1_L_o_reg[18]/NET0131  & ~n281 ;
  assign n1193 = ~n1191 & ~n1192 ;
  assign n1194 = n1190 & ~n1193 ;
  assign n1195 = ~n1190 & n1193 ;
  assign n1196 = ~n1194 & ~n1195 ;
  assign n1197 = \rd1_R_o_reg[8]/NET0131  & ~n281 ;
  assign n1198 = \data_i[59]_pad  & n281 ;
  assign n1199 = ~n1197 & ~n1198 ;
  assign n1200 = ~n266 & ~n501 ;
  assign n1201 = n266 & ~n433 ;
  assign n1202 = ~n1200 & ~n1201 ;
  assign n1203 = ~decrypt_i_pad & ~n1202 ;
  assign n1204 = n250 & ~n439 ;
  assign n1205 = n266 & ~n675 ;
  assign n1206 = ~n772 & ~n1205 ;
  assign n1207 = ~n1204 & n1206 ;
  assign n1208 = decrypt_i_pad & ~n1207 ;
  assign n1209 = ~n1203 & ~n1208 ;
  assign n1210 = ~n266 & ~n634 ;
  assign n1211 = ~n1205 & ~n1210 ;
  assign n1212 = ~decrypt_i_pad & ~n1211 ;
  assign n1213 = ~n648 & ~n679 ;
  assign n1214 = n292 & ~n1213 ;
  assign n1215 = ~n640 & ~n812 ;
  assign n1216 = ~n1214 & n1215 ;
  assign n1217 = decrypt_i_pad & ~n1216 ;
  assign n1218 = ~n1212 & ~n1217 ;
  assign n1219 = ~n266 & ~n323 ;
  assign n1220 = ~n1050 & ~n1219 ;
  assign n1221 = ~decrypt_i_pad & ~n1220 ;
  assign n1222 = ~n493 & ~n1201 ;
  assign n1223 = ~n1083 & n1222 ;
  assign n1224 = decrypt_i_pad & ~n1223 ;
  assign n1225 = ~n1221 & ~n1224 ;
  assign n1264 = \rd1_R_o_reg[23]/NET0131  & ~n281 ;
  assign n1265 = \data_i[5]_pad  & n281 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = n731 & n1266 ;
  assign n1268 = ~n731 & ~n1266 ;
  assign n1269 = ~n1267 & ~n1268 ;
  assign n1259 = n1063 & ~n1070 ;
  assign n1260 = ~n1063 & n1070 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1240 = ~n1079 & n1082 ;
  assign n1241 = n1079 & ~n1082 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = ~n266 & ~n348 ;
  assign n1244 = n266 & ~n696 ;
  assign n1245 = ~n1243 & ~n1244 ;
  assign n1246 = ~decrypt_i_pad & ~n1245 ;
  assign n1247 = n292 & ~n454 ;
  assign n1248 = ~n340 & ~n472 ;
  assign n1249 = ~n1247 & n1248 ;
  assign n1250 = decrypt_i_pad & ~n1249 ;
  assign n1251 = ~n1246 & ~n1250 ;
  assign n1252 = \rd1_R_o_reg[27]/NET0131  & ~n281 ;
  assign n1253 = \data_i[39]_pad  & n281 ;
  assign n1254 = ~n1252 & ~n1253 ;
  assign n1255 = ~n1251 & n1254 ;
  assign n1256 = n1251 & ~n1254 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1270 = n1242 & n1257 ;
  assign n1271 = ~n1261 & n1270 ;
  assign n1226 = ~n266 & ~n568 ;
  assign n1227 = ~n727 & ~n1226 ;
  assign n1228 = ~decrypt_i_pad & ~n1227 ;
  assign n1229 = n292 & ~n622 ;
  assign n1230 = ~n560 & ~n974 ;
  assign n1231 = ~n1229 & n1230 ;
  assign n1232 = decrypt_i_pad & ~n1231 ;
  assign n1233 = ~n1228 & ~n1232 ;
  assign n1234 = \rd1_R_o_reg[25]/NET0131  & ~n281 ;
  assign n1235 = \data_i[55]_pad  & n281 ;
  assign n1236 = ~n1234 & ~n1235 ;
  assign n1237 = ~n1233 & n1236 ;
  assign n1238 = n1233 & ~n1236 ;
  assign n1239 = ~n1237 & ~n1238 ;
  assign n1272 = ~n1239 & ~n1242 ;
  assign n1273 = ~n1257 & n1272 ;
  assign n1274 = ~n1271 & ~n1273 ;
  assign n1275 = n1239 & n1242 ;
  assign n1277 = n1261 & ~n1275 ;
  assign n1276 = ~n1261 & n1275 ;
  assign n1278 = ~n1257 & ~n1276 ;
  assign n1279 = ~n1277 & n1278 ;
  assign n1280 = n1274 & ~n1279 ;
  assign n1281 = n1269 & ~n1280 ;
  assign n1282 = n1261 & n1270 ;
  assign n1283 = ~n1239 & n1282 ;
  assign n1284 = ~n1281 & ~n1283 ;
  assign n1285 = n266 & ~n484 ;
  assign n1286 = ~n266 & ~n480 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1288 = ~decrypt_i_pad & ~n1287 ;
  assign n1290 = n292 & ~n733 ;
  assign n1289 = n266 & ~n605 ;
  assign n1291 = ~n515 & ~n1289 ;
  assign n1292 = ~n1290 & n1291 ;
  assign n1293 = decrypt_i_pad & ~n1292 ;
  assign n1294 = ~n1288 & ~n1293 ;
  assign n1295 = \rd1_R_o_reg[24]/NET0131  & ~n281 ;
  assign n1296 = \data_i[63]_pad  & n281 ;
  assign n1297 = ~n1295 & ~n1296 ;
  assign n1298 = ~n1294 & n1297 ;
  assign n1299 = n1294 & ~n1297 ;
  assign n1300 = ~n1298 & ~n1299 ;
  assign n1301 = ~n1284 & ~n1300 ;
  assign n1310 = ~n1275 & ~n1300 ;
  assign n1302 = n1242 & ~n1261 ;
  assign n1309 = ~n1242 & ~n1257 ;
  assign n1311 = ~n1302 & ~n1309 ;
  assign n1312 = n1310 & n1311 ;
  assign n1303 = n1239 & ~n1257 ;
  assign n1304 = n1302 & n1303 ;
  assign n1305 = ~n1257 & n1300 ;
  assign n1306 = ~n1242 & n1261 ;
  assign n1307 = ~n1302 & ~n1306 ;
  assign n1308 = n1305 & ~n1307 ;
  assign n1313 = ~n1304 & ~n1308 ;
  assign n1314 = ~n1312 & n1313 ;
  assign n1315 = ~n1269 & ~n1314 ;
  assign n1322 = ~n1239 & n1257 ;
  assign n1323 = n1302 & n1322 ;
  assign n1317 = ~n1239 & n1261 ;
  assign n1324 = ~n1317 & ~n1322 ;
  assign n1325 = ~n1302 & ~n1303 ;
  assign n1326 = n1324 & n1325 ;
  assign n1327 = ~n1323 & ~n1326 ;
  assign n1328 = n1300 & ~n1327 ;
  assign n1258 = ~n1242 & n1257 ;
  assign n1262 = n1258 & n1261 ;
  assign n1263 = n1239 & n1262 ;
  assign n1316 = n1262 & n1300 ;
  assign n1318 = n1305 & n1317 ;
  assign n1319 = n1242 & n1318 ;
  assign n1320 = ~n1316 & ~n1319 ;
  assign n1321 = n1269 & ~n1320 ;
  assign n1329 = ~n1263 & ~n1321 ;
  assign n1330 = ~n1328 & n1329 ;
  assign n1331 = ~n1315 & n1330 ;
  assign n1332 = ~n1301 & n1331 ;
  assign n1333 = ~\data_i[14]_pad  & n281 ;
  assign n1334 = ~\rd1_L_o_reg[30]/NET0131  & ~n281 ;
  assign n1335 = ~n1333 & ~n1334 ;
  assign n1336 = n1332 & ~n1335 ;
  assign n1337 = ~n1332 & n1335 ;
  assign n1338 = ~n1336 & ~n1337 ;
  assign n1339 = n266 & ~n1072 ;
  assign n1340 = ~n266 & ~n925 ;
  assign n1341 = ~n1339 & ~n1340 ;
  assign n1342 = ~decrypt_i_pad & ~n1341 ;
  assign n1343 = n292 & ~n758 ;
  assign n1344 = ~n716 & ~n945 ;
  assign n1345 = ~n1343 & n1344 ;
  assign n1346 = decrypt_i_pad & ~n1345 ;
  assign n1347 = ~n1342 & ~n1346 ;
  assign n1348 = ~n266 & ~n1027 ;
  assign n1349 = ~n851 & ~n1348 ;
  assign n1350 = ~decrypt_i_pad & ~n1349 ;
  assign n1351 = ~n284 & n292 ;
  assign n1352 = ~n290 & ~n1056 ;
  assign n1353 = ~n1351 & n1352 ;
  assign n1354 = decrypt_i_pad & ~n1353 ;
  assign n1355 = ~n1350 & ~n1354 ;
  assign n1368 = n908 & ~n936 ;
  assign n1369 = n895 & n1368 ;
  assign n1383 = ~n992 & ~n1369 ;
  assign n1384 = ~n958 & ~n1383 ;
  assign n1385 = n937 & n961 ;
  assign n1386 = ~n1384 & ~n1385 ;
  assign n1387 = n901 & ~n908 ;
  assign n1388 = n958 & ~n1387 ;
  assign n1389 = ~n938 & ~n993 ;
  assign n1390 = n1388 & n1389 ;
  assign n1391 = n901 & n1004 ;
  assign n1392 = ~n1390 & ~n1391 ;
  assign n1393 = n1386 & n1392 ;
  assign n1394 = ~n987 & ~n1393 ;
  assign n1356 = ~n901 & n938 ;
  assign n1357 = n895 & n1356 ;
  assign n1358 = n908 & n993 ;
  assign n1359 = ~n992 & ~n1358 ;
  assign n1360 = ~n895 & n1359 ;
  assign n1361 = ~n941 & n958 ;
  assign n1362 = ~n1360 & n1361 ;
  assign n1363 = ~n1357 & ~n1362 ;
  assign n1364 = n987 & ~n1363 ;
  assign n1379 = n902 & n937 ;
  assign n1380 = ~n1004 & ~n1379 ;
  assign n1381 = ~n1003 & n1380 ;
  assign n1382 = ~n958 & ~n1381 ;
  assign n1365 = ~n901 & n936 ;
  assign n1366 = n895 & n958 ;
  assign n1367 = n1365 & n1366 ;
  assign n1370 = n901 & n1369 ;
  assign n1371 = ~n1367 & ~n1370 ;
  assign n1372 = n908 & ~n1371 ;
  assign n1373 = n937 & ~n958 ;
  assign n1374 = n1008 & n1373 ;
  assign n1375 = ~n961 & ~n1368 ;
  assign n1376 = ~n958 & n987 ;
  assign n1377 = ~n993 & n1376 ;
  assign n1378 = ~n1375 & n1377 ;
  assign n1395 = ~n1374 & ~n1378 ;
  assign n1396 = ~n1372 & n1395 ;
  assign n1397 = ~n1382 & n1396 ;
  assign n1398 = ~n1364 & n1397 ;
  assign n1399 = ~n1394 & n1398 ;
  assign n1400 = ~\data_i[12]_pad  & n281 ;
  assign n1401 = ~\rd1_L_o_reg[22]/NET0131  & ~n281 ;
  assign n1402 = ~n1400 & ~n1401 ;
  assign n1403 = n1399 & ~n1402 ;
  assign n1404 = ~n1399 & n1402 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = ~n266 & ~n546 ;
  assign n1407 = ~n285 & ~n1406 ;
  assign n1408 = ~decrypt_i_pad & ~n1407 ;
  assign n1409 = n292 & ~n310 ;
  assign n1410 = ~n413 & ~n1054 ;
  assign n1411 = ~n1409 & n1410 ;
  assign n1412 = decrypt_i_pad & ~n1411 ;
  assign n1413 = ~n1408 & ~n1412 ;
  assign n1414 = n780 & ~n1413 ;
  assign n1415 = ~n780 & n1413 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = n376 & ~n411 ;
  assign n1418 = ~n376 & n411 ;
  assign n1419 = ~n1417 & ~n1418 ;
  assign n1420 = n1199 & ~n1209 ;
  assign n1421 = ~n1199 & n1209 ;
  assign n1422 = ~n1420 & ~n1421 ;
  assign n1427 = \rd1_R_o_reg[6]/NET0131  & ~n281 ;
  assign n1428 = \data_i[9]_pad  & n281 ;
  assign n1429 = ~n1427 & ~n1428 ;
  assign n1430 = ~n663 & n1429 ;
  assign n1431 = n663 & ~n1429 ;
  assign n1432 = ~n1430 & ~n1431 ;
  assign n1458 = ~n1422 & ~n1432 ;
  assign n1423 = ~n427 & n688 ;
  assign n1424 = n427 & ~n688 ;
  assign n1425 = ~n1423 & ~n1424 ;
  assign n1426 = ~n1422 & ~n1425 ;
  assign n1435 = \rd1_R_o_reg[5]/NET0131  & ~n281 ;
  assign n1436 = \data_i[17]_pad  & n281 ;
  assign n1437 = ~n1435 & ~n1436 ;
  assign n1438 = ~n1355 & n1437 ;
  assign n1439 = n1355 & ~n1437 ;
  assign n1440 = ~n1438 & ~n1439 ;
  assign n1468 = n1425 & ~n1432 ;
  assign n1469 = n1440 & n1468 ;
  assign n1470 = ~n1426 & ~n1469 ;
  assign n1471 = ~n1458 & ~n1470 ;
  assign n1472 = n1422 & n1425 ;
  assign n1473 = ~n1426 & ~n1472 ;
  assign n1452 = n1422 & n1432 ;
  assign n1474 = ~n1440 & ~n1452 ;
  assign n1475 = n1473 & n1474 ;
  assign n1476 = ~n1471 & ~n1475 ;
  assign n1477 = n1419 & ~n1476 ;
  assign n1453 = ~n1425 & n1440 ;
  assign n1466 = ~n1422 & n1453 ;
  assign n1467 = n1432 & n1466 ;
  assign n1441 = ~n1422 & n1432 ;
  assign n1448 = n1422 & ~n1432 ;
  assign n1478 = ~n1441 & ~n1448 ;
  assign n1479 = ~n1419 & ~n1453 ;
  assign n1480 = n1478 & n1479 ;
  assign n1481 = ~n1467 & ~n1480 ;
  assign n1482 = ~n1477 & n1481 ;
  assign n1483 = n1416 & ~n1482 ;
  assign n1433 = n1426 & ~n1432 ;
  assign n1434 = n1419 & n1433 ;
  assign n1443 = n1426 & n1432 ;
  assign n1442 = n1425 & ~n1441 ;
  assign n1444 = n1440 & ~n1442 ;
  assign n1445 = ~n1443 & n1444 ;
  assign n1446 = ~n1434 & ~n1445 ;
  assign n1447 = ~n1416 & ~n1446 ;
  assign n1460 = ~n1416 & ~n1419 ;
  assign n1462 = ~n1440 & n1443 ;
  assign n1449 = ~n1425 & n1448 ;
  assign n1454 = n1425 & ~n1440 ;
  assign n1461 = n1422 & n1454 ;
  assign n1463 = ~n1449 & ~n1461 ;
  assign n1464 = ~n1462 & n1463 ;
  assign n1465 = n1460 & ~n1464 ;
  assign n1455 = ~n1453 & ~n1454 ;
  assign n1450 = ~n1419 & n1440 ;
  assign n1456 = ~n1450 & n1452 ;
  assign n1457 = ~n1455 & n1456 ;
  assign n1451 = n1449 & n1450 ;
  assign n1459 = n1454 & n1458 ;
  assign n1484 = ~n1451 & ~n1459 ;
  assign n1485 = ~n1457 & n1484 ;
  assign n1486 = ~n1465 & n1485 ;
  assign n1487 = ~n1447 & n1486 ;
  assign n1488 = ~n1483 & n1487 ;
  assign n1489 = ~\data_i[42]_pad  & n281 ;
  assign n1490 = ~\rd1_L_o_reg[10]/NET0131  & ~n281 ;
  assign n1491 = ~n1489 & ~n1490 ;
  assign n1492 = n1488 & ~n1491 ;
  assign n1493 = ~n1488 & n1491 ;
  assign n1494 = ~n1492 & ~n1493 ;
  assign n1496 = n1425 & n1452 ;
  assign n1505 = n1450 & ~n1458 ;
  assign n1506 = ~n1496 & n1505 ;
  assign n1513 = n1419 & ~n1440 ;
  assign n1516 = ~n1448 & ~n1450 ;
  assign n1517 = ~n1513 & ~n1516 ;
  assign n1518 = ~n1506 & n1517 ;
  assign n1511 = n1432 & n1473 ;
  assign n1512 = ~n1450 & n1511 ;
  assign n1514 = ~n1422 & n1425 ;
  assign n1515 = n1513 & n1514 ;
  assign n1519 = ~n1512 & ~n1515 ;
  assign n1520 = ~n1518 & n1519 ;
  assign n1521 = n1416 & ~n1520 ;
  assign n1497 = ~n1422 & n1469 ;
  assign n1498 = n1419 & ~n1496 ;
  assign n1499 = ~n1497 & n1498 ;
  assign n1500 = ~n1419 & ~n1443 ;
  assign n1501 = ~n1459 & n1500 ;
  assign n1502 = ~n1499 & ~n1501 ;
  assign n1503 = ~n1419 & ~n1432 ;
  assign n1504 = n1461 & ~n1503 ;
  assign n1507 = ~n1467 & ~n1504 ;
  assign n1508 = ~n1506 & n1507 ;
  assign n1509 = ~n1502 & n1508 ;
  assign n1510 = ~n1416 & ~n1509 ;
  assign n1495 = ~n1419 & n1467 ;
  assign n1522 = ~n1433 & ~n1511 ;
  assign n1523 = n1513 & ~n1522 ;
  assign n1524 = ~n1495 & ~n1523 ;
  assign n1525 = ~n1510 & n1524 ;
  assign n1526 = ~n1521 & n1525 ;
  assign n1527 = ~\data_i[54]_pad  & n281 ;
  assign n1528 = ~\rd1_L_o_reg[25]/NET0131  & ~n281 ;
  assign n1529 = ~n1527 & ~n1528 ;
  assign n1530 = n1526 & ~n1529 ;
  assign n1531 = ~n1526 & n1529 ;
  assign n1532 = ~n1530 & ~n1531 ;
  assign n1577 = ~n1041 & n1254 ;
  assign n1578 = n1041 & ~n1254 ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1566 = ~n709 & n1063 ;
  assign n1567 = n709 & ~n1063 ;
  assign n1568 = ~n1566 & ~n1567 ;
  assign n1536 = n751 & ~n766 ;
  assign n1537 = ~n751 & n766 ;
  assign n1538 = ~n1536 & ~n1537 ;
  assign n1539 = n250 & ~n598 ;
  assign n1540 = ~n744 & ~n1289 ;
  assign n1541 = ~n1539 & n1540 ;
  assign n1542 = ~decrypt_i_pad & ~n1541 ;
  assign n1543 = n292 & ~n1072 ;
  assign n1544 = ~n741 & ~n946 ;
  assign n1545 = ~n1543 & n1544 ;
  assign n1546 = decrypt_i_pad & ~n1545 ;
  assign n1547 = ~n1542 & ~n1546 ;
  assign n1548 = n859 & ~n1547 ;
  assign n1549 = ~n859 & n1547 ;
  assign n1550 = ~n1548 & ~n1549 ;
  assign n1552 = n666 & ~n1347 ;
  assign n1553 = ~n666 & n1347 ;
  assign n1554 = ~n1552 & ~n1553 ;
  assign n1561 = n1550 & n1554 ;
  assign n1581 = ~n1538 & n1561 ;
  assign n1582 = ~n1550 & n1554 ;
  assign n1583 = n1538 & n1582 ;
  assign n1584 = ~n1581 & ~n1583 ;
  assign n1533 = ~n489 & n492 ;
  assign n1534 = n489 & ~n492 ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1559 = n1550 & ~n1554 ;
  assign n1586 = ~n1535 & ~n1559 ;
  assign n1560 = n1535 & n1559 ;
  assign n1585 = n1535 & n1582 ;
  assign n1587 = ~n1560 & ~n1585 ;
  assign n1588 = ~n1586 & n1587 ;
  assign n1589 = n1584 & ~n1588 ;
  assign n1590 = n1568 & ~n1589 ;
  assign n1591 = ~n1550 & ~n1554 ;
  assign n1592 = n1535 & ~n1538 ;
  assign n1593 = n1591 & n1592 ;
  assign n1594 = ~n1590 & ~n1593 ;
  assign n1595 = n1579 & ~n1594 ;
  assign n1557 = ~n1535 & ~n1538 ;
  assign n1558 = ~n1550 & n1557 ;
  assign n1562 = ~n1535 & n1561 ;
  assign n1563 = ~n1560 & ~n1562 ;
  assign n1564 = n1538 & ~n1563 ;
  assign n1565 = ~n1558 & ~n1564 ;
  assign n1569 = ~n1565 & n1568 ;
  assign n1551 = n1538 & ~n1550 ;
  assign n1555 = n1551 & ~n1554 ;
  assign n1556 = ~n1535 & n1555 ;
  assign n1571 = ~n1535 & n1559 ;
  assign n1570 = n1535 & n1561 ;
  assign n1572 = ~n1551 & ~n1570 ;
  assign n1573 = ~n1571 & n1572 ;
  assign n1574 = ~n1568 & ~n1573 ;
  assign n1575 = ~n1556 & ~n1574 ;
  assign n1576 = ~n1569 & n1575 ;
  assign n1580 = ~n1576 & ~n1579 ;
  assign n1596 = n1568 & n1593 ;
  assign n1599 = ~n1538 & ~n1561 ;
  assign n1597 = n1535 & ~n1550 ;
  assign n1598 = ~n1568 & ~n1597 ;
  assign n1600 = n1579 & ~n1591 ;
  assign n1601 = n1598 & n1600 ;
  assign n1602 = n1599 & n1601 ;
  assign n1605 = ~n1596 & ~n1602 ;
  assign n1603 = n1535 & ~n1584 ;
  assign n1604 = n1556 & ~n1568 ;
  assign n1606 = ~n1603 & ~n1604 ;
  assign n1607 = n1605 & n1606 ;
  assign n1608 = ~n1580 & n1607 ;
  assign n1609 = ~n1595 & n1608 ;
  assign n1610 = ~\data_i[50]_pad  & n281 ;
  assign n1611 = ~\rd1_L_o_reg[9]/NET0131  & ~n281 ;
  assign n1612 = ~n1610 & ~n1611 ;
  assign n1613 = n1609 & ~n1612 ;
  assign n1614 = ~n1609 & n1612 ;
  assign n1615 = ~n1613 & ~n1614 ;
  assign n1619 = n1155 & ~n1218 ;
  assign n1620 = ~n1155 & n1218 ;
  assign n1621 = ~n1619 & ~n1620 ;
  assign n1630 = \rd1_R_o_reg[9]/NET0131  & ~n281 ;
  assign n1631 = \data_i[51]_pad  & n281 ;
  assign n1632 = ~n1630 & ~n1631 ;
  assign n1633 = ~n452 & n1632 ;
  assign n1634 = n452 & ~n1632 ;
  assign n1635 = ~n1633 & ~n1634 ;
  assign n1616 = ~n1032 & n1095 ;
  assign n1617 = n1032 & ~n1095 ;
  assign n1618 = ~n1616 & ~n1617 ;
  assign n1625 = n300 & ~n335 ;
  assign n1626 = ~n300 & n335 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1641 = n1618 & n1627 ;
  assign n1642 = ~n1635 & n1641 ;
  assign n1643 = n1621 & n1642 ;
  assign n1622 = ~n1618 & n1621 ;
  assign n1623 = n1618 & ~n1621 ;
  assign n1624 = ~n1622 & ~n1623 ;
  assign n1628 = n1624 & n1627 ;
  assign n1629 = n1621 & ~n1627 ;
  assign n1636 = ~n1629 & n1635 ;
  assign n1637 = ~n1628 & n1636 ;
  assign n1638 = ~n534 & n1199 ;
  assign n1639 = n534 & ~n1199 ;
  assign n1640 = ~n1638 & ~n1639 ;
  assign n1644 = ~n1637 & ~n1640 ;
  assign n1645 = ~n1643 & n1644 ;
  assign n1648 = ~n1618 & ~n1627 ;
  assign n1649 = ~n1635 & ~n1648 ;
  assign n1650 = ~n1641 & n1649 ;
  assign n1646 = n1621 & ~n1635 ;
  assign n1647 = n1628 & ~n1646 ;
  assign n1651 = n1640 & ~n1647 ;
  assign n1652 = ~n1650 & n1651 ;
  assign n1653 = ~n1645 & ~n1652 ;
  assign n1654 = n1623 & ~n1627 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = n688 & ~n1225 ;
  assign n1657 = ~n688 & n1225 ;
  assign n1658 = ~n1656 & ~n1657 ;
  assign n1659 = ~n1655 & ~n1658 ;
  assign n1662 = ~n1618 & ~n1621 ;
  assign n1663 = ~n1627 & n1662 ;
  assign n1660 = n1622 & n1635 ;
  assign n1661 = n1623 & n1627 ;
  assign n1664 = ~n1660 & ~n1661 ;
  assign n1665 = ~n1663 & n1664 ;
  assign n1666 = ~n1642 & n1665 ;
  assign n1667 = n1640 & ~n1666 ;
  assign n1668 = n1629 & n1635 ;
  assign n1669 = n1640 & ~n1668 ;
  assign n1670 = n1618 & n1635 ;
  assign n1671 = n1621 & n1670 ;
  assign n1672 = n1627 & n1662 ;
  assign n1673 = ~n1629 & ~n1672 ;
  assign n1674 = ~n1671 & n1673 ;
  assign n1675 = ~n1669 & ~n1674 ;
  assign n1676 = ~n1667 & ~n1675 ;
  assign n1677 = n1658 & ~n1676 ;
  assign n1678 = ~n1627 & ~n1635 ;
  assign n1679 = ~n1624 & n1678 ;
  assign n1680 = ~n1640 & n1679 ;
  assign n1681 = ~n1635 & n1662 ;
  assign n1682 = ~n1660 & ~n1681 ;
  assign n1683 = ~n1627 & ~n1682 ;
  assign n1684 = n1640 & n1683 ;
  assign n1685 = ~n1680 & ~n1684 ;
  assign n1686 = ~n1677 & n1685 ;
  assign n1687 = ~n1659 & n1686 ;
  assign n1688 = ~\data_i[32]_pad  & n281 ;
  assign n1689 = ~\rd1_L_o_reg[3]/NET0131  & ~n281 ;
  assign n1690 = ~n1688 & ~n1689 ;
  assign n1691 = n1687 & ~n1690 ;
  assign n1692 = ~n1687 & n1690 ;
  assign n1693 = ~n1691 & ~n1692 ;
  assign n1715 = n1538 & ~n1559 ;
  assign n1716 = ~n1582 & n1715 ;
  assign n1717 = ~n1535 & n1716 ;
  assign n1718 = n1538 & n1560 ;
  assign n1719 = n1554 & n1592 ;
  assign n1705 = ~n1538 & n1582 ;
  assign n1720 = ~n1568 & ~n1705 ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1722 = ~n1718 & n1721 ;
  assign n1723 = ~n1554 & n1592 ;
  assign n1724 = n1568 & ~n1591 ;
  assign n1725 = ~n1597 & n1724 ;
  assign n1726 = ~n1723 & n1725 ;
  assign n1727 = ~n1722 & ~n1726 ;
  assign n1728 = ~n1717 & ~n1727 ;
  assign n1729 = n1579 & ~n1728 ;
  assign n1698 = n1538 & n1570 ;
  assign n1694 = ~n1535 & n1582 ;
  assign n1695 = n1538 & n1694 ;
  assign n1696 = ~n1538 & n1559 ;
  assign n1697 = ~n1554 & n1557 ;
  assign n1699 = ~n1696 & ~n1697 ;
  assign n1700 = ~n1695 & n1699 ;
  assign n1701 = ~n1698 & n1700 ;
  assign n1702 = ~n1568 & ~n1701 ;
  assign n1706 = n1535 & n1538 ;
  assign n1707 = ~n1554 & n1706 ;
  assign n1708 = ~n1705 & ~n1707 ;
  assign n1709 = n1568 & ~n1708 ;
  assign n1703 = n1538 & ~n1554 ;
  assign n1704 = n1597 & n1703 ;
  assign n1710 = n1550 & n1557 ;
  assign n1711 = ~n1704 & ~n1710 ;
  assign n1712 = ~n1709 & n1711 ;
  assign n1713 = ~n1702 & n1712 ;
  assign n1714 = ~n1579 & ~n1713 ;
  assign n1731 = ~n1555 & ~n1562 ;
  assign n1732 = n1568 & ~n1731 ;
  assign n1730 = n1535 & n1705 ;
  assign n1733 = ~n1535 & ~n1568 ;
  assign n1734 = n1696 & n1733 ;
  assign n1735 = ~n1730 & ~n1734 ;
  assign n1736 = ~n1732 & n1735 ;
  assign n1737 = ~n1714 & n1736 ;
  assign n1738 = ~n1729 & n1737 ;
  assign n1739 = ~\data_i[48]_pad  & n281 ;
  assign n1740 = ~\rd1_L_o_reg[1]/NET0131  & ~n281 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = n1738 & ~n1741 ;
  assign n1743 = ~n1738 & n1741 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1745 = n1105 & ~n1109 ;
  assign n1746 = n1137 & ~n1745 ;
  assign n1750 = ~n1098 & ~n1110 ;
  assign n1747 = n1109 & ~n1126 ;
  assign n1748 = ~n1101 & n1747 ;
  assign n1749 = n1126 & ~n1138 ;
  assign n1751 = ~n1748 & ~n1749 ;
  assign n1752 = n1750 & n1751 ;
  assign n1753 = ~n1746 & ~n1752 ;
  assign n1754 = n1126 & n1129 ;
  assign n1755 = ~n1753 & ~n1754 ;
  assign n1756 = n1158 & ~n1755 ;
  assign n1766 = n1101 & n1139 ;
  assign n1767 = ~n1168 & ~n1766 ;
  assign n1768 = ~n1158 & ~n1767 ;
  assign n1759 = n1106 & n1747 ;
  assign n1769 = ~n1109 & n1766 ;
  assign n1770 = ~n1759 & ~n1769 ;
  assign n1771 = ~n1768 & n1770 ;
  assign n1772 = n1098 & ~n1771 ;
  assign n1758 = ~n1098 & n1161 ;
  assign n1760 = ~n1143 & ~n1758 ;
  assign n1761 = ~n1759 & n1760 ;
  assign n1757 = ~n1098 & n1180 ;
  assign n1762 = ~n1165 & ~n1757 ;
  assign n1763 = n1761 & n1762 ;
  assign n1764 = ~n1158 & ~n1763 ;
  assign n1765 = ~n1098 & n1185 ;
  assign n1773 = ~n1764 & ~n1765 ;
  assign n1774 = ~n1772 & n1773 ;
  assign n1775 = ~n1756 & n1774 ;
  assign n1776 = ~\data_i[22]_pad  & n281 ;
  assign n1777 = ~\rd1_L_o_reg[29]/NET0131  & ~n281 ;
  assign n1778 = ~n1776 & ~n1777 ;
  assign n1779 = n1775 & ~n1778 ;
  assign n1780 = ~n1775 & n1778 ;
  assign n1781 = ~n1779 & ~n1780 ;
  assign n1785 = n1419 & ~n1448 ;
  assign n1794 = n1454 & ~n1785 ;
  assign n1795 = n1416 & ~n1467 ;
  assign n1796 = ~n1794 & n1795 ;
  assign n1786 = ~n1425 & ~n1440 ;
  assign n1803 = n1478 & n1786 ;
  assign n1804 = ~n1469 & ~n1803 ;
  assign n1805 = n1796 & n1804 ;
  assign n1787 = ~n1514 & ~n1786 ;
  assign n1788 = n1785 & n1787 ;
  assign n1789 = ~n1416 & ~n1788 ;
  assign n1802 = ~n1475 & n1789 ;
  assign n1806 = n1419 & ~n1802 ;
  assign n1807 = ~n1805 & n1806 ;
  assign n1797 = n1422 & ~n1468 ;
  assign n1798 = ~n1786 & n1797 ;
  assign n1799 = n1796 & ~n1798 ;
  assign n1790 = n1425 & n1478 ;
  assign n1791 = ~n1449 & ~n1453 ;
  assign n1792 = ~n1790 & n1791 ;
  assign n1793 = n1789 & ~n1792 ;
  assign n1800 = ~n1419 & ~n1793 ;
  assign n1801 = ~n1799 & n1800 ;
  assign n1782 = ~n1419 & ~n1440 ;
  assign n1783 = ~n1454 & ~n1782 ;
  assign n1784 = n1441 & ~n1783 ;
  assign n1808 = ~n1451 & ~n1784 ;
  assign n1809 = ~n1801 & n1808 ;
  assign n1810 = ~n1807 & n1809 ;
  assign n1811 = ~\data_i[56]_pad  & n281 ;
  assign n1812 = ~\rd1_L_o_reg[0]/NET0131  & ~n281 ;
  assign n1813 = ~n1811 & ~n1812 ;
  assign n1814 = n1810 & ~n1813 ;
  assign n1815 = ~n1810 & n1813 ;
  assign n1816 = ~n1814 & ~n1815 ;
  assign n1817 = ~n1126 & n1129 ;
  assign n1818 = n1098 & ~n1147 ;
  assign n1819 = ~n1817 & n1818 ;
  assign n1820 = n1104 & n1160 ;
  assign n1821 = ~n1098 & ~n1820 ;
  assign n1822 = ~n1759 & n1821 ;
  assign n1823 = ~n1819 & ~n1822 ;
  assign n1824 = ~n1110 & ~n1138 ;
  assign n1825 = n1126 & ~n1824 ;
  assign n1826 = ~n1158 & ~n1765 ;
  assign n1827 = ~n1825 & n1826 ;
  assign n1828 = ~n1823 & n1827 ;
  assign n1833 = n1158 & ~n1169 ;
  assign n1829 = n1098 & n1185 ;
  assign n1834 = ~n1757 & ~n1829 ;
  assign n1830 = ~n1142 & ~n1172 ;
  assign n1831 = n1106 & ~n1830 ;
  assign n1832 = ~n1139 & n1758 ;
  assign n1835 = ~n1831 & ~n1832 ;
  assign n1836 = n1834 & n1835 ;
  assign n1837 = n1833 & n1836 ;
  assign n1838 = ~n1828 & ~n1837 ;
  assign n1839 = n1098 & ~n1164 ;
  assign n1840 = ~n1101 & n1135 ;
  assign n1841 = ~n1098 & ~n1840 ;
  assign n1842 = ~n1754 & n1841 ;
  assign n1843 = ~n1769 & n1842 ;
  assign n1844 = ~n1839 & ~n1843 ;
  assign n1845 = ~n1838 & ~n1844 ;
  assign n1846 = ~\data_i[62]_pad  & n281 ;
  assign n1847 = ~\rd1_L_o_reg[24]/NET0131  & ~n281 ;
  assign n1848 = ~n1846 & ~n1847 ;
  assign n1849 = n1845 & ~n1848 ;
  assign n1850 = ~n1845 & n1848 ;
  assign n1851 = ~n1849 & ~n1850 ;
  assign n1852 = ~n266 & ~n622 ;
  assign n1853 = ~n562 & ~n1852 ;
  assign n1854 = ~decrypt_i_pad & ~n1853 ;
  assign n1855 = n292 & ~n704 ;
  assign n1856 = ~n972 & ~n1244 ;
  assign n1857 = ~n1855 & n1856 ;
  assign n1858 = decrypt_i_pad & ~n1857 ;
  assign n1859 = ~n1854 & ~n1858 ;
  assign n1860 = \rd1_R_o_reg[21]/NET0131  & ~n281 ;
  assign n1861 = \data_i[21]_pad  & n281 ;
  assign n1862 = ~n1860 & ~n1861 ;
  assign n1863 = ~n1859 & n1862 ;
  assign n1864 = n1859 & ~n1862 ;
  assign n1865 = ~n1863 & ~n1864 ;
  assign n1866 = ~n470 & n933 ;
  assign n1867 = n470 & ~n933 ;
  assign n1868 = ~n1866 & ~n1867 ;
  assign n1869 = ~n1865 & n1868 ;
  assign n1870 = ~n522 & n1297 ;
  assign n1871 = n522 & ~n1297 ;
  assign n1872 = ~n1870 & ~n1871 ;
  assign n1873 = ~n266 & ~n758 ;
  assign n1874 = ~n919 & ~n1873 ;
  assign n1875 = ~decrypt_i_pad & ~n1874 ;
  assign n1876 = n292 & ~n722 ;
  assign n1877 = ~n580 & ~n714 ;
  assign n1878 = ~n1876 & n1877 ;
  assign n1879 = decrypt_i_pad & ~n1878 ;
  assign n1880 = ~n1875 & ~n1879 ;
  assign n1881 = \rd1_R_o_reg[22]/NET0131  & ~n281 ;
  assign n1882 = \data_i[13]_pad  & n281 ;
  assign n1883 = ~n1881 & ~n1882 ;
  assign n1884 = ~n1880 & n1883 ;
  assign n1885 = n1880 & ~n1883 ;
  assign n1886 = ~n1884 & ~n1885 ;
  assign n1887 = n1872 & n1886 ;
  assign n1888 = ~n748 & n1266 ;
  assign n1889 = n748 & ~n1266 ;
  assign n1890 = ~n1888 & ~n1889 ;
  assign n1891 = n1872 & ~n1890 ;
  assign n1892 = ~n1872 & n1890 ;
  assign n1893 = ~n1891 & ~n1892 ;
  assign n1894 = ~n1886 & n1893 ;
  assign n1895 = ~n1887 & ~n1894 ;
  assign n1896 = n1869 & ~n1895 ;
  assign n1897 = ~n1865 & ~n1886 ;
  assign n1898 = n1865 & n1886 ;
  assign n1899 = ~n1897 & ~n1898 ;
  assign n1900 = ~n1891 & ~n1899 ;
  assign n1901 = n1872 & ~n1897 ;
  assign n1902 = ~n1868 & ~n1901 ;
  assign n1903 = ~n1900 & n1902 ;
  assign n1907 = n1865 & ~n1872 ;
  assign n1910 = n1886 & n1907 ;
  assign n1911 = n1868 & n1910 ;
  assign n1904 = ~n585 & n905 ;
  assign n1905 = n585 & ~n905 ;
  assign n1906 = ~n1904 & ~n1905 ;
  assign n1908 = n1890 & n1907 ;
  assign n1909 = ~n1886 & n1908 ;
  assign n1912 = n1906 & ~n1909 ;
  assign n1913 = ~n1911 & n1912 ;
  assign n1914 = ~n1903 & n1913 ;
  assign n1915 = ~n1896 & n1914 ;
  assign n1919 = ~n1872 & ~n1886 ;
  assign n1920 = ~n1887 & ~n1919 ;
  assign n1921 = ~n1890 & ~n1907 ;
  assign n1922 = ~n1920 & n1921 ;
  assign n1923 = n1872 & n1890 ;
  assign n1924 = ~n1865 & n1923 ;
  assign n1925 = ~n1910 & ~n1924 ;
  assign n1926 = ~n1922 & n1925 ;
  assign n1927 = ~n1868 & ~n1926 ;
  assign n1916 = n1865 & ~n1890 ;
  assign n1917 = ~n1886 & n1916 ;
  assign n1918 = n1872 & n1917 ;
  assign n1928 = ~n1906 & ~n1918 ;
  assign n1929 = ~n1927 & n1928 ;
  assign n1930 = ~n1915 & ~n1929 ;
  assign n1931 = n1906 & ~n1918 ;
  assign n1933 = ~n1907 & ~n1923 ;
  assign n1934 = n1920 & n1933 ;
  assign n1932 = ~n1865 & n1892 ;
  assign n1935 = ~n1917 & ~n1932 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = ~n1931 & ~n1936 ;
  assign n1938 = n1898 & n1923 ;
  assign n1939 = n1868 & ~n1938 ;
  assign n1940 = ~n1937 & n1939 ;
  assign n1941 = ~n1865 & n1890 ;
  assign n1942 = ~n1916 & ~n1941 ;
  assign n1943 = n1887 & ~n1942 ;
  assign n1944 = ~n1868 & ~n1909 ;
  assign n1945 = ~n1943 & n1944 ;
  assign n1946 = ~n1940 & ~n1945 ;
  assign n1947 = ~n1930 & ~n1946 ;
  assign n1948 = ~\data_i[58]_pad  & n281 ;
  assign n1949 = ~\rd1_L_o_reg[8]/NET0131  & ~n281 ;
  assign n1950 = ~n1948 & ~n1949 ;
  assign n1951 = n1947 & ~n1950 ;
  assign n1952 = ~n1947 & n1950 ;
  assign n1953 = ~n1951 & ~n1952 ;
  assign n1959 = n1239 & n1261 ;
  assign n1960 = ~n1258 & ~n1959 ;
  assign n1961 = ~n1263 & ~n1960 ;
  assign n1957 = ~n1239 & ~n1257 ;
  assign n1958 = n1302 & n1957 ;
  assign n1962 = ~n1300 & ~n1958 ;
  assign n1963 = ~n1961 & n1962 ;
  assign n1964 = ~n1262 & n1300 ;
  assign n1965 = ~n1276 & n1964 ;
  assign n1966 = n1274 & n1965 ;
  assign n1967 = ~n1963 & ~n1966 ;
  assign n1968 = n1269 & ~n1967 ;
  assign n1972 = n1261 & ~n1309 ;
  assign n1973 = ~n1324 & ~n1972 ;
  assign n1970 = ~n1261 & n1303 ;
  assign n1971 = ~n1300 & ~n1970 ;
  assign n1974 = ~n1263 & n1971 ;
  assign n1975 = ~n1973 & n1974 ;
  assign n1977 = ~n1257 & ~n1272 ;
  assign n1978 = ~n1275 & n1977 ;
  assign n1976 = n1258 & ~n1261 ;
  assign n1979 = n1300 & ~n1976 ;
  assign n1980 = ~n1978 & n1979 ;
  assign n1981 = ~n1975 & ~n1980 ;
  assign n1954 = n1239 & ~n1300 ;
  assign n1969 = n1282 & ~n1954 ;
  assign n1982 = ~n1269 & ~n1969 ;
  assign n1983 = ~n1981 & n1982 ;
  assign n1984 = ~n1968 & ~n1983 ;
  assign n1955 = ~n1257 & n1307 ;
  assign n1956 = n1954 & n1955 ;
  assign n1985 = ~n1319 & ~n1956 ;
  assign n1986 = ~n1984 & n1985 ;
  assign n1987 = ~\data_i[36]_pad  & n281 ;
  assign n1988 = ~\rd1_L_o_reg[19]/NET0131  & ~n281 ;
  assign n1989 = ~n1987 & ~n1988 ;
  assign n1990 = n1986 & ~n1989 ;
  assign n1991 = ~n1986 & n1989 ;
  assign n1992 = ~n1990 & ~n1991 ;
  assign n2015 = ~n1627 & n1670 ;
  assign n2016 = ~n1621 & n2015 ;
  assign n2017 = n1640 & ~n1642 ;
  assign n2018 = ~n2016 & n2017 ;
  assign n2019 = n1618 & n1678 ;
  assign n2004 = n1618 & n1629 ;
  assign n2020 = ~n1640 & ~n2004 ;
  assign n2021 = ~n2019 & n2020 ;
  assign n2022 = ~n2018 & ~n2021 ;
  assign n2005 = ~n1635 & n2004 ;
  assign n2023 = ~n1683 & ~n2005 ;
  assign n2024 = ~n2022 & n2023 ;
  assign n2025 = ~n1658 & ~n2024 ;
  assign n2006 = ~n1648 & ~n1661 ;
  assign n2007 = n1635 & ~n2006 ;
  assign n2008 = n1622 & n1627 ;
  assign n2009 = ~n1635 & n2008 ;
  assign n2010 = ~n2005 & ~n2009 ;
  assign n2011 = ~n2007 & n2010 ;
  assign n2012 = ~n1640 & ~n2011 ;
  assign n1994 = ~n1671 & ~n1679 ;
  assign n1995 = n1640 & ~n1994 ;
  assign n1996 = n1635 & n1662 ;
  assign n1997 = ~n1661 & ~n1996 ;
  assign n1998 = ~n1640 & ~n1997 ;
  assign n1993 = n1635 & n1641 ;
  assign n1999 = n1635 & n1663 ;
  assign n2000 = ~n1993 & ~n1999 ;
  assign n2001 = ~n1998 & n2000 ;
  assign n2002 = ~n1995 & n2001 ;
  assign n2003 = n1658 & ~n2002 ;
  assign n2013 = n1627 & n1640 ;
  assign n2014 = ~n1682 & n2013 ;
  assign n2026 = ~n2003 & ~n2014 ;
  assign n2027 = ~n2012 & n2026 ;
  assign n2028 = ~n2025 & n2027 ;
  assign n2029 = ~\data_i[20]_pad  & n281 ;
  assign n2030 = ~\rd1_L_o_reg[21]/NET0131  & ~n281 ;
  assign n2031 = ~n2029 & ~n2030 ;
  assign n2032 = n2028 & ~n2031 ;
  assign n2033 = ~n2028 & n2031 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2046 = ~n942 & ~n1004 ;
  assign n2045 = n895 & ~n960 ;
  assign n2047 = ~n958 & ~n2045 ;
  assign n2048 = n2046 & n2047 ;
  assign n2044 = n908 & n989 ;
  assign n2049 = ~n987 & ~n1374 ;
  assign n2050 = ~n2044 & n2049 ;
  assign n2051 = ~n2048 & n2050 ;
  assign n2055 = n987 & ~n1006 ;
  assign n2052 = n895 & ~n1359 ;
  assign n2053 = ~n1010 & ~n1356 ;
  assign n2054 = ~n958 & ~n2053 ;
  assign n2056 = ~n2052 & ~n2054 ;
  assign n2057 = n2055 & n2056 ;
  assign n2058 = ~n2051 & ~n2057 ;
  assign n2040 = n941 & ~n1387 ;
  assign n2035 = ~n895 & ~n995 ;
  assign n2036 = n895 & n901 ;
  assign n2037 = ~n936 & n2036 ;
  assign n2038 = ~n1356 & ~n2037 ;
  assign n2039 = ~n987 & ~n2038 ;
  assign n2041 = ~n2035 & ~n2039 ;
  assign n2042 = ~n2040 & n2041 ;
  assign n2043 = n958 & ~n2042 ;
  assign n2059 = ~n895 & n1365 ;
  assign n2060 = ~n990 & ~n2059 ;
  assign n2061 = n908 & ~n2060 ;
  assign n2062 = ~n2043 & ~n2061 ;
  assign n2063 = ~n2058 & n2062 ;
  assign n2064 = ~\data_i[26]_pad  & n281 ;
  assign n2065 = ~\rd1_L_o_reg[12]/NET0131  & ~n281 ;
  assign n2066 = ~n2064 & ~n2065 ;
  assign n2067 = n2063 & ~n2066 ;
  assign n2068 = ~n2063 & n2066 ;
  assign n2069 = ~n2067 & ~n2068 ;
  assign n2076 = ~n1872 & n1897 ;
  assign n2074 = n1865 & n1923 ;
  assign n2075 = ~n1890 & n1919 ;
  assign n2077 = ~n2074 & ~n2075 ;
  assign n2078 = ~n2076 & n2077 ;
  assign n2079 = ~n1868 & ~n2078 ;
  assign n2070 = n1893 & n1898 ;
  assign n2071 = ~n1890 & n1920 ;
  assign n2072 = ~n1909 & ~n2071 ;
  assign n2073 = n1868 & ~n2072 ;
  assign n2080 = ~n2070 & ~n2073 ;
  assign n2081 = ~n2079 & n2080 ;
  assign n2082 = ~n1906 & ~n2081 ;
  assign n2087 = ~n1872 & ~n1942 ;
  assign n2086 = n1872 & n1942 ;
  assign n2088 = ~n1868 & ~n2086 ;
  assign n2089 = ~n2087 & n2088 ;
  assign n2083 = n1886 & n1892 ;
  assign n2084 = n1865 & n2083 ;
  assign n2085 = n1868 & n1894 ;
  assign n2090 = ~n2084 & ~n2085 ;
  assign n2091 = ~n2089 & n2090 ;
  assign n2092 = n1906 & ~n2091 ;
  assign n2093 = ~n1865 & n1887 ;
  assign n2094 = ~n1890 & n2093 ;
  assign n2095 = n1869 & n1890 ;
  assign n2096 = n1920 & n2095 ;
  assign n2097 = ~n2094 & ~n2096 ;
  assign n2098 = ~n2092 & n2097 ;
  assign n2099 = ~n2082 & n2098 ;
  assign n2100 = ~\data_i[60]_pad  & n281 ;
  assign n2101 = ~\rd1_L_o_reg[16]/NET0131  & ~n281 ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2103 = n2099 & ~n2102 ;
  assign n2104 = ~n2099 & n2102 ;
  assign n2105 = ~n2103 & ~n2104 ;
  assign n2121 = ~n783 & ~n803 ;
  assign n2122 = ~n825 & ~n2121 ;
  assign n2123 = n822 & ~n869 ;
  assign n2124 = ~n2122 & n2123 ;
  assign n2120 = ~n799 & n868 ;
  assign n2116 = n799 & ~n822 ;
  assign n2117 = ~n839 & ~n2116 ;
  assign n2118 = ~n783 & n837 ;
  assign n2119 = ~n2117 & n2118 ;
  assign n2125 = n862 & ~n2119 ;
  assign n2126 = ~n2120 & n2125 ;
  assign n2127 = ~n2124 & n2126 ;
  assign n2128 = ~n829 & ~n831 ;
  assign n2129 = ~n799 & ~n837 ;
  assign n2130 = ~n2128 & n2129 ;
  assign n2131 = n822 & n837 ;
  assign n2132 = n2121 & n2131 ;
  assign n2133 = ~n862 & ~n2132 ;
  assign n2134 = ~n2130 & n2133 ;
  assign n2135 = n827 & n2134 ;
  assign n2136 = ~n2127 & ~n2135 ;
  assign n2106 = n804 & n822 ;
  assign n2107 = n822 & n825 ;
  assign n2108 = ~n2106 & ~n2107 ;
  assign n2109 = n783 & n828 ;
  assign n2110 = n837 & ~n2109 ;
  assign n2111 = n2108 & n2110 ;
  assign n2112 = ~n822 & n831 ;
  assign n2113 = ~n837 & ~n870 ;
  assign n2114 = ~n2112 & n2113 ;
  assign n2115 = ~n2111 & ~n2114 ;
  assign n2137 = ~n783 & n839 ;
  assign n2138 = ~n822 & n2137 ;
  assign n2139 = ~n2115 & ~n2138 ;
  assign n2140 = ~n2136 & n2139 ;
  assign n2141 = ~\data_i[52]_pad  & n281 ;
  assign n2142 = ~\rd1_L_o_reg[17]/NET0131  & ~n281 ;
  assign n2143 = ~n2141 & ~n2142 ;
  assign n2144 = n2140 & ~n2143 ;
  assign n2145 = ~n2140 & n2143 ;
  assign n2146 = ~n2144 & ~n2145 ;
  assign n2148 = ~n1419 & ~n1454 ;
  assign n2149 = ~n1466 & n2148 ;
  assign n2150 = n1416 & ~n2149 ;
  assign n2147 = ~n1432 & n1466 ;
  assign n2151 = ~n1460 & ~n1511 ;
  assign n2152 = ~n2147 & n2151 ;
  assign n2153 = ~n2150 & n2152 ;
  assign n2157 = ~n1416 & n1419 ;
  assign n2158 = ~n1462 & ~n2157 ;
  assign n2154 = ~n1416 & ~n1786 ;
  assign n2155 = ~n1419 & ~n2154 ;
  assign n2156 = ~n1432 & n1473 ;
  assign n2159 = ~n2155 & ~n2156 ;
  assign n2160 = n2158 & n2159 ;
  assign n2161 = ~n2153 & ~n2160 ;
  assign n2162 = n1419 & n1440 ;
  assign n2163 = n1472 & n2162 ;
  assign n2164 = n1452 & n1782 ;
  assign n2165 = ~n2163 & ~n2164 ;
  assign n2166 = ~n1495 & n2165 ;
  assign n2167 = ~n2161 & n2166 ;
  assign n2168 = ~\data_i[28]_pad  & n281 ;
  assign n2169 = ~\rd1_L_o_reg[20]/NET0131  & ~n281 ;
  assign n2170 = ~n2168 & ~n2169 ;
  assign n2171 = n2167 & ~n2170 ;
  assign n2172 = ~n2167 & n2170 ;
  assign n2173 = ~n2171 & ~n2172 ;
  assign n2174 = ~n1571 & ~n1581 ;
  assign n2175 = n1598 & n2174 ;
  assign n2176 = n1535 & n1696 ;
  assign n2177 = n1568 & ~n1716 ;
  assign n2178 = ~n2176 & n2177 ;
  assign n2179 = ~n2175 & ~n2178 ;
  assign n2180 = n1579 & ~n2179 ;
  assign n2181 = n1550 & n1706 ;
  assign n2182 = ~n1560 & ~n2181 ;
  assign n2183 = ~n1568 & ~n2182 ;
  assign n2188 = ~n1579 & ~n1718 ;
  assign n2189 = ~n2183 & n2188 ;
  assign n2184 = n1568 & n1592 ;
  assign n2185 = ~n1733 & ~n2184 ;
  assign n2186 = ~n1550 & ~n2185 ;
  assign n2187 = n1568 & ~n1584 ;
  assign n2190 = ~n2186 & ~n2187 ;
  assign n2191 = n2189 & n2190 ;
  assign n2192 = ~n2180 & ~n2191 ;
  assign n2193 = ~n1695 & ~n1704 ;
  assign n2194 = ~n1568 & ~n2193 ;
  assign n2195 = ~n1535 & n1568 ;
  assign n2196 = ~n1599 & n2195 ;
  assign n2197 = ~n1715 & n2196 ;
  assign n2198 = ~n2194 & ~n2197 ;
  assign n2199 = ~n2192 & n2198 ;
  assign n2200 = ~\data_i[4]_pad  & n281 ;
  assign n2201 = ~\rd1_L_o_reg[23]/NET0131  & ~n281 ;
  assign n2202 = ~n2200 & ~n2201 ;
  assign n2203 = n2199 & ~n2202 ;
  assign n2204 = ~n2199 & n2202 ;
  assign n2205 = ~n2203 & ~n2204 ;
  assign n2212 = n1622 & ~n1635 ;
  assign n2213 = ~n1654 & ~n2212 ;
  assign n2214 = ~n1671 & n2213 ;
  assign n2215 = ~n1640 & ~n2214 ;
  assign n2219 = ~n1635 & ~n2006 ;
  assign n2216 = n1629 & n1640 ;
  assign n2217 = ~n1670 & n2216 ;
  assign n2218 = n1635 & n1672 ;
  assign n2220 = ~n2217 & ~n2218 ;
  assign n2221 = ~n2219 & n2220 ;
  assign n2222 = ~n2215 & n2221 ;
  assign n2223 = ~n1658 & ~n2222 ;
  assign n2206 = n1624 & n1649 ;
  assign n2207 = ~n2007 & ~n2206 ;
  assign n2208 = n1658 & ~n2207 ;
  assign n2209 = ~n1635 & n1654 ;
  assign n2210 = ~n2208 & ~n2209 ;
  assign n2211 = ~n1640 & ~n2210 ;
  assign n2224 = n1621 & n1627 ;
  assign n2225 = ~n2015 & ~n2224 ;
  assign n2226 = n1640 & ~n2225 ;
  assign n2227 = n1635 & n2008 ;
  assign n2228 = ~n2226 & ~n2227 ;
  assign n2229 = n1658 & ~n2228 ;
  assign n2230 = n1618 & n2224 ;
  assign n2231 = n1635 & ~n2230 ;
  assign n2232 = n1640 & ~n1649 ;
  assign n2233 = ~n2231 & n2232 ;
  assign n2234 = ~n2229 & ~n2233 ;
  assign n2235 = ~n2211 & n2234 ;
  assign n2236 = ~n2223 & n2235 ;
  assign n2237 = ~\data_i[30]_pad  & n281 ;
  assign n2238 = ~\rd1_L_o_reg[28]/NET0131  & ~n281 ;
  assign n2239 = ~n2237 & ~n2238 ;
  assign n2240 = n2236 & ~n2239 ;
  assign n2241 = ~n2236 & n2239 ;
  assign n2242 = ~n2240 & ~n2241 ;
  assign n2258 = ~n1585 & ~n1697 ;
  assign n2259 = ~n1568 & ~n2258 ;
  assign n2260 = n1568 & n1581 ;
  assign n2261 = ~n1564 & ~n2260 ;
  assign n2262 = ~n2259 & n2261 ;
  assign n2263 = ~n1579 & ~n2262 ;
  assign n2247 = ~n1538 & ~n1585 ;
  assign n2248 = ~n1551 & n1568 ;
  assign n2249 = ~n2247 & n2248 ;
  assign n2250 = ~n1704 & ~n2176 ;
  assign n2251 = ~n2249 & n2250 ;
  assign n2252 = n1579 & ~n2251 ;
  assign n2243 = ~n1570 & ~n1694 ;
  assign n2244 = n1579 & ~n2243 ;
  assign n2245 = ~n1698 & ~n2244 ;
  assign n2246 = ~n1568 & ~n2245 ;
  assign n2253 = ~n1560 & ~n1707 ;
  assign n2254 = n1568 & ~n2253 ;
  assign n2255 = ~n1538 & ~n1591 ;
  assign n2256 = ~n1703 & n2195 ;
  assign n2257 = ~n2255 & n2256 ;
  assign n2264 = ~n1604 & ~n2257 ;
  assign n2265 = ~n2254 & n2264 ;
  assign n2266 = ~n2246 & n2265 ;
  assign n2267 = ~n2252 & n2266 ;
  assign n2268 = ~n2263 & n2267 ;
  assign n2269 = ~\data_i[2]_pad  & n281 ;
  assign n2270 = ~\rd1_L_o_reg[15]/NET0131  & ~n281 ;
  assign n2271 = ~n2269 & ~n2270 ;
  assign n2272 = n2268 & ~n2271 ;
  assign n2273 = ~n2268 & n2271 ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = ~n1261 & ~n1322 ;
  assign n2279 = ~n1303 & n2275 ;
  assign n2280 = ~n1257 & n1261 ;
  assign n2281 = n1242 & n2280 ;
  assign n2282 = ~n2279 & ~n2281 ;
  assign n2283 = ~n1300 & ~n2282 ;
  assign n2276 = n1300 & ~n1317 ;
  assign n2277 = ~n2275 & n2276 ;
  assign n2284 = n1257 & n2277 ;
  assign n2285 = ~n1308 & ~n2284 ;
  assign n2286 = ~n2283 & n2285 ;
  assign n2287 = n1269 & ~n2286 ;
  assign n2291 = ~n1282 & ~n1324 ;
  assign n2292 = n1239 & ~n2280 ;
  assign n2293 = ~n1271 & n2292 ;
  assign n2294 = ~n2291 & ~n2293 ;
  assign n2295 = n1300 & ~n2294 ;
  assign n2288 = ~n1242 & n1317 ;
  assign n2289 = ~n1282 & ~n2288 ;
  assign n2290 = n1971 & n2289 ;
  assign n2296 = ~n1269 & ~n2290 ;
  assign n2297 = ~n2295 & n2296 ;
  assign n2298 = n1239 & n1976 ;
  assign n2299 = n1261 & n1322 ;
  assign n2300 = ~n2298 & ~n2299 ;
  assign n2301 = ~n1300 & ~n2300 ;
  assign n2278 = ~n1242 & n2277 ;
  assign n2302 = ~n1958 & ~n2278 ;
  assign n2303 = ~n2301 & n2302 ;
  assign n2304 = ~n2297 & n2303 ;
  assign n2305 = ~n2287 & n2304 ;
  assign n2306 = ~\data_i[24]_pad  & n281 ;
  assign n2307 = ~\rd1_L_o_reg[4]/NET0131  & ~n281 ;
  assign n2308 = ~n2306 & ~n2307 ;
  assign n2309 = n2305 & ~n2308 ;
  assign n2310 = ~n2305 & n2308 ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2312 = ~n1160 & n1173 ;
  assign n2313 = ~n1098 & ~n1109 ;
  assign n2314 = n1820 & ~n2313 ;
  assign n2315 = ~n1158 & ~n2314 ;
  assign n2316 = ~n1754 & n2315 ;
  assign n2317 = ~n2312 & n2316 ;
  assign n2319 = ~n1110 & ~n1135 ;
  assign n2320 = n1098 & ~n2319 ;
  assign n2318 = ~n1098 & n1147 ;
  assign n2321 = ~n1136 & n1158 ;
  assign n2322 = ~n1817 & n2321 ;
  assign n2323 = ~n2318 & n2322 ;
  assign n2324 = ~n2320 & n2323 ;
  assign n2325 = ~n2317 & ~n2324 ;
  assign n2326 = ~n1143 & ~n1148 ;
  assign n2327 = ~n1098 & ~n2326 ;
  assign n2331 = ~n1110 & ~n1149 ;
  assign n2332 = ~n1098 & ~n1158 ;
  assign n2333 = ~n2331 & n2332 ;
  assign n2329 = ~n1105 & ~n1106 ;
  assign n2330 = n1173 & n2329 ;
  assign n2328 = n1181 & n1745 ;
  assign n2334 = ~n1769 & ~n2328 ;
  assign n2335 = ~n2330 & n2334 ;
  assign n2336 = ~n2333 & n2335 ;
  assign n2337 = ~n2327 & n2336 ;
  assign n2338 = ~n2325 & n2337 ;
  assign n2339 = ~\data_i[0]_pad  & n281 ;
  assign n2340 = ~\rd1_L_o_reg[7]/NET0131  & ~n281 ;
  assign n2341 = ~n2339 & ~n2340 ;
  assign n2342 = n2338 & ~n2341 ;
  assign n2343 = ~n2338 & n2341 ;
  assign n2344 = ~n2342 & ~n2343 ;
  assign n2345 = n1886 & ~n1893 ;
  assign n2346 = ~n1894 & ~n2345 ;
  assign n2349 = ~n1906 & n2346 ;
  assign n2347 = n1906 & ~n1907 ;
  assign n2348 = ~n2346 & n2347 ;
  assign n2350 = ~n1890 & n1910 ;
  assign n2351 = ~n1909 & ~n2350 ;
  assign n2352 = ~n2348 & n2351 ;
  assign n2353 = ~n2349 & n2352 ;
  assign n2354 = ~n1868 & ~n2353 ;
  assign n2355 = ~n2083 & ~n2086 ;
  assign n2356 = n1868 & ~n2355 ;
  assign n2357 = n1865 & n2075 ;
  assign n2358 = ~n2356 & ~n2357 ;
  assign n2359 = ~n1906 & ~n2358 ;
  assign n2360 = n1906 & ~n1942 ;
  assign n2361 = ~n2083 & n2360 ;
  assign n2362 = ~n2084 & ~n2361 ;
  assign n2363 = n1868 & ~n2362 ;
  assign n2364 = ~n2359 & ~n2363 ;
  assign n2365 = ~n2354 & n2364 ;
  assign n2366 = ~\data_i[46]_pad  & n281 ;
  assign n2367 = ~\rd1_L_o_reg[26]/NET0131  & ~n281 ;
  assign n2368 = ~n2366 & ~n2367 ;
  assign n2369 = n2365 & ~n2368 ;
  assign n2370 = ~n2365 & n2368 ;
  assign n2371 = ~n2369 & ~n2370 ;
  assign n2376 = ~n1908 & ~n2075 ;
  assign n2377 = ~n2093 & n2376 ;
  assign n2378 = ~n1868 & ~n2377 ;
  assign n2372 = ~n1886 & n2074 ;
  assign n2373 = ~n1897 & ~n2074 ;
  assign n2374 = ~n2071 & n2373 ;
  assign n2375 = n1868 & ~n2374 ;
  assign n2379 = ~n2372 & ~n2375 ;
  assign n2380 = ~n2378 & n2379 ;
  assign n2381 = n1906 & ~n2380 ;
  assign n2384 = n1865 & ~n1906 ;
  assign n2385 = ~n1923 & n2384 ;
  assign n2386 = ~n1920 & n2385 ;
  assign n2382 = ~n1887 & ~n1892 ;
  assign n2383 = ~n1916 & n2382 ;
  assign n2387 = n1868 & ~n2383 ;
  assign n2388 = ~n2386 & n2387 ;
  assign n2389 = n1890 & ~n1899 ;
  assign n2390 = ~n1897 & n2071 ;
  assign n2391 = ~n2389 & ~n2390 ;
  assign n2392 = ~n1906 & ~n2391 ;
  assign n2393 = ~n1868 & ~n2094 ;
  assign n2394 = ~n2392 & n2393 ;
  assign n2395 = ~n2388 & ~n2394 ;
  assign n2396 = ~n2381 & ~n2395 ;
  assign n2397 = ~\data_i[40]_pad  & n281 ;
  assign n2398 = ~\rd1_L_o_reg[2]/NET0131  & ~n281 ;
  assign n2399 = ~n2397 & ~n2398 ;
  assign n2400 = n2396 & ~n2399 ;
  assign n2401 = ~n2396 & n2399 ;
  assign n2402 = ~n2400 & ~n2401 ;
  assign n2406 = ~n1300 & ~n1323 ;
  assign n2405 = n1257 & n1959 ;
  assign n2407 = ~n1955 & ~n2405 ;
  assign n2408 = n2406 & n2407 ;
  assign n2409 = n1300 & ~n1304 ;
  assign n2410 = ~n2288 & n2409 ;
  assign n2411 = ~n2408 & ~n2410 ;
  assign n2404 = ~n1242 & n1970 ;
  assign n2403 = ~n1277 & ~n2275 ;
  assign n2412 = n1269 & ~n2403 ;
  assign n2413 = ~n2404 & n2412 ;
  assign n2414 = ~n2411 & n2413 ;
  assign n2415 = ~n1309 & ~n1322 ;
  assign n2416 = ~n2280 & n2415 ;
  assign n2417 = n1300 & ~n2416 ;
  assign n2418 = ~n1282 & ~n1309 ;
  assign n2419 = n2406 & n2418 ;
  assign n2420 = ~n2417 & ~n2419 ;
  assign n2421 = ~n1269 & ~n1318 ;
  assign n2422 = ~n2298 & n2421 ;
  assign n2423 = ~n2420 & n2422 ;
  assign n2424 = ~n2414 & ~n2423 ;
  assign n2425 = ~\data_i[10]_pad  & n281 ;
  assign n2426 = ~\rd1_L_o_reg[14]/NET0131  & ~n281 ;
  assign n2427 = ~n2425 & ~n2426 ;
  assign n2428 = n2424 & ~n2427 ;
  assign n2429 = ~n2424 & n2427 ;
  assign n2430 = ~n2428 & ~n2429 ;
  assign n2439 = ~n1002 & n2046 ;
  assign n2440 = n958 & ~n2439 ;
  assign n2435 = ~n901 & n941 ;
  assign n2436 = ~n939 & n2036 ;
  assign n2437 = ~n1358 & ~n2436 ;
  assign n2438 = ~n958 & ~n2437 ;
  assign n2441 = ~n2435 & ~n2438 ;
  assign n2442 = ~n2440 & n2441 ;
  assign n2443 = ~n987 & ~n2442 ;
  assign n2431 = n995 & n2046 ;
  assign n2432 = ~n958 & ~n2431 ;
  assign n2433 = n1371 & ~n2432 ;
  assign n2434 = n987 & ~n2433 ;
  assign n2444 = ~n1386 & ~n2036 ;
  assign n2445 = ~n902 & ~n991 ;
  assign n2446 = n1388 & ~n2445 ;
  assign n2447 = ~n2444 & ~n2446 ;
  assign n2448 = ~n2434 & n2447 ;
  assign n2449 = ~n2443 & n2448 ;
  assign n2450 = ~\data_i[6]_pad  & n281 ;
  assign n2451 = ~\rd1_L_o_reg[31]/NET0131  & ~n281 ;
  assign n2452 = ~n2450 & ~n2451 ;
  assign n2453 = n2449 & ~n2452 ;
  assign n2454 = ~n2449 & n2452 ;
  assign n2455 = ~n2453 & ~n2454 ;
  assign n2462 = n837 & n862 ;
  assign n2476 = ~n803 & n2116 ;
  assign n2477 = ~n866 & ~n2476 ;
  assign n2478 = n862 & ~n2477 ;
  assign n2479 = ~n831 & n876 ;
  assign n2480 = ~n866 & ~n2479 ;
  assign n2481 = n837 & ~n2480 ;
  assign n2482 = ~n2478 & ~n2481 ;
  assign n2483 = ~n2462 & ~n2482 ;
  assign n2468 = n783 & n866 ;
  assign n2456 = n799 & n870 ;
  assign n2469 = n837 & ~n2456 ;
  assign n2470 = ~n2468 & n2469 ;
  assign n2471 = ~n2109 & ~n2137 ;
  assign n2472 = n822 & ~n2471 ;
  assign n2473 = ~n825 & ~n837 ;
  assign n2474 = ~n2472 & n2473 ;
  assign n2475 = ~n2470 & ~n2474 ;
  assign n2458 = ~n800 & ~n824 ;
  assign n2459 = ~n804 & ~n822 ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = ~n2138 & ~n2460 ;
  assign n2463 = ~n2461 & n2462 ;
  assign n2464 = ~n804 & ~n868 ;
  assign n2465 = ~n2137 & n2464 ;
  assign n2466 = ~n837 & ~n862 ;
  assign n2467 = ~n2465 & n2466 ;
  assign n2457 = ~n862 & n2456 ;
  assign n2484 = ~n2106 & ~n2457 ;
  assign n2485 = ~n2467 & n2484 ;
  assign n2486 = ~n2463 & n2485 ;
  assign n2487 = ~n2475 & n2486 ;
  assign n2488 = ~n2483 & n2487 ;
  assign n2489 = ~\data_i[34]_pad  & n281 ;
  assign n2490 = ~\rd1_L_o_reg[11]/NET0131  & ~n281 ;
  assign n2491 = ~n2489 & ~n2490 ;
  assign n2492 = n2488 & ~n2491 ;
  assign n2493 = ~n2488 & n2491 ;
  assign n2494 = ~n2492 & ~n2493 ;
  assign n2495 = n800 & n875 ;
  assign n2496 = n837 & ~n2495 ;
  assign n2497 = ~n823 & n2496 ;
  assign n2498 = ~n2107 & ~n2138 ;
  assign n2499 = n2497 & n2498 ;
  assign n2500 = ~n837 & ~n866 ;
  assign n2501 = ~n2106 & n2500 ;
  assign n2502 = ~n2499 & ~n2501 ;
  assign n2505 = n822 & n2137 ;
  assign n2506 = ~n2109 & ~n2476 ;
  assign n2507 = ~n2505 & n2506 ;
  assign n2508 = ~n837 & ~n2507 ;
  assign n2503 = n783 & ~n828 ;
  assign n2504 = n2131 & n2503 ;
  assign n2509 = ~n862 & ~n2468 ;
  assign n2510 = ~n2504 & n2509 ;
  assign n2511 = n2108 & n2510 ;
  assign n2512 = ~n2508 & n2511 ;
  assign n2513 = n799 & n822 ;
  assign n2514 = n2121 & n2513 ;
  assign n2520 = n862 & ~n2514 ;
  assign n2521 = ~n826 & n2520 ;
  assign n2515 = n783 & ~n837 ;
  assign n2516 = n822 & ~n839 ;
  assign n2517 = n2515 & ~n2516 ;
  assign n2518 = n822 & n828 ;
  assign n2519 = ~n2515 & n2518 ;
  assign n2522 = ~n2517 & ~n2519 ;
  assign n2523 = n2521 & n2522 ;
  assign n2524 = ~n2512 & ~n2523 ;
  assign n2525 = ~n2502 & ~n2524 ;
  assign n2526 = ~\data_i[38]_pad  & n281 ;
  assign n2527 = ~\rd1_L_o_reg[27]/NET0131  & ~n281 ;
  assign n2528 = ~n2526 & ~n2527 ;
  assign n2529 = n2525 & ~n2528 ;
  assign n2530 = ~n2525 & n2528 ;
  assign n2531 = ~n2529 & ~n2530 ;
  assign n2532 = ~n1672 & ~n2004 ;
  assign n2543 = ~n1635 & ~n2532 ;
  assign n2544 = ~n1640 & ~n1682 ;
  assign n2545 = ~n2216 & ~n2544 ;
  assign n2546 = ~n2543 & n2545 ;
  assign n2547 = ~n1658 & ~n2546 ;
  assign n2537 = ~n2212 & ~n2230 ;
  assign n2538 = ~n1640 & ~n2537 ;
  assign n2535 = ~n1663 & ~n2008 ;
  assign n2536 = n1640 & ~n2535 ;
  assign n2539 = ~n1999 & ~n2209 ;
  assign n2540 = ~n2536 & n2539 ;
  assign n2541 = ~n2538 & n2540 ;
  assign n2542 = n1658 & ~n2541 ;
  assign n2533 = n1635 & n1640 ;
  assign n2534 = ~n2532 & n2533 ;
  assign n2548 = ~n1623 & ~n1993 ;
  assign n2549 = ~n1635 & ~n1640 ;
  assign n2550 = ~n2533 & ~n2549 ;
  assign n2551 = ~n2548 & n2550 ;
  assign n2552 = ~n2534 & ~n2551 ;
  assign n2553 = ~n2542 & n2552 ;
  assign n2554 = ~n2547 & n2553 ;
  assign n2555 = ~\data_i[18]_pad  & n281 ;
  assign n2556 = ~\rd1_L_o_reg[13]/NET0131  & ~n281 ;
  assign n2557 = ~n2555 & ~n2556 ;
  assign n2558 = n2554 & ~n2557 ;
  assign n2559 = ~n2554 & n2557 ;
  assign n2560 = ~n2558 & ~n2559 ;
  assign n2561 = ~n440 & ~n1087 ;
  assign n2562 = ~n1204 & n2561 ;
  assign n2563 = ~decrypt_i_pad & ~n2562 ;
  assign n2564 = n292 & ~n675 ;
  assign n2565 = ~n635 & ~n773 ;
  assign n2566 = ~n2564 & n2565 ;
  assign n2567 = decrypt_i_pad & ~n2566 ;
  assign n2568 = ~n2563 & ~n2567 ;
  assign n2569 = ~n266 & ~n389 ;
  assign n2570 = ~n652 & ~n2569 ;
  assign n2571 = ~decrypt_i_pad & ~n2570 ;
  assign n2572 = n292 & ~n524 ;
  assign n2573 = ~n381 & ~n1112 ;
  assign n2574 = ~n2572 & n2573 ;
  assign n2575 = decrypt_i_pad & ~n2574 ;
  assign n2576 = ~n2571 & ~n2575 ;
  assign n2577 = ~n266 & ~n368 ;
  assign n2578 = ~n689 & ~n2577 ;
  assign n2579 = ~decrypt_i_pad & ~n2578 ;
  assign n2580 = n292 & ~n464 ;
  assign n2581 = ~n360 & ~n1285 ;
  assign n2582 = ~n2580 & n2581 ;
  assign n2583 = decrypt_i_pad & ~n2582 ;
  assign n2584 = ~n2579 & ~n2583 ;
  assign n2585 = ~n726 & ~n950 ;
  assign n2586 = ~n762 & n2585 ;
  assign n2587 = ~decrypt_i_pad & ~n2586 ;
  assign n2588 = n292 & ~n612 ;
  assign n2589 = ~n576 & ~n1034 ;
  assign n2590 = ~n2588 & n2589 ;
  assign n2591 = decrypt_i_pad & ~n2590 ;
  assign n2592 = ~n2587 & ~n2591 ;
  assign n2593 = ~n540 & ~n1026 ;
  assign n2594 = ~n1351 & n2593 ;
  assign n2595 = ~decrypt_i_pad & ~n2594 ;
  assign n2596 = ~n545 & ~n789 ;
  assign n2597 = ~n1055 & n2596 ;
  assign n2598 = decrypt_i_pad & ~n2597 ;
  assign n2599 = ~n2595 & ~n2598 ;
  assign n2600 = ~n266 & ~n605 ;
  assign n2601 = n266 & ~n733 ;
  assign n2602 = ~n2600 & ~n2601 ;
  assign n2603 = ~decrypt_i_pad & ~n2602 ;
  assign n2604 = n292 & ~n742 ;
  assign n2605 = ~n1339 & ~n1539 ;
  assign n2606 = ~n2604 & n2605 ;
  assign n2607 = decrypt_i_pad & ~n2606 ;
  assign n2608 = ~n2603 & ~n2607 ;
  assign n2609 = ~n465 & ~n485 ;
  assign n2610 = ~n510 & n2609 ;
  assign n2611 = ~decrypt_i_pad & ~n2610 ;
  assign n2612 = n292 & ~n516 ;
  assign n2613 = ~n479 & ~n2601 ;
  assign n2614 = ~n2612 & n2613 ;
  assign n2615 = decrypt_i_pad & ~n2614 ;
  assign n2616 = ~n2611 & ~n2615 ;
  assign n2617 = ~n266 & ~n1213 ;
  assign n2618 = ~n767 & ~n2617 ;
  assign n2619 = ~decrypt_i_pad & ~n2618 ;
  assign n2620 = ~n390 & ~n657 ;
  assign n2621 = ~n811 & n2620 ;
  assign n2622 = decrypt_i_pad & ~n2621 ;
  assign n2623 = ~n2619 & ~n2622 ;
  assign n2624 = \data_ready_reg/NET0131  & \stage1_iter_reg[0]/NET0131  ;
  assign n2625 = ~load_i_pad & ~n2624 ;
  assign n2626 = n250 & ~n2625 ;
  assign n2627 = ~\stage1_iter_reg[0]/NET0131  & ~n250 ;
  assign n2628 = ~n263 & n2627 ;
  assign n2629 = ~n2626 & ~n2628 ;
  assign n2630 = ~\stage1_iter_reg[3]/NET0131  & ~n262 ;
  assign n2631 = ~n263 & ~n2630 ;
  assign n2632 = ~\stage1_iter_reg[2]/NET0131  & ~n254 ;
  assign n2633 = ~n262 & ~n2632 ;
  assign n2634 = ~\data_ready_reg/NET0131  & ~n250 ;
  assign n2635 = ~n281 & ~n2634 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g10087/_0_  = n252 ;
  assign \g10220/_1_  = n255 ;
  assign \g11117/_0_  = ~n297 ;
  assign \g11124/_0_  = ~n300 ;
  assign \g11125/_0_  = ~n335 ;
  assign \g11170/_0_  = ~n373 ;
  assign \g11182/_0_  = ~n376 ;
  assign \g11184/_0_  = ~n411 ;
  assign \g11378/_0_  = ~n427 ;
  assign \g11393/_0_  = ~n452 ;
  assign \g11415/_0_  = ~n470 ;
  assign \g11432/_0_  = ~n489 ;
  assign \g11433/_0_  = ~n492 ;
  assign \g11453/_0_  = ~n506 ;
  assign \g11500/_0_  = ~n522 ;
  assign \g11588/_0_  = ~n534 ;
  assign \g11607/_0_  = ~n551 ;
  assign \g11616/_0_  = ~n585 ;
  assign \g11625/_0_  = ~n588 ;
  assign \g11641_dup/_0_  = ~n610 ;
  assign \g11648/_0_  = ~n628 ;
  assign \g11655/_0_  = ~n663 ;
  assign \g11683/_0_  = ~n666 ;
  assign \g11689/_2_  = ~n669 ;
  assign \g11694/_0_  = ~n685 ;
  assign \g11748/_0_  = ~n688 ;
  assign \g11880/_0_  = ~n709 ;
  assign \g11962/_1_  = n731 ;
  assign \g12016/_0_  = ~n748 ;
  assign \g12038/_0_  = ~n751 ;
  assign \g12039/_0_  = ~n766 ;
  assign \g12094/_0_  = ~n889 ;
  assign \g12100/_0_  = ~n777 ;
  assign \g12132/_0_  = ~n1022 ;
  assign \g12151/_0_  = ~n1032 ;
  assign \g12251/_0_  = ~n1041 ;
  assign \g12279/_0_  = ~n1049 ;
  assign \g12288/_0_  = ~n984 ;
  assign \g12290/_0_  = ~n1060 ;
  assign \g12311/_0_  = ~n1063 ;
  assign \g12313/_0_  = ~n1070 ;
  assign \g12356/_0_  = ~n1079 ;
  assign \g12357/_0_  = ~n1082 ;
  assign \g12427/_0_  = n1196 ;
  assign \g12441/_0_  = ~n1199 ;
  assign \g12442/_0_  = ~n1209 ;
  assign \g12480/_0_  = ~n1092 ;
  assign \g12485/_0_  = ~n1095 ;
  assign \g12506/_0_  = ~n892 ;
  assign \g12544/_0_  = ~n1218 ;
  assign \g12549/_2_  = ~n1225 ;
  assign \g12614/_0_  = n1338 ;
  assign \g12678/_0_  = ~n1123 ;
  assign \g12680/_0_  = ~n1120 ;
  assign \g12748/_0_  = ~n1347 ;
  assign \g15/_0_  = ~n1355 ;
  assign \g25/_0_  = ~n1294 ;
  assign \g31/_0_  = n1405 ;
  assign \g6843/_0_  = n1494 ;
  assign \g6861/_0_  = n1532 ;
  assign \g6863/_0_  = n1615 ;
  assign \g6865/_0_  = ~n1693 ;
  assign \g6887/_0_  = n1744 ;
  assign \g6888/_0_  = n1781 ;
  assign \g6889/_0_  = n1816 ;
  assign \g6890/_0_  = n1851 ;
  assign \g6891/_0_  = n1953 ;
  assign \g6892/_0_  = ~n1992 ;
  assign \g6893/_0_  = ~n2034 ;
  assign \g6894/_0_  = ~n2069 ;
  assign \g6922/_0_  = n2105 ;
  assign \g6923/_0_  = n2146 ;
  assign \g6924/_3_  = n2173 ;
  assign \g6926/_0_  = n2205 ;
  assign \g6927/_0_  = n2242 ;
  assign \g6928/_0_  = n2274 ;
  assign \g6931/_0_  = n2311 ;
  assign \g6933/_0_  = n2344 ;
  assign \g6967/_0_  = n2371 ;
  assign \g6968/_0_  = n2402 ;
  assign \g6969/_0_  = ~n2430 ;
  assign \g6974/_0_  = ~n2455 ;
  assign \g6975/_0_  = n2494 ;
  assign \g6976/_3_  = ~n2531 ;
  assign \g7006/_3_  = n2560 ;
  assign \g8882/_0_  = ~n1859 ;
  assign \g8883/_0_  = ~n2568 ;
  assign \g8884/_0_  = ~n2576 ;
  assign \g8895/_0_  = ~n856 ;
  assign \g8896/_0_  = ~n2584 ;
  assign \g8898/_0_  = ~n793 ;
  assign \g8900/_2_  = ~n981 ;
  assign \g8902/_0_  = ~n2592 ;
  assign \g8907/_0_  = ~n1251 ;
  assign \g8911/_0_  = ~n2599 ;
  assign \g8924/_0_  = ~n2608 ;
  assign \g8927/_0_  = ~n1547 ;
  assign \g8929/_2_  = ~n1413 ;
  assign \g8967/_0_  = ~n955 ;
  assign \g8969/_0_  = ~n1880 ;
  assign \g8973/_2_  = ~n816 ;
  assign \g8987/_0_  = ~n1233 ;
  assign \g8989/_0_  = ~n2616 ;
  assign \g8991/_0_  = ~n930 ;
  assign \g8996/_0_  = ~n2623 ;
  assign \g9099/_0_  = ~n2629 ;
  assign \g9543/_1_  = n2631 ;
  assign \g9751/_1_  = n2633 ;
  assign \g9755/_0_  = n2635 ;
  assign \g9786/_0_  = ~n1437 ;
  assign \g9794/_0_  = ~n933 ;
  assign \g9817/_0_  = ~n1266 ;
  assign \g9836/_0_  = ~n1155 ;
  assign \g9859/_0_  = ~n905 ;
  assign \g9862/_0_  = ~n819 ;
  assign \g9867/_0_  = ~n1429 ;
  assign \g9869/_0_  = ~n1883 ;
  assign \g9876/_0_  = ~n1297 ;
  assign \g9887/_0_  = ~n796 ;
  assign \g9895/_0_  = ~n859 ;
  assign \g9897/_0_  = ~n780 ;
  assign \g9908/_0_  = ~n1236 ;
  assign \g9910/_0_  = ~n1632 ;
  assign \g9915/_0_  = ~n1254 ;
  assign \g9938/_0_  = ~n898 ;
  assign \g9970/_0_  = ~n1862 ;
endmodule
