module top( \a0_pad  , a_pad , b_pad , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , \f0_pad  , f_pad , \g0_pad  , g_pad , \h0_pad  , h_pad , \i0_pad  , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \j0_pad  , \k0_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input b_pad ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \j0_pad  ;
  output \k0_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  wire n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 ;
  assign n35 = c_pad & d_pad ;
  assign n36 = ~c_pad & ~d_pad ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = \i0_pad  & ~n37 ;
  assign n39 = \h0_pad  & n37 ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = e_pad & ~h_pad ;
  assign n42 = ~e_pad & h_pad ;
  assign n43 = ~n41 & ~n42 ;
  assign n48 = ~c_pad & g_pad ;
  assign n49 = ~d_pad & f_pad ;
  assign n50 = n48 & ~n49 ;
  assign n51 = ~n48 & n49 ;
  assign n52 = ~n50 & ~n51 ;
  assign n54 = ~n43 & n52 ;
  assign n53 = n43 & ~n52 ;
  assign n55 = ~b_pad & ~n53 ;
  assign n56 = ~n54 & n55 ;
  assign n45 = ~n37 & n43 ;
  assign n44 = n37 & ~n43 ;
  assign n46 = b_pad & ~n44 ;
  assign n47 = ~n45 & n46 ;
  assign n57 = i_pad & ~j_pad ;
  assign n58 = ~n47 & n57 ;
  assign n59 = ~n56 & n58 ;
  assign n60 = ~q_pad & ~v_pad ;
  assign n61 = ~p_pad & ~u_pad ;
  assign n65 = ~n60 & ~n61 ;
  assign n64 = ~s_pad & ~x_pad ;
  assign n62 = ~r_pad & ~w_pad ;
  assign n63 = ~t_pad & ~y_pad ;
  assign n66 = ~n62 & ~n63 ;
  assign n67 = ~n64 & n66 ;
  assign n68 = n65 & n67 ;
  assign n69 = ~\a0_pad  & b_pad ;
  assign n70 = z_pad & n69 ;
  assign n71 = ~n35 & n70 ;
  assign n72 = ~n68 & n71 ;
  assign n73 = ~\c0_pad  & n72 ;
  assign n74 = ~\c0_pad  & ~\d0_pad  ;
  assign n75 = \c0_pad  & \d0_pad  ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = n72 & n76 ;
  assign n78 = \e0_pad  & n75 ;
  assign n79 = ~\e0_pad  & ~n75 ;
  assign n80 = ~n78 & ~n79 ;
  assign n81 = n72 & n80 ;
  assign n82 = ~\f0_pad  & ~n78 ;
  assign n83 = \f0_pad  & n78 ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = n72 & n84 ;
  assign n86 = \g0_pad  & ~n78 ;
  assign n87 = ~\f0_pad  & ~\g0_pad  ;
  assign n88 = \f0_pad  & \g0_pad  ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = n78 & n89 ;
  assign n91 = ~n86 & ~n90 ;
  assign n92 = n72 & n91 ;
  assign n99 = s_pad & t_pad ;
  assign n100 = r_pad & n99 ;
  assign n129 = ~l_pad & n100 ;
  assign n130 = ~q_pad & ~n129 ;
  assign n131 = ~m_pad & n99 ;
  assign n132 = ~n_pad & t_pad ;
  assign n108 = o_pad & ~t_pad ;
  assign n133 = s_pad & ~n108 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = r_pad & ~n134 ;
  assign n136 = ~n131 & ~n135 ;
  assign n137 = ~n130 & ~n136 ;
  assign n138 = p_pad & ~n137 ;
  assign n106 = q_pad & r_pad ;
  assign n139 = ~p_pad & n99 ;
  assign n140 = n106 & n139 ;
  assign n141 = ~n138 & ~n140 ;
  assign n124 = ~s_pad & ~t_pad ;
  assign n125 = ~r_pad & ~n99 ;
  assign n126 = ~n124 & ~n125 ;
  assign n127 = q_pad & n126 ;
  assign n128 = ~n100 & ~n127 ;
  assign n93 = \e0_pad  & ~n74 ;
  assign n94 = ~\f0_pad  & ~n93 ;
  assign n95 = \f0_pad  & n93 ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = \g0_pad  & n96 ;
  assign n142 = ~k_pad & n99 ;
  assign n143 = n106 & n142 ;
  assign n144 = \h0_pad  & ~n143 ;
  assign n145 = n97 & n144 ;
  assign n146 = ~n128 & n145 ;
  assign n147 = ~n141 & n146 ;
  assign n111 = n_pad & r_pad ;
  assign n112 = ~s_pad & n111 ;
  assign n113 = m_pad & ~r_pad ;
  assign n114 = s_pad & n113 ;
  assign n115 = ~n112 & ~n114 ;
  assign n116 = p_pad & q_pad ;
  assign n117 = t_pad & n116 ;
  assign n118 = ~n115 & n117 ;
  assign n101 = k_pad & ~p_pad ;
  assign n102 = l_pad & ~q_pad ;
  assign n103 = ~n101 & ~n102 ;
  assign n98 = ~p_pad & ~q_pad ;
  assign n104 = ~n98 & n100 ;
  assign n105 = ~n103 & n104 ;
  assign n107 = s_pad & n106 ;
  assign n109 = p_pad & n108 ;
  assign n110 = n107 & n109 ;
  assign n119 = ~n105 & ~n110 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = n97 & ~n120 ;
  assign n122 = ~\h0_pad  & ~n121 ;
  assign n123 = ~\a0_pad  & a_pad ;
  assign n148 = ~n122 & n123 ;
  assign n149 = ~n147 & n148 ;
  assign n150 = q_pad & ~n136 ;
  assign n151 = n88 & n93 ;
  assign n152 = ~n129 & n151 ;
  assign n153 = ~n128 & n152 ;
  assign n154 = ~n150 & n153 ;
  assign n155 = q_pad & ~n131 ;
  assign n156 = n126 & n155 ;
  assign n157 = ~n135 & n156 ;
  assign n158 = n100 & n102 ;
  assign n159 = ~n157 & ~n158 ;
  assign n160 = n87 & ~n93 ;
  assign n161 = ~n159 & n160 ;
  assign n162 = ~n154 & ~n161 ;
  assign n163 = p_pad & ~n162 ;
  assign n164 = ~n89 & ~n96 ;
  assign n165 = t_pad & n101 ;
  assign n166 = n107 & n165 ;
  assign n167 = n164 & n166 ;
  assign n168 = ~\i0_pad  & ~n167 ;
  assign n169 = ~n163 & n168 ;
  assign n170 = \i0_pad  & ~n143 ;
  assign n171 = ~n128 & n170 ;
  assign n172 = n164 & n171 ;
  assign n173 = ~n141 & n172 ;
  assign n174 = n123 & ~n173 ;
  assign n175 = ~n169 & n174 ;
  assign \j0_pad  = ~\h0_pad  ;
  assign \k0_pad  = n40 ;
  assign \l0_pad  = n59 ;
  assign \m0_pad  = n73 ;
  assign \n0_pad  = n77 ;
  assign \o0_pad  = n81 ;
  assign \p0_pad  = n85 ;
  assign \q0_pad  = ~n92 ;
  assign \r0_pad  = n149 ;
  assign \s0_pad  = n175 ;
endmodule
