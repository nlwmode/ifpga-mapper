module top( \C_0_pad  , \C_1_pad  , \C_2_pad  , \C_3_pad  , \C_4_pad  , \C_5_pad  , \C_6_pad  , \C_7_pad  , \C_8_pad  , \P_0_pad  , \X_1_reg/NET0131  , \X_2_reg/NET0131  , \X_3_reg/NET0131  , \X_4_reg/NET0131  , \X_5_reg/NET0131  , \X_6_reg/NET0131  , \X_7_reg/NET0131  , \X_8_reg/NET0131  , \X_8_reg/P0001  , Z_pad , \_al_n0  , \_al_n1  , \g320/_0_  , \g322/_1_  , \g329/_0_  , \g334/_0_  , \g342/_0_  , \g347/_0_  , \g353/_0_  , \g362/_0_  );
  input \C_0_pad  ;
  input \C_1_pad  ;
  input \C_2_pad  ;
  input \C_3_pad  ;
  input \C_4_pad  ;
  input \C_5_pad  ;
  input \C_6_pad  ;
  input \C_7_pad  ;
  input \C_8_pad  ;
  input \P_0_pad  ;
  input \X_1_reg/NET0131  ;
  input \X_2_reg/NET0131  ;
  input \X_3_reg/NET0131  ;
  input \X_4_reg/NET0131  ;
  input \X_5_reg/NET0131  ;
  input \X_6_reg/NET0131  ;
  input \X_7_reg/NET0131  ;
  input \X_8_reg/NET0131  ;
  output \X_8_reg/P0001  ;
  output Z_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g320/_0_  ;
  output \g322/_1_  ;
  output \g329/_0_  ;
  output \g334/_0_  ;
  output \g342/_0_  ;
  output \g347/_0_  ;
  output \g353/_0_  ;
  output \g362/_0_  ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 ;
  assign n19 = ~\X_1_reg/NET0131  & ~\X_2_reg/NET0131  ;
  assign n20 = ~\X_3_reg/NET0131  & ~\X_4_reg/NET0131  ;
  assign n21 = n19 & n20 ;
  assign n22 = \C_5_pad  & \X_5_reg/NET0131  ;
  assign n23 = n21 & n22 ;
  assign n24 = ~\C_0_pad  & ~n23 ;
  assign n25 = \P_0_pad  & ~n24 ;
  assign n42 = \C_3_pad  & \X_3_reg/NET0131  ;
  assign n43 = \C_4_pad  & ~\X_3_reg/NET0131  ;
  assign n44 = \X_4_reg/NET0131  & n43 ;
  assign n45 = ~n42 & ~n44 ;
  assign n39 = \P_0_pad  & ~\X_1_reg/NET0131  ;
  assign n46 = ~\X_2_reg/NET0131  & n39 ;
  assign n47 = ~n45 & n46 ;
  assign n27 = \C_7_pad  & \X_7_reg/NET0131  ;
  assign n28 = \C_8_pad  & ~\X_7_reg/NET0131  ;
  assign n29 = \X_8_reg/NET0131  & n28 ;
  assign n30 = ~n27 & ~n29 ;
  assign n26 = \P_0_pad  & ~\X_5_reg/NET0131  ;
  assign n31 = ~\X_6_reg/NET0131  & n26 ;
  assign n32 = n21 & n31 ;
  assign n33 = ~n30 & n32 ;
  assign n34 = \C_6_pad  & \X_6_reg/NET0131  ;
  assign n35 = n26 & n34 ;
  assign n36 = n21 & n35 ;
  assign n37 = \P_0_pad  & \X_1_reg/NET0131  ;
  assign n38 = \C_1_pad  & n37 ;
  assign n40 = \C_2_pad  & \X_2_reg/NET0131  ;
  assign n41 = n39 & n40 ;
  assign n48 = ~n38 & ~n41 ;
  assign n49 = ~n36 & n48 ;
  assign n50 = ~n33 & n49 ;
  assign n51 = ~n47 & n50 ;
  assign n52 = ~n25 & n51 ;
  assign n53 = \X_2_reg/NET0131  & n37 ;
  assign n54 = \X_3_reg/NET0131  & n53 ;
  assign n55 = \X_4_reg/NET0131  & n54 ;
  assign n56 = \X_5_reg/NET0131  & \X_6_reg/NET0131  ;
  assign n57 = n55 & n56 ;
  assign n58 = \X_7_reg/NET0131  & n57 ;
  assign n59 = ~\X_7_reg/NET0131  & ~n57 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = \X_5_reg/NET0131  & n55 ;
  assign n62 = ~\X_6_reg/NET0131  & ~n61 ;
  assign n63 = ~n57 & ~n62 ;
  assign n64 = ~\X_4_reg/NET0131  & ~n54 ;
  assign n65 = ~n55 & ~n64 ;
  assign n66 = ~\X_5_reg/NET0131  & ~n55 ;
  assign n67 = ~n61 & ~n66 ;
  assign n68 = ~\X_3_reg/NET0131  & ~n53 ;
  assign n69 = ~n54 & ~n68 ;
  assign n70 = ~\X_2_reg/NET0131  & ~n37 ;
  assign n71 = ~n53 & ~n70 ;
  assign n72 = ~\P_0_pad  & \X_1_reg/NET0131  ;
  assign n73 = ~n39 & ~n72 ;
  assign \X_8_reg/P0001  = ~\X_8_reg/NET0131  ;
  assign Z_pad = ~n52 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g320/_0_  = n60 ;
  assign \g322/_1_  = n58 ;
  assign \g329/_0_  = n63 ;
  assign \g334/_0_  = n65 ;
  assign \g342/_0_  = n67 ;
  assign \g347/_0_  = n69 ;
  assign \g353/_0_  = n71 ;
  assign \g362/_0_  = ~n73 ;
endmodule
