module top (\cont_reg[0]/NET0131 , \cont_reg[1]/NET0131 , \cont_reg[2]/NET0131 , \cont_reg[3]/NET0131 , \cont_reg[4]/NET0131 , \cont_reg[5]/NET0131 , \cont_reg[6]/NET0131 , \cont_reg[7]/NET0131 , \mar_reg[0]/NET0131 , \mar_reg[1]/NET0131 , \mar_reg[2]/NET0131 , \mar_reg[3]/NET0131 , \punti_retta[3]_pad , \punti_retta[4]_pad , \punti_retta[6]_pad , \punti_retta[7]_pad , \punti_retta_reg[0]/NET0131 , \punti_retta_reg[1]/NET0131 , \punti_retta_reg[2]/NET0131 , \punti_retta_reg[5]/NET0131 , start_pad, \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , \stato_reg[2]/NET0131 , \t_reg[1]/NET0131 , \t_reg[2]/NET0131 , \t_reg[3]/NET0131 , \t_reg[4]/NET0131 , \t_reg[5]/NET0131 , \t_reg[6]/NET0131 , \x_reg[0]/NET0131 , \x_reg[1]/NET0131 , \x_reg[2]/NET0131 , \x_reg[3]/NET0131 , \x_reg[4]/NET0131 , \x_reg[5]/NET0131 , \x_reg[6]/NET0131 , \x_reg[7]/NET0131 , \y_reg[0]/NET0131 , \y_reg[1]/NET0131 , \y_reg[2]/NET0131 , \y_reg[3]/NET0131 , \_al_n0 , \_al_n1 , \g2119/_0_ , \g2123/_0_ , \g2129/_0_ , \g2133/_0_ , \g2136/_0_ , \g2140/_0_ , \g2141/_0_ , \g2151/_0_ , \g2152/_0_ , \g2166/_0_ , \g2167/_0_ , \g2180/_0_ , \g2181/_0_ , \g2199/_0_ , \g2225/_0_ , \g2227/_0_ , \g2242/_0_ , \g2243/_0_ , \g2272/_0_ , \g2273/_0_ , \g2274/_0_ , \g2275/_0_ , \g2284/_0_ , \g2289/_0_ , \g2303/_0_ , \g2304/_0_ , \g2308/_0_ , \g2309/_0_ , \g2310/_0_ , \g2311/_0_ , \g2312/_0_ , \g2346/_0_ , \g2973/_0_ , \g2984/_0_ , \g3052/_0_ , \g3176/_0_ , \g3277/_0_ , \g3306/_0_ , \g3366/_0_ , \g3371/_0_ , \g3398/_0_ );
	input \cont_reg[0]/NET0131  ;
	input \cont_reg[1]/NET0131  ;
	input \cont_reg[2]/NET0131  ;
	input \cont_reg[3]/NET0131  ;
	input \cont_reg[4]/NET0131  ;
	input \cont_reg[5]/NET0131  ;
	input \cont_reg[6]/NET0131  ;
	input \cont_reg[7]/NET0131  ;
	input \mar_reg[0]/NET0131  ;
	input \mar_reg[1]/NET0131  ;
	input \mar_reg[2]/NET0131  ;
	input \mar_reg[3]/NET0131  ;
	input \punti_retta[3]_pad  ;
	input \punti_retta[4]_pad  ;
	input \punti_retta[6]_pad  ;
	input \punti_retta[7]_pad  ;
	input \punti_retta_reg[0]/NET0131  ;
	input \punti_retta_reg[1]/NET0131  ;
	input \punti_retta_reg[2]/NET0131  ;
	input \punti_retta_reg[5]/NET0131  ;
	input start_pad ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	input \stato_reg[2]/NET0131  ;
	input \t_reg[1]/NET0131  ;
	input \t_reg[2]/NET0131  ;
	input \t_reg[3]/NET0131  ;
	input \t_reg[4]/NET0131  ;
	input \t_reg[5]/NET0131  ;
	input \t_reg[6]/NET0131  ;
	input \x_reg[0]/NET0131  ;
	input \x_reg[1]/NET0131  ;
	input \x_reg[2]/NET0131  ;
	input \x_reg[3]/NET0131  ;
	input \x_reg[4]/NET0131  ;
	input \x_reg[5]/NET0131  ;
	input \x_reg[6]/NET0131  ;
	input \x_reg[7]/NET0131  ;
	input \y_reg[0]/NET0131  ;
	input \y_reg[1]/NET0131  ;
	input \y_reg[2]/NET0131  ;
	input \y_reg[3]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g2119/_0_  ;
	output \g2123/_0_  ;
	output \g2129/_0_  ;
	output \g2133/_0_  ;
	output \g2136/_0_  ;
	output \g2140/_0_  ;
	output \g2141/_0_  ;
	output \g2151/_0_  ;
	output \g2152/_0_  ;
	output \g2166/_0_  ;
	output \g2167/_0_  ;
	output \g2180/_0_  ;
	output \g2181/_0_  ;
	output \g2199/_0_  ;
	output \g2225/_0_  ;
	output \g2227/_0_  ;
	output \g2242/_0_  ;
	output \g2243/_0_  ;
	output \g2272/_0_  ;
	output \g2273/_0_  ;
	output \g2274/_0_  ;
	output \g2275/_0_  ;
	output \g2284/_0_  ;
	output \g2289/_0_  ;
	output \g2303/_0_  ;
	output \g2304/_0_  ;
	output \g2308/_0_  ;
	output \g2309/_0_  ;
	output \g2310/_0_  ;
	output \g2311/_0_  ;
	output \g2312/_0_  ;
	output \g2346/_0_  ;
	output \g2973/_0_  ;
	output \g2984/_0_  ;
	output \g3052/_0_  ;
	output \g3176/_0_  ;
	output \g3277/_0_  ;
	output \g3306/_0_  ;
	output \g3366/_0_  ;
	output \g3371/_0_  ;
	output \g3398/_0_  ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\stato_reg[2]/NET0131 ,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\x_reg[0]/NET0131 ,
		\x_reg[1]/NET0131 ,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\x_reg[2]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\x_reg[4]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\x_reg[6]/NET0131 ,
		\x_reg[7]/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w45_,
		_w46_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\cont_reg[2]/NET0131 ,
		\cont_reg[3]/NET0131 ,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w51_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\cont_reg[4]/NET0131 ,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\cont_reg[5]/NET0131 ,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\mar_reg[2]/NET0131 ,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\mar_reg[3]/NET0131 ,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		_w57_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w44_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		\cont_reg[6]/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		_w44_,
		_w61_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\stato_reg[0]/NET0131 ,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		start_pad,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w66_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w67_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\cont_reg[6]/NET0131 ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		_w64_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w63_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\cont_reg[4]/NET0131 ,
		_w55_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w56_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w60_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\cont_reg[4]/NET0131 ,
		_w60_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w44_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w76_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		\cont_reg[4]/NET0131 ,
		_w70_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\cont_reg[7]/NET0131 ,
		_w70_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\cont_reg[7]/NET0131 ,
		_w60_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\cont_reg[5]/NET0131 ,
		\cont_reg[6]/NET0131 ,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w56_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\cont_reg[7]/NET0131 ,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\cont_reg[7]/NET0131 ,
		_w85_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w60_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		_w44_,
		_w83_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w82_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		start_pad,
		_w66_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w69_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		start_pad,
		_w60_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		_w44_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		_w94_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\punti_retta[6]_pad ,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\cont_reg[6]/NET0131 ,
		_w57_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w44_,
		_w95_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w85_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w99_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w98_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\cont_reg[3]/NET0131 ,
		_w70_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\cont_reg[3]/NET0131 ,
		_w60_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\cont_reg[0]/NET0131 ,
		_w51_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\cont_reg[1]/NET0131 ,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\cont_reg[2]/NET0131 ,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\cont_reg[3]/NET0131 ,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w55_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w60_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w44_,
		_w105_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w111_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w104_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\punti_retta_reg[2]/NET0131 ,
		_w94_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\punti_retta_reg[2]/NET0131 ,
		_w60_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\punti_retta_reg[2]/NET0131 ,
		start_pad,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\cont_reg[2]/NET0131 ,
		_w107_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w108_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		start_pad,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		_w60_,
		_w117_,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		_w44_,
		_w116_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w115_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\punti_retta_reg[5]/NET0131 ,
		_w60_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\punti_retta_reg[5]/NET0131 ,
		start_pad,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		\cont_reg[5]/NET0131 ,
		_w56_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w57_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		start_pad,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w60_,
		_w127_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		_w44_,
		_w126_,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\punti_retta_reg[5]/NET0131 ,
		_w94_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w134_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		\cont_reg[0]/NET0131 ,
		_w51_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w106_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		_w95_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		_w44_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w94_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\punti_retta_reg[0]/NET0131 ,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w95_,
		_w140_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\punti_retta_reg[1]/NET0131 ,
		_w97_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\cont_reg[1]/NET0131 ,
		_w106_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		_w100_,
		_w107_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		_w146_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w145_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w60_,
		_w129_,
		_w150_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		\cont_reg[5]/NET0131 ,
		_w60_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		_w44_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w150_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		\cont_reg[5]/NET0131 ,
		_w70_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w60_,
		_w119_,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		\cont_reg[2]/NET0131 ,
		_w60_,
		_w157_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		_w44_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w156_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\cont_reg[2]/NET0131 ,
		_w70_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		_w60_,
		_w106_,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		_w44_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		_w70_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\cont_reg[1]/NET0131 ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\cont_reg[1]/NET0131 ,
		_w44_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w162_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w165_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w60_,
		_w138_,
		_w169_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\cont_reg[0]/NET0131 ,
		_w60_,
		_w170_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		_w44_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w169_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\cont_reg[0]/NET0131 ,
		_w70_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w172_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\stato_reg[0]/NET0131 ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w60_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w44_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		_w59_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\mar_reg[3]/NET0131 ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		_w181_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		_w67_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w178_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w180_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w44_,
		_w176_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\mar_reg[0]/NET0131 ,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w44_,
		_w60_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\mar_reg[0]/NET0131 ,
		_w184_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w188_,
		_w189_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w190_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		\stato_reg[0]/NET0131 ,
		_w181_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\t_reg[1]/NET0131 ,
		\x_reg[1]/NET0131 ,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\t_reg[1]/NET0131 ,
		\x_reg[1]/NET0131 ,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w193_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		\stato_reg[0]/NET0131 ,
		_w175_,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\mar_reg[3]/NET0131 ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		\mar_reg[0]/NET0131 ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\mar_reg[2]/NET0131 ,
		\mar_reg[3]/NET0131 ,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name160 (
		\mar_reg[1]/NET0131 ,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		\mar_reg[0]/NET0131 ,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w201_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		_w198_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w65_,
		_w187_,
		_w207_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		\x_reg[1]/NET0131 ,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\stato_reg[0]/NET0131 ,
		_w181_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\x_reg[0]/NET0131 ,
		\y_reg[0]/NET0131 ,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\x_reg[1]/NET0131 ,
		\y_reg[1]/NET0131 ,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		\x_reg[1]/NET0131 ,
		\y_reg[1]/NET0131 ,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w211_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w210_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w210_,
		_w213_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		_w209_,
		_w214_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w197_,
		_w206_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w208_,
		_w217_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w218_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w58_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		_w187_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\mar_reg[1]/NET0131 ,
		_w184_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w189_,
		_w223_,
		_w225_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		\mar_reg[2]/NET0131 ,
		_w58_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w59_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		_w187_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		\mar_reg[2]/NET0131 ,
		_w184_,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w189_,
		_w229_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		\mar_reg[3]/NET0131 ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w200_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		_w198_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		_w193_,
		_w207_,
		_w237_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		\x_reg[0]/NET0131 ,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		\x_reg[0]/NET0131 ,
		\y_reg[0]/NET0131 ,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w210_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w209_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w236_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		_w238_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name201 (
		_w193_,
		_w205_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		\stato_reg[2]/NET0131 ,
		_w43_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		_w209_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		\y_reg[1]/NET0131 ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w244_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		\stato_reg[0]/NET0131 ,
		_w68_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w60_,
		_w68_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w65_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		start_pad,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w249_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		_w68_,
		_w95_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w198_,
		_w209_,
		_w255_
	);
	LUT2 #(
		.INIT('h4)
	) name213 (
		_w93_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w254_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\x_reg[5]/NET0131 ,
		_w176_,
		_w258_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\stato_reg[1]/NET0131 ,
		_w44_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w198_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		\t_reg[6]/NET0131 ,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w258_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\x_reg[4]/NET0131 ,
		_w176_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\t_reg[5]/NET0131 ,
		_w260_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\mar_reg[0]/NET0131 ,
		_w234_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w200_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		_w193_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		\y_reg[2]/NET0131 ,
		_w246_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w268_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w201_,
		_w266_,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		_w193_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		\y_reg[3]/NET0131 ,
		_w246_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		start_pad,
		_w250_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w176_,
		_w181_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\x_reg[0]/NET0131 ,
		_w176_,
		_w278_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\t_reg[1]/NET0131 ,
		_w260_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\x_reg[1]/NET0131 ,
		_w176_,
		_w281_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		\t_reg[2]/NET0131 ,
		_w260_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		\x_reg[2]/NET0131 ,
		_w176_,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\t_reg[3]/NET0131 ,
		_w260_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		\x_reg[3]/NET0131 ,
		_w176_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\t_reg[4]/NET0131 ,
		_w260_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w193_,
		_w235_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		\y_reg[0]/NET0131 ,
		_w246_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\punti_retta[4]_pad ,
		_w94_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\punti_retta[4]_pad ,
		_w60_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		\punti_retta[4]_pad ,
		start_pad,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		start_pad,
		_w75_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		_w60_,
		_w295_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name255 (
		_w296_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w44_,
		_w294_,
		_w299_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w293_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		\x_reg[6]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		\x_reg[5]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		\x_reg[4]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\x_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		\x_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w210_,
		_w211_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w212_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		_w306_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w305_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\x_reg[3]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w310_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		_w304_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w302_,
		_w303_,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		_w313_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		\x_reg[5]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\x_reg[4]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\x_reg[3]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		\x_reg[6]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w316_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w319_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w315_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		_w209_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		\t_reg[6]/NET0131 ,
		\x_reg[6]/NET0131 ,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\t_reg[5]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		\t_reg[5]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		\t_reg[4]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		\t_reg[2]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		_w194_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\t_reg[2]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		\t_reg[3]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w332_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		\t_reg[3]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		\t_reg[4]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w335_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		_w334_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w328_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w327_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w325_,
		_w326_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		\t_reg[6]/NET0131 ,
		\x_reg[6]/NET0131 ,
		_w343_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		_w193_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w342_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		\x_reg[7]/NET0131 ,
		_w207_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		_w198_,
		_w271_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		_w345_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w324_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		\x_reg[2]/NET0131 ,
		_w207_,
		_w351_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		_w198_,
		_w267_,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w329_,
		_w331_,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w194_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w194_,
		_w353_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name313 (
		_w193_,
		_w354_,
		_w356_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w305_,
		_w306_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w308_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w308_,
		_w358_,
		_w360_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		_w209_,
		_w359_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w360_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w351_,
		_w352_,
		_w363_
	);
	LUT2 #(
		.INIT('h4)
	) name321 (
		_w357_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		_w362_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		\x_reg[3]/NET0131 ,
		_w207_,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w333_,
		_w335_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		_w332_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w332_,
		_w367_,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		_w193_,
		_w368_,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w311_,
		_w318_,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		_w310_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		_w310_,
		_w372_,
		_w374_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		_w209_,
		_w373_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w374_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w347_,
		_w366_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w371_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w376_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w303_,
		_w316_,
		_w380_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		_w313_,
		_w319_,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		_w380_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		_w380_,
		_w381_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		_w209_,
		_w382_,
		_w384_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\x_reg[5]/NET0131 ,
		_w207_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w326_,
		_w327_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w339_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w326_,
		_w340_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		_w193_,
		_w388_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		_w389_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w347_,
		_w386_,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h4)
	) name351 (
		_w385_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		start_pad,
		_w88_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		\punti_retta[7]_pad ,
		start_pad,
		_w396_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		_w60_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w395_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		\punti_retta[7]_pad ,
		_w60_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		_w44_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		_w398_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\punti_retta[7]_pad ,
		_w94_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		\x_reg[6]/NET0131 ,
		_w207_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w325_,
		_w343_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w331_,
		_w335_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name364 (
		_w330_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w333_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w336_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w327_,
		_w328_,
		_w410_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		_w409_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w326_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		_w405_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w405_,
		_w412_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w193_,
		_w413_,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		_w414_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w304_,
		_w311_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w309_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		_w305_,
		_w311_,
		_w419_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		_w319_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		_w304_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w418_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w303_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w316_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w302_,
		_w320_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name384 (
		_w424_,
		_w425_,
		_w427_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		_w209_,
		_w426_,
		_w428_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w427_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w347_,
		_w404_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w416_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		_w429_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		\punti_retta[3]_pad ,
		_w94_,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		start_pad,
		_w110_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\punti_retta[3]_pad ,
		start_pad,
		_w435_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		_w60_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		_w434_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		\punti_retta[3]_pad ,
		_w60_,
		_w438_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w44_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w437_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w433_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		\x_reg[4]/NET0131 ,
		_w207_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w304_,
		_w317_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w312_,
		_w318_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w443_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		_w443_,
		_w444_,
		_w446_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		_w209_,
		_w445_,
		_w447_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w446_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w328_,
		_w336_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w408_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w408_,
		_w449_,
		_w451_
	);
	LUT2 #(
		.INIT('h2)
	) name409 (
		_w193_,
		_w450_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name410 (
		_w451_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w347_,
		_w442_,
		_w454_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w453_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		_w448_,
		_w455_,
		_w456_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g2119/_0_  = _w73_ ;
	assign \g2123/_0_  = _w81_ ;
	assign \g2129/_0_  = _w92_ ;
	assign \g2133/_0_  = _w103_ ;
	assign \g2136/_0_  = _w114_ ;
	assign \g2140/_0_  = _w125_ ;
	assign \g2141/_0_  = _w136_ ;
	assign \g2151/_0_  = _w144_ ;
	assign \g2152/_0_  = _w149_ ;
	assign \g2166/_0_  = _w155_ ;
	assign \g2167/_0_  = _w161_ ;
	assign \g2180/_0_  = _w168_ ;
	assign \g2181/_0_  = _w174_ ;
	assign \g2199/_0_  = _w186_ ;
	assign \g2225/_0_  = _w192_ ;
	assign \g2227/_0_  = _w220_ ;
	assign \g2242/_0_  = _w226_ ;
	assign \g2243/_0_  = _w232_ ;
	assign \g2272/_0_  = _w243_ ;
	assign \g2273/_0_  = _w248_ ;
	assign \g2274/_0_  = _w253_ ;
	assign \g2275/_0_  = _w257_ ;
	assign \g2284/_0_  = _w262_ ;
	assign \g2289/_0_  = _w265_ ;
	assign \g2303/_0_  = _w270_ ;
	assign \g2304/_0_  = _w274_ ;
	assign \g2308/_0_  = _w277_ ;
	assign \g2309/_0_  = _w280_ ;
	assign \g2310/_0_  = _w283_ ;
	assign \g2311/_0_  = _w286_ ;
	assign \g2312/_0_  = _w289_ ;
	assign \g2346/_0_  = _w292_ ;
	assign \g2973/_0_  = _w301_ ;
	assign \g2984/_0_  = _w350_ ;
	assign \g3052/_0_  = _w365_ ;
	assign \g3176/_0_  = _w379_ ;
	assign \g3277/_0_  = _w394_ ;
	assign \g3306/_0_  = _w403_ ;
	assign \g3366/_0_  = _w432_ ;
	assign \g3371/_0_  = _w441_ ;
	assign \g3398/_0_  = _w456_ ;
endmodule;