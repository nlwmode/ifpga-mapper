module top (\v0_pad , \v10_reg/NET0131 , \v11_reg/NET0131 , \v12_reg/NET0131 , \v1_pad , \v2_pad , \v3_pad , \v4_pad , \v5_pad , \v6_pad , \v7_reg/NET0131 , \v8_reg/NET0131 , \v9_reg/NET0131 , \_al_n0 , \_al_n1 , \g528/_2_ , \g534/_0_ , \g535/_0_ , \g537/_0_ , \g560/_3_ , \g722/_0_ , \g754/_0_ , \v13_D_10_pad , \v13_D_11_pad , \v13_D_12_pad , \v13_D_6_pad , \v13_D_7_pad , \v13_D_9_pad );
	input \v0_pad  ;
	input \v10_reg/NET0131  ;
	input \v11_reg/NET0131  ;
	input \v12_reg/NET0131  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input \v5_pad  ;
	input \v6_pad  ;
	input \v7_reg/NET0131  ;
	input \v8_reg/NET0131  ;
	input \v9_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g528/_2_  ;
	output \g534/_0_  ;
	output \g535/_0_  ;
	output \g537/_0_  ;
	output \g560/_3_  ;
	output \g722/_0_  ;
	output \g754/_0_  ;
	output \v13_D_10_pad  ;
	output \v13_D_11_pad  ;
	output \v13_D_12_pad  ;
	output \v13_D_6_pad  ;
	output \v13_D_7_pad  ;
	output \v13_D_9_pad  ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w15_
	);
	LUT4 #(
		.INIT('h0100)
	) name1 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w16_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w17_
	);
	LUT3 #(
		.INIT('h01)
	) name3 (
		\v0_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w18_
	);
	LUT3 #(
		.INIT('hd0)
	) name4 (
		\v10_reg/NET0131 ,
		_w16_,
		_w18_,
		_w19_
	);
	LUT3 #(
		.INIT('h02)
	) name5 (
		\v1_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w20_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w21_
	);
	LUT3 #(
		.INIT('h02)
	) name7 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w22_
	);
	LUT3 #(
		.INIT('ha8)
	) name8 (
		_w20_,
		_w21_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		_w24_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w25_
	);
	LUT4 #(
		.INIT('h0010)
	) name11 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w25_,
		_w26_,
		_w27_
	);
	LUT3 #(
		.INIT('hef)
	) name13 (
		_w19_,
		_w23_,
		_w27_,
		_w28_
	);
	LUT3 #(
		.INIT('h02)
	) name14 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w29_
	);
	LUT4 #(
		.INIT('h0010)
	) name15 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v1_pad ,
		\v5_pad ,
		_w30_
	);
	LUT3 #(
		.INIT('h15)
	) name16 (
		_w26_,
		_w29_,
		_w30_,
		_w31_
	);
	LUT3 #(
		.INIT('ha8)
	) name17 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w32_
	);
	LUT3 #(
		.INIT('ha2)
	) name18 (
		\v0_pad ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w33_
	);
	LUT4 #(
		.INIT('h3331)
	) name19 (
		_w17_,
		_w25_,
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h7)
	) name20 (
		_w31_,
		_w34_,
		_w35_
	);
	LUT4 #(
		.INIT('h0008)
	) name21 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w36_
	);
	LUT3 #(
		.INIT('h10)
	) name22 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w37_
	);
	LUT3 #(
		.INIT('h20)
	) name23 (
		\v3_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w39_
	);
	LUT4 #(
		.INIT('h2000)
	) name25 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w40_
	);
	LUT4 #(
		.INIT('h0015)
	) name26 (
		_w36_,
		_w37_,
		_w38_,
		_w40_,
		_w41_
	);
	LUT4 #(
		.INIT('h0002)
	) name27 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT4 #(
		.INIT('h0100)
	) name29 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v4_pad ,
		\v8_reg/NET0131 ,
		_w44_
	);
	LUT3 #(
		.INIT('h2a)
	) name30 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w45_
	);
	LUT4 #(
		.INIT('h4440)
	) name31 (
		\v12_reg/NET0131 ,
		_w42_,
		_w44_,
		_w45_,
		_w46_
	);
	LUT4 #(
		.INIT('h0001)
	) name32 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w47_
	);
	LUT4 #(
		.INIT('h0008)
	) name33 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT4 #(
		.INIT('h4000)
	) name35 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w50_
	);
	LUT3 #(
		.INIT('h31)
	) name36 (
		\v2_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\v11_reg/NET0131 ,
		\v4_pad ,
		_w52_
	);
	LUT3 #(
		.INIT('h45)
	) name38 (
		_w50_,
		_w51_,
		_w52_,
		_w53_
	);
	LUT4 #(
		.INIT('h0e04)
	) name39 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w54_
	);
	LUT4 #(
		.INIT('h0080)
	) name40 (
		\v11_reg/NET0131 ,
		\v5_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w55_
	);
	LUT4 #(
		.INIT('h0400)
	) name41 (
		\v2_pad ,
		\v3_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w56_
	);
	LUT3 #(
		.INIT('h01)
	) name42 (
		_w54_,
		_w55_,
		_w56_,
		_w57_
	);
	LUT4 #(
		.INIT('hccc8)
	) name43 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		_w42_,
		_w58_,
		_w59_
	);
	LUT3 #(
		.INIT('h70)
	) name45 (
		_w53_,
		_w57_,
		_w59_,
		_w60_
	);
	LUT3 #(
		.INIT('h54)
	) name46 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w44_,
		_w61_
	);
	LUT4 #(
		.INIT('h0010)
	) name47 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w62_
	);
	LUT3 #(
		.INIT('h23)
	) name48 (
		\v5_pad ,
		_w62_,
		_w36_,
		_w63_
	);
	LUT3 #(
		.INIT('h8a)
	) name49 (
		_w42_,
		_w61_,
		_w63_,
		_w64_
	);
	LUT3 #(
		.INIT('h4c)
	) name50 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v5_pad ,
		_w65_
	);
	LUT3 #(
		.INIT('h10)
	) name51 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w66_
	);
	LUT3 #(
		.INIT('h20)
	) name52 (
		_w20_,
		_w65_,
		_w66_,
		_w67_
	);
	LUT4 #(
		.INIT('hfca8)
	) name53 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w68_
	);
	LUT3 #(
		.INIT('ha2)
	) name54 (
		\v9_reg/NET0131 ,
		_w24_,
		_w68_,
		_w69_
	);
	LUT4 #(
		.INIT('h444c)
	) name55 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w70_
	);
	LUT4 #(
		.INIT('h54fe)
	) name56 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v4_pad ,
		\v7_reg/NET0131 ,
		_w71_
	);
	LUT4 #(
		.INIT('hafab)
	) name57 (
		\v10_reg/NET0131 ,
		_w39_,
		_w70_,
		_w71_,
		_w72_
	);
	LUT4 #(
		.INIT('h5f13)
	) name58 (
		_w22_,
		_w24_,
		_w29_,
		_w68_,
		_w73_
	);
	LUT3 #(
		.INIT('h15)
	) name59 (
		_w69_,
		_w72_,
		_w73_,
		_w74_
	);
	LUT4 #(
		.INIT('h4000)
	) name60 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w47_,
		_w75_,
		_w76_
	);
	LUT3 #(
		.INIT('h80)
	) name62 (
		\v5_pad ,
		_w42_,
		_w36_,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\v3_pad ,
		\v8_reg/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name64 (
		\v2_pad ,
		\v3_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\v4_pad ,
		\v7_reg/NET0131 ,
		_w80_
	);
	LUT4 #(
		.INIT('h8880)
	) name66 (
		_w15_,
		_w42_,
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('he)
	) name67 (
		_w77_,
		_w81_,
		_w82_
	);
	LUT3 #(
		.INIT('h08)
	) name68 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w83_
	);
	LUT4 #(
		.INIT('h4440)
	) name69 (
		\v12_reg/NET0131 ,
		_w42_,
		_w44_,
		_w83_,
		_w84_
	);
	LUT3 #(
		.INIT('h08)
	) name70 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w85_
	);
	LUT3 #(
		.INIT('h10)
	) name71 (
		\v10_reg/NET0131 ,
		\v1_pad ,
		\v4_pad ,
		_w86_
	);
	LUT4 #(
		.INIT('h0001)
	) name72 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w87_
	);
	LUT4 #(
		.INIT('hec00)
	) name73 (
		_w78_,
		_w85_,
		_w86_,
		_w87_,
		_w88_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g528/_2_  = _w28_ ;
	assign \g534/_0_  = _w35_ ;
	assign \g535/_0_  = _w43_ ;
	assign \g537/_0_  = _w46_ ;
	assign \g560/_3_  = _w49_ ;
	assign \g722/_0_  = _w60_ ;
	assign \g754/_0_  = _w64_ ;
	assign \v13_D_10_pad  = _w67_ ;
	assign \v13_D_11_pad  = _w74_ ;
	assign \v13_D_12_pad  = _w76_ ;
	assign \v13_D_6_pad  = _w82_ ;
	assign \v13_D_7_pad  = _w84_ ;
	assign \v13_D_9_pad  = _w88_ ;
endmodule;