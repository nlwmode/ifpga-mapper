module top (\pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 , \pi135 , \pi136 , \pi137 , \pi138 , \pi139 , \pi140 , \pi141 , \pi142 , \pi143 , \pi144 , \pi145 , \pi146 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 , \po128 , \po129 , \po130 , \po131 , \po132 , \po133 , \po134 , \po135 , \po136 , \po137 , \po138 , \po139 , \po140 , \po141 );
	input \pi000  ;
	input \pi001  ;
	input \pi002  ;
	input \pi003  ;
	input \pi004  ;
	input \pi005  ;
	input \pi006  ;
	input \pi007  ;
	input \pi008  ;
	input \pi009  ;
	input \pi010  ;
	input \pi011  ;
	input \pi012  ;
	input \pi013  ;
	input \pi014  ;
	input \pi015  ;
	input \pi016  ;
	input \pi017  ;
	input \pi018  ;
	input \pi019  ;
	input \pi020  ;
	input \pi021  ;
	input \pi022  ;
	input \pi023  ;
	input \pi024  ;
	input \pi025  ;
	input \pi026  ;
	input \pi027  ;
	input \pi028  ;
	input \pi029  ;
	input \pi030  ;
	input \pi031  ;
	input \pi032  ;
	input \pi033  ;
	input \pi034  ;
	input \pi035  ;
	input \pi036  ;
	input \pi037  ;
	input \pi038  ;
	input \pi039  ;
	input \pi040  ;
	input \pi041  ;
	input \pi042  ;
	input \pi043  ;
	input \pi044  ;
	input \pi045  ;
	input \pi046  ;
	input \pi047  ;
	input \pi048  ;
	input \pi049  ;
	input \pi050  ;
	input \pi051  ;
	input \pi052  ;
	input \pi053  ;
	input \pi054  ;
	input \pi055  ;
	input \pi056  ;
	input \pi057  ;
	input \pi058  ;
	input \pi059  ;
	input \pi060  ;
	input \pi061  ;
	input \pi062  ;
	input \pi063  ;
	input \pi064  ;
	input \pi065  ;
	input \pi066  ;
	input \pi067  ;
	input \pi068  ;
	input \pi069  ;
	input \pi070  ;
	input \pi071  ;
	input \pi072  ;
	input \pi073  ;
	input \pi074  ;
	input \pi075  ;
	input \pi076  ;
	input \pi077  ;
	input \pi078  ;
	input \pi079  ;
	input \pi080  ;
	input \pi081  ;
	input \pi082  ;
	input \pi083  ;
	input \pi084  ;
	input \pi085  ;
	input \pi086  ;
	input \pi087  ;
	input \pi088  ;
	input \pi089  ;
	input \pi090  ;
	input \pi091  ;
	input \pi092  ;
	input \pi093  ;
	input \pi094  ;
	input \pi095  ;
	input \pi096  ;
	input \pi097  ;
	input \pi098  ;
	input \pi099  ;
	input \pi100  ;
	input \pi101  ;
	input \pi102  ;
	input \pi103  ;
	input \pi104  ;
	input \pi105  ;
	input \pi106  ;
	input \pi107  ;
	input \pi108  ;
	input \pi109  ;
	input \pi110  ;
	input \pi111  ;
	input \pi112  ;
	input \pi113  ;
	input \pi114  ;
	input \pi115  ;
	input \pi116  ;
	input \pi117  ;
	input \pi118  ;
	input \pi119  ;
	input \pi120  ;
	input \pi121  ;
	input \pi122  ;
	input \pi123  ;
	input \pi124  ;
	input \pi125  ;
	input \pi126  ;
	input \pi127  ;
	input \pi128  ;
	input \pi129  ;
	input \pi130  ;
	input \pi131  ;
	input \pi132  ;
	input \pi133  ;
	input \pi134  ;
	input \pi135  ;
	input \pi136  ;
	input \pi137  ;
	input \pi138  ;
	input \pi139  ;
	input \pi140  ;
	input \pi141  ;
	input \pi142  ;
	input \pi143  ;
	input \pi144  ;
	input \pi145  ;
	input \pi146  ;
	output \po000  ;
	output \po001  ;
	output \po002  ;
	output \po003  ;
	output \po004  ;
	output \po005  ;
	output \po006  ;
	output \po007  ;
	output \po008  ;
	output \po009  ;
	output \po010  ;
	output \po011  ;
	output \po012  ;
	output \po013  ;
	output \po014  ;
	output \po015  ;
	output \po016  ;
	output \po017  ;
	output \po018  ;
	output \po019  ;
	output \po020  ;
	output \po021  ;
	output \po022  ;
	output \po023  ;
	output \po024  ;
	output \po025  ;
	output \po026  ;
	output \po027  ;
	output \po028  ;
	output \po029  ;
	output \po030  ;
	output \po031  ;
	output \po032  ;
	output \po033  ;
	output \po034  ;
	output \po035  ;
	output \po036  ;
	output \po037  ;
	output \po038  ;
	output \po039  ;
	output \po040  ;
	output \po041  ;
	output \po042  ;
	output \po043  ;
	output \po044  ;
	output \po045  ;
	output \po046  ;
	output \po047  ;
	output \po048  ;
	output \po049  ;
	output \po050  ;
	output \po051  ;
	output \po052  ;
	output \po053  ;
	output \po054  ;
	output \po055  ;
	output \po056  ;
	output \po057  ;
	output \po058  ;
	output \po059  ;
	output \po060  ;
	output \po061  ;
	output \po062  ;
	output \po063  ;
	output \po064  ;
	output \po065  ;
	output \po066  ;
	output \po067  ;
	output \po068  ;
	output \po069  ;
	output \po070  ;
	output \po071  ;
	output \po072  ;
	output \po073  ;
	output \po074  ;
	output \po075  ;
	output \po076  ;
	output \po077  ;
	output \po078  ;
	output \po079  ;
	output \po080  ;
	output \po081  ;
	output \po082  ;
	output \po083  ;
	output \po084  ;
	output \po085  ;
	output \po086  ;
	output \po087  ;
	output \po088  ;
	output \po089  ;
	output \po090  ;
	output \po091  ;
	output \po092  ;
	output \po093  ;
	output \po094  ;
	output \po095  ;
	output \po096  ;
	output \po097  ;
	output \po098  ;
	output \po099  ;
	output \po100  ;
	output \po101  ;
	output \po102  ;
	output \po103  ;
	output \po104  ;
	output \po105  ;
	output \po106  ;
	output \po107  ;
	output \po108  ;
	output \po109  ;
	output \po110  ;
	output \po111  ;
	output \po112  ;
	output \po113  ;
	output \po114  ;
	output \po115  ;
	output \po116  ;
	output \po117  ;
	output \po118  ;
	output \po119  ;
	output \po120  ;
	output \po121  ;
	output \po122  ;
	output \po123  ;
	output \po124  ;
	output \po125  ;
	output \po126  ;
	output \po127  ;
	output \po128  ;
	output \po129  ;
	output \po130  ;
	output \po131  ;
	output \po132  ;
	output \po133  ;
	output \po134  ;
	output \po135  ;
	output \po136  ;
	output \po137  ;
	output \po138  ;
	output \po139  ;
	output \po140  ;
	output \po141  ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\pi003 ,
		\pi129 ,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\pi000 ,
		\pi054 ,
		_w150_
	);
	LUT3 #(
		.INIT('h01)
	) name2 (
		\pi004 ,
		\pi016 ,
		\pi019 ,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\pi017 ,
		\pi018 ,
		_w152_
	);
	LUT4 #(
		.INIT('h0001)
	) name4 (
		\pi005 ,
		\pi006 ,
		\pi012 ,
		\pi022 ,
		_w153_
	);
	LUT3 #(
		.INIT('h80)
	) name5 (
		_w151_,
		_w152_,
		_w153_,
		_w154_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		\pi007 ,
		\pi013 ,
		\pi014 ,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\pi009 ,
		\pi011 ,
		_w156_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		\pi008 ,
		\pi009 ,
		\pi011 ,
		\pi021 ,
		_w157_
	);
	LUT3 #(
		.INIT('h40)
	) name9 (
		\pi000 ,
		_w155_,
		_w157_,
		_w158_
	);
	LUT3 #(
		.INIT('h10)
	) name10 (
		\pi009 ,
		\pi011 ,
		\pi054 ,
		_w159_
	);
	LUT4 #(
		.INIT('h0010)
	) name11 (
		\pi005 ,
		\pi022 ,
		\pi054 ,
		\pi056 ,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT4 #(
		.INIT('h1500)
	) name13 (
		_w150_,
		_w154_,
		_w158_,
		_w161_,
		_w162_
	);
	LUT4 #(
		.INIT('h0001)
	) name14 (
		\pi007 ,
		\pi008 ,
		\pi013 ,
		\pi021 ,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\pi010 ,
		\pi014 ,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT4 #(
		.INIT('hfce0)
	) name17 (
		\pi007 ,
		\pi008 ,
		\pi013 ,
		\pi021 ,
		_w166_
	);
	LUT4 #(
		.INIT('h0051)
	) name18 (
		\pi010 ,
		\pi014 ,
		_w163_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('h5576)
	) name19 (
		\pi007 ,
		\pi008 ,
		\pi013 ,
		\pi021 ,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		\pi014 ,
		_w168_,
		_w169_
	);
	LUT4 #(
		.INIT('h7757)
	) name21 (
		_w154_,
		_w165_,
		_w167_,
		_w169_,
		_w170_
	);
	LUT3 #(
		.INIT('h0e)
	) name22 (
		\pi005 ,
		\pi022 ,
		\pi056 ,
		_w171_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		_w156_,
		_w171_,
		_w172_
	);
	LUT4 #(
		.INIT('h1500)
	) name24 (
		_w150_,
		_w154_,
		_w158_,
		_w172_,
		_w173_
	);
	LUT4 #(
		.INIT('hfddd)
	) name25 (
		_w149_,
		_w162_,
		_w170_,
		_w173_,
		_w174_
	);
	LUT3 #(
		.INIT('h45)
	) name26 (
		\pi001 ,
		\pi017 ,
		\pi054 ,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\pi010 ,
		\pi022 ,
		_w176_
	);
	LUT3 #(
		.INIT('h01)
	) name28 (
		\pi010 ,
		\pi013 ,
		\pi022 ,
		_w177_
	);
	LUT3 #(
		.INIT('h01)
	) name29 (
		\pi008 ,
		\pi011 ,
		\pi021 ,
		_w178_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\pi014 ,
		\pi018 ,
		_w179_
	);
	LUT3 #(
		.INIT('h80)
	) name31 (
		_w177_,
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\pi005 ,
		\pi006 ,
		_w181_
	);
	LUT4 #(
		.INIT('h0001)
	) name33 (
		\pi005 ,
		\pi006 ,
		\pi007 ,
		\pi012 ,
		_w182_
	);
	LUT3 #(
		.INIT('h40)
	) name34 (
		\pi001 ,
		_w151_,
		_w182_,
		_w183_
	);
	LUT4 #(
		.INIT('ha888)
	) name35 (
		_w149_,
		_w175_,
		_w180_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\pi009 ,
		\pi013 ,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w182_,
		_w185_,
		_w186_
	);
	LUT3 #(
		.INIT('h80)
	) name38 (
		_w151_,
		_w152_,
		_w178_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\pi010 ,
		\pi014 ,
		_w188_
	);
	LUT4 #(
		.INIT('h0100)
	) name40 (
		\pi010 ,
		\pi014 ,
		\pi022 ,
		\pi054 ,
		_w189_
	);
	LUT3 #(
		.INIT('hd0)
	) name41 (
		\pi013 ,
		_w182_,
		_w189_,
		_w190_
	);
	LUT3 #(
		.INIT('h40)
	) name42 (
		_w186_,
		_w187_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\pi013 ,
		_w182_,
		_w192_
	);
	LUT4 #(
		.INIT('hfac8)
	) name44 (
		\pi005 ,
		\pi006 ,
		\pi007 ,
		\pi012 ,
		_w193_
	);
	LUT4 #(
		.INIT('heee0)
	) name45 (
		\pi005 ,
		\pi006 ,
		\pi007 ,
		\pi012 ,
		_w194_
	);
	LUT3 #(
		.INIT('h01)
	) name46 (
		\pi009 ,
		_w193_,
		_w194_,
		_w195_
	);
	LUT3 #(
		.INIT('ha8)
	) name47 (
		_w149_,
		_w192_,
		_w195_,
		_w196_
	);
	LUT3 #(
		.INIT('h15)
	) name48 (
		_w184_,
		_w191_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\pi122 ,
		\pi127 ,
		_w198_
	);
	LUT3 #(
		.INIT('h15)
	) name50 (
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w199_
	);
	LUT4 #(
		.INIT('h0111)
	) name51 (
		\pi065 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\pi042 ,
		\pi044 ,
		_w201_
	);
	LUT4 #(
		.INIT('h0001)
	) name53 (
		\pi038 ,
		\pi040 ,
		\pi042 ,
		\pi044 ,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\pi046 ,
		\pi050 ,
		_w203_
	);
	LUT3 #(
		.INIT('h01)
	) name55 (
		\pi041 ,
		\pi043 ,
		\pi047 ,
		_w204_
	);
	LUT4 #(
		.INIT('h0001)
	) name56 (
		\pi041 ,
		\pi043 ,
		\pi047 ,
		\pi048 ,
		_w205_
	);
	LUT3 #(
		.INIT('h80)
	) name57 (
		_w202_,
		_w203_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\pi002 ,
		\pi020 ,
		_w207_
	);
	LUT4 #(
		.INIT('h0001)
	) name59 (
		\pi002 ,
		\pi015 ,
		\pi020 ,
		\pi049 ,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\pi024 ,
		\pi045 ,
		_w209_
	);
	LUT4 #(
		.INIT('h0111)
	) name61 (
		\pi024 ,
		\pi045 ,
		\pi122 ,
		\pi127 ,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w208_,
		_w210_,
		_w211_
	);
	LUT3 #(
		.INIT('h40)
	) name63 (
		\pi065 ,
		_w208_,
		_w210_,
		_w212_
	);
	LUT3 #(
		.INIT('h15)
	) name64 (
		_w200_,
		_w206_,
		_w212_,
		_w213_
	);
	LUT3 #(
		.INIT('h40)
	) name65 (
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w214_
	);
	LUT4 #(
		.INIT('h2000)
	) name66 (
		\pi002 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\pi045 ,
		\pi048 ,
		_w216_
	);
	LUT4 #(
		.INIT('h8000)
	) name68 (
		_w202_,
		_w203_,
		_w204_,
		_w216_,
		_w217_
	);
	LUT4 #(
		.INIT('h0001)
	) name69 (
		\pi015 ,
		\pi020 ,
		\pi024 ,
		\pi049 ,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\pi002 ,
		\pi082 ,
		_w219_
	);
	LUT4 #(
		.INIT('h4055)
	) name71 (
		_w215_,
		_w217_,
		_w218_,
		_w219_,
		_w220_
	);
	LUT3 #(
		.INIT('h15)
	) name72 (
		\pi129 ,
		_w213_,
		_w220_,
		_w221_
	);
	LUT4 #(
		.INIT('h0002)
	) name73 (
		\pi000 ,
		\pi113 ,
		\pi123 ,
		\pi129 ,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\pi009 ,
		\pi014 ,
		_w223_
	);
	LUT4 #(
		.INIT('h0001)
	) name75 (
		\pi007 ,
		\pi009 ,
		\pi012 ,
		\pi014 ,
		_w224_
	);
	LUT3 #(
		.INIT('h80)
	) name76 (
		_w177_,
		_w181_,
		_w224_,
		_w225_
	);
	LUT3 #(
		.INIT('h01)
	) name77 (
		\pi061 ,
		\pi118 ,
		\pi129 ,
		_w226_
	);
	LUT4 #(
		.INIT('hdfcc)
	) name78 (
		_w187_,
		_w222_,
		_w225_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\pi004 ,
		\pi054 ,
		_w228_
	);
	LUT4 #(
		.INIT('h0100)
	) name80 (
		\pi008 ,
		\pi011 ,
		\pi021 ,
		\pi054 ,
		_w229_
	);
	LUT3 #(
		.INIT('h80)
	) name81 (
		_w151_,
		_w152_,
		_w229_,
		_w230_
	);
	LUT3 #(
		.INIT('h02)
	) name82 (
		\pi010 ,
		\pi014 ,
		\pi022 ,
		_w231_
	);
	LUT3 #(
		.INIT('h80)
	) name83 (
		_w182_,
		_w185_,
		_w231_,
		_w232_
	);
	LUT4 #(
		.INIT('ha888)
	) name84 (
		_w149_,
		_w228_,
		_w230_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\pi005 ,
		\pi054 ,
		_w234_
	);
	LUT4 #(
		.INIT('h0001)
	) name86 (
		\pi008 ,
		\pi011 ,
		\pi017 ,
		\pi021 ,
		_w235_
	);
	LUT4 #(
		.INIT('h4000)
	) name87 (
		\pi059 ,
		_w177_,
		_w223_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		\pi016 ,
		\pi054 ,
		_w237_
	);
	LUT4 #(
		.INIT('h0001)
	) name89 (
		\pi004 ,
		\pi018 ,
		\pi019 ,
		\pi029 ,
		_w238_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\pi025 ,
		\pi028 ,
		_w239_
	);
	LUT4 #(
		.INIT('h8000)
	) name91 (
		_w182_,
		_w237_,
		_w238_,
		_w239_,
		_w240_
	);
	LUT4 #(
		.INIT('ha888)
	) name92 (
		_w149_,
		_w234_,
		_w236_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\pi006 ,
		\pi054 ,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\pi025 ,
		\pi028 ,
		_w243_
	);
	LUT4 #(
		.INIT('h8000)
	) name95 (
		_w182_,
		_w237_,
		_w238_,
		_w243_,
		_w244_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name96 (
		_w149_,
		_w236_,
		_w242_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\pi007 ,
		\pi054 ,
		_w246_
	);
	LUT4 #(
		.INIT('h0100)
	) name98 (
		\pi004 ,
		\pi016 ,
		\pi019 ,
		\pi054 ,
		_w247_
	);
	LUT4 #(
		.INIT('h8000)
	) name99 (
		_w177_,
		_w181_,
		_w224_,
		_w247_,
		_w248_
	);
	LUT3 #(
		.INIT('h01)
	) name100 (
		\pi011 ,
		\pi017 ,
		\pi018 ,
		_w249_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\pi008 ,
		\pi021 ,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w249_,
		_w250_,
		_w251_
	);
	LUT4 #(
		.INIT('ha888)
	) name103 (
		_w149_,
		_w246_,
		_w248_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		\pi008 ,
		\pi054 ,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\pi008 ,
		\pi021 ,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w249_,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name107 (
		_w149_,
		_w248_,
		_w253_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\pi009 ,
		\pi054 ,
		_w257_
	);
	LUT4 #(
		.INIT('h0001)
	) name109 (
		\pi008 ,
		\pi017 ,
		\pi018 ,
		\pi021 ,
		_w258_
	);
	LUT3 #(
		.INIT('h40)
	) name110 (
		\pi013 ,
		_w182_,
		_w258_,
		_w259_
	);
	LUT3 #(
		.INIT('h04)
	) name111 (
		\pi009 ,
		\pi011 ,
		\pi014 ,
		_w260_
	);
	LUT3 #(
		.INIT('h80)
	) name112 (
		_w176_,
		_w247_,
		_w260_,
		_w261_
	);
	LUT4 #(
		.INIT('ha888)
	) name113 (
		_w149_,
		_w257_,
		_w259_,
		_w261_,
		_w262_
	);
	LUT4 #(
		.INIT('h0004)
	) name114 (
		\pi003 ,
		\pi010 ,
		\pi054 ,
		\pi129 ,
		_w263_
	);
	LUT4 #(
		.INIT('h4000)
	) name115 (
		\pi009 ,
		_w176_,
		_w247_,
		_w258_,
		_w264_
	);
	LUT3 #(
		.INIT('h10)
	) name116 (
		\pi011 ,
		\pi013 ,
		\pi014 ,
		_w265_
	);
	LUT3 #(
		.INIT('h80)
	) name117 (
		_w149_,
		_w182_,
		_w265_,
		_w266_
	);
	LUT3 #(
		.INIT('hea)
	) name118 (
		_w263_,
		_w264_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\pi011 ,
		\pi054 ,
		_w268_
	);
	LUT3 #(
		.INIT('h10)
	) name120 (
		\pi009 ,
		\pi011 ,
		\pi022 ,
		_w269_
	);
	LUT3 #(
		.INIT('h80)
	) name121 (
		_w188_,
		_w247_,
		_w269_,
		_w270_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name122 (
		_w149_,
		_w259_,
		_w268_,
		_w270_,
		_w271_
	);
	LUT4 #(
		.INIT('h0004)
	) name123 (
		\pi003 ,
		\pi012 ,
		\pi054 ,
		\pi129 ,
		_w272_
	);
	LUT3 #(
		.INIT('h80)
	) name124 (
		\pi018 ,
		_w149_,
		_w235_,
		_w273_
	);
	LUT3 #(
		.INIT('hec)
	) name125 (
		_w248_,
		_w272_,
		_w273_,
		_w274_
	);
	LUT4 #(
		.INIT('h0004)
	) name126 (
		\pi003 ,
		\pi013 ,
		\pi054 ,
		\pi129 ,
		_w275_
	);
	LUT3 #(
		.INIT('h01)
	) name127 (
		\pi005 ,
		\pi006 ,
		\pi018 ,
		_w276_
	);
	LUT4 #(
		.INIT('h8000)
	) name128 (
		_w177_,
		_w224_,
		_w247_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\pi025 ,
		\pi028 ,
		_w278_
	);
	LUT4 #(
		.INIT('h0010)
	) name130 (
		\pi025 ,
		\pi028 ,
		\pi029 ,
		\pi059 ,
		_w279_
	);
	LUT3 #(
		.INIT('h80)
	) name131 (
		_w149_,
		_w235_,
		_w279_,
		_w280_
	);
	LUT3 #(
		.INIT('hea)
	) name132 (
		_w275_,
		_w277_,
		_w280_,
		_w281_
	);
	LUT4 #(
		.INIT('h0004)
	) name133 (
		\pi003 ,
		\pi014 ,
		\pi054 ,
		\pi129 ,
		_w282_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		\pi011 ,
		\pi013 ,
		_w283_
	);
	LUT4 #(
		.INIT('h8000)
	) name135 (
		_w151_,
		_w182_,
		_w189_,
		_w283_,
		_w284_
	);
	LUT3 #(
		.INIT('h40)
	) name136 (
		\pi009 ,
		_w149_,
		_w258_,
		_w285_
	);
	LUT3 #(
		.INIT('hea)
	) name137 (
		_w282_,
		_w284_,
		_w285_,
		_w286_
	);
	LUT3 #(
		.INIT('h01)
	) name138 (
		\pi015 ,
		\pi024 ,
		\pi049 ,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w207_,
		_w287_,
		_w288_
	);
	LUT3 #(
		.INIT('h80)
	) name140 (
		\pi082 ,
		_w217_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		\pi024 ,
		\pi049 ,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\pi015 ,
		\pi082 ,
		_w291_
	);
	LUT3 #(
		.INIT('h70)
	) name143 (
		_w217_,
		_w290_,
		_w291_,
		_w292_
	);
	LUT4 #(
		.INIT('h2000)
	) name144 (
		\pi015 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w293_
	);
	LUT3 #(
		.INIT('h15)
	) name145 (
		\pi070 ,
		\pi122 ,
		\pi127 ,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w293_,
		_w294_,
		_w295_
	);
	LUT4 #(
		.INIT('hcccc)
	) name147 (
		\pi015 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w296_
	);
	LUT4 #(
		.INIT('h080f)
	) name148 (
		_w217_,
		_w287_,
		_w295_,
		_w296_,
		_w297_
	);
	LUT4 #(
		.INIT('h5554)
	) name149 (
		\pi129 ,
		_w289_,
		_w292_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\pi016 ,
		\pi054 ,
		_w299_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		\pi005 ,
		\pi006 ,
		_w300_
	);
	LUT3 #(
		.INIT('h80)
	) name152 (
		_w177_,
		_w224_,
		_w300_,
		_w301_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name153 (
		_w149_,
		_w230_,
		_w299_,
		_w301_,
		_w302_
	);
	LUT4 #(
		.INIT('h0004)
	) name154 (
		\pi003 ,
		\pi017 ,
		\pi054 ,
		\pi129 ,
		_w303_
	);
	LUT3 #(
		.INIT('h40)
	) name155 (
		\pi029 ,
		\pi054 ,
		\pi059 ,
		_w304_
	);
	LUT3 #(
		.INIT('h80)
	) name156 (
		_w149_,
		_w278_,
		_w304_,
		_w305_
	);
	LUT4 #(
		.INIT('hf8f0)
	) name157 (
		_w187_,
		_w225_,
		_w303_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\pi018 ,
		\pi054 ,
		_w307_
	);
	LUT3 #(
		.INIT('h80)
	) name159 (
		_w177_,
		_w223_,
		_w235_,
		_w308_
	);
	LUT4 #(
		.INIT('h0004)
	) name160 (
		\pi004 ,
		\pi016 ,
		\pi018 ,
		\pi019 ,
		_w309_
	);
	LUT3 #(
		.INIT('h80)
	) name161 (
		\pi054 ,
		_w182_,
		_w309_,
		_w310_
	);
	LUT4 #(
		.INIT('ha888)
	) name162 (
		_w149_,
		_w307_,
		_w308_,
		_w310_,
		_w311_
	);
	LUT4 #(
		.INIT('h0004)
	) name163 (
		\pi003 ,
		\pi019 ,
		\pi054 ,
		\pi129 ,
		_w312_
	);
	LUT4 #(
		.INIT('h0010)
	) name164 (
		\pi008 ,
		\pi011 ,
		\pi017 ,
		\pi021 ,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w149_,
		_w313_,
		_w314_
	);
	LUT3 #(
		.INIT('hec)
	) name166 (
		_w277_,
		_w312_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\pi020 ,
		\pi082 ,
		_w316_
	);
	LUT3 #(
		.INIT('h20)
	) name168 (
		\pi002 ,
		\pi020 ,
		\pi082 ,
		_w317_
	);
	LUT4 #(
		.INIT('h078f)
	) name169 (
		_w217_,
		_w287_,
		_w316_,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('h2000)
	) name170 (
		\pi020 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w319_
	);
	LUT3 #(
		.INIT('h15)
	) name171 (
		\pi071 ,
		\pi122 ,
		\pi127 ,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w319_,
		_w320_,
		_w321_
	);
	LUT4 #(
		.INIT('hcccc)
	) name173 (
		\pi020 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w322_
	);
	LUT4 #(
		.INIT('h080f)
	) name174 (
		_w217_,
		_w218_,
		_w321_,
		_w322_,
		_w323_
	);
	LUT3 #(
		.INIT('h51)
	) name175 (
		\pi129 ,
		_w318_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\pi021 ,
		\pi054 ,
		_w325_
	);
	LUT4 #(
		.INIT('h0100)
	) name177 (
		\pi004 ,
		\pi016 ,
		\pi018 ,
		\pi019 ,
		_w326_
	);
	LUT3 #(
		.INIT('h80)
	) name178 (
		\pi054 ,
		_w182_,
		_w326_,
		_w327_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name179 (
		_w149_,
		_w308_,
		_w325_,
		_w327_,
		_w328_
	);
	LUT4 #(
		.INIT('h0004)
	) name180 (
		\pi003 ,
		\pi022 ,
		\pi054 ,
		\pi129 ,
		_w329_
	);
	LUT4 #(
		.INIT('h0002)
	) name181 (
		\pi005 ,
		\pi006 ,
		\pi011 ,
		\pi012 ,
		_w330_
	);
	LUT3 #(
		.INIT('h80)
	) name182 (
		_w149_,
		_w155_,
		_w330_,
		_w331_
	);
	LUT3 #(
		.INIT('hec)
	) name183 (
		_w264_,
		_w329_,
		_w331_,
		_w332_
	);
	LUT4 #(
		.INIT('h00b0)
	) name184 (
		\pi023 ,
		\pi055 ,
		\pi061 ,
		\pi129 ,
		_w333_
	);
	LUT3 #(
		.INIT('h2a)
	) name185 (
		\pi063 ,
		\pi122 ,
		\pi127 ,
		_w334_
	);
	LUT4 #(
		.INIT('h0222)
	) name186 (
		\pi063 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w208_,
		_w334_,
		_w336_
	);
	LUT3 #(
		.INIT('h13)
	) name188 (
		_w217_,
		_w335_,
		_w336_,
		_w337_
	);
	LUT4 #(
		.INIT('h5010)
	) name189 (
		\pi024 ,
		\pi082 ,
		_w198_,
		_w208_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		\pi024 ,
		\pi082 ,
		_w339_
	);
	LUT3 #(
		.INIT('h23)
	) name191 (
		_w217_,
		_w338_,
		_w339_,
		_w340_
	);
	LUT3 #(
		.INIT('h10)
	) name192 (
		\pi046 ,
		\pi050 ,
		\pi082 ,
		_w341_
	);
	LUT3 #(
		.INIT('h02)
	) name193 (
		\pi024 ,
		\pi045 ,
		\pi048 ,
		_w342_
	);
	LUT4 #(
		.INIT('h8000)
	) name194 (
		_w202_,
		_w204_,
		_w341_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\pi129 ,
		_w343_,
		_w344_
	);
	LUT3 #(
		.INIT('h80)
	) name196 (
		_w337_,
		_w340_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h9)
	) name197 (
		\pi053 ,
		\pi058 ,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\pi053 ,
		\pi058 ,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		\pi096 ,
		\pi110 ,
		_w348_
	);
	LUT3 #(
		.INIT('h54)
	) name200 (
		\pi085 ,
		\pi096 ,
		\pi110 ,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name201 (
		\pi085 ,
		\pi116 ,
		_w350_
	);
	LUT3 #(
		.INIT('hc4)
	) name202 (
		\pi085 ,
		\pi100 ,
		\pi116 ,
		_w351_
	);
	LUT3 #(
		.INIT('h08)
	) name203 (
		\pi025 ,
		\pi085 ,
		\pi116 ,
		_w352_
	);
	LUT4 #(
		.INIT('h5510)
	) name204 (
		\pi027 ,
		_w349_,
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		\pi026 ,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		\pi025 ,
		\pi116 ,
		_w355_
	);
	LUT4 #(
		.INIT('h0100)
	) name207 (
		\pi039 ,
		\pi051 ,
		\pi052 ,
		\pi116 ,
		_w356_
	);
	LUT3 #(
		.INIT('ha8)
	) name208 (
		\pi027 ,
		_w355_,
		_w356_,
		_w357_
	);
	LUT3 #(
		.INIT('h01)
	) name209 (
		\pi039 ,
		\pi051 ,
		\pi052 ,
		_w358_
	);
	LUT4 #(
		.INIT('haaa8)
	) name210 (
		\pi027 ,
		\pi039 ,
		\pi051 ,
		\pi052 ,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\pi025 ,
		\pi110 ,
		_w360_
	);
	LUT4 #(
		.INIT('h0002)
	) name212 (
		\pi025 ,
		\pi095 ,
		\pi097 ,
		\pi100 ,
		_w361_
	);
	LUT3 #(
		.INIT('h54)
	) name213 (
		_w359_,
		_w360_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\pi026 ,
		\pi085 ,
		_w363_
	);
	LUT3 #(
		.INIT('he0)
	) name215 (
		_w357_,
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\pi026 ,
		\pi085 ,
		_w365_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w356_,
		_w365_,
		_w366_
	);
	LUT3 #(
		.INIT('h32)
	) name218 (
		\pi025 ,
		\pi027 ,
		\pi116 ,
		_w367_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name219 (
		_w346_,
		_w356_,
		_w365_,
		_w367_,
		_w368_
	);
	LUT4 #(
		.INIT('h5455)
	) name220 (
		_w347_,
		_w354_,
		_w364_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		\pi053 ,
		\pi058 ,
		_w370_
	);
	LUT4 #(
		.INIT('h0001)
	) name222 (
		\pi003 ,
		\pi053 ,
		\pi058 ,
		\pi129 ,
		_w371_
	);
	LUT3 #(
		.INIT('h01)
	) name223 (
		\pi026 ,
		\pi027 ,
		\pi085 ,
		_w372_
	);
	LUT4 #(
		.INIT('h0004)
	) name224 (
		\pi003 ,
		\pi025 ,
		\pi116 ,
		\pi129 ,
		_w373_
	);
	LUT3 #(
		.INIT('h15)
	) name225 (
		_w371_,
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		_w369_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		\pi026 ,
		\pi116 ,
		_w376_
	);
	LUT3 #(
		.INIT('h04)
	) name228 (
		_w349_,
		_w351_,
		_w376_,
		_w377_
	);
	LUT3 #(
		.INIT('h01)
	) name229 (
		\pi027 ,
		\pi053 ,
		\pi058 ,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w149_,
		_w378_,
		_w379_
	);
	LUT3 #(
		.INIT('he0)
	) name231 (
		_w366_,
		_w377_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		\pi027 ,
		\pi085 ,
		_w381_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w356_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\pi085 ,
		\pi116 ,
		_w383_
	);
	LUT4 #(
		.INIT('h0004)
	) name235 (
		\pi085 ,
		\pi095 ,
		\pi096 ,
		\pi110 ,
		_w384_
	);
	LUT3 #(
		.INIT('h13)
	) name236 (
		\pi027 ,
		\pi100 ,
		\pi116 ,
		_w385_
	);
	LUT3 #(
		.INIT('he0)
	) name237 (
		_w383_,
		_w384_,
		_w385_,
		_w386_
	);
	LUT3 #(
		.INIT('h01)
	) name238 (
		\pi003 ,
		\pi026 ,
		\pi129 ,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w370_,
		_w387_,
		_w388_
	);
	LUT3 #(
		.INIT('he0)
	) name240 (
		_w382_,
		_w386_,
		_w388_,
		_w389_
	);
	LUT3 #(
		.INIT('h08)
	) name241 (
		\pi028 ,
		\pi053 ,
		\pi116 ,
		_w390_
	);
	LUT3 #(
		.INIT('h40)
	) name242 (
		\pi058 ,
		_w372_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h6)
	) name243 (
		\pi026 ,
		\pi027 ,
		_w392_
	);
	LUT4 #(
		.INIT('h0060)
	) name244 (
		\pi026 ,
		\pi027 ,
		\pi028 ,
		\pi116 ,
		_w393_
	);
	LUT4 #(
		.INIT('h5554)
	) name245 (
		\pi026 ,
		\pi039 ,
		\pi051 ,
		\pi052 ,
		_w394_
	);
	LUT4 #(
		.INIT('h0001)
	) name246 (
		\pi027 ,
		\pi039 ,
		\pi051 ,
		\pi052 ,
		_w395_
	);
	LUT3 #(
		.INIT('h01)
	) name247 (
		\pi095 ,
		\pi097 ,
		\pi100 ,
		_w396_
	);
	LUT4 #(
		.INIT('h00fe)
	) name248 (
		\pi095 ,
		\pi097 ,
		\pi100 ,
		\pi110 ,
		_w397_
	);
	LUT4 #(
		.INIT('h00a8)
	) name249 (
		\pi028 ,
		_w394_,
		_w395_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w393_,
		_w398_,
		_w399_
	);
	LUT3 #(
		.INIT('h04)
	) name251 (
		\pi026 ,
		\pi095 ,
		\pi100 ,
		_w400_
	);
	LUT4 #(
		.INIT('h135f)
	) name252 (
		\pi026 ,
		_w348_,
		_w356_,
		_w400_,
		_w401_
	);
	LUT3 #(
		.INIT('h40)
	) name253 (
		\pi026 ,
		\pi027 ,
		\pi116 ,
		_w402_
	);
	LUT3 #(
		.INIT('h45)
	) name254 (
		\pi085 ,
		_w358_,
		_w402_,
		_w403_
	);
	LUT3 #(
		.INIT('he0)
	) name255 (
		\pi027 ,
		_w401_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		\pi053 ,
		\pi085 ,
		_w405_
	);
	LUT4 #(
		.INIT('h1110)
	) name257 (
		\pi026 ,
		\pi027 ,
		\pi028 ,
		\pi116 ,
		_w406_
	);
	LUT3 #(
		.INIT('h15)
	) name258 (
		\pi053 ,
		\pi100 ,
		\pi116 ,
		_w407_
	);
	LUT4 #(
		.INIT('h5444)
	) name259 (
		\pi058 ,
		_w405_,
		_w406_,
		_w407_,
		_w408_
	);
	LUT4 #(
		.INIT('h4055)
	) name260 (
		_w391_,
		_w399_,
		_w404_,
		_w408_,
		_w409_
	);
	LUT3 #(
		.INIT('h01)
	) name261 (
		\pi026 ,
		\pi053 ,
		\pi085 ,
		_w410_
	);
	LUT4 #(
		.INIT('h0040)
	) name262 (
		\pi027 ,
		\pi028 ,
		\pi058 ,
		\pi116 ,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w410_,
		_w411_,
		_w412_
	);
	LUT3 #(
		.INIT('ha2)
	) name264 (
		_w149_,
		_w409_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		\pi029 ,
		\pi116 ,
		_w414_
	);
	LUT4 #(
		.INIT('h0008)
	) name266 (
		\pi026 ,
		\pi029 ,
		\pi085 ,
		\pi116 ,
		_w415_
	);
	LUT3 #(
		.INIT('h2a)
	) name267 (
		\pi026 ,
		_w378_,
		_w415_,
		_w416_
	);
	LUT3 #(
		.INIT('h02)
	) name268 (
		\pi027 ,
		\pi053 ,
		\pi058 ,
		_w417_
	);
	LUT3 #(
		.INIT('h40)
	) name269 (
		\pi085 ,
		_w414_,
		_w417_,
		_w418_
	);
	LUT4 #(
		.INIT('h0c44)
	) name270 (
		\pi029 ,
		\pi058 ,
		\pi097 ,
		\pi116 ,
		_w419_
	);
	LUT4 #(
		.INIT('h0008)
	) name271 (
		\pi029 ,
		\pi053 ,
		\pi058 ,
		\pi116 ,
		_w420_
	);
	LUT3 #(
		.INIT('h0e)
	) name272 (
		\pi053 ,
		_w419_,
		_w420_,
		_w421_
	);
	LUT4 #(
		.INIT('h0001)
	) name273 (
		\pi095 ,
		\pi096 ,
		\pi100 ,
		\pi110 ,
		_w422_
	);
	LUT3 #(
		.INIT('h15)
	) name274 (
		\pi058 ,
		\pi097 ,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\pi029 ,
		\pi110 ,
		_w424_
	);
	LUT4 #(
		.INIT('h0002)
	) name276 (
		\pi029 ,
		\pi095 ,
		\pi097 ,
		\pi100 ,
		_w425_
	);
	LUT3 #(
		.INIT('h01)
	) name277 (
		_w420_,
		_w424_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		\pi027 ,
		\pi085 ,
		_w427_
	);
	LUT4 #(
		.INIT('h1500)
	) name279 (
		_w421_,
		_w423_,
		_w426_,
		_w427_,
		_w428_
	);
	LUT3 #(
		.INIT('h08)
	) name280 (
		\pi029 ,
		\pi085 ,
		\pi116 ,
		_w429_
	);
	LUT3 #(
		.INIT('h57)
	) name281 (
		_w378_,
		_w415_,
		_w429_,
		_w430_
	);
	LUT4 #(
		.INIT('h5455)
	) name282 (
		_w416_,
		_w418_,
		_w428_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		_w149_,
		_w431_,
		_w432_
	);
	LUT4 #(
		.INIT('h0305)
	) name284 (
		\pi030 ,
		\pi060 ,
		\pi106 ,
		\pi109 ,
		_w433_
	);
	LUT3 #(
		.INIT('h0b)
	) name285 (
		\pi088 ,
		\pi106 ,
		\pi129 ,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w433_,
		_w434_,
		_w435_
	);
	LUT4 #(
		.INIT('h0503)
	) name287 (
		\pi030 ,
		\pi031 ,
		\pi106 ,
		\pi109 ,
		_w436_
	);
	LUT3 #(
		.INIT('h0b)
	) name288 (
		\pi089 ,
		\pi106 ,
		\pi129 ,
		_w437_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w436_,
		_w437_,
		_w438_
	);
	LUT4 #(
		.INIT('h0503)
	) name290 (
		\pi031 ,
		\pi032 ,
		\pi106 ,
		\pi109 ,
		_w439_
	);
	LUT3 #(
		.INIT('h0b)
	) name291 (
		\pi099 ,
		\pi106 ,
		\pi129 ,
		_w440_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		_w439_,
		_w440_,
		_w441_
	);
	LUT4 #(
		.INIT('h0503)
	) name293 (
		\pi032 ,
		\pi033 ,
		\pi106 ,
		\pi109 ,
		_w442_
	);
	LUT3 #(
		.INIT('h0b)
	) name294 (
		\pi090 ,
		\pi106 ,
		\pi129 ,
		_w443_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		_w442_,
		_w443_,
		_w444_
	);
	LUT4 #(
		.INIT('h0503)
	) name296 (
		\pi033 ,
		\pi034 ,
		\pi106 ,
		\pi109 ,
		_w445_
	);
	LUT3 #(
		.INIT('h0b)
	) name297 (
		\pi091 ,
		\pi106 ,
		\pi129 ,
		_w446_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w445_,
		_w446_,
		_w447_
	);
	LUT4 #(
		.INIT('h0503)
	) name299 (
		\pi034 ,
		\pi035 ,
		\pi106 ,
		\pi109 ,
		_w448_
	);
	LUT3 #(
		.INIT('h0b)
	) name300 (
		\pi092 ,
		\pi106 ,
		\pi129 ,
		_w449_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w448_,
		_w449_,
		_w450_
	);
	LUT4 #(
		.INIT('h0503)
	) name302 (
		\pi035 ,
		\pi036 ,
		\pi106 ,
		\pi109 ,
		_w451_
	);
	LUT3 #(
		.INIT('h0b)
	) name303 (
		\pi098 ,
		\pi106 ,
		\pi129 ,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w451_,
		_w452_,
		_w453_
	);
	LUT4 #(
		.INIT('h0503)
	) name305 (
		\pi036 ,
		\pi037 ,
		\pi106 ,
		\pi109 ,
		_w454_
	);
	LUT3 #(
		.INIT('h0b)
	) name306 (
		\pi093 ,
		\pi106 ,
		\pi129 ,
		_w455_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w454_,
		_w455_,
		_w456_
	);
	LUT3 #(
		.INIT('h01)
	) name308 (
		\pi024 ,
		\pi045 ,
		\pi048 ,
		_w457_
	);
	LUT4 #(
		.INIT('h8000)
	) name309 (
		_w203_,
		_w204_,
		_w208_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		\pi082 ,
		_w202_,
		_w459_
	);
	LUT4 #(
		.INIT('h0100)
	) name311 (
		\pi040 ,
		\pi042 ,
		\pi044 ,
		\pi082 ,
		_w460_
	);
	LUT4 #(
		.INIT('ha888)
	) name312 (
		\pi038 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w461_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT3 #(
		.INIT('h15)
	) name314 (
		\pi074 ,
		\pi122 ,
		\pi127 ,
		_w463_
	);
	LUT3 #(
		.INIT('hd0)
	) name315 (
		\pi082 ,
		_w202_,
		_w463_,
		_w464_
	);
	LUT4 #(
		.INIT('h000b)
	) name316 (
		_w458_,
		_w459_,
		_w462_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		\pi129 ,
		_w465_,
		_w466_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name318 (
		\pi039 ,
		\pi051 ,
		\pi052 ,
		\pi109 ,
		_w467_
	);
	LUT4 #(
		.INIT('h0100)
	) name319 (
		\pi039 ,
		\pi051 ,
		\pi052 ,
		\pi109 ,
		_w468_
	);
	LUT4 #(
		.INIT('h3332)
	) name320 (
		\pi106 ,
		\pi129 ,
		_w467_,
		_w468_,
		_w469_
	);
	LUT3 #(
		.INIT('he0)
	) name321 (
		\pi042 ,
		\pi044 ,
		\pi082 ,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w198_,
		_w470_,
		_w471_
	);
	LUT3 #(
		.INIT('h01)
	) name323 (
		\pi038 ,
		\pi046 ,
		\pi050 ,
		_w472_
	);
	LUT4 #(
		.INIT('h8000)
	) name324 (
		_w204_,
		_w208_,
		_w457_,
		_w472_,
		_w473_
	);
	LUT3 #(
		.INIT('h10)
	) name325 (
		\pi042 ,
		\pi044 ,
		\pi082 ,
		_w474_
	);
	LUT4 #(
		.INIT('h1011)
	) name326 (
		\pi040 ,
		_w471_,
		_w473_,
		_w474_,
		_w475_
	);
	LUT3 #(
		.INIT('h2a)
	) name327 (
		\pi073 ,
		\pi122 ,
		\pi127 ,
		_w476_
	);
	LUT4 #(
		.INIT('h0222)
	) name328 (
		\pi073 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w201_,
		_w476_,
		_w478_
	);
	LUT4 #(
		.INIT('h0200)
	) name330 (
		\pi040 ,
		\pi042 ,
		\pi044 ,
		\pi082 ,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		\pi129 ,
		_w479_,
		_w480_
	);
	LUT4 #(
		.INIT('h1300)
	) name332 (
		_w473_,
		_w477_,
		_w478_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w475_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		\pi043 ,
		\pi047 ,
		_w483_
	);
	LUT3 #(
		.INIT('h80)
	) name335 (
		_w208_,
		_w457_,
		_w483_,
		_w484_
	);
	LUT4 #(
		.INIT('h0100)
	) name336 (
		\pi041 ,
		\pi046 ,
		\pi050 ,
		\pi082 ,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w202_,
		_w485_,
		_w486_
	);
	LUT4 #(
		.INIT('ha888)
	) name338 (
		\pi041 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w487_
	);
	LUT3 #(
		.INIT('h70)
	) name339 (
		_w202_,
		_w341_,
		_w487_,
		_w488_
	);
	LUT3 #(
		.INIT('h01)
	) name340 (
		\pi041 ,
		\pi046 ,
		\pi050 ,
		_w489_
	);
	LUT3 #(
		.INIT('h15)
	) name341 (
		\pi076 ,
		\pi122 ,
		\pi127 ,
		_w490_
	);
	LUT4 #(
		.INIT('hd500)
	) name342 (
		\pi082 ,
		_w202_,
		_w489_,
		_w490_,
		_w491_
	);
	LUT4 #(
		.INIT('h000b)
	) name343 (
		_w484_,
		_w486_,
		_w488_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		\pi129 ,
		_w492_,
		_w493_
	);
	LUT3 #(
		.INIT('h15)
	) name345 (
		\pi072 ,
		\pi122 ,
		\pi127 ,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w470_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('h0001)
	) name347 (
		\pi038 ,
		\pi040 ,
		\pi046 ,
		\pi050 ,
		_w496_
	);
	LUT4 #(
		.INIT('h8000)
	) name348 (
		_w204_,
		_w208_,
		_w457_,
		_w496_,
		_w497_
	);
	LUT3 #(
		.INIT('h8a)
	) name349 (
		\pi042 ,
		\pi044 ,
		\pi082 ,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w199_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('h0031)
	) name351 (
		_w474_,
		_w495_,
		_w497_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		\pi129 ,
		_w500_,
		_w501_
	);
	LUT3 #(
		.INIT('h40)
	) name353 (
		\pi047 ,
		_w208_,
		_w457_,
		_w502_
	);
	LUT4 #(
		.INIT('h0001)
	) name354 (
		\pi041 ,
		\pi043 ,
		\pi046 ,
		\pi050 ,
		_w503_
	);
	LUT3 #(
		.INIT('h80)
	) name355 (
		\pi082 ,
		_w202_,
		_w503_,
		_w504_
	);
	LUT4 #(
		.INIT('ha888)
	) name356 (
		\pi043 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w505_
	);
	LUT3 #(
		.INIT('h70)
	) name357 (
		_w202_,
		_w485_,
		_w505_,
		_w506_
	);
	LUT3 #(
		.INIT('h15)
	) name358 (
		\pi077 ,
		\pi122 ,
		\pi127 ,
		_w507_
	);
	LUT4 #(
		.INIT('hd500)
	) name359 (
		\pi082 ,
		_w202_,
		_w503_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('h000b)
	) name360 (
		_w502_,
		_w504_,
		_w506_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		\pi129 ,
		_w509_,
		_w510_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name362 (
		\pi044 ,
		\pi067 ,
		\pi122 ,
		\pi127 ,
		_w511_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\pi082 ,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h4)
	) name364 (
		\pi042 ,
		_w511_,
		_w513_
	);
	LUT3 #(
		.INIT('h07)
	) name365 (
		\pi044 ,
		\pi082 ,
		\pi129 ,
		_w514_
	);
	LUT4 #(
		.INIT('h1300)
	) name366 (
		_w497_,
		_w512_,
		_w513_,
		_w514_,
		_w515_
	);
	LUT4 #(
		.INIT('h2000)
	) name367 (
		\pi045 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		\pi045 ,
		\pi082 ,
		_w517_
	);
	LUT4 #(
		.INIT('h7f00)
	) name369 (
		_w202_,
		_w203_,
		_w205_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w516_,
		_w518_,
		_w519_
	);
	LUT3 #(
		.INIT('h15)
	) name371 (
		\pi068 ,
		\pi122 ,
		\pi127 ,
		_w520_
	);
	LUT4 #(
		.INIT('h0073)
	) name372 (
		\pi024 ,
		\pi082 ,
		_w208_,
		_w520_,
		_w521_
	);
	LUT3 #(
		.INIT('h0d)
	) name373 (
		\pi082 ,
		_w217_,
		_w521_,
		_w522_
	);
	LUT3 #(
		.INIT('h51)
	) name374 (
		\pi129 ,
		_w519_,
		_w522_,
		_w523_
	);
	LUT4 #(
		.INIT('h0111)
	) name375 (
		\pi075 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		\pi050 ,
		\pi082 ,
		_w525_
	);
	LUT4 #(
		.INIT('ha888)
	) name377 (
		\pi046 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w526_
	);
	LUT4 #(
		.INIT('h2033)
	) name378 (
		_w202_,
		_w524_,
		_w525_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\pi129 ,
		_w527_,
		_w528_
	);
	LUT3 #(
		.INIT('h15)
	) name380 (
		\pi075 ,
		\pi122 ,
		\pi127 ,
		_w529_
	);
	LUT4 #(
		.INIT('h3222)
	) name381 (
		\pi075 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w530_
	);
	LUT4 #(
		.INIT('h0080)
	) name382 (
		_w204_,
		_w208_,
		_w457_,
		_w529_,
		_w531_
	);
	LUT3 #(
		.INIT('h40)
	) name383 (
		\pi129 ,
		_w202_,
		_w203_,
		_w532_
	);
	LUT3 #(
		.INIT('h10)
	) name384 (
		_w530_,
		_w531_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('he)
	) name385 (
		_w528_,
		_w533_,
		_w534_
	);
	LUT3 #(
		.INIT('h15)
	) name386 (
		\pi064 ,
		\pi122 ,
		\pi127 ,
		_w535_
	);
	LUT4 #(
		.INIT('h00d5)
	) name387 (
		\pi082 ,
		_w208_,
		_w457_,
		_w535_,
		_w536_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name388 (
		\pi082 ,
		_w202_,
		_w203_,
		_w204_,
		_w537_
	);
	LUT4 #(
		.INIT('h2000)
	) name389 (
		\pi047 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\pi047 ,
		\pi082 ,
		_w539_
	);
	LUT4 #(
		.INIT('h080f)
	) name391 (
		_w202_,
		_w503_,
		_w538_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('h0155)
	) name392 (
		\pi129 ,
		_w536_,
		_w537_,
		_w540_,
		_w541_
	);
	LUT4 #(
		.INIT('h0080)
	) name393 (
		_w202_,
		_w203_,
		_w204_,
		_w214_,
		_w542_
	);
	LUT3 #(
		.INIT('h02)
	) name394 (
		\pi048 ,
		_w199_,
		_w542_,
		_w543_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name395 (
		\pi082 ,
		_w202_,
		_w203_,
		_w205_,
		_w544_
	);
	LUT3 #(
		.INIT('h15)
	) name396 (
		\pi062 ,
		\pi122 ,
		\pi127 ,
		_w545_
	);
	LUT4 #(
		.INIT('h00d5)
	) name397 (
		\pi082 ,
		_w208_,
		_w209_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w544_,
		_w546_,
		_w547_
	);
	LUT3 #(
		.INIT('h54)
	) name399 (
		\pi129 ,
		_w543_,
		_w547_,
		_w548_
	);
	LUT3 #(
		.INIT('h0d)
	) name400 (
		\pi082 ,
		_w208_,
		_w214_,
		_w549_
	);
	LUT4 #(
		.INIT('h4555)
	) name401 (
		\pi024 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w550_
	);
	LUT4 #(
		.INIT('h020a)
	) name402 (
		\pi049 ,
		_w217_,
		_w549_,
		_w550_,
		_w551_
	);
	LUT3 #(
		.INIT('h15)
	) name403 (
		\pi069 ,
		\pi122 ,
		\pi127 ,
		_w552_
	);
	LUT3 #(
		.INIT('h0d)
	) name404 (
		\pi082 ,
		_w208_,
		_w552_,
		_w553_
	);
	LUT4 #(
		.INIT('h00d5)
	) name405 (
		\pi082 ,
		_w217_,
		_w290_,
		_w553_,
		_w554_
	);
	LUT3 #(
		.INIT('h54)
	) name406 (
		\pi129 ,
		_w551_,
		_w554_,
		_w555_
	);
	LUT3 #(
		.INIT('h31)
	) name407 (
		\pi082 ,
		_w198_,
		_w202_,
		_w556_
	);
	LUT4 #(
		.INIT('h0001)
	) name408 (
		\pi041 ,
		\pi043 ,
		\pi046 ,
		\pi047 ,
		_w557_
	);
	LUT3 #(
		.INIT('h80)
	) name409 (
		_w208_,
		_w457_,
		_w557_,
		_w558_
	);
	LUT4 #(
		.INIT('h1011)
	) name410 (
		\pi050 ,
		_w556_,
		_w558_,
		_w459_,
		_w559_
	);
	LUT3 #(
		.INIT('h2a)
	) name411 (
		\pi066 ,
		\pi122 ,
		\pi127 ,
		_w560_
	);
	LUT4 #(
		.INIT('h0222)
	) name412 (
		\pi066 ,
		\pi082 ,
		\pi122 ,
		\pi127 ,
		_w561_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w202_,
		_w560_,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\pi050 ,
		\pi082 ,
		_w563_
	);
	LUT3 #(
		.INIT('h15)
	) name415 (
		\pi129 ,
		_w202_,
		_w563_,
		_w564_
	);
	LUT4 #(
		.INIT('h1300)
	) name416 (
		_w558_,
		_w561_,
		_w562_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		_w559_,
		_w565_,
		_w566_
	);
	LUT4 #(
		.INIT('h00de)
	) name418 (
		\pi051 ,
		\pi106 ,
		\pi109 ,
		\pi129 ,
		_w567_
	);
	LUT4 #(
		.INIT('h0603)
	) name419 (
		\pi051 ,
		\pi052 ,
		\pi106 ,
		\pi109 ,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		\pi129 ,
		_w568_,
		_w569_
	);
	LUT3 #(
		.INIT('hb1)
	) name421 (
		\pi053 ,
		\pi097 ,
		\pi116 ,
		_w570_
	);
	LUT3 #(
		.INIT('h31)
	) name422 (
		\pi053 ,
		\pi058 ,
		\pi116 ,
		_w571_
	);
	LUT3 #(
		.INIT('h23)
	) name423 (
		_w422_,
		_w570_,
		_w571_,
		_w572_
	);
	LUT4 #(
		.INIT('h0051)
	) name424 (
		\pi003 ,
		\pi058 ,
		\pi116 ,
		\pi129 ,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w372_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w572_,
		_w574_,
		_w575_
	);
	LUT4 #(
		.INIT('h00ea)
	) name427 (
		\pi082 ,
		\pi122 ,
		\pi127 ,
		\pi129 ,
		_w576_
	);
	LUT3 #(
		.INIT('h8f)
	) name428 (
		_w206_,
		_w211_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('he)
	) name429 (
		\pi123 ,
		\pi129 ,
		_w578_
	);
	LUT4 #(
		.INIT('h0002)
	) name430 (
		\pi114 ,
		\pi122 ,
		\pi123 ,
		\pi129 ,
		_w579_
	);
	LUT3 #(
		.INIT('h04)
	) name431 (
		\pi026 ,
		\pi037 ,
		\pi058 ,
		_w580_
	);
	LUT4 #(
		.INIT('h9fbf)
	) name432 (
		\pi026 ,
		\pi058 ,
		\pi094 ,
		\pi116 ,
		_w581_
	);
	LUT4 #(
		.INIT('h500c)
	) name433 (
		\pi026 ,
		\pi037 ,
		\pi058 ,
		\pi116 ,
		_w582_
	);
	LUT4 #(
		.INIT('h2232)
	) name434 (
		\pi053 ,
		_w580_,
		_w581_,
		_w582_,
		_w583_
	);
	LUT4 #(
		.INIT('h0004)
	) name435 (
		\pi026 ,
		\pi037 ,
		\pi053 ,
		\pi058 ,
		_w584_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		\pi085 ,
		_w584_,
		_w585_
	);
	LUT3 #(
		.INIT('h01)
	) name437 (
		\pi003 ,
		\pi027 ,
		\pi129 ,
		_w586_
	);
	LUT4 #(
		.INIT('h0001)
	) name438 (
		\pi003 ,
		\pi053 ,
		\pi085 ,
		\pi129 ,
		_w587_
	);
	LUT3 #(
		.INIT('h13)
	) name439 (
		_w580_,
		_w586_,
		_w587_,
		_w588_
	);
	LUT3 #(
		.INIT('h01)
	) name440 (
		_w583_,
		_w585_,
		_w588_,
		_w589_
	);
	LUT3 #(
		.INIT('h80)
	) name441 (
		\pi058 ,
		\pi060 ,
		\pi116 ,
		_w590_
	);
	LUT3 #(
		.INIT('h40)
	) name442 (
		\pi027 ,
		_w410_,
		_w590_,
		_w591_
	);
	LUT4 #(
		.INIT('h0001)
	) name443 (
		\pi026 ,
		\pi053 ,
		\pi085 ,
		\pi116 ,
		_w592_
	);
	LUT4 #(
		.INIT('h0107)
	) name444 (
		\pi026 ,
		\pi053 ,
		\pi058 ,
		\pi085 ,
		_w593_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		\pi027 ,
		\pi057 ,
		_w594_
	);
	LUT3 #(
		.INIT('he0)
	) name446 (
		_w592_,
		_w593_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		\pi057 ,
		\pi058 ,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w410_,
		_w596_,
		_w597_
	);
	LUT4 #(
		.INIT('haaa8)
	) name449 (
		_w149_,
		_w591_,
		_w595_,
		_w597_,
		_w598_
	);
	LUT4 #(
		.INIT('h0010)
	) name450 (
		\pi026 ,
		\pi027 ,
		\pi058 ,
		\pi116 ,
		_w599_
	);
	LUT3 #(
		.INIT('h06)
	) name451 (
		\pi026 ,
		\pi027 ,
		\pi058 ,
		_w600_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name452 (
		_w356_,
		_w587_,
		_w599_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		\pi059 ,
		\pi116 ,
		_w602_
	);
	LUT4 #(
		.INIT('h0008)
	) name454 (
		\pi026 ,
		\pi059 ,
		\pi085 ,
		\pi116 ,
		_w603_
	);
	LUT3 #(
		.INIT('h80)
	) name455 (
		_w149_,
		_w378_,
		_w603_,
		_w604_
	);
	LUT3 #(
		.INIT('h02)
	) name456 (
		\pi059 ,
		\pi085 ,
		\pi116 ,
		_w605_
	);
	LUT3 #(
		.INIT('h2a)
	) name457 (
		\pi027 ,
		_w370_,
		_w605_,
		_w606_
	);
	LUT4 #(
		.INIT('h0060)
	) name458 (
		\pi053 ,
		\pi058 ,
		\pi059 ,
		\pi116 ,
		_w607_
	);
	LUT2 #(
		.INIT('h4)
	) name459 (
		\pi085 ,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		\pi059 ,
		\pi110 ,
		_w609_
	);
	LUT4 #(
		.INIT('h0001)
	) name461 (
		\pi059 ,
		\pi095 ,
		\pi097 ,
		\pi100 ,
		_w610_
	);
	LUT3 #(
		.INIT('h02)
	) name462 (
		_w370_,
		_w609_,
		_w610_,
		_w611_
	);
	LUT3 #(
		.INIT('h51)
	) name463 (
		\pi085 ,
		_w348_,
		_w396_,
		_w612_
	);
	LUT4 #(
		.INIT('h1fff)
	) name464 (
		\pi027 ,
		\pi085 ,
		_w370_,
		_w602_,
		_w613_
	);
	LUT4 #(
		.INIT('h1500)
	) name465 (
		_w608_,
		_w611_,
		_w612_,
		_w613_,
		_w614_
	);
	LUT4 #(
		.INIT('hccce)
	) name466 (
		_w387_,
		_w604_,
		_w606_,
		_w614_,
		_w615_
	);
	LUT4 #(
		.INIT('haba8)
	) name467 (
		\pi060 ,
		\pi117 ,
		\pi122 ,
		\pi123 ,
		_w616_
	);
	LUT4 #(
		.INIT('h0010)
	) name468 (
		\pi114 ,
		\pi122 ,
		\pi123 ,
		\pi129 ,
		_w617_
	);
	LUT4 #(
		.INIT('h0080)
	) name469 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi138 ,
		_w618_
	);
	LUT3 #(
		.INIT('h20)
	) name470 (
		\pi136 ,
		\pi137 ,
		\pi140 ,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		\pi062 ,
		\pi129 ,
		_w620_
	);
	LUT3 #(
		.INIT('h04)
	) name472 (
		\pi129 ,
		\pi136 ,
		\pi137 ,
		_w621_
	);
	LUT4 #(
		.INIT('h8d8f)
	) name473 (
		_w618_,
		_w619_,
		_w620_,
		_w621_,
		_w622_
	);
	LUT3 #(
		.INIT('h20)
	) name474 (
		\pi136 ,
		\pi137 ,
		\pi142 ,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name475 (
		\pi063 ,
		\pi129 ,
		_w624_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name476 (
		_w618_,
		_w621_,
		_w623_,
		_w624_,
		_w625_
	);
	LUT3 #(
		.INIT('h20)
	) name477 (
		\pi136 ,
		\pi137 ,
		\pi139 ,
		_w626_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		\pi064 ,
		\pi129 ,
		_w627_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name479 (
		_w618_,
		_w621_,
		_w626_,
		_w627_,
		_w628_
	);
	LUT3 #(
		.INIT('h20)
	) name480 (
		\pi136 ,
		\pi137 ,
		\pi146 ,
		_w629_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		\pi065 ,
		\pi129 ,
		_w630_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name482 (
		_w618_,
		_w621_,
		_w629_,
		_w630_,
		_w631_
	);
	LUT3 #(
		.INIT('h10)
	) name483 (
		\pi136 ,
		\pi137 ,
		\pi143 ,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\pi066 ,
		\pi129 ,
		_w633_
	);
	LUT3 #(
		.INIT('h01)
	) name485 (
		\pi129 ,
		\pi136 ,
		\pi137 ,
		_w634_
	);
	LUT4 #(
		.INIT('h8d8f)
	) name486 (
		_w618_,
		_w632_,
		_w633_,
		_w634_,
		_w635_
	);
	LUT3 #(
		.INIT('h10)
	) name487 (
		\pi136 ,
		\pi137 ,
		\pi139 ,
		_w636_
	);
	LUT2 #(
		.INIT('h2)
	) name488 (
		\pi067 ,
		\pi129 ,
		_w637_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name489 (
		_w618_,
		_w634_,
		_w636_,
		_w637_,
		_w638_
	);
	LUT3 #(
		.INIT('h20)
	) name490 (
		\pi136 ,
		\pi137 ,
		\pi141 ,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		\pi068 ,
		\pi129 ,
		_w640_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name492 (
		_w618_,
		_w621_,
		_w639_,
		_w640_,
		_w641_
	);
	LUT3 #(
		.INIT('h20)
	) name493 (
		\pi136 ,
		\pi137 ,
		\pi143 ,
		_w642_
	);
	LUT2 #(
		.INIT('h2)
	) name494 (
		\pi069 ,
		\pi129 ,
		_w643_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name495 (
		_w618_,
		_w621_,
		_w642_,
		_w643_,
		_w644_
	);
	LUT3 #(
		.INIT('h20)
	) name496 (
		\pi136 ,
		\pi137 ,
		\pi144 ,
		_w645_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		\pi070 ,
		\pi129 ,
		_w646_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name498 (
		_w618_,
		_w621_,
		_w645_,
		_w646_,
		_w647_
	);
	LUT3 #(
		.INIT('h20)
	) name499 (
		\pi136 ,
		\pi137 ,
		\pi145 ,
		_w648_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		\pi071 ,
		\pi129 ,
		_w649_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name501 (
		_w618_,
		_w621_,
		_w648_,
		_w649_,
		_w650_
	);
	LUT3 #(
		.INIT('h10)
	) name502 (
		\pi136 ,
		\pi137 ,
		\pi140 ,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name503 (
		\pi072 ,
		\pi129 ,
		_w652_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name504 (
		_w618_,
		_w634_,
		_w651_,
		_w652_,
		_w653_
	);
	LUT3 #(
		.INIT('h10)
	) name505 (
		\pi136 ,
		\pi137 ,
		\pi141 ,
		_w654_
	);
	LUT2 #(
		.INIT('h2)
	) name506 (
		\pi073 ,
		\pi129 ,
		_w655_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name507 (
		_w618_,
		_w634_,
		_w654_,
		_w655_,
		_w656_
	);
	LUT3 #(
		.INIT('h10)
	) name508 (
		\pi136 ,
		\pi137 ,
		\pi142 ,
		_w657_
	);
	LUT2 #(
		.INIT('h2)
	) name509 (
		\pi074 ,
		\pi129 ,
		_w658_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name510 (
		_w618_,
		_w634_,
		_w657_,
		_w658_,
		_w659_
	);
	LUT3 #(
		.INIT('h10)
	) name511 (
		\pi136 ,
		\pi137 ,
		\pi144 ,
		_w660_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		\pi075 ,
		\pi129 ,
		_w661_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name513 (
		_w618_,
		_w634_,
		_w660_,
		_w661_,
		_w662_
	);
	LUT3 #(
		.INIT('h10)
	) name514 (
		\pi136 ,
		\pi137 ,
		\pi145 ,
		_w663_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		\pi076 ,
		\pi129 ,
		_w664_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name516 (
		_w618_,
		_w634_,
		_w663_,
		_w664_,
		_w665_
	);
	LUT3 #(
		.INIT('h10)
	) name517 (
		\pi136 ,
		\pi137 ,
		\pi146 ,
		_w666_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		\pi077 ,
		\pi129 ,
		_w667_
	);
	LUT4 #(
		.INIT('ha0f7)
	) name519 (
		_w618_,
		_w634_,
		_w666_,
		_w667_,
		_w668_
	);
	LUT3 #(
		.INIT('h04)
	) name520 (
		\pi136 ,
		\pi137 ,
		\pi142 ,
		_w669_
	);
	LUT2 #(
		.INIT('h2)
	) name521 (
		\pi078 ,
		\pi129 ,
		_w670_
	);
	LUT3 #(
		.INIT('h10)
	) name522 (
		\pi129 ,
		\pi136 ,
		\pi137 ,
		_w671_
	);
	LUT4 #(
		.INIT('h7270)
	) name523 (
		_w618_,
		_w669_,
		_w670_,
		_w671_,
		_w672_
	);
	LUT3 #(
		.INIT('h04)
	) name524 (
		\pi136 ,
		\pi137 ,
		\pi143 ,
		_w673_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\pi079 ,
		\pi129 ,
		_w674_
	);
	LUT4 #(
		.INIT('h5f08)
	) name526 (
		_w618_,
		_w671_,
		_w673_,
		_w674_,
		_w675_
	);
	LUT3 #(
		.INIT('h04)
	) name527 (
		\pi136 ,
		\pi137 ,
		\pi144 ,
		_w676_
	);
	LUT2 #(
		.INIT('h2)
	) name528 (
		\pi080 ,
		\pi129 ,
		_w677_
	);
	LUT4 #(
		.INIT('h5f08)
	) name529 (
		_w618_,
		_w671_,
		_w676_,
		_w677_,
		_w678_
	);
	LUT3 #(
		.INIT('h04)
	) name530 (
		\pi136 ,
		\pi137 ,
		\pi145 ,
		_w679_
	);
	LUT2 #(
		.INIT('h2)
	) name531 (
		\pi081 ,
		\pi129 ,
		_w680_
	);
	LUT4 #(
		.INIT('h5f08)
	) name532 (
		_w618_,
		_w671_,
		_w679_,
		_w680_,
		_w681_
	);
	LUT3 #(
		.INIT('h04)
	) name533 (
		\pi136 ,
		\pi137 ,
		\pi146 ,
		_w682_
	);
	LUT2 #(
		.INIT('h2)
	) name534 (
		\pi082 ,
		\pi129 ,
		_w683_
	);
	LUT4 #(
		.INIT('h5f08)
	) name535 (
		_w618_,
		_w671_,
		_w682_,
		_w683_,
		_w684_
	);
	LUT4 #(
		.INIT('h0080)
	) name536 (
		\pi031 ,
		\pi136 ,
		\pi137 ,
		\pi138 ,
		_w685_
	);
	LUT3 #(
		.INIT('h32)
	) name537 (
		\pi087 ,
		\pi136 ,
		\pi138 ,
		_w686_
	);
	LUT3 #(
		.INIT('h4c)
	) name538 (
		\pi115 ,
		\pi137 ,
		\pi138 ,
		_w687_
	);
	LUT3 #(
		.INIT('h15)
	) name539 (
		_w685_,
		_w686_,
		_w687_,
		_w688_
	);
	LUT4 #(
		.INIT('hc050)
	) name540 (
		\pi062 ,
		\pi089 ,
		\pi136 ,
		\pi138 ,
		_w689_
	);
	LUT4 #(
		.INIT('h0c05)
	) name541 (
		\pi072 ,
		\pi119 ,
		\pi136 ,
		\pi138 ,
		_w690_
	);
	LUT3 #(
		.INIT('h54)
	) name542 (
		\pi137 ,
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('hd)
	) name543 (
		_w688_,
		_w691_,
		_w692_
	);
	LUT3 #(
		.INIT('h04)
	) name544 (
		\pi136 ,
		\pi137 ,
		\pi141 ,
		_w693_
	);
	LUT2 #(
		.INIT('h2)
	) name545 (
		\pi084 ,
		\pi129 ,
		_w694_
	);
	LUT4 #(
		.INIT('h5f08)
	) name546 (
		_w618_,
		_w671_,
		_w693_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		\pi085 ,
		\pi110 ,
		_w696_
	);
	LUT3 #(
		.INIT('h04)
	) name548 (
		\pi085 ,
		\pi096 ,
		\pi110 ,
		_w697_
	);
	LUT3 #(
		.INIT('h45)
	) name549 (
		_w350_,
		_w396_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		_w378_,
		_w387_,
		_w699_
	);
	LUT2 #(
		.INIT('h4)
	) name551 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT3 #(
		.INIT('h04)
	) name552 (
		\pi136 ,
		\pi137 ,
		\pi139 ,
		_w701_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		\pi086 ,
		\pi129 ,
		_w702_
	);
	LUT4 #(
		.INIT('h5f08)
	) name554 (
		_w618_,
		_w671_,
		_w701_,
		_w702_,
		_w703_
	);
	LUT3 #(
		.INIT('h04)
	) name555 (
		\pi136 ,
		\pi137 ,
		\pi140 ,
		_w704_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		\pi087 ,
		\pi129 ,
		_w705_
	);
	LUT4 #(
		.INIT('h5f08)
	) name557 (
		_w618_,
		_w671_,
		_w704_,
		_w705_,
		_w706_
	);
	LUT3 #(
		.INIT('h80)
	) name558 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		_w707_
	);
	LUT3 #(
		.INIT('h08)
	) name559 (
		\pi136 ,
		\pi137 ,
		\pi138 ,
		_w708_
	);
	LUT3 #(
		.INIT('h15)
	) name560 (
		\pi088 ,
		_w707_,
		_w708_,
		_w709_
	);
	LUT4 #(
		.INIT('h0080)
	) name561 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi139 ,
		_w710_
	);
	LUT3 #(
		.INIT('h15)
	) name562 (
		\pi129 ,
		_w708_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w709_,
		_w711_,
		_w712_
	);
	LUT3 #(
		.INIT('h15)
	) name564 (
		\pi089 ,
		_w707_,
		_w708_,
		_w713_
	);
	LUT4 #(
		.INIT('h0080)
	) name565 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi140 ,
		_w714_
	);
	LUT3 #(
		.INIT('h15)
	) name566 (
		\pi129 ,
		_w708_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h4)
	) name567 (
		_w713_,
		_w715_,
		_w716_
	);
	LUT3 #(
		.INIT('h15)
	) name568 (
		\pi090 ,
		_w707_,
		_w708_,
		_w717_
	);
	LUT4 #(
		.INIT('h0080)
	) name569 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi142 ,
		_w718_
	);
	LUT3 #(
		.INIT('h15)
	) name570 (
		\pi129 ,
		_w708_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w717_,
		_w719_,
		_w720_
	);
	LUT3 #(
		.INIT('h15)
	) name572 (
		\pi091 ,
		_w707_,
		_w708_,
		_w721_
	);
	LUT4 #(
		.INIT('h0080)
	) name573 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi143 ,
		_w722_
	);
	LUT3 #(
		.INIT('h15)
	) name574 (
		\pi129 ,
		_w708_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w721_,
		_w723_,
		_w724_
	);
	LUT3 #(
		.INIT('h15)
	) name576 (
		\pi092 ,
		_w707_,
		_w708_,
		_w725_
	);
	LUT4 #(
		.INIT('h0080)
	) name577 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi144 ,
		_w726_
	);
	LUT3 #(
		.INIT('h15)
	) name578 (
		\pi129 ,
		_w708_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h4)
	) name579 (
		_w725_,
		_w727_,
		_w728_
	);
	LUT3 #(
		.INIT('h15)
	) name580 (
		\pi093 ,
		_w707_,
		_w708_,
		_w729_
	);
	LUT4 #(
		.INIT('h0080)
	) name581 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi146 ,
		_w730_
	);
	LUT3 #(
		.INIT('h15)
	) name582 (
		\pi129 ,
		_w708_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w729_,
		_w731_,
		_w732_
	);
	LUT4 #(
		.INIT('h0200)
	) name584 (
		\pi082 ,
		\pi136 ,
		\pi137 ,
		\pi138 ,
		_w733_
	);
	LUT3 #(
		.INIT('h15)
	) name585 (
		\pi094 ,
		_w707_,
		_w733_,
		_w734_
	);
	LUT3 #(
		.INIT('h15)
	) name586 (
		\pi129 ,
		_w718_,
		_w733_,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		_w734_,
		_w735_,
		_w736_
	);
	LUT4 #(
		.INIT('h8000)
	) name588 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi143 ,
		_w737_
	);
	LUT3 #(
		.INIT('h40)
	) name589 (
		\pi129 ,
		_w733_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		\pi003 ,
		\pi110 ,
		_w739_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		\pi095 ,
		\pi129 ,
		_w740_
	);
	LUT4 #(
		.INIT('h7200)
	) name592 (
		_w707_,
		_w733_,
		_w739_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('he)
	) name593 (
		_w738_,
		_w741_,
		_w742_
	);
	LUT4 #(
		.INIT('h8000)
	) name594 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi146 ,
		_w743_
	);
	LUT3 #(
		.INIT('h40)
	) name595 (
		\pi129 ,
		_w733_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		\pi096 ,
		\pi129 ,
		_w745_
	);
	LUT4 #(
		.INIT('h7200)
	) name597 (
		_w707_,
		_w733_,
		_w739_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('he)
	) name598 (
		_w744_,
		_w746_,
		_w747_
	);
	LUT4 #(
		.INIT('h8000)
	) name599 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi145 ,
		_w748_
	);
	LUT3 #(
		.INIT('h40)
	) name600 (
		\pi129 ,
		_w733_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		\pi097 ,
		\pi129 ,
		_w750_
	);
	LUT4 #(
		.INIT('h7200)
	) name602 (
		_w707_,
		_w733_,
		_w739_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('he)
	) name603 (
		_w749_,
		_w751_,
		_w752_
	);
	LUT3 #(
		.INIT('h15)
	) name604 (
		\pi098 ,
		_w707_,
		_w708_,
		_w753_
	);
	LUT4 #(
		.INIT('h0080)
	) name605 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi145 ,
		_w754_
	);
	LUT3 #(
		.INIT('h15)
	) name606 (
		\pi129 ,
		_w708_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w753_,
		_w755_,
		_w756_
	);
	LUT3 #(
		.INIT('h15)
	) name608 (
		\pi099 ,
		_w707_,
		_w708_,
		_w757_
	);
	LUT4 #(
		.INIT('h0080)
	) name609 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi141 ,
		_w758_
	);
	LUT3 #(
		.INIT('h15)
	) name610 (
		\pi129 ,
		_w708_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		_w757_,
		_w759_,
		_w760_
	);
	LUT4 #(
		.INIT('h8000)
	) name612 (
		\pi131 ,
		\pi132 ,
		\pi133 ,
		\pi144 ,
		_w761_
	);
	LUT3 #(
		.INIT('h40)
	) name613 (
		\pi129 ,
		_w733_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h2)
	) name614 (
		\pi100 ,
		\pi129 ,
		_w763_
	);
	LUT4 #(
		.INIT('h7200)
	) name615 (
		_w707_,
		_w733_,
		_w739_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('he)
	) name616 (
		_w762_,
		_w764_,
		_w765_
	);
	LUT4 #(
		.INIT('h0080)
	) name617 (
		\pi037 ,
		\pi136 ,
		\pi137 ,
		\pi138 ,
		_w766_
	);
	LUT3 #(
		.INIT('h32)
	) name618 (
		\pi082 ,
		\pi136 ,
		\pi138 ,
		_w767_
	);
	LUT3 #(
		.INIT('h8c)
	) name619 (
		\pi096 ,
		\pi137 ,
		\pi138 ,
		_w768_
	);
	LUT3 #(
		.INIT('h15)
	) name620 (
		_w766_,
		_w767_,
		_w768_,
		_w769_
	);
	LUT4 #(
		.INIT('hc050)
	) name621 (
		\pi065 ,
		\pi093 ,
		\pi136 ,
		\pi138 ,
		_w770_
	);
	LUT4 #(
		.INIT('h0c05)
	) name622 (
		\pi077 ,
		\pi124 ,
		\pi136 ,
		\pi138 ,
		_w771_
	);
	LUT3 #(
		.INIT('h54)
	) name623 (
		\pi137 ,
		_w770_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('hd)
	) name624 (
		_w769_,
		_w772_,
		_w773_
	);
	LUT4 #(
		.INIT('hf35f)
	) name625 (
		\pi091 ,
		\pi095 ,
		\pi136 ,
		\pi137 ,
		_w774_
	);
	LUT4 #(
		.INIT('hac00)
	) name626 (
		\pi034 ,
		\pi079 ,
		\pi136 ,
		\pi137 ,
		_w775_
	);
	LUT4 #(
		.INIT('h0035)
	) name627 (
		\pi066 ,
		\pi069 ,
		\pi136 ,
		\pi137 ,
		_w776_
	);
	LUT4 #(
		.INIT('h7772)
	) name628 (
		\pi138 ,
		_w774_,
		_w775_,
		_w776_,
		_w777_
	);
	LUT4 #(
		.INIT('hf35f)
	) name629 (
		\pi090 ,
		\pi094 ,
		\pi136 ,
		\pi137 ,
		_w778_
	);
	LUT4 #(
		.INIT('hac00)
	) name630 (
		\pi033 ,
		\pi078 ,
		\pi136 ,
		\pi137 ,
		_w779_
	);
	LUT4 #(
		.INIT('h0053)
	) name631 (
		\pi063 ,
		\pi074 ,
		\pi136 ,
		\pi137 ,
		_w780_
	);
	LUT4 #(
		.INIT('h7772)
	) name632 (
		\pi138 ,
		_w778_,
		_w779_,
		_w780_,
		_w781_
	);
	LUT4 #(
		.INIT('hfc5f)
	) name633 (
		\pi099 ,
		\pi112 ,
		\pi136 ,
		\pi137 ,
		_w782_
	);
	LUT4 #(
		.INIT('hac00)
	) name634 (
		\pi032 ,
		\pi084 ,
		\pi136 ,
		\pi137 ,
		_w783_
	);
	LUT4 #(
		.INIT('h0053)
	) name635 (
		\pi068 ,
		\pi073 ,
		\pi136 ,
		\pi137 ,
		_w784_
	);
	LUT4 #(
		.INIT('h7772)
	) name636 (
		\pi138 ,
		_w782_,
		_w783_,
		_w784_,
		_w785_
	);
	LUT4 #(
		.INIT('h0080)
	) name637 (
		\pi035 ,
		\pi136 ,
		\pi137 ,
		\pi138 ,
		_w786_
	);
	LUT3 #(
		.INIT('h32)
	) name638 (
		\pi080 ,
		\pi136 ,
		\pi138 ,
		_w787_
	);
	LUT3 #(
		.INIT('h8c)
	) name639 (
		\pi100 ,
		\pi137 ,
		\pi138 ,
		_w788_
	);
	LUT3 #(
		.INIT('h15)
	) name640 (
		_w786_,
		_w787_,
		_w788_,
		_w789_
	);
	LUT4 #(
		.INIT('hc050)
	) name641 (
		\pi070 ,
		\pi092 ,
		\pi136 ,
		\pi138 ,
		_w790_
	);
	LUT4 #(
		.INIT('h0c05)
	) name642 (
		\pi075 ,
		\pi125 ,
		\pi136 ,
		\pi138 ,
		_w791_
	);
	LUT3 #(
		.INIT('h54)
	) name643 (
		\pi137 ,
		_w790_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('hd)
	) name644 (
		_w789_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('h0040)
	) name645 (
		\pi003 ,
		\pi085 ,
		\pi116 ,
		\pi129 ,
		_w794_
	);
	LUT4 #(
		.INIT('h0001)
	) name646 (
		\pi026 ,
		\pi027 ,
		\pi053 ,
		\pi058 ,
		_w795_
	);
	LUT4 #(
		.INIT('h2000)
	) name647 (
		_w149_,
		_w396_,
		_w696_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('he)
	) name648 (
		_w794_,
		_w796_,
		_w797_
	);
	LUT4 #(
		.INIT('h0080)
	) name649 (
		\pi036 ,
		\pi136 ,
		\pi137 ,
		\pi138 ,
		_w798_
	);
	LUT3 #(
		.INIT('h32)
	) name650 (
		\pi081 ,
		\pi136 ,
		\pi138 ,
		_w799_
	);
	LUT3 #(
		.INIT('h8c)
	) name651 (
		\pi097 ,
		\pi137 ,
		\pi138 ,
		_w800_
	);
	LUT3 #(
		.INIT('h15)
	) name652 (
		_w798_,
		_w799_,
		_w800_,
		_w801_
	);
	LUT4 #(
		.INIT('hc050)
	) name653 (
		\pi071 ,
		\pi098 ,
		\pi136 ,
		\pi138 ,
		_w802_
	);
	LUT4 #(
		.INIT('h0a03)
	) name654 (
		\pi023 ,
		\pi076 ,
		\pi136 ,
		\pi138 ,
		_w803_
	);
	LUT3 #(
		.INIT('h54)
	) name655 (
		\pi137 ,
		_w802_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('hd)
	) name656 (
		_w801_,
		_w804_,
		_w805_
	);
	LUT4 #(
		.INIT('h0080)
	) name657 (
		\pi030 ,
		\pi136 ,
		\pi137 ,
		\pi138 ,
		_w806_
	);
	LUT3 #(
		.INIT('h32)
	) name658 (
		\pi086 ,
		\pi136 ,
		\pi138 ,
		_w807_
	);
	LUT3 #(
		.INIT('h8c)
	) name659 (
		\pi111 ,
		\pi137 ,
		\pi138 ,
		_w808_
	);
	LUT3 #(
		.INIT('h15)
	) name660 (
		_w806_,
		_w807_,
		_w808_,
		_w809_
	);
	LUT4 #(
		.INIT('hc050)
	) name661 (
		\pi064 ,
		\pi088 ,
		\pi136 ,
		\pi138 ,
		_w810_
	);
	LUT4 #(
		.INIT('h0c05)
	) name662 (
		\pi067 ,
		\pi120 ,
		\pi136 ,
		\pi138 ,
		_w811_
	);
	LUT3 #(
		.INIT('h54)
	) name663 (
		\pi137 ,
		_w810_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('hd)
	) name664 (
		_w809_,
		_w812_,
		_w813_
	);
	LUT4 #(
		.INIT('h0001)
	) name665 (
		\pi026 ,
		\pi039 ,
		\pi051 ,
		\pi052 ,
		_w814_
	);
	LUT3 #(
		.INIT('h04)
	) name666 (
		\pi003 ,
		\pi116 ,
		\pi129 ,
		_w815_
	);
	LUT3 #(
		.INIT('h20)
	) name667 (
		_w392_,
		_w814_,
		_w815_,
		_w816_
	);
	LUT3 #(
		.INIT('hd9)
	) name668 (
		\pi053 ,
		\pi058 ,
		\pi097 ,
		_w817_
	);
	LUT2 #(
		.INIT('h2)
	) name669 (
		_w815_,
		_w817_,
		_w818_
	);
	LUT4 #(
		.INIT('h4000)
	) name670 (
		\pi129 ,
		\pi131 ,
		\pi132 ,
		\pi133 ,
		_w819_
	);
	LUT4 #(
		.INIT('hca00)
	) name671 (
		\pi111 ,
		\pi139 ,
		_w733_,
		_w819_,
		_w820_
	);
	LUT4 #(
		.INIT('hc500)
	) name672 (
		\pi112 ,
		\pi141 ,
		_w733_,
		_w819_,
		_w821_
	);
	LUT3 #(
		.INIT('h10)
	) name673 (
		\pi011 ,
		\pi022 ,
		\pi054 ,
		_w822_
	);
	LUT4 #(
		.INIT('h0045)
	) name674 (
		\pi003 ,
		\pi054 ,
		\pi113 ,
		\pi129 ,
		_w823_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		_w822_,
		_w823_,
		_w824_
	);
	LUT4 #(
		.INIT('hc500)
	) name676 (
		\pi115 ,
		\pi140 ,
		_w733_,
		_w819_,
		_w825_
	);
	LUT4 #(
		.INIT('h0001)
	) name677 (
		\pi004 ,
		\pi007 ,
		\pi009 ,
		\pi012 ,
		_w826_
	);
	LUT3 #(
		.INIT('h04)
	) name678 (
		\pi003 ,
		\pi054 ,
		\pi129 ,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		_w826_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('hd)
	) name680 (
		\pi122 ,
		\pi129 ,
		_w829_
	);
	LUT3 #(
		.INIT('h0e)
	) name681 (
		\pi054 ,
		\pi118 ,
		\pi129 ,
		_w830_
	);
	LUT3 #(
		.INIT('hd0)
	) name682 (
		\pi054 ,
		_w279_,
		_w830_,
		_w831_
	);
	LUT3 #(
		.INIT('h0e)
	) name683 (
		\pi095 ,
		\pi100 ,
		\pi129 ,
		_w832_
	);
	LUT3 #(
		.INIT('h01)
	) name684 (
		\pi003 ,
		\pi110 ,
		\pi120 ,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		\pi111 ,
		\pi129 ,
		_w834_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		_w833_,
		_w834_,
		_w835_
	);
	LUT3 #(
		.INIT('h08)
	) name687 (
		\pi081 ,
		\pi120 ,
		\pi129 ,
		_w836_
	);
	LUT2 #(
		.INIT('he)
	) name688 (
		\pi129 ,
		\pi134 ,
		_w837_
	);
	LUT2 #(
		.INIT('he)
	) name689 (
		\pi129 ,
		\pi135 ,
		_w838_
	);
	LUT2 #(
		.INIT('h2)
	) name690 (
		\pi057 ,
		\pi129 ,
		_w839_
	);
	LUT4 #(
		.INIT('h00ba)
	) name691 (
		\pi003 ,
		\pi096 ,
		\pi125 ,
		\pi129 ,
		_w840_
	);
	LUT3 #(
		.INIT('h40)
	) name692 (
		\pi126 ,
		\pi132 ,
		\pi133 ,
		_w841_
	);
	assign \po000  = \pi108 ;
	assign \po001  = \pi083 ;
	assign \po002  = \pi104 ;
	assign \po003  = \pi103 ;
	assign \po004  = \pi102 ;
	assign \po005  = \pi105 ;
	assign \po006  = \pi107 ;
	assign \po007  = \pi101 ;
	assign \po008  = \pi126 ;
	assign \po009  = \pi121 ;
	assign \po010  = \pi001 ;
	assign \po011  = \pi000 ;
	assign \po012  = 1'b1;
	assign \po013  = \pi130 ;
	assign \po014  = \pi128 ;
	assign \po015  = _w174_ ;
	assign \po016  = _w197_ ;
	assign \po017  = _w221_ ;
	assign \po018  = _w227_ ;
	assign \po019  = _w233_ ;
	assign \po020  = _w241_ ;
	assign \po021  = _w245_ ;
	assign \po022  = _w252_ ;
	assign \po023  = _w256_ ;
	assign \po024  = _w262_ ;
	assign \po025  = _w267_ ;
	assign \po026  = _w271_ ;
	assign \po027  = _w274_ ;
	assign \po028  = _w281_ ;
	assign \po029  = _w286_ ;
	assign \po030  = _w298_ ;
	assign \po031  = _w302_ ;
	assign \po032  = _w306_ ;
	assign \po033  = _w311_ ;
	assign \po034  = _w315_ ;
	assign \po035  = _w324_ ;
	assign \po036  = _w328_ ;
	assign \po037  = _w332_ ;
	assign \po038  = _w333_ ;
	assign \po039  = _w345_ ;
	assign \po040  = _w375_ ;
	assign \po041  = _w380_ ;
	assign \po042  = _w389_ ;
	assign \po043  = _w413_ ;
	assign \po044  = _w432_ ;
	assign \po045  = _w435_ ;
	assign \po046  = _w438_ ;
	assign \po047  = _w441_ ;
	assign \po048  = _w444_ ;
	assign \po049  = _w447_ ;
	assign \po050  = _w450_ ;
	assign \po051  = _w453_ ;
	assign \po052  = _w456_ ;
	assign \po053  = _w466_ ;
	assign \po054  = _w469_ ;
	assign \po055  = _w482_ ;
	assign \po056  = _w493_ ;
	assign \po057  = _w501_ ;
	assign \po058  = _w510_ ;
	assign \po059  = _w515_ ;
	assign \po060  = _w523_ ;
	assign \po061  = _w534_ ;
	assign \po062  = _w541_ ;
	assign \po063  = _w548_ ;
	assign \po064  = _w555_ ;
	assign \po065  = _w566_ ;
	assign \po066  = _w567_ ;
	assign \po067  = _w569_ ;
	assign \po068  = _w575_ ;
	assign \po069  = _w577_ ;
	assign \po070  = _w579_ ;
	assign \po071  = _w589_ ;
	assign \po072  = _w598_ ;
	assign \po073  = _w601_ ;
	assign \po074  = _w615_ ;
	assign \po075  = _w616_ ;
	assign \po076  = _w617_ ;
	assign \po077  = _w622_ ;
	assign \po078  = _w625_ ;
	assign \po079  = _w628_ ;
	assign \po080  = _w631_ ;
	assign \po081  = _w635_ ;
	assign \po082  = _w638_ ;
	assign \po083  = _w641_ ;
	assign \po084  = _w644_ ;
	assign \po085  = _w647_ ;
	assign \po086  = _w650_ ;
	assign \po087  = _w653_ ;
	assign \po088  = _w656_ ;
	assign \po089  = _w659_ ;
	assign \po090  = _w662_ ;
	assign \po091  = _w665_ ;
	assign \po092  = _w668_ ;
	assign \po093  = _w672_ ;
	assign \po094  = _w675_ ;
	assign \po095  = _w678_ ;
	assign \po096  = _w681_ ;
	assign \po097  = _w684_ ;
	assign \po098  = _w692_ ;
	assign \po099  = _w695_ ;
	assign \po100  = _w700_ ;
	assign \po101  = _w703_ ;
	assign \po102  = _w706_ ;
	assign \po103  = _w712_ ;
	assign \po104  = _w716_ ;
	assign \po105  = _w720_ ;
	assign \po106  = _w724_ ;
	assign \po107  = _w728_ ;
	assign \po108  = _w732_ ;
	assign \po109  = _w736_ ;
	assign \po110  = _w742_ ;
	assign \po111  = _w747_ ;
	assign \po112  = _w752_ ;
	assign \po113  = _w756_ ;
	assign \po114  = _w760_ ;
	assign \po115  = _w765_ ;
	assign \po116  = _w773_ ;
	assign \po117  = _w777_ ;
	assign \po118  = _w781_ ;
	assign \po119  = _w785_ ;
	assign \po120  = _w793_ ;
	assign \po121  = _w797_ ;
	assign \po122  = _w805_ ;
	assign \po123  = _w813_ ;
	assign \po124  = _w816_ ;
	assign \po125  = _w818_ ;
	assign \po126  = _w820_ ;
	assign \po127  = _w821_ ;
	assign \po128  = _w824_ ;
	assign \po129  = _w578_ ;
	assign \po130  = _w825_ ;
	assign \po131  = _w828_ ;
	assign \po132  = _w829_ ;
	assign \po133  = _w831_ ;
	assign \po134  = _w832_ ;
	assign \po135  = _w835_ ;
	assign \po136  = _w836_ ;
	assign \po137  = _w837_ ;
	assign \po138  = _w838_ ;
	assign \po139  = _w839_ ;
	assign \po140  = _w840_ ;
	assign \po141  = _w841_ ;
endmodule;