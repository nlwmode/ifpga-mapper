module top (\totalcoeffs[0] , \totalcoeffs[1] , \totalcoeffs[2] , \totalcoeffs[3] , \totalcoeffs[4] , \ctable[0] , \ctable[1] , \ctable[2] , \trailingones[0] , \trailingones[1] , \coeff_token[0] , \coeff_token[1] , \coeff_token[2] , \coeff_token[3] , \coeff_token[4] , \coeff_token[5] , \ctoken_len[0] , \ctoken_len[1] , \ctoken_len[2] , \ctoken_len[3] , \ctoken_len[4] );
	input \totalcoeffs[0]  ;
	input \totalcoeffs[1]  ;
	input \totalcoeffs[2]  ;
	input \totalcoeffs[3]  ;
	input \totalcoeffs[4]  ;
	input \ctable[0]  ;
	input \ctable[1]  ;
	input \ctable[2]  ;
	input \trailingones[0]  ;
	input \trailingones[1]  ;
	output \coeff_token[0]  ;
	output \coeff_token[1]  ;
	output \coeff_token[2]  ;
	output \coeff_token[3]  ;
	output \coeff_token[4]  ;
	output \coeff_token[5]  ;
	output \ctoken_len[0]  ;
	output \ctoken_len[1]  ;
	output \ctoken_len[2]  ;
	output \ctoken_len[3]  ;
	output \ctoken_len[4]  ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w14_ ;
	wire _w13_ ;
	wire _w12_ ;
	wire _w11_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\ctable[0] ,
		\ctable[2] ,
		_w11_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\trailingones[0] ,
		_w11_,
		_w12_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\totalcoeffs[0] ,
		\totalcoeffs[1] ,
		_w13_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\totalcoeffs[2] ,
		\trailingones[1] ,
		_w14_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		_w13_,
		_w14_,
		_w15_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w12_,
		_w15_,
		_w16_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\ctable[2] ,
		\trailingones[1] ,
		_w17_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w12_,
		_w17_,
		_w18_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\totalcoeffs[1] ,
		_w18_,
		_w19_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\totalcoeffs[1] ,
		\ctable[2] ,
		_w20_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\ctable[0] ,
		\trailingones[1] ,
		_w21_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w20_,
		_w21_,
		_w22_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w19_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\totalcoeffs[0] ,
		\totalcoeffs[2] ,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w23_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w16_,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\totalcoeffs[3] ,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\totalcoeffs[3] ,
		\ctable[0] ,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\totalcoeffs[0] ,
		\trailingones[1] ,
		_w29_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\totalcoeffs[1] ,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\totalcoeffs[1] ,
		\trailingones[1] ,
		_w31_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		_w28_,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w30_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\totalcoeffs[0] ,
		\trailingones[1] ,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\totalcoeffs[1] ,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\totalcoeffs[1] ,
		\trailingones[1] ,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\ctable[2] ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w35_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w33_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\totalcoeffs[2] ,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\totalcoeffs[2] ,
		\totalcoeffs[3] ,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\trailingones[1] ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\totalcoeffs[0] ,
		\totalcoeffs[3] ,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\totalcoeffs[1] ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\totalcoeffs[1] ,
		\totalcoeffs[3] ,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		\totalcoeffs[0] ,
		\ctable[0] ,
		_w47_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		\totalcoeffs[0] ,
		\totalcoeffs[1] ,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\totalcoeffs[2] ,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w47_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\trailingones[1] ,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w45_,
		_w46_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\ctable[2] ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w40_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\trailingones[0] ,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w27_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\ctable[1] ,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\totalcoeffs[1] ,
		_w29_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\trailingones[0] ,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w14_,
		_w48_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\totalcoeffs[3] ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\totalcoeffs[2] ,
		\trailingones[1] ,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\totalcoeffs[1] ,
		\trailingones[1] ,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		\totalcoeffs[2] ,
		\ctable[1] ,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\totalcoeffs[3] ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		_w65_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w64_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\trailingones[0] ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\totalcoeffs[1] ,
		\trailingones[0] ,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\totalcoeffs[2] ,
		\totalcoeffs[3] ,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w31_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w71_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\totalcoeffs[0] ,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w63_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w70_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\ctable[0] ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\totalcoeffs[2] ,
		_w34_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\ctable[1] ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\totalcoeffs[3] ,
		_w30_,
		_w81_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		_w79_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\ctable[0] ,
		_w80_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\totalcoeffs[0] ,
		\totalcoeffs[2] ,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w31_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\ctable[0] ,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\ctable[1] ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w29_,
		_w34_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\totalcoeffs[1] ,
		\ctable[0] ,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\totalcoeffs[2] ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w89_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w88_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\totalcoeffs[3] ,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\totalcoeffs[2] ,
		_w36_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w64_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\totalcoeffs[0] ,
		\totalcoeffs[3] ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\ctable[1] ,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w96_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w84_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w94_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\trailingones[0] ,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\trailingones[0] ,
		_w65_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		\totalcoeffs[3] ,
		_w85_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w78_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w102_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\ctable[2] ,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w58_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\totalcoeffs[4] ,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\totalcoeffs[1] ,
		\totalcoeffs[3] ,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\ctable[1] ,
		\trailingones[0] ,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\ctable[0] ,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		\totalcoeffs[4] ,
		\trailingones[0] ,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\ctable[1] ,
		\trailingones[1] ,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		_w113_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\ctable[1] ,
		\trailingones[1] ,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\totalcoeffs[4] ,
		\trailingones[1] ,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\ctable[0] ,
		\ctable[1] ,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\trailingones[0] ,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w120_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w117_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		\ctable[2] ,
		_w85_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w111_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w124_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w110_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w14_,
		_w112_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\trailingones[0] ,
		\trailingones[1] ,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w47_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		\ctable[0] ,
		\trailingones[0] ,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\ctable[1] ,
		\trailingones[1] ,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\ctable[1] ,
		\trailingones[0] ,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\totalcoeffs[0] ,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w134_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w131_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		\totalcoeffs[2] ,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\ctable[1] ,
		\trailingones[0] ,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		\totalcoeffs[0] ,
		\ctable[1] ,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\totalcoeffs[2] ,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		_w132_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w140_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		\trailingones[1] ,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w139_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\totalcoeffs[1] ,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\totalcoeffs[2] ,
		\trailingones[1] ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\totalcoeffs[0] ,
		\trailingones[0] ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\totalcoeffs[0] ,
		\trailingones[0] ,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w64_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w150_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		\ctable[0] ,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\totalcoeffs[0] ,
		_w134_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\trailingones[0] ,
		\trailingones[1] ,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\trailingones[0] ,
		\trailingones[1] ,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\ctable[0] ,
		\trailingones[0] ,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		\ctable[1] ,
		\trailingones[1] ,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w158_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w155_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\totalcoeffs[2] ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w154_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\totalcoeffs[1] ,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w129_,
		_w147_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\totalcoeffs[4] ,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		\totalcoeffs[2] ,
		_w13_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w114_,
		_w159_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\ctable[1] ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w119_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		_w160_,
		_w170_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w173_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w169_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\totalcoeffs[3] ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\totalcoeffs[1] ,
		\trailingones[0] ,
		_w178_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		\totalcoeffs[2] ,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\totalcoeffs[1] ,
		\trailingones[0] ,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\ctable[1] ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w179_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\totalcoeffs[3] ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\totalcoeffs[0] ,
		\trailingones[0] ,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\totalcoeffs[0] ,
		\totalcoeffs[1] ,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\totalcoeffs[1] ,
		\ctable[1] ,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\totalcoeffs[2] ,
		_w184_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w185_,
		_w186_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w187_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w183_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\ctable[0] ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		\totalcoeffs[3] ,
		\trailingones[0] ,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		\totalcoeffs[2] ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\totalcoeffs[0] ,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		\totalcoeffs[2] ,
		\trailingones[0] ,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\ctable[0] ,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\totalcoeffs[3] ,
		\trailingones[0] ,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w132_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\totalcoeffs[0] ,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w196_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		\totalcoeffs[1] ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		\totalcoeffs[2] ,
		\trailingones[0] ,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\totalcoeffs[0] ,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\totalcoeffs[0] ,
		\ctable[0] ,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w47_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w203_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		\totalcoeffs[1] ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w194_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w201_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		\ctable[1] ,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		\trailingones[1] ,
		_w191_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\totalcoeffs[1] ,
		\totalcoeffs[2] ,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\totalcoeffs[3] ,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w159_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		\totalcoeffs[1] ,
		\totalcoeffs[3] ,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w195_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w90_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		\totalcoeffs[0] ,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\ctable[0] ,
		_w214_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w41_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w219_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		\ctable[1] ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		\trailingones[1] ,
		_w215_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\totalcoeffs[4] ,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		_w212_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w177_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		\ctable[2] ,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		\ctable[1] ,
		_w28_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w36_,
		_w202_,
		_w231_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		_w79_,
		_w185_,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\totalcoeffs[2] ,
		_w13_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\trailingones[0] ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name224 (
		_w232_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w231_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		\ctable[2] ,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w15_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		\totalcoeffs[4] ,
		_w230_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		_w238_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w229_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w158_,
		_w178_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		\totalcoeffs[2] ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		\trailingones[1] ,
		_w151_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		\ctable[0] ,
		_w156_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		\ctable[0] ,
		_w64_,
		_w247_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		\totalcoeffs[1] ,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w246_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w243_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		\totalcoeffs[3] ,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w42_,
		_w180_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\ctable[0] ,
		_w216_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		\totalcoeffs[2] ,
		_w156_,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		_w252_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\totalcoeffs[0] ,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w251_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\ctable[1] ,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\ctable[1] ,
		_w31_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w36_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\trailingones[0] ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		\totalcoeffs[1] ,
		\trailingones[1] ,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w65_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		_w197_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w262_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		\totalcoeffs[2] ,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		\trailingones[0] ,
		_w14_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\totalcoeffs[2] ,
		_w263_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w180_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		\ctable[1] ,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\totalcoeffs[2] ,
		_w156_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w268_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w271_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\totalcoeffs[3] ,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w267_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		_w204_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w259_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\totalcoeffs[4] ,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		\totalcoeffs[2] ,
		_w111_,
		_w280_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		\ctable[1] ,
		\trailingones[0] ,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w157_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		\ctable[0] ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		_w280_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		\totalcoeffs[4] ,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\totalcoeffs[1] ,
		\trailingones[0] ,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		\ctable[1] ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		\trailingones[1] ,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		\totalcoeffs[2] ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		\trailingones[0] ,
		_w31_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		\totalcoeffs[3] ,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		\totalcoeffs[3] ,
		_w202_,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		\ctable[0] ,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		\totalcoeffs[2] ,
		\ctable[0] ,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		\totalcoeffs[3] ,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		\trailingones[0] ,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w294_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		\totalcoeffs[1] ,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		\ctable[0] ,
		\ctable[1] ,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		\totalcoeffs[3] ,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w178_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w299_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\trailingones[1] ,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		\totalcoeffs[3] ,
		\trailingones[1] ,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w46_,
		_w130_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		\ctable[1] ,
		_w305_,
		_w307_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\totalcoeffs[1] ,
		_w305_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w281_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\totalcoeffs[2] ,
		_w112_,
		_w311_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		\totalcoeffs[1] ,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		\ctable[0] ,
		_w193_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name303 (
		_w312_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\totalcoeffs[4] ,
		_w308_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w310_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		_w314_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w292_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		_w304_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		\totalcoeffs[0] ,
		_w285_,
		_w320_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w319_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w279_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		\ctable[2] ,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		\ctable[2] ,
		_w157_,
		_w324_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		\totalcoeffs[0] ,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w30_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w34_,
		_w178_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w326_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		\ctable[0] ,
		\ctable[1] ,
		_w329_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		\totalcoeffs[4] ,
		_w41_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w329_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h4)
	) name321 (
		_w328_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w323_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		\trailingones[1] ,
		_w300_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w286_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\totalcoeffs[3] ,
		_w65_,
		_w336_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		\totalcoeffs[1] ,
		_w295_,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		\ctable[1] ,
		_w41_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w337_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\ctable[0] ,
		\trailingones[1] ,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w156_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		\totalcoeffs[2] ,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		\totalcoeffs[3] ,
		_w281_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		\totalcoeffs[1] ,
		_w113_,
		_w345_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		\totalcoeffs[0] ,
		_w336_,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w339_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		_w346_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w186_,
		_w196_,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w301_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		\trailingones[1] ,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		\ctable[0] ,
		_w130_,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		\totalcoeffs[3] ,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		\totalcoeffs[2] ,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		\totalcoeffs[3] ,
		\trailingones[0] ,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		\ctable[1] ,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		\totalcoeffs[3] ,
		\ctable[0] ,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w357_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\ctable[0] ,
		\trailingones[0] ,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		\totalcoeffs[2] ,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\totalcoeffs[2] ,
		_w198_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		\trailingones[1] ,
		_w361_,
		_w363_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w355_,
		_w359_,
		_w365_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w364_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name356 (
		\totalcoeffs[1] ,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		\totalcoeffs[0] ,
		_w352_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w349_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		\totalcoeffs[3] ,
		\ctable[1] ,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		\totalcoeffs[2] ,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h4)
	) name362 (
		_w41_,
		_w300_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\trailingones[1] ,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w334_,
		_w371_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		\trailingones[0] ,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w375_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\totalcoeffs[1] ,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w21_,
		_w140_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		\totalcoeffs[2] ,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		\ctable[1] ,
		_w340_,
		_w382_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w263_,
		_w360_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		_w382_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w381_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\totalcoeffs[3] ,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w335_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w379_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w370_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\totalcoeffs[4] ,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		\totalcoeffs[3] ,
		\totalcoeffs[4] ,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w170_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w121_,
		_w329_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		\ctable[0] ,
		_w157_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w393_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w392_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w390_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\ctable[2] ,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		\totalcoeffs[4] ,
		_w233_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		\totalcoeffs[3] ,
		\totalcoeffs[4] ,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w391_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		_w170_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w399_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h4)
	) name393 (
		\ctable[2] ,
		_w121_,
		_w404_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		_w403_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w170_,
		_w400_,
		_w406_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w392_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		_w404_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w121_,
		_w392_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		\ctable[2] ,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h2)
	) name400 (
		\ctable[2] ,
		\trailingones[1] ,
		_w411_
	);
	LUT2 #(
		.INIT('h2)
	) name401 (
		\trailingones[0] ,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		\totalcoeffs[1] ,
		\totalcoeffs[2] ,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w412_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w95_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		\totalcoeffs[0] ,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		\totalcoeffs[1] ,
		_w244_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w156_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		\totalcoeffs[2] ,
		\ctable[2] ,
		_w419_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		_w418_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w416_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		_w230_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		\totalcoeffs[0] ,
		\totalcoeffs[2] ,
		_w423_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		_w71_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		_w66_,
		_w151_,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		\trailingones[1] ,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		\totalcoeffs[1] ,
		_w156_,
		_w428_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\totalcoeffs[0] ,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		_w36_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		\totalcoeffs[0] ,
		\ctable[1] ,
		_w431_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w178_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w213_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		_w264_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w430_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\ctable[0] ,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		_w36_,
		_w149_,
		_w437_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w204_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w427_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		_w436_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		\totalcoeffs[3] ,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		\totalcoeffs[1] ,
		\ctable[0] ,
		_w442_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		\totalcoeffs[2] ,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		_w115_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		\ctable[0] ,
		_w263_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w444_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		\totalcoeffs[0] ,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w21_,
		_w423_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w447_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		\trailingones[0] ,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\trailingones[1] ,
		_w423_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w103_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		\ctable[0] ,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		\totalcoeffs[2] ,
		\trailingones[0] ,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w195_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w64_,
		_w148_,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		\ctable[1] ,
		_w455_,
		_w457_
	);
	LUT2 #(
		.INIT('h4)
	) name447 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w453_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w450_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		\totalcoeffs[3] ,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		\totalcoeffs[2] ,
		_w156_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w244_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		\ctable[1] ,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		\totalcoeffs[2] ,
		\ctable[0] ,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w89_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		\ctable[1] ,
		_w295_,
		_w467_
	);
	LUT2 #(
		.INIT('h2)
	) name457 (
		_w29_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w466_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		\trailingones[0] ,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		\totalcoeffs[1] ,
		_w464_,
		_w471_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		_w470_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		_w29_,
		_w454_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\trailingones[0] ,
		_w204_,
		_w474_
	);
	LUT2 #(
		.INIT('h2)
	) name464 (
		_w148_,
		_w431_,
		_w475_
	);
	LUT2 #(
		.INIT('h4)
	) name465 (
		_w474_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		\totalcoeffs[1] ,
		_w473_,
		_w477_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w476_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w472_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w441_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		_w461_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		\ctable[2] ,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w422_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		\totalcoeffs[4] ,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w410_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w115_,
		_w197_,
		_w486_
	);
	LUT2 #(
		.INIT('h2)
	) name476 (
		\totalcoeffs[3] ,
		_w157_,
		_w487_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w151_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		\ctable[1] ,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		\trailingones[0] ,
		_w305_,
		_w490_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		_w489_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		\totalcoeffs[2] ,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w184_,
		_w371_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w281_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\trailingones[1] ,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		\trailingones[0] ,
		_w133_,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		\totalcoeffs[0] ,
		_w371_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w118_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w496_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w495_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		\totalcoeffs[2] ,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w486_,
		_w492_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name492 (
		_w501_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		\totalcoeffs[1] ,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h2)
	) name494 (
		_w141_,
		_w158_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		\ctable[1] ,
		_w157_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		_w79_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w505_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h2)
	) name498 (
		\totalcoeffs[3] ,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		\totalcoeffs[0] ,
		_w195_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\ctable[1] ,
		_w151_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w510_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		\trailingones[1] ,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		\ctable[1] ,
		_w197_,
		_w514_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		_w462_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w513_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		_w509_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		\totalcoeffs[1] ,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name508 (
		\trailingones[1] ,
		_w66_,
		_w519_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		_w356_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		_w518_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w504_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		\ctable[0] ,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		\totalcoeffs[0] ,
		_w456_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		\trailingones[1] ,
		_w47_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w524_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\trailingones[0] ,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\totalcoeffs[2] ,
		_w353_,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w527_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		\totalcoeffs[3] ,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		\totalcoeffs[3] ,
		\ctable[0] ,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w14_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		\totalcoeffs[2] ,
		_w149_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w157_,
		_w532_,
		_w534_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w533_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w530_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h2)
	) name526 (
		\totalcoeffs[1] ,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		_w43_,
		_w272_,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		\totalcoeffs[2] ,
		\totalcoeffs[3] ,
		_w539_
	);
	LUT2 #(
		.INIT('h2)
	) name529 (
		_w158_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		\totalcoeffs[2] ,
		_w43_,
		_w541_
	);
	LUT2 #(
		.INIT('h2)
	) name531 (
		\ctable[0] ,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		_w540_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w538_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		\totalcoeffs[1] ,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		\trailingones[0] ,
		_w340_,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name536 (
		_w539_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w545_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		_w537_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\ctable[1] ,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w523_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		\ctable[2] ,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name542 (
		_w158_,
		_w423_,
		_w553_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		_w203_,
		_w411_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w553_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		_w28_,
		_w186_,
		_w556_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w555_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w552_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		\totalcoeffs[4] ,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		\ctable[0] ,
		\ctable[2] ,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		_w392_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name551 (
		\ctable[1] ,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w559_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		_w28_,
		_w48_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w90_,
		_w358_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		\totalcoeffs[2] ,
		_w97_,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		_w565_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w564_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h2)
	) name558 (
		\trailingones[0] ,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		\ctable[0] ,
		_w184_,
		_w570_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		_w213_,
		_w531_,
		_w571_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w570_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w569_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		\trailingones[1] ,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w295_,
		_w531_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		\totalcoeffs[1] ,
		_w293_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h4)
	) name567 (
		_w47_,
		_w202_,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w216_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w577_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h2)
	) name570 (
		\trailingones[1] ,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w264_,
		_w442_,
		_w582_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		_w72_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w65_,
		_w465_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w309_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name575 (
		\totalcoeffs[0] ,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		\totalcoeffs[2] ,
		_w65_,
		_w587_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w305_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		_w565_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w583_,
		_w586_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		\trailingones[0] ,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w574_,
		_w581_,
		_w593_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		\ctable[1] ,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w36_,
		_w184_,
		_w596_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		_w260_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		\totalcoeffs[2] ,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		\ctable[1] ,
		_w71_,
		_w599_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		_w429_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name590 (
		_w358_,
		_w598_,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		_w600_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w595_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		\ctable[2] ,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		\totalcoeffs[0] ,
		_w455_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w203_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		\trailingones[1] ,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		\trailingones[0] ,
		_w451_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		_w607_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		\totalcoeffs[1] ,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h8)
	) name600 (
		_w263_,
		_w510_,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		_w610_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		_w230_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w604_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		\totalcoeffs[4] ,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w561_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		\totalcoeffs[4] ,
		_w280_,
		_w617_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w329_,
		_w391_,
		_w618_
	);
	LUT2 #(
		.INIT('h2)
	) name608 (
		_w184_,
		_w382_,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name609 (
		\totalcoeffs[3] ,
		_w133_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w619_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		\totalcoeffs[2] ,
		_w618_,
		_w622_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w621_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		\totalcoeffs[3] ,
		_w394_,
		_w624_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		_w462_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w623_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		\totalcoeffs[1] ,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		_w372_,
		_w394_,
		_w628_
	);
	LUT2 #(
		.INIT('h2)
	) name618 (
		_w21_,
		_w184_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		\totalcoeffs[3] ,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w29_,
		_w135_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w630_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		\totalcoeffs[2] ,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		\ctable[1] ,
		_w546_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		\totalcoeffs[3] ,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		_w628_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		_w633_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name627 (
		\totalcoeffs[1] ,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h8)
	) name628 (
		_w204_,
		_w372_,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		\ctable[2] ,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w428_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		\ctable[2] ,
		_w280_,
		_w642_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		\totalcoeffs[0] ,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		\ctable[0] ,
		_w72_,
		_w644_
	);
	LUT2 #(
		.INIT('h2)
	) name634 (
		\ctable[1] ,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h2)
	) name635 (
		\ctable[2] ,
		_w72_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w617_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w645_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w643_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		_w641_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		_w627_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		_w638_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		\trailingones[0] ,
		_w30_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\totalcoeffs[2] ,
		_w400_,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name644 (
		_w35_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w653_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		_w392_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name647 (
		\ctable[2] ,
		_w329_,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name648 (
		_w657_,
		_w658_,
		_w659_
	);
	assign \coeff_token[0]  = _w128_ ;
	assign \coeff_token[1]  = _w241_ ;
	assign \coeff_token[2]  = _w333_ ;
	assign \coeff_token[3]  = _w398_ ;
	assign \coeff_token[4]  = _w405_ ;
	assign \coeff_token[5]  = _w408_ ;
	assign \ctoken_len[0]  = _w485_ ;
	assign \ctoken_len[1]  = _w563_ ;
	assign \ctoken_len[2]  = _w616_ ;
	assign \ctoken_len[3]  = _w652_ ;
	assign \ctoken_len[4]  = _w659_ ;
endmodule;