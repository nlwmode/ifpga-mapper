module top (\a0_pad , a_pad, b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad );
	input \a0_pad  ;
	input a_pad ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		c_pad,
		d_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		c_pad,
		d_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\i0_pad ,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\h0_pad ,
		_w37_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		e_pad,
		h_pad,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		e_pad,
		h_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		_w37_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		_w37_,
		_w43_,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		b_pad,
		_w44_,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		c_pad,
		g_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		d_pad,
		f_pad,
		_w49_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w48_,
		_w49_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		_w43_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w43_,
		_w52_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		b_pad,
		_w53_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		i_pad,
		j_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w47_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		_w56_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		q_pad,
		v_pad,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		p_pad,
		u_pad,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		r_pad,
		w_pad,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		t_pad,
		y_pad,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		s_pad,
		x_pad,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w60_,
		_w61_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w62_,
		_w63_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w64_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w65_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\a0_pad ,
		b_pad,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		z_pad,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w35_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		_w68_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\c0_pad ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\c0_pad ,
		\d0_pad ,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\c0_pad ,
		\d0_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w74_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w72_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\e0_pad ,
		_w75_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\e0_pad ,
		_w75_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w72_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\f0_pad ,
		_w78_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\f0_pad ,
		_w78_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w72_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\g0_pad ,
		_w78_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\f0_pad ,
		\g0_pad ,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\f0_pad ,
		\g0_pad ,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w87_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w78_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w86_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w72_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\e0_pad ,
		_w74_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\f0_pad ,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\f0_pad ,
		_w93_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\g0_pad ,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		p_pad,
		q_pad,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		s_pad,
		t_pad,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		r_pad,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		k_pad,
		p_pad,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		l_pad,
		q_pad,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w98_,
		_w100_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		q_pad,
		r_pad,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		s_pad,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		o_pad,
		t_pad,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		p_pad,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w107_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		n_pad,
		r_pad,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		s_pad,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		m_pad,
		r_pad,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		s_pad,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w112_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		p_pad,
		q_pad,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		t_pad,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w115_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w105_,
		_w110_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		_w97_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\h0_pad ,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		\a0_pad ,
		a_pad,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		s_pad,
		t_pad,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		r_pad,
		_w99_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w124_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		q_pad,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w100_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		l_pad,
		_w100_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		q_pad,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		m_pad,
		_w99_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		n_pad,
		t_pad,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		s_pad,
		_w108_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		r_pad,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w131_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w130_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		p_pad,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		p_pad,
		_w99_,
		_w139_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w106_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w138_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		k_pad,
		_w99_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w106_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\h0_pad ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w97_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w128_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w141_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w122_,
		_w123_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w147_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		q_pad,
		_w136_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w88_,
		_w93_,
		_w151_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w129_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w128_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		_w150_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		q_pad,
		_w131_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w126_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		_w135_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w100_,
		_w102_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		_w87_,
		_w93_,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w154_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		p_pad,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w89_,
		_w96_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		t_pad,
		_w101_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w107_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w164_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\i0_pad ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w163_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		\i0_pad ,
		_w143_,
		_w170_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w128_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w164_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		_w141_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		_w123_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w169_,
		_w174_,
		_w175_
	);
	assign \j0_pad  = \h0_pad ;
	assign \k0_pad  = _w40_ ;
	assign \l0_pad  = _w59_ ;
	assign \m0_pad  = _w73_ ;
	assign \n0_pad  = _w77_ ;
	assign \o0_pad  = _w81_ ;
	assign \p0_pad  = _w85_ ;
	assign \q0_pad  = _w92_ ;
	assign \r0_pad  = _w149_ ;
	assign \s0_pad  = _w175_ ;
endmodule;