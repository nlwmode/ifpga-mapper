module top (\106GAT(15)_pad , \113GAT(16)_pad , \120GAT(17)_pad , \127GAT(18)_pad , \134GAT(19)_pad , \141GAT(20)_pad , \148GAT(21)_pad , \155GAT(22)_pad , \15GAT(2)_pad , \162GAT(23)_pad , \169GAT(24)_pad , \176GAT(25)_pad , \183GAT(26)_pad , \190GAT(27)_pad , \197GAT(28)_pad , \1GAT(0)_pad , \204GAT(29)_pad , \211GAT(30)_pad , \218GAT(31)_pad , \225GAT(32)_pad , \226GAT(33)_pad , \227GAT(34)_pad , \228GAT(35)_pad , \229GAT(36)_pad , \22GAT(3)_pad , \230GAT(37)_pad , \231GAT(38)_pad , \232GAT(39)_pad , \233GAT(40)_pad , \29GAT(4)_pad , \36GAT(5)_pad , \43GAT(6)_pad , \50GAT(7)_pad , \57GAT(8)_pad , \64GAT(9)_pad , \71GAT(10)_pad , \78GAT(11)_pad , \85GAT(12)_pad , \8GAT(1)_pad , \92GAT(13)_pad , \99GAT(14)_pad , \1324GAT(583)_pad , \1325GAT(579)_pad , \1326GAT(575)_pad , \1327GAT(571)_pad , \1328GAT(584)_pad , \1329GAT(580)_pad , \1330GAT(576)_pad , \1331GAT(572)_pad , \1332GAT(585)_pad , \1333GAT(581)_pad , \1334GAT(577)_pad , \1335GAT(573)_pad , \1336GAT(586)_pad , \1337GAT(582)_pad , \1338GAT(578)_pad , \1339GAT(574)_pad , \1340GAT(567)_pad , \1341GAT(563)_pad , \1342GAT(559)_pad , \1343GAT(555)_pad , \1344GAT(568)_pad , \1345GAT(564)_pad , \1346GAT(560)_pad , \1347GAT(556)_pad , \1348GAT(569)_pad , \1349GAT(565)_pad , \1350GAT(561)_pad , \1351GAT(557)_pad , \1352GAT(570)_pad , \1353GAT(566)_pad , \1354GAT(562)_pad , \1355GAT(558)_pad );
	input \106GAT(15)_pad  ;
	input \113GAT(16)_pad  ;
	input \120GAT(17)_pad  ;
	input \127GAT(18)_pad  ;
	input \134GAT(19)_pad  ;
	input \141GAT(20)_pad  ;
	input \148GAT(21)_pad  ;
	input \155GAT(22)_pad  ;
	input \15GAT(2)_pad  ;
	input \162GAT(23)_pad  ;
	input \169GAT(24)_pad  ;
	input \176GAT(25)_pad  ;
	input \183GAT(26)_pad  ;
	input \190GAT(27)_pad  ;
	input \197GAT(28)_pad  ;
	input \1GAT(0)_pad  ;
	input \204GAT(29)_pad  ;
	input \211GAT(30)_pad  ;
	input \218GAT(31)_pad  ;
	input \225GAT(32)_pad  ;
	input \226GAT(33)_pad  ;
	input \227GAT(34)_pad  ;
	input \228GAT(35)_pad  ;
	input \229GAT(36)_pad  ;
	input \22GAT(3)_pad  ;
	input \230GAT(37)_pad  ;
	input \231GAT(38)_pad  ;
	input \232GAT(39)_pad  ;
	input \233GAT(40)_pad  ;
	input \29GAT(4)_pad  ;
	input \36GAT(5)_pad  ;
	input \43GAT(6)_pad  ;
	input \50GAT(7)_pad  ;
	input \57GAT(8)_pad  ;
	input \64GAT(9)_pad  ;
	input \71GAT(10)_pad  ;
	input \78GAT(11)_pad  ;
	input \85GAT(12)_pad  ;
	input \8GAT(1)_pad  ;
	input \92GAT(13)_pad  ;
	input \99GAT(14)_pad  ;
	output \1324GAT(583)_pad  ;
	output \1325GAT(579)_pad  ;
	output \1326GAT(575)_pad  ;
	output \1327GAT(571)_pad  ;
	output \1328GAT(584)_pad  ;
	output \1329GAT(580)_pad  ;
	output \1330GAT(576)_pad  ;
	output \1331GAT(572)_pad  ;
	output \1332GAT(585)_pad  ;
	output \1333GAT(581)_pad  ;
	output \1334GAT(577)_pad  ;
	output \1335GAT(573)_pad  ;
	output \1336GAT(586)_pad  ;
	output \1337GAT(582)_pad  ;
	output \1338GAT(578)_pad  ;
	output \1339GAT(574)_pad  ;
	output \1340GAT(567)_pad  ;
	output \1341GAT(563)_pad  ;
	output \1342GAT(559)_pad  ;
	output \1343GAT(555)_pad  ;
	output \1344GAT(568)_pad  ;
	output \1345GAT(564)_pad  ;
	output \1346GAT(560)_pad  ;
	output \1347GAT(556)_pad  ;
	output \1348GAT(569)_pad  ;
	output \1349GAT(565)_pad  ;
	output \1350GAT(561)_pad  ;
	output \1351GAT(557)_pad  ;
	output \1352GAT(570)_pad  ;
	output \1353GAT(566)_pad  ;
	output \1354GAT(562)_pad  ;
	output \1355GAT(558)_pad  ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	LUT4 #(
		.INIT('h9669)
	) name0 (
		\169GAT(24)_pad ,
		\176GAT(25)_pad ,
		\183GAT(26)_pad ,
		\190GAT(27)_pad ,
		_w43_
	);
	LUT3 #(
		.INIT('h87)
	) name1 (
		\226GAT(33)_pad ,
		\233GAT(40)_pad ,
		\64GAT(9)_pad ,
		_w44_
	);
	LUT2 #(
		.INIT('h9)
	) name2 (
		\36GAT(5)_pad ,
		\8GAT(1)_pad ,
		_w45_
	);
	LUT3 #(
		.INIT('h96)
	) name3 (
		_w43_,
		_w44_,
		_w45_,
		_w46_
	);
	LUT4 #(
		.INIT('h6996)
	) name4 (
		\197GAT(28)_pad ,
		\204GAT(29)_pad ,
		\211GAT(30)_pad ,
		\218GAT(31)_pad ,
		_w47_
	);
	LUT2 #(
		.INIT('h9)
	) name5 (
		\92GAT(13)_pad ,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h6)
	) name6 (
		_w46_,
		_w48_,
		_w49_
	);
	LUT4 #(
		.INIT('h9669)
	) name7 (
		\113GAT(16)_pad ,
		\120GAT(17)_pad ,
		\127GAT(18)_pad ,
		\134GAT(19)_pad ,
		_w50_
	);
	LUT4 #(
		.INIT('h6a95)
	) name8 (
		\15GAT(2)_pad ,
		\227GAT(34)_pad ,
		\233GAT(40)_pad ,
		\43GAT(6)_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h9)
	) name9 (
		\71GAT(10)_pad ,
		\99GAT(14)_pad ,
		_w52_
	);
	LUT4 #(
		.INIT('h6996)
	) name10 (
		_w43_,
		_w50_,
		_w51_,
		_w52_,
		_w53_
	);
	LUT3 #(
		.INIT('h87)
	) name11 (
		\225GAT(32)_pad ,
		\233GAT(40)_pad ,
		\57GAT(8)_pad ,
		_w54_
	);
	LUT2 #(
		.INIT('h9)
	) name12 (
		\1GAT(0)_pad ,
		\29GAT(4)_pad ,
		_w55_
	);
	LUT3 #(
		.INIT('h96)
	) name13 (
		_w50_,
		_w54_,
		_w55_,
		_w56_
	);
	LUT4 #(
		.INIT('h9669)
	) name14 (
		\141GAT(20)_pad ,
		\148GAT(21)_pad ,
		\155GAT(22)_pad ,
		\162GAT(23)_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h9)
	) name15 (
		\85GAT(12)_pad ,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\228GAT(35)_pad ,
		\233GAT(40)_pad ,
		_w59_
	);
	LUT4 #(
		.INIT('h9669)
	) name17 (
		\106GAT(15)_pad ,
		\22GAT(3)_pad ,
		\50GAT(7)_pad ,
		\78GAT(11)_pad ,
		_w60_
	);
	LUT4 #(
		.INIT('h9669)
	) name18 (
		_w47_,
		_w57_,
		_w59_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h60)
	) name19 (
		_w56_,
		_w58_,
		_w61_,
		_w62_
	);
	LUT3 #(
		.INIT('h90)
	) name20 (
		_w56_,
		_w58_,
		_w61_,
		_w63_
	);
	LUT4 #(
		.INIT('h8e9f)
	) name21 (
		_w49_,
		_w53_,
		_w62_,
		_w63_,
		_w64_
	);
	LUT4 #(
		.INIT('h0990)
	) name22 (
		_w46_,
		_w48_,
		_w56_,
		_w58_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w53_,
		_w61_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w65_,
		_w66_,
		_w67_
	);
	LUT4 #(
		.INIT('h9669)
	) name25 (
		\106GAT(15)_pad ,
		\85GAT(12)_pad ,
		\92GAT(13)_pad ,
		\99GAT(14)_pad ,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\230GAT(37)_pad ,
		\233GAT(40)_pad ,
		_w69_
	);
	LUT2 #(
		.INIT('h9)
	) name27 (
		_w68_,
		_w69_,
		_w70_
	);
	LUT4 #(
		.INIT('h9669)
	) name28 (
		\57GAT(8)_pad ,
		\64GAT(9)_pad ,
		\71GAT(10)_pad ,
		\78GAT(11)_pad ,
		_w71_
	);
	LUT2 #(
		.INIT('h6)
	) name29 (
		\120GAT(17)_pad ,
		\148GAT(21)_pad ,
		_w72_
	);
	LUT2 #(
		.INIT('h9)
	) name30 (
		\176GAT(25)_pad ,
		\204GAT(29)_pad ,
		_w73_
	);
	LUT3 #(
		.INIT('h69)
	) name31 (
		_w71_,
		_w72_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h6)
	) name32 (
		_w70_,
		_w74_,
		_w75_
	);
	LUT4 #(
		.INIT('h9669)
	) name33 (
		\29GAT(4)_pad ,
		\36GAT(5)_pad ,
		\43GAT(6)_pad ,
		\50GAT(7)_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h9)
	) name34 (
		\113GAT(16)_pad ,
		\141GAT(20)_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h9)
	) name35 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT4 #(
		.INIT('h9669)
	) name36 (
		\15GAT(2)_pad ,
		\1GAT(0)_pad ,
		\22GAT(3)_pad ,
		\8GAT(1)_pad ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\229GAT(36)_pad ,
		\233GAT(40)_pad ,
		_w80_
	);
	LUT2 #(
		.INIT('h9)
	) name38 (
		\169GAT(24)_pad ,
		\197GAT(28)_pad ,
		_w81_
	);
	LUT3 #(
		.INIT('h69)
	) name39 (
		_w79_,
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h6)
	) name40 (
		_w78_,
		_w82_,
		_w83_
	);
	LUT4 #(
		.INIT('h0660)
	) name41 (
		_w70_,
		_w74_,
		_w78_,
		_w82_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\232GAT(39)_pad ,
		\233GAT(40)_pad ,
		_w85_
	);
	LUT4 #(
		.INIT('h9669)
	) name43 (
		\134GAT(19)_pad ,
		\162GAT(23)_pad ,
		\190GAT(27)_pad ,
		\218GAT(31)_pad ,
		_w86_
	);
	LUT4 #(
		.INIT('h9669)
	) name44 (
		_w68_,
		_w76_,
		_w85_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\231GAT(38)_pad ,
		\233GAT(40)_pad ,
		_w88_
	);
	LUT4 #(
		.INIT('h6996)
	) name46 (
		\127GAT(18)_pad ,
		\155GAT(22)_pad ,
		\183GAT(26)_pad ,
		\211GAT(30)_pad ,
		_w89_
	);
	LUT4 #(
		.INIT('h9669)
	) name47 (
		_w71_,
		_w79_,
		_w88_,
		_w89_,
		_w90_
	);
	LUT4 #(
		.INIT('h0009)
	) name48 (
		_w56_,
		_w58_,
		_w87_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w84_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('h59aa)
	) name50 (
		\1GAT(0)_pad ,
		_w64_,
		_w67_,
		_w92_,
		_w93_
	);
	LUT4 #(
		.INIT('h0006)
	) name51 (
		_w46_,
		_w48_,
		_w87_,
		_w90_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w84_,
		_w94_,
		_w95_
	);
	LUT4 #(
		.INIT('h59aa)
	) name53 (
		\8GAT(1)_pad ,
		_w64_,
		_w67_,
		_w95_,
		_w96_
	);
	LUT3 #(
		.INIT('h02)
	) name54 (
		_w53_,
		_w87_,
		_w90_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w84_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h59aa)
	) name56 (
		\15GAT(2)_pad ,
		_w64_,
		_w67_,
		_w98_,
		_w99_
	);
	LUT3 #(
		.INIT('h01)
	) name57 (
		_w61_,
		_w87_,
		_w90_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w84_,
		_w100_,
		_w101_
	);
	LUT4 #(
		.INIT('h59aa)
	) name59 (
		\22GAT(3)_pad ,
		_w64_,
		_w67_,
		_w101_,
		_w102_
	);
	LUT3 #(
		.INIT('h90)
	) name60 (
		_w56_,
		_w58_,
		_w87_,
		_w103_
	);
	LUT3 #(
		.INIT('h80)
	) name61 (
		_w84_,
		_w90_,
		_w103_,
		_w104_
	);
	LUT4 #(
		.INIT('h59aa)
	) name62 (
		\29GAT(4)_pad ,
		_w64_,
		_w67_,
		_w104_,
		_w105_
	);
	LUT3 #(
		.INIT('h60)
	) name63 (
		_w46_,
		_w48_,
		_w87_,
		_w106_
	);
	LUT3 #(
		.INIT('h80)
	) name64 (
		_w84_,
		_w90_,
		_w106_,
		_w107_
	);
	LUT4 #(
		.INIT('h59aa)
	) name65 (
		\36GAT(5)_pad ,
		_w64_,
		_w67_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w53_,
		_w87_,
		_w109_
	);
	LUT3 #(
		.INIT('h80)
	) name67 (
		_w84_,
		_w90_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('h59aa)
	) name68 (
		\43GAT(6)_pad ,
		_w64_,
		_w67_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w61_,
		_w87_,
		_w112_
	);
	LUT3 #(
		.INIT('h80)
	) name70 (
		_w84_,
		_w90_,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('h59aa)
	) name71 (
		\50GAT(7)_pad ,
		_w64_,
		_w67_,
		_w113_,
		_w114_
	);
	LUT4 #(
		.INIT('h9009)
	) name72 (
		_w70_,
		_w74_,
		_w78_,
		_w82_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w91_,
		_w115_,
		_w116_
	);
	LUT4 #(
		.INIT('h59aa)
	) name74 (
		\57GAT(8)_pad ,
		_w64_,
		_w67_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w94_,
		_w115_,
		_w118_
	);
	LUT4 #(
		.INIT('h59aa)
	) name76 (
		\64GAT(9)_pad ,
		_w64_,
		_w67_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w97_,
		_w115_,
		_w120_
	);
	LUT4 #(
		.INIT('h59aa)
	) name78 (
		\71GAT(10)_pad ,
		_w64_,
		_w67_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w100_,
		_w115_,
		_w122_
	);
	LUT4 #(
		.INIT('h59aa)
	) name80 (
		\78GAT(11)_pad ,
		_w64_,
		_w67_,
		_w122_,
		_w123_
	);
	LUT3 #(
		.INIT('h80)
	) name81 (
		_w90_,
		_w103_,
		_w115_,
		_w124_
	);
	LUT4 #(
		.INIT('h59aa)
	) name82 (
		\85GAT(12)_pad ,
		_w64_,
		_w67_,
		_w124_,
		_w125_
	);
	LUT3 #(
		.INIT('h80)
	) name83 (
		_w90_,
		_w106_,
		_w115_,
		_w126_
	);
	LUT4 #(
		.INIT('h59aa)
	) name84 (
		\92GAT(13)_pad ,
		_w64_,
		_w67_,
		_w126_,
		_w127_
	);
	LUT3 #(
		.INIT('h80)
	) name85 (
		_w90_,
		_w109_,
		_w115_,
		_w128_
	);
	LUT4 #(
		.INIT('h59aa)
	) name86 (
		\99GAT(14)_pad ,
		_w64_,
		_w67_,
		_w128_,
		_w129_
	);
	LUT3 #(
		.INIT('h80)
	) name87 (
		_w90_,
		_w112_,
		_w115_,
		_w130_
	);
	LUT4 #(
		.INIT('h59aa)
	) name88 (
		\106GAT(15)_pad ,
		_w64_,
		_w67_,
		_w130_,
		_w131_
	);
	LUT4 #(
		.INIT('hf6fd)
	) name89 (
		_w75_,
		_w83_,
		_w87_,
		_w90_,
		_w132_
	);
	LUT4 #(
		.INIT('h6006)
	) name90 (
		_w70_,
		_w74_,
		_w78_,
		_w82_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w87_,
		_w90_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w53_,
		_w61_,
		_w136_
	);
	LUT4 #(
		.INIT('h9009)
	) name94 (
		_w46_,
		_w48_,
		_w56_,
		_w58_,
		_w137_
	);
	LUT3 #(
		.INIT('h80)
	) name95 (
		_w83_,
		_w136_,
		_w137_,
		_w138_
	);
	LUT4 #(
		.INIT('h59aa)
	) name96 (
		\113GAT(16)_pad ,
		_w132_,
		_w135_,
		_w138_,
		_w139_
	);
	LUT3 #(
		.INIT('h40)
	) name97 (
		_w75_,
		_w136_,
		_w137_,
		_w140_
	);
	LUT4 #(
		.INIT('h59aa)
	) name98 (
		\120GAT(17)_pad ,
		_w132_,
		_w135_,
		_w140_,
		_w141_
	);
	LUT3 #(
		.INIT('h40)
	) name99 (
		_w90_,
		_w136_,
		_w137_,
		_w142_
	);
	LUT4 #(
		.INIT('h59aa)
	) name100 (
		\127GAT(18)_pad ,
		_w132_,
		_w135_,
		_w142_,
		_w143_
	);
	LUT3 #(
		.INIT('h80)
	) name101 (
		_w87_,
		_w136_,
		_w137_,
		_w144_
	);
	LUT4 #(
		.INIT('h59aa)
	) name102 (
		\134GAT(19)_pad ,
		_w132_,
		_w135_,
		_w144_,
		_w145_
	);
	LUT3 #(
		.INIT('h14)
	) name103 (
		_w61_,
		_w78_,
		_w82_,
		_w146_
	);
	LUT3 #(
		.INIT('h40)
	) name104 (
		_w53_,
		_w137_,
		_w146_,
		_w147_
	);
	LUT4 #(
		.INIT('h59aa)
	) name105 (
		\141GAT(20)_pad ,
		_w132_,
		_w135_,
		_w147_,
		_w148_
	);
	LUT3 #(
		.INIT('h41)
	) name106 (
		_w61_,
		_w70_,
		_w74_,
		_w149_
	);
	LUT3 #(
		.INIT('h40)
	) name107 (
		_w53_,
		_w137_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h59aa)
	) name108 (
		\148GAT(21)_pad ,
		_w132_,
		_w135_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w61_,
		_w90_,
		_w152_
	);
	LUT3 #(
		.INIT('h40)
	) name110 (
		_w53_,
		_w137_,
		_w152_,
		_w153_
	);
	LUT4 #(
		.INIT('h59aa)
	) name111 (
		\155GAT(22)_pad ,
		_w132_,
		_w135_,
		_w153_,
		_w154_
	);
	LUT3 #(
		.INIT('h40)
	) name112 (
		_w53_,
		_w112_,
		_w137_,
		_w155_
	);
	LUT4 #(
		.INIT('h59aa)
	) name113 (
		\162GAT(23)_pad ,
		_w132_,
		_w135_,
		_w155_,
		_w156_
	);
	LUT4 #(
		.INIT('h0660)
	) name114 (
		_w46_,
		_w48_,
		_w56_,
		_w58_,
		_w157_
	);
	LUT3 #(
		.INIT('h80)
	) name115 (
		_w83_,
		_w136_,
		_w157_,
		_w158_
	);
	LUT4 #(
		.INIT('h59aa)
	) name116 (
		\169GAT(24)_pad ,
		_w132_,
		_w135_,
		_w158_,
		_w159_
	);
	LUT3 #(
		.INIT('h40)
	) name117 (
		_w75_,
		_w136_,
		_w157_,
		_w160_
	);
	LUT4 #(
		.INIT('h59aa)
	) name118 (
		\176GAT(25)_pad ,
		_w132_,
		_w135_,
		_w160_,
		_w161_
	);
	LUT3 #(
		.INIT('h40)
	) name119 (
		_w90_,
		_w136_,
		_w157_,
		_w162_
	);
	LUT4 #(
		.INIT('h59aa)
	) name120 (
		\183GAT(26)_pad ,
		_w132_,
		_w135_,
		_w162_,
		_w163_
	);
	LUT3 #(
		.INIT('h80)
	) name121 (
		_w87_,
		_w136_,
		_w157_,
		_w164_
	);
	LUT4 #(
		.INIT('h59aa)
	) name122 (
		\190GAT(27)_pad ,
		_w132_,
		_w135_,
		_w164_,
		_w165_
	);
	LUT3 #(
		.INIT('h40)
	) name123 (
		_w53_,
		_w146_,
		_w157_,
		_w166_
	);
	LUT4 #(
		.INIT('h59aa)
	) name124 (
		\197GAT(28)_pad ,
		_w132_,
		_w135_,
		_w166_,
		_w167_
	);
	LUT3 #(
		.INIT('h40)
	) name125 (
		_w53_,
		_w149_,
		_w157_,
		_w168_
	);
	LUT4 #(
		.INIT('h59aa)
	) name126 (
		\204GAT(29)_pad ,
		_w132_,
		_w135_,
		_w168_,
		_w169_
	);
	LUT3 #(
		.INIT('h40)
	) name127 (
		_w53_,
		_w152_,
		_w157_,
		_w170_
	);
	LUT4 #(
		.INIT('h59aa)
	) name128 (
		\211GAT(30)_pad ,
		_w132_,
		_w135_,
		_w170_,
		_w171_
	);
	LUT3 #(
		.INIT('h40)
	) name129 (
		_w53_,
		_w112_,
		_w157_,
		_w172_
	);
	LUT4 #(
		.INIT('h59aa)
	) name130 (
		\218GAT(31)_pad ,
		_w132_,
		_w135_,
		_w172_,
		_w173_
	);
	assign \1324GAT(583)_pad  = _w93_ ;
	assign \1325GAT(579)_pad  = _w96_ ;
	assign \1326GAT(575)_pad  = _w99_ ;
	assign \1327GAT(571)_pad  = _w102_ ;
	assign \1328GAT(584)_pad  = _w105_ ;
	assign \1329GAT(580)_pad  = _w108_ ;
	assign \1330GAT(576)_pad  = _w111_ ;
	assign \1331GAT(572)_pad  = _w114_ ;
	assign \1332GAT(585)_pad  = _w117_ ;
	assign \1333GAT(581)_pad  = _w119_ ;
	assign \1334GAT(577)_pad  = _w121_ ;
	assign \1335GAT(573)_pad  = _w123_ ;
	assign \1336GAT(586)_pad  = _w125_ ;
	assign \1337GAT(582)_pad  = _w127_ ;
	assign \1338GAT(578)_pad  = _w129_ ;
	assign \1339GAT(574)_pad  = _w131_ ;
	assign \1340GAT(567)_pad  = _w139_ ;
	assign \1341GAT(563)_pad  = _w141_ ;
	assign \1342GAT(559)_pad  = _w143_ ;
	assign \1343GAT(555)_pad  = _w145_ ;
	assign \1344GAT(568)_pad  = _w148_ ;
	assign \1345GAT(564)_pad  = _w151_ ;
	assign \1346GAT(560)_pad  = _w154_ ;
	assign \1347GAT(556)_pad  = _w156_ ;
	assign \1348GAT(569)_pad  = _w159_ ;
	assign \1349GAT(565)_pad  = _w161_ ;
	assign \1350GAT(561)_pad  = _w163_ ;
	assign \1351GAT(557)_pad  = _w165_ ;
	assign \1352GAT(570)_pad  = _w167_ ;
	assign \1353GAT(566)_pad  = _w169_ ;
	assign \1354GAT(562)_pad  = _w171_ ;
	assign \1355GAT(558)_pad  = _w173_ ;
endmodule;