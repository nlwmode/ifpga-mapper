module top( ACCRPY_pad , \BULL0_pad  , \BULL1_pad  , \BULL2_pad  , \BULL3_pad  , \BULL4_pad  , \BULL5_pad  , \BULL6_pad  , CAPSD_pad , \CAT0_pad  , \CAT1_pad  , \CAT2_pad  , \CAT3_pad  , \CAT4_pad  , \CAT5_pad  , COMPPAR_pad , \DEL1_pad  , END_pad , FBI_pad , \IBT0_pad  , \IBT1_pad  , \IBT2_pad  , ICLR_pad , KBG_N_pad , LSD_pad , MARSSR_pad , MMERR_pad , ORWD_N_pad , OVACC_pad , OWL_N_pad , \PLUTO0_pad  , \PLUTO1_pad  , \PLUTO2_pad  , \PLUTO3_pad  , \PLUTO4_pad  , \PLUTO5_pad  , PY_pad , RATR_pad , SDO_pad , \STAR0_pad  , \STAR1_pad  , \STAR2_pad  , \STAR3_pad  , VACC_pad , VERR_N_pad , VLENESR_pad , \VST1_pad  , VSUMESR_pad , WATCH_pad , ACCRPY_P_pad , \BULL0_P_pad  , \BULL1_P_pad  , \BULL2_P_pad  , \BULL3_P_pad  , \BULL4_P_pad  , \BULL5_P_pad  , \BULL6_P_pad  , COMPPAR_P_pad , \DEL1_P_pad  , END_P_pad , KBG_F_pad , LSD_P_pad , MARSSR_P_pad , ORWD_F_pad , OVACC_P_pad , OWL_F_pad , \PLUTO0_P_pad  , \PLUTO1_P_pad  , \PLUTO2_P_pad  , \PLUTO3_P_pad  , \PLUTO4_P_pad  , \PLUTO5_P_pad  , PY_P_pad , RATR_P_pad , \STAR0_P_pad  , \STAR1_P_pad  , \STAR2_P_pad  , \STAR3_P_pad  , VERR_F_pad , VLENESR_P_pad , \VST0_P_pad  , \VST1_P_pad  , VSUMESR_P_pad , WATCH_P_pad , \n1022  );
  input ACCRPY_pad ;
  input \BULL0_pad  ;
  input \BULL1_pad  ;
  input \BULL2_pad  ;
  input \BULL3_pad  ;
  input \BULL4_pad  ;
  input \BULL5_pad  ;
  input \BULL6_pad  ;
  input CAPSD_pad ;
  input \CAT0_pad  ;
  input \CAT1_pad  ;
  input \CAT2_pad  ;
  input \CAT3_pad  ;
  input \CAT4_pad  ;
  input \CAT5_pad  ;
  input COMPPAR_pad ;
  input \DEL1_pad  ;
  input END_pad ;
  input FBI_pad ;
  input \IBT0_pad  ;
  input \IBT1_pad  ;
  input \IBT2_pad  ;
  input ICLR_pad ;
  input KBG_N_pad ;
  input LSD_pad ;
  input MARSSR_pad ;
  input MMERR_pad ;
  input ORWD_N_pad ;
  input OVACC_pad ;
  input OWL_N_pad ;
  input \PLUTO0_pad  ;
  input \PLUTO1_pad  ;
  input \PLUTO2_pad  ;
  input \PLUTO3_pad  ;
  input \PLUTO4_pad  ;
  input \PLUTO5_pad  ;
  input PY_pad ;
  input RATR_pad ;
  input SDO_pad ;
  input \STAR0_pad  ;
  input \STAR1_pad  ;
  input \STAR2_pad  ;
  input \STAR3_pad  ;
  input VACC_pad ;
  input VERR_N_pad ;
  input VLENESR_pad ;
  input \VST1_pad  ;
  input VSUMESR_pad ;
  input WATCH_pad ;
  output ACCRPY_P_pad ;
  output \BULL0_P_pad  ;
  output \BULL1_P_pad  ;
  output \BULL2_P_pad  ;
  output \BULL3_P_pad  ;
  output \BULL4_P_pad  ;
  output \BULL5_P_pad  ;
  output \BULL6_P_pad  ;
  output COMPPAR_P_pad ;
  output \DEL1_P_pad  ;
  output END_P_pad ;
  output KBG_F_pad ;
  output LSD_P_pad ;
  output MARSSR_P_pad ;
  output ORWD_F_pad ;
  output OVACC_P_pad ;
  output OWL_F_pad ;
  output \PLUTO0_P_pad  ;
  output \PLUTO1_P_pad  ;
  output \PLUTO2_P_pad  ;
  output \PLUTO3_P_pad  ;
  output \PLUTO4_P_pad  ;
  output \PLUTO5_P_pad  ;
  output PY_P_pad ;
  output RATR_P_pad ;
  output \STAR0_P_pad  ;
  output \STAR1_P_pad  ;
  output \STAR2_P_pad  ;
  output \STAR3_P_pad  ;
  output VERR_F_pad ;
  output VLENESR_P_pad ;
  output \VST0_P_pad  ;
  output \VST1_P_pad  ;
  output VSUMESR_P_pad ;
  output WATCH_P_pad ;
  output \n1022  ;
  wire n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 ;
  assign n50 = \CAT3_pad  & \IBT0_pad  ;
  assign n51 = \CAT2_pad  & ~\IBT0_pad  ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = \IBT2_pad  & WATCH_pad ;
  assign n54 = ~\IBT1_pad  & n53 ;
  assign n55 = n52 & n54 ;
  assign n56 = \CAT5_pad  & \IBT0_pad  ;
  assign n57 = \CAT4_pad  & ~\IBT0_pad  ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = \IBT1_pad  & n53 ;
  assign n60 = n58 & n59 ;
  assign n61 = ~n55 & ~n60 ;
  assign n62 = \IBT1_pad  & ~\IBT2_pad  ;
  assign n63 = \CAT1_pad  & \IBT0_pad  ;
  assign n64 = n62 & ~n63 ;
  assign n65 = \CAT0_pad  & ~\IBT0_pad  ;
  assign n66 = WATCH_pad & ~n65 ;
  assign n67 = n64 & n66 ;
  assign n68 = \STAR0_pad  & \STAR1_pad  ;
  assign n69 = FBI_pad & ~\STAR2_pad  ;
  assign n70 = n68 & n69 ;
  assign n71 = ~n67 & n70 ;
  assign n72 = n61 & n71 ;
  assign n73 = ~ACCRPY_pad & ~n72 ;
  assign n74 = OWL_N_pad & ~n73 ;
  assign n75 = \BULL0_pad  & ~WATCH_pad ;
  assign n76 = ~\BULL0_pad  & WATCH_pad ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = OWL_N_pad & ~n77 ;
  assign n79 = \BULL0_pad  & \BULL1_pad  ;
  assign n80 = WATCH_pad & n79 ;
  assign n81 = \BULL1_pad  & ~OWL_N_pad ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = OWL_N_pad & WATCH_pad ;
  assign n84 = \BULL0_pad  & n83 ;
  assign n85 = ~\BULL1_pad  & ~n84 ;
  assign n86 = n82 & ~n85 ;
  assign n87 = ~\BULL2_pad  & ~n80 ;
  assign n88 = \BULL2_pad  & WATCH_pad ;
  assign n89 = n79 & n88 ;
  assign n90 = OWL_N_pad & ~n89 ;
  assign n91 = ~n87 & n90 ;
  assign n92 = \BULL3_pad  & OWL_N_pad ;
  assign n93 = ~n89 & n92 ;
  assign n94 = ~\BULL3_pad  & OWL_N_pad ;
  assign n95 = n89 & n94 ;
  assign n96 = ~n93 & ~n95 ;
  assign n97 = \BULL3_pad  & n89 ;
  assign n98 = \BULL4_pad  & OWL_N_pad ;
  assign n99 = ~n97 & n98 ;
  assign n100 = ~\BULL4_pad  & n92 ;
  assign n101 = n89 & n100 ;
  assign n102 = ~n99 & ~n101 ;
  assign n103 = \BULL5_pad  & OWL_N_pad ;
  assign n104 = ~n97 & n103 ;
  assign n105 = \BULL4_pad  & \BULL5_pad  ;
  assign n106 = ~\BULL4_pad  & ~\BULL5_pad  ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = n92 & n107 ;
  assign n109 = n89 & n108 ;
  assign n110 = ~n104 & ~n109 ;
  assign n111 = \BULL2_pad  & \BULL3_pad  ;
  assign n112 = n105 & n111 ;
  assign n113 = \BULL6_pad  & ~n112 ;
  assign n114 = \BULL6_pad  & OWL_N_pad ;
  assign n115 = ~n80 & n114 ;
  assign n116 = ~n113 & ~n115 ;
  assign n117 = \BULL3_pad  & ~\BULL6_pad  ;
  assign n118 = n105 & n117 ;
  assign n119 = n89 & n118 ;
  assign n120 = n116 & ~n119 ;
  assign n121 = OWL_N_pad & ~n120 ;
  assign n122 = \DEL1_pad  & FBI_pad ;
  assign n123 = COMPPAR_pad & OWL_N_pad ;
  assign n124 = ~n122 & n123 ;
  assign n125 = ~COMPPAR_pad & OWL_N_pad ;
  assign n126 = n122 & n125 ;
  assign n127 = ~n124 & ~n126 ;
  assign n128 = CAPSD_pad & ~ICLR_pad ;
  assign n129 = ~END_pad & ~n72 ;
  assign n130 = OWL_N_pad & ~n129 ;
  assign n131 = n61 & ~n67 ;
  assign n132 = ~\STAR2_pad  & \STAR3_pad  ;
  assign n133 = FBI_pad & n132 ;
  assign n134 = n68 & n133 ;
  assign n135 = ~n131 & n134 ;
  assign n136 = ~\STAR2_pad  & n68 ;
  assign n137 = FBI_pad & ~n136 ;
  assign n138 = ~n67 & n137 ;
  assign n139 = n61 & n138 ;
  assign n140 = KBG_N_pad & ~n139 ;
  assign n141 = ~n135 & n140 ;
  assign n142 = OWL_N_pad & ~n141 ;
  assign n143 = LSD_pad & OWL_N_pad ;
  assign n144 = ~n134 & n143 ;
  assign n145 = FBI_pad & ~\STAR3_pad  ;
  assign n146 = ~n143 & n145 ;
  assign n147 = n136 & n146 ;
  assign n148 = n83 & n147 ;
  assign n149 = ~n144 & ~n148 ;
  assign n150 = ~\IBT1_pad  & \IBT2_pad  ;
  assign n151 = n52 & n150 ;
  assign n152 = \IBT1_pad  & \IBT2_pad  ;
  assign n153 = n58 & n152 ;
  assign n154 = ~n151 & ~n153 ;
  assign n155 = n64 & ~n65 ;
  assign n156 = ~n144 & ~n155 ;
  assign n157 = n154 & n156 ;
  assign n158 = ~n149 & ~n157 ;
  assign n159 = ~\BULL5_pad  & \BULL6_pad  ;
  assign n160 = ~\BULL3_pad  & \BULL4_pad  ;
  assign n161 = n159 & n160 ;
  assign n162 = \BULL1_pad  & ~\BULL2_pad  ;
  assign n163 = n76 & n162 ;
  assign n164 = n161 & n163 ;
  assign n165 = ~MARSSR_pad & ~n164 ;
  assign n166 = OWL_N_pad & ~n165 ;
  assign n167 = ~ICLR_pad & VACC_pad ;
  assign n168 = ~END_pad & ~ICLR_pad ;
  assign n169 = KBG_N_pad & n168 ;
  assign n170 = ~n164 & n169 ;
  assign n171 = OWL_N_pad & \PLUTO0_pad  ;
  assign n172 = ~\IBT0_pad  & OWL_N_pad ;
  assign n173 = n62 & n172 ;
  assign n174 = ~n171 & ~n173 ;
  assign n175 = KBG_N_pad & ~n164 ;
  assign n176 = ~MMERR_pad & ~SDO_pad ;
  assign n177 = COMPPAR_pad & ~\VST1_pad  ;
  assign n178 = ~n176 & n177 ;
  assign n179 = END_pad & ~n178 ;
  assign n180 = ~n171 & ~n179 ;
  assign n181 = n175 & n180 ;
  assign n182 = ~n174 & ~n181 ;
  assign n183 = OWL_N_pad & \PLUTO1_pad  ;
  assign n184 = n175 & ~n179 ;
  assign n185 = \IBT0_pad  & OWL_N_pad ;
  assign n186 = n62 & n185 ;
  assign n187 = ~n184 & n186 ;
  assign n188 = ~n183 & ~n187 ;
  assign n189 = OWL_N_pad & \PLUTO2_pad  ;
  assign n190 = \IBT2_pad  & n172 ;
  assign n191 = ~\IBT1_pad  & n190 ;
  assign n192 = ~n184 & n191 ;
  assign n193 = ~n189 & ~n192 ;
  assign n194 = OWL_N_pad & \PLUTO3_pad  ;
  assign n195 = n150 & n185 ;
  assign n196 = ~n184 & n195 ;
  assign n197 = ~n194 & ~n196 ;
  assign n198 = OWL_N_pad & \PLUTO4_pad  ;
  assign n199 = \IBT1_pad  & n190 ;
  assign n200 = ~n184 & n199 ;
  assign n201 = ~n198 & ~n200 ;
  assign n202 = OWL_N_pad & \PLUTO5_pad  ;
  assign n203 = n152 & n185 ;
  assign n204 = ~n184 & n203 ;
  assign n205 = ~n202 & ~n204 ;
  assign n206 = ~FBI_pad & PY_pad ;
  assign n207 = ~n122 & ~n206 ;
  assign n208 = ~ICLR_pad & ~n207 ;
  assign n209 = COMPPAR_pad & ~RATR_pad ;
  assign n210 = ~n176 & n209 ;
  assign n211 = ~END_pad & ~RATR_pad ;
  assign n212 = OWL_N_pad & ~n211 ;
  assign n213 = ~n210 & n212 ;
  assign n214 = ~FBI_pad & OWL_N_pad ;
  assign n215 = \STAR0_pad  & ~n214 ;
  assign n216 = ~ORWD_N_pad & \STAR0_pad  ;
  assign n217 = ~n215 & ~n216 ;
  assign n218 = ~n67 & ~n215 ;
  assign n219 = n61 & n218 ;
  assign n220 = ~n217 & ~n219 ;
  assign n221 = FBI_pad & OWL_N_pad ;
  assign n222 = ~ORWD_N_pad & OWL_N_pad ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = ~n67 & ~n221 ;
  assign n225 = n61 & n224 ;
  assign n226 = ~n223 & ~n225 ;
  assign n227 = ~\STAR0_pad  & ~n226 ;
  assign n228 = ~n220 & ~n227 ;
  assign n229 = ~FBI_pad & ORWD_N_pad ;
  assign n230 = ~FBI_pad & ~n67 ;
  assign n231 = n61 & n230 ;
  assign n232 = ~n229 & ~n231 ;
  assign n233 = n68 & n232 ;
  assign n234 = OWL_N_pad & \STAR1_pad  ;
  assign n235 = ~n220 & n234 ;
  assign n236 = ~n233 & n235 ;
  assign n237 = \STAR0_pad  & ~\STAR1_pad  ;
  assign n238 = n226 & n237 ;
  assign n239 = ~n236 & ~n238 ;
  assign n240 = OWL_N_pad & \STAR2_pad  ;
  assign n241 = ~n233 & n240 ;
  assign n242 = n136 & n226 ;
  assign n243 = ~n241 & ~n242 ;
  assign n244 = \STAR2_pad  & n68 ;
  assign n245 = n232 & n244 ;
  assign n246 = OWL_N_pad & \STAR3_pad  ;
  assign n247 = ~n245 & n246 ;
  assign n248 = OWL_N_pad & ~\STAR3_pad  ;
  assign n249 = FBI_pad & \STAR2_pad  ;
  assign n250 = n68 & n249 ;
  assign n251 = ~ORWD_N_pad & n244 ;
  assign n252 = ~n131 & n251 ;
  assign n253 = ~n250 & ~n252 ;
  assign n254 = n248 & ~n253 ;
  assign n255 = ~n247 & ~n254 ;
  assign n256 = VERR_N_pad & ~n164 ;
  assign n257 = ~n139 & n256 ;
  assign n258 = ~n135 & n257 ;
  assign n259 = OWL_N_pad & ~n258 ;
  assign n260 = KBG_N_pad & ~VLENESR_pad ;
  assign n261 = OWL_N_pad & ~n260 ;
  assign n262 = FBI_pad & ~ICLR_pad ;
  assign n263 = \VST1_pad  & n262 ;
  assign n264 = ~FBI_pad & ~ICLR_pad ;
  assign n265 = SDO_pad & n264 ;
  assign n266 = ~n263 & ~n265 ;
  assign n267 = \VST1_pad  & n264 ;
  assign n268 = PY_pad & n262 ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = END_pad & \VST1_pad  ;
  assign n271 = ~VSUMESR_pad & ~n270 ;
  assign n272 = OWL_N_pad & ~n271 ;
  assign n273 = OVACC_pad & ~VACC_pad ;
  assign n274 = ~WATCH_pad & ~n273 ;
  assign n275 = OWL_N_pad & ~n274 ;
  assign n276 = ~n67 & n136 ;
  assign n277 = n61 & n276 ;
  assign n278 = n226 & ~n277 ;
  assign ACCRPY_P_pad = n74 ;
  assign \BULL0_P_pad  = n78 ;
  assign \BULL1_P_pad  = n86 ;
  assign \BULL2_P_pad  = n91 ;
  assign \BULL3_P_pad  = ~n96 ;
  assign \BULL4_P_pad  = ~n102 ;
  assign \BULL5_P_pad  = ~n110 ;
  assign \BULL6_P_pad  = n121 ;
  assign COMPPAR_P_pad = ~n127 ;
  assign \DEL1_P_pad  = n128 ;
  assign END_P_pad = n130 ;
  assign KBG_F_pad = ~n142 ;
  assign LSD_P_pad = n158 ;
  assign MARSSR_P_pad = n166 ;
  assign ORWD_F_pad = n131 ;
  assign OVACC_P_pad = n167 ;
  assign OWL_F_pad = n170 ;
  assign \PLUTO0_P_pad  = n182 ;
  assign \PLUTO1_P_pad  = ~n188 ;
  assign \PLUTO2_P_pad  = ~n193 ;
  assign \PLUTO3_P_pad  = ~n197 ;
  assign \PLUTO4_P_pad  = ~n201 ;
  assign \PLUTO5_P_pad  = ~n205 ;
  assign PY_P_pad = n208 ;
  assign RATR_P_pad = n213 ;
  assign \STAR0_P_pad  = n228 ;
  assign \STAR1_P_pad  = ~n239 ;
  assign \STAR2_P_pad  = ~n243 ;
  assign \STAR3_P_pad  = ~n255 ;
  assign VERR_F_pad = ~n259 ;
  assign VLENESR_P_pad = n261 ;
  assign \VST0_P_pad  = ~n266 ;
  assign \VST1_P_pad  = ~n269 ;
  assign VSUMESR_P_pad = n272 ;
  assign WATCH_P_pad = n275 ;
  assign \n1022  = n278 ;
endmodule
