module top (\IC0(32)_pad , \IC1(33)_pad , \IC2(34)_pad , \IC3(35)_pad , \IC4(36)_pad , \IC5(37)_pad , \IC6(38)_pad , \IC7(39)_pad , \ID0(0)_pad , \ID1(1)_pad , \ID10(10)_pad , \ID11(11)_pad , \ID12(12)_pad , \ID13(13)_pad , \ID14(14)_pad , \ID15(15)_pad , \ID16(16)_pad , \ID17(17)_pad , \ID18(18)_pad , \ID19(19)_pad , \ID2(2)_pad , \ID20(20)_pad , \ID21(21)_pad , \ID22(22)_pad , \ID23(23)_pad , \ID24(24)_pad , \ID25(25)_pad , \ID26(26)_pad , \ID27(27)_pad , \ID28(28)_pad , \ID29(29)_pad , \ID3(3)_pad , \ID30(30)_pad , \ID31(31)_pad , \ID4(4)_pad , \ID5(5)_pad , \ID6(6)_pad , \ID7(7)_pad , \ID8(8)_pad , \ID9(9)_pad , \R(40)_pad , \OD0(242)_pad , \OD1(241)_pad , \OD10(232)_pad , \OD11(231)_pad , \OD12(230)_pad , \OD13(229)_pad , \OD14(228)_pad , \OD15(227)_pad , \OD16(226)_pad , \OD17(225)_pad , \OD18(224)_pad , \OD19(223)_pad , \OD2(240)_pad , \OD20(222)_pad , \OD21(221)_pad , \OD22(220)_pad , \OD23(219)_pad , \OD24(218)_pad , \OD25(217)_pad , \OD26(216)_pad , \OD27(215)_pad , \OD28(214)_pad , \OD29(213)_pad , \OD3(239)_pad , \OD30(212)_pad , \OD31(211)_pad , \OD4(238)_pad , \OD5(237)_pad , \OD6(236)_pad , \OD7(235)_pad , \OD8(234)_pad , \OD9(233)_pad );
	input \IC0(32)_pad  ;
	input \IC1(33)_pad  ;
	input \IC2(34)_pad  ;
	input \IC3(35)_pad  ;
	input \IC4(36)_pad  ;
	input \IC5(37)_pad  ;
	input \IC6(38)_pad  ;
	input \IC7(39)_pad  ;
	input \ID0(0)_pad  ;
	input \ID1(1)_pad  ;
	input \ID10(10)_pad  ;
	input \ID11(11)_pad  ;
	input \ID12(12)_pad  ;
	input \ID13(13)_pad  ;
	input \ID14(14)_pad  ;
	input \ID15(15)_pad  ;
	input \ID16(16)_pad  ;
	input \ID17(17)_pad  ;
	input \ID18(18)_pad  ;
	input \ID19(19)_pad  ;
	input \ID2(2)_pad  ;
	input \ID20(20)_pad  ;
	input \ID21(21)_pad  ;
	input \ID22(22)_pad  ;
	input \ID23(23)_pad  ;
	input \ID24(24)_pad  ;
	input \ID25(25)_pad  ;
	input \ID26(26)_pad  ;
	input \ID27(27)_pad  ;
	input \ID28(28)_pad  ;
	input \ID29(29)_pad  ;
	input \ID3(3)_pad  ;
	input \ID30(30)_pad  ;
	input \ID31(31)_pad  ;
	input \ID4(4)_pad  ;
	input \ID5(5)_pad  ;
	input \ID6(6)_pad  ;
	input \ID7(7)_pad  ;
	input \ID8(8)_pad  ;
	input \ID9(9)_pad  ;
	input \R(40)_pad  ;
	output \OD0(242)_pad  ;
	output \OD1(241)_pad  ;
	output \OD10(232)_pad  ;
	output \OD11(231)_pad  ;
	output \OD12(230)_pad  ;
	output \OD13(229)_pad  ;
	output \OD14(228)_pad  ;
	output \OD15(227)_pad  ;
	output \OD16(226)_pad  ;
	output \OD17(225)_pad  ;
	output \OD18(224)_pad  ;
	output \OD19(223)_pad  ;
	output \OD2(240)_pad  ;
	output \OD20(222)_pad  ;
	output \OD21(221)_pad  ;
	output \OD22(220)_pad  ;
	output \OD23(219)_pad  ;
	output \OD24(218)_pad  ;
	output \OD25(217)_pad  ;
	output \OD26(216)_pad  ;
	output \OD27(215)_pad  ;
	output \OD28(214)_pad  ;
	output \OD29(213)_pad  ;
	output \OD3(239)_pad  ;
	output \OD30(212)_pad  ;
	output \OD31(211)_pad  ;
	output \OD4(238)_pad  ;
	output \OD5(237)_pad  ;
	output \OD6(236)_pad  ;
	output \OD7(235)_pad  ;
	output \OD8(234)_pad  ;
	output \OD9(233)_pad  ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	LUT4 #(
		.INIT('h9669)
	) name0 (
		\ID20(20)_pad ,
		\ID21(21)_pad ,
		\ID22(22)_pad ,
		\ID23(23)_pad ,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\IC0(32)_pad ,
		\R(40)_pad ,
		_w44_
	);
	LUT4 #(
		.INIT('h9669)
	) name2 (
		\ID16(16)_pad ,
		\ID17(17)_pad ,
		\ID18(18)_pad ,
		\ID19(19)_pad ,
		_w45_
	);
	LUT4 #(
		.INIT('h9669)
	) name3 (
		\ID0(0)_pad ,
		\ID12(12)_pad ,
		\ID4(4)_pad ,
		\ID8(8)_pad ,
		_w46_
	);
	LUT4 #(
		.INIT('h6996)
	) name4 (
		_w43_,
		_w44_,
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\IC3(35)_pad ,
		\R(40)_pad ,
		_w48_
	);
	LUT2 #(
		.INIT('h9)
	) name6 (
		_w43_,
		_w48_,
		_w49_
	);
	LUT3 #(
		.INIT('h96)
	) name7 (
		\ID11(11)_pad ,
		\ID15(15)_pad ,
		\ID3(3)_pad ,
		_w50_
	);
	LUT4 #(
		.INIT('h9669)
	) name8 (
		\ID28(28)_pad ,
		\ID29(29)_pad ,
		\ID30(30)_pad ,
		\ID31(31)_pad ,
		_w51_
	);
	LUT3 #(
		.INIT('h96)
	) name9 (
		\ID7(7)_pad ,
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h6)
	) name10 (
		_w49_,
		_w52_,
		_w53_
	);
	LUT4 #(
		.INIT('h6996)
	) name11 (
		\ID24(24)_pad ,
		\ID25(25)_pad ,
		\ID26(26)_pad ,
		\ID27(27)_pad ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\IC2(34)_pad ,
		\R(40)_pad ,
		_w55_
	);
	LUT4 #(
		.INIT('h9669)
	) name13 (
		\ID10(10)_pad ,
		\ID14(14)_pad ,
		\ID2(2)_pad ,
		\ID6(6)_pad ,
		_w56_
	);
	LUT4 #(
		.INIT('h6996)
	) name14 (
		_w45_,
		_w54_,
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\IC1(33)_pad ,
		\R(40)_pad ,
		_w58_
	);
	LUT4 #(
		.INIT('h9669)
	) name16 (
		\ID1(1)_pad ,
		\ID13(13)_pad ,
		\ID5(5)_pad ,
		\ID9(9)_pad ,
		_w59_
	);
	LUT4 #(
		.INIT('h6996)
	) name17 (
		_w51_,
		_w58_,
		_w54_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w47_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h01)
	) name19 (
		_w47_,
		_w60_,
		_w57_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		_w47_,
		_w60_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w47_,
		_w60_,
		_w64_
	);
	LUT3 #(
		.INIT('h08)
	) name22 (
		_w47_,
		_w60_,
		_w57_,
		_w65_
	);
	LUT3 #(
		.INIT('hd6)
	) name23 (
		_w47_,
		_w60_,
		_w57_,
		_w66_
	);
	LUT3 #(
		.INIT('h09)
	) name24 (
		_w49_,
		_w52_,
		_w57_,
		_w67_
	);
	LUT4 #(
		.INIT('h31f5)
	) name25 (
		_w53_,
		_w63_,
		_w66_,
		_w67_,
		_w68_
	);
	LUT4 #(
		.INIT('h9669)
	) name26 (
		\ID4(4)_pad ,
		\ID5(5)_pad ,
		\ID6(6)_pad ,
		\ID7(7)_pad ,
		_w69_
	);
	LUT4 #(
		.INIT('h6996)
	) name27 (
		\ID12(12)_pad ,
		\ID13(13)_pad ,
		\ID14(14)_pad ,
		\ID15(15)_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h9)
	) name28 (
		\ID19(19)_pad ,
		\ID31(31)_pad ,
		_w71_
	);
	LUT3 #(
		.INIT('h93)
	) name29 (
		\IC7(39)_pad ,
		\ID27(27)_pad ,
		\R(40)_pad ,
		_w72_
	);
	LUT4 #(
		.INIT('h9669)
	) name30 (
		\ID23(23)_pad ,
		_w70_,
		_w71_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h6)
	) name31 (
		_w69_,
		_w73_,
		_w74_
	);
	LUT4 #(
		.INIT('h6996)
	) name32 (
		\ID0(0)_pad ,
		\ID1(1)_pad ,
		\ID2(2)_pad ,
		\ID3(3)_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\IC6(38)_pad ,
		\R(40)_pad ,
		_w76_
	);
	LUT4 #(
		.INIT('h9669)
	) name34 (
		\ID10(10)_pad ,
		\ID11(11)_pad ,
		\ID8(8)_pad ,
		\ID9(9)_pad ,
		_w77_
	);
	LUT4 #(
		.INIT('h9669)
	) name35 (
		\ID18(18)_pad ,
		\ID22(22)_pad ,
		\ID26(26)_pad ,
		\ID30(30)_pad ,
		_w78_
	);
	LUT4 #(
		.INIT('h9669)
	) name36 (
		_w75_,
		_w76_,
		_w77_,
		_w78_,
		_w79_
	);
	LUT3 #(
		.INIT('h09)
	) name37 (
		_w69_,
		_w73_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\IC5(37)_pad ,
		\R(40)_pad ,
		_w81_
	);
	LUT4 #(
		.INIT('h9669)
	) name39 (
		\ID17(17)_pad ,
		\ID21(21)_pad ,
		\ID25(25)_pad ,
		\ID29(29)_pad ,
		_w82_
	);
	LUT4 #(
		.INIT('h6996)
	) name40 (
		_w70_,
		_w77_,
		_w81_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\IC4(36)_pad ,
		\R(40)_pad ,
		_w84_
	);
	LUT4 #(
		.INIT('h9669)
	) name42 (
		\ID16(16)_pad ,
		\ID20(20)_pad ,
		\ID24(24)_pad ,
		\ID28(28)_pad ,
		_w85_
	);
	LUT4 #(
		.INIT('h6996)
	) name43 (
		_w69_,
		_w75_,
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w83_,
		_w86_,
		_w87_
	);
	LUT4 #(
		.INIT('h1000)
	) name45 (
		_w47_,
		_w68_,
		_w80_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h6)
	) name46 (
		\ID0(0)_pad ,
		_w88_,
		_w89_
	);
	LUT4 #(
		.INIT('h2000)
	) name47 (
		_w60_,
		_w68_,
		_w80_,
		_w87_,
		_w90_
	);
	LUT2 #(
		.INIT('h6)
	) name48 (
		\ID1(1)_pad ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		_w83_,
		_w86_,
		_w92_
	);
	LUT4 #(
		.INIT('h2000)
	) name50 (
		_w57_,
		_w68_,
		_w80_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h6)
	) name51 (
		\ID10(10)_pad ,
		_w93_,
		_w94_
	);
	LUT4 #(
		.INIT('h1000)
	) name52 (
		_w53_,
		_w68_,
		_w80_,
		_w92_,
		_w95_
	);
	LUT2 #(
		.INIT('h6)
	) name53 (
		\ID11(11)_pad ,
		_w95_,
		_w96_
	);
	LUT3 #(
		.INIT('h08)
	) name54 (
		_w79_,
		_w83_,
		_w86_,
		_w97_
	);
	LUT4 #(
		.INIT('h0400)
	) name55 (
		_w47_,
		_w74_,
		_w68_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h6)
	) name56 (
		\ID12(12)_pad ,
		_w98_,
		_w99_
	);
	LUT4 #(
		.INIT('h0800)
	) name57 (
		_w74_,
		_w60_,
		_w68_,
		_w97_,
		_w100_
	);
	LUT2 #(
		.INIT('h6)
	) name58 (
		\ID13(13)_pad ,
		_w100_,
		_w101_
	);
	LUT4 #(
		.INIT('h0800)
	) name59 (
		_w74_,
		_w57_,
		_w68_,
		_w97_,
		_w102_
	);
	LUT2 #(
		.INIT('h6)
	) name60 (
		\ID14(14)_pad ,
		_w102_,
		_w103_
	);
	LUT4 #(
		.INIT('h0200)
	) name61 (
		_w74_,
		_w53_,
		_w68_,
		_w97_,
		_w104_
	);
	LUT2 #(
		.INIT('h6)
	) name62 (
		\ID15(15)_pad ,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w83_,
		_w86_,
		_w106_
	);
	LUT3 #(
		.INIT('h20)
	) name64 (
		_w79_,
		_w83_,
		_w86_,
		_w107_
	);
	LUT3 #(
		.INIT('hd6)
	) name65 (
		_w79_,
		_w83_,
		_w86_,
		_w108_
	);
	LUT3 #(
		.INIT('h60)
	) name66 (
		_w69_,
		_w73_,
		_w79_,
		_w109_
	);
	LUT4 #(
		.INIT('h32fa)
	) name67 (
		_w74_,
		_w106_,
		_w108_,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('h60)
	) name68 (
		_w49_,
		_w52_,
		_w57_,
		_w111_
	);
	LUT4 #(
		.INIT('h0800)
	) name69 (
		_w61_,
		_w86_,
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h6)
	) name70 (
		\ID16(16)_pad ,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('h0800)
	) name71 (
		_w61_,
		_w83_,
		_w110_,
		_w111_,
		_w114_
	);
	LUT2 #(
		.INIT('h6)
	) name72 (
		\ID17(17)_pad ,
		_w114_,
		_w115_
	);
	LUT4 #(
		.INIT('h0400)
	) name73 (
		_w79_,
		_w61_,
		_w110_,
		_w111_,
		_w116_
	);
	LUT2 #(
		.INIT('h6)
	) name74 (
		\ID18(18)_pad ,
		_w116_,
		_w117_
	);
	LUT4 #(
		.INIT('h0800)
	) name75 (
		_w74_,
		_w61_,
		_w110_,
		_w111_,
		_w118_
	);
	LUT2 #(
		.INIT('h6)
	) name76 (
		\ID19(19)_pad ,
		_w118_,
		_w119_
	);
	LUT4 #(
		.INIT('h2000)
	) name77 (
		_w57_,
		_w68_,
		_w80_,
		_w87_,
		_w120_
	);
	LUT2 #(
		.INIT('h6)
	) name78 (
		\ID2(2)_pad ,
		_w120_,
		_w121_
	);
	LUT4 #(
		.INIT('h0040)
	) name79 (
		_w53_,
		_w62_,
		_w86_,
		_w110_,
		_w122_
	);
	LUT2 #(
		.INIT('h6)
	) name80 (
		\ID20(20)_pad ,
		_w122_,
		_w123_
	);
	LUT4 #(
		.INIT('h0040)
	) name81 (
		_w53_,
		_w62_,
		_w83_,
		_w110_,
		_w124_
	);
	LUT2 #(
		.INIT('h6)
	) name82 (
		\ID21(21)_pad ,
		_w124_,
		_w125_
	);
	LUT4 #(
		.INIT('h0010)
	) name83 (
		_w79_,
		_w53_,
		_w62_,
		_w110_,
		_w126_
	);
	LUT2 #(
		.INIT('h6)
	) name84 (
		\ID22(22)_pad ,
		_w126_,
		_w127_
	);
	LUT4 #(
		.INIT('h0020)
	) name85 (
		_w74_,
		_w53_,
		_w62_,
		_w110_,
		_w128_
	);
	LUT2 #(
		.INIT('h6)
	) name86 (
		\ID23(23)_pad ,
		_w128_,
		_w129_
	);
	LUT4 #(
		.INIT('h0800)
	) name87 (
		_w64_,
		_w86_,
		_w110_,
		_w111_,
		_w130_
	);
	LUT2 #(
		.INIT('h6)
	) name88 (
		\ID24(24)_pad ,
		_w130_,
		_w131_
	);
	LUT4 #(
		.INIT('h0800)
	) name89 (
		_w64_,
		_w83_,
		_w110_,
		_w111_,
		_w132_
	);
	LUT2 #(
		.INIT('h6)
	) name90 (
		\ID25(25)_pad ,
		_w132_,
		_w133_
	);
	LUT4 #(
		.INIT('h0400)
	) name91 (
		_w79_,
		_w64_,
		_w110_,
		_w111_,
		_w134_
	);
	LUT2 #(
		.INIT('h6)
	) name92 (
		\ID26(26)_pad ,
		_w134_,
		_w135_
	);
	LUT4 #(
		.INIT('h0800)
	) name93 (
		_w74_,
		_w64_,
		_w110_,
		_w111_,
		_w136_
	);
	LUT2 #(
		.INIT('h6)
	) name94 (
		\ID27(27)_pad ,
		_w136_,
		_w137_
	);
	LUT4 #(
		.INIT('h0040)
	) name95 (
		_w53_,
		_w65_,
		_w86_,
		_w110_,
		_w138_
	);
	LUT2 #(
		.INIT('h6)
	) name96 (
		\ID28(28)_pad ,
		_w138_,
		_w139_
	);
	LUT4 #(
		.INIT('h0040)
	) name97 (
		_w53_,
		_w65_,
		_w83_,
		_w110_,
		_w140_
	);
	LUT2 #(
		.INIT('h6)
	) name98 (
		\ID29(29)_pad ,
		_w140_,
		_w141_
	);
	LUT4 #(
		.INIT('h1000)
	) name99 (
		_w53_,
		_w68_,
		_w80_,
		_w87_,
		_w142_
	);
	LUT2 #(
		.INIT('h6)
	) name100 (
		\ID3(3)_pad ,
		_w142_,
		_w143_
	);
	LUT4 #(
		.INIT('h0010)
	) name101 (
		_w79_,
		_w53_,
		_w65_,
		_w110_,
		_w144_
	);
	LUT2 #(
		.INIT('h6)
	) name102 (
		\ID30(30)_pad ,
		_w144_,
		_w145_
	);
	LUT4 #(
		.INIT('h0020)
	) name103 (
		_w74_,
		_w53_,
		_w65_,
		_w110_,
		_w146_
	);
	LUT2 #(
		.INIT('h6)
	) name104 (
		\ID31(31)_pad ,
		_w146_,
		_w147_
	);
	LUT4 #(
		.INIT('h0400)
	) name105 (
		_w47_,
		_w74_,
		_w68_,
		_w107_,
		_w148_
	);
	LUT2 #(
		.INIT('h6)
	) name106 (
		\ID4(4)_pad ,
		_w148_,
		_w149_
	);
	LUT4 #(
		.INIT('h0800)
	) name107 (
		_w74_,
		_w60_,
		_w68_,
		_w107_,
		_w150_
	);
	LUT2 #(
		.INIT('h6)
	) name108 (
		\ID5(5)_pad ,
		_w150_,
		_w151_
	);
	LUT4 #(
		.INIT('h0800)
	) name109 (
		_w74_,
		_w57_,
		_w68_,
		_w107_,
		_w152_
	);
	LUT2 #(
		.INIT('h6)
	) name110 (
		\ID6(6)_pad ,
		_w152_,
		_w153_
	);
	LUT4 #(
		.INIT('h0200)
	) name111 (
		_w74_,
		_w53_,
		_w68_,
		_w107_,
		_w154_
	);
	LUT2 #(
		.INIT('h6)
	) name112 (
		\ID7(7)_pad ,
		_w154_,
		_w155_
	);
	LUT4 #(
		.INIT('h1000)
	) name113 (
		_w47_,
		_w68_,
		_w80_,
		_w92_,
		_w156_
	);
	LUT2 #(
		.INIT('h6)
	) name114 (
		\ID8(8)_pad ,
		_w156_,
		_w157_
	);
	LUT4 #(
		.INIT('h2000)
	) name115 (
		_w60_,
		_w68_,
		_w80_,
		_w92_,
		_w158_
	);
	LUT2 #(
		.INIT('h6)
	) name116 (
		\ID9(9)_pad ,
		_w158_,
		_w159_
	);
	assign \OD0(242)_pad  = _w89_ ;
	assign \OD1(241)_pad  = _w91_ ;
	assign \OD10(232)_pad  = _w94_ ;
	assign \OD11(231)_pad  = _w96_ ;
	assign \OD12(230)_pad  = _w99_ ;
	assign \OD13(229)_pad  = _w101_ ;
	assign \OD14(228)_pad  = _w103_ ;
	assign \OD15(227)_pad  = _w105_ ;
	assign \OD16(226)_pad  = _w113_ ;
	assign \OD17(225)_pad  = _w115_ ;
	assign \OD18(224)_pad  = _w117_ ;
	assign \OD19(223)_pad  = _w119_ ;
	assign \OD2(240)_pad  = _w121_ ;
	assign \OD20(222)_pad  = _w123_ ;
	assign \OD21(221)_pad  = _w125_ ;
	assign \OD22(220)_pad  = _w127_ ;
	assign \OD23(219)_pad  = _w129_ ;
	assign \OD24(218)_pad  = _w131_ ;
	assign \OD25(217)_pad  = _w133_ ;
	assign \OD26(216)_pad  = _w135_ ;
	assign \OD27(215)_pad  = _w137_ ;
	assign \OD28(214)_pad  = _w139_ ;
	assign \OD29(213)_pad  = _w141_ ;
	assign \OD3(239)_pad  = _w143_ ;
	assign \OD30(212)_pad  = _w145_ ;
	assign \OD31(211)_pad  = _w147_ ;
	assign \OD4(238)_pad  = _w149_ ;
	assign \OD5(237)_pad  = _w151_ ;
	assign \OD6(236)_pad  = _w153_ ;
	assign \OD7(235)_pad  = _w155_ ;
	assign \OD8(234)_pad  = _w157_ ;
	assign \OD9(233)_pad  = _w159_ ;
endmodule;