module top (\100(38)_pad , \103(39)_pad , \106(40)_pad , \109(41)_pad , \11(2)_pad , \112(42)_pad , \113(43)_pad , \114(44)_pad , \115(45)_pad , \116(46)_pad , \117(47)_pad , \118(48)_pad , \119(49)_pad , \120(50)_pad , \121(51)_pad , \122(52)_pad , \123(53)_pad , \126(54)_pad , \127(55)_pad , \128(56)_pad , \129(57)_pad , \130(58)_pad , \131(59)_pad , \132(60)_pad , \135(61)_pad , \136(62)_pad , \14(3)_pad , \140(64)_pad , \144(354)_pad , \145(66)_pad , \146(67)_pad , \149(68)_pad , \1497(156)_pad , \152(69)_pad , \155(70)_pad , \158(71)_pad , \161(72)_pad , \164(73)_pad , \167(74)_pad , \1689(157)_pad , \1690(158)_pad , \1691(159)_pad , \1694(160)_pad , \17(4)_pad , \170(75)_pad , \173(76)_pad , \176(77)_pad , \179(78)_pad , \182(79)_pad , \185(80)_pad , \188(81)_pad , \191(82)_pad , \194(83)_pad , \197(84)_pad , \20(5)_pad , \200(85)_pad , \203(86)_pad , \206(87)_pad , \209(88)_pad , \210(89)_pad , \217(90)_pad , \2174(161)_pad , \218(91)_pad , \225(92)_pad , \226(93)_pad , \23(6)_pad , \233(94)_pad , \234(95)_pad , \2358(162)_pad , \24(7)_pad , \241(96)_pad , \242(97)_pad , \245(98)_pad , \248(99)_pad , \25(8)_pad , \251(100)_pad , \254(101)_pad , \257(102)_pad , \26(9)_pad , \264(103)_pad , \265(104)_pad , \27(10)_pad , \272(105)_pad , \273(106)_pad , \280(107)_pad , \281(108)_pad , \2824(163)_pad , \288(109)_pad , \289(110)_pad , \292(111)_pad , \298(299)_pad , \302(114)_pad , \307(115)_pad , \308(116)_pad , \31(11)_pad , \315(117)_pad , \316(118)_pad , \323(119)_pad , \324(120)_pad , \331(121)_pad , \332(122)_pad , \335(123)_pad , \338(124)_pad , \34(12)_pad , \341(125)_pad , \348(126)_pad , \351(127)_pad , \3546(165)_pad , \3548(166)_pad , \3550(167)_pad , \3552(168)_pad , \358(128)_pad , \361(129)_pad , \366(130)_pad , \369(131)_pad , \37(13)_pad , \3717(169)_pad , \372(132)_pad , \3724(170)_pad , \373(133)_pad , \374(134)_pad , \386(135)_pad , \389(136)_pad , \4(1)_pad , \40(14)_pad , \400(137)_pad , \4087(171)_pad , \4088(172)_pad , \4089(173)_pad , \4090(174)_pad , \4091(175)_pad , \4092(176)_pad , \411(138)_pad , \4115(177)_pad , \422(139)_pad , \43(15)_pad , \435(140)_pad , \446(141)_pad , \457(142)_pad , \46(16)_pad , \468(143)_pad , \479(144)_pad , \49(17)_pad , \490(145)_pad , \503(146)_pad , \514(147)_pad , \52(18)_pad , \523(148)_pad , \53(19)_pad , \534(149)_pad , \54(20)_pad , \545(150)_pad , \552(152)_pad , \556(153)_pad , \559(154)_pad , \562(155)_pad , \61(21)_pad , \64(22)_pad , \67(23)_pad , \70(24)_pad , \73(25)_pad , \76(26)_pad , \79(27)_pad , \80(28)_pad , \81(29)_pad , \82(30)_pad , \83(31)_pad , \86(32)_pad , \87(33)_pad , \88(34)_pad , \889(734)_pad , \892(408)_pad , \91(35)_pad , \926(624)_pad , \94(36)_pad , \97(37)_pad , \973(202)_pad , \993(850)_pad , \1000(2168)_pad , \1002(1920)_pad , \1004(1977)_pad , \588(1696)_pad , \593(733)_pad , \598(1623)_pad , \599(269)_pad , \600(259)_pad , \601(220)_pad , \604(223)_pad , \606(407)_pad , \611(275)_pad , \612(263)_pad , \615(1750)_pad , \618(1925)_pad , \621(1893)_pad , \626(1752)_pad , \632(1692)_pad , \634(665)_pad , \636(1280)_pad , \639(1275)_pad , \642(2222)_pad , \645(2271)_pad , \648(2295)_pad , \651(2314)_pad , \654(2315)_pad , \656(621)_pad , \658(2483)_pad , \661(2178)_pad , \664(2223)_pad , \667(2224)_pad , \670(2225)_pad , \673(1276)_pad , \676(2229)_pad , \679(2272)_pad , \682(2296)_pad , \685(2316)_pad , \688(2317)_pad , \690(2484)_pad , \693(2179)_pad , \696(2226)_pad , \699(2227)_pad , \702(2228)_pad , \704(1281)_pad , \707(1277)_pad , \712(2297)_pad , \715(1278)_pad , \722(2131)_pad , \727(2298)_pad , \732(2300)_pad , \737(2279)_pad , \742(2238)_pad , \747(2187)_pad , \752(2189)_pad , \757(2190)_pad , \762(2184)_pad , \767(2479)_pad , \772(2299)_pad , \777(2278)_pad , \782(2239)_pad , \787(2186)_pad , \792(2188)_pad , \797(2191)_pad , \802(2183)_pad , \807(2480)_pad , \809(655)_pad , \810(356)_pad , \813(2260)_pad , \815(627)_pad , \820(1283)_pad , \822(1933)_pad , \824(2274)_pad , \826(2275)_pad , \828(2233)_pad , \830(2182)_pad , \832(2133)_pad , \834(2123)_pad , \836(2128)_pad , \838(2064)_pad , \843(2455)_pad , \845(845)_pad , \847(465)_pad , \848(330)_pad , \849(219)_pad , \850(217)_pad , \851(218)_pad , \854(2268)_pad , \859(2132)_pad , \861(2070)_pad , \863(2276)_pad , \865(2277)_pad , \867(2237)_pad , \869(2181)_pad , \871(2127)_pad , \873(2124)_pad , \875(2125)_pad , \877(2126)_pad , \882(2456)_pad , \998(2163)_pad , \u2023_syn_3 , \u2095_syn_3 , \u2109_syn_3 , \u2318_syn_3 , \u3086_syn_3 );
	input \100(38)_pad  ;
	input \103(39)_pad  ;
	input \106(40)_pad  ;
	input \109(41)_pad  ;
	input \11(2)_pad  ;
	input \112(42)_pad  ;
	input \113(43)_pad  ;
	input \114(44)_pad  ;
	input \115(45)_pad  ;
	input \116(46)_pad  ;
	input \117(47)_pad  ;
	input \118(48)_pad  ;
	input \119(49)_pad  ;
	input \120(50)_pad  ;
	input \121(51)_pad  ;
	input \122(52)_pad  ;
	input \123(53)_pad  ;
	input \126(54)_pad  ;
	input \127(55)_pad  ;
	input \128(56)_pad  ;
	input \129(57)_pad  ;
	input \130(58)_pad  ;
	input \131(59)_pad  ;
	input \132(60)_pad  ;
	input \135(61)_pad  ;
	input \136(62)_pad  ;
	input \14(3)_pad  ;
	input \140(64)_pad  ;
	input \144(354)_pad  ;
	input \145(66)_pad  ;
	input \146(67)_pad  ;
	input \149(68)_pad  ;
	input \1497(156)_pad  ;
	input \152(69)_pad  ;
	input \155(70)_pad  ;
	input \158(71)_pad  ;
	input \161(72)_pad  ;
	input \164(73)_pad  ;
	input \167(74)_pad  ;
	input \1689(157)_pad  ;
	input \1690(158)_pad  ;
	input \1691(159)_pad  ;
	input \1694(160)_pad  ;
	input \17(4)_pad  ;
	input \170(75)_pad  ;
	input \173(76)_pad  ;
	input \176(77)_pad  ;
	input \179(78)_pad  ;
	input \182(79)_pad  ;
	input \185(80)_pad  ;
	input \188(81)_pad  ;
	input \191(82)_pad  ;
	input \194(83)_pad  ;
	input \197(84)_pad  ;
	input \20(5)_pad  ;
	input \200(85)_pad  ;
	input \203(86)_pad  ;
	input \206(87)_pad  ;
	input \209(88)_pad  ;
	input \210(89)_pad  ;
	input \217(90)_pad  ;
	input \2174(161)_pad  ;
	input \218(91)_pad  ;
	input \225(92)_pad  ;
	input \226(93)_pad  ;
	input \23(6)_pad  ;
	input \233(94)_pad  ;
	input \234(95)_pad  ;
	input \2358(162)_pad  ;
	input \24(7)_pad  ;
	input \241(96)_pad  ;
	input \242(97)_pad  ;
	input \245(98)_pad  ;
	input \248(99)_pad  ;
	input \25(8)_pad  ;
	input \251(100)_pad  ;
	input \254(101)_pad  ;
	input \257(102)_pad  ;
	input \26(9)_pad  ;
	input \264(103)_pad  ;
	input \265(104)_pad  ;
	input \27(10)_pad  ;
	input \272(105)_pad  ;
	input \273(106)_pad  ;
	input \280(107)_pad  ;
	input \281(108)_pad  ;
	input \2824(163)_pad  ;
	input \288(109)_pad  ;
	input \289(110)_pad  ;
	input \292(111)_pad  ;
	input \298(299)_pad  ;
	input \302(114)_pad  ;
	input \307(115)_pad  ;
	input \308(116)_pad  ;
	input \31(11)_pad  ;
	input \315(117)_pad  ;
	input \316(118)_pad  ;
	input \323(119)_pad  ;
	input \324(120)_pad  ;
	input \331(121)_pad  ;
	input \332(122)_pad  ;
	input \335(123)_pad  ;
	input \338(124)_pad  ;
	input \34(12)_pad  ;
	input \341(125)_pad  ;
	input \348(126)_pad  ;
	input \351(127)_pad  ;
	input \3546(165)_pad  ;
	input \3548(166)_pad  ;
	input \3550(167)_pad  ;
	input \3552(168)_pad  ;
	input \358(128)_pad  ;
	input \361(129)_pad  ;
	input \366(130)_pad  ;
	input \369(131)_pad  ;
	input \37(13)_pad  ;
	input \3717(169)_pad  ;
	input \372(132)_pad  ;
	input \3724(170)_pad  ;
	input \373(133)_pad  ;
	input \374(134)_pad  ;
	input \386(135)_pad  ;
	input \389(136)_pad  ;
	input \4(1)_pad  ;
	input \40(14)_pad  ;
	input \400(137)_pad  ;
	input \4087(171)_pad  ;
	input \4088(172)_pad  ;
	input \4089(173)_pad  ;
	input \4090(174)_pad  ;
	input \4091(175)_pad  ;
	input \4092(176)_pad  ;
	input \411(138)_pad  ;
	input \4115(177)_pad  ;
	input \422(139)_pad  ;
	input \43(15)_pad  ;
	input \435(140)_pad  ;
	input \446(141)_pad  ;
	input \457(142)_pad  ;
	input \46(16)_pad  ;
	input \468(143)_pad  ;
	input \479(144)_pad  ;
	input \49(17)_pad  ;
	input \490(145)_pad  ;
	input \503(146)_pad  ;
	input \514(147)_pad  ;
	input \52(18)_pad  ;
	input \523(148)_pad  ;
	input \53(19)_pad  ;
	input \534(149)_pad  ;
	input \54(20)_pad  ;
	input \545(150)_pad  ;
	input \552(152)_pad  ;
	input \556(153)_pad  ;
	input \559(154)_pad  ;
	input \562(155)_pad  ;
	input \61(21)_pad  ;
	input \64(22)_pad  ;
	input \67(23)_pad  ;
	input \70(24)_pad  ;
	input \73(25)_pad  ;
	input \76(26)_pad  ;
	input \79(27)_pad  ;
	input \80(28)_pad  ;
	input \81(29)_pad  ;
	input \82(30)_pad  ;
	input \83(31)_pad  ;
	input \86(32)_pad  ;
	input \87(33)_pad  ;
	input \88(34)_pad  ;
	input \889(734)_pad  ;
	input \892(408)_pad  ;
	input \91(35)_pad  ;
	input \926(624)_pad  ;
	input \94(36)_pad  ;
	input \97(37)_pad  ;
	input \973(202)_pad  ;
	input \993(850)_pad  ;
	output \1000(2168)_pad  ;
	output \1002(1920)_pad  ;
	output \1004(1977)_pad  ;
	output \588(1696)_pad  ;
	output \593(733)_pad  ;
	output \598(1623)_pad  ;
	output \599(269)_pad  ;
	output \600(259)_pad  ;
	output \601(220)_pad  ;
	output \604(223)_pad  ;
	output \606(407)_pad  ;
	output \611(275)_pad  ;
	output \612(263)_pad  ;
	output \615(1750)_pad  ;
	output \618(1925)_pad  ;
	output \621(1893)_pad  ;
	output \626(1752)_pad  ;
	output \632(1692)_pad  ;
	output \634(665)_pad  ;
	output \636(1280)_pad  ;
	output \639(1275)_pad  ;
	output \642(2222)_pad  ;
	output \645(2271)_pad  ;
	output \648(2295)_pad  ;
	output \651(2314)_pad  ;
	output \654(2315)_pad  ;
	output \656(621)_pad  ;
	output \658(2483)_pad  ;
	output \661(2178)_pad  ;
	output \664(2223)_pad  ;
	output \667(2224)_pad  ;
	output \670(2225)_pad  ;
	output \673(1276)_pad  ;
	output \676(2229)_pad  ;
	output \679(2272)_pad  ;
	output \682(2296)_pad  ;
	output \685(2316)_pad  ;
	output \688(2317)_pad  ;
	output \690(2484)_pad  ;
	output \693(2179)_pad  ;
	output \696(2226)_pad  ;
	output \699(2227)_pad  ;
	output \702(2228)_pad  ;
	output \704(1281)_pad  ;
	output \707(1277)_pad  ;
	output \712(2297)_pad  ;
	output \715(1278)_pad  ;
	output \722(2131)_pad  ;
	output \727(2298)_pad  ;
	output \732(2300)_pad  ;
	output \737(2279)_pad  ;
	output \742(2238)_pad  ;
	output \747(2187)_pad  ;
	output \752(2189)_pad  ;
	output \757(2190)_pad  ;
	output \762(2184)_pad  ;
	output \767(2479)_pad  ;
	output \772(2299)_pad  ;
	output \777(2278)_pad  ;
	output \782(2239)_pad  ;
	output \787(2186)_pad  ;
	output \792(2188)_pad  ;
	output \797(2191)_pad  ;
	output \802(2183)_pad  ;
	output \807(2480)_pad  ;
	output \809(655)_pad  ;
	output \810(356)_pad  ;
	output \813(2260)_pad  ;
	output \815(627)_pad  ;
	output \820(1283)_pad  ;
	output \822(1933)_pad  ;
	output \824(2274)_pad  ;
	output \826(2275)_pad  ;
	output \828(2233)_pad  ;
	output \830(2182)_pad  ;
	output \832(2133)_pad  ;
	output \834(2123)_pad  ;
	output \836(2128)_pad  ;
	output \838(2064)_pad  ;
	output \843(2455)_pad  ;
	output \845(845)_pad  ;
	output \847(465)_pad  ;
	output \848(330)_pad  ;
	output \849(219)_pad  ;
	output \850(217)_pad  ;
	output \851(218)_pad  ;
	output \854(2268)_pad  ;
	output \859(2132)_pad  ;
	output \861(2070)_pad  ;
	output \863(2276)_pad  ;
	output \865(2277)_pad  ;
	output \867(2237)_pad  ;
	output \869(2181)_pad  ;
	output \871(2127)_pad  ;
	output \873(2124)_pad  ;
	output \875(2125)_pad  ;
	output \877(2126)_pad  ;
	output \882(2456)_pad  ;
	output \998(2163)_pad  ;
	output \u2023_syn_3  ;
	output \u2095_syn_3  ;
	output \u2109_syn_3  ;
	output \u2318_syn_3  ;
	output \u3086_syn_3  ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w422_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w417_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w237_ ;
	wire _w367_ ;
	wire _w110_ ;
	wire _w651_ ;
	wire _w236_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w363_ ;
	wire _w106_ ;
	wire _w647_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w219_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w191_ ;
	wire _w223_ ;
	wire _w421_ ;
	wire _w164_ ;
	wire _w705_ ;
	wire _w291_ ;
	wire _w224_ ;
	wire _w332_ ;
	wire _w75_ ;
	wire _w616_ ;
	wire _w202_ ;
	wire _w193_ ;
	wire _w220_ ;
	wire _w418_ ;
	wire _w161_ ;
	wire _w702_ ;
	wire _w288_ ;
	wire _w218_ ;
	wire _w416_ ;
	wire _w159_ ;
	wire _w700_ ;
	wire _w286_ ;
	wire _w238_ ;
	wire _w377_ ;
	wire _w120_ ;
	wire _w661_ ;
	wire _w247_ ;
	wire _w207_ ;
	wire _w182_ ;
	wire _w235_ ;
	wire _w374_ ;
	wire _w117_ ;
	wire _w658_ ;
	wire _w244_ ;
	wire _w204_ ;
	wire _w228_ ;
	wire _w197_ ;
	wire _w184_ ;
	wire _w192_ ;
	wire _w225_ ;
	wire _w423_ ;
	wire _w166_ ;
	wire _w707_ ;
	wire _w293_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w196_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w203_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w208_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w287_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w292_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w701_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w706_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\245(98)_pad ,
		_w75_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\338(124)_pad ,
		_w106_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\348(126)_pad ,
		_w110_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\358(128)_pad ,
		_w117_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\366(130)_pad ,
		_w120_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\545(150)_pad ,
		_w159_
	);
	LUT1 #(
		.INIT('h1)
	) name6 (
		\552(152)_pad ,
		_w161_
	);
	LUT1 #(
		.INIT('h1)
	) name7 (
		\559(154)_pad ,
		_w164_
	);
	LUT1 #(
		.INIT('h1)
	) name8 (
		\562(155)_pad ,
		_w166_
	);
	LUT1 #(
		.INIT('h1)
	) name9 (
		\889(734)_pad ,
		_w182_
	);
	LUT1 #(
		.INIT('h1)
	) name10 (
		\892(408)_pad ,
		_w184_
	);
	LUT3 #(
		.INIT('h35)
	) name11 (
		\226(93)_pad ,
		\233(94)_pad ,
		\335(123)_pad ,
		_w191_
	);
	LUT3 #(
		.INIT('h35)
	) name12 (
		\257(102)_pad ,
		\264(103)_pad ,
		\335(123)_pad ,
		_w192_
	);
	LUT3 #(
		.INIT('h35)
	) name13 (
		\273(106)_pad ,
		\280(107)_pad ,
		\335(123)_pad ,
		_w193_
	);
	LUT3 #(
		.INIT('h69)
	) name14 (
		_w191_,
		_w192_,
		_w193_,
		_w194_
	);
	LUT3 #(
		.INIT('h35)
	) name15 (
		\234(95)_pad ,
		\241(96)_pad ,
		\335(123)_pad ,
		_w195_
	);
	LUT3 #(
		.INIT('h35)
	) name16 (
		\281(108)_pad ,
		\288(109)_pad ,
		\335(123)_pad ,
		_w196_
	);
	LUT2 #(
		.INIT('h9)
	) name17 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT3 #(
		.INIT('h35)
	) name18 (
		\265(104)_pad ,
		\272(105)_pad ,
		\335(123)_pad ,
		_w198_
	);
	LUT3 #(
		.INIT('h35)
	) name19 (
		\210(89)_pad ,
		\217(90)_pad ,
		\335(123)_pad ,
		_w199_
	);
	LUT3 #(
		.INIT('hca)
	) name20 (
		\289(110)_pad ,
		\292(111)_pad ,
		\335(123)_pad ,
		_w200_
	);
	LUT3 #(
		.INIT('h69)
	) name21 (
		_w198_,
		_w199_,
		_w200_,
		_w201_
	);
	LUT3 #(
		.INIT('h35)
	) name22 (
		\218(91)_pad ,
		\225(92)_pad ,
		\335(123)_pad ,
		_w202_
	);
	LUT3 #(
		.INIT('h35)
	) name23 (
		\206(87)_pad ,
		\209(88)_pad ,
		\335(123)_pad ,
		_w203_
	);
	LUT2 #(
		.INIT('h9)
	) name24 (
		_w202_,
		_w203_,
		_w204_
	);
	LUT4 #(
		.INIT('h9669)
	) name25 (
		_w194_,
		_w197_,
		_w201_,
		_w204_,
		_w205_
	);
	LUT4 #(
		.INIT('h6996)
	) name26 (
		\316(118)_pad ,
		\324(120)_pad ,
		\341(125)_pad ,
		\369(131)_pad ,
		_w206_
	);
	LUT3 #(
		.INIT('h96)
	) name27 (
		\298(299)_pad ,
		\308(116)_pad ,
		\361(129)_pad ,
		_w207_
	);
	LUT2 #(
		.INIT('h9)
	) name28 (
		\302(114)_pad ,
		\351(127)_pad ,
		_w208_
	);
	LUT3 #(
		.INIT('h69)
	) name29 (
		_w206_,
		_w207_,
		_w208_,
		_w209_
	);
	LUT3 #(
		.INIT('h96)
	) name30 (
		_w206_,
		_w207_,
		_w208_,
		_w210_
	);
	LUT4 #(
		.INIT('h6996)
	) name31 (
		\206(87)_pad ,
		\218(91)_pad ,
		\281(108)_pad ,
		\289(110)_pad ,
		_w211_
	);
	LUT4 #(
		.INIT('h9669)
	) name32 (
		\210(89)_pad ,
		\257(102)_pad ,
		\265(104)_pad ,
		\273(106)_pad ,
		_w212_
	);
	LUT2 #(
		.INIT('h9)
	) name33 (
		\226(93)_pad ,
		\234(95)_pad ,
		_w213_
	);
	LUT3 #(
		.INIT('h69)
	) name34 (
		_w211_,
		_w212_,
		_w213_,
		_w214_
	);
	LUT3 #(
		.INIT('h96)
	) name35 (
		_w211_,
		_w212_,
		_w213_,
		_w215_
	);
	LUT4 #(
		.INIT('hca00)
	) name36 (
		\281(108)_pad ,
		\288(109)_pad ,
		\335(123)_pad ,
		\374(134)_pad ,
		_w216_
	);
	LUT4 #(
		.INIT('h0035)
	) name37 (
		\281(108)_pad ,
		\288(109)_pad ,
		\335(123)_pad ,
		\374(134)_pad ,
		_w217_
	);
	LUT4 #(
		.INIT('h35ca)
	) name38 (
		\281(108)_pad ,
		\288(109)_pad ,
		\335(123)_pad ,
		\374(134)_pad ,
		_w218_
	);
	LUT4 #(
		.INIT('hca00)
	) name39 (
		\273(106)_pad ,
		\280(107)_pad ,
		\335(123)_pad ,
		\411(138)_pad ,
		_w219_
	);
	LUT4 #(
		.INIT('h0035)
	) name40 (
		\273(106)_pad ,
		\280(107)_pad ,
		\335(123)_pad ,
		\411(138)_pad ,
		_w220_
	);
	LUT4 #(
		.INIT('h35ca)
	) name41 (
		\273(106)_pad ,
		\280(107)_pad ,
		\335(123)_pad ,
		\411(138)_pad ,
		_w221_
	);
	LUT4 #(
		.INIT('hca00)
	) name42 (
		\265(104)_pad ,
		\272(105)_pad ,
		\335(123)_pad ,
		\400(137)_pad ,
		_w222_
	);
	LUT4 #(
		.INIT('h0035)
	) name43 (
		\265(104)_pad ,
		\272(105)_pad ,
		\335(123)_pad ,
		\400(137)_pad ,
		_w223_
	);
	LUT4 #(
		.INIT('h35ca)
	) name44 (
		\265(104)_pad ,
		\272(105)_pad ,
		\335(123)_pad ,
		\400(137)_pad ,
		_w224_
	);
	LUT3 #(
		.INIT('h80)
	) name45 (
		_w218_,
		_w221_,
		_w224_,
		_w225_
	);
	LUT4 #(
		.INIT('h35ca)
	) name46 (
		\234(95)_pad ,
		\241(96)_pad ,
		\335(123)_pad ,
		\435(140)_pad ,
		_w226_
	);
	LUT4 #(
		.INIT('hca00)
	) name47 (
		\257(102)_pad ,
		\264(103)_pad ,
		\335(123)_pad ,
		\389(136)_pad ,
		_w227_
	);
	LUT4 #(
		.INIT('h0035)
	) name48 (
		\257(102)_pad ,
		\264(103)_pad ,
		\335(123)_pad ,
		\389(136)_pad ,
		_w228_
	);
	LUT4 #(
		.INIT('h35ca)
	) name49 (
		\257(102)_pad ,
		\264(103)_pad ,
		\335(123)_pad ,
		\389(136)_pad ,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w226_,
		_w229_,
		_w230_
	);
	LUT4 #(
		.INIT('hca00)
	) name51 (
		\226(93)_pad ,
		\233(94)_pad ,
		\335(123)_pad ,
		\422(139)_pad ,
		_w231_
	);
	LUT4 #(
		.INIT('h35ca)
	) name52 (
		\218(91)_pad ,
		\225(92)_pad ,
		\335(123)_pad ,
		\468(143)_pad ,
		_w232_
	);
	LUT4 #(
		.INIT('h0035)
	) name53 (
		\226(93)_pad ,
		\233(94)_pad ,
		\335(123)_pad ,
		\422(139)_pad ,
		_w233_
	);
	LUT3 #(
		.INIT('h90)
	) name54 (
		\422(139)_pad ,
		_w191_,
		_w232_,
		_w234_
	);
	LUT4 #(
		.INIT('hca00)
	) name55 (
		\206(87)_pad ,
		\209(88)_pad ,
		\335(123)_pad ,
		\446(141)_pad ,
		_w235_
	);
	LUT4 #(
		.INIT('h0035)
	) name56 (
		\206(87)_pad ,
		\209(88)_pad ,
		\335(123)_pad ,
		\446(141)_pad ,
		_w236_
	);
	LUT4 #(
		.INIT('h35ca)
	) name57 (
		\206(87)_pad ,
		\209(88)_pad ,
		\335(123)_pad ,
		\446(141)_pad ,
		_w237_
	);
	LUT4 #(
		.INIT('hca00)
	) name58 (
		\210(89)_pad ,
		\217(90)_pad ,
		\335(123)_pad ,
		\457(142)_pad ,
		_w238_
	);
	LUT4 #(
		.INIT('h0035)
	) name59 (
		\210(89)_pad ,
		\217(90)_pad ,
		\335(123)_pad ,
		\457(142)_pad ,
		_w239_
	);
	LUT4 #(
		.INIT('h35ca)
	) name60 (
		\210(89)_pad ,
		\217(90)_pad ,
		\335(123)_pad ,
		\457(142)_pad ,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w237_,
		_w240_,
		_w241_
	);
	LUT4 #(
		.INIT('h8000)
	) name62 (
		_w234_,
		_w225_,
		_w230_,
		_w241_,
		_w242_
	);
	LUT4 #(
		.INIT('hac00)
	) name63 (
		\248(99)_pad ,
		\251(100)_pad ,
		\316(118)_pad ,
		\490(145)_pad ,
		_w243_
	);
	LUT4 #(
		.INIT('h0053)
	) name64 (
		\242(97)_pad ,
		\254(101)_pad ,
		\316(118)_pad ,
		\490(145)_pad ,
		_w244_
	);
	LUT4 #(
		.INIT('hac00)
	) name65 (
		\248(99)_pad ,
		\251(100)_pad ,
		\308(116)_pad ,
		\479(144)_pad ,
		_w245_
	);
	LUT4 #(
		.INIT('h0053)
	) name66 (
		\242(97)_pad ,
		\254(101)_pad ,
		\308(116)_pad ,
		\479(144)_pad ,
		_w246_
	);
	LUT4 #(
		.INIT('heee0)
	) name67 (
		_w243_,
		_w244_,
		_w245_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h1b00)
	) name68 (
		\341(125)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\523(148)_pad ,
		_w248_
	);
	LUT4 #(
		.INIT('h00d8)
	) name69 (
		\341(125)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\523(148)_pad ,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w248_,
		_w249_,
		_w250_
	);
	LUT3 #(
		.INIT('h53)
	) name71 (
		\242(97)_pad ,
		\254(101)_pad ,
		\298(299)_pad ,
		_w251_
	);
	LUT3 #(
		.INIT('h53)
	) name72 (
		\248(99)_pad ,
		\251(100)_pad ,
		\302(114)_pad ,
		_w252_
	);
	LUT3 #(
		.INIT('h53)
	) name73 (
		\248(99)_pad ,
		\251(100)_pad ,
		\361(129)_pad ,
		_w253_
	);
	LUT3 #(
		.INIT('hc5)
	) name74 (
		\3546(165)_pad ,
		\3552(168)_pad ,
		\514(147)_pad ,
		_w254_
	);
	LUT4 #(
		.INIT('h0004)
	) name75 (
		_w253_,
		_w251_,
		_w252_,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('h1b00)
	) name76 (
		\324(120)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\503(146)_pad ,
		_w256_
	);
	LUT4 #(
		.INIT('h00d8)
	) name77 (
		\324(120)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\503(146)_pad ,
		_w257_
	);
	LUT4 #(
		.INIT('h1b00)
	) name78 (
		\351(127)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\534(149)_pad ,
		_w258_
	);
	LUT4 #(
		.INIT('h00d8)
	) name79 (
		\351(127)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\534(149)_pad ,
		_w259_
	);
	LUT4 #(
		.INIT('heee0)
	) name80 (
		_w256_,
		_w257_,
		_w258_,
		_w259_,
		_w260_
	);
	LUT4 #(
		.INIT('h2000)
	) name81 (
		_w247_,
		_w250_,
		_w255_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\552(152)_pad ,
		\562(155)_pad ,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\332(122)_pad ,
		\338(124)_pad ,
		_w263_
	);
	LUT3 #(
		.INIT('h2d)
	) name84 (
		\332(122)_pad ,
		\338(124)_pad ,
		\514(147)_pad ,
		_w264_
	);
	LUT3 #(
		.INIT('h1b)
	) name85 (
		\332(122)_pad ,
		\341(125)_pad ,
		\348(126)_pad ,
		_w265_
	);
	LUT4 #(
		.INIT('he400)
	) name86 (
		\332(122)_pad ,
		\341(125)_pad ,
		\348(126)_pad ,
		\523(148)_pad ,
		_w266_
	);
	LUT4 #(
		.INIT('h001b)
	) name87 (
		\332(122)_pad ,
		\341(125)_pad ,
		\348(126)_pad ,
		\523(148)_pad ,
		_w267_
	);
	LUT4 #(
		.INIT('h1be4)
	) name88 (
		\332(122)_pad ,
		\341(125)_pad ,
		\348(126)_pad ,
		\523(148)_pad ,
		_w268_
	);
	LUT3 #(
		.INIT('h1b)
	) name89 (
		\332(122)_pad ,
		\351(127)_pad ,
		\358(128)_pad ,
		_w269_
	);
	LUT4 #(
		.INIT('he400)
	) name90 (
		\332(122)_pad ,
		\351(127)_pad ,
		\358(128)_pad ,
		\534(149)_pad ,
		_w270_
	);
	LUT4 #(
		.INIT('h001b)
	) name91 (
		\332(122)_pad ,
		\351(127)_pad ,
		\358(128)_pad ,
		\534(149)_pad ,
		_w271_
	);
	LUT4 #(
		.INIT('h1be4)
	) name92 (
		\332(122)_pad ,
		\351(127)_pad ,
		\358(128)_pad ,
		\534(149)_pad ,
		_w272_
	);
	LUT3 #(
		.INIT('h1b)
	) name93 (
		\332(122)_pad ,
		\361(129)_pad ,
		\366(130)_pad ,
		_w273_
	);
	LUT4 #(
		.INIT('h8000)
	) name94 (
		_w264_,
		_w268_,
		_w272_,
		_w273_,
		_w274_
	);
	LUT3 #(
		.INIT('hca)
	) name95 (
		\324(120)_pad ,
		\331(121)_pad ,
		\332(122)_pad ,
		_w275_
	);
	LUT4 #(
		.INIT('h35ca)
	) name96 (
		\324(120)_pad ,
		\331(121)_pad ,
		\332(122)_pad ,
		\503(146)_pad ,
		_w276_
	);
	LUT3 #(
		.INIT('h1d)
	) name97 (
		\298(299)_pad ,
		\332(122)_pad ,
		\889(734)_pad ,
		_w277_
	);
	LUT3 #(
		.INIT('h35)
	) name98 (
		\302(114)_pad ,
		\307(115)_pad ,
		\332(122)_pad ,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT3 #(
		.INIT('h35)
	) name100 (
		\308(116)_pad ,
		\315(117)_pad ,
		\332(122)_pad ,
		_w280_
	);
	LUT4 #(
		.INIT('h35ca)
	) name101 (
		\308(116)_pad ,
		\315(117)_pad ,
		\332(122)_pad ,
		\479(144)_pad ,
		_w281_
	);
	LUT3 #(
		.INIT('h35)
	) name102 (
		\316(118)_pad ,
		\323(119)_pad ,
		\332(122)_pad ,
		_w282_
	);
	LUT4 #(
		.INIT('hca00)
	) name103 (
		\316(118)_pad ,
		\323(119)_pad ,
		\332(122)_pad ,
		\490(145)_pad ,
		_w283_
	);
	LUT4 #(
		.INIT('h0035)
	) name104 (
		\316(118)_pad ,
		\323(119)_pad ,
		\332(122)_pad ,
		\490(145)_pad ,
		_w284_
	);
	LUT4 #(
		.INIT('h35ca)
	) name105 (
		\316(118)_pad ,
		\323(119)_pad ,
		\332(122)_pad ,
		\490(145)_pad ,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w281_,
		_w285_,
		_w286_
	);
	LUT4 #(
		.INIT('h8000)
	) name107 (
		_w277_,
		_w278_,
		_w281_,
		_w285_,
		_w287_
	);
	LUT3 #(
		.INIT('h80)
	) name108 (
		_w274_,
		_w276_,
		_w287_,
		_w288_
	);
	LUT4 #(
		.INIT('h3110)
	) name109 (
		\534(149)_pad ,
		_w266_,
		_w269_,
		_w273_,
		_w289_
	);
	LUT4 #(
		.INIT('h222b)
	) name110 (
		\514(147)_pad ,
		_w263_,
		_w267_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('he080)
	) name111 (
		\503(146)_pad ,
		_w275_,
		_w287_,
		_w290_,
		_w291_
	);
	LUT3 #(
		.INIT('h4d)
	) name112 (
		\479(144)_pad ,
		_w280_,
		_w283_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w279_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('hb)
	) name114 (
		_w291_,
		_w293_,
		_w294_
	);
	LUT3 #(
		.INIT('h4d)
	) name115 (
		\468(143)_pad ,
		_w202_,
		_w231_,
		_w295_
	);
	LUT4 #(
		.INIT('h004d)
	) name116 (
		\468(143)_pad ,
		_w202_,
		_w231_,
		_w238_,
		_w296_
	);
	LUT4 #(
		.INIT('h004d)
	) name117 (
		\411(138)_pad ,
		_w193_,
		_w216_,
		_w222_,
		_w297_
	);
	LUT4 #(
		.INIT('hddd4)
	) name118 (
		\389(136)_pad ,
		_w192_,
		_w223_,
		_w297_,
		_w298_
	);
	LUT4 #(
		.INIT('h20b0)
	) name119 (
		\435(140)_pad ,
		_w195_,
		_w234_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w236_,
		_w239_,
		_w300_
	);
	LUT4 #(
		.INIT('hfbaa)
	) name121 (
		_w235_,
		_w296_,
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\373(133)_pad ,
		\993(850)_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		\2358(162)_pad ,
		\87(33)_pad ,
		_w303_
	);
	LUT2 #(
		.INIT('h7)
	) name124 (
		\27(10)_pad ,
		\31(11)_pad ,
		_w304_
	);
	LUT4 #(
		.INIT('hc080)
	) name125 (
		\2358(162)_pad ,
		\27(10)_pad ,
		\31(11)_pad ,
		\86(32)_pad ,
		_w305_
	);
	LUT2 #(
		.INIT('hb)
	) name126 (
		_w303_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\2358(162)_pad ,
		\25(8)_pad ,
		_w307_
	);
	LUT4 #(
		.INIT('hb000)
	) name128 (
		\2358(162)_pad ,
		\24(7)_pad ,
		\27(10)_pad ,
		\31(11)_pad ,
		_w308_
	);
	LUT3 #(
		.INIT('h8a)
	) name129 (
		\144(354)_pad ,
		_w307_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w311_
	);
	LUT4 #(
		.INIT('h8000)
	) name132 (
		\54(20)_pad ,
		_w268_,
		_w272_,
		_w273_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w264_,
		_w312_,
		_w313_
	);
	LUT3 #(
		.INIT('h56)
	) name134 (
		_w276_,
		_w290_,
		_w313_,
		_w314_
	);
	LUT4 #(
		.INIT('h5060)
	) name135 (
		_w276_,
		_w290_,
		_w311_,
		_w313_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w316_
	);
	LUT3 #(
		.INIT('h40)
	) name137 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		\52(18)_pad ,
		_w317_
	);
	LUT4 #(
		.INIT('h00ef)
	) name138 (
		_w256_,
		_w257_,
		_w316_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w315_,
		_w318_,
		_w319_
	);
	LUT3 #(
		.INIT('h8a)
	) name140 (
		_w310_,
		_w315_,
		_w318_,
		_w320_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w321_
	);
	LUT4 #(
		.INIT('h8000)
	) name142 (
		\4(1)_pad ,
		_w218_,
		_w221_,
		_w224_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w229_,
		_w322_,
		_w323_
	);
	LUT3 #(
		.INIT('ha6)
	) name144 (
		_w226_,
		_w298_,
		_w323_,
		_w324_
	);
	LUT4 #(
		.INIT('h5090)
	) name145 (
		_w226_,
		_w298_,
		_w311_,
		_w323_,
		_w325_
	);
	LUT4 #(
		.INIT('h1b00)
	) name146 (
		\234(95)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\435(140)_pad ,
		_w326_
	);
	LUT4 #(
		.INIT('h00d8)
	) name147 (
		\234(95)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\435(140)_pad ,
		_w327_
	);
	LUT3 #(
		.INIT('h20)
	) name148 (
		\122(52)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w328_
	);
	LUT4 #(
		.INIT('h00fd)
	) name149 (
		_w316_,
		_w326_,
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w325_,
		_w329_,
		_w330_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name151 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		\170(75)_pad ,
		\200(85)_pad ,
		_w331_
	);
	LUT4 #(
		.INIT('h7500)
	) name152 (
		_w321_,
		_w325_,
		_w329_,
		_w331_,
		_w332_
	);
	LUT3 #(
		.INIT('h8a)
	) name153 (
		\926(624)_pad ,
		_w320_,
		_w332_,
		_w333_
	);
	LUT4 #(
		.INIT('h1117)
	) name154 (
		\503(146)_pad ,
		_w275_,
		_w290_,
		_w313_,
		_w334_
	);
	LUT3 #(
		.INIT('h20)
	) name155 (
		\112(42)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w335_
	);
	LUT4 #(
		.INIT('h00ef)
	) name156 (
		_w243_,
		_w244_,
		_w316_,
		_w335_,
		_w336_
	);
	LUT4 #(
		.INIT('h7b00)
	) name157 (
		_w285_,
		_w311_,
		_w334_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		_w310_,
		_w337_,
		_w338_
	);
	LUT4 #(
		.INIT('h35ca)
	) name159 (
		\226(93)_pad ,
		\233(94)_pad ,
		\335(123)_pad ,
		\422(139)_pad ,
		_w339_
	);
	LUT4 #(
		.INIT('hbb2b)
	) name160 (
		\435(140)_pad ,
		_w195_,
		_w298_,
		_w323_,
		_w340_
	);
	LUT4 #(
		.INIT('h1b00)
	) name161 (
		\226(93)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\422(139)_pad ,
		_w341_
	);
	LUT4 #(
		.INIT('h00d8)
	) name162 (
		\226(93)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\422(139)_pad ,
		_w342_
	);
	LUT3 #(
		.INIT('h20)
	) name163 (
		\113(43)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w343_
	);
	LUT4 #(
		.INIT('h00fd)
	) name164 (
		_w316_,
		_w341_,
		_w342_,
		_w343_,
		_w344_
	);
	LUT4 #(
		.INIT('hd700)
	) name165 (
		_w311_,
		_w339_,
		_w340_,
		_w344_,
		_w345_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name166 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		\173(76)_pad ,
		\203(86)_pad ,
		_w346_
	);
	LUT3 #(
		.INIT('hd0)
	) name167 (
		_w321_,
		_w345_,
		_w346_,
		_w347_
	);
	LUT3 #(
		.INIT('h8a)
	) name168 (
		\926(624)_pad ,
		_w338_,
		_w347_,
		_w348_
	);
	LUT3 #(
		.INIT('h40)
	) name169 (
		_w281_,
		_w285_,
		_w334_,
		_w349_
	);
	LUT2 #(
		.INIT('h9)
	) name170 (
		_w281_,
		_w284_,
		_w350_
	);
	LUT4 #(
		.INIT('hcc80)
	) name171 (
		_w285_,
		_w311_,
		_w334_,
		_w350_,
		_w351_
	);
	LUT3 #(
		.INIT('h20)
	) name172 (
		\116(46)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w352_
	);
	LUT4 #(
		.INIT('h00ef)
	) name173 (
		_w245_,
		_w246_,
		_w316_,
		_w352_,
		_w353_
	);
	LUT3 #(
		.INIT('hb0)
	) name174 (
		_w349_,
		_w351_,
		_w353_,
		_w354_
	);
	LUT4 #(
		.INIT('h20aa)
	) name175 (
		_w310_,
		_w349_,
		_w351_,
		_w353_,
		_w355_
	);
	LUT2 #(
		.INIT('h9)
	) name176 (
		_w232_,
		_w233_,
		_w356_
	);
	LUT4 #(
		.INIT('ha208)
	) name177 (
		_w311_,
		_w339_,
		_w340_,
		_w356_,
		_w357_
	);
	LUT4 #(
		.INIT('h1b00)
	) name178 (
		\218(91)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\468(143)_pad ,
		_w358_
	);
	LUT4 #(
		.INIT('h00d8)
	) name179 (
		\218(91)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\468(143)_pad ,
		_w359_
	);
	LUT3 #(
		.INIT('h40)
	) name180 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		\53(19)_pad ,
		_w360_
	);
	LUT4 #(
		.INIT('h00fd)
	) name181 (
		_w316_,
		_w358_,
		_w359_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w357_,
		_w361_,
		_w362_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name183 (
		\167(74)_pad ,
		\1689(157)_pad ,
		\1690(158)_pad ,
		\197(84)_pad ,
		_w363_
	);
	LUT4 #(
		.INIT('h7500)
	) name184 (
		_w321_,
		_w357_,
		_w361_,
		_w363_,
		_w364_
	);
	LUT3 #(
		.INIT('h8a)
	) name185 (
		\926(624)_pad ,
		_w355_,
		_w364_,
		_w365_
	);
	LUT3 #(
		.INIT('hc4)
	) name186 (
		_w286_,
		_w292_,
		_w334_,
		_w366_
	);
	LUT4 #(
		.INIT('ha020)
	) name187 (
		_w278_,
		_w286_,
		_w292_,
		_w334_,
		_w367_
	);
	LUT4 #(
		.INIT('h5a9a)
	) name188 (
		_w278_,
		_w286_,
		_w292_,
		_w334_,
		_w368_
	);
	LUT3 #(
		.INIT('h20)
	) name189 (
		\121(51)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w369_
	);
	LUT3 #(
		.INIT('h07)
	) name190 (
		_w252_,
		_w316_,
		_w369_,
		_w370_
	);
	LUT3 #(
		.INIT('hd0)
	) name191 (
		_w311_,
		_w368_,
		_w370_,
		_w371_
	);
	LUT4 #(
		.INIT('h08cc)
	) name192 (
		_w311_,
		_w310_,
		_w368_,
		_w370_,
		_w372_
	);
	LUT3 #(
		.INIT('hd4)
	) name193 (
		\468(143)_pad ,
		_w202_,
		_w233_,
		_w373_
	);
	LUT4 #(
		.INIT('haa59)
	) name194 (
		_w240_,
		_w295_,
		_w340_,
		_w373_,
		_w374_
	);
	LUT4 #(
		.INIT('h1b00)
	) name195 (
		\210(89)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\457(142)_pad ,
		_w375_
	);
	LUT4 #(
		.INIT('h00d8)
	) name196 (
		\210(89)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\457(142)_pad ,
		_w376_
	);
	LUT3 #(
		.INIT('h20)
	) name197 (
		\114(44)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w377_
	);
	LUT4 #(
		.INIT('h00fd)
	) name198 (
		_w316_,
		_w375_,
		_w376_,
		_w377_,
		_w378_
	);
	LUT3 #(
		.INIT('h70)
	) name199 (
		_w311_,
		_w374_,
		_w378_,
		_w379_
	);
	LUT4 #(
		.INIT('h80aa)
	) name200 (
		_w321_,
		_w311_,
		_w374_,
		_w378_,
		_w380_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name201 (
		\164(73)_pad ,
		\1689(157)_pad ,
		\1690(158)_pad ,
		\194(83)_pad ,
		_w381_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name202 (
		\926(624)_pad ,
		_w380_,
		_w372_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h6)
	) name203 (
		_w277_,
		_w367_,
		_w383_
	);
	LUT3 #(
		.INIT('h20)
	) name204 (
		\123(53)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w384_
	);
	LUT3 #(
		.INIT('h0b)
	) name205 (
		_w251_,
		_w316_,
		_w384_,
		_w385_
	);
	LUT4 #(
		.INIT('h7b00)
	) name206 (
		_w277_,
		_w311_,
		_w367_,
		_w385_,
		_w386_
	);
	LUT3 #(
		.INIT('h23)
	) name207 (
		_w234_,
		_w239_,
		_w296_,
		_w387_
	);
	LUT4 #(
		.INIT('h59aa)
	) name208 (
		_w237_,
		_w296_,
		_w340_,
		_w387_,
		_w388_
	);
	LUT4 #(
		.INIT('hd800)
	) name209 (
		\206(87)_pad ,
		\248(99)_pad ,
		\251(100)_pad ,
		\446(141)_pad ,
		_w389_
	);
	LUT4 #(
		.INIT('h0027)
	) name210 (
		\206(87)_pad ,
		\242(97)_pad ,
		\254(101)_pad ,
		\446(141)_pad ,
		_w390_
	);
	LUT3 #(
		.INIT('h20)
	) name211 (
		\115(45)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w391_
	);
	LUT4 #(
		.INIT('h00fd)
	) name212 (
		_w316_,
		_w389_,
		_w390_,
		_w391_,
		_w392_
	);
	LUT3 #(
		.INIT('h70)
	) name213 (
		_w311_,
		_w388_,
		_w392_,
		_w393_
	);
	LUT4 #(
		.INIT('h80aa)
	) name214 (
		_w321_,
		_w311_,
		_w388_,
		_w392_,
		_w394_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name215 (
		\161(72)_pad ,
		\1689(157)_pad ,
		\1690(158)_pad ,
		\191(82)_pad ,
		_w395_
	);
	LUT4 #(
		.INIT('h3100)
	) name216 (
		_w310_,
		_w394_,
		_w386_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h2)
	) name217 (
		\926(624)_pad ,
		_w396_,
		_w397_
	);
	LUT3 #(
		.INIT('h7f)
	) name218 (
		\140(64)_pad ,
		\27(10)_pad ,
		\31(11)_pad ,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\4092(176)_pad ,
		\97(37)_pad ,
		_w399_
	);
	LUT2 #(
		.INIT('h6)
	) name220 (
		_w226_,
		_w229_,
		_w400_
	);
	LUT3 #(
		.INIT('h42)
	) name221 (
		\411(138)_pad ,
		_w193_,
		_w216_,
		_w401_
	);
	LUT4 #(
		.INIT('h2224)
	) name222 (
		\389(136)_pad ,
		_w192_,
		_w223_,
		_w297_,
		_w402_
	);
	LUT2 #(
		.INIT('h9)
	) name223 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT4 #(
		.INIT('h0c0d)
	) name224 (
		_w223_,
		_w225_,
		_w228_,
		_w297_,
		_w404_
	);
	LUT4 #(
		.INIT('h0302)
	) name225 (
		_w223_,
		_w225_,
		_w227_,
		_w297_,
		_w405_
	);
	LUT3 #(
		.INIT('h24)
	) name226 (
		\411(138)_pad ,
		_w193_,
		_w217_,
		_w406_
	);
	LUT4 #(
		.INIT('h02a8)
	) name227 (
		_w218_,
		_w404_,
		_w405_,
		_w406_,
		_w407_
	);
	LUT4 #(
		.INIT('h41e9)
	) name228 (
		\1497(156)_pad ,
		_w218_,
		_w403_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h6)
	) name229 (
		_w221_,
		_w224_,
		_w409_
	);
	LUT3 #(
		.INIT('h80)
	) name230 (
		\1497(156)_pad ,
		_w225_,
		_w230_,
		_w410_
	);
	LUT4 #(
		.INIT('h00d4)
	) name231 (
		\435(140)_pad ,
		_w195_,
		_w298_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('hb4d2)
	) name232 (
		\457(142)_pad ,
		_w199_,
		_w237_,
		_w295_,
		_w412_
	);
	LUT2 #(
		.INIT('h6)
	) name233 (
		_w356_,
		_w412_,
		_w413_
	);
	LUT4 #(
		.INIT('h6996)
	) name234 (
		_w231_,
		_w232_,
		_w237_,
		_w240_,
		_w414_
	);
	LUT4 #(
		.INIT('h00dc)
	) name235 (
		_w234_,
		_w239_,
		_w296_,
		_w373_,
		_w415_
	);
	LUT4 #(
		.INIT('h6f00)
	) name236 (
		\422(139)_pad ,
		_w191_,
		_w232_,
		_w238_,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w295_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w415_,
		_w417_,
		_w418_
	);
	LUT4 #(
		.INIT('hd88d)
	) name239 (
		_w411_,
		_w413_,
		_w414_,
		_w418_,
		_w419_
	);
	LUT4 #(
		.INIT('h9669)
	) name240 (
		_w400_,
		_w408_,
		_w409_,
		_w419_,
		_w420_
	);
	LUT4 #(
		.INIT('hd800)
	) name241 (
		\234(95)_pad ,
		\248(99)_pad ,
		\251(100)_pad ,
		\435(140)_pad ,
		_w421_
	);
	LUT4 #(
		.INIT('h0027)
	) name242 (
		\234(95)_pad ,
		\242(97)_pad ,
		\254(101)_pad ,
		\435(140)_pad ,
		_w422_
	);
	LUT4 #(
		.INIT('hd800)
	) name243 (
		\226(93)_pad ,
		\248(99)_pad ,
		\251(100)_pad ,
		\422(139)_pad ,
		_w423_
	);
	LUT4 #(
		.INIT('h0027)
	) name244 (
		\226(93)_pad ,
		\242(97)_pad ,
		\254(101)_pad ,
		\422(139)_pad ,
		_w424_
	);
	LUT4 #(
		.INIT('heee1)
	) name245 (
		_w421_,
		_w422_,
		_w423_,
		_w424_,
		_w425_
	);
	LUT4 #(
		.INIT('hd800)
	) name246 (
		\210(89)_pad ,
		\248(99)_pad ,
		\251(100)_pad ,
		\457(142)_pad ,
		_w426_
	);
	LUT4 #(
		.INIT('h0027)
	) name247 (
		\210(89)_pad ,
		\242(97)_pad ,
		\254(101)_pad ,
		\457(142)_pad ,
		_w427_
	);
	LUT4 #(
		.INIT('heee1)
	) name248 (
		_w389_,
		_w390_,
		_w426_,
		_w427_,
		_w428_
	);
	LUT4 #(
		.INIT('hd800)
	) name249 (
		\218(91)_pad ,
		\248(99)_pad ,
		\251(100)_pad ,
		\468(143)_pad ,
		_w429_
	);
	LUT4 #(
		.INIT('h0027)
	) name250 (
		\218(91)_pad ,
		\242(97)_pad ,
		\254(101)_pad ,
		\468(143)_pad ,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w429_,
		_w430_,
		_w431_
	);
	LUT3 #(
		.INIT('h69)
	) name252 (
		_w425_,
		_w428_,
		_w431_,
		_w432_
	);
	LUT4 #(
		.INIT('hac00)
	) name253 (
		\248(99)_pad ,
		\251(100)_pad ,
		\257(102)_pad ,
		\389(136)_pad ,
		_w433_
	);
	LUT4 #(
		.INIT('h0053)
	) name254 (
		\242(97)_pad ,
		\254(101)_pad ,
		\257(102)_pad ,
		\389(136)_pad ,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w433_,
		_w434_,
		_w435_
	);
	LUT4 #(
		.INIT('hac00)
	) name256 (
		\248(99)_pad ,
		\251(100)_pad ,
		\281(108)_pad ,
		\374(134)_pad ,
		_w436_
	);
	LUT4 #(
		.INIT('h0053)
	) name257 (
		\242(97)_pad ,
		\254(101)_pad ,
		\281(108)_pad ,
		\374(134)_pad ,
		_w437_
	);
	LUT4 #(
		.INIT('hac00)
	) name258 (
		\248(99)_pad ,
		\251(100)_pad ,
		\273(106)_pad ,
		\411(138)_pad ,
		_w438_
	);
	LUT4 #(
		.INIT('h0053)
	) name259 (
		\242(97)_pad ,
		\254(101)_pad ,
		\273(106)_pad ,
		\411(138)_pad ,
		_w439_
	);
	LUT4 #(
		.INIT('heee1)
	) name260 (
		_w436_,
		_w437_,
		_w438_,
		_w439_,
		_w440_
	);
	LUT4 #(
		.INIT('hac00)
	) name261 (
		\248(99)_pad ,
		\251(100)_pad ,
		\265(104)_pad ,
		\400(137)_pad ,
		_w441_
	);
	LUT4 #(
		.INIT('h0053)
	) name262 (
		\242(97)_pad ,
		\254(101)_pad ,
		\265(104)_pad ,
		\400(137)_pad ,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w441_,
		_w442_,
		_w443_
	);
	LUT3 #(
		.INIT('h69)
	) name264 (
		_w435_,
		_w440_,
		_w443_,
		_w444_
	);
	LUT4 #(
		.INIT('h2332)
	) name265 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w432_,
		_w444_,
		_w445_
	);
	LUT4 #(
		.INIT('h2033)
	) name266 (
		\4091(175)_pad ,
		_w399_,
		_w420_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\4092(176)_pad ,
		\94(36)_pad ,
		_w447_
	);
	LUT4 #(
		.INIT('h9669)
	) name268 (
		_w264_,
		_w268_,
		_w272_,
		_w276_,
		_w448_
	);
	LUT3 #(
		.INIT('h24)
	) name269 (
		\523(148)_pad ,
		_w265_,
		_w271_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w274_,
		_w449_,
		_w450_
	);
	LUT4 #(
		.INIT('h0415)
	) name271 (
		_w273_,
		_w290_,
		_w449_,
		_w450_,
		_w451_
	);
	LUT4 #(
		.INIT('ha280)
	) name272 (
		_w273_,
		_w290_,
		_w449_,
		_w450_,
		_w452_
	);
	LUT4 #(
		.INIT('h2224)
	) name273 (
		\514(147)_pad ,
		_w263_,
		_w267_,
		_w289_,
		_w453_
	);
	LUT3 #(
		.INIT('h48)
	) name274 (
		_w270_,
		_w273_,
		_w453_,
		_w454_
	);
	LUT4 #(
		.INIT('h5746)
	) name275 (
		\2174(161)_pad ,
		_w451_,
		_w452_,
		_w454_,
		_w455_
	);
	LUT3 #(
		.INIT('h80)
	) name276 (
		\2174(161)_pad ,
		_w274_,
		_w276_,
		_w456_
	);
	LUT4 #(
		.INIT('h0017)
	) name277 (
		\503(146)_pad ,
		_w275_,
		_w290_,
		_w456_,
		_w457_
	);
	LUT4 #(
		.INIT('h2302)
	) name278 (
		\479(144)_pad ,
		_w278_,
		_w280_,
		_w283_,
		_w458_
	);
	LUT3 #(
		.INIT('h96)
	) name279 (
		_w277_,
		_w350_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h6)
	) name280 (
		_w281_,
		_w283_,
		_w460_
	);
	LUT4 #(
		.INIT('h0223)
	) name281 (
		\479(144)_pad ,
		_w278_,
		_w280_,
		_w284_,
		_w461_
	);
	LUT3 #(
		.INIT('h69)
	) name282 (
		_w277_,
		_w460_,
		_w461_,
		_w462_
	);
	LUT3 #(
		.INIT('hd8)
	) name283 (
		_w457_,
		_w459_,
		_w462_,
		_w463_
	);
	LUT4 #(
		.INIT('h2882)
	) name284 (
		\4091(175)_pad ,
		_w448_,
		_w455_,
		_w463_,
		_w464_
	);
	LUT3 #(
		.INIT('hc5)
	) name285 (
		\242(97)_pad ,
		\248(99)_pad ,
		\514(147)_pad ,
		_w465_
	);
	LUT2 #(
		.INIT('h9)
	) name286 (
		_w251_,
		_w252_,
		_w466_
	);
	LUT4 #(
		.INIT('h111e)
	) name287 (
		_w243_,
		_w244_,
		_w245_,
		_w246_,
		_w467_
	);
	LUT3 #(
		.INIT('h69)
	) name288 (
		_w465_,
		_w466_,
		_w467_,
		_w468_
	);
	LUT4 #(
		.INIT('hac00)
	) name289 (
		\248(99)_pad ,
		\251(100)_pad ,
		\324(120)_pad ,
		\503(146)_pad ,
		_w469_
	);
	LUT4 #(
		.INIT('h0053)
	) name290 (
		\242(97)_pad ,
		\254(101)_pad ,
		\324(120)_pad ,
		\503(146)_pad ,
		_w470_
	);
	LUT3 #(
		.INIT('h56)
	) name291 (
		_w253_,
		_w469_,
		_w470_,
		_w471_
	);
	LUT4 #(
		.INIT('hac00)
	) name292 (
		\248(99)_pad ,
		\251(100)_pad ,
		\341(125)_pad ,
		\523(148)_pad ,
		_w472_
	);
	LUT4 #(
		.INIT('h0053)
	) name293 (
		\242(97)_pad ,
		\254(101)_pad ,
		\341(125)_pad ,
		\523(148)_pad ,
		_w473_
	);
	LUT4 #(
		.INIT('hac00)
	) name294 (
		\248(99)_pad ,
		\251(100)_pad ,
		\351(127)_pad ,
		\534(149)_pad ,
		_w474_
	);
	LUT4 #(
		.INIT('h0053)
	) name295 (
		\242(97)_pad ,
		\254(101)_pad ,
		\351(127)_pad ,
		\534(149)_pad ,
		_w475_
	);
	LUT4 #(
		.INIT('heee1)
	) name296 (
		_w472_,
		_w473_,
		_w474_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h6)
	) name297 (
		_w471_,
		_w476_,
		_w477_
	);
	LUT4 #(
		.INIT('h3223)
	) name298 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w468_,
		_w477_,
		_w478_
	);
	LUT4 #(
		.INIT('h8a88)
	) name299 (
		_w310_,
		_w447_,
		_w464_,
		_w478_,
		_w479_
	);
	LUT4 #(
		.INIT('h37bf)
	) name300 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		\176(77)_pad ,
		\179(78)_pad ,
		_w480_
	);
	LUT4 #(
		.INIT('h0d00)
	) name301 (
		_w321_,
		_w446_,
		_w479_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('hd)
	) name302 (
		\926(624)_pad ,
		_w481_,
		_w482_
	);
	LUT3 #(
		.INIT('h60)
	) name303 (
		\4(1)_pad ,
		_w218_,
		_w311_,
		_w483_
	);
	LUT4 #(
		.INIT('h1b00)
	) name304 (
		\281(108)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\374(134)_pad ,
		_w484_
	);
	LUT4 #(
		.INIT('h00d8)
	) name305 (
		\281(108)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\374(134)_pad ,
		_w485_
	);
	LUT3 #(
		.INIT('h20)
	) name306 (
		\117(47)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w486_
	);
	LUT4 #(
		.INIT('h00fd)
	) name307 (
		_w316_,
		_w484_,
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		_w483_,
		_w487_,
		_w488_
	);
	LUT3 #(
		.INIT('h8a)
	) name309 (
		_w321_,
		_w483_,
		_w487_,
		_w489_
	);
	LUT4 #(
		.INIT('h001b)
	) name310 (
		\332(122)_pad ,
		\361(129)_pad ,
		\366(130)_pad ,
		\54(20)_pad ,
		_w490_
	);
	LUT4 #(
		.INIT('h1be4)
	) name311 (
		\332(122)_pad ,
		\361(129)_pad ,
		\366(130)_pad ,
		\54(20)_pad ,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		_w311_,
		_w491_,
		_w492_
	);
	LUT3 #(
		.INIT('h20)
	) name313 (
		\131(59)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w493_
	);
	LUT3 #(
		.INIT('h07)
	) name314 (
		_w253_,
		_w316_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w492_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('h37bf)
	) name316 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		\182(79)_pad ,
		\185(80)_pad ,
		_w496_
	);
	LUT4 #(
		.INIT('h7500)
	) name317 (
		_w310_,
		_w492_,
		_w494_,
		_w496_,
		_w497_
	);
	LUT3 #(
		.INIT('h8a)
	) name318 (
		\926(624)_pad ,
		_w489_,
		_w497_,
		_w498_
	);
	LUT4 #(
		.INIT('h718e)
	) name319 (
		\374(134)_pad ,
		\4(1)_pad ,
		_w196_,
		_w221_,
		_w499_
	);
	LUT4 #(
		.INIT('h1b00)
	) name320 (
		\273(106)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\411(138)_pad ,
		_w500_
	);
	LUT4 #(
		.INIT('h00d8)
	) name321 (
		\273(106)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\411(138)_pad ,
		_w501_
	);
	LUT3 #(
		.INIT('h20)
	) name322 (
		\126(54)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w502_
	);
	LUT4 #(
		.INIT('h00fd)
	) name323 (
		_w316_,
		_w500_,
		_w501_,
		_w502_,
		_w503_
	);
	LUT3 #(
		.INIT('h70)
	) name324 (
		_w311_,
		_w499_,
		_w503_,
		_w504_
	);
	LUT4 #(
		.INIT('h80aa)
	) name325 (
		_w321_,
		_w311_,
		_w499_,
		_w503_,
		_w505_
	);
	LUT4 #(
		.INIT('h9060)
	) name326 (
		\534(149)_pad ,
		_w269_,
		_w311_,
		_w490_,
		_w506_
	);
	LUT3 #(
		.INIT('h20)
	) name327 (
		\129(57)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w507_
	);
	LUT4 #(
		.INIT('h00ef)
	) name328 (
		_w258_,
		_w259_,
		_w316_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w506_,
		_w508_,
		_w509_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name330 (
		\158(71)_pad ,
		\1689(157)_pad ,
		\1690(158)_pad ,
		\188(81)_pad ,
		_w510_
	);
	LUT4 #(
		.INIT('h7500)
	) name331 (
		_w310_,
		_w506_,
		_w508_,
		_w510_,
		_w511_
	);
	LUT3 #(
		.INIT('h8a)
	) name332 (
		\926(624)_pad ,
		_w505_,
		_w511_,
		_w512_
	);
	LUT4 #(
		.INIT('h008e)
	) name333 (
		\374(134)_pad ,
		\4(1)_pad ,
		_w196_,
		_w220_,
		_w513_
	);
	LUT3 #(
		.INIT('h36)
	) name334 (
		_w219_,
		_w224_,
		_w513_,
		_w514_
	);
	LUT4 #(
		.INIT('h3060)
	) name335 (
		_w219_,
		_w224_,
		_w311_,
		_w513_,
		_w515_
	);
	LUT4 #(
		.INIT('h1b00)
	) name336 (
		\265(104)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\400(137)_pad ,
		_w516_
	);
	LUT4 #(
		.INIT('h00d8)
	) name337 (
		\265(104)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\400(137)_pad ,
		_w517_
	);
	LUT3 #(
		.INIT('h20)
	) name338 (
		\127(55)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w518_
	);
	LUT4 #(
		.INIT('h00fd)
	) name339 (
		_w316_,
		_w516_,
		_w517_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		_w515_,
		_w519_,
		_w520_
	);
	LUT3 #(
		.INIT('h8a)
	) name341 (
		_w321_,
		_w515_,
		_w519_,
		_w521_
	);
	LUT4 #(
		.INIT('h399c)
	) name342 (
		\534(149)_pad ,
		_w268_,
		_w269_,
		_w490_,
		_w522_
	);
	LUT3 #(
		.INIT('h20)
	) name343 (
		\119(49)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w523_
	);
	LUT4 #(
		.INIT('h00ef)
	) name344 (
		_w248_,
		_w249_,
		_w316_,
		_w523_,
		_w524_
	);
	LUT3 #(
		.INIT('hd0)
	) name345 (
		_w311_,
		_w522_,
		_w524_,
		_w525_
	);
	LUT4 #(
		.INIT('h08cc)
	) name346 (
		_w311_,
		_w310_,
		_w522_,
		_w524_,
		_w526_
	);
	LUT4 #(
		.INIT('h53ff)
	) name347 (
		\152(69)_pad ,
		\155(70)_pad ,
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		_w526_,
		_w527_,
		_w528_
	);
	LUT3 #(
		.INIT('h8a)
	) name349 (
		\926(624)_pad ,
		_w521_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('hcc36)
	) name350 (
		_w223_,
		_w229_,
		_w297_,
		_w322_,
		_w530_
	);
	LUT4 #(
		.INIT('h1b00)
	) name351 (
		\257(102)_pad ,
		\3550(167)_pad ,
		\3552(168)_pad ,
		\389(136)_pad ,
		_w531_
	);
	LUT4 #(
		.INIT('h00d8)
	) name352 (
		\257(102)_pad ,
		\3546(165)_pad ,
		\3548(166)_pad ,
		\389(136)_pad ,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w531_,
		_w532_,
		_w533_
	);
	LUT3 #(
		.INIT('h20)
	) name354 (
		\128(56)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w534_
	);
	LUT4 #(
		.INIT('h00fd)
	) name355 (
		_w316_,
		_w531_,
		_w532_,
		_w534_,
		_w535_
	);
	LUT3 #(
		.INIT('hd0)
	) name356 (
		_w311_,
		_w530_,
		_w535_,
		_w536_
	);
	LUT4 #(
		.INIT('h08aa)
	) name357 (
		_w321_,
		_w311_,
		_w530_,
		_w535_,
		_w537_
	);
	LUT4 #(
		.INIT('haa56)
	) name358 (
		_w264_,
		_w267_,
		_w289_,
		_w312_,
		_w538_
	);
	LUT3 #(
		.INIT('h20)
	) name359 (
		\130(58)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w539_
	);
	LUT3 #(
		.INIT('h07)
	) name360 (
		_w254_,
		_w316_,
		_w539_,
		_w540_
	);
	LUT3 #(
		.INIT('hd0)
	) name361 (
		_w311_,
		_w538_,
		_w540_,
		_w541_
	);
	LUT4 #(
		.INIT('h08cc)
	) name362 (
		_w311_,
		_w310_,
		_w538_,
		_w540_,
		_w542_
	);
	LUT4 #(
		.INIT('h53ff)
	) name363 (
		\146(67)_pad ,
		\149(68)_pad ,
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w543_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name364 (
		\926(624)_pad ,
		_w542_,
		_w537_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\2358(162)_pad ,
		\81(29)_pad ,
		_w545_
	);
	LUT4 #(
		.INIT('hb000)
	) name366 (
		\2358(162)_pad ,
		\26(9)_pad ,
		\27(10)_pad ,
		\31(11)_pad ,
		_w546_
	);
	LUT3 #(
		.INIT('h8a)
	) name367 (
		\144(354)_pad ,
		_w545_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w548_
	);
	LUT3 #(
		.INIT('hb0)
	) name369 (
		_w315_,
		_w318_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w550_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name371 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		\170(75)_pad ,
		\200(85)_pad ,
		_w551_
	);
	LUT4 #(
		.INIT('h4f00)
	) name372 (
		_w325_,
		_w329_,
		_w550_,
		_w551_,
		_w552_
	);
	LUT3 #(
		.INIT('h8a)
	) name373 (
		\926(624)_pad ,
		_w549_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w337_,
		_w548_,
		_w554_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name375 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		\173(76)_pad ,
		\203(86)_pad ,
		_w555_
	);
	LUT3 #(
		.INIT('hb0)
	) name376 (
		_w345_,
		_w550_,
		_w555_,
		_w556_
	);
	LUT3 #(
		.INIT('h8a)
	) name377 (
		\926(624)_pad ,
		_w554_,
		_w556_,
		_w557_
	);
	LUT4 #(
		.INIT('h4f00)
	) name378 (
		_w349_,
		_w351_,
		_w353_,
		_w548_,
		_w558_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name379 (
		\167(74)_pad ,
		\1691(159)_pad ,
		\1694(160)_pad ,
		\197(84)_pad ,
		_w559_
	);
	LUT4 #(
		.INIT('h4f00)
	) name380 (
		_w357_,
		_w361_,
		_w550_,
		_w559_,
		_w560_
	);
	LUT3 #(
		.INIT('h8a)
	) name381 (
		\926(624)_pad ,
		_w558_,
		_w560_,
		_w561_
	);
	LUT4 #(
		.INIT('h2f00)
	) name382 (
		_w311_,
		_w368_,
		_w370_,
		_w548_,
		_w562_
	);
	LUT4 #(
		.INIT('h8f00)
	) name383 (
		_w311_,
		_w374_,
		_w378_,
		_w550_,
		_w563_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name384 (
		\164(73)_pad ,
		\1691(159)_pad ,
		\1694(160)_pad ,
		\194(83)_pad ,
		_w564_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name385 (
		\926(624)_pad ,
		_w563_,
		_w562_,
		_w564_,
		_w565_
	);
	LUT4 #(
		.INIT('h8f00)
	) name386 (
		_w311_,
		_w388_,
		_w392_,
		_w550_,
		_w566_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name387 (
		\161(72)_pad ,
		\1691(159)_pad ,
		\1694(160)_pad ,
		\191(82)_pad ,
		_w567_
	);
	LUT4 #(
		.INIT('h0b00)
	) name388 (
		_w386_,
		_w548_,
		_w566_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		\926(624)_pad ,
		_w568_,
		_w569_
	);
	LUT4 #(
		.INIT('hba00)
	) name390 (
		_w447_,
		_w464_,
		_w478_,
		_w548_,
		_w570_
	);
	LUT4 #(
		.INIT('h37bf)
	) name391 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		\176(77)_pad ,
		\179(78)_pad ,
		_w571_
	);
	LUT4 #(
		.INIT('h0b00)
	) name392 (
		_w446_,
		_w550_,
		_w570_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('hd)
	) name393 (
		\926(624)_pad ,
		_w572_,
		_w573_
	);
	LUT3 #(
		.INIT('hb0)
	) name394 (
		_w483_,
		_w487_,
		_w550_,
		_w574_
	);
	LUT4 #(
		.INIT('h37bf)
	) name395 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		\182(79)_pad ,
		\185(80)_pad ,
		_w575_
	);
	LUT4 #(
		.INIT('h4f00)
	) name396 (
		_w492_,
		_w494_,
		_w548_,
		_w575_,
		_w576_
	);
	LUT3 #(
		.INIT('h8a)
	) name397 (
		\926(624)_pad ,
		_w574_,
		_w576_,
		_w577_
	);
	LUT4 #(
		.INIT('h8f00)
	) name398 (
		_w311_,
		_w499_,
		_w503_,
		_w550_,
		_w578_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name399 (
		\158(71)_pad ,
		\1691(159)_pad ,
		\1694(160)_pad ,
		\188(81)_pad ,
		_w579_
	);
	LUT4 #(
		.INIT('h4f00)
	) name400 (
		_w506_,
		_w508_,
		_w548_,
		_w579_,
		_w580_
	);
	LUT3 #(
		.INIT('h8a)
	) name401 (
		\926(624)_pad ,
		_w578_,
		_w580_,
		_w581_
	);
	LUT3 #(
		.INIT('hb0)
	) name402 (
		_w515_,
		_w519_,
		_w550_,
		_w582_
	);
	LUT4 #(
		.INIT('h2f00)
	) name403 (
		_w311_,
		_w522_,
		_w524_,
		_w548_,
		_w583_
	);
	LUT4 #(
		.INIT('h53ff)
	) name404 (
		\152(69)_pad ,
		\155(70)_pad ,
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w584_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT3 #(
		.INIT('h8a)
	) name406 (
		\926(624)_pad ,
		_w582_,
		_w585_,
		_w586_
	);
	LUT4 #(
		.INIT('h2f00)
	) name407 (
		_w311_,
		_w530_,
		_w535_,
		_w550_,
		_w587_
	);
	LUT4 #(
		.INIT('h2f00)
	) name408 (
		_w311_,
		_w538_,
		_w540_,
		_w548_,
		_w588_
	);
	LUT4 #(
		.INIT('h53ff)
	) name409 (
		\146(67)_pad ,
		\149(68)_pad ,
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w589_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name410 (
		\926(624)_pad ,
		_w588_,
		_w587_,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		\2358(162)_pad ,
		\34(12)_pad ,
		_w591_
	);
	LUT4 #(
		.INIT('hc080)
	) name412 (
		\2358(162)_pad ,
		\27(10)_pad ,
		\31(11)_pad ,
		\88(34)_pad ,
		_w592_
	);
	LUT2 #(
		.INIT('hb)
	) name413 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\23(6)_pad ,
		\2358(162)_pad ,
		_w594_
	);
	LUT4 #(
		.INIT('h80c0)
	) name415 (
		\2358(162)_pad ,
		\27(10)_pad ,
		\31(11)_pad ,
		\79(27)_pad ,
		_w595_
	);
	LUT3 #(
		.INIT('h8a)
	) name416 (
		\144(354)_pad ,
		_w594_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w597_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w598_
	);
	LUT4 #(
		.INIT('h8f00)
	) name419 (
		_w311_,
		_w388_,
		_w392_,
		_w598_,
		_w599_
	);
	LUT4 #(
		.INIT('h53ff)
	) name420 (
		\106(40)_pad ,
		\109(41)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w600_
	);
	LUT4 #(
		.INIT('hdcff)
	) name421 (
		_w386_,
		_w599_,
		_w597_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\2358(162)_pad ,
		\80(28)_pad ,
		_w602_
	);
	LUT4 #(
		.INIT('h80c0)
	) name423 (
		\2358(162)_pad ,
		\27(10)_pad ,
		\31(11)_pad ,
		\82(30)_pad ,
		_w603_
	);
	LUT3 #(
		.INIT('h8a)
	) name424 (
		\144(354)_pad ,
		_w602_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w605_
	);
	LUT3 #(
		.INIT('hb0)
	) name426 (
		_w483_,
		_w487_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w607_
	);
	LUT4 #(
		.INIT('h37f7)
	) name428 (
		\11(2)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		\61(21)_pad ,
		_w608_
	);
	LUT4 #(
		.INIT('h4f00)
	) name429 (
		_w492_,
		_w494_,
		_w607_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('hb)
	) name430 (
		_w606_,
		_w609_,
		_w610_
	);
	LUT4 #(
		.INIT('h8f00)
	) name431 (
		_w311_,
		_w388_,
		_w392_,
		_w605_,
		_w611_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name432 (
		\106(40)_pad ,
		\109(41)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w612_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name433 (
		_w386_,
		_w607_,
		_w611_,
		_w612_,
		_w613_
	);
	LUT4 #(
		.INIT('h2f00)
	) name434 (
		_w311_,
		_w368_,
		_w370_,
		_w607_,
		_w614_
	);
	LUT4 #(
		.INIT('h8f00)
	) name435 (
		_w311_,
		_w374_,
		_w378_,
		_w605_,
		_w615_
	);
	LUT4 #(
		.INIT('h57df)
	) name436 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		\46(16)_pad ,
		\49(17)_pad ,
		_w616_
	);
	LUT3 #(
		.INIT('hef)
	) name437 (
		_w615_,
		_w614_,
		_w616_,
		_w617_
	);
	LUT4 #(
		.INIT('h4f00)
	) name438 (
		_w349_,
		_w351_,
		_w353_,
		_w607_,
		_w618_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name439 (
		\100(38)_pad ,
		\103(39)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w619_
	);
	LUT4 #(
		.INIT('h4f00)
	) name440 (
		_w357_,
		_w361_,
		_w605_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('hb)
	) name441 (
		_w618_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w337_,
		_w607_,
		_w622_
	);
	LUT4 #(
		.INIT('h737f)
	) name443 (
		\40(14)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		\91(35)_pad ,
		_w623_
	);
	LUT3 #(
		.INIT('hb0)
	) name444 (
		_w345_,
		_w605_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('hb)
	) name445 (
		_w622_,
		_w624_,
		_w625_
	);
	LUT3 #(
		.INIT('hb0)
	) name446 (
		_w315_,
		_w318_,
		_w607_,
		_w626_
	);
	LUT4 #(
		.INIT('h737f)
	) name447 (
		\37(13)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		\43(15)_pad ,
		_w627_
	);
	LUT4 #(
		.INIT('h4f00)
	) name448 (
		_w325_,
		_w329_,
		_w605_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('hb)
	) name449 (
		_w626_,
		_w628_,
		_w629_
	);
	LUT4 #(
		.INIT('h2f00)
	) name450 (
		_w311_,
		_w530_,
		_w535_,
		_w605_,
		_w630_
	);
	LUT4 #(
		.INIT('h2f00)
	) name451 (
		_w311_,
		_w538_,
		_w540_,
		_w607_,
		_w631_
	);
	LUT4 #(
		.INIT('h737f)
	) name452 (
		\20(5)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		\76(26)_pad ,
		_w632_
	);
	LUT3 #(
		.INIT('hef)
	) name453 (
		_w631_,
		_w630_,
		_w632_,
		_w633_
	);
	LUT3 #(
		.INIT('hb0)
	) name454 (
		_w515_,
		_w519_,
		_w605_,
		_w634_
	);
	LUT4 #(
		.INIT('h2f00)
	) name455 (
		_w311_,
		_w522_,
		_w524_,
		_w607_,
		_w635_
	);
	LUT4 #(
		.INIT('h737f)
	) name456 (
		\17(4)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		\73(25)_pad ,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('hb)
	) name458 (
		_w634_,
		_w637_,
		_w638_
	);
	LUT4 #(
		.INIT('h8f00)
	) name459 (
		_w311_,
		_w499_,
		_w503_,
		_w605_,
		_w639_
	);
	LUT4 #(
		.INIT('h57df)
	) name460 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		\67(23)_pad ,
		\70(24)_pad ,
		_w640_
	);
	LUT4 #(
		.INIT('h4f00)
	) name461 (
		_w506_,
		_w508_,
		_w607_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('hb)
	) name462 (
		_w639_,
		_w641_,
		_w642_
	);
	LUT4 #(
		.INIT('hba00)
	) name463 (
		_w447_,
		_w464_,
		_w478_,
		_w607_,
		_w643_
	);
	LUT4 #(
		.INIT('h37f7)
	) name464 (
		\14(3)_pad ,
		\4087(171)_pad ,
		\4088(172)_pad ,
		\64(22)_pad ,
		_w644_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name465 (
		_w446_,
		_w605_,
		_w643_,
		_w644_,
		_w645_
	);
	LUT4 #(
		.INIT('h2f00)
	) name466 (
		_w311_,
		_w368_,
		_w370_,
		_w597_,
		_w646_
	);
	LUT4 #(
		.INIT('h8f00)
	) name467 (
		_w311_,
		_w374_,
		_w378_,
		_w598_,
		_w647_
	);
	LUT4 #(
		.INIT('h37bf)
	) name468 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		\46(16)_pad ,
		\49(17)_pad ,
		_w648_
	);
	LUT3 #(
		.INIT('hef)
	) name469 (
		_w647_,
		_w646_,
		_w648_,
		_w649_
	);
	LUT4 #(
		.INIT('h4f00)
	) name470 (
		_w349_,
		_w351_,
		_w353_,
		_w597_,
		_w650_
	);
	LUT4 #(
		.INIT('h35ff)
	) name471 (
		\100(38)_pad ,
		\103(39)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w651_
	);
	LUT4 #(
		.INIT('h4f00)
	) name472 (
		_w357_,
		_w361_,
		_w598_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('hb)
	) name473 (
		_w650_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		_w337_,
		_w597_,
		_w654_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name475 (
		\40(14)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		\91(35)_pad ,
		_w655_
	);
	LUT3 #(
		.INIT('hb0)
	) name476 (
		_w345_,
		_w598_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('hb)
	) name477 (
		_w654_,
		_w656_,
		_w657_
	);
	LUT3 #(
		.INIT('hb0)
	) name478 (
		_w315_,
		_w318_,
		_w597_,
		_w658_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name479 (
		\37(13)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		\43(15)_pad ,
		_w659_
	);
	LUT4 #(
		.INIT('h4f00)
	) name480 (
		_w325_,
		_w329_,
		_w598_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('hb)
	) name481 (
		_w658_,
		_w660_,
		_w661_
	);
	LUT4 #(
		.INIT('h2f00)
	) name482 (
		_w311_,
		_w530_,
		_w535_,
		_w598_,
		_w662_
	);
	LUT4 #(
		.INIT('h2f00)
	) name483 (
		_w311_,
		_w538_,
		_w540_,
		_w597_,
		_w663_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name484 (
		\20(5)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		\76(26)_pad ,
		_w664_
	);
	LUT3 #(
		.INIT('hef)
	) name485 (
		_w663_,
		_w662_,
		_w664_,
		_w665_
	);
	LUT3 #(
		.INIT('hb0)
	) name486 (
		_w515_,
		_w519_,
		_w598_,
		_w666_
	);
	LUT4 #(
		.INIT('h2f00)
	) name487 (
		_w311_,
		_w522_,
		_w524_,
		_w597_,
		_w667_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name488 (
		\17(4)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		\73(25)_pad ,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('hb)
	) name490 (
		_w666_,
		_w669_,
		_w670_
	);
	LUT4 #(
		.INIT('h8f00)
	) name491 (
		_w311_,
		_w499_,
		_w503_,
		_w598_,
		_w671_
	);
	LUT4 #(
		.INIT('h37bf)
	) name492 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		\67(23)_pad ,
		\70(24)_pad ,
		_w672_
	);
	LUT4 #(
		.INIT('h4f00)
	) name493 (
		_w506_,
		_w508_,
		_w597_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('hb)
	) name494 (
		_w671_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('hba00)
	) name495 (
		_w447_,
		_w464_,
		_w478_,
		_w597_,
		_w675_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name496 (
		\14(3)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		\64(22)_pad ,
		_w676_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name497 (
		_w446_,
		_w598_,
		_w675_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\144(354)_pad ,
		\145(66)_pad ,
		_w678_
	);
	LUT2 #(
		.INIT('h9)
	) name499 (
		\132(60)_pad ,
		_w367_,
		_w679_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		\136(62)_pad ,
		\973(202)_pad ,
		_w680_
	);
	LUT3 #(
		.INIT('h7f)
	) name501 (
		\27(10)_pad ,
		\31(11)_pad ,
		\83(31)_pad ,
		_w681_
	);
	LUT4 #(
		.INIT('h2882)
	) name502 (
		_w311_,
		_w448_,
		_w455_,
		_w463_,
		_w682_
	);
	LUT4 #(
		.INIT('h8998)
	) name503 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w468_,
		_w477_,
		_w683_
	);
	LUT3 #(
		.INIT('h20)
	) name504 (
		\120(50)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w683_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('hb)
	) name506 (
		_w682_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('hd)
	) name507 (
		\27(10)_pad ,
		\2824(163)_pad ,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\386(135)_pad ,
		\556(153)_pad ,
		_w688_
	);
	LUT2 #(
		.INIT('h7)
	) name509 (
		\386(135)_pad ,
		\556(153)_pad ,
		_w689_
	);
	LUT3 #(
		.INIT('h1b)
	) name510 (
		\332(122)_pad ,
		\369(131)_pad ,
		\372(132)_pad ,
		_w690_
	);
	LUT4 #(
		.INIT('h9669)
	) name511 (
		_w265_,
		_w278_,
		_w280_,
		_w690_,
		_w691_
	);
	LUT4 #(
		.INIT('h9669)
	) name512 (
		_w269_,
		_w273_,
		_w277_,
		_w282_,
		_w692_
	);
	LUT4 #(
		.INIT('h35c5)
	) name513 (
		\324(120)_pad ,
		\331(121)_pad ,
		\332(122)_pad ,
		\338(124)_pad ,
		_w693_
	);
	LUT3 #(
		.INIT('h69)
	) name514 (
		_w691_,
		_w692_,
		_w693_,
		_w694_
	);
	LUT3 #(
		.INIT('h96)
	) name515 (
		_w691_,
		_w692_,
		_w693_,
		_w695_
	);
	LUT4 #(
		.INIT('h8000)
	) name516 (
		\245(98)_pad ,
		\552(152)_pad ,
		\559(154)_pad ,
		\562(155)_pad ,
		_w696_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		_w688_,
		_w696_,
		_w697_
	);
	LUT3 #(
		.INIT('h80)
	) name518 (
		_w209_,
		_w214_,
		_w697_,
		_w698_
	);
	LUT3 #(
		.INIT('h40)
	) name519 (
		_w205_,
		_w694_,
		_w698_,
		_w699_
	);
	LUT3 #(
		.INIT('hb0)
	) name520 (
		_w483_,
		_w487_,
		_w598_,
		_w700_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name521 (
		\11(2)_pad ,
		\4089(173)_pad ,
		\4090(174)_pad ,
		\61(21)_pad ,
		_w701_
	);
	LUT4 #(
		.INIT('h4f00)
	) name522 (
		_w492_,
		_w494_,
		_w597_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('hb)
	) name523 (
		_w700_,
		_w702_,
		_w703_
	);
	LUT4 #(
		.INIT('h9889)
	) name524 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w432_,
		_w444_,
		_w704_
	);
	LUT3 #(
		.INIT('h20)
	) name525 (
		\118(48)_pad ,
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w704_,
		_w705_,
		_w706_
	);
	LUT3 #(
		.INIT('h8f)
	) name527 (
		_w311_,
		_w420_,
		_w706_,
		_w707_
	);
	LUT3 #(
		.INIT('hc4)
	) name528 (
		\123(53)_pad ,
		\3717(169)_pad ,
		\3724(170)_pad ,
		_w708_
	);
	LUT4 #(
		.INIT('h7d00)
	) name529 (
		\3724(170)_pad ,
		_w277_,
		_w367_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h8)
	) name530 (
		\135(61)_pad ,
		\4115(177)_pad ,
		_w710_
	);
	LUT4 #(
		.INIT('h56a6)
	) name531 (
		\132(60)_pad ,
		\298(299)_pad ,
		\332(122)_pad ,
		\889(734)_pad ,
		_w711_
	);
	LUT4 #(
		.INIT('h5410)
	) name532 (
		\3717(169)_pad ,
		\3724(170)_pad ,
		_w251_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w710_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		_w709_,
		_w713_,
		_w714_
	);
	LUT4 #(
		.INIT('h2814)
	) name535 (
		\4(1)_pad ,
		_w232_,
		_w233_,
		_w218_,
		_w715_
	);
	LUT2 #(
		.INIT('h4)
	) name536 (
		_w499_,
		_w715_,
		_w716_
	);
	LUT3 #(
		.INIT('h40)
	) name537 (
		_w514_,
		_w530_,
		_w716_,
		_w717_
	);
	LUT4 #(
		.INIT('h8200)
	) name538 (
		_w324_,
		_w339_,
		_w340_,
		_w717_,
		_w718_
	);
	LUT3 #(
		.INIT('h10)
	) name539 (
		_w374_,
		_w388_,
		_w718_,
		_w719_
	);
	LUT4 #(
		.INIT('h2800)
	) name540 (
		_w272_,
		_w281_,
		_w284_,
		_w491_,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		_w522_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h8)
	) name542 (
		_w538_,
		_w721_,
		_w722_
	);
	LUT4 #(
		.INIT('h1200)
	) name543 (
		_w285_,
		_w314_,
		_w334_,
		_w722_,
		_w723_
	);
	LUT4 #(
		.INIT('h2800)
	) name544 (
		_w277_,
		_w278_,
		_w366_,
		_w723_,
		_w724_
	);
	LUT4 #(
		.INIT('heee0)
	) name545 (
		_w500_,
		_w501_,
		_w516_,
		_w517_,
		_w725_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w533_,
		_w725_,
		_w726_
	);
	LUT4 #(
		.INIT('heee0)
	) name547 (
		_w326_,
		_w327_,
		_w341_,
		_w342_,
		_w727_
	);
	LUT4 #(
		.INIT('heee0)
	) name548 (
		_w358_,
		_w359_,
		_w375_,
		_w376_,
		_w728_
	);
	LUT4 #(
		.INIT('heee0)
	) name549 (
		_w389_,
		_w390_,
		_w484_,
		_w485_,
		_w729_
	);
	LUT3 #(
		.INIT('h80)
	) name550 (
		_w727_,
		_w728_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		_w726_,
		_w730_,
		_w731_
	);
	assign \1000(2168)_pad  = _w205_ ;
	assign \1002(1920)_pad  = _w210_ ;
	assign \1004(1977)_pad  = _w215_ ;
	assign \588(1696)_pad  = _w242_ ;
	assign \593(733)_pad  = _w182_ ;
	assign \598(1623)_pad  = _w261_ ;
	assign \599(269)_pad  = _w110_ ;
	assign \600(259)_pad  = _w120_ ;
	assign \601(220)_pad  = _w262_ ;
	assign \604(223)_pad  = _w159_ ;
	assign \606(407)_pad  = _w184_ ;
	assign \611(275)_pad  = _w106_ ;
	assign \612(263)_pad  = _w117_ ;
	assign \615(1750)_pad  = _w288_ ;
	assign \618(1925)_pad  = _w294_ ;
	assign \621(1893)_pad  = _w301_ ;
	assign \626(1752)_pad  = _w288_ ;
	assign \632(1692)_pad  = _w242_ ;
	assign \634(665)_pad  = _w302_ ;
	assign \636(1280)_pad  = _w306_ ;
	assign \639(1275)_pad  = _w309_ ;
	assign \642(2222)_pad  = _w333_ ;
	assign \645(2271)_pad  = _w348_ ;
	assign \648(2295)_pad  = _w365_ ;
	assign \651(2314)_pad  = _w382_ ;
	assign \654(2315)_pad  = _w397_ ;
	assign \656(621)_pad  = _w398_ ;
	assign \658(2483)_pad  = _w482_ ;
	assign \661(2178)_pad  = _w498_ ;
	assign \664(2223)_pad  = _w512_ ;
	assign \667(2224)_pad  = _w529_ ;
	assign \670(2225)_pad  = _w544_ ;
	assign \673(1276)_pad  = _w547_ ;
	assign \676(2229)_pad  = _w553_ ;
	assign \679(2272)_pad  = _w557_ ;
	assign \682(2296)_pad  = _w561_ ;
	assign \685(2316)_pad  = _w565_ ;
	assign \688(2317)_pad  = _w569_ ;
	assign \690(2484)_pad  = _w573_ ;
	assign \693(2179)_pad  = _w577_ ;
	assign \696(2226)_pad  = _w581_ ;
	assign \699(2227)_pad  = _w586_ ;
	assign \702(2228)_pad  = _w590_ ;
	assign \704(1281)_pad  = _w593_ ;
	assign \707(1277)_pad  = _w596_ ;
	assign \712(2297)_pad  = _w601_ ;
	assign \715(1278)_pad  = _w604_ ;
	assign \722(2131)_pad  = _w610_ ;
	assign \727(2298)_pad  = _w613_ ;
	assign \732(2300)_pad  = _w617_ ;
	assign \737(2279)_pad  = _w621_ ;
	assign \742(2238)_pad  = _w625_ ;
	assign \747(2187)_pad  = _w629_ ;
	assign \752(2189)_pad  = _w633_ ;
	assign \757(2190)_pad  = _w638_ ;
	assign \762(2184)_pad  = _w642_ ;
	assign \767(2479)_pad  = _w645_ ;
	assign \772(2299)_pad  = _w649_ ;
	assign \777(2278)_pad  = _w653_ ;
	assign \782(2239)_pad  = _w657_ ;
	assign \787(2186)_pad  = _w661_ ;
	assign \792(2188)_pad  = _w665_ ;
	assign \797(2191)_pad  = _w670_ ;
	assign \802(2183)_pad  = _w674_ ;
	assign \807(2480)_pad  = _w677_ ;
	assign \809(655)_pad  = _w304_ ;
	assign \810(356)_pad  = _w678_ ;
	assign \813(2260)_pad  = _w679_ ;
	assign \815(627)_pad  = _w680_ ;
	assign \820(1283)_pad  = _w681_ ;
	assign \822(1933)_pad  = _w495_ ;
	assign \824(2274)_pad  = _w386_ ;
	assign \826(2275)_pad  = _w371_ ;
	assign \828(2233)_pad  = _w354_ ;
	assign \830(2182)_pad  = _w337_ ;
	assign \832(2133)_pad  = _w319_ ;
	assign \834(2123)_pad  = _w541_ ;
	assign \836(2128)_pad  = _w525_ ;
	assign \838(2064)_pad  = _w509_ ;
	assign \843(2455)_pad  = _w686_ ;
	assign \845(845)_pad  = _w687_ ;
	assign \847(465)_pad  = _w689_ ;
	assign \848(330)_pad  = _w75_ ;
	assign \849(219)_pad  = _w161_ ;
	assign \850(217)_pad  = _w166_ ;
	assign \851(218)_pad  = _w164_ ;
	assign \854(2268)_pad  = _w699_ ;
	assign \859(2132)_pad  = _w703_ ;
	assign \861(2070)_pad  = _w488_ ;
	assign \863(2276)_pad  = _w393_ ;
	assign \865(2277)_pad  = _w379_ ;
	assign \867(2237)_pad  = _w362_ ;
	assign \869(2181)_pad  = _w345_ ;
	assign \871(2127)_pad  = _w330_ ;
	assign \873(2124)_pad  = _w536_ ;
	assign \875(2125)_pad  = _w520_ ;
	assign \877(2126)_pad  = _w504_ ;
	assign \882(2456)_pad  = _w707_ ;
	assign \998(2163)_pad  = _w695_ ;
	assign \u2023_syn_3  = _w714_ ;
	assign \u2095_syn_3  = _w719_ ;
	assign \u2109_syn_3  = _w724_ ;
	assign \u2318_syn_3  = _w383_ ;
	assign \u3086_syn_3  = _w731_ ;
endmodule;